
module compare_N16384_CC8 ( clk, rst, x, y, g );
  input [2047:0] x;
  input [2047:0] y;
  input clk, rst;
  output g;
  wire   ci, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240;

  DFF ci_reg ( .D(g), .CLK(clk), .RST(rst), .I(1'b1), .Q(ci) );
  XOR U2052 ( .A(y[3]), .B(n10227), .Z(n10228) );
  XOR U2053 ( .A(y[7]), .B(n10211), .Z(n10212) );
  XOR U2054 ( .A(y[11]), .B(n10195), .Z(n10196) );
  XOR U2055 ( .A(y[15]), .B(n10179), .Z(n10180) );
  XOR U2056 ( .A(y[19]), .B(n10163), .Z(n10164) );
  XOR U2057 ( .A(y[23]), .B(n10147), .Z(n10148) );
  XOR U2058 ( .A(y[27]), .B(n10131), .Z(n10132) );
  XOR U2059 ( .A(y[31]), .B(n10115), .Z(n10116) );
  XOR U2060 ( .A(y[35]), .B(n10099), .Z(n10100) );
  XOR U2061 ( .A(y[39]), .B(n10083), .Z(n10084) );
  XOR U2062 ( .A(y[43]), .B(n10067), .Z(n10068) );
  XOR U2063 ( .A(y[47]), .B(n10051), .Z(n10052) );
  XOR U2064 ( .A(y[51]), .B(n10035), .Z(n10036) );
  XOR U2065 ( .A(y[55]), .B(n10019), .Z(n10020) );
  XOR U2066 ( .A(y[59]), .B(n10003), .Z(n10004) );
  XOR U2067 ( .A(y[63]), .B(n9987), .Z(n9988) );
  XOR U2068 ( .A(y[67]), .B(n9971), .Z(n9972) );
  XOR U2069 ( .A(y[71]), .B(n9955), .Z(n9956) );
  XOR U2070 ( .A(y[75]), .B(n9939), .Z(n9940) );
  XOR U2071 ( .A(y[79]), .B(n9923), .Z(n9924) );
  XOR U2072 ( .A(y[83]), .B(n9907), .Z(n9908) );
  XOR U2073 ( .A(y[87]), .B(n9891), .Z(n9892) );
  XOR U2074 ( .A(y[91]), .B(n9875), .Z(n9876) );
  XOR U2075 ( .A(y[95]), .B(n9859), .Z(n9860) );
  XOR U2076 ( .A(y[99]), .B(n9843), .Z(n9844) );
  XOR U2077 ( .A(y[103]), .B(n9827), .Z(n9828) );
  XOR U2078 ( .A(y[107]), .B(n9811), .Z(n9812) );
  XOR U2079 ( .A(y[111]), .B(n9795), .Z(n9796) );
  XOR U2080 ( .A(y[115]), .B(n9779), .Z(n9780) );
  XOR U2081 ( .A(y[119]), .B(n9763), .Z(n9764) );
  XOR U2082 ( .A(y[123]), .B(n9747), .Z(n9748) );
  XOR U2083 ( .A(y[127]), .B(n9731), .Z(n9732) );
  XOR U2084 ( .A(y[131]), .B(n9715), .Z(n9716) );
  XOR U2085 ( .A(y[135]), .B(n9699), .Z(n9700) );
  XOR U2086 ( .A(y[139]), .B(n9683), .Z(n9684) );
  XOR U2087 ( .A(y[143]), .B(n9667), .Z(n9668) );
  XOR U2088 ( .A(y[147]), .B(n9651), .Z(n9652) );
  XOR U2089 ( .A(y[151]), .B(n9635), .Z(n9636) );
  XOR U2090 ( .A(y[155]), .B(n9619), .Z(n9620) );
  XOR U2091 ( .A(y[159]), .B(n9603), .Z(n9604) );
  XOR U2092 ( .A(y[163]), .B(n9587), .Z(n9588) );
  XOR U2093 ( .A(y[167]), .B(n9571), .Z(n9572) );
  XOR U2094 ( .A(y[171]), .B(n9555), .Z(n9556) );
  XOR U2095 ( .A(y[175]), .B(n9539), .Z(n9540) );
  XOR U2096 ( .A(y[179]), .B(n9523), .Z(n9524) );
  XOR U2097 ( .A(y[183]), .B(n9507), .Z(n9508) );
  XOR U2098 ( .A(y[187]), .B(n9491), .Z(n9492) );
  XOR U2099 ( .A(y[191]), .B(n9475), .Z(n9476) );
  XOR U2100 ( .A(y[195]), .B(n9459), .Z(n9460) );
  XOR U2101 ( .A(y[199]), .B(n9443), .Z(n9444) );
  XOR U2102 ( .A(y[203]), .B(n9427), .Z(n9428) );
  XOR U2103 ( .A(y[207]), .B(n9411), .Z(n9412) );
  XOR U2104 ( .A(y[211]), .B(n9395), .Z(n9396) );
  XOR U2105 ( .A(y[215]), .B(n9379), .Z(n9380) );
  XOR U2106 ( .A(y[219]), .B(n9363), .Z(n9364) );
  XOR U2107 ( .A(y[223]), .B(n9347), .Z(n9348) );
  XOR U2108 ( .A(y[227]), .B(n9331), .Z(n9332) );
  XOR U2109 ( .A(y[231]), .B(n9315), .Z(n9316) );
  XOR U2110 ( .A(y[235]), .B(n9299), .Z(n9300) );
  XOR U2111 ( .A(y[239]), .B(n9283), .Z(n9284) );
  XOR U2112 ( .A(y[243]), .B(n9267), .Z(n9268) );
  XOR U2113 ( .A(y[247]), .B(n9251), .Z(n9252) );
  XOR U2114 ( .A(y[251]), .B(n9235), .Z(n9236) );
  XOR U2115 ( .A(y[255]), .B(n9219), .Z(n9220) );
  XOR U2116 ( .A(y[259]), .B(n9203), .Z(n9204) );
  XOR U2117 ( .A(y[263]), .B(n9187), .Z(n9188) );
  XOR U2118 ( .A(y[267]), .B(n9171), .Z(n9172) );
  XOR U2119 ( .A(y[271]), .B(n9155), .Z(n9156) );
  XOR U2120 ( .A(y[275]), .B(n9139), .Z(n9140) );
  XOR U2121 ( .A(y[279]), .B(n9123), .Z(n9124) );
  XOR U2122 ( .A(y[283]), .B(n9107), .Z(n9108) );
  XOR U2123 ( .A(y[287]), .B(n9091), .Z(n9092) );
  XOR U2124 ( .A(y[291]), .B(n9075), .Z(n9076) );
  XOR U2125 ( .A(y[295]), .B(n9059), .Z(n9060) );
  XOR U2126 ( .A(y[299]), .B(n9043), .Z(n9044) );
  XOR U2127 ( .A(y[303]), .B(n9027), .Z(n9028) );
  XOR U2128 ( .A(y[307]), .B(n9011), .Z(n9012) );
  XOR U2129 ( .A(y[311]), .B(n8995), .Z(n8996) );
  XOR U2130 ( .A(y[315]), .B(n8979), .Z(n8980) );
  XOR U2131 ( .A(y[319]), .B(n8963), .Z(n8964) );
  XOR U2132 ( .A(y[323]), .B(n8947), .Z(n8948) );
  XOR U2133 ( .A(y[327]), .B(n8931), .Z(n8932) );
  XOR U2134 ( .A(y[331]), .B(n8915), .Z(n8916) );
  XOR U2135 ( .A(y[335]), .B(n8899), .Z(n8900) );
  XOR U2136 ( .A(y[339]), .B(n8883), .Z(n8884) );
  XOR U2137 ( .A(y[343]), .B(n8867), .Z(n8868) );
  XOR U2138 ( .A(y[347]), .B(n8851), .Z(n8852) );
  XOR U2139 ( .A(y[351]), .B(n8835), .Z(n8836) );
  XOR U2140 ( .A(y[355]), .B(n8819), .Z(n8820) );
  XOR U2141 ( .A(y[359]), .B(n8803), .Z(n8804) );
  XOR U2142 ( .A(y[363]), .B(n8787), .Z(n8788) );
  XOR U2143 ( .A(y[367]), .B(n8771), .Z(n8772) );
  XOR U2144 ( .A(y[371]), .B(n8755), .Z(n8756) );
  XOR U2145 ( .A(y[375]), .B(n8739), .Z(n8740) );
  XOR U2146 ( .A(y[379]), .B(n8723), .Z(n8724) );
  XOR U2147 ( .A(y[383]), .B(n8707), .Z(n8708) );
  XOR U2148 ( .A(y[387]), .B(n8691), .Z(n8692) );
  XOR U2149 ( .A(y[391]), .B(n8675), .Z(n8676) );
  XOR U2150 ( .A(y[395]), .B(n8659), .Z(n8660) );
  XOR U2151 ( .A(y[399]), .B(n8643), .Z(n8644) );
  XOR U2152 ( .A(y[403]), .B(n8627), .Z(n8628) );
  XOR U2153 ( .A(y[407]), .B(n8611), .Z(n8612) );
  XOR U2154 ( .A(y[411]), .B(n8595), .Z(n8596) );
  XOR U2155 ( .A(y[415]), .B(n8579), .Z(n8580) );
  XOR U2156 ( .A(y[419]), .B(n8563), .Z(n8564) );
  XOR U2157 ( .A(y[423]), .B(n8547), .Z(n8548) );
  XOR U2158 ( .A(y[427]), .B(n8531), .Z(n8532) );
  XOR U2159 ( .A(y[431]), .B(n8515), .Z(n8516) );
  XOR U2160 ( .A(y[435]), .B(n8499), .Z(n8500) );
  XOR U2161 ( .A(y[439]), .B(n8483), .Z(n8484) );
  XOR U2162 ( .A(y[443]), .B(n8467), .Z(n8468) );
  XOR U2163 ( .A(y[447]), .B(n8451), .Z(n8452) );
  XOR U2164 ( .A(y[451]), .B(n8435), .Z(n8436) );
  XOR U2165 ( .A(y[455]), .B(n8419), .Z(n8420) );
  XOR U2166 ( .A(y[459]), .B(n8403), .Z(n8404) );
  XOR U2167 ( .A(y[463]), .B(n8387), .Z(n8388) );
  XOR U2168 ( .A(y[467]), .B(n8371), .Z(n8372) );
  XOR U2169 ( .A(y[471]), .B(n8355), .Z(n8356) );
  XOR U2170 ( .A(y[475]), .B(n8339), .Z(n8340) );
  XOR U2171 ( .A(y[479]), .B(n8323), .Z(n8324) );
  XOR U2172 ( .A(y[483]), .B(n8307), .Z(n8308) );
  XOR U2173 ( .A(y[487]), .B(n8291), .Z(n8292) );
  XOR U2174 ( .A(y[491]), .B(n8275), .Z(n8276) );
  XOR U2175 ( .A(y[495]), .B(n8259), .Z(n8260) );
  XOR U2176 ( .A(y[499]), .B(n8243), .Z(n8244) );
  XOR U2177 ( .A(y[503]), .B(n8227), .Z(n8228) );
  XOR U2178 ( .A(y[507]), .B(n8211), .Z(n8212) );
  XOR U2179 ( .A(y[511]), .B(n8195), .Z(n8196) );
  XOR U2180 ( .A(y[515]), .B(n8179), .Z(n8180) );
  XOR U2181 ( .A(y[519]), .B(n8163), .Z(n8164) );
  XOR U2182 ( .A(y[523]), .B(n8147), .Z(n8148) );
  XOR U2183 ( .A(y[527]), .B(n8131), .Z(n8132) );
  XOR U2184 ( .A(y[531]), .B(n8115), .Z(n8116) );
  XOR U2185 ( .A(y[535]), .B(n8099), .Z(n8100) );
  XOR U2186 ( .A(y[539]), .B(n8083), .Z(n8084) );
  XOR U2187 ( .A(y[543]), .B(n8067), .Z(n8068) );
  XOR U2188 ( .A(y[547]), .B(n8051), .Z(n8052) );
  XOR U2189 ( .A(y[551]), .B(n8035), .Z(n8036) );
  XOR U2190 ( .A(y[555]), .B(n8019), .Z(n8020) );
  XOR U2191 ( .A(y[559]), .B(n8003), .Z(n8004) );
  XOR U2192 ( .A(y[563]), .B(n7987), .Z(n7988) );
  XOR U2193 ( .A(y[567]), .B(n7971), .Z(n7972) );
  XOR U2194 ( .A(y[571]), .B(n7955), .Z(n7956) );
  XOR U2195 ( .A(y[575]), .B(n7939), .Z(n7940) );
  XOR U2196 ( .A(y[579]), .B(n7923), .Z(n7924) );
  XOR U2197 ( .A(y[583]), .B(n7907), .Z(n7908) );
  XOR U2198 ( .A(y[587]), .B(n7891), .Z(n7892) );
  XOR U2199 ( .A(y[591]), .B(n7875), .Z(n7876) );
  XOR U2200 ( .A(y[595]), .B(n7859), .Z(n7860) );
  XOR U2201 ( .A(y[599]), .B(n7843), .Z(n7844) );
  XOR U2202 ( .A(y[603]), .B(n7827), .Z(n7828) );
  XOR U2203 ( .A(y[607]), .B(n7811), .Z(n7812) );
  XOR U2204 ( .A(y[611]), .B(n7795), .Z(n7796) );
  XOR U2205 ( .A(y[615]), .B(n7779), .Z(n7780) );
  XOR U2206 ( .A(y[619]), .B(n7763), .Z(n7764) );
  XOR U2207 ( .A(y[623]), .B(n7747), .Z(n7748) );
  XOR U2208 ( .A(y[627]), .B(n7731), .Z(n7732) );
  XOR U2209 ( .A(y[631]), .B(n7715), .Z(n7716) );
  XOR U2210 ( .A(y[635]), .B(n7699), .Z(n7700) );
  XOR U2211 ( .A(y[639]), .B(n7683), .Z(n7684) );
  XOR U2212 ( .A(y[643]), .B(n7667), .Z(n7668) );
  XOR U2213 ( .A(y[647]), .B(n7651), .Z(n7652) );
  XOR U2214 ( .A(y[651]), .B(n7635), .Z(n7636) );
  XOR U2215 ( .A(y[655]), .B(n7619), .Z(n7620) );
  XOR U2216 ( .A(y[659]), .B(n7603), .Z(n7604) );
  XOR U2217 ( .A(y[663]), .B(n7587), .Z(n7588) );
  XOR U2218 ( .A(y[667]), .B(n7571), .Z(n7572) );
  XOR U2219 ( .A(y[671]), .B(n7555), .Z(n7556) );
  XOR U2220 ( .A(y[675]), .B(n7539), .Z(n7540) );
  XOR U2221 ( .A(y[679]), .B(n7523), .Z(n7524) );
  XOR U2222 ( .A(y[683]), .B(n7507), .Z(n7508) );
  XOR U2223 ( .A(y[687]), .B(n7491), .Z(n7492) );
  XOR U2224 ( .A(y[691]), .B(n7475), .Z(n7476) );
  XOR U2225 ( .A(y[695]), .B(n7459), .Z(n7460) );
  XOR U2226 ( .A(y[699]), .B(n7443), .Z(n7444) );
  XOR U2227 ( .A(y[703]), .B(n7427), .Z(n7428) );
  XOR U2228 ( .A(y[707]), .B(n7411), .Z(n7412) );
  XOR U2229 ( .A(y[711]), .B(n7395), .Z(n7396) );
  XOR U2230 ( .A(y[715]), .B(n7379), .Z(n7380) );
  XOR U2231 ( .A(y[719]), .B(n7363), .Z(n7364) );
  XOR U2232 ( .A(y[723]), .B(n7347), .Z(n7348) );
  XOR U2233 ( .A(y[727]), .B(n7331), .Z(n7332) );
  XOR U2234 ( .A(y[731]), .B(n7315), .Z(n7316) );
  XOR U2235 ( .A(y[735]), .B(n7299), .Z(n7300) );
  XOR U2236 ( .A(y[739]), .B(n7283), .Z(n7284) );
  XOR U2237 ( .A(y[743]), .B(n7267), .Z(n7268) );
  XOR U2238 ( .A(y[747]), .B(n7251), .Z(n7252) );
  XOR U2239 ( .A(y[751]), .B(n7235), .Z(n7236) );
  XOR U2240 ( .A(y[755]), .B(n7219), .Z(n7220) );
  XOR U2241 ( .A(y[759]), .B(n7203), .Z(n7204) );
  XOR U2242 ( .A(y[763]), .B(n7187), .Z(n7188) );
  XOR U2243 ( .A(y[767]), .B(n7171), .Z(n7172) );
  XOR U2244 ( .A(y[771]), .B(n7155), .Z(n7156) );
  XOR U2245 ( .A(y[775]), .B(n7139), .Z(n7140) );
  XOR U2246 ( .A(y[779]), .B(n7123), .Z(n7124) );
  XOR U2247 ( .A(y[783]), .B(n7107), .Z(n7108) );
  XOR U2248 ( .A(y[787]), .B(n7091), .Z(n7092) );
  XOR U2249 ( .A(y[791]), .B(n7075), .Z(n7076) );
  XOR U2250 ( .A(y[795]), .B(n7059), .Z(n7060) );
  XOR U2251 ( .A(y[799]), .B(n7043), .Z(n7044) );
  XOR U2252 ( .A(y[803]), .B(n7027), .Z(n7028) );
  XOR U2253 ( .A(y[807]), .B(n7011), .Z(n7012) );
  XOR U2254 ( .A(y[811]), .B(n6995), .Z(n6996) );
  XOR U2255 ( .A(y[815]), .B(n6979), .Z(n6980) );
  XOR U2256 ( .A(y[819]), .B(n6963), .Z(n6964) );
  XOR U2257 ( .A(y[823]), .B(n6947), .Z(n6948) );
  XOR U2258 ( .A(y[827]), .B(n6931), .Z(n6932) );
  XOR U2259 ( .A(y[831]), .B(n6915), .Z(n6916) );
  XOR U2260 ( .A(y[835]), .B(n6899), .Z(n6900) );
  XOR U2261 ( .A(y[839]), .B(n6883), .Z(n6884) );
  XOR U2262 ( .A(y[843]), .B(n6867), .Z(n6868) );
  XOR U2263 ( .A(y[847]), .B(n6851), .Z(n6852) );
  XOR U2264 ( .A(y[851]), .B(n6835), .Z(n6836) );
  XOR U2265 ( .A(y[855]), .B(n6819), .Z(n6820) );
  XOR U2266 ( .A(y[859]), .B(n6803), .Z(n6804) );
  XOR U2267 ( .A(y[863]), .B(n6787), .Z(n6788) );
  XOR U2268 ( .A(y[867]), .B(n6771), .Z(n6772) );
  XOR U2269 ( .A(y[871]), .B(n6755), .Z(n6756) );
  XOR U2270 ( .A(y[875]), .B(n6739), .Z(n6740) );
  XOR U2271 ( .A(y[879]), .B(n6723), .Z(n6724) );
  XOR U2272 ( .A(y[883]), .B(n6707), .Z(n6708) );
  XOR U2273 ( .A(y[887]), .B(n6691), .Z(n6692) );
  XOR U2274 ( .A(y[891]), .B(n6675), .Z(n6676) );
  XOR U2275 ( .A(y[895]), .B(n6659), .Z(n6660) );
  XOR U2276 ( .A(y[899]), .B(n6643), .Z(n6644) );
  XOR U2277 ( .A(y[903]), .B(n6627), .Z(n6628) );
  XOR U2278 ( .A(y[907]), .B(n6611), .Z(n6612) );
  XOR U2279 ( .A(y[911]), .B(n6595), .Z(n6596) );
  XOR U2280 ( .A(y[915]), .B(n6579), .Z(n6580) );
  XOR U2281 ( .A(y[919]), .B(n6563), .Z(n6564) );
  XOR U2282 ( .A(y[923]), .B(n6547), .Z(n6548) );
  XOR U2283 ( .A(y[927]), .B(n6531), .Z(n6532) );
  XOR U2284 ( .A(y[931]), .B(n6515), .Z(n6516) );
  XOR U2285 ( .A(y[935]), .B(n6499), .Z(n6500) );
  XOR U2286 ( .A(y[939]), .B(n6483), .Z(n6484) );
  XOR U2287 ( .A(y[943]), .B(n6467), .Z(n6468) );
  XOR U2288 ( .A(y[947]), .B(n6451), .Z(n6452) );
  XOR U2289 ( .A(y[951]), .B(n6435), .Z(n6436) );
  XOR U2290 ( .A(y[955]), .B(n6419), .Z(n6420) );
  XOR U2291 ( .A(y[959]), .B(n6403), .Z(n6404) );
  XOR U2292 ( .A(y[963]), .B(n6387), .Z(n6388) );
  XOR U2293 ( .A(y[967]), .B(n6371), .Z(n6372) );
  XOR U2294 ( .A(y[971]), .B(n6355), .Z(n6356) );
  XOR U2295 ( .A(y[975]), .B(n6339), .Z(n6340) );
  XOR U2296 ( .A(y[979]), .B(n6323), .Z(n6324) );
  XOR U2297 ( .A(y[983]), .B(n6307), .Z(n6308) );
  XOR U2298 ( .A(y[987]), .B(n6291), .Z(n6292) );
  XOR U2299 ( .A(y[991]), .B(n6275), .Z(n6276) );
  XOR U2300 ( .A(y[995]), .B(n6259), .Z(n6260) );
  XOR U2301 ( .A(y[999]), .B(n6243), .Z(n6244) );
  XOR U2302 ( .A(y[1003]), .B(n6227), .Z(n6228) );
  XOR U2303 ( .A(y[1007]), .B(n6211), .Z(n6212) );
  XOR U2304 ( .A(y[1011]), .B(n6195), .Z(n6196) );
  XOR U2305 ( .A(y[1015]), .B(n6179), .Z(n6180) );
  XOR U2306 ( .A(y[1019]), .B(n6163), .Z(n6164) );
  XOR U2307 ( .A(y[1023]), .B(n6147), .Z(n6148) );
  XOR U2308 ( .A(y[1027]), .B(n6131), .Z(n6132) );
  XOR U2309 ( .A(y[1031]), .B(n6115), .Z(n6116) );
  XOR U2310 ( .A(y[1035]), .B(n6099), .Z(n6100) );
  XOR U2311 ( .A(y[1039]), .B(n6083), .Z(n6084) );
  XOR U2312 ( .A(y[1043]), .B(n6067), .Z(n6068) );
  XOR U2313 ( .A(y[1047]), .B(n6051), .Z(n6052) );
  XOR U2314 ( .A(y[1051]), .B(n6035), .Z(n6036) );
  XOR U2315 ( .A(y[1055]), .B(n6019), .Z(n6020) );
  XOR U2316 ( .A(y[1059]), .B(n6003), .Z(n6004) );
  XOR U2317 ( .A(y[1063]), .B(n5987), .Z(n5988) );
  XOR U2318 ( .A(y[1067]), .B(n5971), .Z(n5972) );
  XOR U2319 ( .A(y[1071]), .B(n5955), .Z(n5956) );
  XOR U2320 ( .A(y[1075]), .B(n5939), .Z(n5940) );
  XOR U2321 ( .A(y[1079]), .B(n5923), .Z(n5924) );
  XOR U2322 ( .A(y[1083]), .B(n5907), .Z(n5908) );
  XOR U2323 ( .A(y[1087]), .B(n5891), .Z(n5892) );
  XOR U2324 ( .A(y[1091]), .B(n5875), .Z(n5876) );
  XOR U2325 ( .A(y[1095]), .B(n5859), .Z(n5860) );
  XOR U2326 ( .A(y[1099]), .B(n5843), .Z(n5844) );
  XOR U2327 ( .A(y[1103]), .B(n5827), .Z(n5828) );
  XOR U2328 ( .A(y[1107]), .B(n5811), .Z(n5812) );
  XOR U2329 ( .A(y[1111]), .B(n5795), .Z(n5796) );
  XOR U2330 ( .A(y[1115]), .B(n5779), .Z(n5780) );
  XOR U2331 ( .A(y[1119]), .B(n5763), .Z(n5764) );
  XOR U2332 ( .A(y[1123]), .B(n5747), .Z(n5748) );
  XOR U2333 ( .A(y[1127]), .B(n5731), .Z(n5732) );
  XOR U2334 ( .A(y[1131]), .B(n5715), .Z(n5716) );
  XOR U2335 ( .A(y[1135]), .B(n5699), .Z(n5700) );
  XOR U2336 ( .A(y[1139]), .B(n5683), .Z(n5684) );
  XOR U2337 ( .A(y[1143]), .B(n5667), .Z(n5668) );
  XOR U2338 ( .A(y[1147]), .B(n5651), .Z(n5652) );
  XOR U2339 ( .A(y[1151]), .B(n5635), .Z(n5636) );
  XOR U2340 ( .A(y[1155]), .B(n5619), .Z(n5620) );
  XOR U2341 ( .A(y[1159]), .B(n5603), .Z(n5604) );
  XOR U2342 ( .A(y[1163]), .B(n5587), .Z(n5588) );
  XOR U2343 ( .A(y[1167]), .B(n5571), .Z(n5572) );
  XOR U2344 ( .A(y[1171]), .B(n5555), .Z(n5556) );
  XOR U2345 ( .A(y[1175]), .B(n5539), .Z(n5540) );
  XOR U2346 ( .A(y[1179]), .B(n5523), .Z(n5524) );
  XOR U2347 ( .A(y[1183]), .B(n5507), .Z(n5508) );
  XOR U2348 ( .A(y[1187]), .B(n5491), .Z(n5492) );
  XOR U2349 ( .A(y[1191]), .B(n5475), .Z(n5476) );
  XOR U2350 ( .A(y[1195]), .B(n5459), .Z(n5460) );
  XOR U2351 ( .A(y[1199]), .B(n5443), .Z(n5444) );
  XOR U2352 ( .A(y[1203]), .B(n5427), .Z(n5428) );
  XOR U2353 ( .A(y[1207]), .B(n5411), .Z(n5412) );
  XOR U2354 ( .A(y[1211]), .B(n5395), .Z(n5396) );
  XOR U2355 ( .A(y[1215]), .B(n5379), .Z(n5380) );
  XOR U2356 ( .A(y[1219]), .B(n5363), .Z(n5364) );
  XOR U2357 ( .A(y[1223]), .B(n5347), .Z(n5348) );
  XOR U2358 ( .A(y[1227]), .B(n5331), .Z(n5332) );
  XOR U2359 ( .A(y[1231]), .B(n5315), .Z(n5316) );
  XOR U2360 ( .A(y[1235]), .B(n5299), .Z(n5300) );
  XOR U2361 ( .A(y[1239]), .B(n5283), .Z(n5284) );
  XOR U2362 ( .A(y[1243]), .B(n5267), .Z(n5268) );
  XOR U2363 ( .A(y[1247]), .B(n5251), .Z(n5252) );
  XOR U2364 ( .A(y[1251]), .B(n5235), .Z(n5236) );
  XOR U2365 ( .A(y[1255]), .B(n5219), .Z(n5220) );
  XOR U2366 ( .A(y[1259]), .B(n5203), .Z(n5204) );
  XOR U2367 ( .A(y[1263]), .B(n5187), .Z(n5188) );
  XOR U2368 ( .A(y[1267]), .B(n5171), .Z(n5172) );
  XOR U2369 ( .A(y[1271]), .B(n5155), .Z(n5156) );
  XOR U2370 ( .A(y[1275]), .B(n5139), .Z(n5140) );
  XOR U2371 ( .A(y[1279]), .B(n5123), .Z(n5124) );
  XOR U2372 ( .A(y[1283]), .B(n5107), .Z(n5108) );
  XOR U2373 ( .A(y[1287]), .B(n5091), .Z(n5092) );
  XOR U2374 ( .A(y[1291]), .B(n5075), .Z(n5076) );
  XOR U2375 ( .A(y[1295]), .B(n5059), .Z(n5060) );
  XOR U2376 ( .A(y[1299]), .B(n5043), .Z(n5044) );
  XOR U2377 ( .A(y[1303]), .B(n5027), .Z(n5028) );
  XOR U2378 ( .A(y[1307]), .B(n5011), .Z(n5012) );
  XOR U2379 ( .A(y[1311]), .B(n4995), .Z(n4996) );
  XOR U2380 ( .A(y[1315]), .B(n4979), .Z(n4980) );
  XOR U2381 ( .A(y[1319]), .B(n4963), .Z(n4964) );
  XOR U2382 ( .A(y[1323]), .B(n4947), .Z(n4948) );
  XOR U2383 ( .A(y[1327]), .B(n4931), .Z(n4932) );
  XOR U2384 ( .A(y[1331]), .B(n4915), .Z(n4916) );
  XOR U2385 ( .A(y[1335]), .B(n4899), .Z(n4900) );
  XOR U2386 ( .A(y[1339]), .B(n4883), .Z(n4884) );
  XOR U2387 ( .A(y[1343]), .B(n4867), .Z(n4868) );
  XOR U2388 ( .A(y[1347]), .B(n4851), .Z(n4852) );
  XOR U2389 ( .A(y[1351]), .B(n4835), .Z(n4836) );
  XOR U2390 ( .A(y[1355]), .B(n4819), .Z(n4820) );
  XOR U2391 ( .A(y[1359]), .B(n4803), .Z(n4804) );
  XOR U2392 ( .A(y[1363]), .B(n4787), .Z(n4788) );
  XOR U2393 ( .A(y[1367]), .B(n4771), .Z(n4772) );
  XOR U2394 ( .A(y[1371]), .B(n4755), .Z(n4756) );
  XOR U2395 ( .A(y[1375]), .B(n4739), .Z(n4740) );
  XOR U2396 ( .A(y[1379]), .B(n4723), .Z(n4724) );
  XOR U2397 ( .A(y[1383]), .B(n4707), .Z(n4708) );
  XOR U2398 ( .A(y[1387]), .B(n4691), .Z(n4692) );
  XOR U2399 ( .A(y[1391]), .B(n4675), .Z(n4676) );
  XOR U2400 ( .A(y[1395]), .B(n4659), .Z(n4660) );
  XOR U2401 ( .A(y[1399]), .B(n4643), .Z(n4644) );
  XOR U2402 ( .A(y[1403]), .B(n4627), .Z(n4628) );
  XOR U2403 ( .A(y[1407]), .B(n4611), .Z(n4612) );
  XOR U2404 ( .A(y[1411]), .B(n4595), .Z(n4596) );
  XOR U2405 ( .A(y[1415]), .B(n4579), .Z(n4580) );
  XOR U2406 ( .A(y[1419]), .B(n4563), .Z(n4564) );
  XOR U2407 ( .A(y[1423]), .B(n4547), .Z(n4548) );
  XOR U2408 ( .A(y[1427]), .B(n4531), .Z(n4532) );
  XOR U2409 ( .A(y[1431]), .B(n4515), .Z(n4516) );
  XOR U2410 ( .A(y[1435]), .B(n4499), .Z(n4500) );
  XOR U2411 ( .A(y[1439]), .B(n4483), .Z(n4484) );
  XOR U2412 ( .A(y[1443]), .B(n4467), .Z(n4468) );
  XOR U2413 ( .A(y[1447]), .B(n4451), .Z(n4452) );
  XOR U2414 ( .A(y[1451]), .B(n4435), .Z(n4436) );
  XOR U2415 ( .A(y[1455]), .B(n4419), .Z(n4420) );
  XOR U2416 ( .A(y[1459]), .B(n4403), .Z(n4404) );
  XOR U2417 ( .A(y[1463]), .B(n4387), .Z(n4388) );
  XOR U2418 ( .A(y[1467]), .B(n4371), .Z(n4372) );
  XOR U2419 ( .A(y[1471]), .B(n4355), .Z(n4356) );
  XOR U2420 ( .A(y[1475]), .B(n4339), .Z(n4340) );
  XOR U2421 ( .A(y[1479]), .B(n4323), .Z(n4324) );
  XOR U2422 ( .A(y[1483]), .B(n4307), .Z(n4308) );
  XOR U2423 ( .A(y[1487]), .B(n4291), .Z(n4292) );
  XOR U2424 ( .A(y[1491]), .B(n4275), .Z(n4276) );
  XOR U2425 ( .A(y[1495]), .B(n4259), .Z(n4260) );
  XOR U2426 ( .A(y[1499]), .B(n4243), .Z(n4244) );
  XOR U2427 ( .A(y[1503]), .B(n4227), .Z(n4228) );
  XOR U2428 ( .A(y[1507]), .B(n4211), .Z(n4212) );
  XOR U2429 ( .A(y[1511]), .B(n4195), .Z(n4196) );
  XOR U2430 ( .A(y[1515]), .B(n4179), .Z(n4180) );
  XOR U2431 ( .A(y[1519]), .B(n4163), .Z(n4164) );
  XOR U2432 ( .A(y[1523]), .B(n4147), .Z(n4148) );
  XOR U2433 ( .A(y[1527]), .B(n4131), .Z(n4132) );
  XOR U2434 ( .A(y[1531]), .B(n4115), .Z(n4116) );
  XOR U2435 ( .A(y[1535]), .B(n4099), .Z(n4100) );
  XOR U2436 ( .A(y[1539]), .B(n4083), .Z(n4084) );
  XOR U2437 ( .A(y[1543]), .B(n4067), .Z(n4068) );
  XOR U2438 ( .A(y[1547]), .B(n4051), .Z(n4052) );
  XOR U2439 ( .A(y[1551]), .B(n4035), .Z(n4036) );
  XOR U2440 ( .A(y[1555]), .B(n4019), .Z(n4020) );
  XOR U2441 ( .A(y[1559]), .B(n4003), .Z(n4004) );
  XOR U2442 ( .A(y[1563]), .B(n3987), .Z(n3988) );
  XOR U2443 ( .A(y[1567]), .B(n3971), .Z(n3972) );
  XOR U2444 ( .A(y[1571]), .B(n3955), .Z(n3956) );
  XOR U2445 ( .A(y[1575]), .B(n3939), .Z(n3940) );
  XOR U2446 ( .A(y[1579]), .B(n3923), .Z(n3924) );
  XOR U2447 ( .A(y[1583]), .B(n3907), .Z(n3908) );
  XOR U2448 ( .A(y[1587]), .B(n3891), .Z(n3892) );
  XOR U2449 ( .A(y[1591]), .B(n3875), .Z(n3876) );
  XOR U2450 ( .A(y[1595]), .B(n3859), .Z(n3860) );
  XOR U2451 ( .A(y[1599]), .B(n3843), .Z(n3844) );
  XOR U2452 ( .A(y[1603]), .B(n3827), .Z(n3828) );
  XOR U2453 ( .A(y[1607]), .B(n3811), .Z(n3812) );
  XOR U2454 ( .A(y[1611]), .B(n3795), .Z(n3796) );
  XOR U2455 ( .A(y[1615]), .B(n3779), .Z(n3780) );
  XOR U2456 ( .A(y[1619]), .B(n3763), .Z(n3764) );
  XOR U2457 ( .A(y[1623]), .B(n3747), .Z(n3748) );
  XOR U2458 ( .A(y[1627]), .B(n3731), .Z(n3732) );
  XOR U2459 ( .A(y[1631]), .B(n3715), .Z(n3716) );
  XOR U2460 ( .A(y[1635]), .B(n3699), .Z(n3700) );
  XOR U2461 ( .A(y[1639]), .B(n3683), .Z(n3684) );
  XOR U2462 ( .A(y[1643]), .B(n3667), .Z(n3668) );
  XOR U2463 ( .A(y[1647]), .B(n3651), .Z(n3652) );
  XOR U2464 ( .A(y[1651]), .B(n3635), .Z(n3636) );
  XOR U2465 ( .A(y[1655]), .B(n3619), .Z(n3620) );
  XOR U2466 ( .A(y[1659]), .B(n3603), .Z(n3604) );
  XOR U2467 ( .A(y[1663]), .B(n3587), .Z(n3588) );
  XOR U2468 ( .A(y[1667]), .B(n3571), .Z(n3572) );
  XOR U2469 ( .A(y[1671]), .B(n3555), .Z(n3556) );
  XOR U2470 ( .A(y[1675]), .B(n3539), .Z(n3540) );
  XOR U2471 ( .A(y[1679]), .B(n3523), .Z(n3524) );
  XOR U2472 ( .A(y[1683]), .B(n3507), .Z(n3508) );
  XOR U2473 ( .A(y[1687]), .B(n3491), .Z(n3492) );
  XOR U2474 ( .A(y[1691]), .B(n3475), .Z(n3476) );
  XOR U2475 ( .A(y[1695]), .B(n3459), .Z(n3460) );
  XOR U2476 ( .A(y[1699]), .B(n3443), .Z(n3444) );
  XOR U2477 ( .A(y[1703]), .B(n3427), .Z(n3428) );
  XOR U2478 ( .A(y[1707]), .B(n3411), .Z(n3412) );
  XOR U2479 ( .A(y[1711]), .B(n3395), .Z(n3396) );
  XOR U2480 ( .A(y[1715]), .B(n3379), .Z(n3380) );
  XOR U2481 ( .A(y[1719]), .B(n3363), .Z(n3364) );
  XOR U2482 ( .A(y[1723]), .B(n3347), .Z(n3348) );
  XOR U2483 ( .A(y[1727]), .B(n3331), .Z(n3332) );
  XOR U2484 ( .A(y[1731]), .B(n3315), .Z(n3316) );
  XOR U2485 ( .A(y[1735]), .B(n3299), .Z(n3300) );
  XOR U2486 ( .A(y[1739]), .B(n3283), .Z(n3284) );
  XOR U2487 ( .A(y[1743]), .B(n3267), .Z(n3268) );
  XOR U2488 ( .A(y[1747]), .B(n3251), .Z(n3252) );
  XOR U2489 ( .A(y[1751]), .B(n3235), .Z(n3236) );
  XOR U2490 ( .A(y[1755]), .B(n3219), .Z(n3220) );
  XOR U2491 ( .A(y[1759]), .B(n3203), .Z(n3204) );
  XOR U2492 ( .A(y[1763]), .B(n3187), .Z(n3188) );
  XOR U2493 ( .A(y[1767]), .B(n3171), .Z(n3172) );
  XOR U2494 ( .A(y[1771]), .B(n3155), .Z(n3156) );
  XOR U2495 ( .A(y[1775]), .B(n3139), .Z(n3140) );
  XOR U2496 ( .A(y[1779]), .B(n3123), .Z(n3124) );
  XOR U2497 ( .A(y[1783]), .B(n3107), .Z(n3108) );
  XOR U2498 ( .A(y[1787]), .B(n3091), .Z(n3092) );
  XOR U2499 ( .A(y[1791]), .B(n3075), .Z(n3076) );
  XOR U2500 ( .A(y[1795]), .B(n3059), .Z(n3060) );
  XOR U2501 ( .A(y[1799]), .B(n3043), .Z(n3044) );
  XOR U2502 ( .A(y[1803]), .B(n3027), .Z(n3028) );
  XOR U2503 ( .A(y[1807]), .B(n3011), .Z(n3012) );
  XOR U2504 ( .A(y[1811]), .B(n2995), .Z(n2996) );
  XOR U2505 ( .A(y[1815]), .B(n2979), .Z(n2980) );
  XOR U2506 ( .A(y[1819]), .B(n2963), .Z(n2964) );
  XOR U2507 ( .A(y[1823]), .B(n2947), .Z(n2948) );
  XOR U2508 ( .A(y[1827]), .B(n2931), .Z(n2932) );
  XOR U2509 ( .A(y[1831]), .B(n2915), .Z(n2916) );
  XOR U2510 ( .A(y[1835]), .B(n2899), .Z(n2900) );
  XOR U2511 ( .A(y[1839]), .B(n2883), .Z(n2884) );
  XOR U2512 ( .A(y[1843]), .B(n2867), .Z(n2868) );
  XOR U2513 ( .A(y[1847]), .B(n2851), .Z(n2852) );
  XOR U2514 ( .A(y[1851]), .B(n2835), .Z(n2836) );
  XOR U2515 ( .A(y[1855]), .B(n2819), .Z(n2820) );
  XOR U2516 ( .A(y[1859]), .B(n2803), .Z(n2804) );
  XOR U2517 ( .A(y[1863]), .B(n2787), .Z(n2788) );
  XOR U2518 ( .A(y[1867]), .B(n2771), .Z(n2772) );
  XOR U2519 ( .A(y[1871]), .B(n2755), .Z(n2756) );
  XOR U2520 ( .A(y[1875]), .B(n2739), .Z(n2740) );
  XOR U2521 ( .A(y[1879]), .B(n2723), .Z(n2724) );
  XOR U2522 ( .A(y[1883]), .B(n2707), .Z(n2708) );
  XOR U2523 ( .A(y[1887]), .B(n2691), .Z(n2692) );
  XOR U2524 ( .A(y[1891]), .B(n2675), .Z(n2676) );
  XOR U2525 ( .A(y[1895]), .B(n2659), .Z(n2660) );
  XOR U2526 ( .A(y[1899]), .B(n2643), .Z(n2644) );
  XOR U2527 ( .A(y[1903]), .B(n2627), .Z(n2628) );
  XOR U2528 ( .A(y[1907]), .B(n2611), .Z(n2612) );
  XOR U2529 ( .A(y[1911]), .B(n2595), .Z(n2596) );
  XOR U2530 ( .A(y[1915]), .B(n2579), .Z(n2580) );
  XOR U2531 ( .A(y[1919]), .B(n2563), .Z(n2564) );
  XOR U2532 ( .A(y[1923]), .B(n2547), .Z(n2548) );
  XOR U2533 ( .A(y[1927]), .B(n2531), .Z(n2532) );
  XOR U2534 ( .A(y[1931]), .B(n2515), .Z(n2516) );
  XOR U2535 ( .A(y[1935]), .B(n2499), .Z(n2500) );
  XOR U2536 ( .A(y[1939]), .B(n2483), .Z(n2484) );
  XOR U2537 ( .A(y[1943]), .B(n2467), .Z(n2468) );
  XOR U2538 ( .A(y[1947]), .B(n2451), .Z(n2452) );
  XOR U2539 ( .A(y[1951]), .B(n2435), .Z(n2436) );
  XOR U2540 ( .A(y[1955]), .B(n2419), .Z(n2420) );
  XOR U2541 ( .A(y[1959]), .B(n2403), .Z(n2404) );
  XOR U2542 ( .A(y[1963]), .B(n2387), .Z(n2388) );
  XOR U2543 ( .A(y[1967]), .B(n2371), .Z(n2372) );
  XOR U2544 ( .A(y[1971]), .B(n2355), .Z(n2356) );
  XOR U2545 ( .A(y[1975]), .B(n2339), .Z(n2340) );
  XOR U2546 ( .A(y[1979]), .B(n2323), .Z(n2324) );
  XOR U2547 ( .A(y[1983]), .B(n2307), .Z(n2308) );
  XOR U2548 ( .A(y[1987]), .B(n2291), .Z(n2292) );
  XOR U2549 ( .A(y[1991]), .B(n2275), .Z(n2276) );
  XOR U2550 ( .A(y[1995]), .B(n2259), .Z(n2260) );
  XOR U2551 ( .A(y[1999]), .B(n2243), .Z(n2244) );
  XOR U2552 ( .A(y[2003]), .B(n2227), .Z(n2228) );
  XOR U2553 ( .A(y[2007]), .B(n2211), .Z(n2212) );
  XOR U2554 ( .A(y[2011]), .B(n2195), .Z(n2196) );
  XOR U2555 ( .A(y[2015]), .B(n2179), .Z(n2180) );
  XOR U2556 ( .A(y[2019]), .B(n2163), .Z(n2164) );
  XOR U2557 ( .A(y[2023]), .B(n2147), .Z(n2148) );
  XOR U2558 ( .A(y[2027]), .B(n2131), .Z(n2132) );
  XOR U2559 ( .A(y[2031]), .B(n2115), .Z(n2116) );
  XOR U2560 ( .A(y[2035]), .B(n2099), .Z(n2100) );
  XOR U2561 ( .A(y[2039]), .B(n2083), .Z(n2084) );
  XOR U2562 ( .A(y[2043]), .B(n2067), .Z(n2068) );
  XOR U2563 ( .A(y[4]), .B(n10223), .Z(n10224) );
  XOR U2564 ( .A(y[8]), .B(n10207), .Z(n10208) );
  XOR U2565 ( .A(y[12]), .B(n10191), .Z(n10192) );
  XOR U2566 ( .A(y[16]), .B(n10175), .Z(n10176) );
  XOR U2567 ( .A(y[20]), .B(n10159), .Z(n10160) );
  XOR U2568 ( .A(y[24]), .B(n10143), .Z(n10144) );
  XOR U2569 ( .A(y[28]), .B(n10127), .Z(n10128) );
  XOR U2570 ( .A(y[32]), .B(n10111), .Z(n10112) );
  XOR U2571 ( .A(y[36]), .B(n10095), .Z(n10096) );
  XOR U2572 ( .A(y[40]), .B(n10079), .Z(n10080) );
  XOR U2573 ( .A(y[44]), .B(n10063), .Z(n10064) );
  XOR U2574 ( .A(y[48]), .B(n10047), .Z(n10048) );
  XOR U2575 ( .A(y[52]), .B(n10031), .Z(n10032) );
  XOR U2576 ( .A(y[56]), .B(n10015), .Z(n10016) );
  XOR U2577 ( .A(y[60]), .B(n9999), .Z(n10000) );
  XOR U2578 ( .A(y[64]), .B(n9983), .Z(n9984) );
  XOR U2579 ( .A(y[68]), .B(n9967), .Z(n9968) );
  XOR U2580 ( .A(y[72]), .B(n9951), .Z(n9952) );
  XOR U2581 ( .A(y[76]), .B(n9935), .Z(n9936) );
  XOR U2582 ( .A(y[80]), .B(n9919), .Z(n9920) );
  XOR U2583 ( .A(y[84]), .B(n9903), .Z(n9904) );
  XOR U2584 ( .A(y[88]), .B(n9887), .Z(n9888) );
  XOR U2585 ( .A(y[92]), .B(n9871), .Z(n9872) );
  XOR U2586 ( .A(y[96]), .B(n9855), .Z(n9856) );
  XOR U2587 ( .A(y[100]), .B(n9839), .Z(n9840) );
  XOR U2588 ( .A(y[104]), .B(n9823), .Z(n9824) );
  XOR U2589 ( .A(y[108]), .B(n9807), .Z(n9808) );
  XOR U2590 ( .A(y[112]), .B(n9791), .Z(n9792) );
  XOR U2591 ( .A(y[116]), .B(n9775), .Z(n9776) );
  XOR U2592 ( .A(y[120]), .B(n9759), .Z(n9760) );
  XOR U2593 ( .A(y[124]), .B(n9743), .Z(n9744) );
  XOR U2594 ( .A(y[128]), .B(n9727), .Z(n9728) );
  XOR U2595 ( .A(y[132]), .B(n9711), .Z(n9712) );
  XOR U2596 ( .A(y[136]), .B(n9695), .Z(n9696) );
  XOR U2597 ( .A(y[140]), .B(n9679), .Z(n9680) );
  XOR U2598 ( .A(y[144]), .B(n9663), .Z(n9664) );
  XOR U2599 ( .A(y[148]), .B(n9647), .Z(n9648) );
  XOR U2600 ( .A(y[152]), .B(n9631), .Z(n9632) );
  XOR U2601 ( .A(y[156]), .B(n9615), .Z(n9616) );
  XOR U2602 ( .A(y[160]), .B(n9599), .Z(n9600) );
  XOR U2603 ( .A(y[164]), .B(n9583), .Z(n9584) );
  XOR U2604 ( .A(y[168]), .B(n9567), .Z(n9568) );
  XOR U2605 ( .A(y[172]), .B(n9551), .Z(n9552) );
  XOR U2606 ( .A(y[176]), .B(n9535), .Z(n9536) );
  XOR U2607 ( .A(y[180]), .B(n9519), .Z(n9520) );
  XOR U2608 ( .A(y[184]), .B(n9503), .Z(n9504) );
  XOR U2609 ( .A(y[188]), .B(n9487), .Z(n9488) );
  XOR U2610 ( .A(y[192]), .B(n9471), .Z(n9472) );
  XOR U2611 ( .A(y[196]), .B(n9455), .Z(n9456) );
  XOR U2612 ( .A(y[200]), .B(n9439), .Z(n9440) );
  XOR U2613 ( .A(y[204]), .B(n9423), .Z(n9424) );
  XOR U2614 ( .A(y[208]), .B(n9407), .Z(n9408) );
  XOR U2615 ( .A(y[212]), .B(n9391), .Z(n9392) );
  XOR U2616 ( .A(y[216]), .B(n9375), .Z(n9376) );
  XOR U2617 ( .A(y[220]), .B(n9359), .Z(n9360) );
  XOR U2618 ( .A(y[224]), .B(n9343), .Z(n9344) );
  XOR U2619 ( .A(y[228]), .B(n9327), .Z(n9328) );
  XOR U2620 ( .A(y[232]), .B(n9311), .Z(n9312) );
  XOR U2621 ( .A(y[236]), .B(n9295), .Z(n9296) );
  XOR U2622 ( .A(y[240]), .B(n9279), .Z(n9280) );
  XOR U2623 ( .A(y[244]), .B(n9263), .Z(n9264) );
  XOR U2624 ( .A(y[248]), .B(n9247), .Z(n9248) );
  XOR U2625 ( .A(y[252]), .B(n9231), .Z(n9232) );
  XOR U2626 ( .A(y[256]), .B(n9215), .Z(n9216) );
  XOR U2627 ( .A(y[260]), .B(n9199), .Z(n9200) );
  XOR U2628 ( .A(y[264]), .B(n9183), .Z(n9184) );
  XOR U2629 ( .A(y[268]), .B(n9167), .Z(n9168) );
  XOR U2630 ( .A(y[272]), .B(n9151), .Z(n9152) );
  XOR U2631 ( .A(y[276]), .B(n9135), .Z(n9136) );
  XOR U2632 ( .A(y[280]), .B(n9119), .Z(n9120) );
  XOR U2633 ( .A(y[284]), .B(n9103), .Z(n9104) );
  XOR U2634 ( .A(y[288]), .B(n9087), .Z(n9088) );
  XOR U2635 ( .A(y[292]), .B(n9071), .Z(n9072) );
  XOR U2636 ( .A(y[296]), .B(n9055), .Z(n9056) );
  XOR U2637 ( .A(y[300]), .B(n9039), .Z(n9040) );
  XOR U2638 ( .A(y[304]), .B(n9023), .Z(n9024) );
  XOR U2639 ( .A(y[308]), .B(n9007), .Z(n9008) );
  XOR U2640 ( .A(y[312]), .B(n8991), .Z(n8992) );
  XOR U2641 ( .A(y[316]), .B(n8975), .Z(n8976) );
  XOR U2642 ( .A(y[320]), .B(n8959), .Z(n8960) );
  XOR U2643 ( .A(y[324]), .B(n8943), .Z(n8944) );
  XOR U2644 ( .A(y[328]), .B(n8927), .Z(n8928) );
  XOR U2645 ( .A(y[332]), .B(n8911), .Z(n8912) );
  XOR U2646 ( .A(y[336]), .B(n8895), .Z(n8896) );
  XOR U2647 ( .A(y[340]), .B(n8879), .Z(n8880) );
  XOR U2648 ( .A(y[344]), .B(n8863), .Z(n8864) );
  XOR U2649 ( .A(y[348]), .B(n8847), .Z(n8848) );
  XOR U2650 ( .A(y[352]), .B(n8831), .Z(n8832) );
  XOR U2651 ( .A(y[356]), .B(n8815), .Z(n8816) );
  XOR U2652 ( .A(y[360]), .B(n8799), .Z(n8800) );
  XOR U2653 ( .A(y[364]), .B(n8783), .Z(n8784) );
  XOR U2654 ( .A(y[368]), .B(n8767), .Z(n8768) );
  XOR U2655 ( .A(y[372]), .B(n8751), .Z(n8752) );
  XOR U2656 ( .A(y[376]), .B(n8735), .Z(n8736) );
  XOR U2657 ( .A(y[380]), .B(n8719), .Z(n8720) );
  XOR U2658 ( .A(y[384]), .B(n8703), .Z(n8704) );
  XOR U2659 ( .A(y[388]), .B(n8687), .Z(n8688) );
  XOR U2660 ( .A(y[392]), .B(n8671), .Z(n8672) );
  XOR U2661 ( .A(y[396]), .B(n8655), .Z(n8656) );
  XOR U2662 ( .A(y[400]), .B(n8639), .Z(n8640) );
  XOR U2663 ( .A(y[404]), .B(n8623), .Z(n8624) );
  XOR U2664 ( .A(y[408]), .B(n8607), .Z(n8608) );
  XOR U2665 ( .A(y[412]), .B(n8591), .Z(n8592) );
  XOR U2666 ( .A(y[416]), .B(n8575), .Z(n8576) );
  XOR U2667 ( .A(y[420]), .B(n8559), .Z(n8560) );
  XOR U2668 ( .A(y[424]), .B(n8543), .Z(n8544) );
  XOR U2669 ( .A(y[428]), .B(n8527), .Z(n8528) );
  XOR U2670 ( .A(y[432]), .B(n8511), .Z(n8512) );
  XOR U2671 ( .A(y[436]), .B(n8495), .Z(n8496) );
  XOR U2672 ( .A(y[440]), .B(n8479), .Z(n8480) );
  XOR U2673 ( .A(y[444]), .B(n8463), .Z(n8464) );
  XOR U2674 ( .A(y[448]), .B(n8447), .Z(n8448) );
  XOR U2675 ( .A(y[452]), .B(n8431), .Z(n8432) );
  XOR U2676 ( .A(y[456]), .B(n8415), .Z(n8416) );
  XOR U2677 ( .A(y[460]), .B(n8399), .Z(n8400) );
  XOR U2678 ( .A(y[464]), .B(n8383), .Z(n8384) );
  XOR U2679 ( .A(y[468]), .B(n8367), .Z(n8368) );
  XOR U2680 ( .A(y[472]), .B(n8351), .Z(n8352) );
  XOR U2681 ( .A(y[476]), .B(n8335), .Z(n8336) );
  XOR U2682 ( .A(y[480]), .B(n8319), .Z(n8320) );
  XOR U2683 ( .A(y[484]), .B(n8303), .Z(n8304) );
  XOR U2684 ( .A(y[488]), .B(n8287), .Z(n8288) );
  XOR U2685 ( .A(y[492]), .B(n8271), .Z(n8272) );
  XOR U2686 ( .A(y[496]), .B(n8255), .Z(n8256) );
  XOR U2687 ( .A(y[500]), .B(n8239), .Z(n8240) );
  XOR U2688 ( .A(y[504]), .B(n8223), .Z(n8224) );
  XOR U2689 ( .A(y[508]), .B(n8207), .Z(n8208) );
  XOR U2690 ( .A(y[512]), .B(n8191), .Z(n8192) );
  XOR U2691 ( .A(y[516]), .B(n8175), .Z(n8176) );
  XOR U2692 ( .A(y[520]), .B(n8159), .Z(n8160) );
  XOR U2693 ( .A(y[524]), .B(n8143), .Z(n8144) );
  XOR U2694 ( .A(y[528]), .B(n8127), .Z(n8128) );
  XOR U2695 ( .A(y[532]), .B(n8111), .Z(n8112) );
  XOR U2696 ( .A(y[536]), .B(n8095), .Z(n8096) );
  XOR U2697 ( .A(y[540]), .B(n8079), .Z(n8080) );
  XOR U2698 ( .A(y[544]), .B(n8063), .Z(n8064) );
  XOR U2699 ( .A(y[548]), .B(n8047), .Z(n8048) );
  XOR U2700 ( .A(y[552]), .B(n8031), .Z(n8032) );
  XOR U2701 ( .A(y[556]), .B(n8015), .Z(n8016) );
  XOR U2702 ( .A(y[560]), .B(n7999), .Z(n8000) );
  XOR U2703 ( .A(y[564]), .B(n7983), .Z(n7984) );
  XOR U2704 ( .A(y[568]), .B(n7967), .Z(n7968) );
  XOR U2705 ( .A(y[572]), .B(n7951), .Z(n7952) );
  XOR U2706 ( .A(y[576]), .B(n7935), .Z(n7936) );
  XOR U2707 ( .A(y[580]), .B(n7919), .Z(n7920) );
  XOR U2708 ( .A(y[584]), .B(n7903), .Z(n7904) );
  XOR U2709 ( .A(y[588]), .B(n7887), .Z(n7888) );
  XOR U2710 ( .A(y[592]), .B(n7871), .Z(n7872) );
  XOR U2711 ( .A(y[596]), .B(n7855), .Z(n7856) );
  XOR U2712 ( .A(y[600]), .B(n7839), .Z(n7840) );
  XOR U2713 ( .A(y[604]), .B(n7823), .Z(n7824) );
  XOR U2714 ( .A(y[608]), .B(n7807), .Z(n7808) );
  XOR U2715 ( .A(y[612]), .B(n7791), .Z(n7792) );
  XOR U2716 ( .A(y[616]), .B(n7775), .Z(n7776) );
  XOR U2717 ( .A(y[620]), .B(n7759), .Z(n7760) );
  XOR U2718 ( .A(y[624]), .B(n7743), .Z(n7744) );
  XOR U2719 ( .A(y[628]), .B(n7727), .Z(n7728) );
  XOR U2720 ( .A(y[632]), .B(n7711), .Z(n7712) );
  XOR U2721 ( .A(y[636]), .B(n7695), .Z(n7696) );
  XOR U2722 ( .A(y[640]), .B(n7679), .Z(n7680) );
  XOR U2723 ( .A(y[644]), .B(n7663), .Z(n7664) );
  XOR U2724 ( .A(y[648]), .B(n7647), .Z(n7648) );
  XOR U2725 ( .A(y[652]), .B(n7631), .Z(n7632) );
  XOR U2726 ( .A(y[656]), .B(n7615), .Z(n7616) );
  XOR U2727 ( .A(y[660]), .B(n7599), .Z(n7600) );
  XOR U2728 ( .A(y[664]), .B(n7583), .Z(n7584) );
  XOR U2729 ( .A(y[668]), .B(n7567), .Z(n7568) );
  XOR U2730 ( .A(y[672]), .B(n7551), .Z(n7552) );
  XOR U2731 ( .A(y[676]), .B(n7535), .Z(n7536) );
  XOR U2732 ( .A(y[680]), .B(n7519), .Z(n7520) );
  XOR U2733 ( .A(y[684]), .B(n7503), .Z(n7504) );
  XOR U2734 ( .A(y[688]), .B(n7487), .Z(n7488) );
  XOR U2735 ( .A(y[692]), .B(n7471), .Z(n7472) );
  XOR U2736 ( .A(y[696]), .B(n7455), .Z(n7456) );
  XOR U2737 ( .A(y[700]), .B(n7439), .Z(n7440) );
  XOR U2738 ( .A(y[704]), .B(n7423), .Z(n7424) );
  XOR U2739 ( .A(y[708]), .B(n7407), .Z(n7408) );
  XOR U2740 ( .A(y[712]), .B(n7391), .Z(n7392) );
  XOR U2741 ( .A(y[716]), .B(n7375), .Z(n7376) );
  XOR U2742 ( .A(y[720]), .B(n7359), .Z(n7360) );
  XOR U2743 ( .A(y[724]), .B(n7343), .Z(n7344) );
  XOR U2744 ( .A(y[728]), .B(n7327), .Z(n7328) );
  XOR U2745 ( .A(y[732]), .B(n7311), .Z(n7312) );
  XOR U2746 ( .A(y[736]), .B(n7295), .Z(n7296) );
  XOR U2747 ( .A(y[740]), .B(n7279), .Z(n7280) );
  XOR U2748 ( .A(y[744]), .B(n7263), .Z(n7264) );
  XOR U2749 ( .A(y[748]), .B(n7247), .Z(n7248) );
  XOR U2750 ( .A(y[752]), .B(n7231), .Z(n7232) );
  XOR U2751 ( .A(y[756]), .B(n7215), .Z(n7216) );
  XOR U2752 ( .A(y[760]), .B(n7199), .Z(n7200) );
  XOR U2753 ( .A(y[764]), .B(n7183), .Z(n7184) );
  XOR U2754 ( .A(y[768]), .B(n7167), .Z(n7168) );
  XOR U2755 ( .A(y[772]), .B(n7151), .Z(n7152) );
  XOR U2756 ( .A(y[776]), .B(n7135), .Z(n7136) );
  XOR U2757 ( .A(y[780]), .B(n7119), .Z(n7120) );
  XOR U2758 ( .A(y[784]), .B(n7103), .Z(n7104) );
  XOR U2759 ( .A(y[788]), .B(n7087), .Z(n7088) );
  XOR U2760 ( .A(y[792]), .B(n7071), .Z(n7072) );
  XOR U2761 ( .A(y[796]), .B(n7055), .Z(n7056) );
  XOR U2762 ( .A(y[800]), .B(n7039), .Z(n7040) );
  XOR U2763 ( .A(y[804]), .B(n7023), .Z(n7024) );
  XOR U2764 ( .A(y[808]), .B(n7007), .Z(n7008) );
  XOR U2765 ( .A(y[812]), .B(n6991), .Z(n6992) );
  XOR U2766 ( .A(y[816]), .B(n6975), .Z(n6976) );
  XOR U2767 ( .A(y[820]), .B(n6959), .Z(n6960) );
  XOR U2768 ( .A(y[824]), .B(n6943), .Z(n6944) );
  XOR U2769 ( .A(y[828]), .B(n6927), .Z(n6928) );
  XOR U2770 ( .A(y[832]), .B(n6911), .Z(n6912) );
  XOR U2771 ( .A(y[836]), .B(n6895), .Z(n6896) );
  XOR U2772 ( .A(y[840]), .B(n6879), .Z(n6880) );
  XOR U2773 ( .A(y[844]), .B(n6863), .Z(n6864) );
  XOR U2774 ( .A(y[848]), .B(n6847), .Z(n6848) );
  XOR U2775 ( .A(y[852]), .B(n6831), .Z(n6832) );
  XOR U2776 ( .A(y[856]), .B(n6815), .Z(n6816) );
  XOR U2777 ( .A(y[860]), .B(n6799), .Z(n6800) );
  XOR U2778 ( .A(y[864]), .B(n6783), .Z(n6784) );
  XOR U2779 ( .A(y[868]), .B(n6767), .Z(n6768) );
  XOR U2780 ( .A(y[872]), .B(n6751), .Z(n6752) );
  XOR U2781 ( .A(y[876]), .B(n6735), .Z(n6736) );
  XOR U2782 ( .A(y[880]), .B(n6719), .Z(n6720) );
  XOR U2783 ( .A(y[884]), .B(n6703), .Z(n6704) );
  XOR U2784 ( .A(y[888]), .B(n6687), .Z(n6688) );
  XOR U2785 ( .A(y[892]), .B(n6671), .Z(n6672) );
  XOR U2786 ( .A(y[896]), .B(n6655), .Z(n6656) );
  XOR U2787 ( .A(y[900]), .B(n6639), .Z(n6640) );
  XOR U2788 ( .A(y[904]), .B(n6623), .Z(n6624) );
  XOR U2789 ( .A(y[908]), .B(n6607), .Z(n6608) );
  XOR U2790 ( .A(y[912]), .B(n6591), .Z(n6592) );
  XOR U2791 ( .A(y[916]), .B(n6575), .Z(n6576) );
  XOR U2792 ( .A(y[920]), .B(n6559), .Z(n6560) );
  XOR U2793 ( .A(y[924]), .B(n6543), .Z(n6544) );
  XOR U2794 ( .A(y[928]), .B(n6527), .Z(n6528) );
  XOR U2795 ( .A(y[932]), .B(n6511), .Z(n6512) );
  XOR U2796 ( .A(y[936]), .B(n6495), .Z(n6496) );
  XOR U2797 ( .A(y[940]), .B(n6479), .Z(n6480) );
  XOR U2798 ( .A(y[944]), .B(n6463), .Z(n6464) );
  XOR U2799 ( .A(y[948]), .B(n6447), .Z(n6448) );
  XOR U2800 ( .A(y[952]), .B(n6431), .Z(n6432) );
  XOR U2801 ( .A(y[956]), .B(n6415), .Z(n6416) );
  XOR U2802 ( .A(y[960]), .B(n6399), .Z(n6400) );
  XOR U2803 ( .A(y[964]), .B(n6383), .Z(n6384) );
  XOR U2804 ( .A(y[968]), .B(n6367), .Z(n6368) );
  XOR U2805 ( .A(y[972]), .B(n6351), .Z(n6352) );
  XOR U2806 ( .A(y[976]), .B(n6335), .Z(n6336) );
  XOR U2807 ( .A(y[980]), .B(n6319), .Z(n6320) );
  XOR U2808 ( .A(y[984]), .B(n6303), .Z(n6304) );
  XOR U2809 ( .A(y[988]), .B(n6287), .Z(n6288) );
  XOR U2810 ( .A(y[992]), .B(n6271), .Z(n6272) );
  XOR U2811 ( .A(y[996]), .B(n6255), .Z(n6256) );
  XOR U2812 ( .A(y[1000]), .B(n6239), .Z(n6240) );
  XOR U2813 ( .A(y[1004]), .B(n6223), .Z(n6224) );
  XOR U2814 ( .A(y[1008]), .B(n6207), .Z(n6208) );
  XOR U2815 ( .A(y[1012]), .B(n6191), .Z(n6192) );
  XOR U2816 ( .A(y[1016]), .B(n6175), .Z(n6176) );
  XOR U2817 ( .A(y[1020]), .B(n6159), .Z(n6160) );
  XOR U2818 ( .A(y[1024]), .B(n6143), .Z(n6144) );
  XOR U2819 ( .A(y[1028]), .B(n6127), .Z(n6128) );
  XOR U2820 ( .A(y[1032]), .B(n6111), .Z(n6112) );
  XOR U2821 ( .A(y[1036]), .B(n6095), .Z(n6096) );
  XOR U2822 ( .A(y[1040]), .B(n6079), .Z(n6080) );
  XOR U2823 ( .A(y[1044]), .B(n6063), .Z(n6064) );
  XOR U2824 ( .A(y[1048]), .B(n6047), .Z(n6048) );
  XOR U2825 ( .A(y[1052]), .B(n6031), .Z(n6032) );
  XOR U2826 ( .A(y[1056]), .B(n6015), .Z(n6016) );
  XOR U2827 ( .A(y[1060]), .B(n5999), .Z(n6000) );
  XOR U2828 ( .A(y[1064]), .B(n5983), .Z(n5984) );
  XOR U2829 ( .A(y[1068]), .B(n5967), .Z(n5968) );
  XOR U2830 ( .A(y[1072]), .B(n5951), .Z(n5952) );
  XOR U2831 ( .A(y[1076]), .B(n5935), .Z(n5936) );
  XOR U2832 ( .A(y[1080]), .B(n5919), .Z(n5920) );
  XOR U2833 ( .A(y[1084]), .B(n5903), .Z(n5904) );
  XOR U2834 ( .A(y[1088]), .B(n5887), .Z(n5888) );
  XOR U2835 ( .A(y[1092]), .B(n5871), .Z(n5872) );
  XOR U2836 ( .A(y[1096]), .B(n5855), .Z(n5856) );
  XOR U2837 ( .A(y[1100]), .B(n5839), .Z(n5840) );
  XOR U2838 ( .A(y[1104]), .B(n5823), .Z(n5824) );
  XOR U2839 ( .A(y[1108]), .B(n5807), .Z(n5808) );
  XOR U2840 ( .A(y[1112]), .B(n5791), .Z(n5792) );
  XOR U2841 ( .A(y[1116]), .B(n5775), .Z(n5776) );
  XOR U2842 ( .A(y[1120]), .B(n5759), .Z(n5760) );
  XOR U2843 ( .A(y[1124]), .B(n5743), .Z(n5744) );
  XOR U2844 ( .A(y[1128]), .B(n5727), .Z(n5728) );
  XOR U2845 ( .A(y[1132]), .B(n5711), .Z(n5712) );
  XOR U2846 ( .A(y[1136]), .B(n5695), .Z(n5696) );
  XOR U2847 ( .A(y[1140]), .B(n5679), .Z(n5680) );
  XOR U2848 ( .A(y[1144]), .B(n5663), .Z(n5664) );
  XOR U2849 ( .A(y[1148]), .B(n5647), .Z(n5648) );
  XOR U2850 ( .A(y[1152]), .B(n5631), .Z(n5632) );
  XOR U2851 ( .A(y[1156]), .B(n5615), .Z(n5616) );
  XOR U2852 ( .A(y[1160]), .B(n5599), .Z(n5600) );
  XOR U2853 ( .A(y[1164]), .B(n5583), .Z(n5584) );
  XOR U2854 ( .A(y[1168]), .B(n5567), .Z(n5568) );
  XOR U2855 ( .A(y[1172]), .B(n5551), .Z(n5552) );
  XOR U2856 ( .A(y[1176]), .B(n5535), .Z(n5536) );
  XOR U2857 ( .A(y[1180]), .B(n5519), .Z(n5520) );
  XOR U2858 ( .A(y[1184]), .B(n5503), .Z(n5504) );
  XOR U2859 ( .A(y[1188]), .B(n5487), .Z(n5488) );
  XOR U2860 ( .A(y[1192]), .B(n5471), .Z(n5472) );
  XOR U2861 ( .A(y[1196]), .B(n5455), .Z(n5456) );
  XOR U2862 ( .A(y[1200]), .B(n5439), .Z(n5440) );
  XOR U2863 ( .A(y[1204]), .B(n5423), .Z(n5424) );
  XOR U2864 ( .A(y[1208]), .B(n5407), .Z(n5408) );
  XOR U2865 ( .A(y[1212]), .B(n5391), .Z(n5392) );
  XOR U2866 ( .A(y[1216]), .B(n5375), .Z(n5376) );
  XOR U2867 ( .A(y[1220]), .B(n5359), .Z(n5360) );
  XOR U2868 ( .A(y[1224]), .B(n5343), .Z(n5344) );
  XOR U2869 ( .A(y[1228]), .B(n5327), .Z(n5328) );
  XOR U2870 ( .A(y[1232]), .B(n5311), .Z(n5312) );
  XOR U2871 ( .A(y[1236]), .B(n5295), .Z(n5296) );
  XOR U2872 ( .A(y[1240]), .B(n5279), .Z(n5280) );
  XOR U2873 ( .A(y[1244]), .B(n5263), .Z(n5264) );
  XOR U2874 ( .A(y[1248]), .B(n5247), .Z(n5248) );
  XOR U2875 ( .A(y[1252]), .B(n5231), .Z(n5232) );
  XOR U2876 ( .A(y[1256]), .B(n5215), .Z(n5216) );
  XOR U2877 ( .A(y[1260]), .B(n5199), .Z(n5200) );
  XOR U2878 ( .A(y[1264]), .B(n5183), .Z(n5184) );
  XOR U2879 ( .A(y[1268]), .B(n5167), .Z(n5168) );
  XOR U2880 ( .A(y[1272]), .B(n5151), .Z(n5152) );
  XOR U2881 ( .A(y[1276]), .B(n5135), .Z(n5136) );
  XOR U2882 ( .A(y[1280]), .B(n5119), .Z(n5120) );
  XOR U2883 ( .A(y[1284]), .B(n5103), .Z(n5104) );
  XOR U2884 ( .A(y[1288]), .B(n5087), .Z(n5088) );
  XOR U2885 ( .A(y[1292]), .B(n5071), .Z(n5072) );
  XOR U2886 ( .A(y[1296]), .B(n5055), .Z(n5056) );
  XOR U2887 ( .A(y[1300]), .B(n5039), .Z(n5040) );
  XOR U2888 ( .A(y[1304]), .B(n5023), .Z(n5024) );
  XOR U2889 ( .A(y[1308]), .B(n5007), .Z(n5008) );
  XOR U2890 ( .A(y[1312]), .B(n4991), .Z(n4992) );
  XOR U2891 ( .A(y[1316]), .B(n4975), .Z(n4976) );
  XOR U2892 ( .A(y[1320]), .B(n4959), .Z(n4960) );
  XOR U2893 ( .A(y[1324]), .B(n4943), .Z(n4944) );
  XOR U2894 ( .A(y[1328]), .B(n4927), .Z(n4928) );
  XOR U2895 ( .A(y[1332]), .B(n4911), .Z(n4912) );
  XOR U2896 ( .A(y[1336]), .B(n4895), .Z(n4896) );
  XOR U2897 ( .A(y[1340]), .B(n4879), .Z(n4880) );
  XOR U2898 ( .A(y[1344]), .B(n4863), .Z(n4864) );
  XOR U2899 ( .A(y[1348]), .B(n4847), .Z(n4848) );
  XOR U2900 ( .A(y[1352]), .B(n4831), .Z(n4832) );
  XOR U2901 ( .A(y[1356]), .B(n4815), .Z(n4816) );
  XOR U2902 ( .A(y[1360]), .B(n4799), .Z(n4800) );
  XOR U2903 ( .A(y[1364]), .B(n4783), .Z(n4784) );
  XOR U2904 ( .A(y[1368]), .B(n4767), .Z(n4768) );
  XOR U2905 ( .A(y[1372]), .B(n4751), .Z(n4752) );
  XOR U2906 ( .A(y[1376]), .B(n4735), .Z(n4736) );
  XOR U2907 ( .A(y[1380]), .B(n4719), .Z(n4720) );
  XOR U2908 ( .A(y[1384]), .B(n4703), .Z(n4704) );
  XOR U2909 ( .A(y[1388]), .B(n4687), .Z(n4688) );
  XOR U2910 ( .A(y[1392]), .B(n4671), .Z(n4672) );
  XOR U2911 ( .A(y[1396]), .B(n4655), .Z(n4656) );
  XOR U2912 ( .A(y[1400]), .B(n4639), .Z(n4640) );
  XOR U2913 ( .A(y[1404]), .B(n4623), .Z(n4624) );
  XOR U2914 ( .A(y[1408]), .B(n4607), .Z(n4608) );
  XOR U2915 ( .A(y[1412]), .B(n4591), .Z(n4592) );
  XOR U2916 ( .A(y[1416]), .B(n4575), .Z(n4576) );
  XOR U2917 ( .A(y[1420]), .B(n4559), .Z(n4560) );
  XOR U2918 ( .A(y[1424]), .B(n4543), .Z(n4544) );
  XOR U2919 ( .A(y[1428]), .B(n4527), .Z(n4528) );
  XOR U2920 ( .A(y[1432]), .B(n4511), .Z(n4512) );
  XOR U2921 ( .A(y[1436]), .B(n4495), .Z(n4496) );
  XOR U2922 ( .A(y[1440]), .B(n4479), .Z(n4480) );
  XOR U2923 ( .A(y[1444]), .B(n4463), .Z(n4464) );
  XOR U2924 ( .A(y[1448]), .B(n4447), .Z(n4448) );
  XOR U2925 ( .A(y[1452]), .B(n4431), .Z(n4432) );
  XOR U2926 ( .A(y[1456]), .B(n4415), .Z(n4416) );
  XOR U2927 ( .A(y[1460]), .B(n4399), .Z(n4400) );
  XOR U2928 ( .A(y[1464]), .B(n4383), .Z(n4384) );
  XOR U2929 ( .A(y[1468]), .B(n4367), .Z(n4368) );
  XOR U2930 ( .A(y[1472]), .B(n4351), .Z(n4352) );
  XOR U2931 ( .A(y[1476]), .B(n4335), .Z(n4336) );
  XOR U2932 ( .A(y[1480]), .B(n4319), .Z(n4320) );
  XOR U2933 ( .A(y[1484]), .B(n4303), .Z(n4304) );
  XOR U2934 ( .A(y[1488]), .B(n4287), .Z(n4288) );
  XOR U2935 ( .A(y[1492]), .B(n4271), .Z(n4272) );
  XOR U2936 ( .A(y[1496]), .B(n4255), .Z(n4256) );
  XOR U2937 ( .A(y[1500]), .B(n4239), .Z(n4240) );
  XOR U2938 ( .A(y[1504]), .B(n4223), .Z(n4224) );
  XOR U2939 ( .A(y[1508]), .B(n4207), .Z(n4208) );
  XOR U2940 ( .A(y[1512]), .B(n4191), .Z(n4192) );
  XOR U2941 ( .A(y[1516]), .B(n4175), .Z(n4176) );
  XOR U2942 ( .A(y[1520]), .B(n4159), .Z(n4160) );
  XOR U2943 ( .A(y[1524]), .B(n4143), .Z(n4144) );
  XOR U2944 ( .A(y[1528]), .B(n4127), .Z(n4128) );
  XOR U2945 ( .A(y[1532]), .B(n4111), .Z(n4112) );
  XOR U2946 ( .A(y[1536]), .B(n4095), .Z(n4096) );
  XOR U2947 ( .A(y[1540]), .B(n4079), .Z(n4080) );
  XOR U2948 ( .A(y[1544]), .B(n4063), .Z(n4064) );
  XOR U2949 ( .A(y[1548]), .B(n4047), .Z(n4048) );
  XOR U2950 ( .A(y[1552]), .B(n4031), .Z(n4032) );
  XOR U2951 ( .A(y[1556]), .B(n4015), .Z(n4016) );
  XOR U2952 ( .A(y[1560]), .B(n3999), .Z(n4000) );
  XOR U2953 ( .A(y[1564]), .B(n3983), .Z(n3984) );
  XOR U2954 ( .A(y[1568]), .B(n3967), .Z(n3968) );
  XOR U2955 ( .A(y[1572]), .B(n3951), .Z(n3952) );
  XOR U2956 ( .A(y[1576]), .B(n3935), .Z(n3936) );
  XOR U2957 ( .A(y[1580]), .B(n3919), .Z(n3920) );
  XOR U2958 ( .A(y[1584]), .B(n3903), .Z(n3904) );
  XOR U2959 ( .A(y[1588]), .B(n3887), .Z(n3888) );
  XOR U2960 ( .A(y[1592]), .B(n3871), .Z(n3872) );
  XOR U2961 ( .A(y[1596]), .B(n3855), .Z(n3856) );
  XOR U2962 ( .A(y[1600]), .B(n3839), .Z(n3840) );
  XOR U2963 ( .A(y[1604]), .B(n3823), .Z(n3824) );
  XOR U2964 ( .A(y[1608]), .B(n3807), .Z(n3808) );
  XOR U2965 ( .A(y[1612]), .B(n3791), .Z(n3792) );
  XOR U2966 ( .A(y[1616]), .B(n3775), .Z(n3776) );
  XOR U2967 ( .A(y[1620]), .B(n3759), .Z(n3760) );
  XOR U2968 ( .A(y[1624]), .B(n3743), .Z(n3744) );
  XOR U2969 ( .A(y[1628]), .B(n3727), .Z(n3728) );
  XOR U2970 ( .A(y[1632]), .B(n3711), .Z(n3712) );
  XOR U2971 ( .A(y[1636]), .B(n3695), .Z(n3696) );
  XOR U2972 ( .A(y[1640]), .B(n3679), .Z(n3680) );
  XOR U2973 ( .A(y[1644]), .B(n3663), .Z(n3664) );
  XOR U2974 ( .A(y[1648]), .B(n3647), .Z(n3648) );
  XOR U2975 ( .A(y[1652]), .B(n3631), .Z(n3632) );
  XOR U2976 ( .A(y[1656]), .B(n3615), .Z(n3616) );
  XOR U2977 ( .A(y[1660]), .B(n3599), .Z(n3600) );
  XOR U2978 ( .A(y[1664]), .B(n3583), .Z(n3584) );
  XOR U2979 ( .A(y[1668]), .B(n3567), .Z(n3568) );
  XOR U2980 ( .A(y[1672]), .B(n3551), .Z(n3552) );
  XOR U2981 ( .A(y[1676]), .B(n3535), .Z(n3536) );
  XOR U2982 ( .A(y[1680]), .B(n3519), .Z(n3520) );
  XOR U2983 ( .A(y[1684]), .B(n3503), .Z(n3504) );
  XOR U2984 ( .A(y[1688]), .B(n3487), .Z(n3488) );
  XOR U2985 ( .A(y[1692]), .B(n3471), .Z(n3472) );
  XOR U2986 ( .A(y[1696]), .B(n3455), .Z(n3456) );
  XOR U2987 ( .A(y[1700]), .B(n3439), .Z(n3440) );
  XOR U2988 ( .A(y[1704]), .B(n3423), .Z(n3424) );
  XOR U2989 ( .A(y[1708]), .B(n3407), .Z(n3408) );
  XOR U2990 ( .A(y[1712]), .B(n3391), .Z(n3392) );
  XOR U2991 ( .A(y[1716]), .B(n3375), .Z(n3376) );
  XOR U2992 ( .A(y[1720]), .B(n3359), .Z(n3360) );
  XOR U2993 ( .A(y[1724]), .B(n3343), .Z(n3344) );
  XOR U2994 ( .A(y[1728]), .B(n3327), .Z(n3328) );
  XOR U2995 ( .A(y[1732]), .B(n3311), .Z(n3312) );
  XOR U2996 ( .A(y[1736]), .B(n3295), .Z(n3296) );
  XOR U2997 ( .A(y[1740]), .B(n3279), .Z(n3280) );
  XOR U2998 ( .A(y[1744]), .B(n3263), .Z(n3264) );
  XOR U2999 ( .A(y[1748]), .B(n3247), .Z(n3248) );
  XOR U3000 ( .A(y[1752]), .B(n3231), .Z(n3232) );
  XOR U3001 ( .A(y[1756]), .B(n3215), .Z(n3216) );
  XOR U3002 ( .A(y[1760]), .B(n3199), .Z(n3200) );
  XOR U3003 ( .A(y[1764]), .B(n3183), .Z(n3184) );
  XOR U3004 ( .A(y[1768]), .B(n3167), .Z(n3168) );
  XOR U3005 ( .A(y[1772]), .B(n3151), .Z(n3152) );
  XOR U3006 ( .A(y[1776]), .B(n3135), .Z(n3136) );
  XOR U3007 ( .A(y[1780]), .B(n3119), .Z(n3120) );
  XOR U3008 ( .A(y[1784]), .B(n3103), .Z(n3104) );
  XOR U3009 ( .A(y[1788]), .B(n3087), .Z(n3088) );
  XOR U3010 ( .A(y[1792]), .B(n3071), .Z(n3072) );
  XOR U3011 ( .A(y[1796]), .B(n3055), .Z(n3056) );
  XOR U3012 ( .A(y[1800]), .B(n3039), .Z(n3040) );
  XOR U3013 ( .A(y[1804]), .B(n3023), .Z(n3024) );
  XOR U3014 ( .A(y[1808]), .B(n3007), .Z(n3008) );
  XOR U3015 ( .A(y[1812]), .B(n2991), .Z(n2992) );
  XOR U3016 ( .A(y[1816]), .B(n2975), .Z(n2976) );
  XOR U3017 ( .A(y[1820]), .B(n2959), .Z(n2960) );
  XOR U3018 ( .A(y[1824]), .B(n2943), .Z(n2944) );
  XOR U3019 ( .A(y[1828]), .B(n2927), .Z(n2928) );
  XOR U3020 ( .A(y[1832]), .B(n2911), .Z(n2912) );
  XOR U3021 ( .A(y[1836]), .B(n2895), .Z(n2896) );
  XOR U3022 ( .A(y[1840]), .B(n2879), .Z(n2880) );
  XOR U3023 ( .A(y[1844]), .B(n2863), .Z(n2864) );
  XOR U3024 ( .A(y[1848]), .B(n2847), .Z(n2848) );
  XOR U3025 ( .A(y[1852]), .B(n2831), .Z(n2832) );
  XOR U3026 ( .A(y[1856]), .B(n2815), .Z(n2816) );
  XOR U3027 ( .A(y[1860]), .B(n2799), .Z(n2800) );
  XOR U3028 ( .A(y[1864]), .B(n2783), .Z(n2784) );
  XOR U3029 ( .A(y[1868]), .B(n2767), .Z(n2768) );
  XOR U3030 ( .A(y[1872]), .B(n2751), .Z(n2752) );
  XOR U3031 ( .A(y[1876]), .B(n2735), .Z(n2736) );
  XOR U3032 ( .A(y[1880]), .B(n2719), .Z(n2720) );
  XOR U3033 ( .A(y[1884]), .B(n2703), .Z(n2704) );
  XOR U3034 ( .A(y[1888]), .B(n2687), .Z(n2688) );
  XOR U3035 ( .A(y[1892]), .B(n2671), .Z(n2672) );
  XOR U3036 ( .A(y[1896]), .B(n2655), .Z(n2656) );
  XOR U3037 ( .A(y[1900]), .B(n2639), .Z(n2640) );
  XOR U3038 ( .A(y[1904]), .B(n2623), .Z(n2624) );
  XOR U3039 ( .A(y[1908]), .B(n2607), .Z(n2608) );
  XOR U3040 ( .A(y[1912]), .B(n2591), .Z(n2592) );
  XOR U3041 ( .A(y[1916]), .B(n2575), .Z(n2576) );
  XOR U3042 ( .A(y[1920]), .B(n2559), .Z(n2560) );
  XOR U3043 ( .A(y[1924]), .B(n2543), .Z(n2544) );
  XOR U3044 ( .A(y[1928]), .B(n2527), .Z(n2528) );
  XOR U3045 ( .A(y[1932]), .B(n2511), .Z(n2512) );
  XOR U3046 ( .A(y[1936]), .B(n2495), .Z(n2496) );
  XOR U3047 ( .A(y[1940]), .B(n2479), .Z(n2480) );
  XOR U3048 ( .A(y[1944]), .B(n2463), .Z(n2464) );
  XOR U3049 ( .A(y[1948]), .B(n2447), .Z(n2448) );
  XOR U3050 ( .A(y[1952]), .B(n2431), .Z(n2432) );
  XOR U3051 ( .A(y[1956]), .B(n2415), .Z(n2416) );
  XOR U3052 ( .A(y[1960]), .B(n2399), .Z(n2400) );
  XOR U3053 ( .A(y[1964]), .B(n2383), .Z(n2384) );
  XOR U3054 ( .A(y[1968]), .B(n2367), .Z(n2368) );
  XOR U3055 ( .A(y[1972]), .B(n2351), .Z(n2352) );
  XOR U3056 ( .A(y[1976]), .B(n2335), .Z(n2336) );
  XOR U3057 ( .A(y[1980]), .B(n2319), .Z(n2320) );
  XOR U3058 ( .A(y[1984]), .B(n2303), .Z(n2304) );
  XOR U3059 ( .A(y[1988]), .B(n2287), .Z(n2288) );
  XOR U3060 ( .A(y[1992]), .B(n2271), .Z(n2272) );
  XOR U3061 ( .A(y[1996]), .B(n2255), .Z(n2256) );
  XOR U3062 ( .A(y[2000]), .B(n2239), .Z(n2240) );
  XOR U3063 ( .A(y[2004]), .B(n2223), .Z(n2224) );
  XOR U3064 ( .A(y[2008]), .B(n2207), .Z(n2208) );
  XOR U3065 ( .A(y[2012]), .B(n2191), .Z(n2192) );
  XOR U3066 ( .A(y[2016]), .B(n2175), .Z(n2176) );
  XOR U3067 ( .A(y[2020]), .B(n2159), .Z(n2160) );
  XOR U3068 ( .A(y[2024]), .B(n2143), .Z(n2144) );
  XOR U3069 ( .A(y[2028]), .B(n2127), .Z(n2128) );
  XOR U3070 ( .A(y[2032]), .B(n2111), .Z(n2112) );
  XOR U3071 ( .A(y[2036]), .B(n2095), .Z(n2096) );
  XOR U3072 ( .A(y[2040]), .B(n2079), .Z(n2080) );
  XOR U3073 ( .A(y[2044]), .B(n2063), .Z(n2064) );
  XOR U3074 ( .A(y[5]), .B(n10219), .Z(n10220) );
  XOR U3075 ( .A(y[9]), .B(n10203), .Z(n10204) );
  XOR U3076 ( .A(y[13]), .B(n10187), .Z(n10188) );
  XOR U3077 ( .A(y[17]), .B(n10171), .Z(n10172) );
  XOR U3078 ( .A(y[21]), .B(n10155), .Z(n10156) );
  XOR U3079 ( .A(y[25]), .B(n10139), .Z(n10140) );
  XOR U3080 ( .A(y[29]), .B(n10123), .Z(n10124) );
  XOR U3081 ( .A(y[33]), .B(n10107), .Z(n10108) );
  XOR U3082 ( .A(y[37]), .B(n10091), .Z(n10092) );
  XOR U3083 ( .A(y[41]), .B(n10075), .Z(n10076) );
  XOR U3084 ( .A(y[45]), .B(n10059), .Z(n10060) );
  XOR U3085 ( .A(y[49]), .B(n10043), .Z(n10044) );
  XOR U3086 ( .A(y[53]), .B(n10027), .Z(n10028) );
  XOR U3087 ( .A(y[57]), .B(n10011), .Z(n10012) );
  XOR U3088 ( .A(y[61]), .B(n9995), .Z(n9996) );
  XOR U3089 ( .A(y[65]), .B(n9979), .Z(n9980) );
  XOR U3090 ( .A(y[69]), .B(n9963), .Z(n9964) );
  XOR U3091 ( .A(y[73]), .B(n9947), .Z(n9948) );
  XOR U3092 ( .A(y[77]), .B(n9931), .Z(n9932) );
  XOR U3093 ( .A(y[81]), .B(n9915), .Z(n9916) );
  XOR U3094 ( .A(y[85]), .B(n9899), .Z(n9900) );
  XOR U3095 ( .A(y[89]), .B(n9883), .Z(n9884) );
  XOR U3096 ( .A(y[93]), .B(n9867), .Z(n9868) );
  XOR U3097 ( .A(y[97]), .B(n9851), .Z(n9852) );
  XOR U3098 ( .A(y[101]), .B(n9835), .Z(n9836) );
  XOR U3099 ( .A(y[105]), .B(n9819), .Z(n9820) );
  XOR U3100 ( .A(y[109]), .B(n9803), .Z(n9804) );
  XOR U3101 ( .A(y[113]), .B(n9787), .Z(n9788) );
  XOR U3102 ( .A(y[117]), .B(n9771), .Z(n9772) );
  XOR U3103 ( .A(y[121]), .B(n9755), .Z(n9756) );
  XOR U3104 ( .A(y[125]), .B(n9739), .Z(n9740) );
  XOR U3105 ( .A(y[129]), .B(n9723), .Z(n9724) );
  XOR U3106 ( .A(y[133]), .B(n9707), .Z(n9708) );
  XOR U3107 ( .A(y[137]), .B(n9691), .Z(n9692) );
  XOR U3108 ( .A(y[141]), .B(n9675), .Z(n9676) );
  XOR U3109 ( .A(y[145]), .B(n9659), .Z(n9660) );
  XOR U3110 ( .A(y[149]), .B(n9643), .Z(n9644) );
  XOR U3111 ( .A(y[153]), .B(n9627), .Z(n9628) );
  XOR U3112 ( .A(y[157]), .B(n9611), .Z(n9612) );
  XOR U3113 ( .A(y[161]), .B(n9595), .Z(n9596) );
  XOR U3114 ( .A(y[165]), .B(n9579), .Z(n9580) );
  XOR U3115 ( .A(y[169]), .B(n9563), .Z(n9564) );
  XOR U3116 ( .A(y[173]), .B(n9547), .Z(n9548) );
  XOR U3117 ( .A(y[177]), .B(n9531), .Z(n9532) );
  XOR U3118 ( .A(y[181]), .B(n9515), .Z(n9516) );
  XOR U3119 ( .A(y[185]), .B(n9499), .Z(n9500) );
  XOR U3120 ( .A(y[189]), .B(n9483), .Z(n9484) );
  XOR U3121 ( .A(y[193]), .B(n9467), .Z(n9468) );
  XOR U3122 ( .A(y[197]), .B(n9451), .Z(n9452) );
  XOR U3123 ( .A(y[201]), .B(n9435), .Z(n9436) );
  XOR U3124 ( .A(y[205]), .B(n9419), .Z(n9420) );
  XOR U3125 ( .A(y[209]), .B(n9403), .Z(n9404) );
  XOR U3126 ( .A(y[213]), .B(n9387), .Z(n9388) );
  XOR U3127 ( .A(y[217]), .B(n9371), .Z(n9372) );
  XOR U3128 ( .A(y[221]), .B(n9355), .Z(n9356) );
  XOR U3129 ( .A(y[225]), .B(n9339), .Z(n9340) );
  XOR U3130 ( .A(y[229]), .B(n9323), .Z(n9324) );
  XOR U3131 ( .A(y[233]), .B(n9307), .Z(n9308) );
  XOR U3132 ( .A(y[237]), .B(n9291), .Z(n9292) );
  XOR U3133 ( .A(y[241]), .B(n9275), .Z(n9276) );
  XOR U3134 ( .A(y[245]), .B(n9259), .Z(n9260) );
  XOR U3135 ( .A(y[249]), .B(n9243), .Z(n9244) );
  XOR U3136 ( .A(y[253]), .B(n9227), .Z(n9228) );
  XOR U3137 ( .A(y[257]), .B(n9211), .Z(n9212) );
  XOR U3138 ( .A(y[261]), .B(n9195), .Z(n9196) );
  XOR U3139 ( .A(y[265]), .B(n9179), .Z(n9180) );
  XOR U3140 ( .A(y[269]), .B(n9163), .Z(n9164) );
  XOR U3141 ( .A(y[273]), .B(n9147), .Z(n9148) );
  XOR U3142 ( .A(y[277]), .B(n9131), .Z(n9132) );
  XOR U3143 ( .A(y[281]), .B(n9115), .Z(n9116) );
  XOR U3144 ( .A(y[285]), .B(n9099), .Z(n9100) );
  XOR U3145 ( .A(y[289]), .B(n9083), .Z(n9084) );
  XOR U3146 ( .A(y[293]), .B(n9067), .Z(n9068) );
  XOR U3147 ( .A(y[297]), .B(n9051), .Z(n9052) );
  XOR U3148 ( .A(y[301]), .B(n9035), .Z(n9036) );
  XOR U3149 ( .A(y[305]), .B(n9019), .Z(n9020) );
  XOR U3150 ( .A(y[309]), .B(n9003), .Z(n9004) );
  XOR U3151 ( .A(y[313]), .B(n8987), .Z(n8988) );
  XOR U3152 ( .A(y[317]), .B(n8971), .Z(n8972) );
  XOR U3153 ( .A(y[321]), .B(n8955), .Z(n8956) );
  XOR U3154 ( .A(y[325]), .B(n8939), .Z(n8940) );
  XOR U3155 ( .A(y[329]), .B(n8923), .Z(n8924) );
  XOR U3156 ( .A(y[333]), .B(n8907), .Z(n8908) );
  XOR U3157 ( .A(y[337]), .B(n8891), .Z(n8892) );
  XOR U3158 ( .A(y[341]), .B(n8875), .Z(n8876) );
  XOR U3159 ( .A(y[345]), .B(n8859), .Z(n8860) );
  XOR U3160 ( .A(y[349]), .B(n8843), .Z(n8844) );
  XOR U3161 ( .A(y[353]), .B(n8827), .Z(n8828) );
  XOR U3162 ( .A(y[357]), .B(n8811), .Z(n8812) );
  XOR U3163 ( .A(y[361]), .B(n8795), .Z(n8796) );
  XOR U3164 ( .A(y[365]), .B(n8779), .Z(n8780) );
  XOR U3165 ( .A(y[369]), .B(n8763), .Z(n8764) );
  XOR U3166 ( .A(y[373]), .B(n8747), .Z(n8748) );
  XOR U3167 ( .A(y[377]), .B(n8731), .Z(n8732) );
  XOR U3168 ( .A(y[381]), .B(n8715), .Z(n8716) );
  XOR U3169 ( .A(y[385]), .B(n8699), .Z(n8700) );
  XOR U3170 ( .A(y[389]), .B(n8683), .Z(n8684) );
  XOR U3171 ( .A(y[393]), .B(n8667), .Z(n8668) );
  XOR U3172 ( .A(y[397]), .B(n8651), .Z(n8652) );
  XOR U3173 ( .A(y[401]), .B(n8635), .Z(n8636) );
  XOR U3174 ( .A(y[405]), .B(n8619), .Z(n8620) );
  XOR U3175 ( .A(y[409]), .B(n8603), .Z(n8604) );
  XOR U3176 ( .A(y[413]), .B(n8587), .Z(n8588) );
  XOR U3177 ( .A(y[417]), .B(n8571), .Z(n8572) );
  XOR U3178 ( .A(y[421]), .B(n8555), .Z(n8556) );
  XOR U3179 ( .A(y[425]), .B(n8539), .Z(n8540) );
  XOR U3180 ( .A(y[429]), .B(n8523), .Z(n8524) );
  XOR U3181 ( .A(y[433]), .B(n8507), .Z(n8508) );
  XOR U3182 ( .A(y[437]), .B(n8491), .Z(n8492) );
  XOR U3183 ( .A(y[441]), .B(n8475), .Z(n8476) );
  XOR U3184 ( .A(y[445]), .B(n8459), .Z(n8460) );
  XOR U3185 ( .A(y[449]), .B(n8443), .Z(n8444) );
  XOR U3186 ( .A(y[453]), .B(n8427), .Z(n8428) );
  XOR U3187 ( .A(y[457]), .B(n8411), .Z(n8412) );
  XOR U3188 ( .A(y[461]), .B(n8395), .Z(n8396) );
  XOR U3189 ( .A(y[465]), .B(n8379), .Z(n8380) );
  XOR U3190 ( .A(y[469]), .B(n8363), .Z(n8364) );
  XOR U3191 ( .A(y[473]), .B(n8347), .Z(n8348) );
  XOR U3192 ( .A(y[477]), .B(n8331), .Z(n8332) );
  XOR U3193 ( .A(y[481]), .B(n8315), .Z(n8316) );
  XOR U3194 ( .A(y[485]), .B(n8299), .Z(n8300) );
  XOR U3195 ( .A(y[489]), .B(n8283), .Z(n8284) );
  XOR U3196 ( .A(y[493]), .B(n8267), .Z(n8268) );
  XOR U3197 ( .A(y[497]), .B(n8251), .Z(n8252) );
  XOR U3198 ( .A(y[501]), .B(n8235), .Z(n8236) );
  XOR U3199 ( .A(y[505]), .B(n8219), .Z(n8220) );
  XOR U3200 ( .A(y[509]), .B(n8203), .Z(n8204) );
  XOR U3201 ( .A(y[513]), .B(n8187), .Z(n8188) );
  XOR U3202 ( .A(y[517]), .B(n8171), .Z(n8172) );
  XOR U3203 ( .A(y[521]), .B(n8155), .Z(n8156) );
  XOR U3204 ( .A(y[525]), .B(n8139), .Z(n8140) );
  XOR U3205 ( .A(y[529]), .B(n8123), .Z(n8124) );
  XOR U3206 ( .A(y[533]), .B(n8107), .Z(n8108) );
  XOR U3207 ( .A(y[537]), .B(n8091), .Z(n8092) );
  XOR U3208 ( .A(y[541]), .B(n8075), .Z(n8076) );
  XOR U3209 ( .A(y[545]), .B(n8059), .Z(n8060) );
  XOR U3210 ( .A(y[549]), .B(n8043), .Z(n8044) );
  XOR U3211 ( .A(y[553]), .B(n8027), .Z(n8028) );
  XOR U3212 ( .A(y[557]), .B(n8011), .Z(n8012) );
  XOR U3213 ( .A(y[561]), .B(n7995), .Z(n7996) );
  XOR U3214 ( .A(y[565]), .B(n7979), .Z(n7980) );
  XOR U3215 ( .A(y[569]), .B(n7963), .Z(n7964) );
  XOR U3216 ( .A(y[573]), .B(n7947), .Z(n7948) );
  XOR U3217 ( .A(y[577]), .B(n7931), .Z(n7932) );
  XOR U3218 ( .A(y[581]), .B(n7915), .Z(n7916) );
  XOR U3219 ( .A(y[585]), .B(n7899), .Z(n7900) );
  XOR U3220 ( .A(y[589]), .B(n7883), .Z(n7884) );
  XOR U3221 ( .A(y[593]), .B(n7867), .Z(n7868) );
  XOR U3222 ( .A(y[597]), .B(n7851), .Z(n7852) );
  XOR U3223 ( .A(y[601]), .B(n7835), .Z(n7836) );
  XOR U3224 ( .A(y[605]), .B(n7819), .Z(n7820) );
  XOR U3225 ( .A(y[609]), .B(n7803), .Z(n7804) );
  XOR U3226 ( .A(y[613]), .B(n7787), .Z(n7788) );
  XOR U3227 ( .A(y[617]), .B(n7771), .Z(n7772) );
  XOR U3228 ( .A(y[621]), .B(n7755), .Z(n7756) );
  XOR U3229 ( .A(y[625]), .B(n7739), .Z(n7740) );
  XOR U3230 ( .A(y[629]), .B(n7723), .Z(n7724) );
  XOR U3231 ( .A(y[633]), .B(n7707), .Z(n7708) );
  XOR U3232 ( .A(y[637]), .B(n7691), .Z(n7692) );
  XOR U3233 ( .A(y[641]), .B(n7675), .Z(n7676) );
  XOR U3234 ( .A(y[645]), .B(n7659), .Z(n7660) );
  XOR U3235 ( .A(y[649]), .B(n7643), .Z(n7644) );
  XOR U3236 ( .A(y[653]), .B(n7627), .Z(n7628) );
  XOR U3237 ( .A(y[657]), .B(n7611), .Z(n7612) );
  XOR U3238 ( .A(y[661]), .B(n7595), .Z(n7596) );
  XOR U3239 ( .A(y[665]), .B(n7579), .Z(n7580) );
  XOR U3240 ( .A(y[669]), .B(n7563), .Z(n7564) );
  XOR U3241 ( .A(y[673]), .B(n7547), .Z(n7548) );
  XOR U3242 ( .A(y[677]), .B(n7531), .Z(n7532) );
  XOR U3243 ( .A(y[681]), .B(n7515), .Z(n7516) );
  XOR U3244 ( .A(y[685]), .B(n7499), .Z(n7500) );
  XOR U3245 ( .A(y[689]), .B(n7483), .Z(n7484) );
  XOR U3246 ( .A(y[693]), .B(n7467), .Z(n7468) );
  XOR U3247 ( .A(y[697]), .B(n7451), .Z(n7452) );
  XOR U3248 ( .A(y[701]), .B(n7435), .Z(n7436) );
  XOR U3249 ( .A(y[705]), .B(n7419), .Z(n7420) );
  XOR U3250 ( .A(y[709]), .B(n7403), .Z(n7404) );
  XOR U3251 ( .A(y[713]), .B(n7387), .Z(n7388) );
  XOR U3252 ( .A(y[717]), .B(n7371), .Z(n7372) );
  XOR U3253 ( .A(y[721]), .B(n7355), .Z(n7356) );
  XOR U3254 ( .A(y[725]), .B(n7339), .Z(n7340) );
  XOR U3255 ( .A(y[729]), .B(n7323), .Z(n7324) );
  XOR U3256 ( .A(y[733]), .B(n7307), .Z(n7308) );
  XOR U3257 ( .A(y[737]), .B(n7291), .Z(n7292) );
  XOR U3258 ( .A(y[741]), .B(n7275), .Z(n7276) );
  XOR U3259 ( .A(y[745]), .B(n7259), .Z(n7260) );
  XOR U3260 ( .A(y[749]), .B(n7243), .Z(n7244) );
  XOR U3261 ( .A(y[753]), .B(n7227), .Z(n7228) );
  XOR U3262 ( .A(y[757]), .B(n7211), .Z(n7212) );
  XOR U3263 ( .A(y[761]), .B(n7195), .Z(n7196) );
  XOR U3264 ( .A(y[765]), .B(n7179), .Z(n7180) );
  XOR U3265 ( .A(y[769]), .B(n7163), .Z(n7164) );
  XOR U3266 ( .A(y[773]), .B(n7147), .Z(n7148) );
  XOR U3267 ( .A(y[777]), .B(n7131), .Z(n7132) );
  XOR U3268 ( .A(y[781]), .B(n7115), .Z(n7116) );
  XOR U3269 ( .A(y[785]), .B(n7099), .Z(n7100) );
  XOR U3270 ( .A(y[789]), .B(n7083), .Z(n7084) );
  XOR U3271 ( .A(y[793]), .B(n7067), .Z(n7068) );
  XOR U3272 ( .A(y[797]), .B(n7051), .Z(n7052) );
  XOR U3273 ( .A(y[801]), .B(n7035), .Z(n7036) );
  XOR U3274 ( .A(y[805]), .B(n7019), .Z(n7020) );
  XOR U3275 ( .A(y[809]), .B(n7003), .Z(n7004) );
  XOR U3276 ( .A(y[813]), .B(n6987), .Z(n6988) );
  XOR U3277 ( .A(y[817]), .B(n6971), .Z(n6972) );
  XOR U3278 ( .A(y[821]), .B(n6955), .Z(n6956) );
  XOR U3279 ( .A(y[825]), .B(n6939), .Z(n6940) );
  XOR U3280 ( .A(y[829]), .B(n6923), .Z(n6924) );
  XOR U3281 ( .A(y[833]), .B(n6907), .Z(n6908) );
  XOR U3282 ( .A(y[837]), .B(n6891), .Z(n6892) );
  XOR U3283 ( .A(y[841]), .B(n6875), .Z(n6876) );
  XOR U3284 ( .A(y[845]), .B(n6859), .Z(n6860) );
  XOR U3285 ( .A(y[849]), .B(n6843), .Z(n6844) );
  XOR U3286 ( .A(y[853]), .B(n6827), .Z(n6828) );
  XOR U3287 ( .A(y[857]), .B(n6811), .Z(n6812) );
  XOR U3288 ( .A(y[861]), .B(n6795), .Z(n6796) );
  XOR U3289 ( .A(y[865]), .B(n6779), .Z(n6780) );
  XOR U3290 ( .A(y[869]), .B(n6763), .Z(n6764) );
  XOR U3291 ( .A(y[873]), .B(n6747), .Z(n6748) );
  XOR U3292 ( .A(y[877]), .B(n6731), .Z(n6732) );
  XOR U3293 ( .A(y[881]), .B(n6715), .Z(n6716) );
  XOR U3294 ( .A(y[885]), .B(n6699), .Z(n6700) );
  XOR U3295 ( .A(y[889]), .B(n6683), .Z(n6684) );
  XOR U3296 ( .A(y[893]), .B(n6667), .Z(n6668) );
  XOR U3297 ( .A(y[897]), .B(n6651), .Z(n6652) );
  XOR U3298 ( .A(y[901]), .B(n6635), .Z(n6636) );
  XOR U3299 ( .A(y[905]), .B(n6619), .Z(n6620) );
  XOR U3300 ( .A(y[909]), .B(n6603), .Z(n6604) );
  XOR U3301 ( .A(y[913]), .B(n6587), .Z(n6588) );
  XOR U3302 ( .A(y[917]), .B(n6571), .Z(n6572) );
  XOR U3303 ( .A(y[921]), .B(n6555), .Z(n6556) );
  XOR U3304 ( .A(y[925]), .B(n6539), .Z(n6540) );
  XOR U3305 ( .A(y[929]), .B(n6523), .Z(n6524) );
  XOR U3306 ( .A(y[933]), .B(n6507), .Z(n6508) );
  XOR U3307 ( .A(y[937]), .B(n6491), .Z(n6492) );
  XOR U3308 ( .A(y[941]), .B(n6475), .Z(n6476) );
  XOR U3309 ( .A(y[945]), .B(n6459), .Z(n6460) );
  XOR U3310 ( .A(y[949]), .B(n6443), .Z(n6444) );
  XOR U3311 ( .A(y[953]), .B(n6427), .Z(n6428) );
  XOR U3312 ( .A(y[957]), .B(n6411), .Z(n6412) );
  XOR U3313 ( .A(y[961]), .B(n6395), .Z(n6396) );
  XOR U3314 ( .A(y[965]), .B(n6379), .Z(n6380) );
  XOR U3315 ( .A(y[969]), .B(n6363), .Z(n6364) );
  XOR U3316 ( .A(y[973]), .B(n6347), .Z(n6348) );
  XOR U3317 ( .A(y[977]), .B(n6331), .Z(n6332) );
  XOR U3318 ( .A(y[981]), .B(n6315), .Z(n6316) );
  XOR U3319 ( .A(y[985]), .B(n6299), .Z(n6300) );
  XOR U3320 ( .A(y[989]), .B(n6283), .Z(n6284) );
  XOR U3321 ( .A(y[993]), .B(n6267), .Z(n6268) );
  XOR U3322 ( .A(y[997]), .B(n6251), .Z(n6252) );
  XOR U3323 ( .A(y[1001]), .B(n6235), .Z(n6236) );
  XOR U3324 ( .A(y[1005]), .B(n6219), .Z(n6220) );
  XOR U3325 ( .A(y[1009]), .B(n6203), .Z(n6204) );
  XOR U3326 ( .A(y[1013]), .B(n6187), .Z(n6188) );
  XOR U3327 ( .A(y[1017]), .B(n6171), .Z(n6172) );
  XOR U3328 ( .A(y[1021]), .B(n6155), .Z(n6156) );
  XOR U3329 ( .A(y[1025]), .B(n6139), .Z(n6140) );
  XOR U3330 ( .A(y[1029]), .B(n6123), .Z(n6124) );
  XOR U3331 ( .A(y[1033]), .B(n6107), .Z(n6108) );
  XOR U3332 ( .A(y[1037]), .B(n6091), .Z(n6092) );
  XOR U3333 ( .A(y[1041]), .B(n6075), .Z(n6076) );
  XOR U3334 ( .A(y[1045]), .B(n6059), .Z(n6060) );
  XOR U3335 ( .A(y[1049]), .B(n6043), .Z(n6044) );
  XOR U3336 ( .A(y[1053]), .B(n6027), .Z(n6028) );
  XOR U3337 ( .A(y[1057]), .B(n6011), .Z(n6012) );
  XOR U3338 ( .A(y[1061]), .B(n5995), .Z(n5996) );
  XOR U3339 ( .A(y[1065]), .B(n5979), .Z(n5980) );
  XOR U3340 ( .A(y[1069]), .B(n5963), .Z(n5964) );
  XOR U3341 ( .A(y[1073]), .B(n5947), .Z(n5948) );
  XOR U3342 ( .A(y[1077]), .B(n5931), .Z(n5932) );
  XOR U3343 ( .A(y[1081]), .B(n5915), .Z(n5916) );
  XOR U3344 ( .A(y[1085]), .B(n5899), .Z(n5900) );
  XOR U3345 ( .A(y[1089]), .B(n5883), .Z(n5884) );
  XOR U3346 ( .A(y[1093]), .B(n5867), .Z(n5868) );
  XOR U3347 ( .A(y[1097]), .B(n5851), .Z(n5852) );
  XOR U3348 ( .A(y[1101]), .B(n5835), .Z(n5836) );
  XOR U3349 ( .A(y[1105]), .B(n5819), .Z(n5820) );
  XOR U3350 ( .A(y[1109]), .B(n5803), .Z(n5804) );
  XOR U3351 ( .A(y[1113]), .B(n5787), .Z(n5788) );
  XOR U3352 ( .A(y[1117]), .B(n5771), .Z(n5772) );
  XOR U3353 ( .A(y[1121]), .B(n5755), .Z(n5756) );
  XOR U3354 ( .A(y[1125]), .B(n5739), .Z(n5740) );
  XOR U3355 ( .A(y[1129]), .B(n5723), .Z(n5724) );
  XOR U3356 ( .A(y[1133]), .B(n5707), .Z(n5708) );
  XOR U3357 ( .A(y[1137]), .B(n5691), .Z(n5692) );
  XOR U3358 ( .A(y[1141]), .B(n5675), .Z(n5676) );
  XOR U3359 ( .A(y[1145]), .B(n5659), .Z(n5660) );
  XOR U3360 ( .A(y[1149]), .B(n5643), .Z(n5644) );
  XOR U3361 ( .A(y[1153]), .B(n5627), .Z(n5628) );
  XOR U3362 ( .A(y[1157]), .B(n5611), .Z(n5612) );
  XOR U3363 ( .A(y[1161]), .B(n5595), .Z(n5596) );
  XOR U3364 ( .A(y[1165]), .B(n5579), .Z(n5580) );
  XOR U3365 ( .A(y[1169]), .B(n5563), .Z(n5564) );
  XOR U3366 ( .A(y[1173]), .B(n5547), .Z(n5548) );
  XOR U3367 ( .A(y[1177]), .B(n5531), .Z(n5532) );
  XOR U3368 ( .A(y[1181]), .B(n5515), .Z(n5516) );
  XOR U3369 ( .A(y[1185]), .B(n5499), .Z(n5500) );
  XOR U3370 ( .A(y[1189]), .B(n5483), .Z(n5484) );
  XOR U3371 ( .A(y[1193]), .B(n5467), .Z(n5468) );
  XOR U3372 ( .A(y[1197]), .B(n5451), .Z(n5452) );
  XOR U3373 ( .A(y[1201]), .B(n5435), .Z(n5436) );
  XOR U3374 ( .A(y[1205]), .B(n5419), .Z(n5420) );
  XOR U3375 ( .A(y[1209]), .B(n5403), .Z(n5404) );
  XOR U3376 ( .A(y[1213]), .B(n5387), .Z(n5388) );
  XOR U3377 ( .A(y[1217]), .B(n5371), .Z(n5372) );
  XOR U3378 ( .A(y[1221]), .B(n5355), .Z(n5356) );
  XOR U3379 ( .A(y[1225]), .B(n5339), .Z(n5340) );
  XOR U3380 ( .A(y[1229]), .B(n5323), .Z(n5324) );
  XOR U3381 ( .A(y[1233]), .B(n5307), .Z(n5308) );
  XOR U3382 ( .A(y[1237]), .B(n5291), .Z(n5292) );
  XOR U3383 ( .A(y[1241]), .B(n5275), .Z(n5276) );
  XOR U3384 ( .A(y[1245]), .B(n5259), .Z(n5260) );
  XOR U3385 ( .A(y[1249]), .B(n5243), .Z(n5244) );
  XOR U3386 ( .A(y[1253]), .B(n5227), .Z(n5228) );
  XOR U3387 ( .A(y[1257]), .B(n5211), .Z(n5212) );
  XOR U3388 ( .A(y[1261]), .B(n5195), .Z(n5196) );
  XOR U3389 ( .A(y[1265]), .B(n5179), .Z(n5180) );
  XOR U3390 ( .A(y[1269]), .B(n5163), .Z(n5164) );
  XOR U3391 ( .A(y[1273]), .B(n5147), .Z(n5148) );
  XOR U3392 ( .A(y[1277]), .B(n5131), .Z(n5132) );
  XOR U3393 ( .A(y[1281]), .B(n5115), .Z(n5116) );
  XOR U3394 ( .A(y[1285]), .B(n5099), .Z(n5100) );
  XOR U3395 ( .A(y[1289]), .B(n5083), .Z(n5084) );
  XOR U3396 ( .A(y[1293]), .B(n5067), .Z(n5068) );
  XOR U3397 ( .A(y[1297]), .B(n5051), .Z(n5052) );
  XOR U3398 ( .A(y[1301]), .B(n5035), .Z(n5036) );
  XOR U3399 ( .A(y[1305]), .B(n5019), .Z(n5020) );
  XOR U3400 ( .A(y[1309]), .B(n5003), .Z(n5004) );
  XOR U3401 ( .A(y[1313]), .B(n4987), .Z(n4988) );
  XOR U3402 ( .A(y[1317]), .B(n4971), .Z(n4972) );
  XOR U3403 ( .A(y[1321]), .B(n4955), .Z(n4956) );
  XOR U3404 ( .A(y[1325]), .B(n4939), .Z(n4940) );
  XOR U3405 ( .A(y[1329]), .B(n4923), .Z(n4924) );
  XOR U3406 ( .A(y[1333]), .B(n4907), .Z(n4908) );
  XOR U3407 ( .A(y[1337]), .B(n4891), .Z(n4892) );
  XOR U3408 ( .A(y[1341]), .B(n4875), .Z(n4876) );
  XOR U3409 ( .A(y[1345]), .B(n4859), .Z(n4860) );
  XOR U3410 ( .A(y[1349]), .B(n4843), .Z(n4844) );
  XOR U3411 ( .A(y[1353]), .B(n4827), .Z(n4828) );
  XOR U3412 ( .A(y[1357]), .B(n4811), .Z(n4812) );
  XOR U3413 ( .A(y[1361]), .B(n4795), .Z(n4796) );
  XOR U3414 ( .A(y[1365]), .B(n4779), .Z(n4780) );
  XOR U3415 ( .A(y[1369]), .B(n4763), .Z(n4764) );
  XOR U3416 ( .A(y[1373]), .B(n4747), .Z(n4748) );
  XOR U3417 ( .A(y[1377]), .B(n4731), .Z(n4732) );
  XOR U3418 ( .A(y[1381]), .B(n4715), .Z(n4716) );
  XOR U3419 ( .A(y[1385]), .B(n4699), .Z(n4700) );
  XOR U3420 ( .A(y[1389]), .B(n4683), .Z(n4684) );
  XOR U3421 ( .A(y[1393]), .B(n4667), .Z(n4668) );
  XOR U3422 ( .A(y[1397]), .B(n4651), .Z(n4652) );
  XOR U3423 ( .A(y[1401]), .B(n4635), .Z(n4636) );
  XOR U3424 ( .A(y[1405]), .B(n4619), .Z(n4620) );
  XOR U3425 ( .A(y[1409]), .B(n4603), .Z(n4604) );
  XOR U3426 ( .A(y[1413]), .B(n4587), .Z(n4588) );
  XOR U3427 ( .A(y[1417]), .B(n4571), .Z(n4572) );
  XOR U3428 ( .A(y[1421]), .B(n4555), .Z(n4556) );
  XOR U3429 ( .A(y[1425]), .B(n4539), .Z(n4540) );
  XOR U3430 ( .A(y[1429]), .B(n4523), .Z(n4524) );
  XOR U3431 ( .A(y[1433]), .B(n4507), .Z(n4508) );
  XOR U3432 ( .A(y[1437]), .B(n4491), .Z(n4492) );
  XOR U3433 ( .A(y[1441]), .B(n4475), .Z(n4476) );
  XOR U3434 ( .A(y[1445]), .B(n4459), .Z(n4460) );
  XOR U3435 ( .A(y[1449]), .B(n4443), .Z(n4444) );
  XOR U3436 ( .A(y[1453]), .B(n4427), .Z(n4428) );
  XOR U3437 ( .A(y[1457]), .B(n4411), .Z(n4412) );
  XOR U3438 ( .A(y[1461]), .B(n4395), .Z(n4396) );
  XOR U3439 ( .A(y[1465]), .B(n4379), .Z(n4380) );
  XOR U3440 ( .A(y[1469]), .B(n4363), .Z(n4364) );
  XOR U3441 ( .A(y[1473]), .B(n4347), .Z(n4348) );
  XOR U3442 ( .A(y[1477]), .B(n4331), .Z(n4332) );
  XOR U3443 ( .A(y[1481]), .B(n4315), .Z(n4316) );
  XOR U3444 ( .A(y[1485]), .B(n4299), .Z(n4300) );
  XOR U3445 ( .A(y[1489]), .B(n4283), .Z(n4284) );
  XOR U3446 ( .A(y[1493]), .B(n4267), .Z(n4268) );
  XOR U3447 ( .A(y[1497]), .B(n4251), .Z(n4252) );
  XOR U3448 ( .A(y[1501]), .B(n4235), .Z(n4236) );
  XOR U3449 ( .A(y[1505]), .B(n4219), .Z(n4220) );
  XOR U3450 ( .A(y[1509]), .B(n4203), .Z(n4204) );
  XOR U3451 ( .A(y[1513]), .B(n4187), .Z(n4188) );
  XOR U3452 ( .A(y[1517]), .B(n4171), .Z(n4172) );
  XOR U3453 ( .A(y[1521]), .B(n4155), .Z(n4156) );
  XOR U3454 ( .A(y[1525]), .B(n4139), .Z(n4140) );
  XOR U3455 ( .A(y[1529]), .B(n4123), .Z(n4124) );
  XOR U3456 ( .A(y[1533]), .B(n4107), .Z(n4108) );
  XOR U3457 ( .A(y[1537]), .B(n4091), .Z(n4092) );
  XOR U3458 ( .A(y[1541]), .B(n4075), .Z(n4076) );
  XOR U3459 ( .A(y[1545]), .B(n4059), .Z(n4060) );
  XOR U3460 ( .A(y[1549]), .B(n4043), .Z(n4044) );
  XOR U3461 ( .A(y[1553]), .B(n4027), .Z(n4028) );
  XOR U3462 ( .A(y[1557]), .B(n4011), .Z(n4012) );
  XOR U3463 ( .A(y[1561]), .B(n3995), .Z(n3996) );
  XOR U3464 ( .A(y[1565]), .B(n3979), .Z(n3980) );
  XOR U3465 ( .A(y[1569]), .B(n3963), .Z(n3964) );
  XOR U3466 ( .A(y[1573]), .B(n3947), .Z(n3948) );
  XOR U3467 ( .A(y[1577]), .B(n3931), .Z(n3932) );
  XOR U3468 ( .A(y[1581]), .B(n3915), .Z(n3916) );
  XOR U3469 ( .A(y[1585]), .B(n3899), .Z(n3900) );
  XOR U3470 ( .A(y[1589]), .B(n3883), .Z(n3884) );
  XOR U3471 ( .A(y[1593]), .B(n3867), .Z(n3868) );
  XOR U3472 ( .A(y[1597]), .B(n3851), .Z(n3852) );
  XOR U3473 ( .A(y[1601]), .B(n3835), .Z(n3836) );
  XOR U3474 ( .A(y[1605]), .B(n3819), .Z(n3820) );
  XOR U3475 ( .A(y[1609]), .B(n3803), .Z(n3804) );
  XOR U3476 ( .A(y[1613]), .B(n3787), .Z(n3788) );
  XOR U3477 ( .A(y[1617]), .B(n3771), .Z(n3772) );
  XOR U3478 ( .A(y[1621]), .B(n3755), .Z(n3756) );
  XOR U3479 ( .A(y[1625]), .B(n3739), .Z(n3740) );
  XOR U3480 ( .A(y[1629]), .B(n3723), .Z(n3724) );
  XOR U3481 ( .A(y[1633]), .B(n3707), .Z(n3708) );
  XOR U3482 ( .A(y[1637]), .B(n3691), .Z(n3692) );
  XOR U3483 ( .A(y[1641]), .B(n3675), .Z(n3676) );
  XOR U3484 ( .A(y[1645]), .B(n3659), .Z(n3660) );
  XOR U3485 ( .A(y[1649]), .B(n3643), .Z(n3644) );
  XOR U3486 ( .A(y[1653]), .B(n3627), .Z(n3628) );
  XOR U3487 ( .A(y[1657]), .B(n3611), .Z(n3612) );
  XOR U3488 ( .A(y[1661]), .B(n3595), .Z(n3596) );
  XOR U3489 ( .A(y[1665]), .B(n3579), .Z(n3580) );
  XOR U3490 ( .A(y[1669]), .B(n3563), .Z(n3564) );
  XOR U3491 ( .A(y[1673]), .B(n3547), .Z(n3548) );
  XOR U3492 ( .A(y[1677]), .B(n3531), .Z(n3532) );
  XOR U3493 ( .A(y[1681]), .B(n3515), .Z(n3516) );
  XOR U3494 ( .A(y[1685]), .B(n3499), .Z(n3500) );
  XOR U3495 ( .A(y[1689]), .B(n3483), .Z(n3484) );
  XOR U3496 ( .A(y[1693]), .B(n3467), .Z(n3468) );
  XOR U3497 ( .A(y[1697]), .B(n3451), .Z(n3452) );
  XOR U3498 ( .A(y[1701]), .B(n3435), .Z(n3436) );
  XOR U3499 ( .A(y[1705]), .B(n3419), .Z(n3420) );
  XOR U3500 ( .A(y[1709]), .B(n3403), .Z(n3404) );
  XOR U3501 ( .A(y[1713]), .B(n3387), .Z(n3388) );
  XOR U3502 ( .A(y[1717]), .B(n3371), .Z(n3372) );
  XOR U3503 ( .A(y[1721]), .B(n3355), .Z(n3356) );
  XOR U3504 ( .A(y[1725]), .B(n3339), .Z(n3340) );
  XOR U3505 ( .A(y[1729]), .B(n3323), .Z(n3324) );
  XOR U3506 ( .A(y[1733]), .B(n3307), .Z(n3308) );
  XOR U3507 ( .A(y[1737]), .B(n3291), .Z(n3292) );
  XOR U3508 ( .A(y[1741]), .B(n3275), .Z(n3276) );
  XOR U3509 ( .A(y[1745]), .B(n3259), .Z(n3260) );
  XOR U3510 ( .A(y[1749]), .B(n3243), .Z(n3244) );
  XOR U3511 ( .A(y[1753]), .B(n3227), .Z(n3228) );
  XOR U3512 ( .A(y[1757]), .B(n3211), .Z(n3212) );
  XOR U3513 ( .A(y[1761]), .B(n3195), .Z(n3196) );
  XOR U3514 ( .A(y[1765]), .B(n3179), .Z(n3180) );
  XOR U3515 ( .A(y[1769]), .B(n3163), .Z(n3164) );
  XOR U3516 ( .A(y[1773]), .B(n3147), .Z(n3148) );
  XOR U3517 ( .A(y[1777]), .B(n3131), .Z(n3132) );
  XOR U3518 ( .A(y[1781]), .B(n3115), .Z(n3116) );
  XOR U3519 ( .A(y[1785]), .B(n3099), .Z(n3100) );
  XOR U3520 ( .A(y[1789]), .B(n3083), .Z(n3084) );
  XOR U3521 ( .A(y[1793]), .B(n3067), .Z(n3068) );
  XOR U3522 ( .A(y[1797]), .B(n3051), .Z(n3052) );
  XOR U3523 ( .A(y[1801]), .B(n3035), .Z(n3036) );
  XOR U3524 ( .A(y[1805]), .B(n3019), .Z(n3020) );
  XOR U3525 ( .A(y[1809]), .B(n3003), .Z(n3004) );
  XOR U3526 ( .A(y[1813]), .B(n2987), .Z(n2988) );
  XOR U3527 ( .A(y[1817]), .B(n2971), .Z(n2972) );
  XOR U3528 ( .A(y[1821]), .B(n2955), .Z(n2956) );
  XOR U3529 ( .A(y[1825]), .B(n2939), .Z(n2940) );
  XOR U3530 ( .A(y[1829]), .B(n2923), .Z(n2924) );
  XOR U3531 ( .A(y[1833]), .B(n2907), .Z(n2908) );
  XOR U3532 ( .A(y[1837]), .B(n2891), .Z(n2892) );
  XOR U3533 ( .A(y[1841]), .B(n2875), .Z(n2876) );
  XOR U3534 ( .A(y[1845]), .B(n2859), .Z(n2860) );
  XOR U3535 ( .A(y[1849]), .B(n2843), .Z(n2844) );
  XOR U3536 ( .A(y[1853]), .B(n2827), .Z(n2828) );
  XOR U3537 ( .A(y[1857]), .B(n2811), .Z(n2812) );
  XOR U3538 ( .A(y[1861]), .B(n2795), .Z(n2796) );
  XOR U3539 ( .A(y[1865]), .B(n2779), .Z(n2780) );
  XOR U3540 ( .A(y[1869]), .B(n2763), .Z(n2764) );
  XOR U3541 ( .A(y[1873]), .B(n2747), .Z(n2748) );
  XOR U3542 ( .A(y[1877]), .B(n2731), .Z(n2732) );
  XOR U3543 ( .A(y[1881]), .B(n2715), .Z(n2716) );
  XOR U3544 ( .A(y[1885]), .B(n2699), .Z(n2700) );
  XOR U3545 ( .A(y[1889]), .B(n2683), .Z(n2684) );
  XOR U3546 ( .A(y[1893]), .B(n2667), .Z(n2668) );
  XOR U3547 ( .A(y[1897]), .B(n2651), .Z(n2652) );
  XOR U3548 ( .A(y[1901]), .B(n2635), .Z(n2636) );
  XOR U3549 ( .A(y[1905]), .B(n2619), .Z(n2620) );
  XOR U3550 ( .A(y[1909]), .B(n2603), .Z(n2604) );
  XOR U3551 ( .A(y[1913]), .B(n2587), .Z(n2588) );
  XOR U3552 ( .A(y[1917]), .B(n2571), .Z(n2572) );
  XOR U3553 ( .A(y[1921]), .B(n2555), .Z(n2556) );
  XOR U3554 ( .A(y[1925]), .B(n2539), .Z(n2540) );
  XOR U3555 ( .A(y[1929]), .B(n2523), .Z(n2524) );
  XOR U3556 ( .A(y[1933]), .B(n2507), .Z(n2508) );
  XOR U3557 ( .A(y[1937]), .B(n2491), .Z(n2492) );
  XOR U3558 ( .A(y[1941]), .B(n2475), .Z(n2476) );
  XOR U3559 ( .A(y[1945]), .B(n2459), .Z(n2460) );
  XOR U3560 ( .A(y[1949]), .B(n2443), .Z(n2444) );
  XOR U3561 ( .A(y[1953]), .B(n2427), .Z(n2428) );
  XOR U3562 ( .A(y[1957]), .B(n2411), .Z(n2412) );
  XOR U3563 ( .A(y[1961]), .B(n2395), .Z(n2396) );
  XOR U3564 ( .A(y[1965]), .B(n2379), .Z(n2380) );
  XOR U3565 ( .A(y[1969]), .B(n2363), .Z(n2364) );
  XOR U3566 ( .A(y[1973]), .B(n2347), .Z(n2348) );
  XOR U3567 ( .A(y[1977]), .B(n2331), .Z(n2332) );
  XOR U3568 ( .A(y[1981]), .B(n2315), .Z(n2316) );
  XOR U3569 ( .A(y[1985]), .B(n2299), .Z(n2300) );
  XOR U3570 ( .A(y[1989]), .B(n2283), .Z(n2284) );
  XOR U3571 ( .A(y[1993]), .B(n2267), .Z(n2268) );
  XOR U3572 ( .A(y[1997]), .B(n2251), .Z(n2252) );
  XOR U3573 ( .A(y[2001]), .B(n2235), .Z(n2236) );
  XOR U3574 ( .A(y[2005]), .B(n2219), .Z(n2220) );
  XOR U3575 ( .A(y[2009]), .B(n2203), .Z(n2204) );
  XOR U3576 ( .A(y[2013]), .B(n2187), .Z(n2188) );
  XOR U3577 ( .A(y[2017]), .B(n2171), .Z(n2172) );
  XOR U3578 ( .A(y[2021]), .B(n2155), .Z(n2156) );
  XOR U3579 ( .A(y[2025]), .B(n2139), .Z(n2140) );
  XOR U3580 ( .A(y[2029]), .B(n2123), .Z(n2124) );
  XOR U3581 ( .A(y[2033]), .B(n2107), .Z(n2108) );
  XOR U3582 ( .A(y[2037]), .B(n2091), .Z(n2092) );
  XOR U3583 ( .A(y[2041]), .B(n2075), .Z(n2076) );
  XOR U3584 ( .A(y[2045]), .B(n2059), .Z(n2060) );
  XOR U3585 ( .A(y[2]), .B(n10231), .Z(n10232) );
  XOR U3586 ( .A(y[6]), .B(n10215), .Z(n10216) );
  XOR U3587 ( .A(y[10]), .B(n10199), .Z(n10200) );
  XOR U3588 ( .A(y[14]), .B(n10183), .Z(n10184) );
  XOR U3589 ( .A(y[18]), .B(n10167), .Z(n10168) );
  XOR U3590 ( .A(y[22]), .B(n10151), .Z(n10152) );
  XOR U3591 ( .A(y[26]), .B(n10135), .Z(n10136) );
  XOR U3592 ( .A(y[30]), .B(n10119), .Z(n10120) );
  XOR U3593 ( .A(y[34]), .B(n10103), .Z(n10104) );
  XOR U3594 ( .A(y[38]), .B(n10087), .Z(n10088) );
  XOR U3595 ( .A(y[42]), .B(n10071), .Z(n10072) );
  XOR U3596 ( .A(y[46]), .B(n10055), .Z(n10056) );
  XOR U3597 ( .A(y[50]), .B(n10039), .Z(n10040) );
  XOR U3598 ( .A(y[54]), .B(n10023), .Z(n10024) );
  XOR U3599 ( .A(y[58]), .B(n10007), .Z(n10008) );
  XOR U3600 ( .A(y[62]), .B(n9991), .Z(n9992) );
  XOR U3601 ( .A(y[66]), .B(n9975), .Z(n9976) );
  XOR U3602 ( .A(y[70]), .B(n9959), .Z(n9960) );
  XOR U3603 ( .A(y[74]), .B(n9943), .Z(n9944) );
  XOR U3604 ( .A(y[78]), .B(n9927), .Z(n9928) );
  XOR U3605 ( .A(y[82]), .B(n9911), .Z(n9912) );
  XOR U3606 ( .A(y[86]), .B(n9895), .Z(n9896) );
  XOR U3607 ( .A(y[90]), .B(n9879), .Z(n9880) );
  XOR U3608 ( .A(y[94]), .B(n9863), .Z(n9864) );
  XOR U3609 ( .A(y[98]), .B(n9847), .Z(n9848) );
  XOR U3610 ( .A(y[102]), .B(n9831), .Z(n9832) );
  XOR U3611 ( .A(y[106]), .B(n9815), .Z(n9816) );
  XOR U3612 ( .A(y[110]), .B(n9799), .Z(n9800) );
  XOR U3613 ( .A(y[114]), .B(n9783), .Z(n9784) );
  XOR U3614 ( .A(y[118]), .B(n9767), .Z(n9768) );
  XOR U3615 ( .A(y[122]), .B(n9751), .Z(n9752) );
  XOR U3616 ( .A(y[126]), .B(n9735), .Z(n9736) );
  XOR U3617 ( .A(y[130]), .B(n9719), .Z(n9720) );
  XOR U3618 ( .A(y[134]), .B(n9703), .Z(n9704) );
  XOR U3619 ( .A(y[138]), .B(n9687), .Z(n9688) );
  XOR U3620 ( .A(y[142]), .B(n9671), .Z(n9672) );
  XOR U3621 ( .A(y[146]), .B(n9655), .Z(n9656) );
  XOR U3622 ( .A(y[150]), .B(n9639), .Z(n9640) );
  XOR U3623 ( .A(y[154]), .B(n9623), .Z(n9624) );
  XOR U3624 ( .A(y[158]), .B(n9607), .Z(n9608) );
  XOR U3625 ( .A(y[162]), .B(n9591), .Z(n9592) );
  XOR U3626 ( .A(y[166]), .B(n9575), .Z(n9576) );
  XOR U3627 ( .A(y[170]), .B(n9559), .Z(n9560) );
  XOR U3628 ( .A(y[174]), .B(n9543), .Z(n9544) );
  XOR U3629 ( .A(y[178]), .B(n9527), .Z(n9528) );
  XOR U3630 ( .A(y[182]), .B(n9511), .Z(n9512) );
  XOR U3631 ( .A(y[186]), .B(n9495), .Z(n9496) );
  XOR U3632 ( .A(y[190]), .B(n9479), .Z(n9480) );
  XOR U3633 ( .A(y[194]), .B(n9463), .Z(n9464) );
  XOR U3634 ( .A(y[198]), .B(n9447), .Z(n9448) );
  XOR U3635 ( .A(y[202]), .B(n9431), .Z(n9432) );
  XOR U3636 ( .A(y[206]), .B(n9415), .Z(n9416) );
  XOR U3637 ( .A(y[210]), .B(n9399), .Z(n9400) );
  XOR U3638 ( .A(y[214]), .B(n9383), .Z(n9384) );
  XOR U3639 ( .A(y[218]), .B(n9367), .Z(n9368) );
  XOR U3640 ( .A(y[222]), .B(n9351), .Z(n9352) );
  XOR U3641 ( .A(y[226]), .B(n9335), .Z(n9336) );
  XOR U3642 ( .A(y[230]), .B(n9319), .Z(n9320) );
  XOR U3643 ( .A(y[234]), .B(n9303), .Z(n9304) );
  XOR U3644 ( .A(y[238]), .B(n9287), .Z(n9288) );
  XOR U3645 ( .A(y[242]), .B(n9271), .Z(n9272) );
  XOR U3646 ( .A(y[246]), .B(n9255), .Z(n9256) );
  XOR U3647 ( .A(y[250]), .B(n9239), .Z(n9240) );
  XOR U3648 ( .A(y[254]), .B(n9223), .Z(n9224) );
  XOR U3649 ( .A(y[258]), .B(n9207), .Z(n9208) );
  XOR U3650 ( .A(y[262]), .B(n9191), .Z(n9192) );
  XOR U3651 ( .A(y[266]), .B(n9175), .Z(n9176) );
  XOR U3652 ( .A(y[270]), .B(n9159), .Z(n9160) );
  XOR U3653 ( .A(y[274]), .B(n9143), .Z(n9144) );
  XOR U3654 ( .A(y[278]), .B(n9127), .Z(n9128) );
  XOR U3655 ( .A(y[282]), .B(n9111), .Z(n9112) );
  XOR U3656 ( .A(y[286]), .B(n9095), .Z(n9096) );
  XOR U3657 ( .A(y[290]), .B(n9079), .Z(n9080) );
  XOR U3658 ( .A(y[294]), .B(n9063), .Z(n9064) );
  XOR U3659 ( .A(y[298]), .B(n9047), .Z(n9048) );
  XOR U3660 ( .A(y[302]), .B(n9031), .Z(n9032) );
  XOR U3661 ( .A(y[306]), .B(n9015), .Z(n9016) );
  XOR U3662 ( .A(y[310]), .B(n8999), .Z(n9000) );
  XOR U3663 ( .A(y[314]), .B(n8983), .Z(n8984) );
  XOR U3664 ( .A(y[318]), .B(n8967), .Z(n8968) );
  XOR U3665 ( .A(y[322]), .B(n8951), .Z(n8952) );
  XOR U3666 ( .A(y[326]), .B(n8935), .Z(n8936) );
  XOR U3667 ( .A(y[330]), .B(n8919), .Z(n8920) );
  XOR U3668 ( .A(y[334]), .B(n8903), .Z(n8904) );
  XOR U3669 ( .A(y[338]), .B(n8887), .Z(n8888) );
  XOR U3670 ( .A(y[342]), .B(n8871), .Z(n8872) );
  XOR U3671 ( .A(y[346]), .B(n8855), .Z(n8856) );
  XOR U3672 ( .A(y[350]), .B(n8839), .Z(n8840) );
  XOR U3673 ( .A(y[354]), .B(n8823), .Z(n8824) );
  XOR U3674 ( .A(y[358]), .B(n8807), .Z(n8808) );
  XOR U3675 ( .A(y[362]), .B(n8791), .Z(n8792) );
  XOR U3676 ( .A(y[366]), .B(n8775), .Z(n8776) );
  XOR U3677 ( .A(y[370]), .B(n8759), .Z(n8760) );
  XOR U3678 ( .A(y[374]), .B(n8743), .Z(n8744) );
  XOR U3679 ( .A(y[378]), .B(n8727), .Z(n8728) );
  XOR U3680 ( .A(y[382]), .B(n8711), .Z(n8712) );
  XOR U3681 ( .A(y[386]), .B(n8695), .Z(n8696) );
  XOR U3682 ( .A(y[390]), .B(n8679), .Z(n8680) );
  XOR U3683 ( .A(y[394]), .B(n8663), .Z(n8664) );
  XOR U3684 ( .A(y[398]), .B(n8647), .Z(n8648) );
  XOR U3685 ( .A(y[402]), .B(n8631), .Z(n8632) );
  XOR U3686 ( .A(y[406]), .B(n8615), .Z(n8616) );
  XOR U3687 ( .A(y[410]), .B(n8599), .Z(n8600) );
  XOR U3688 ( .A(y[414]), .B(n8583), .Z(n8584) );
  XOR U3689 ( .A(y[418]), .B(n8567), .Z(n8568) );
  XOR U3690 ( .A(y[422]), .B(n8551), .Z(n8552) );
  XOR U3691 ( .A(y[426]), .B(n8535), .Z(n8536) );
  XOR U3692 ( .A(y[430]), .B(n8519), .Z(n8520) );
  XOR U3693 ( .A(y[434]), .B(n8503), .Z(n8504) );
  XOR U3694 ( .A(y[438]), .B(n8487), .Z(n8488) );
  XOR U3695 ( .A(y[442]), .B(n8471), .Z(n8472) );
  XOR U3696 ( .A(y[446]), .B(n8455), .Z(n8456) );
  XOR U3697 ( .A(y[450]), .B(n8439), .Z(n8440) );
  XOR U3698 ( .A(y[454]), .B(n8423), .Z(n8424) );
  XOR U3699 ( .A(y[458]), .B(n8407), .Z(n8408) );
  XOR U3700 ( .A(y[462]), .B(n8391), .Z(n8392) );
  XOR U3701 ( .A(y[466]), .B(n8375), .Z(n8376) );
  XOR U3702 ( .A(y[470]), .B(n8359), .Z(n8360) );
  XOR U3703 ( .A(y[474]), .B(n8343), .Z(n8344) );
  XOR U3704 ( .A(y[478]), .B(n8327), .Z(n8328) );
  XOR U3705 ( .A(y[482]), .B(n8311), .Z(n8312) );
  XOR U3706 ( .A(y[486]), .B(n8295), .Z(n8296) );
  XOR U3707 ( .A(y[490]), .B(n8279), .Z(n8280) );
  XOR U3708 ( .A(y[494]), .B(n8263), .Z(n8264) );
  XOR U3709 ( .A(y[498]), .B(n8247), .Z(n8248) );
  XOR U3710 ( .A(y[502]), .B(n8231), .Z(n8232) );
  XOR U3711 ( .A(y[506]), .B(n8215), .Z(n8216) );
  XOR U3712 ( .A(y[510]), .B(n8199), .Z(n8200) );
  XOR U3713 ( .A(y[514]), .B(n8183), .Z(n8184) );
  XOR U3714 ( .A(y[518]), .B(n8167), .Z(n8168) );
  XOR U3715 ( .A(y[522]), .B(n8151), .Z(n8152) );
  XOR U3716 ( .A(y[526]), .B(n8135), .Z(n8136) );
  XOR U3717 ( .A(y[530]), .B(n8119), .Z(n8120) );
  XOR U3718 ( .A(y[534]), .B(n8103), .Z(n8104) );
  XOR U3719 ( .A(y[538]), .B(n8087), .Z(n8088) );
  XOR U3720 ( .A(y[542]), .B(n8071), .Z(n8072) );
  XOR U3721 ( .A(y[546]), .B(n8055), .Z(n8056) );
  XOR U3722 ( .A(y[550]), .B(n8039), .Z(n8040) );
  XOR U3723 ( .A(y[554]), .B(n8023), .Z(n8024) );
  XOR U3724 ( .A(y[558]), .B(n8007), .Z(n8008) );
  XOR U3725 ( .A(y[562]), .B(n7991), .Z(n7992) );
  XOR U3726 ( .A(y[566]), .B(n7975), .Z(n7976) );
  XOR U3727 ( .A(y[570]), .B(n7959), .Z(n7960) );
  XOR U3728 ( .A(y[574]), .B(n7943), .Z(n7944) );
  XOR U3729 ( .A(y[578]), .B(n7927), .Z(n7928) );
  XOR U3730 ( .A(y[582]), .B(n7911), .Z(n7912) );
  XOR U3731 ( .A(y[586]), .B(n7895), .Z(n7896) );
  XOR U3732 ( .A(y[590]), .B(n7879), .Z(n7880) );
  XOR U3733 ( .A(y[594]), .B(n7863), .Z(n7864) );
  XOR U3734 ( .A(y[598]), .B(n7847), .Z(n7848) );
  XOR U3735 ( .A(y[602]), .B(n7831), .Z(n7832) );
  XOR U3736 ( .A(y[606]), .B(n7815), .Z(n7816) );
  XOR U3737 ( .A(y[610]), .B(n7799), .Z(n7800) );
  XOR U3738 ( .A(y[614]), .B(n7783), .Z(n7784) );
  XOR U3739 ( .A(y[618]), .B(n7767), .Z(n7768) );
  XOR U3740 ( .A(y[622]), .B(n7751), .Z(n7752) );
  XOR U3741 ( .A(y[626]), .B(n7735), .Z(n7736) );
  XOR U3742 ( .A(y[630]), .B(n7719), .Z(n7720) );
  XOR U3743 ( .A(y[634]), .B(n7703), .Z(n7704) );
  XOR U3744 ( .A(y[638]), .B(n7687), .Z(n7688) );
  XOR U3745 ( .A(y[642]), .B(n7671), .Z(n7672) );
  XOR U3746 ( .A(y[646]), .B(n7655), .Z(n7656) );
  XOR U3747 ( .A(y[650]), .B(n7639), .Z(n7640) );
  XOR U3748 ( .A(y[654]), .B(n7623), .Z(n7624) );
  XOR U3749 ( .A(y[658]), .B(n7607), .Z(n7608) );
  XOR U3750 ( .A(y[662]), .B(n7591), .Z(n7592) );
  XOR U3751 ( .A(y[666]), .B(n7575), .Z(n7576) );
  XOR U3752 ( .A(y[670]), .B(n7559), .Z(n7560) );
  XOR U3753 ( .A(y[674]), .B(n7543), .Z(n7544) );
  XOR U3754 ( .A(y[678]), .B(n7527), .Z(n7528) );
  XOR U3755 ( .A(y[682]), .B(n7511), .Z(n7512) );
  XOR U3756 ( .A(y[686]), .B(n7495), .Z(n7496) );
  XOR U3757 ( .A(y[690]), .B(n7479), .Z(n7480) );
  XOR U3758 ( .A(y[694]), .B(n7463), .Z(n7464) );
  XOR U3759 ( .A(y[698]), .B(n7447), .Z(n7448) );
  XOR U3760 ( .A(y[702]), .B(n7431), .Z(n7432) );
  XOR U3761 ( .A(y[706]), .B(n7415), .Z(n7416) );
  XOR U3762 ( .A(y[710]), .B(n7399), .Z(n7400) );
  XOR U3763 ( .A(y[714]), .B(n7383), .Z(n7384) );
  XOR U3764 ( .A(y[718]), .B(n7367), .Z(n7368) );
  XOR U3765 ( .A(y[722]), .B(n7351), .Z(n7352) );
  XOR U3766 ( .A(y[726]), .B(n7335), .Z(n7336) );
  XOR U3767 ( .A(y[730]), .B(n7319), .Z(n7320) );
  XOR U3768 ( .A(y[734]), .B(n7303), .Z(n7304) );
  XOR U3769 ( .A(y[738]), .B(n7287), .Z(n7288) );
  XOR U3770 ( .A(y[742]), .B(n7271), .Z(n7272) );
  XOR U3771 ( .A(y[746]), .B(n7255), .Z(n7256) );
  XOR U3772 ( .A(y[750]), .B(n7239), .Z(n7240) );
  XOR U3773 ( .A(y[754]), .B(n7223), .Z(n7224) );
  XOR U3774 ( .A(y[758]), .B(n7207), .Z(n7208) );
  XOR U3775 ( .A(y[762]), .B(n7191), .Z(n7192) );
  XOR U3776 ( .A(y[766]), .B(n7175), .Z(n7176) );
  XOR U3777 ( .A(y[770]), .B(n7159), .Z(n7160) );
  XOR U3778 ( .A(y[774]), .B(n7143), .Z(n7144) );
  XOR U3779 ( .A(y[778]), .B(n7127), .Z(n7128) );
  XOR U3780 ( .A(y[782]), .B(n7111), .Z(n7112) );
  XOR U3781 ( .A(y[786]), .B(n7095), .Z(n7096) );
  XOR U3782 ( .A(y[790]), .B(n7079), .Z(n7080) );
  XOR U3783 ( .A(y[794]), .B(n7063), .Z(n7064) );
  XOR U3784 ( .A(y[798]), .B(n7047), .Z(n7048) );
  XOR U3785 ( .A(y[802]), .B(n7031), .Z(n7032) );
  XOR U3786 ( .A(y[806]), .B(n7015), .Z(n7016) );
  XOR U3787 ( .A(y[810]), .B(n6999), .Z(n7000) );
  XOR U3788 ( .A(y[814]), .B(n6983), .Z(n6984) );
  XOR U3789 ( .A(y[818]), .B(n6967), .Z(n6968) );
  XOR U3790 ( .A(y[822]), .B(n6951), .Z(n6952) );
  XOR U3791 ( .A(y[826]), .B(n6935), .Z(n6936) );
  XOR U3792 ( .A(y[830]), .B(n6919), .Z(n6920) );
  XOR U3793 ( .A(y[834]), .B(n6903), .Z(n6904) );
  XOR U3794 ( .A(y[838]), .B(n6887), .Z(n6888) );
  XOR U3795 ( .A(y[842]), .B(n6871), .Z(n6872) );
  XOR U3796 ( .A(y[846]), .B(n6855), .Z(n6856) );
  XOR U3797 ( .A(y[850]), .B(n6839), .Z(n6840) );
  XOR U3798 ( .A(y[854]), .B(n6823), .Z(n6824) );
  XOR U3799 ( .A(y[858]), .B(n6807), .Z(n6808) );
  XOR U3800 ( .A(y[862]), .B(n6791), .Z(n6792) );
  XOR U3801 ( .A(y[866]), .B(n6775), .Z(n6776) );
  XOR U3802 ( .A(y[870]), .B(n6759), .Z(n6760) );
  XOR U3803 ( .A(y[874]), .B(n6743), .Z(n6744) );
  XOR U3804 ( .A(y[878]), .B(n6727), .Z(n6728) );
  XOR U3805 ( .A(y[882]), .B(n6711), .Z(n6712) );
  XOR U3806 ( .A(y[886]), .B(n6695), .Z(n6696) );
  XOR U3807 ( .A(y[890]), .B(n6679), .Z(n6680) );
  XOR U3808 ( .A(y[894]), .B(n6663), .Z(n6664) );
  XOR U3809 ( .A(y[898]), .B(n6647), .Z(n6648) );
  XOR U3810 ( .A(y[902]), .B(n6631), .Z(n6632) );
  XOR U3811 ( .A(y[906]), .B(n6615), .Z(n6616) );
  XOR U3812 ( .A(y[910]), .B(n6599), .Z(n6600) );
  XOR U3813 ( .A(y[914]), .B(n6583), .Z(n6584) );
  XOR U3814 ( .A(y[918]), .B(n6567), .Z(n6568) );
  XOR U3815 ( .A(y[922]), .B(n6551), .Z(n6552) );
  XOR U3816 ( .A(y[926]), .B(n6535), .Z(n6536) );
  XOR U3817 ( .A(y[930]), .B(n6519), .Z(n6520) );
  XOR U3818 ( .A(y[934]), .B(n6503), .Z(n6504) );
  XOR U3819 ( .A(y[938]), .B(n6487), .Z(n6488) );
  XOR U3820 ( .A(y[942]), .B(n6471), .Z(n6472) );
  XOR U3821 ( .A(y[946]), .B(n6455), .Z(n6456) );
  XOR U3822 ( .A(y[950]), .B(n6439), .Z(n6440) );
  XOR U3823 ( .A(y[954]), .B(n6423), .Z(n6424) );
  XOR U3824 ( .A(y[958]), .B(n6407), .Z(n6408) );
  XOR U3825 ( .A(y[962]), .B(n6391), .Z(n6392) );
  XOR U3826 ( .A(y[966]), .B(n6375), .Z(n6376) );
  XOR U3827 ( .A(y[970]), .B(n6359), .Z(n6360) );
  XOR U3828 ( .A(y[974]), .B(n6343), .Z(n6344) );
  XOR U3829 ( .A(y[978]), .B(n6327), .Z(n6328) );
  XOR U3830 ( .A(y[982]), .B(n6311), .Z(n6312) );
  XOR U3831 ( .A(y[986]), .B(n6295), .Z(n6296) );
  XOR U3832 ( .A(y[990]), .B(n6279), .Z(n6280) );
  XOR U3833 ( .A(y[994]), .B(n6263), .Z(n6264) );
  XOR U3834 ( .A(y[998]), .B(n6247), .Z(n6248) );
  XOR U3835 ( .A(y[1002]), .B(n6231), .Z(n6232) );
  XOR U3836 ( .A(y[1006]), .B(n6215), .Z(n6216) );
  XOR U3837 ( .A(y[1010]), .B(n6199), .Z(n6200) );
  XOR U3838 ( .A(y[1014]), .B(n6183), .Z(n6184) );
  XOR U3839 ( .A(y[1018]), .B(n6167), .Z(n6168) );
  XOR U3840 ( .A(y[1022]), .B(n6151), .Z(n6152) );
  XOR U3841 ( .A(y[1026]), .B(n6135), .Z(n6136) );
  XOR U3842 ( .A(y[1030]), .B(n6119), .Z(n6120) );
  XOR U3843 ( .A(y[1034]), .B(n6103), .Z(n6104) );
  XOR U3844 ( .A(y[1038]), .B(n6087), .Z(n6088) );
  XOR U3845 ( .A(y[1042]), .B(n6071), .Z(n6072) );
  XOR U3846 ( .A(y[1046]), .B(n6055), .Z(n6056) );
  XOR U3847 ( .A(y[1050]), .B(n6039), .Z(n6040) );
  XOR U3848 ( .A(y[1054]), .B(n6023), .Z(n6024) );
  XOR U3849 ( .A(y[1058]), .B(n6007), .Z(n6008) );
  XOR U3850 ( .A(y[1062]), .B(n5991), .Z(n5992) );
  XOR U3851 ( .A(y[1066]), .B(n5975), .Z(n5976) );
  XOR U3852 ( .A(y[1070]), .B(n5959), .Z(n5960) );
  XOR U3853 ( .A(y[1074]), .B(n5943), .Z(n5944) );
  XOR U3854 ( .A(y[1078]), .B(n5927), .Z(n5928) );
  XOR U3855 ( .A(y[1082]), .B(n5911), .Z(n5912) );
  XOR U3856 ( .A(y[1086]), .B(n5895), .Z(n5896) );
  XOR U3857 ( .A(y[1090]), .B(n5879), .Z(n5880) );
  XOR U3858 ( .A(y[1094]), .B(n5863), .Z(n5864) );
  XOR U3859 ( .A(y[1098]), .B(n5847), .Z(n5848) );
  XOR U3860 ( .A(y[1102]), .B(n5831), .Z(n5832) );
  XOR U3861 ( .A(y[1106]), .B(n5815), .Z(n5816) );
  XOR U3862 ( .A(y[1110]), .B(n5799), .Z(n5800) );
  XOR U3863 ( .A(y[1114]), .B(n5783), .Z(n5784) );
  XOR U3864 ( .A(y[1118]), .B(n5767), .Z(n5768) );
  XOR U3865 ( .A(y[1122]), .B(n5751), .Z(n5752) );
  XOR U3866 ( .A(y[1126]), .B(n5735), .Z(n5736) );
  XOR U3867 ( .A(y[1130]), .B(n5719), .Z(n5720) );
  XOR U3868 ( .A(y[1134]), .B(n5703), .Z(n5704) );
  XOR U3869 ( .A(y[1138]), .B(n5687), .Z(n5688) );
  XOR U3870 ( .A(y[1142]), .B(n5671), .Z(n5672) );
  XOR U3871 ( .A(y[1146]), .B(n5655), .Z(n5656) );
  XOR U3872 ( .A(y[1150]), .B(n5639), .Z(n5640) );
  XOR U3873 ( .A(y[1154]), .B(n5623), .Z(n5624) );
  XOR U3874 ( .A(y[1158]), .B(n5607), .Z(n5608) );
  XOR U3875 ( .A(y[1162]), .B(n5591), .Z(n5592) );
  XOR U3876 ( .A(y[1166]), .B(n5575), .Z(n5576) );
  XOR U3877 ( .A(y[1170]), .B(n5559), .Z(n5560) );
  XOR U3878 ( .A(y[1174]), .B(n5543), .Z(n5544) );
  XOR U3879 ( .A(y[1178]), .B(n5527), .Z(n5528) );
  XOR U3880 ( .A(y[1182]), .B(n5511), .Z(n5512) );
  XOR U3881 ( .A(y[1186]), .B(n5495), .Z(n5496) );
  XOR U3882 ( .A(y[1190]), .B(n5479), .Z(n5480) );
  XOR U3883 ( .A(y[1194]), .B(n5463), .Z(n5464) );
  XOR U3884 ( .A(y[1198]), .B(n5447), .Z(n5448) );
  XOR U3885 ( .A(y[1202]), .B(n5431), .Z(n5432) );
  XOR U3886 ( .A(y[1206]), .B(n5415), .Z(n5416) );
  XOR U3887 ( .A(y[1210]), .B(n5399), .Z(n5400) );
  XOR U3888 ( .A(y[1214]), .B(n5383), .Z(n5384) );
  XOR U3889 ( .A(y[1218]), .B(n5367), .Z(n5368) );
  XOR U3890 ( .A(y[1222]), .B(n5351), .Z(n5352) );
  XOR U3891 ( .A(y[1226]), .B(n5335), .Z(n5336) );
  XOR U3892 ( .A(y[1230]), .B(n5319), .Z(n5320) );
  XOR U3893 ( .A(y[1234]), .B(n5303), .Z(n5304) );
  XOR U3894 ( .A(y[1238]), .B(n5287), .Z(n5288) );
  XOR U3895 ( .A(y[1242]), .B(n5271), .Z(n5272) );
  XOR U3896 ( .A(y[1246]), .B(n5255), .Z(n5256) );
  XOR U3897 ( .A(y[1250]), .B(n5239), .Z(n5240) );
  XOR U3898 ( .A(y[1254]), .B(n5223), .Z(n5224) );
  XOR U3899 ( .A(y[1258]), .B(n5207), .Z(n5208) );
  XOR U3900 ( .A(y[1262]), .B(n5191), .Z(n5192) );
  XOR U3901 ( .A(y[1266]), .B(n5175), .Z(n5176) );
  XOR U3902 ( .A(y[1270]), .B(n5159), .Z(n5160) );
  XOR U3903 ( .A(y[1274]), .B(n5143), .Z(n5144) );
  XOR U3904 ( .A(y[1278]), .B(n5127), .Z(n5128) );
  XOR U3905 ( .A(y[1282]), .B(n5111), .Z(n5112) );
  XOR U3906 ( .A(y[1286]), .B(n5095), .Z(n5096) );
  XOR U3907 ( .A(y[1290]), .B(n5079), .Z(n5080) );
  XOR U3908 ( .A(y[1294]), .B(n5063), .Z(n5064) );
  XOR U3909 ( .A(y[1298]), .B(n5047), .Z(n5048) );
  XOR U3910 ( .A(y[1302]), .B(n5031), .Z(n5032) );
  XOR U3911 ( .A(y[1306]), .B(n5015), .Z(n5016) );
  XOR U3912 ( .A(y[1310]), .B(n4999), .Z(n5000) );
  XOR U3913 ( .A(y[1314]), .B(n4983), .Z(n4984) );
  XOR U3914 ( .A(y[1318]), .B(n4967), .Z(n4968) );
  XOR U3915 ( .A(y[1322]), .B(n4951), .Z(n4952) );
  XOR U3916 ( .A(y[1326]), .B(n4935), .Z(n4936) );
  XOR U3917 ( .A(y[1330]), .B(n4919), .Z(n4920) );
  XOR U3918 ( .A(y[1334]), .B(n4903), .Z(n4904) );
  XOR U3919 ( .A(y[1338]), .B(n4887), .Z(n4888) );
  XOR U3920 ( .A(y[1342]), .B(n4871), .Z(n4872) );
  XOR U3921 ( .A(y[1346]), .B(n4855), .Z(n4856) );
  XOR U3922 ( .A(y[1350]), .B(n4839), .Z(n4840) );
  XOR U3923 ( .A(y[1354]), .B(n4823), .Z(n4824) );
  XOR U3924 ( .A(y[1358]), .B(n4807), .Z(n4808) );
  XOR U3925 ( .A(y[1362]), .B(n4791), .Z(n4792) );
  XOR U3926 ( .A(y[1366]), .B(n4775), .Z(n4776) );
  XOR U3927 ( .A(y[1370]), .B(n4759), .Z(n4760) );
  XOR U3928 ( .A(y[1374]), .B(n4743), .Z(n4744) );
  XOR U3929 ( .A(y[1378]), .B(n4727), .Z(n4728) );
  XOR U3930 ( .A(y[1382]), .B(n4711), .Z(n4712) );
  XOR U3931 ( .A(y[1386]), .B(n4695), .Z(n4696) );
  XOR U3932 ( .A(y[1390]), .B(n4679), .Z(n4680) );
  XOR U3933 ( .A(y[1394]), .B(n4663), .Z(n4664) );
  XOR U3934 ( .A(y[1398]), .B(n4647), .Z(n4648) );
  XOR U3935 ( .A(y[1402]), .B(n4631), .Z(n4632) );
  XOR U3936 ( .A(y[1406]), .B(n4615), .Z(n4616) );
  XOR U3937 ( .A(y[1410]), .B(n4599), .Z(n4600) );
  XOR U3938 ( .A(y[1414]), .B(n4583), .Z(n4584) );
  XOR U3939 ( .A(y[1418]), .B(n4567), .Z(n4568) );
  XOR U3940 ( .A(y[1422]), .B(n4551), .Z(n4552) );
  XOR U3941 ( .A(y[1426]), .B(n4535), .Z(n4536) );
  XOR U3942 ( .A(y[1430]), .B(n4519), .Z(n4520) );
  XOR U3943 ( .A(y[1434]), .B(n4503), .Z(n4504) );
  XOR U3944 ( .A(y[1438]), .B(n4487), .Z(n4488) );
  XOR U3945 ( .A(y[1442]), .B(n4471), .Z(n4472) );
  XOR U3946 ( .A(y[1446]), .B(n4455), .Z(n4456) );
  XOR U3947 ( .A(y[1450]), .B(n4439), .Z(n4440) );
  XOR U3948 ( .A(y[1454]), .B(n4423), .Z(n4424) );
  XOR U3949 ( .A(y[1458]), .B(n4407), .Z(n4408) );
  XOR U3950 ( .A(y[1462]), .B(n4391), .Z(n4392) );
  XOR U3951 ( .A(y[1466]), .B(n4375), .Z(n4376) );
  XOR U3952 ( .A(y[1470]), .B(n4359), .Z(n4360) );
  XOR U3953 ( .A(y[1474]), .B(n4343), .Z(n4344) );
  XOR U3954 ( .A(y[1478]), .B(n4327), .Z(n4328) );
  XOR U3955 ( .A(y[1482]), .B(n4311), .Z(n4312) );
  XOR U3956 ( .A(y[1486]), .B(n4295), .Z(n4296) );
  XOR U3957 ( .A(y[1490]), .B(n4279), .Z(n4280) );
  XOR U3958 ( .A(y[1494]), .B(n4263), .Z(n4264) );
  XOR U3959 ( .A(y[1498]), .B(n4247), .Z(n4248) );
  XOR U3960 ( .A(y[1502]), .B(n4231), .Z(n4232) );
  XOR U3961 ( .A(y[1506]), .B(n4215), .Z(n4216) );
  XOR U3962 ( .A(y[1510]), .B(n4199), .Z(n4200) );
  XOR U3963 ( .A(y[1514]), .B(n4183), .Z(n4184) );
  XOR U3964 ( .A(y[1518]), .B(n4167), .Z(n4168) );
  XOR U3965 ( .A(y[1522]), .B(n4151), .Z(n4152) );
  XOR U3966 ( .A(y[1526]), .B(n4135), .Z(n4136) );
  XOR U3967 ( .A(y[1530]), .B(n4119), .Z(n4120) );
  XOR U3968 ( .A(y[1534]), .B(n4103), .Z(n4104) );
  XOR U3969 ( .A(y[1538]), .B(n4087), .Z(n4088) );
  XOR U3970 ( .A(y[1542]), .B(n4071), .Z(n4072) );
  XOR U3971 ( .A(y[1546]), .B(n4055), .Z(n4056) );
  XOR U3972 ( .A(y[1550]), .B(n4039), .Z(n4040) );
  XOR U3973 ( .A(y[1554]), .B(n4023), .Z(n4024) );
  XOR U3974 ( .A(y[1558]), .B(n4007), .Z(n4008) );
  XOR U3975 ( .A(y[1562]), .B(n3991), .Z(n3992) );
  XOR U3976 ( .A(y[1566]), .B(n3975), .Z(n3976) );
  XOR U3977 ( .A(y[1570]), .B(n3959), .Z(n3960) );
  XOR U3978 ( .A(y[1574]), .B(n3943), .Z(n3944) );
  XOR U3979 ( .A(y[1578]), .B(n3927), .Z(n3928) );
  XOR U3980 ( .A(y[1582]), .B(n3911), .Z(n3912) );
  XOR U3981 ( .A(y[1586]), .B(n3895), .Z(n3896) );
  XOR U3982 ( .A(y[1590]), .B(n3879), .Z(n3880) );
  XOR U3983 ( .A(y[1594]), .B(n3863), .Z(n3864) );
  XOR U3984 ( .A(y[1598]), .B(n3847), .Z(n3848) );
  XOR U3985 ( .A(y[1602]), .B(n3831), .Z(n3832) );
  XOR U3986 ( .A(y[1606]), .B(n3815), .Z(n3816) );
  XOR U3987 ( .A(y[1610]), .B(n3799), .Z(n3800) );
  XOR U3988 ( .A(y[1614]), .B(n3783), .Z(n3784) );
  XOR U3989 ( .A(y[1618]), .B(n3767), .Z(n3768) );
  XOR U3990 ( .A(y[1622]), .B(n3751), .Z(n3752) );
  XOR U3991 ( .A(y[1626]), .B(n3735), .Z(n3736) );
  XOR U3992 ( .A(y[1630]), .B(n3719), .Z(n3720) );
  XOR U3993 ( .A(y[1634]), .B(n3703), .Z(n3704) );
  XOR U3994 ( .A(y[1638]), .B(n3687), .Z(n3688) );
  XOR U3995 ( .A(y[1642]), .B(n3671), .Z(n3672) );
  XOR U3996 ( .A(y[1646]), .B(n3655), .Z(n3656) );
  XOR U3997 ( .A(y[1650]), .B(n3639), .Z(n3640) );
  XOR U3998 ( .A(y[1654]), .B(n3623), .Z(n3624) );
  XOR U3999 ( .A(y[1658]), .B(n3607), .Z(n3608) );
  XOR U4000 ( .A(y[1662]), .B(n3591), .Z(n3592) );
  XOR U4001 ( .A(y[1666]), .B(n3575), .Z(n3576) );
  XOR U4002 ( .A(y[1670]), .B(n3559), .Z(n3560) );
  XOR U4003 ( .A(y[1674]), .B(n3543), .Z(n3544) );
  XOR U4004 ( .A(y[1678]), .B(n3527), .Z(n3528) );
  XOR U4005 ( .A(y[1682]), .B(n3511), .Z(n3512) );
  XOR U4006 ( .A(y[1686]), .B(n3495), .Z(n3496) );
  XOR U4007 ( .A(y[1690]), .B(n3479), .Z(n3480) );
  XOR U4008 ( .A(y[1694]), .B(n3463), .Z(n3464) );
  XOR U4009 ( .A(y[1698]), .B(n3447), .Z(n3448) );
  XOR U4010 ( .A(y[1702]), .B(n3431), .Z(n3432) );
  XOR U4011 ( .A(y[1706]), .B(n3415), .Z(n3416) );
  XOR U4012 ( .A(y[1710]), .B(n3399), .Z(n3400) );
  XOR U4013 ( .A(y[1714]), .B(n3383), .Z(n3384) );
  XOR U4014 ( .A(y[1718]), .B(n3367), .Z(n3368) );
  XOR U4015 ( .A(y[1722]), .B(n3351), .Z(n3352) );
  XOR U4016 ( .A(y[1726]), .B(n3335), .Z(n3336) );
  XOR U4017 ( .A(y[1730]), .B(n3319), .Z(n3320) );
  XOR U4018 ( .A(y[1734]), .B(n3303), .Z(n3304) );
  XOR U4019 ( .A(y[1738]), .B(n3287), .Z(n3288) );
  XOR U4020 ( .A(y[1742]), .B(n3271), .Z(n3272) );
  XOR U4021 ( .A(y[1746]), .B(n3255), .Z(n3256) );
  XOR U4022 ( .A(y[1750]), .B(n3239), .Z(n3240) );
  XOR U4023 ( .A(y[1754]), .B(n3223), .Z(n3224) );
  XOR U4024 ( .A(y[1758]), .B(n3207), .Z(n3208) );
  XOR U4025 ( .A(y[1762]), .B(n3191), .Z(n3192) );
  XOR U4026 ( .A(y[1766]), .B(n3175), .Z(n3176) );
  XOR U4027 ( .A(y[1770]), .B(n3159), .Z(n3160) );
  XOR U4028 ( .A(y[1774]), .B(n3143), .Z(n3144) );
  XOR U4029 ( .A(y[1778]), .B(n3127), .Z(n3128) );
  XOR U4030 ( .A(y[1782]), .B(n3111), .Z(n3112) );
  XOR U4031 ( .A(y[1786]), .B(n3095), .Z(n3096) );
  XOR U4032 ( .A(y[1790]), .B(n3079), .Z(n3080) );
  XOR U4033 ( .A(y[1794]), .B(n3063), .Z(n3064) );
  XOR U4034 ( .A(y[1798]), .B(n3047), .Z(n3048) );
  XOR U4035 ( .A(y[1802]), .B(n3031), .Z(n3032) );
  XOR U4036 ( .A(y[1806]), .B(n3015), .Z(n3016) );
  XOR U4037 ( .A(y[1810]), .B(n2999), .Z(n3000) );
  XOR U4038 ( .A(y[1814]), .B(n2983), .Z(n2984) );
  XOR U4039 ( .A(y[1818]), .B(n2967), .Z(n2968) );
  XOR U4040 ( .A(y[1822]), .B(n2951), .Z(n2952) );
  XOR U4041 ( .A(y[1826]), .B(n2935), .Z(n2936) );
  XOR U4042 ( .A(y[1830]), .B(n2919), .Z(n2920) );
  XOR U4043 ( .A(y[1834]), .B(n2903), .Z(n2904) );
  XOR U4044 ( .A(y[1838]), .B(n2887), .Z(n2888) );
  XOR U4045 ( .A(y[1842]), .B(n2871), .Z(n2872) );
  XOR U4046 ( .A(y[1846]), .B(n2855), .Z(n2856) );
  XOR U4047 ( .A(y[1850]), .B(n2839), .Z(n2840) );
  XOR U4048 ( .A(y[1854]), .B(n2823), .Z(n2824) );
  XOR U4049 ( .A(y[1858]), .B(n2807), .Z(n2808) );
  XOR U4050 ( .A(y[1862]), .B(n2791), .Z(n2792) );
  XOR U4051 ( .A(y[1866]), .B(n2775), .Z(n2776) );
  XOR U4052 ( .A(y[1870]), .B(n2759), .Z(n2760) );
  XOR U4053 ( .A(y[1874]), .B(n2743), .Z(n2744) );
  XOR U4054 ( .A(y[1878]), .B(n2727), .Z(n2728) );
  XOR U4055 ( .A(y[1882]), .B(n2711), .Z(n2712) );
  XOR U4056 ( .A(y[1886]), .B(n2695), .Z(n2696) );
  XOR U4057 ( .A(y[1890]), .B(n2679), .Z(n2680) );
  XOR U4058 ( .A(y[1894]), .B(n2663), .Z(n2664) );
  XOR U4059 ( .A(y[1898]), .B(n2647), .Z(n2648) );
  XOR U4060 ( .A(y[1902]), .B(n2631), .Z(n2632) );
  XOR U4061 ( .A(y[1906]), .B(n2615), .Z(n2616) );
  XOR U4062 ( .A(y[1910]), .B(n2599), .Z(n2600) );
  XOR U4063 ( .A(y[1914]), .B(n2583), .Z(n2584) );
  XOR U4064 ( .A(y[1918]), .B(n2567), .Z(n2568) );
  XOR U4065 ( .A(y[1922]), .B(n2551), .Z(n2552) );
  XOR U4066 ( .A(y[1926]), .B(n2535), .Z(n2536) );
  XOR U4067 ( .A(y[1930]), .B(n2519), .Z(n2520) );
  XOR U4068 ( .A(y[1934]), .B(n2503), .Z(n2504) );
  XOR U4069 ( .A(y[1938]), .B(n2487), .Z(n2488) );
  XOR U4070 ( .A(y[1942]), .B(n2471), .Z(n2472) );
  XOR U4071 ( .A(y[1946]), .B(n2455), .Z(n2456) );
  XOR U4072 ( .A(y[1950]), .B(n2439), .Z(n2440) );
  XOR U4073 ( .A(y[1954]), .B(n2423), .Z(n2424) );
  XOR U4074 ( .A(y[1958]), .B(n2407), .Z(n2408) );
  XOR U4075 ( .A(y[1962]), .B(n2391), .Z(n2392) );
  XOR U4076 ( .A(y[1966]), .B(n2375), .Z(n2376) );
  XOR U4077 ( .A(y[1970]), .B(n2359), .Z(n2360) );
  XOR U4078 ( .A(y[1974]), .B(n2343), .Z(n2344) );
  XOR U4079 ( .A(y[1978]), .B(n2327), .Z(n2328) );
  XOR U4080 ( .A(y[1982]), .B(n2311), .Z(n2312) );
  XOR U4081 ( .A(y[1986]), .B(n2295), .Z(n2296) );
  XOR U4082 ( .A(y[1990]), .B(n2279), .Z(n2280) );
  XOR U4083 ( .A(y[1994]), .B(n2263), .Z(n2264) );
  XOR U4084 ( .A(y[1998]), .B(n2247), .Z(n2248) );
  XOR U4085 ( .A(y[2002]), .B(n2231), .Z(n2232) );
  XOR U4086 ( .A(y[2006]), .B(n2215), .Z(n2216) );
  XOR U4087 ( .A(y[2010]), .B(n2199), .Z(n2200) );
  XOR U4088 ( .A(y[2014]), .B(n2183), .Z(n2184) );
  XOR U4089 ( .A(y[2018]), .B(n2167), .Z(n2168) );
  XOR U4090 ( .A(y[2022]), .B(n2151), .Z(n2152) );
  XOR U4091 ( .A(y[2026]), .B(n2135), .Z(n2136) );
  XOR U4092 ( .A(y[2030]), .B(n2119), .Z(n2120) );
  XOR U4093 ( .A(y[2034]), .B(n2103), .Z(n2104) );
  XOR U4094 ( .A(y[2038]), .B(n2087), .Z(n2088) );
  XOR U4095 ( .A(y[2042]), .B(n2071), .Z(n2072) );
  XOR U4096 ( .A(y[2046]), .B(n2055), .Z(n2056) );
  XOR U4097 ( .A(n2050), .B(n2051), .Z(g) );
  AND U4098 ( .A(n2052), .B(n2053), .Z(n2050) );
  XOR U4099 ( .A(x[2047]), .B(n2051), .Z(n2053) );
  XNOR U4100 ( .A(y[2047]), .B(n2051), .Z(n2052) );
  XNOR U4101 ( .A(n2054), .B(n2055), .Z(n2051) );
  AND U4102 ( .A(n2056), .B(n2057), .Z(n2054) );
  XNOR U4103 ( .A(x[2046]), .B(n2055), .Z(n2057) );
  XOR U4104 ( .A(n2058), .B(n2059), .Z(n2055) );
  AND U4105 ( .A(n2060), .B(n2061), .Z(n2058) );
  XNOR U4106 ( .A(x[2045]), .B(n2059), .Z(n2061) );
  XOR U4107 ( .A(n2062), .B(n2063), .Z(n2059) );
  AND U4108 ( .A(n2064), .B(n2065), .Z(n2062) );
  XNOR U4109 ( .A(x[2044]), .B(n2063), .Z(n2065) );
  XOR U4110 ( .A(n2066), .B(n2067), .Z(n2063) );
  AND U4111 ( .A(n2068), .B(n2069), .Z(n2066) );
  XNOR U4112 ( .A(x[2043]), .B(n2067), .Z(n2069) );
  XOR U4113 ( .A(n2070), .B(n2071), .Z(n2067) );
  AND U4114 ( .A(n2072), .B(n2073), .Z(n2070) );
  XNOR U4115 ( .A(x[2042]), .B(n2071), .Z(n2073) );
  XOR U4116 ( .A(n2074), .B(n2075), .Z(n2071) );
  AND U4117 ( .A(n2076), .B(n2077), .Z(n2074) );
  XNOR U4118 ( .A(x[2041]), .B(n2075), .Z(n2077) );
  XOR U4119 ( .A(n2078), .B(n2079), .Z(n2075) );
  AND U4120 ( .A(n2080), .B(n2081), .Z(n2078) );
  XNOR U4121 ( .A(x[2040]), .B(n2079), .Z(n2081) );
  XOR U4122 ( .A(n2082), .B(n2083), .Z(n2079) );
  AND U4123 ( .A(n2084), .B(n2085), .Z(n2082) );
  XNOR U4124 ( .A(x[2039]), .B(n2083), .Z(n2085) );
  XOR U4125 ( .A(n2086), .B(n2087), .Z(n2083) );
  AND U4126 ( .A(n2088), .B(n2089), .Z(n2086) );
  XNOR U4127 ( .A(x[2038]), .B(n2087), .Z(n2089) );
  XOR U4128 ( .A(n2090), .B(n2091), .Z(n2087) );
  AND U4129 ( .A(n2092), .B(n2093), .Z(n2090) );
  XNOR U4130 ( .A(x[2037]), .B(n2091), .Z(n2093) );
  XOR U4131 ( .A(n2094), .B(n2095), .Z(n2091) );
  AND U4132 ( .A(n2096), .B(n2097), .Z(n2094) );
  XNOR U4133 ( .A(x[2036]), .B(n2095), .Z(n2097) );
  XOR U4134 ( .A(n2098), .B(n2099), .Z(n2095) );
  AND U4135 ( .A(n2100), .B(n2101), .Z(n2098) );
  XNOR U4136 ( .A(x[2035]), .B(n2099), .Z(n2101) );
  XOR U4137 ( .A(n2102), .B(n2103), .Z(n2099) );
  AND U4138 ( .A(n2104), .B(n2105), .Z(n2102) );
  XNOR U4139 ( .A(x[2034]), .B(n2103), .Z(n2105) );
  XOR U4140 ( .A(n2106), .B(n2107), .Z(n2103) );
  AND U4141 ( .A(n2108), .B(n2109), .Z(n2106) );
  XNOR U4142 ( .A(x[2033]), .B(n2107), .Z(n2109) );
  XOR U4143 ( .A(n2110), .B(n2111), .Z(n2107) );
  AND U4144 ( .A(n2112), .B(n2113), .Z(n2110) );
  XNOR U4145 ( .A(x[2032]), .B(n2111), .Z(n2113) );
  XOR U4146 ( .A(n2114), .B(n2115), .Z(n2111) );
  AND U4147 ( .A(n2116), .B(n2117), .Z(n2114) );
  XNOR U4148 ( .A(x[2031]), .B(n2115), .Z(n2117) );
  XOR U4149 ( .A(n2118), .B(n2119), .Z(n2115) );
  AND U4150 ( .A(n2120), .B(n2121), .Z(n2118) );
  XNOR U4151 ( .A(x[2030]), .B(n2119), .Z(n2121) );
  XOR U4152 ( .A(n2122), .B(n2123), .Z(n2119) );
  AND U4153 ( .A(n2124), .B(n2125), .Z(n2122) );
  XNOR U4154 ( .A(x[2029]), .B(n2123), .Z(n2125) );
  XOR U4155 ( .A(n2126), .B(n2127), .Z(n2123) );
  AND U4156 ( .A(n2128), .B(n2129), .Z(n2126) );
  XNOR U4157 ( .A(x[2028]), .B(n2127), .Z(n2129) );
  XOR U4158 ( .A(n2130), .B(n2131), .Z(n2127) );
  AND U4159 ( .A(n2132), .B(n2133), .Z(n2130) );
  XNOR U4160 ( .A(x[2027]), .B(n2131), .Z(n2133) );
  XOR U4161 ( .A(n2134), .B(n2135), .Z(n2131) );
  AND U4162 ( .A(n2136), .B(n2137), .Z(n2134) );
  XNOR U4163 ( .A(x[2026]), .B(n2135), .Z(n2137) );
  XOR U4164 ( .A(n2138), .B(n2139), .Z(n2135) );
  AND U4165 ( .A(n2140), .B(n2141), .Z(n2138) );
  XNOR U4166 ( .A(x[2025]), .B(n2139), .Z(n2141) );
  XOR U4167 ( .A(n2142), .B(n2143), .Z(n2139) );
  AND U4168 ( .A(n2144), .B(n2145), .Z(n2142) );
  XNOR U4169 ( .A(x[2024]), .B(n2143), .Z(n2145) );
  XOR U4170 ( .A(n2146), .B(n2147), .Z(n2143) );
  AND U4171 ( .A(n2148), .B(n2149), .Z(n2146) );
  XNOR U4172 ( .A(x[2023]), .B(n2147), .Z(n2149) );
  XOR U4173 ( .A(n2150), .B(n2151), .Z(n2147) );
  AND U4174 ( .A(n2152), .B(n2153), .Z(n2150) );
  XNOR U4175 ( .A(x[2022]), .B(n2151), .Z(n2153) );
  XOR U4176 ( .A(n2154), .B(n2155), .Z(n2151) );
  AND U4177 ( .A(n2156), .B(n2157), .Z(n2154) );
  XNOR U4178 ( .A(x[2021]), .B(n2155), .Z(n2157) );
  XOR U4179 ( .A(n2158), .B(n2159), .Z(n2155) );
  AND U4180 ( .A(n2160), .B(n2161), .Z(n2158) );
  XNOR U4181 ( .A(x[2020]), .B(n2159), .Z(n2161) );
  XOR U4182 ( .A(n2162), .B(n2163), .Z(n2159) );
  AND U4183 ( .A(n2164), .B(n2165), .Z(n2162) );
  XNOR U4184 ( .A(x[2019]), .B(n2163), .Z(n2165) );
  XOR U4185 ( .A(n2166), .B(n2167), .Z(n2163) );
  AND U4186 ( .A(n2168), .B(n2169), .Z(n2166) );
  XNOR U4187 ( .A(x[2018]), .B(n2167), .Z(n2169) );
  XOR U4188 ( .A(n2170), .B(n2171), .Z(n2167) );
  AND U4189 ( .A(n2172), .B(n2173), .Z(n2170) );
  XNOR U4190 ( .A(x[2017]), .B(n2171), .Z(n2173) );
  XOR U4191 ( .A(n2174), .B(n2175), .Z(n2171) );
  AND U4192 ( .A(n2176), .B(n2177), .Z(n2174) );
  XNOR U4193 ( .A(x[2016]), .B(n2175), .Z(n2177) );
  XOR U4194 ( .A(n2178), .B(n2179), .Z(n2175) );
  AND U4195 ( .A(n2180), .B(n2181), .Z(n2178) );
  XNOR U4196 ( .A(x[2015]), .B(n2179), .Z(n2181) );
  XOR U4197 ( .A(n2182), .B(n2183), .Z(n2179) );
  AND U4198 ( .A(n2184), .B(n2185), .Z(n2182) );
  XNOR U4199 ( .A(x[2014]), .B(n2183), .Z(n2185) );
  XOR U4200 ( .A(n2186), .B(n2187), .Z(n2183) );
  AND U4201 ( .A(n2188), .B(n2189), .Z(n2186) );
  XNOR U4202 ( .A(x[2013]), .B(n2187), .Z(n2189) );
  XOR U4203 ( .A(n2190), .B(n2191), .Z(n2187) );
  AND U4204 ( .A(n2192), .B(n2193), .Z(n2190) );
  XNOR U4205 ( .A(x[2012]), .B(n2191), .Z(n2193) );
  XOR U4206 ( .A(n2194), .B(n2195), .Z(n2191) );
  AND U4207 ( .A(n2196), .B(n2197), .Z(n2194) );
  XNOR U4208 ( .A(x[2011]), .B(n2195), .Z(n2197) );
  XOR U4209 ( .A(n2198), .B(n2199), .Z(n2195) );
  AND U4210 ( .A(n2200), .B(n2201), .Z(n2198) );
  XNOR U4211 ( .A(x[2010]), .B(n2199), .Z(n2201) );
  XOR U4212 ( .A(n2202), .B(n2203), .Z(n2199) );
  AND U4213 ( .A(n2204), .B(n2205), .Z(n2202) );
  XNOR U4214 ( .A(x[2009]), .B(n2203), .Z(n2205) );
  XOR U4215 ( .A(n2206), .B(n2207), .Z(n2203) );
  AND U4216 ( .A(n2208), .B(n2209), .Z(n2206) );
  XNOR U4217 ( .A(x[2008]), .B(n2207), .Z(n2209) );
  XOR U4218 ( .A(n2210), .B(n2211), .Z(n2207) );
  AND U4219 ( .A(n2212), .B(n2213), .Z(n2210) );
  XNOR U4220 ( .A(x[2007]), .B(n2211), .Z(n2213) );
  XOR U4221 ( .A(n2214), .B(n2215), .Z(n2211) );
  AND U4222 ( .A(n2216), .B(n2217), .Z(n2214) );
  XNOR U4223 ( .A(x[2006]), .B(n2215), .Z(n2217) );
  XOR U4224 ( .A(n2218), .B(n2219), .Z(n2215) );
  AND U4225 ( .A(n2220), .B(n2221), .Z(n2218) );
  XNOR U4226 ( .A(x[2005]), .B(n2219), .Z(n2221) );
  XOR U4227 ( .A(n2222), .B(n2223), .Z(n2219) );
  AND U4228 ( .A(n2224), .B(n2225), .Z(n2222) );
  XNOR U4229 ( .A(x[2004]), .B(n2223), .Z(n2225) );
  XOR U4230 ( .A(n2226), .B(n2227), .Z(n2223) );
  AND U4231 ( .A(n2228), .B(n2229), .Z(n2226) );
  XNOR U4232 ( .A(x[2003]), .B(n2227), .Z(n2229) );
  XOR U4233 ( .A(n2230), .B(n2231), .Z(n2227) );
  AND U4234 ( .A(n2232), .B(n2233), .Z(n2230) );
  XNOR U4235 ( .A(x[2002]), .B(n2231), .Z(n2233) );
  XOR U4236 ( .A(n2234), .B(n2235), .Z(n2231) );
  AND U4237 ( .A(n2236), .B(n2237), .Z(n2234) );
  XNOR U4238 ( .A(x[2001]), .B(n2235), .Z(n2237) );
  XOR U4239 ( .A(n2238), .B(n2239), .Z(n2235) );
  AND U4240 ( .A(n2240), .B(n2241), .Z(n2238) );
  XNOR U4241 ( .A(x[2000]), .B(n2239), .Z(n2241) );
  XOR U4242 ( .A(n2242), .B(n2243), .Z(n2239) );
  AND U4243 ( .A(n2244), .B(n2245), .Z(n2242) );
  XNOR U4244 ( .A(x[1999]), .B(n2243), .Z(n2245) );
  XOR U4245 ( .A(n2246), .B(n2247), .Z(n2243) );
  AND U4246 ( .A(n2248), .B(n2249), .Z(n2246) );
  XNOR U4247 ( .A(x[1998]), .B(n2247), .Z(n2249) );
  XOR U4248 ( .A(n2250), .B(n2251), .Z(n2247) );
  AND U4249 ( .A(n2252), .B(n2253), .Z(n2250) );
  XNOR U4250 ( .A(x[1997]), .B(n2251), .Z(n2253) );
  XOR U4251 ( .A(n2254), .B(n2255), .Z(n2251) );
  AND U4252 ( .A(n2256), .B(n2257), .Z(n2254) );
  XNOR U4253 ( .A(x[1996]), .B(n2255), .Z(n2257) );
  XOR U4254 ( .A(n2258), .B(n2259), .Z(n2255) );
  AND U4255 ( .A(n2260), .B(n2261), .Z(n2258) );
  XNOR U4256 ( .A(x[1995]), .B(n2259), .Z(n2261) );
  XOR U4257 ( .A(n2262), .B(n2263), .Z(n2259) );
  AND U4258 ( .A(n2264), .B(n2265), .Z(n2262) );
  XNOR U4259 ( .A(x[1994]), .B(n2263), .Z(n2265) );
  XOR U4260 ( .A(n2266), .B(n2267), .Z(n2263) );
  AND U4261 ( .A(n2268), .B(n2269), .Z(n2266) );
  XNOR U4262 ( .A(x[1993]), .B(n2267), .Z(n2269) );
  XOR U4263 ( .A(n2270), .B(n2271), .Z(n2267) );
  AND U4264 ( .A(n2272), .B(n2273), .Z(n2270) );
  XNOR U4265 ( .A(x[1992]), .B(n2271), .Z(n2273) );
  XOR U4266 ( .A(n2274), .B(n2275), .Z(n2271) );
  AND U4267 ( .A(n2276), .B(n2277), .Z(n2274) );
  XNOR U4268 ( .A(x[1991]), .B(n2275), .Z(n2277) );
  XOR U4269 ( .A(n2278), .B(n2279), .Z(n2275) );
  AND U4270 ( .A(n2280), .B(n2281), .Z(n2278) );
  XNOR U4271 ( .A(x[1990]), .B(n2279), .Z(n2281) );
  XOR U4272 ( .A(n2282), .B(n2283), .Z(n2279) );
  AND U4273 ( .A(n2284), .B(n2285), .Z(n2282) );
  XNOR U4274 ( .A(x[1989]), .B(n2283), .Z(n2285) );
  XOR U4275 ( .A(n2286), .B(n2287), .Z(n2283) );
  AND U4276 ( .A(n2288), .B(n2289), .Z(n2286) );
  XNOR U4277 ( .A(x[1988]), .B(n2287), .Z(n2289) );
  XOR U4278 ( .A(n2290), .B(n2291), .Z(n2287) );
  AND U4279 ( .A(n2292), .B(n2293), .Z(n2290) );
  XNOR U4280 ( .A(x[1987]), .B(n2291), .Z(n2293) );
  XOR U4281 ( .A(n2294), .B(n2295), .Z(n2291) );
  AND U4282 ( .A(n2296), .B(n2297), .Z(n2294) );
  XNOR U4283 ( .A(x[1986]), .B(n2295), .Z(n2297) );
  XOR U4284 ( .A(n2298), .B(n2299), .Z(n2295) );
  AND U4285 ( .A(n2300), .B(n2301), .Z(n2298) );
  XNOR U4286 ( .A(x[1985]), .B(n2299), .Z(n2301) );
  XOR U4287 ( .A(n2302), .B(n2303), .Z(n2299) );
  AND U4288 ( .A(n2304), .B(n2305), .Z(n2302) );
  XNOR U4289 ( .A(x[1984]), .B(n2303), .Z(n2305) );
  XOR U4290 ( .A(n2306), .B(n2307), .Z(n2303) );
  AND U4291 ( .A(n2308), .B(n2309), .Z(n2306) );
  XNOR U4292 ( .A(x[1983]), .B(n2307), .Z(n2309) );
  XOR U4293 ( .A(n2310), .B(n2311), .Z(n2307) );
  AND U4294 ( .A(n2312), .B(n2313), .Z(n2310) );
  XNOR U4295 ( .A(x[1982]), .B(n2311), .Z(n2313) );
  XOR U4296 ( .A(n2314), .B(n2315), .Z(n2311) );
  AND U4297 ( .A(n2316), .B(n2317), .Z(n2314) );
  XNOR U4298 ( .A(x[1981]), .B(n2315), .Z(n2317) );
  XOR U4299 ( .A(n2318), .B(n2319), .Z(n2315) );
  AND U4300 ( .A(n2320), .B(n2321), .Z(n2318) );
  XNOR U4301 ( .A(x[1980]), .B(n2319), .Z(n2321) );
  XOR U4302 ( .A(n2322), .B(n2323), .Z(n2319) );
  AND U4303 ( .A(n2324), .B(n2325), .Z(n2322) );
  XNOR U4304 ( .A(x[1979]), .B(n2323), .Z(n2325) );
  XOR U4305 ( .A(n2326), .B(n2327), .Z(n2323) );
  AND U4306 ( .A(n2328), .B(n2329), .Z(n2326) );
  XNOR U4307 ( .A(x[1978]), .B(n2327), .Z(n2329) );
  XOR U4308 ( .A(n2330), .B(n2331), .Z(n2327) );
  AND U4309 ( .A(n2332), .B(n2333), .Z(n2330) );
  XNOR U4310 ( .A(x[1977]), .B(n2331), .Z(n2333) );
  XOR U4311 ( .A(n2334), .B(n2335), .Z(n2331) );
  AND U4312 ( .A(n2336), .B(n2337), .Z(n2334) );
  XNOR U4313 ( .A(x[1976]), .B(n2335), .Z(n2337) );
  XOR U4314 ( .A(n2338), .B(n2339), .Z(n2335) );
  AND U4315 ( .A(n2340), .B(n2341), .Z(n2338) );
  XNOR U4316 ( .A(x[1975]), .B(n2339), .Z(n2341) );
  XOR U4317 ( .A(n2342), .B(n2343), .Z(n2339) );
  AND U4318 ( .A(n2344), .B(n2345), .Z(n2342) );
  XNOR U4319 ( .A(x[1974]), .B(n2343), .Z(n2345) );
  XOR U4320 ( .A(n2346), .B(n2347), .Z(n2343) );
  AND U4321 ( .A(n2348), .B(n2349), .Z(n2346) );
  XNOR U4322 ( .A(x[1973]), .B(n2347), .Z(n2349) );
  XOR U4323 ( .A(n2350), .B(n2351), .Z(n2347) );
  AND U4324 ( .A(n2352), .B(n2353), .Z(n2350) );
  XNOR U4325 ( .A(x[1972]), .B(n2351), .Z(n2353) );
  XOR U4326 ( .A(n2354), .B(n2355), .Z(n2351) );
  AND U4327 ( .A(n2356), .B(n2357), .Z(n2354) );
  XNOR U4328 ( .A(x[1971]), .B(n2355), .Z(n2357) );
  XOR U4329 ( .A(n2358), .B(n2359), .Z(n2355) );
  AND U4330 ( .A(n2360), .B(n2361), .Z(n2358) );
  XNOR U4331 ( .A(x[1970]), .B(n2359), .Z(n2361) );
  XOR U4332 ( .A(n2362), .B(n2363), .Z(n2359) );
  AND U4333 ( .A(n2364), .B(n2365), .Z(n2362) );
  XNOR U4334 ( .A(x[1969]), .B(n2363), .Z(n2365) );
  XOR U4335 ( .A(n2366), .B(n2367), .Z(n2363) );
  AND U4336 ( .A(n2368), .B(n2369), .Z(n2366) );
  XNOR U4337 ( .A(x[1968]), .B(n2367), .Z(n2369) );
  XOR U4338 ( .A(n2370), .B(n2371), .Z(n2367) );
  AND U4339 ( .A(n2372), .B(n2373), .Z(n2370) );
  XNOR U4340 ( .A(x[1967]), .B(n2371), .Z(n2373) );
  XOR U4341 ( .A(n2374), .B(n2375), .Z(n2371) );
  AND U4342 ( .A(n2376), .B(n2377), .Z(n2374) );
  XNOR U4343 ( .A(x[1966]), .B(n2375), .Z(n2377) );
  XOR U4344 ( .A(n2378), .B(n2379), .Z(n2375) );
  AND U4345 ( .A(n2380), .B(n2381), .Z(n2378) );
  XNOR U4346 ( .A(x[1965]), .B(n2379), .Z(n2381) );
  XOR U4347 ( .A(n2382), .B(n2383), .Z(n2379) );
  AND U4348 ( .A(n2384), .B(n2385), .Z(n2382) );
  XNOR U4349 ( .A(x[1964]), .B(n2383), .Z(n2385) );
  XOR U4350 ( .A(n2386), .B(n2387), .Z(n2383) );
  AND U4351 ( .A(n2388), .B(n2389), .Z(n2386) );
  XNOR U4352 ( .A(x[1963]), .B(n2387), .Z(n2389) );
  XOR U4353 ( .A(n2390), .B(n2391), .Z(n2387) );
  AND U4354 ( .A(n2392), .B(n2393), .Z(n2390) );
  XNOR U4355 ( .A(x[1962]), .B(n2391), .Z(n2393) );
  XOR U4356 ( .A(n2394), .B(n2395), .Z(n2391) );
  AND U4357 ( .A(n2396), .B(n2397), .Z(n2394) );
  XNOR U4358 ( .A(x[1961]), .B(n2395), .Z(n2397) );
  XOR U4359 ( .A(n2398), .B(n2399), .Z(n2395) );
  AND U4360 ( .A(n2400), .B(n2401), .Z(n2398) );
  XNOR U4361 ( .A(x[1960]), .B(n2399), .Z(n2401) );
  XOR U4362 ( .A(n2402), .B(n2403), .Z(n2399) );
  AND U4363 ( .A(n2404), .B(n2405), .Z(n2402) );
  XNOR U4364 ( .A(x[1959]), .B(n2403), .Z(n2405) );
  XOR U4365 ( .A(n2406), .B(n2407), .Z(n2403) );
  AND U4366 ( .A(n2408), .B(n2409), .Z(n2406) );
  XNOR U4367 ( .A(x[1958]), .B(n2407), .Z(n2409) );
  XOR U4368 ( .A(n2410), .B(n2411), .Z(n2407) );
  AND U4369 ( .A(n2412), .B(n2413), .Z(n2410) );
  XNOR U4370 ( .A(x[1957]), .B(n2411), .Z(n2413) );
  XOR U4371 ( .A(n2414), .B(n2415), .Z(n2411) );
  AND U4372 ( .A(n2416), .B(n2417), .Z(n2414) );
  XNOR U4373 ( .A(x[1956]), .B(n2415), .Z(n2417) );
  XOR U4374 ( .A(n2418), .B(n2419), .Z(n2415) );
  AND U4375 ( .A(n2420), .B(n2421), .Z(n2418) );
  XNOR U4376 ( .A(x[1955]), .B(n2419), .Z(n2421) );
  XOR U4377 ( .A(n2422), .B(n2423), .Z(n2419) );
  AND U4378 ( .A(n2424), .B(n2425), .Z(n2422) );
  XNOR U4379 ( .A(x[1954]), .B(n2423), .Z(n2425) );
  XOR U4380 ( .A(n2426), .B(n2427), .Z(n2423) );
  AND U4381 ( .A(n2428), .B(n2429), .Z(n2426) );
  XNOR U4382 ( .A(x[1953]), .B(n2427), .Z(n2429) );
  XOR U4383 ( .A(n2430), .B(n2431), .Z(n2427) );
  AND U4384 ( .A(n2432), .B(n2433), .Z(n2430) );
  XNOR U4385 ( .A(x[1952]), .B(n2431), .Z(n2433) );
  XOR U4386 ( .A(n2434), .B(n2435), .Z(n2431) );
  AND U4387 ( .A(n2436), .B(n2437), .Z(n2434) );
  XNOR U4388 ( .A(x[1951]), .B(n2435), .Z(n2437) );
  XOR U4389 ( .A(n2438), .B(n2439), .Z(n2435) );
  AND U4390 ( .A(n2440), .B(n2441), .Z(n2438) );
  XNOR U4391 ( .A(x[1950]), .B(n2439), .Z(n2441) );
  XOR U4392 ( .A(n2442), .B(n2443), .Z(n2439) );
  AND U4393 ( .A(n2444), .B(n2445), .Z(n2442) );
  XNOR U4394 ( .A(x[1949]), .B(n2443), .Z(n2445) );
  XOR U4395 ( .A(n2446), .B(n2447), .Z(n2443) );
  AND U4396 ( .A(n2448), .B(n2449), .Z(n2446) );
  XNOR U4397 ( .A(x[1948]), .B(n2447), .Z(n2449) );
  XOR U4398 ( .A(n2450), .B(n2451), .Z(n2447) );
  AND U4399 ( .A(n2452), .B(n2453), .Z(n2450) );
  XNOR U4400 ( .A(x[1947]), .B(n2451), .Z(n2453) );
  XOR U4401 ( .A(n2454), .B(n2455), .Z(n2451) );
  AND U4402 ( .A(n2456), .B(n2457), .Z(n2454) );
  XNOR U4403 ( .A(x[1946]), .B(n2455), .Z(n2457) );
  XOR U4404 ( .A(n2458), .B(n2459), .Z(n2455) );
  AND U4405 ( .A(n2460), .B(n2461), .Z(n2458) );
  XNOR U4406 ( .A(x[1945]), .B(n2459), .Z(n2461) );
  XOR U4407 ( .A(n2462), .B(n2463), .Z(n2459) );
  AND U4408 ( .A(n2464), .B(n2465), .Z(n2462) );
  XNOR U4409 ( .A(x[1944]), .B(n2463), .Z(n2465) );
  XOR U4410 ( .A(n2466), .B(n2467), .Z(n2463) );
  AND U4411 ( .A(n2468), .B(n2469), .Z(n2466) );
  XNOR U4412 ( .A(x[1943]), .B(n2467), .Z(n2469) );
  XOR U4413 ( .A(n2470), .B(n2471), .Z(n2467) );
  AND U4414 ( .A(n2472), .B(n2473), .Z(n2470) );
  XNOR U4415 ( .A(x[1942]), .B(n2471), .Z(n2473) );
  XOR U4416 ( .A(n2474), .B(n2475), .Z(n2471) );
  AND U4417 ( .A(n2476), .B(n2477), .Z(n2474) );
  XNOR U4418 ( .A(x[1941]), .B(n2475), .Z(n2477) );
  XOR U4419 ( .A(n2478), .B(n2479), .Z(n2475) );
  AND U4420 ( .A(n2480), .B(n2481), .Z(n2478) );
  XNOR U4421 ( .A(x[1940]), .B(n2479), .Z(n2481) );
  XOR U4422 ( .A(n2482), .B(n2483), .Z(n2479) );
  AND U4423 ( .A(n2484), .B(n2485), .Z(n2482) );
  XNOR U4424 ( .A(x[1939]), .B(n2483), .Z(n2485) );
  XOR U4425 ( .A(n2486), .B(n2487), .Z(n2483) );
  AND U4426 ( .A(n2488), .B(n2489), .Z(n2486) );
  XNOR U4427 ( .A(x[1938]), .B(n2487), .Z(n2489) );
  XOR U4428 ( .A(n2490), .B(n2491), .Z(n2487) );
  AND U4429 ( .A(n2492), .B(n2493), .Z(n2490) );
  XNOR U4430 ( .A(x[1937]), .B(n2491), .Z(n2493) );
  XOR U4431 ( .A(n2494), .B(n2495), .Z(n2491) );
  AND U4432 ( .A(n2496), .B(n2497), .Z(n2494) );
  XNOR U4433 ( .A(x[1936]), .B(n2495), .Z(n2497) );
  XOR U4434 ( .A(n2498), .B(n2499), .Z(n2495) );
  AND U4435 ( .A(n2500), .B(n2501), .Z(n2498) );
  XNOR U4436 ( .A(x[1935]), .B(n2499), .Z(n2501) );
  XOR U4437 ( .A(n2502), .B(n2503), .Z(n2499) );
  AND U4438 ( .A(n2504), .B(n2505), .Z(n2502) );
  XNOR U4439 ( .A(x[1934]), .B(n2503), .Z(n2505) );
  XOR U4440 ( .A(n2506), .B(n2507), .Z(n2503) );
  AND U4441 ( .A(n2508), .B(n2509), .Z(n2506) );
  XNOR U4442 ( .A(x[1933]), .B(n2507), .Z(n2509) );
  XOR U4443 ( .A(n2510), .B(n2511), .Z(n2507) );
  AND U4444 ( .A(n2512), .B(n2513), .Z(n2510) );
  XNOR U4445 ( .A(x[1932]), .B(n2511), .Z(n2513) );
  XOR U4446 ( .A(n2514), .B(n2515), .Z(n2511) );
  AND U4447 ( .A(n2516), .B(n2517), .Z(n2514) );
  XNOR U4448 ( .A(x[1931]), .B(n2515), .Z(n2517) );
  XOR U4449 ( .A(n2518), .B(n2519), .Z(n2515) );
  AND U4450 ( .A(n2520), .B(n2521), .Z(n2518) );
  XNOR U4451 ( .A(x[1930]), .B(n2519), .Z(n2521) );
  XOR U4452 ( .A(n2522), .B(n2523), .Z(n2519) );
  AND U4453 ( .A(n2524), .B(n2525), .Z(n2522) );
  XNOR U4454 ( .A(x[1929]), .B(n2523), .Z(n2525) );
  XOR U4455 ( .A(n2526), .B(n2527), .Z(n2523) );
  AND U4456 ( .A(n2528), .B(n2529), .Z(n2526) );
  XNOR U4457 ( .A(x[1928]), .B(n2527), .Z(n2529) );
  XOR U4458 ( .A(n2530), .B(n2531), .Z(n2527) );
  AND U4459 ( .A(n2532), .B(n2533), .Z(n2530) );
  XNOR U4460 ( .A(x[1927]), .B(n2531), .Z(n2533) );
  XOR U4461 ( .A(n2534), .B(n2535), .Z(n2531) );
  AND U4462 ( .A(n2536), .B(n2537), .Z(n2534) );
  XNOR U4463 ( .A(x[1926]), .B(n2535), .Z(n2537) );
  XOR U4464 ( .A(n2538), .B(n2539), .Z(n2535) );
  AND U4465 ( .A(n2540), .B(n2541), .Z(n2538) );
  XNOR U4466 ( .A(x[1925]), .B(n2539), .Z(n2541) );
  XOR U4467 ( .A(n2542), .B(n2543), .Z(n2539) );
  AND U4468 ( .A(n2544), .B(n2545), .Z(n2542) );
  XNOR U4469 ( .A(x[1924]), .B(n2543), .Z(n2545) );
  XOR U4470 ( .A(n2546), .B(n2547), .Z(n2543) );
  AND U4471 ( .A(n2548), .B(n2549), .Z(n2546) );
  XNOR U4472 ( .A(x[1923]), .B(n2547), .Z(n2549) );
  XOR U4473 ( .A(n2550), .B(n2551), .Z(n2547) );
  AND U4474 ( .A(n2552), .B(n2553), .Z(n2550) );
  XNOR U4475 ( .A(x[1922]), .B(n2551), .Z(n2553) );
  XOR U4476 ( .A(n2554), .B(n2555), .Z(n2551) );
  AND U4477 ( .A(n2556), .B(n2557), .Z(n2554) );
  XNOR U4478 ( .A(x[1921]), .B(n2555), .Z(n2557) );
  XOR U4479 ( .A(n2558), .B(n2559), .Z(n2555) );
  AND U4480 ( .A(n2560), .B(n2561), .Z(n2558) );
  XNOR U4481 ( .A(x[1920]), .B(n2559), .Z(n2561) );
  XOR U4482 ( .A(n2562), .B(n2563), .Z(n2559) );
  AND U4483 ( .A(n2564), .B(n2565), .Z(n2562) );
  XNOR U4484 ( .A(x[1919]), .B(n2563), .Z(n2565) );
  XOR U4485 ( .A(n2566), .B(n2567), .Z(n2563) );
  AND U4486 ( .A(n2568), .B(n2569), .Z(n2566) );
  XNOR U4487 ( .A(x[1918]), .B(n2567), .Z(n2569) );
  XOR U4488 ( .A(n2570), .B(n2571), .Z(n2567) );
  AND U4489 ( .A(n2572), .B(n2573), .Z(n2570) );
  XNOR U4490 ( .A(x[1917]), .B(n2571), .Z(n2573) );
  XOR U4491 ( .A(n2574), .B(n2575), .Z(n2571) );
  AND U4492 ( .A(n2576), .B(n2577), .Z(n2574) );
  XNOR U4493 ( .A(x[1916]), .B(n2575), .Z(n2577) );
  XOR U4494 ( .A(n2578), .B(n2579), .Z(n2575) );
  AND U4495 ( .A(n2580), .B(n2581), .Z(n2578) );
  XNOR U4496 ( .A(x[1915]), .B(n2579), .Z(n2581) );
  XOR U4497 ( .A(n2582), .B(n2583), .Z(n2579) );
  AND U4498 ( .A(n2584), .B(n2585), .Z(n2582) );
  XNOR U4499 ( .A(x[1914]), .B(n2583), .Z(n2585) );
  XOR U4500 ( .A(n2586), .B(n2587), .Z(n2583) );
  AND U4501 ( .A(n2588), .B(n2589), .Z(n2586) );
  XNOR U4502 ( .A(x[1913]), .B(n2587), .Z(n2589) );
  XOR U4503 ( .A(n2590), .B(n2591), .Z(n2587) );
  AND U4504 ( .A(n2592), .B(n2593), .Z(n2590) );
  XNOR U4505 ( .A(x[1912]), .B(n2591), .Z(n2593) );
  XOR U4506 ( .A(n2594), .B(n2595), .Z(n2591) );
  AND U4507 ( .A(n2596), .B(n2597), .Z(n2594) );
  XNOR U4508 ( .A(x[1911]), .B(n2595), .Z(n2597) );
  XOR U4509 ( .A(n2598), .B(n2599), .Z(n2595) );
  AND U4510 ( .A(n2600), .B(n2601), .Z(n2598) );
  XNOR U4511 ( .A(x[1910]), .B(n2599), .Z(n2601) );
  XOR U4512 ( .A(n2602), .B(n2603), .Z(n2599) );
  AND U4513 ( .A(n2604), .B(n2605), .Z(n2602) );
  XNOR U4514 ( .A(x[1909]), .B(n2603), .Z(n2605) );
  XOR U4515 ( .A(n2606), .B(n2607), .Z(n2603) );
  AND U4516 ( .A(n2608), .B(n2609), .Z(n2606) );
  XNOR U4517 ( .A(x[1908]), .B(n2607), .Z(n2609) );
  XOR U4518 ( .A(n2610), .B(n2611), .Z(n2607) );
  AND U4519 ( .A(n2612), .B(n2613), .Z(n2610) );
  XNOR U4520 ( .A(x[1907]), .B(n2611), .Z(n2613) );
  XOR U4521 ( .A(n2614), .B(n2615), .Z(n2611) );
  AND U4522 ( .A(n2616), .B(n2617), .Z(n2614) );
  XNOR U4523 ( .A(x[1906]), .B(n2615), .Z(n2617) );
  XOR U4524 ( .A(n2618), .B(n2619), .Z(n2615) );
  AND U4525 ( .A(n2620), .B(n2621), .Z(n2618) );
  XNOR U4526 ( .A(x[1905]), .B(n2619), .Z(n2621) );
  XOR U4527 ( .A(n2622), .B(n2623), .Z(n2619) );
  AND U4528 ( .A(n2624), .B(n2625), .Z(n2622) );
  XNOR U4529 ( .A(x[1904]), .B(n2623), .Z(n2625) );
  XOR U4530 ( .A(n2626), .B(n2627), .Z(n2623) );
  AND U4531 ( .A(n2628), .B(n2629), .Z(n2626) );
  XNOR U4532 ( .A(x[1903]), .B(n2627), .Z(n2629) );
  XOR U4533 ( .A(n2630), .B(n2631), .Z(n2627) );
  AND U4534 ( .A(n2632), .B(n2633), .Z(n2630) );
  XNOR U4535 ( .A(x[1902]), .B(n2631), .Z(n2633) );
  XOR U4536 ( .A(n2634), .B(n2635), .Z(n2631) );
  AND U4537 ( .A(n2636), .B(n2637), .Z(n2634) );
  XNOR U4538 ( .A(x[1901]), .B(n2635), .Z(n2637) );
  XOR U4539 ( .A(n2638), .B(n2639), .Z(n2635) );
  AND U4540 ( .A(n2640), .B(n2641), .Z(n2638) );
  XNOR U4541 ( .A(x[1900]), .B(n2639), .Z(n2641) );
  XOR U4542 ( .A(n2642), .B(n2643), .Z(n2639) );
  AND U4543 ( .A(n2644), .B(n2645), .Z(n2642) );
  XNOR U4544 ( .A(x[1899]), .B(n2643), .Z(n2645) );
  XOR U4545 ( .A(n2646), .B(n2647), .Z(n2643) );
  AND U4546 ( .A(n2648), .B(n2649), .Z(n2646) );
  XNOR U4547 ( .A(x[1898]), .B(n2647), .Z(n2649) );
  XOR U4548 ( .A(n2650), .B(n2651), .Z(n2647) );
  AND U4549 ( .A(n2652), .B(n2653), .Z(n2650) );
  XNOR U4550 ( .A(x[1897]), .B(n2651), .Z(n2653) );
  XOR U4551 ( .A(n2654), .B(n2655), .Z(n2651) );
  AND U4552 ( .A(n2656), .B(n2657), .Z(n2654) );
  XNOR U4553 ( .A(x[1896]), .B(n2655), .Z(n2657) );
  XOR U4554 ( .A(n2658), .B(n2659), .Z(n2655) );
  AND U4555 ( .A(n2660), .B(n2661), .Z(n2658) );
  XNOR U4556 ( .A(x[1895]), .B(n2659), .Z(n2661) );
  XOR U4557 ( .A(n2662), .B(n2663), .Z(n2659) );
  AND U4558 ( .A(n2664), .B(n2665), .Z(n2662) );
  XNOR U4559 ( .A(x[1894]), .B(n2663), .Z(n2665) );
  XOR U4560 ( .A(n2666), .B(n2667), .Z(n2663) );
  AND U4561 ( .A(n2668), .B(n2669), .Z(n2666) );
  XNOR U4562 ( .A(x[1893]), .B(n2667), .Z(n2669) );
  XOR U4563 ( .A(n2670), .B(n2671), .Z(n2667) );
  AND U4564 ( .A(n2672), .B(n2673), .Z(n2670) );
  XNOR U4565 ( .A(x[1892]), .B(n2671), .Z(n2673) );
  XOR U4566 ( .A(n2674), .B(n2675), .Z(n2671) );
  AND U4567 ( .A(n2676), .B(n2677), .Z(n2674) );
  XNOR U4568 ( .A(x[1891]), .B(n2675), .Z(n2677) );
  XOR U4569 ( .A(n2678), .B(n2679), .Z(n2675) );
  AND U4570 ( .A(n2680), .B(n2681), .Z(n2678) );
  XNOR U4571 ( .A(x[1890]), .B(n2679), .Z(n2681) );
  XOR U4572 ( .A(n2682), .B(n2683), .Z(n2679) );
  AND U4573 ( .A(n2684), .B(n2685), .Z(n2682) );
  XNOR U4574 ( .A(x[1889]), .B(n2683), .Z(n2685) );
  XOR U4575 ( .A(n2686), .B(n2687), .Z(n2683) );
  AND U4576 ( .A(n2688), .B(n2689), .Z(n2686) );
  XNOR U4577 ( .A(x[1888]), .B(n2687), .Z(n2689) );
  XOR U4578 ( .A(n2690), .B(n2691), .Z(n2687) );
  AND U4579 ( .A(n2692), .B(n2693), .Z(n2690) );
  XNOR U4580 ( .A(x[1887]), .B(n2691), .Z(n2693) );
  XOR U4581 ( .A(n2694), .B(n2695), .Z(n2691) );
  AND U4582 ( .A(n2696), .B(n2697), .Z(n2694) );
  XNOR U4583 ( .A(x[1886]), .B(n2695), .Z(n2697) );
  XOR U4584 ( .A(n2698), .B(n2699), .Z(n2695) );
  AND U4585 ( .A(n2700), .B(n2701), .Z(n2698) );
  XNOR U4586 ( .A(x[1885]), .B(n2699), .Z(n2701) );
  XOR U4587 ( .A(n2702), .B(n2703), .Z(n2699) );
  AND U4588 ( .A(n2704), .B(n2705), .Z(n2702) );
  XNOR U4589 ( .A(x[1884]), .B(n2703), .Z(n2705) );
  XOR U4590 ( .A(n2706), .B(n2707), .Z(n2703) );
  AND U4591 ( .A(n2708), .B(n2709), .Z(n2706) );
  XNOR U4592 ( .A(x[1883]), .B(n2707), .Z(n2709) );
  XOR U4593 ( .A(n2710), .B(n2711), .Z(n2707) );
  AND U4594 ( .A(n2712), .B(n2713), .Z(n2710) );
  XNOR U4595 ( .A(x[1882]), .B(n2711), .Z(n2713) );
  XOR U4596 ( .A(n2714), .B(n2715), .Z(n2711) );
  AND U4597 ( .A(n2716), .B(n2717), .Z(n2714) );
  XNOR U4598 ( .A(x[1881]), .B(n2715), .Z(n2717) );
  XOR U4599 ( .A(n2718), .B(n2719), .Z(n2715) );
  AND U4600 ( .A(n2720), .B(n2721), .Z(n2718) );
  XNOR U4601 ( .A(x[1880]), .B(n2719), .Z(n2721) );
  XOR U4602 ( .A(n2722), .B(n2723), .Z(n2719) );
  AND U4603 ( .A(n2724), .B(n2725), .Z(n2722) );
  XNOR U4604 ( .A(x[1879]), .B(n2723), .Z(n2725) );
  XOR U4605 ( .A(n2726), .B(n2727), .Z(n2723) );
  AND U4606 ( .A(n2728), .B(n2729), .Z(n2726) );
  XNOR U4607 ( .A(x[1878]), .B(n2727), .Z(n2729) );
  XOR U4608 ( .A(n2730), .B(n2731), .Z(n2727) );
  AND U4609 ( .A(n2732), .B(n2733), .Z(n2730) );
  XNOR U4610 ( .A(x[1877]), .B(n2731), .Z(n2733) );
  XOR U4611 ( .A(n2734), .B(n2735), .Z(n2731) );
  AND U4612 ( .A(n2736), .B(n2737), .Z(n2734) );
  XNOR U4613 ( .A(x[1876]), .B(n2735), .Z(n2737) );
  XOR U4614 ( .A(n2738), .B(n2739), .Z(n2735) );
  AND U4615 ( .A(n2740), .B(n2741), .Z(n2738) );
  XNOR U4616 ( .A(x[1875]), .B(n2739), .Z(n2741) );
  XOR U4617 ( .A(n2742), .B(n2743), .Z(n2739) );
  AND U4618 ( .A(n2744), .B(n2745), .Z(n2742) );
  XNOR U4619 ( .A(x[1874]), .B(n2743), .Z(n2745) );
  XOR U4620 ( .A(n2746), .B(n2747), .Z(n2743) );
  AND U4621 ( .A(n2748), .B(n2749), .Z(n2746) );
  XNOR U4622 ( .A(x[1873]), .B(n2747), .Z(n2749) );
  XOR U4623 ( .A(n2750), .B(n2751), .Z(n2747) );
  AND U4624 ( .A(n2752), .B(n2753), .Z(n2750) );
  XNOR U4625 ( .A(x[1872]), .B(n2751), .Z(n2753) );
  XOR U4626 ( .A(n2754), .B(n2755), .Z(n2751) );
  AND U4627 ( .A(n2756), .B(n2757), .Z(n2754) );
  XNOR U4628 ( .A(x[1871]), .B(n2755), .Z(n2757) );
  XOR U4629 ( .A(n2758), .B(n2759), .Z(n2755) );
  AND U4630 ( .A(n2760), .B(n2761), .Z(n2758) );
  XNOR U4631 ( .A(x[1870]), .B(n2759), .Z(n2761) );
  XOR U4632 ( .A(n2762), .B(n2763), .Z(n2759) );
  AND U4633 ( .A(n2764), .B(n2765), .Z(n2762) );
  XNOR U4634 ( .A(x[1869]), .B(n2763), .Z(n2765) );
  XOR U4635 ( .A(n2766), .B(n2767), .Z(n2763) );
  AND U4636 ( .A(n2768), .B(n2769), .Z(n2766) );
  XNOR U4637 ( .A(x[1868]), .B(n2767), .Z(n2769) );
  XOR U4638 ( .A(n2770), .B(n2771), .Z(n2767) );
  AND U4639 ( .A(n2772), .B(n2773), .Z(n2770) );
  XNOR U4640 ( .A(x[1867]), .B(n2771), .Z(n2773) );
  XOR U4641 ( .A(n2774), .B(n2775), .Z(n2771) );
  AND U4642 ( .A(n2776), .B(n2777), .Z(n2774) );
  XNOR U4643 ( .A(x[1866]), .B(n2775), .Z(n2777) );
  XOR U4644 ( .A(n2778), .B(n2779), .Z(n2775) );
  AND U4645 ( .A(n2780), .B(n2781), .Z(n2778) );
  XNOR U4646 ( .A(x[1865]), .B(n2779), .Z(n2781) );
  XOR U4647 ( .A(n2782), .B(n2783), .Z(n2779) );
  AND U4648 ( .A(n2784), .B(n2785), .Z(n2782) );
  XNOR U4649 ( .A(x[1864]), .B(n2783), .Z(n2785) );
  XOR U4650 ( .A(n2786), .B(n2787), .Z(n2783) );
  AND U4651 ( .A(n2788), .B(n2789), .Z(n2786) );
  XNOR U4652 ( .A(x[1863]), .B(n2787), .Z(n2789) );
  XOR U4653 ( .A(n2790), .B(n2791), .Z(n2787) );
  AND U4654 ( .A(n2792), .B(n2793), .Z(n2790) );
  XNOR U4655 ( .A(x[1862]), .B(n2791), .Z(n2793) );
  XOR U4656 ( .A(n2794), .B(n2795), .Z(n2791) );
  AND U4657 ( .A(n2796), .B(n2797), .Z(n2794) );
  XNOR U4658 ( .A(x[1861]), .B(n2795), .Z(n2797) );
  XOR U4659 ( .A(n2798), .B(n2799), .Z(n2795) );
  AND U4660 ( .A(n2800), .B(n2801), .Z(n2798) );
  XNOR U4661 ( .A(x[1860]), .B(n2799), .Z(n2801) );
  XOR U4662 ( .A(n2802), .B(n2803), .Z(n2799) );
  AND U4663 ( .A(n2804), .B(n2805), .Z(n2802) );
  XNOR U4664 ( .A(x[1859]), .B(n2803), .Z(n2805) );
  XOR U4665 ( .A(n2806), .B(n2807), .Z(n2803) );
  AND U4666 ( .A(n2808), .B(n2809), .Z(n2806) );
  XNOR U4667 ( .A(x[1858]), .B(n2807), .Z(n2809) );
  XOR U4668 ( .A(n2810), .B(n2811), .Z(n2807) );
  AND U4669 ( .A(n2812), .B(n2813), .Z(n2810) );
  XNOR U4670 ( .A(x[1857]), .B(n2811), .Z(n2813) );
  XOR U4671 ( .A(n2814), .B(n2815), .Z(n2811) );
  AND U4672 ( .A(n2816), .B(n2817), .Z(n2814) );
  XNOR U4673 ( .A(x[1856]), .B(n2815), .Z(n2817) );
  XOR U4674 ( .A(n2818), .B(n2819), .Z(n2815) );
  AND U4675 ( .A(n2820), .B(n2821), .Z(n2818) );
  XNOR U4676 ( .A(x[1855]), .B(n2819), .Z(n2821) );
  XOR U4677 ( .A(n2822), .B(n2823), .Z(n2819) );
  AND U4678 ( .A(n2824), .B(n2825), .Z(n2822) );
  XNOR U4679 ( .A(x[1854]), .B(n2823), .Z(n2825) );
  XOR U4680 ( .A(n2826), .B(n2827), .Z(n2823) );
  AND U4681 ( .A(n2828), .B(n2829), .Z(n2826) );
  XNOR U4682 ( .A(x[1853]), .B(n2827), .Z(n2829) );
  XOR U4683 ( .A(n2830), .B(n2831), .Z(n2827) );
  AND U4684 ( .A(n2832), .B(n2833), .Z(n2830) );
  XNOR U4685 ( .A(x[1852]), .B(n2831), .Z(n2833) );
  XOR U4686 ( .A(n2834), .B(n2835), .Z(n2831) );
  AND U4687 ( .A(n2836), .B(n2837), .Z(n2834) );
  XNOR U4688 ( .A(x[1851]), .B(n2835), .Z(n2837) );
  XOR U4689 ( .A(n2838), .B(n2839), .Z(n2835) );
  AND U4690 ( .A(n2840), .B(n2841), .Z(n2838) );
  XNOR U4691 ( .A(x[1850]), .B(n2839), .Z(n2841) );
  XOR U4692 ( .A(n2842), .B(n2843), .Z(n2839) );
  AND U4693 ( .A(n2844), .B(n2845), .Z(n2842) );
  XNOR U4694 ( .A(x[1849]), .B(n2843), .Z(n2845) );
  XOR U4695 ( .A(n2846), .B(n2847), .Z(n2843) );
  AND U4696 ( .A(n2848), .B(n2849), .Z(n2846) );
  XNOR U4697 ( .A(x[1848]), .B(n2847), .Z(n2849) );
  XOR U4698 ( .A(n2850), .B(n2851), .Z(n2847) );
  AND U4699 ( .A(n2852), .B(n2853), .Z(n2850) );
  XNOR U4700 ( .A(x[1847]), .B(n2851), .Z(n2853) );
  XOR U4701 ( .A(n2854), .B(n2855), .Z(n2851) );
  AND U4702 ( .A(n2856), .B(n2857), .Z(n2854) );
  XNOR U4703 ( .A(x[1846]), .B(n2855), .Z(n2857) );
  XOR U4704 ( .A(n2858), .B(n2859), .Z(n2855) );
  AND U4705 ( .A(n2860), .B(n2861), .Z(n2858) );
  XNOR U4706 ( .A(x[1845]), .B(n2859), .Z(n2861) );
  XOR U4707 ( .A(n2862), .B(n2863), .Z(n2859) );
  AND U4708 ( .A(n2864), .B(n2865), .Z(n2862) );
  XNOR U4709 ( .A(x[1844]), .B(n2863), .Z(n2865) );
  XOR U4710 ( .A(n2866), .B(n2867), .Z(n2863) );
  AND U4711 ( .A(n2868), .B(n2869), .Z(n2866) );
  XNOR U4712 ( .A(x[1843]), .B(n2867), .Z(n2869) );
  XOR U4713 ( .A(n2870), .B(n2871), .Z(n2867) );
  AND U4714 ( .A(n2872), .B(n2873), .Z(n2870) );
  XNOR U4715 ( .A(x[1842]), .B(n2871), .Z(n2873) );
  XOR U4716 ( .A(n2874), .B(n2875), .Z(n2871) );
  AND U4717 ( .A(n2876), .B(n2877), .Z(n2874) );
  XNOR U4718 ( .A(x[1841]), .B(n2875), .Z(n2877) );
  XOR U4719 ( .A(n2878), .B(n2879), .Z(n2875) );
  AND U4720 ( .A(n2880), .B(n2881), .Z(n2878) );
  XNOR U4721 ( .A(x[1840]), .B(n2879), .Z(n2881) );
  XOR U4722 ( .A(n2882), .B(n2883), .Z(n2879) );
  AND U4723 ( .A(n2884), .B(n2885), .Z(n2882) );
  XNOR U4724 ( .A(x[1839]), .B(n2883), .Z(n2885) );
  XOR U4725 ( .A(n2886), .B(n2887), .Z(n2883) );
  AND U4726 ( .A(n2888), .B(n2889), .Z(n2886) );
  XNOR U4727 ( .A(x[1838]), .B(n2887), .Z(n2889) );
  XOR U4728 ( .A(n2890), .B(n2891), .Z(n2887) );
  AND U4729 ( .A(n2892), .B(n2893), .Z(n2890) );
  XNOR U4730 ( .A(x[1837]), .B(n2891), .Z(n2893) );
  XOR U4731 ( .A(n2894), .B(n2895), .Z(n2891) );
  AND U4732 ( .A(n2896), .B(n2897), .Z(n2894) );
  XNOR U4733 ( .A(x[1836]), .B(n2895), .Z(n2897) );
  XOR U4734 ( .A(n2898), .B(n2899), .Z(n2895) );
  AND U4735 ( .A(n2900), .B(n2901), .Z(n2898) );
  XNOR U4736 ( .A(x[1835]), .B(n2899), .Z(n2901) );
  XOR U4737 ( .A(n2902), .B(n2903), .Z(n2899) );
  AND U4738 ( .A(n2904), .B(n2905), .Z(n2902) );
  XNOR U4739 ( .A(x[1834]), .B(n2903), .Z(n2905) );
  XOR U4740 ( .A(n2906), .B(n2907), .Z(n2903) );
  AND U4741 ( .A(n2908), .B(n2909), .Z(n2906) );
  XNOR U4742 ( .A(x[1833]), .B(n2907), .Z(n2909) );
  XOR U4743 ( .A(n2910), .B(n2911), .Z(n2907) );
  AND U4744 ( .A(n2912), .B(n2913), .Z(n2910) );
  XNOR U4745 ( .A(x[1832]), .B(n2911), .Z(n2913) );
  XOR U4746 ( .A(n2914), .B(n2915), .Z(n2911) );
  AND U4747 ( .A(n2916), .B(n2917), .Z(n2914) );
  XNOR U4748 ( .A(x[1831]), .B(n2915), .Z(n2917) );
  XOR U4749 ( .A(n2918), .B(n2919), .Z(n2915) );
  AND U4750 ( .A(n2920), .B(n2921), .Z(n2918) );
  XNOR U4751 ( .A(x[1830]), .B(n2919), .Z(n2921) );
  XOR U4752 ( .A(n2922), .B(n2923), .Z(n2919) );
  AND U4753 ( .A(n2924), .B(n2925), .Z(n2922) );
  XNOR U4754 ( .A(x[1829]), .B(n2923), .Z(n2925) );
  XOR U4755 ( .A(n2926), .B(n2927), .Z(n2923) );
  AND U4756 ( .A(n2928), .B(n2929), .Z(n2926) );
  XNOR U4757 ( .A(x[1828]), .B(n2927), .Z(n2929) );
  XOR U4758 ( .A(n2930), .B(n2931), .Z(n2927) );
  AND U4759 ( .A(n2932), .B(n2933), .Z(n2930) );
  XNOR U4760 ( .A(x[1827]), .B(n2931), .Z(n2933) );
  XOR U4761 ( .A(n2934), .B(n2935), .Z(n2931) );
  AND U4762 ( .A(n2936), .B(n2937), .Z(n2934) );
  XNOR U4763 ( .A(x[1826]), .B(n2935), .Z(n2937) );
  XOR U4764 ( .A(n2938), .B(n2939), .Z(n2935) );
  AND U4765 ( .A(n2940), .B(n2941), .Z(n2938) );
  XNOR U4766 ( .A(x[1825]), .B(n2939), .Z(n2941) );
  XOR U4767 ( .A(n2942), .B(n2943), .Z(n2939) );
  AND U4768 ( .A(n2944), .B(n2945), .Z(n2942) );
  XNOR U4769 ( .A(x[1824]), .B(n2943), .Z(n2945) );
  XOR U4770 ( .A(n2946), .B(n2947), .Z(n2943) );
  AND U4771 ( .A(n2948), .B(n2949), .Z(n2946) );
  XNOR U4772 ( .A(x[1823]), .B(n2947), .Z(n2949) );
  XOR U4773 ( .A(n2950), .B(n2951), .Z(n2947) );
  AND U4774 ( .A(n2952), .B(n2953), .Z(n2950) );
  XNOR U4775 ( .A(x[1822]), .B(n2951), .Z(n2953) );
  XOR U4776 ( .A(n2954), .B(n2955), .Z(n2951) );
  AND U4777 ( .A(n2956), .B(n2957), .Z(n2954) );
  XNOR U4778 ( .A(x[1821]), .B(n2955), .Z(n2957) );
  XOR U4779 ( .A(n2958), .B(n2959), .Z(n2955) );
  AND U4780 ( .A(n2960), .B(n2961), .Z(n2958) );
  XNOR U4781 ( .A(x[1820]), .B(n2959), .Z(n2961) );
  XOR U4782 ( .A(n2962), .B(n2963), .Z(n2959) );
  AND U4783 ( .A(n2964), .B(n2965), .Z(n2962) );
  XNOR U4784 ( .A(x[1819]), .B(n2963), .Z(n2965) );
  XOR U4785 ( .A(n2966), .B(n2967), .Z(n2963) );
  AND U4786 ( .A(n2968), .B(n2969), .Z(n2966) );
  XNOR U4787 ( .A(x[1818]), .B(n2967), .Z(n2969) );
  XOR U4788 ( .A(n2970), .B(n2971), .Z(n2967) );
  AND U4789 ( .A(n2972), .B(n2973), .Z(n2970) );
  XNOR U4790 ( .A(x[1817]), .B(n2971), .Z(n2973) );
  XOR U4791 ( .A(n2974), .B(n2975), .Z(n2971) );
  AND U4792 ( .A(n2976), .B(n2977), .Z(n2974) );
  XNOR U4793 ( .A(x[1816]), .B(n2975), .Z(n2977) );
  XOR U4794 ( .A(n2978), .B(n2979), .Z(n2975) );
  AND U4795 ( .A(n2980), .B(n2981), .Z(n2978) );
  XNOR U4796 ( .A(x[1815]), .B(n2979), .Z(n2981) );
  XOR U4797 ( .A(n2982), .B(n2983), .Z(n2979) );
  AND U4798 ( .A(n2984), .B(n2985), .Z(n2982) );
  XNOR U4799 ( .A(x[1814]), .B(n2983), .Z(n2985) );
  XOR U4800 ( .A(n2986), .B(n2987), .Z(n2983) );
  AND U4801 ( .A(n2988), .B(n2989), .Z(n2986) );
  XNOR U4802 ( .A(x[1813]), .B(n2987), .Z(n2989) );
  XOR U4803 ( .A(n2990), .B(n2991), .Z(n2987) );
  AND U4804 ( .A(n2992), .B(n2993), .Z(n2990) );
  XNOR U4805 ( .A(x[1812]), .B(n2991), .Z(n2993) );
  XOR U4806 ( .A(n2994), .B(n2995), .Z(n2991) );
  AND U4807 ( .A(n2996), .B(n2997), .Z(n2994) );
  XNOR U4808 ( .A(x[1811]), .B(n2995), .Z(n2997) );
  XOR U4809 ( .A(n2998), .B(n2999), .Z(n2995) );
  AND U4810 ( .A(n3000), .B(n3001), .Z(n2998) );
  XNOR U4811 ( .A(x[1810]), .B(n2999), .Z(n3001) );
  XOR U4812 ( .A(n3002), .B(n3003), .Z(n2999) );
  AND U4813 ( .A(n3004), .B(n3005), .Z(n3002) );
  XNOR U4814 ( .A(x[1809]), .B(n3003), .Z(n3005) );
  XOR U4815 ( .A(n3006), .B(n3007), .Z(n3003) );
  AND U4816 ( .A(n3008), .B(n3009), .Z(n3006) );
  XNOR U4817 ( .A(x[1808]), .B(n3007), .Z(n3009) );
  XOR U4818 ( .A(n3010), .B(n3011), .Z(n3007) );
  AND U4819 ( .A(n3012), .B(n3013), .Z(n3010) );
  XNOR U4820 ( .A(x[1807]), .B(n3011), .Z(n3013) );
  XOR U4821 ( .A(n3014), .B(n3015), .Z(n3011) );
  AND U4822 ( .A(n3016), .B(n3017), .Z(n3014) );
  XNOR U4823 ( .A(x[1806]), .B(n3015), .Z(n3017) );
  XOR U4824 ( .A(n3018), .B(n3019), .Z(n3015) );
  AND U4825 ( .A(n3020), .B(n3021), .Z(n3018) );
  XNOR U4826 ( .A(x[1805]), .B(n3019), .Z(n3021) );
  XOR U4827 ( .A(n3022), .B(n3023), .Z(n3019) );
  AND U4828 ( .A(n3024), .B(n3025), .Z(n3022) );
  XNOR U4829 ( .A(x[1804]), .B(n3023), .Z(n3025) );
  XOR U4830 ( .A(n3026), .B(n3027), .Z(n3023) );
  AND U4831 ( .A(n3028), .B(n3029), .Z(n3026) );
  XNOR U4832 ( .A(x[1803]), .B(n3027), .Z(n3029) );
  XOR U4833 ( .A(n3030), .B(n3031), .Z(n3027) );
  AND U4834 ( .A(n3032), .B(n3033), .Z(n3030) );
  XNOR U4835 ( .A(x[1802]), .B(n3031), .Z(n3033) );
  XOR U4836 ( .A(n3034), .B(n3035), .Z(n3031) );
  AND U4837 ( .A(n3036), .B(n3037), .Z(n3034) );
  XNOR U4838 ( .A(x[1801]), .B(n3035), .Z(n3037) );
  XOR U4839 ( .A(n3038), .B(n3039), .Z(n3035) );
  AND U4840 ( .A(n3040), .B(n3041), .Z(n3038) );
  XNOR U4841 ( .A(x[1800]), .B(n3039), .Z(n3041) );
  XOR U4842 ( .A(n3042), .B(n3043), .Z(n3039) );
  AND U4843 ( .A(n3044), .B(n3045), .Z(n3042) );
  XNOR U4844 ( .A(x[1799]), .B(n3043), .Z(n3045) );
  XOR U4845 ( .A(n3046), .B(n3047), .Z(n3043) );
  AND U4846 ( .A(n3048), .B(n3049), .Z(n3046) );
  XNOR U4847 ( .A(x[1798]), .B(n3047), .Z(n3049) );
  XOR U4848 ( .A(n3050), .B(n3051), .Z(n3047) );
  AND U4849 ( .A(n3052), .B(n3053), .Z(n3050) );
  XNOR U4850 ( .A(x[1797]), .B(n3051), .Z(n3053) );
  XOR U4851 ( .A(n3054), .B(n3055), .Z(n3051) );
  AND U4852 ( .A(n3056), .B(n3057), .Z(n3054) );
  XNOR U4853 ( .A(x[1796]), .B(n3055), .Z(n3057) );
  XOR U4854 ( .A(n3058), .B(n3059), .Z(n3055) );
  AND U4855 ( .A(n3060), .B(n3061), .Z(n3058) );
  XNOR U4856 ( .A(x[1795]), .B(n3059), .Z(n3061) );
  XOR U4857 ( .A(n3062), .B(n3063), .Z(n3059) );
  AND U4858 ( .A(n3064), .B(n3065), .Z(n3062) );
  XNOR U4859 ( .A(x[1794]), .B(n3063), .Z(n3065) );
  XOR U4860 ( .A(n3066), .B(n3067), .Z(n3063) );
  AND U4861 ( .A(n3068), .B(n3069), .Z(n3066) );
  XNOR U4862 ( .A(x[1793]), .B(n3067), .Z(n3069) );
  XOR U4863 ( .A(n3070), .B(n3071), .Z(n3067) );
  AND U4864 ( .A(n3072), .B(n3073), .Z(n3070) );
  XNOR U4865 ( .A(x[1792]), .B(n3071), .Z(n3073) );
  XOR U4866 ( .A(n3074), .B(n3075), .Z(n3071) );
  AND U4867 ( .A(n3076), .B(n3077), .Z(n3074) );
  XNOR U4868 ( .A(x[1791]), .B(n3075), .Z(n3077) );
  XOR U4869 ( .A(n3078), .B(n3079), .Z(n3075) );
  AND U4870 ( .A(n3080), .B(n3081), .Z(n3078) );
  XNOR U4871 ( .A(x[1790]), .B(n3079), .Z(n3081) );
  XOR U4872 ( .A(n3082), .B(n3083), .Z(n3079) );
  AND U4873 ( .A(n3084), .B(n3085), .Z(n3082) );
  XNOR U4874 ( .A(x[1789]), .B(n3083), .Z(n3085) );
  XOR U4875 ( .A(n3086), .B(n3087), .Z(n3083) );
  AND U4876 ( .A(n3088), .B(n3089), .Z(n3086) );
  XNOR U4877 ( .A(x[1788]), .B(n3087), .Z(n3089) );
  XOR U4878 ( .A(n3090), .B(n3091), .Z(n3087) );
  AND U4879 ( .A(n3092), .B(n3093), .Z(n3090) );
  XNOR U4880 ( .A(x[1787]), .B(n3091), .Z(n3093) );
  XOR U4881 ( .A(n3094), .B(n3095), .Z(n3091) );
  AND U4882 ( .A(n3096), .B(n3097), .Z(n3094) );
  XNOR U4883 ( .A(x[1786]), .B(n3095), .Z(n3097) );
  XOR U4884 ( .A(n3098), .B(n3099), .Z(n3095) );
  AND U4885 ( .A(n3100), .B(n3101), .Z(n3098) );
  XNOR U4886 ( .A(x[1785]), .B(n3099), .Z(n3101) );
  XOR U4887 ( .A(n3102), .B(n3103), .Z(n3099) );
  AND U4888 ( .A(n3104), .B(n3105), .Z(n3102) );
  XNOR U4889 ( .A(x[1784]), .B(n3103), .Z(n3105) );
  XOR U4890 ( .A(n3106), .B(n3107), .Z(n3103) );
  AND U4891 ( .A(n3108), .B(n3109), .Z(n3106) );
  XNOR U4892 ( .A(x[1783]), .B(n3107), .Z(n3109) );
  XOR U4893 ( .A(n3110), .B(n3111), .Z(n3107) );
  AND U4894 ( .A(n3112), .B(n3113), .Z(n3110) );
  XNOR U4895 ( .A(x[1782]), .B(n3111), .Z(n3113) );
  XOR U4896 ( .A(n3114), .B(n3115), .Z(n3111) );
  AND U4897 ( .A(n3116), .B(n3117), .Z(n3114) );
  XNOR U4898 ( .A(x[1781]), .B(n3115), .Z(n3117) );
  XOR U4899 ( .A(n3118), .B(n3119), .Z(n3115) );
  AND U4900 ( .A(n3120), .B(n3121), .Z(n3118) );
  XNOR U4901 ( .A(x[1780]), .B(n3119), .Z(n3121) );
  XOR U4902 ( .A(n3122), .B(n3123), .Z(n3119) );
  AND U4903 ( .A(n3124), .B(n3125), .Z(n3122) );
  XNOR U4904 ( .A(x[1779]), .B(n3123), .Z(n3125) );
  XOR U4905 ( .A(n3126), .B(n3127), .Z(n3123) );
  AND U4906 ( .A(n3128), .B(n3129), .Z(n3126) );
  XNOR U4907 ( .A(x[1778]), .B(n3127), .Z(n3129) );
  XOR U4908 ( .A(n3130), .B(n3131), .Z(n3127) );
  AND U4909 ( .A(n3132), .B(n3133), .Z(n3130) );
  XNOR U4910 ( .A(x[1777]), .B(n3131), .Z(n3133) );
  XOR U4911 ( .A(n3134), .B(n3135), .Z(n3131) );
  AND U4912 ( .A(n3136), .B(n3137), .Z(n3134) );
  XNOR U4913 ( .A(x[1776]), .B(n3135), .Z(n3137) );
  XOR U4914 ( .A(n3138), .B(n3139), .Z(n3135) );
  AND U4915 ( .A(n3140), .B(n3141), .Z(n3138) );
  XNOR U4916 ( .A(x[1775]), .B(n3139), .Z(n3141) );
  XOR U4917 ( .A(n3142), .B(n3143), .Z(n3139) );
  AND U4918 ( .A(n3144), .B(n3145), .Z(n3142) );
  XNOR U4919 ( .A(x[1774]), .B(n3143), .Z(n3145) );
  XOR U4920 ( .A(n3146), .B(n3147), .Z(n3143) );
  AND U4921 ( .A(n3148), .B(n3149), .Z(n3146) );
  XNOR U4922 ( .A(x[1773]), .B(n3147), .Z(n3149) );
  XOR U4923 ( .A(n3150), .B(n3151), .Z(n3147) );
  AND U4924 ( .A(n3152), .B(n3153), .Z(n3150) );
  XNOR U4925 ( .A(x[1772]), .B(n3151), .Z(n3153) );
  XOR U4926 ( .A(n3154), .B(n3155), .Z(n3151) );
  AND U4927 ( .A(n3156), .B(n3157), .Z(n3154) );
  XNOR U4928 ( .A(x[1771]), .B(n3155), .Z(n3157) );
  XOR U4929 ( .A(n3158), .B(n3159), .Z(n3155) );
  AND U4930 ( .A(n3160), .B(n3161), .Z(n3158) );
  XNOR U4931 ( .A(x[1770]), .B(n3159), .Z(n3161) );
  XOR U4932 ( .A(n3162), .B(n3163), .Z(n3159) );
  AND U4933 ( .A(n3164), .B(n3165), .Z(n3162) );
  XNOR U4934 ( .A(x[1769]), .B(n3163), .Z(n3165) );
  XOR U4935 ( .A(n3166), .B(n3167), .Z(n3163) );
  AND U4936 ( .A(n3168), .B(n3169), .Z(n3166) );
  XNOR U4937 ( .A(x[1768]), .B(n3167), .Z(n3169) );
  XOR U4938 ( .A(n3170), .B(n3171), .Z(n3167) );
  AND U4939 ( .A(n3172), .B(n3173), .Z(n3170) );
  XNOR U4940 ( .A(x[1767]), .B(n3171), .Z(n3173) );
  XOR U4941 ( .A(n3174), .B(n3175), .Z(n3171) );
  AND U4942 ( .A(n3176), .B(n3177), .Z(n3174) );
  XNOR U4943 ( .A(x[1766]), .B(n3175), .Z(n3177) );
  XOR U4944 ( .A(n3178), .B(n3179), .Z(n3175) );
  AND U4945 ( .A(n3180), .B(n3181), .Z(n3178) );
  XNOR U4946 ( .A(x[1765]), .B(n3179), .Z(n3181) );
  XOR U4947 ( .A(n3182), .B(n3183), .Z(n3179) );
  AND U4948 ( .A(n3184), .B(n3185), .Z(n3182) );
  XNOR U4949 ( .A(x[1764]), .B(n3183), .Z(n3185) );
  XOR U4950 ( .A(n3186), .B(n3187), .Z(n3183) );
  AND U4951 ( .A(n3188), .B(n3189), .Z(n3186) );
  XNOR U4952 ( .A(x[1763]), .B(n3187), .Z(n3189) );
  XOR U4953 ( .A(n3190), .B(n3191), .Z(n3187) );
  AND U4954 ( .A(n3192), .B(n3193), .Z(n3190) );
  XNOR U4955 ( .A(x[1762]), .B(n3191), .Z(n3193) );
  XOR U4956 ( .A(n3194), .B(n3195), .Z(n3191) );
  AND U4957 ( .A(n3196), .B(n3197), .Z(n3194) );
  XNOR U4958 ( .A(x[1761]), .B(n3195), .Z(n3197) );
  XOR U4959 ( .A(n3198), .B(n3199), .Z(n3195) );
  AND U4960 ( .A(n3200), .B(n3201), .Z(n3198) );
  XNOR U4961 ( .A(x[1760]), .B(n3199), .Z(n3201) );
  XOR U4962 ( .A(n3202), .B(n3203), .Z(n3199) );
  AND U4963 ( .A(n3204), .B(n3205), .Z(n3202) );
  XNOR U4964 ( .A(x[1759]), .B(n3203), .Z(n3205) );
  XOR U4965 ( .A(n3206), .B(n3207), .Z(n3203) );
  AND U4966 ( .A(n3208), .B(n3209), .Z(n3206) );
  XNOR U4967 ( .A(x[1758]), .B(n3207), .Z(n3209) );
  XOR U4968 ( .A(n3210), .B(n3211), .Z(n3207) );
  AND U4969 ( .A(n3212), .B(n3213), .Z(n3210) );
  XNOR U4970 ( .A(x[1757]), .B(n3211), .Z(n3213) );
  XOR U4971 ( .A(n3214), .B(n3215), .Z(n3211) );
  AND U4972 ( .A(n3216), .B(n3217), .Z(n3214) );
  XNOR U4973 ( .A(x[1756]), .B(n3215), .Z(n3217) );
  XOR U4974 ( .A(n3218), .B(n3219), .Z(n3215) );
  AND U4975 ( .A(n3220), .B(n3221), .Z(n3218) );
  XNOR U4976 ( .A(x[1755]), .B(n3219), .Z(n3221) );
  XOR U4977 ( .A(n3222), .B(n3223), .Z(n3219) );
  AND U4978 ( .A(n3224), .B(n3225), .Z(n3222) );
  XNOR U4979 ( .A(x[1754]), .B(n3223), .Z(n3225) );
  XOR U4980 ( .A(n3226), .B(n3227), .Z(n3223) );
  AND U4981 ( .A(n3228), .B(n3229), .Z(n3226) );
  XNOR U4982 ( .A(x[1753]), .B(n3227), .Z(n3229) );
  XOR U4983 ( .A(n3230), .B(n3231), .Z(n3227) );
  AND U4984 ( .A(n3232), .B(n3233), .Z(n3230) );
  XNOR U4985 ( .A(x[1752]), .B(n3231), .Z(n3233) );
  XOR U4986 ( .A(n3234), .B(n3235), .Z(n3231) );
  AND U4987 ( .A(n3236), .B(n3237), .Z(n3234) );
  XNOR U4988 ( .A(x[1751]), .B(n3235), .Z(n3237) );
  XOR U4989 ( .A(n3238), .B(n3239), .Z(n3235) );
  AND U4990 ( .A(n3240), .B(n3241), .Z(n3238) );
  XNOR U4991 ( .A(x[1750]), .B(n3239), .Z(n3241) );
  XOR U4992 ( .A(n3242), .B(n3243), .Z(n3239) );
  AND U4993 ( .A(n3244), .B(n3245), .Z(n3242) );
  XNOR U4994 ( .A(x[1749]), .B(n3243), .Z(n3245) );
  XOR U4995 ( .A(n3246), .B(n3247), .Z(n3243) );
  AND U4996 ( .A(n3248), .B(n3249), .Z(n3246) );
  XNOR U4997 ( .A(x[1748]), .B(n3247), .Z(n3249) );
  XOR U4998 ( .A(n3250), .B(n3251), .Z(n3247) );
  AND U4999 ( .A(n3252), .B(n3253), .Z(n3250) );
  XNOR U5000 ( .A(x[1747]), .B(n3251), .Z(n3253) );
  XOR U5001 ( .A(n3254), .B(n3255), .Z(n3251) );
  AND U5002 ( .A(n3256), .B(n3257), .Z(n3254) );
  XNOR U5003 ( .A(x[1746]), .B(n3255), .Z(n3257) );
  XOR U5004 ( .A(n3258), .B(n3259), .Z(n3255) );
  AND U5005 ( .A(n3260), .B(n3261), .Z(n3258) );
  XNOR U5006 ( .A(x[1745]), .B(n3259), .Z(n3261) );
  XOR U5007 ( .A(n3262), .B(n3263), .Z(n3259) );
  AND U5008 ( .A(n3264), .B(n3265), .Z(n3262) );
  XNOR U5009 ( .A(x[1744]), .B(n3263), .Z(n3265) );
  XOR U5010 ( .A(n3266), .B(n3267), .Z(n3263) );
  AND U5011 ( .A(n3268), .B(n3269), .Z(n3266) );
  XNOR U5012 ( .A(x[1743]), .B(n3267), .Z(n3269) );
  XOR U5013 ( .A(n3270), .B(n3271), .Z(n3267) );
  AND U5014 ( .A(n3272), .B(n3273), .Z(n3270) );
  XNOR U5015 ( .A(x[1742]), .B(n3271), .Z(n3273) );
  XOR U5016 ( .A(n3274), .B(n3275), .Z(n3271) );
  AND U5017 ( .A(n3276), .B(n3277), .Z(n3274) );
  XNOR U5018 ( .A(x[1741]), .B(n3275), .Z(n3277) );
  XOR U5019 ( .A(n3278), .B(n3279), .Z(n3275) );
  AND U5020 ( .A(n3280), .B(n3281), .Z(n3278) );
  XNOR U5021 ( .A(x[1740]), .B(n3279), .Z(n3281) );
  XOR U5022 ( .A(n3282), .B(n3283), .Z(n3279) );
  AND U5023 ( .A(n3284), .B(n3285), .Z(n3282) );
  XNOR U5024 ( .A(x[1739]), .B(n3283), .Z(n3285) );
  XOR U5025 ( .A(n3286), .B(n3287), .Z(n3283) );
  AND U5026 ( .A(n3288), .B(n3289), .Z(n3286) );
  XNOR U5027 ( .A(x[1738]), .B(n3287), .Z(n3289) );
  XOR U5028 ( .A(n3290), .B(n3291), .Z(n3287) );
  AND U5029 ( .A(n3292), .B(n3293), .Z(n3290) );
  XNOR U5030 ( .A(x[1737]), .B(n3291), .Z(n3293) );
  XOR U5031 ( .A(n3294), .B(n3295), .Z(n3291) );
  AND U5032 ( .A(n3296), .B(n3297), .Z(n3294) );
  XNOR U5033 ( .A(x[1736]), .B(n3295), .Z(n3297) );
  XOR U5034 ( .A(n3298), .B(n3299), .Z(n3295) );
  AND U5035 ( .A(n3300), .B(n3301), .Z(n3298) );
  XNOR U5036 ( .A(x[1735]), .B(n3299), .Z(n3301) );
  XOR U5037 ( .A(n3302), .B(n3303), .Z(n3299) );
  AND U5038 ( .A(n3304), .B(n3305), .Z(n3302) );
  XNOR U5039 ( .A(x[1734]), .B(n3303), .Z(n3305) );
  XOR U5040 ( .A(n3306), .B(n3307), .Z(n3303) );
  AND U5041 ( .A(n3308), .B(n3309), .Z(n3306) );
  XNOR U5042 ( .A(x[1733]), .B(n3307), .Z(n3309) );
  XOR U5043 ( .A(n3310), .B(n3311), .Z(n3307) );
  AND U5044 ( .A(n3312), .B(n3313), .Z(n3310) );
  XNOR U5045 ( .A(x[1732]), .B(n3311), .Z(n3313) );
  XOR U5046 ( .A(n3314), .B(n3315), .Z(n3311) );
  AND U5047 ( .A(n3316), .B(n3317), .Z(n3314) );
  XNOR U5048 ( .A(x[1731]), .B(n3315), .Z(n3317) );
  XOR U5049 ( .A(n3318), .B(n3319), .Z(n3315) );
  AND U5050 ( .A(n3320), .B(n3321), .Z(n3318) );
  XNOR U5051 ( .A(x[1730]), .B(n3319), .Z(n3321) );
  XOR U5052 ( .A(n3322), .B(n3323), .Z(n3319) );
  AND U5053 ( .A(n3324), .B(n3325), .Z(n3322) );
  XNOR U5054 ( .A(x[1729]), .B(n3323), .Z(n3325) );
  XOR U5055 ( .A(n3326), .B(n3327), .Z(n3323) );
  AND U5056 ( .A(n3328), .B(n3329), .Z(n3326) );
  XNOR U5057 ( .A(x[1728]), .B(n3327), .Z(n3329) );
  XOR U5058 ( .A(n3330), .B(n3331), .Z(n3327) );
  AND U5059 ( .A(n3332), .B(n3333), .Z(n3330) );
  XNOR U5060 ( .A(x[1727]), .B(n3331), .Z(n3333) );
  XOR U5061 ( .A(n3334), .B(n3335), .Z(n3331) );
  AND U5062 ( .A(n3336), .B(n3337), .Z(n3334) );
  XNOR U5063 ( .A(x[1726]), .B(n3335), .Z(n3337) );
  XOR U5064 ( .A(n3338), .B(n3339), .Z(n3335) );
  AND U5065 ( .A(n3340), .B(n3341), .Z(n3338) );
  XNOR U5066 ( .A(x[1725]), .B(n3339), .Z(n3341) );
  XOR U5067 ( .A(n3342), .B(n3343), .Z(n3339) );
  AND U5068 ( .A(n3344), .B(n3345), .Z(n3342) );
  XNOR U5069 ( .A(x[1724]), .B(n3343), .Z(n3345) );
  XOR U5070 ( .A(n3346), .B(n3347), .Z(n3343) );
  AND U5071 ( .A(n3348), .B(n3349), .Z(n3346) );
  XNOR U5072 ( .A(x[1723]), .B(n3347), .Z(n3349) );
  XOR U5073 ( .A(n3350), .B(n3351), .Z(n3347) );
  AND U5074 ( .A(n3352), .B(n3353), .Z(n3350) );
  XNOR U5075 ( .A(x[1722]), .B(n3351), .Z(n3353) );
  XOR U5076 ( .A(n3354), .B(n3355), .Z(n3351) );
  AND U5077 ( .A(n3356), .B(n3357), .Z(n3354) );
  XNOR U5078 ( .A(x[1721]), .B(n3355), .Z(n3357) );
  XOR U5079 ( .A(n3358), .B(n3359), .Z(n3355) );
  AND U5080 ( .A(n3360), .B(n3361), .Z(n3358) );
  XNOR U5081 ( .A(x[1720]), .B(n3359), .Z(n3361) );
  XOR U5082 ( .A(n3362), .B(n3363), .Z(n3359) );
  AND U5083 ( .A(n3364), .B(n3365), .Z(n3362) );
  XNOR U5084 ( .A(x[1719]), .B(n3363), .Z(n3365) );
  XOR U5085 ( .A(n3366), .B(n3367), .Z(n3363) );
  AND U5086 ( .A(n3368), .B(n3369), .Z(n3366) );
  XNOR U5087 ( .A(x[1718]), .B(n3367), .Z(n3369) );
  XOR U5088 ( .A(n3370), .B(n3371), .Z(n3367) );
  AND U5089 ( .A(n3372), .B(n3373), .Z(n3370) );
  XNOR U5090 ( .A(x[1717]), .B(n3371), .Z(n3373) );
  XOR U5091 ( .A(n3374), .B(n3375), .Z(n3371) );
  AND U5092 ( .A(n3376), .B(n3377), .Z(n3374) );
  XNOR U5093 ( .A(x[1716]), .B(n3375), .Z(n3377) );
  XOR U5094 ( .A(n3378), .B(n3379), .Z(n3375) );
  AND U5095 ( .A(n3380), .B(n3381), .Z(n3378) );
  XNOR U5096 ( .A(x[1715]), .B(n3379), .Z(n3381) );
  XOR U5097 ( .A(n3382), .B(n3383), .Z(n3379) );
  AND U5098 ( .A(n3384), .B(n3385), .Z(n3382) );
  XNOR U5099 ( .A(x[1714]), .B(n3383), .Z(n3385) );
  XOR U5100 ( .A(n3386), .B(n3387), .Z(n3383) );
  AND U5101 ( .A(n3388), .B(n3389), .Z(n3386) );
  XNOR U5102 ( .A(x[1713]), .B(n3387), .Z(n3389) );
  XOR U5103 ( .A(n3390), .B(n3391), .Z(n3387) );
  AND U5104 ( .A(n3392), .B(n3393), .Z(n3390) );
  XNOR U5105 ( .A(x[1712]), .B(n3391), .Z(n3393) );
  XOR U5106 ( .A(n3394), .B(n3395), .Z(n3391) );
  AND U5107 ( .A(n3396), .B(n3397), .Z(n3394) );
  XNOR U5108 ( .A(x[1711]), .B(n3395), .Z(n3397) );
  XOR U5109 ( .A(n3398), .B(n3399), .Z(n3395) );
  AND U5110 ( .A(n3400), .B(n3401), .Z(n3398) );
  XNOR U5111 ( .A(x[1710]), .B(n3399), .Z(n3401) );
  XOR U5112 ( .A(n3402), .B(n3403), .Z(n3399) );
  AND U5113 ( .A(n3404), .B(n3405), .Z(n3402) );
  XNOR U5114 ( .A(x[1709]), .B(n3403), .Z(n3405) );
  XOR U5115 ( .A(n3406), .B(n3407), .Z(n3403) );
  AND U5116 ( .A(n3408), .B(n3409), .Z(n3406) );
  XNOR U5117 ( .A(x[1708]), .B(n3407), .Z(n3409) );
  XOR U5118 ( .A(n3410), .B(n3411), .Z(n3407) );
  AND U5119 ( .A(n3412), .B(n3413), .Z(n3410) );
  XNOR U5120 ( .A(x[1707]), .B(n3411), .Z(n3413) );
  XOR U5121 ( .A(n3414), .B(n3415), .Z(n3411) );
  AND U5122 ( .A(n3416), .B(n3417), .Z(n3414) );
  XNOR U5123 ( .A(x[1706]), .B(n3415), .Z(n3417) );
  XOR U5124 ( .A(n3418), .B(n3419), .Z(n3415) );
  AND U5125 ( .A(n3420), .B(n3421), .Z(n3418) );
  XNOR U5126 ( .A(x[1705]), .B(n3419), .Z(n3421) );
  XOR U5127 ( .A(n3422), .B(n3423), .Z(n3419) );
  AND U5128 ( .A(n3424), .B(n3425), .Z(n3422) );
  XNOR U5129 ( .A(x[1704]), .B(n3423), .Z(n3425) );
  XOR U5130 ( .A(n3426), .B(n3427), .Z(n3423) );
  AND U5131 ( .A(n3428), .B(n3429), .Z(n3426) );
  XNOR U5132 ( .A(x[1703]), .B(n3427), .Z(n3429) );
  XOR U5133 ( .A(n3430), .B(n3431), .Z(n3427) );
  AND U5134 ( .A(n3432), .B(n3433), .Z(n3430) );
  XNOR U5135 ( .A(x[1702]), .B(n3431), .Z(n3433) );
  XOR U5136 ( .A(n3434), .B(n3435), .Z(n3431) );
  AND U5137 ( .A(n3436), .B(n3437), .Z(n3434) );
  XNOR U5138 ( .A(x[1701]), .B(n3435), .Z(n3437) );
  XOR U5139 ( .A(n3438), .B(n3439), .Z(n3435) );
  AND U5140 ( .A(n3440), .B(n3441), .Z(n3438) );
  XNOR U5141 ( .A(x[1700]), .B(n3439), .Z(n3441) );
  XOR U5142 ( .A(n3442), .B(n3443), .Z(n3439) );
  AND U5143 ( .A(n3444), .B(n3445), .Z(n3442) );
  XNOR U5144 ( .A(x[1699]), .B(n3443), .Z(n3445) );
  XOR U5145 ( .A(n3446), .B(n3447), .Z(n3443) );
  AND U5146 ( .A(n3448), .B(n3449), .Z(n3446) );
  XNOR U5147 ( .A(x[1698]), .B(n3447), .Z(n3449) );
  XOR U5148 ( .A(n3450), .B(n3451), .Z(n3447) );
  AND U5149 ( .A(n3452), .B(n3453), .Z(n3450) );
  XNOR U5150 ( .A(x[1697]), .B(n3451), .Z(n3453) );
  XOR U5151 ( .A(n3454), .B(n3455), .Z(n3451) );
  AND U5152 ( .A(n3456), .B(n3457), .Z(n3454) );
  XNOR U5153 ( .A(x[1696]), .B(n3455), .Z(n3457) );
  XOR U5154 ( .A(n3458), .B(n3459), .Z(n3455) );
  AND U5155 ( .A(n3460), .B(n3461), .Z(n3458) );
  XNOR U5156 ( .A(x[1695]), .B(n3459), .Z(n3461) );
  XOR U5157 ( .A(n3462), .B(n3463), .Z(n3459) );
  AND U5158 ( .A(n3464), .B(n3465), .Z(n3462) );
  XNOR U5159 ( .A(x[1694]), .B(n3463), .Z(n3465) );
  XOR U5160 ( .A(n3466), .B(n3467), .Z(n3463) );
  AND U5161 ( .A(n3468), .B(n3469), .Z(n3466) );
  XNOR U5162 ( .A(x[1693]), .B(n3467), .Z(n3469) );
  XOR U5163 ( .A(n3470), .B(n3471), .Z(n3467) );
  AND U5164 ( .A(n3472), .B(n3473), .Z(n3470) );
  XNOR U5165 ( .A(x[1692]), .B(n3471), .Z(n3473) );
  XOR U5166 ( .A(n3474), .B(n3475), .Z(n3471) );
  AND U5167 ( .A(n3476), .B(n3477), .Z(n3474) );
  XNOR U5168 ( .A(x[1691]), .B(n3475), .Z(n3477) );
  XOR U5169 ( .A(n3478), .B(n3479), .Z(n3475) );
  AND U5170 ( .A(n3480), .B(n3481), .Z(n3478) );
  XNOR U5171 ( .A(x[1690]), .B(n3479), .Z(n3481) );
  XOR U5172 ( .A(n3482), .B(n3483), .Z(n3479) );
  AND U5173 ( .A(n3484), .B(n3485), .Z(n3482) );
  XNOR U5174 ( .A(x[1689]), .B(n3483), .Z(n3485) );
  XOR U5175 ( .A(n3486), .B(n3487), .Z(n3483) );
  AND U5176 ( .A(n3488), .B(n3489), .Z(n3486) );
  XNOR U5177 ( .A(x[1688]), .B(n3487), .Z(n3489) );
  XOR U5178 ( .A(n3490), .B(n3491), .Z(n3487) );
  AND U5179 ( .A(n3492), .B(n3493), .Z(n3490) );
  XNOR U5180 ( .A(x[1687]), .B(n3491), .Z(n3493) );
  XOR U5181 ( .A(n3494), .B(n3495), .Z(n3491) );
  AND U5182 ( .A(n3496), .B(n3497), .Z(n3494) );
  XNOR U5183 ( .A(x[1686]), .B(n3495), .Z(n3497) );
  XOR U5184 ( .A(n3498), .B(n3499), .Z(n3495) );
  AND U5185 ( .A(n3500), .B(n3501), .Z(n3498) );
  XNOR U5186 ( .A(x[1685]), .B(n3499), .Z(n3501) );
  XOR U5187 ( .A(n3502), .B(n3503), .Z(n3499) );
  AND U5188 ( .A(n3504), .B(n3505), .Z(n3502) );
  XNOR U5189 ( .A(x[1684]), .B(n3503), .Z(n3505) );
  XOR U5190 ( .A(n3506), .B(n3507), .Z(n3503) );
  AND U5191 ( .A(n3508), .B(n3509), .Z(n3506) );
  XNOR U5192 ( .A(x[1683]), .B(n3507), .Z(n3509) );
  XOR U5193 ( .A(n3510), .B(n3511), .Z(n3507) );
  AND U5194 ( .A(n3512), .B(n3513), .Z(n3510) );
  XNOR U5195 ( .A(x[1682]), .B(n3511), .Z(n3513) );
  XOR U5196 ( .A(n3514), .B(n3515), .Z(n3511) );
  AND U5197 ( .A(n3516), .B(n3517), .Z(n3514) );
  XNOR U5198 ( .A(x[1681]), .B(n3515), .Z(n3517) );
  XOR U5199 ( .A(n3518), .B(n3519), .Z(n3515) );
  AND U5200 ( .A(n3520), .B(n3521), .Z(n3518) );
  XNOR U5201 ( .A(x[1680]), .B(n3519), .Z(n3521) );
  XOR U5202 ( .A(n3522), .B(n3523), .Z(n3519) );
  AND U5203 ( .A(n3524), .B(n3525), .Z(n3522) );
  XNOR U5204 ( .A(x[1679]), .B(n3523), .Z(n3525) );
  XOR U5205 ( .A(n3526), .B(n3527), .Z(n3523) );
  AND U5206 ( .A(n3528), .B(n3529), .Z(n3526) );
  XNOR U5207 ( .A(x[1678]), .B(n3527), .Z(n3529) );
  XOR U5208 ( .A(n3530), .B(n3531), .Z(n3527) );
  AND U5209 ( .A(n3532), .B(n3533), .Z(n3530) );
  XNOR U5210 ( .A(x[1677]), .B(n3531), .Z(n3533) );
  XOR U5211 ( .A(n3534), .B(n3535), .Z(n3531) );
  AND U5212 ( .A(n3536), .B(n3537), .Z(n3534) );
  XNOR U5213 ( .A(x[1676]), .B(n3535), .Z(n3537) );
  XOR U5214 ( .A(n3538), .B(n3539), .Z(n3535) );
  AND U5215 ( .A(n3540), .B(n3541), .Z(n3538) );
  XNOR U5216 ( .A(x[1675]), .B(n3539), .Z(n3541) );
  XOR U5217 ( .A(n3542), .B(n3543), .Z(n3539) );
  AND U5218 ( .A(n3544), .B(n3545), .Z(n3542) );
  XNOR U5219 ( .A(x[1674]), .B(n3543), .Z(n3545) );
  XOR U5220 ( .A(n3546), .B(n3547), .Z(n3543) );
  AND U5221 ( .A(n3548), .B(n3549), .Z(n3546) );
  XNOR U5222 ( .A(x[1673]), .B(n3547), .Z(n3549) );
  XOR U5223 ( .A(n3550), .B(n3551), .Z(n3547) );
  AND U5224 ( .A(n3552), .B(n3553), .Z(n3550) );
  XNOR U5225 ( .A(x[1672]), .B(n3551), .Z(n3553) );
  XOR U5226 ( .A(n3554), .B(n3555), .Z(n3551) );
  AND U5227 ( .A(n3556), .B(n3557), .Z(n3554) );
  XNOR U5228 ( .A(x[1671]), .B(n3555), .Z(n3557) );
  XOR U5229 ( .A(n3558), .B(n3559), .Z(n3555) );
  AND U5230 ( .A(n3560), .B(n3561), .Z(n3558) );
  XNOR U5231 ( .A(x[1670]), .B(n3559), .Z(n3561) );
  XOR U5232 ( .A(n3562), .B(n3563), .Z(n3559) );
  AND U5233 ( .A(n3564), .B(n3565), .Z(n3562) );
  XNOR U5234 ( .A(x[1669]), .B(n3563), .Z(n3565) );
  XOR U5235 ( .A(n3566), .B(n3567), .Z(n3563) );
  AND U5236 ( .A(n3568), .B(n3569), .Z(n3566) );
  XNOR U5237 ( .A(x[1668]), .B(n3567), .Z(n3569) );
  XOR U5238 ( .A(n3570), .B(n3571), .Z(n3567) );
  AND U5239 ( .A(n3572), .B(n3573), .Z(n3570) );
  XNOR U5240 ( .A(x[1667]), .B(n3571), .Z(n3573) );
  XOR U5241 ( .A(n3574), .B(n3575), .Z(n3571) );
  AND U5242 ( .A(n3576), .B(n3577), .Z(n3574) );
  XNOR U5243 ( .A(x[1666]), .B(n3575), .Z(n3577) );
  XOR U5244 ( .A(n3578), .B(n3579), .Z(n3575) );
  AND U5245 ( .A(n3580), .B(n3581), .Z(n3578) );
  XNOR U5246 ( .A(x[1665]), .B(n3579), .Z(n3581) );
  XOR U5247 ( .A(n3582), .B(n3583), .Z(n3579) );
  AND U5248 ( .A(n3584), .B(n3585), .Z(n3582) );
  XNOR U5249 ( .A(x[1664]), .B(n3583), .Z(n3585) );
  XOR U5250 ( .A(n3586), .B(n3587), .Z(n3583) );
  AND U5251 ( .A(n3588), .B(n3589), .Z(n3586) );
  XNOR U5252 ( .A(x[1663]), .B(n3587), .Z(n3589) );
  XOR U5253 ( .A(n3590), .B(n3591), .Z(n3587) );
  AND U5254 ( .A(n3592), .B(n3593), .Z(n3590) );
  XNOR U5255 ( .A(x[1662]), .B(n3591), .Z(n3593) );
  XOR U5256 ( .A(n3594), .B(n3595), .Z(n3591) );
  AND U5257 ( .A(n3596), .B(n3597), .Z(n3594) );
  XNOR U5258 ( .A(x[1661]), .B(n3595), .Z(n3597) );
  XOR U5259 ( .A(n3598), .B(n3599), .Z(n3595) );
  AND U5260 ( .A(n3600), .B(n3601), .Z(n3598) );
  XNOR U5261 ( .A(x[1660]), .B(n3599), .Z(n3601) );
  XOR U5262 ( .A(n3602), .B(n3603), .Z(n3599) );
  AND U5263 ( .A(n3604), .B(n3605), .Z(n3602) );
  XNOR U5264 ( .A(x[1659]), .B(n3603), .Z(n3605) );
  XOR U5265 ( .A(n3606), .B(n3607), .Z(n3603) );
  AND U5266 ( .A(n3608), .B(n3609), .Z(n3606) );
  XNOR U5267 ( .A(x[1658]), .B(n3607), .Z(n3609) );
  XOR U5268 ( .A(n3610), .B(n3611), .Z(n3607) );
  AND U5269 ( .A(n3612), .B(n3613), .Z(n3610) );
  XNOR U5270 ( .A(x[1657]), .B(n3611), .Z(n3613) );
  XOR U5271 ( .A(n3614), .B(n3615), .Z(n3611) );
  AND U5272 ( .A(n3616), .B(n3617), .Z(n3614) );
  XNOR U5273 ( .A(x[1656]), .B(n3615), .Z(n3617) );
  XOR U5274 ( .A(n3618), .B(n3619), .Z(n3615) );
  AND U5275 ( .A(n3620), .B(n3621), .Z(n3618) );
  XNOR U5276 ( .A(x[1655]), .B(n3619), .Z(n3621) );
  XOR U5277 ( .A(n3622), .B(n3623), .Z(n3619) );
  AND U5278 ( .A(n3624), .B(n3625), .Z(n3622) );
  XNOR U5279 ( .A(x[1654]), .B(n3623), .Z(n3625) );
  XOR U5280 ( .A(n3626), .B(n3627), .Z(n3623) );
  AND U5281 ( .A(n3628), .B(n3629), .Z(n3626) );
  XNOR U5282 ( .A(x[1653]), .B(n3627), .Z(n3629) );
  XOR U5283 ( .A(n3630), .B(n3631), .Z(n3627) );
  AND U5284 ( .A(n3632), .B(n3633), .Z(n3630) );
  XNOR U5285 ( .A(x[1652]), .B(n3631), .Z(n3633) );
  XOR U5286 ( .A(n3634), .B(n3635), .Z(n3631) );
  AND U5287 ( .A(n3636), .B(n3637), .Z(n3634) );
  XNOR U5288 ( .A(x[1651]), .B(n3635), .Z(n3637) );
  XOR U5289 ( .A(n3638), .B(n3639), .Z(n3635) );
  AND U5290 ( .A(n3640), .B(n3641), .Z(n3638) );
  XNOR U5291 ( .A(x[1650]), .B(n3639), .Z(n3641) );
  XOR U5292 ( .A(n3642), .B(n3643), .Z(n3639) );
  AND U5293 ( .A(n3644), .B(n3645), .Z(n3642) );
  XNOR U5294 ( .A(x[1649]), .B(n3643), .Z(n3645) );
  XOR U5295 ( .A(n3646), .B(n3647), .Z(n3643) );
  AND U5296 ( .A(n3648), .B(n3649), .Z(n3646) );
  XNOR U5297 ( .A(x[1648]), .B(n3647), .Z(n3649) );
  XOR U5298 ( .A(n3650), .B(n3651), .Z(n3647) );
  AND U5299 ( .A(n3652), .B(n3653), .Z(n3650) );
  XNOR U5300 ( .A(x[1647]), .B(n3651), .Z(n3653) );
  XOR U5301 ( .A(n3654), .B(n3655), .Z(n3651) );
  AND U5302 ( .A(n3656), .B(n3657), .Z(n3654) );
  XNOR U5303 ( .A(x[1646]), .B(n3655), .Z(n3657) );
  XOR U5304 ( .A(n3658), .B(n3659), .Z(n3655) );
  AND U5305 ( .A(n3660), .B(n3661), .Z(n3658) );
  XNOR U5306 ( .A(x[1645]), .B(n3659), .Z(n3661) );
  XOR U5307 ( .A(n3662), .B(n3663), .Z(n3659) );
  AND U5308 ( .A(n3664), .B(n3665), .Z(n3662) );
  XNOR U5309 ( .A(x[1644]), .B(n3663), .Z(n3665) );
  XOR U5310 ( .A(n3666), .B(n3667), .Z(n3663) );
  AND U5311 ( .A(n3668), .B(n3669), .Z(n3666) );
  XNOR U5312 ( .A(x[1643]), .B(n3667), .Z(n3669) );
  XOR U5313 ( .A(n3670), .B(n3671), .Z(n3667) );
  AND U5314 ( .A(n3672), .B(n3673), .Z(n3670) );
  XNOR U5315 ( .A(x[1642]), .B(n3671), .Z(n3673) );
  XOR U5316 ( .A(n3674), .B(n3675), .Z(n3671) );
  AND U5317 ( .A(n3676), .B(n3677), .Z(n3674) );
  XNOR U5318 ( .A(x[1641]), .B(n3675), .Z(n3677) );
  XOR U5319 ( .A(n3678), .B(n3679), .Z(n3675) );
  AND U5320 ( .A(n3680), .B(n3681), .Z(n3678) );
  XNOR U5321 ( .A(x[1640]), .B(n3679), .Z(n3681) );
  XOR U5322 ( .A(n3682), .B(n3683), .Z(n3679) );
  AND U5323 ( .A(n3684), .B(n3685), .Z(n3682) );
  XNOR U5324 ( .A(x[1639]), .B(n3683), .Z(n3685) );
  XOR U5325 ( .A(n3686), .B(n3687), .Z(n3683) );
  AND U5326 ( .A(n3688), .B(n3689), .Z(n3686) );
  XNOR U5327 ( .A(x[1638]), .B(n3687), .Z(n3689) );
  XOR U5328 ( .A(n3690), .B(n3691), .Z(n3687) );
  AND U5329 ( .A(n3692), .B(n3693), .Z(n3690) );
  XNOR U5330 ( .A(x[1637]), .B(n3691), .Z(n3693) );
  XOR U5331 ( .A(n3694), .B(n3695), .Z(n3691) );
  AND U5332 ( .A(n3696), .B(n3697), .Z(n3694) );
  XNOR U5333 ( .A(x[1636]), .B(n3695), .Z(n3697) );
  XOR U5334 ( .A(n3698), .B(n3699), .Z(n3695) );
  AND U5335 ( .A(n3700), .B(n3701), .Z(n3698) );
  XNOR U5336 ( .A(x[1635]), .B(n3699), .Z(n3701) );
  XOR U5337 ( .A(n3702), .B(n3703), .Z(n3699) );
  AND U5338 ( .A(n3704), .B(n3705), .Z(n3702) );
  XNOR U5339 ( .A(x[1634]), .B(n3703), .Z(n3705) );
  XOR U5340 ( .A(n3706), .B(n3707), .Z(n3703) );
  AND U5341 ( .A(n3708), .B(n3709), .Z(n3706) );
  XNOR U5342 ( .A(x[1633]), .B(n3707), .Z(n3709) );
  XOR U5343 ( .A(n3710), .B(n3711), .Z(n3707) );
  AND U5344 ( .A(n3712), .B(n3713), .Z(n3710) );
  XNOR U5345 ( .A(x[1632]), .B(n3711), .Z(n3713) );
  XOR U5346 ( .A(n3714), .B(n3715), .Z(n3711) );
  AND U5347 ( .A(n3716), .B(n3717), .Z(n3714) );
  XNOR U5348 ( .A(x[1631]), .B(n3715), .Z(n3717) );
  XOR U5349 ( .A(n3718), .B(n3719), .Z(n3715) );
  AND U5350 ( .A(n3720), .B(n3721), .Z(n3718) );
  XNOR U5351 ( .A(x[1630]), .B(n3719), .Z(n3721) );
  XOR U5352 ( .A(n3722), .B(n3723), .Z(n3719) );
  AND U5353 ( .A(n3724), .B(n3725), .Z(n3722) );
  XNOR U5354 ( .A(x[1629]), .B(n3723), .Z(n3725) );
  XOR U5355 ( .A(n3726), .B(n3727), .Z(n3723) );
  AND U5356 ( .A(n3728), .B(n3729), .Z(n3726) );
  XNOR U5357 ( .A(x[1628]), .B(n3727), .Z(n3729) );
  XOR U5358 ( .A(n3730), .B(n3731), .Z(n3727) );
  AND U5359 ( .A(n3732), .B(n3733), .Z(n3730) );
  XNOR U5360 ( .A(x[1627]), .B(n3731), .Z(n3733) );
  XOR U5361 ( .A(n3734), .B(n3735), .Z(n3731) );
  AND U5362 ( .A(n3736), .B(n3737), .Z(n3734) );
  XNOR U5363 ( .A(x[1626]), .B(n3735), .Z(n3737) );
  XOR U5364 ( .A(n3738), .B(n3739), .Z(n3735) );
  AND U5365 ( .A(n3740), .B(n3741), .Z(n3738) );
  XNOR U5366 ( .A(x[1625]), .B(n3739), .Z(n3741) );
  XOR U5367 ( .A(n3742), .B(n3743), .Z(n3739) );
  AND U5368 ( .A(n3744), .B(n3745), .Z(n3742) );
  XNOR U5369 ( .A(x[1624]), .B(n3743), .Z(n3745) );
  XOR U5370 ( .A(n3746), .B(n3747), .Z(n3743) );
  AND U5371 ( .A(n3748), .B(n3749), .Z(n3746) );
  XNOR U5372 ( .A(x[1623]), .B(n3747), .Z(n3749) );
  XOR U5373 ( .A(n3750), .B(n3751), .Z(n3747) );
  AND U5374 ( .A(n3752), .B(n3753), .Z(n3750) );
  XNOR U5375 ( .A(x[1622]), .B(n3751), .Z(n3753) );
  XOR U5376 ( .A(n3754), .B(n3755), .Z(n3751) );
  AND U5377 ( .A(n3756), .B(n3757), .Z(n3754) );
  XNOR U5378 ( .A(x[1621]), .B(n3755), .Z(n3757) );
  XOR U5379 ( .A(n3758), .B(n3759), .Z(n3755) );
  AND U5380 ( .A(n3760), .B(n3761), .Z(n3758) );
  XNOR U5381 ( .A(x[1620]), .B(n3759), .Z(n3761) );
  XOR U5382 ( .A(n3762), .B(n3763), .Z(n3759) );
  AND U5383 ( .A(n3764), .B(n3765), .Z(n3762) );
  XNOR U5384 ( .A(x[1619]), .B(n3763), .Z(n3765) );
  XOR U5385 ( .A(n3766), .B(n3767), .Z(n3763) );
  AND U5386 ( .A(n3768), .B(n3769), .Z(n3766) );
  XNOR U5387 ( .A(x[1618]), .B(n3767), .Z(n3769) );
  XOR U5388 ( .A(n3770), .B(n3771), .Z(n3767) );
  AND U5389 ( .A(n3772), .B(n3773), .Z(n3770) );
  XNOR U5390 ( .A(x[1617]), .B(n3771), .Z(n3773) );
  XOR U5391 ( .A(n3774), .B(n3775), .Z(n3771) );
  AND U5392 ( .A(n3776), .B(n3777), .Z(n3774) );
  XNOR U5393 ( .A(x[1616]), .B(n3775), .Z(n3777) );
  XOR U5394 ( .A(n3778), .B(n3779), .Z(n3775) );
  AND U5395 ( .A(n3780), .B(n3781), .Z(n3778) );
  XNOR U5396 ( .A(x[1615]), .B(n3779), .Z(n3781) );
  XOR U5397 ( .A(n3782), .B(n3783), .Z(n3779) );
  AND U5398 ( .A(n3784), .B(n3785), .Z(n3782) );
  XNOR U5399 ( .A(x[1614]), .B(n3783), .Z(n3785) );
  XOR U5400 ( .A(n3786), .B(n3787), .Z(n3783) );
  AND U5401 ( .A(n3788), .B(n3789), .Z(n3786) );
  XNOR U5402 ( .A(x[1613]), .B(n3787), .Z(n3789) );
  XOR U5403 ( .A(n3790), .B(n3791), .Z(n3787) );
  AND U5404 ( .A(n3792), .B(n3793), .Z(n3790) );
  XNOR U5405 ( .A(x[1612]), .B(n3791), .Z(n3793) );
  XOR U5406 ( .A(n3794), .B(n3795), .Z(n3791) );
  AND U5407 ( .A(n3796), .B(n3797), .Z(n3794) );
  XNOR U5408 ( .A(x[1611]), .B(n3795), .Z(n3797) );
  XOR U5409 ( .A(n3798), .B(n3799), .Z(n3795) );
  AND U5410 ( .A(n3800), .B(n3801), .Z(n3798) );
  XNOR U5411 ( .A(x[1610]), .B(n3799), .Z(n3801) );
  XOR U5412 ( .A(n3802), .B(n3803), .Z(n3799) );
  AND U5413 ( .A(n3804), .B(n3805), .Z(n3802) );
  XNOR U5414 ( .A(x[1609]), .B(n3803), .Z(n3805) );
  XOR U5415 ( .A(n3806), .B(n3807), .Z(n3803) );
  AND U5416 ( .A(n3808), .B(n3809), .Z(n3806) );
  XNOR U5417 ( .A(x[1608]), .B(n3807), .Z(n3809) );
  XOR U5418 ( .A(n3810), .B(n3811), .Z(n3807) );
  AND U5419 ( .A(n3812), .B(n3813), .Z(n3810) );
  XNOR U5420 ( .A(x[1607]), .B(n3811), .Z(n3813) );
  XOR U5421 ( .A(n3814), .B(n3815), .Z(n3811) );
  AND U5422 ( .A(n3816), .B(n3817), .Z(n3814) );
  XNOR U5423 ( .A(x[1606]), .B(n3815), .Z(n3817) );
  XOR U5424 ( .A(n3818), .B(n3819), .Z(n3815) );
  AND U5425 ( .A(n3820), .B(n3821), .Z(n3818) );
  XNOR U5426 ( .A(x[1605]), .B(n3819), .Z(n3821) );
  XOR U5427 ( .A(n3822), .B(n3823), .Z(n3819) );
  AND U5428 ( .A(n3824), .B(n3825), .Z(n3822) );
  XNOR U5429 ( .A(x[1604]), .B(n3823), .Z(n3825) );
  XOR U5430 ( .A(n3826), .B(n3827), .Z(n3823) );
  AND U5431 ( .A(n3828), .B(n3829), .Z(n3826) );
  XNOR U5432 ( .A(x[1603]), .B(n3827), .Z(n3829) );
  XOR U5433 ( .A(n3830), .B(n3831), .Z(n3827) );
  AND U5434 ( .A(n3832), .B(n3833), .Z(n3830) );
  XNOR U5435 ( .A(x[1602]), .B(n3831), .Z(n3833) );
  XOR U5436 ( .A(n3834), .B(n3835), .Z(n3831) );
  AND U5437 ( .A(n3836), .B(n3837), .Z(n3834) );
  XNOR U5438 ( .A(x[1601]), .B(n3835), .Z(n3837) );
  XOR U5439 ( .A(n3838), .B(n3839), .Z(n3835) );
  AND U5440 ( .A(n3840), .B(n3841), .Z(n3838) );
  XNOR U5441 ( .A(x[1600]), .B(n3839), .Z(n3841) );
  XOR U5442 ( .A(n3842), .B(n3843), .Z(n3839) );
  AND U5443 ( .A(n3844), .B(n3845), .Z(n3842) );
  XNOR U5444 ( .A(x[1599]), .B(n3843), .Z(n3845) );
  XOR U5445 ( .A(n3846), .B(n3847), .Z(n3843) );
  AND U5446 ( .A(n3848), .B(n3849), .Z(n3846) );
  XNOR U5447 ( .A(x[1598]), .B(n3847), .Z(n3849) );
  XOR U5448 ( .A(n3850), .B(n3851), .Z(n3847) );
  AND U5449 ( .A(n3852), .B(n3853), .Z(n3850) );
  XNOR U5450 ( .A(x[1597]), .B(n3851), .Z(n3853) );
  XOR U5451 ( .A(n3854), .B(n3855), .Z(n3851) );
  AND U5452 ( .A(n3856), .B(n3857), .Z(n3854) );
  XNOR U5453 ( .A(x[1596]), .B(n3855), .Z(n3857) );
  XOR U5454 ( .A(n3858), .B(n3859), .Z(n3855) );
  AND U5455 ( .A(n3860), .B(n3861), .Z(n3858) );
  XNOR U5456 ( .A(x[1595]), .B(n3859), .Z(n3861) );
  XOR U5457 ( .A(n3862), .B(n3863), .Z(n3859) );
  AND U5458 ( .A(n3864), .B(n3865), .Z(n3862) );
  XNOR U5459 ( .A(x[1594]), .B(n3863), .Z(n3865) );
  XOR U5460 ( .A(n3866), .B(n3867), .Z(n3863) );
  AND U5461 ( .A(n3868), .B(n3869), .Z(n3866) );
  XNOR U5462 ( .A(x[1593]), .B(n3867), .Z(n3869) );
  XOR U5463 ( .A(n3870), .B(n3871), .Z(n3867) );
  AND U5464 ( .A(n3872), .B(n3873), .Z(n3870) );
  XNOR U5465 ( .A(x[1592]), .B(n3871), .Z(n3873) );
  XOR U5466 ( .A(n3874), .B(n3875), .Z(n3871) );
  AND U5467 ( .A(n3876), .B(n3877), .Z(n3874) );
  XNOR U5468 ( .A(x[1591]), .B(n3875), .Z(n3877) );
  XOR U5469 ( .A(n3878), .B(n3879), .Z(n3875) );
  AND U5470 ( .A(n3880), .B(n3881), .Z(n3878) );
  XNOR U5471 ( .A(x[1590]), .B(n3879), .Z(n3881) );
  XOR U5472 ( .A(n3882), .B(n3883), .Z(n3879) );
  AND U5473 ( .A(n3884), .B(n3885), .Z(n3882) );
  XNOR U5474 ( .A(x[1589]), .B(n3883), .Z(n3885) );
  XOR U5475 ( .A(n3886), .B(n3887), .Z(n3883) );
  AND U5476 ( .A(n3888), .B(n3889), .Z(n3886) );
  XNOR U5477 ( .A(x[1588]), .B(n3887), .Z(n3889) );
  XOR U5478 ( .A(n3890), .B(n3891), .Z(n3887) );
  AND U5479 ( .A(n3892), .B(n3893), .Z(n3890) );
  XNOR U5480 ( .A(x[1587]), .B(n3891), .Z(n3893) );
  XOR U5481 ( .A(n3894), .B(n3895), .Z(n3891) );
  AND U5482 ( .A(n3896), .B(n3897), .Z(n3894) );
  XNOR U5483 ( .A(x[1586]), .B(n3895), .Z(n3897) );
  XOR U5484 ( .A(n3898), .B(n3899), .Z(n3895) );
  AND U5485 ( .A(n3900), .B(n3901), .Z(n3898) );
  XNOR U5486 ( .A(x[1585]), .B(n3899), .Z(n3901) );
  XOR U5487 ( .A(n3902), .B(n3903), .Z(n3899) );
  AND U5488 ( .A(n3904), .B(n3905), .Z(n3902) );
  XNOR U5489 ( .A(x[1584]), .B(n3903), .Z(n3905) );
  XOR U5490 ( .A(n3906), .B(n3907), .Z(n3903) );
  AND U5491 ( .A(n3908), .B(n3909), .Z(n3906) );
  XNOR U5492 ( .A(x[1583]), .B(n3907), .Z(n3909) );
  XOR U5493 ( .A(n3910), .B(n3911), .Z(n3907) );
  AND U5494 ( .A(n3912), .B(n3913), .Z(n3910) );
  XNOR U5495 ( .A(x[1582]), .B(n3911), .Z(n3913) );
  XOR U5496 ( .A(n3914), .B(n3915), .Z(n3911) );
  AND U5497 ( .A(n3916), .B(n3917), .Z(n3914) );
  XNOR U5498 ( .A(x[1581]), .B(n3915), .Z(n3917) );
  XOR U5499 ( .A(n3918), .B(n3919), .Z(n3915) );
  AND U5500 ( .A(n3920), .B(n3921), .Z(n3918) );
  XNOR U5501 ( .A(x[1580]), .B(n3919), .Z(n3921) );
  XOR U5502 ( .A(n3922), .B(n3923), .Z(n3919) );
  AND U5503 ( .A(n3924), .B(n3925), .Z(n3922) );
  XNOR U5504 ( .A(x[1579]), .B(n3923), .Z(n3925) );
  XOR U5505 ( .A(n3926), .B(n3927), .Z(n3923) );
  AND U5506 ( .A(n3928), .B(n3929), .Z(n3926) );
  XNOR U5507 ( .A(x[1578]), .B(n3927), .Z(n3929) );
  XOR U5508 ( .A(n3930), .B(n3931), .Z(n3927) );
  AND U5509 ( .A(n3932), .B(n3933), .Z(n3930) );
  XNOR U5510 ( .A(x[1577]), .B(n3931), .Z(n3933) );
  XOR U5511 ( .A(n3934), .B(n3935), .Z(n3931) );
  AND U5512 ( .A(n3936), .B(n3937), .Z(n3934) );
  XNOR U5513 ( .A(x[1576]), .B(n3935), .Z(n3937) );
  XOR U5514 ( .A(n3938), .B(n3939), .Z(n3935) );
  AND U5515 ( .A(n3940), .B(n3941), .Z(n3938) );
  XNOR U5516 ( .A(x[1575]), .B(n3939), .Z(n3941) );
  XOR U5517 ( .A(n3942), .B(n3943), .Z(n3939) );
  AND U5518 ( .A(n3944), .B(n3945), .Z(n3942) );
  XNOR U5519 ( .A(x[1574]), .B(n3943), .Z(n3945) );
  XOR U5520 ( .A(n3946), .B(n3947), .Z(n3943) );
  AND U5521 ( .A(n3948), .B(n3949), .Z(n3946) );
  XNOR U5522 ( .A(x[1573]), .B(n3947), .Z(n3949) );
  XOR U5523 ( .A(n3950), .B(n3951), .Z(n3947) );
  AND U5524 ( .A(n3952), .B(n3953), .Z(n3950) );
  XNOR U5525 ( .A(x[1572]), .B(n3951), .Z(n3953) );
  XOR U5526 ( .A(n3954), .B(n3955), .Z(n3951) );
  AND U5527 ( .A(n3956), .B(n3957), .Z(n3954) );
  XNOR U5528 ( .A(x[1571]), .B(n3955), .Z(n3957) );
  XOR U5529 ( .A(n3958), .B(n3959), .Z(n3955) );
  AND U5530 ( .A(n3960), .B(n3961), .Z(n3958) );
  XNOR U5531 ( .A(x[1570]), .B(n3959), .Z(n3961) );
  XOR U5532 ( .A(n3962), .B(n3963), .Z(n3959) );
  AND U5533 ( .A(n3964), .B(n3965), .Z(n3962) );
  XNOR U5534 ( .A(x[1569]), .B(n3963), .Z(n3965) );
  XOR U5535 ( .A(n3966), .B(n3967), .Z(n3963) );
  AND U5536 ( .A(n3968), .B(n3969), .Z(n3966) );
  XNOR U5537 ( .A(x[1568]), .B(n3967), .Z(n3969) );
  XOR U5538 ( .A(n3970), .B(n3971), .Z(n3967) );
  AND U5539 ( .A(n3972), .B(n3973), .Z(n3970) );
  XNOR U5540 ( .A(x[1567]), .B(n3971), .Z(n3973) );
  XOR U5541 ( .A(n3974), .B(n3975), .Z(n3971) );
  AND U5542 ( .A(n3976), .B(n3977), .Z(n3974) );
  XNOR U5543 ( .A(x[1566]), .B(n3975), .Z(n3977) );
  XOR U5544 ( .A(n3978), .B(n3979), .Z(n3975) );
  AND U5545 ( .A(n3980), .B(n3981), .Z(n3978) );
  XNOR U5546 ( .A(x[1565]), .B(n3979), .Z(n3981) );
  XOR U5547 ( .A(n3982), .B(n3983), .Z(n3979) );
  AND U5548 ( .A(n3984), .B(n3985), .Z(n3982) );
  XNOR U5549 ( .A(x[1564]), .B(n3983), .Z(n3985) );
  XOR U5550 ( .A(n3986), .B(n3987), .Z(n3983) );
  AND U5551 ( .A(n3988), .B(n3989), .Z(n3986) );
  XNOR U5552 ( .A(x[1563]), .B(n3987), .Z(n3989) );
  XOR U5553 ( .A(n3990), .B(n3991), .Z(n3987) );
  AND U5554 ( .A(n3992), .B(n3993), .Z(n3990) );
  XNOR U5555 ( .A(x[1562]), .B(n3991), .Z(n3993) );
  XOR U5556 ( .A(n3994), .B(n3995), .Z(n3991) );
  AND U5557 ( .A(n3996), .B(n3997), .Z(n3994) );
  XNOR U5558 ( .A(x[1561]), .B(n3995), .Z(n3997) );
  XOR U5559 ( .A(n3998), .B(n3999), .Z(n3995) );
  AND U5560 ( .A(n4000), .B(n4001), .Z(n3998) );
  XNOR U5561 ( .A(x[1560]), .B(n3999), .Z(n4001) );
  XOR U5562 ( .A(n4002), .B(n4003), .Z(n3999) );
  AND U5563 ( .A(n4004), .B(n4005), .Z(n4002) );
  XNOR U5564 ( .A(x[1559]), .B(n4003), .Z(n4005) );
  XOR U5565 ( .A(n4006), .B(n4007), .Z(n4003) );
  AND U5566 ( .A(n4008), .B(n4009), .Z(n4006) );
  XNOR U5567 ( .A(x[1558]), .B(n4007), .Z(n4009) );
  XOR U5568 ( .A(n4010), .B(n4011), .Z(n4007) );
  AND U5569 ( .A(n4012), .B(n4013), .Z(n4010) );
  XNOR U5570 ( .A(x[1557]), .B(n4011), .Z(n4013) );
  XOR U5571 ( .A(n4014), .B(n4015), .Z(n4011) );
  AND U5572 ( .A(n4016), .B(n4017), .Z(n4014) );
  XNOR U5573 ( .A(x[1556]), .B(n4015), .Z(n4017) );
  XOR U5574 ( .A(n4018), .B(n4019), .Z(n4015) );
  AND U5575 ( .A(n4020), .B(n4021), .Z(n4018) );
  XNOR U5576 ( .A(x[1555]), .B(n4019), .Z(n4021) );
  XOR U5577 ( .A(n4022), .B(n4023), .Z(n4019) );
  AND U5578 ( .A(n4024), .B(n4025), .Z(n4022) );
  XNOR U5579 ( .A(x[1554]), .B(n4023), .Z(n4025) );
  XOR U5580 ( .A(n4026), .B(n4027), .Z(n4023) );
  AND U5581 ( .A(n4028), .B(n4029), .Z(n4026) );
  XNOR U5582 ( .A(x[1553]), .B(n4027), .Z(n4029) );
  XOR U5583 ( .A(n4030), .B(n4031), .Z(n4027) );
  AND U5584 ( .A(n4032), .B(n4033), .Z(n4030) );
  XNOR U5585 ( .A(x[1552]), .B(n4031), .Z(n4033) );
  XOR U5586 ( .A(n4034), .B(n4035), .Z(n4031) );
  AND U5587 ( .A(n4036), .B(n4037), .Z(n4034) );
  XNOR U5588 ( .A(x[1551]), .B(n4035), .Z(n4037) );
  XOR U5589 ( .A(n4038), .B(n4039), .Z(n4035) );
  AND U5590 ( .A(n4040), .B(n4041), .Z(n4038) );
  XNOR U5591 ( .A(x[1550]), .B(n4039), .Z(n4041) );
  XOR U5592 ( .A(n4042), .B(n4043), .Z(n4039) );
  AND U5593 ( .A(n4044), .B(n4045), .Z(n4042) );
  XNOR U5594 ( .A(x[1549]), .B(n4043), .Z(n4045) );
  XOR U5595 ( .A(n4046), .B(n4047), .Z(n4043) );
  AND U5596 ( .A(n4048), .B(n4049), .Z(n4046) );
  XNOR U5597 ( .A(x[1548]), .B(n4047), .Z(n4049) );
  XOR U5598 ( .A(n4050), .B(n4051), .Z(n4047) );
  AND U5599 ( .A(n4052), .B(n4053), .Z(n4050) );
  XNOR U5600 ( .A(x[1547]), .B(n4051), .Z(n4053) );
  XOR U5601 ( .A(n4054), .B(n4055), .Z(n4051) );
  AND U5602 ( .A(n4056), .B(n4057), .Z(n4054) );
  XNOR U5603 ( .A(x[1546]), .B(n4055), .Z(n4057) );
  XOR U5604 ( .A(n4058), .B(n4059), .Z(n4055) );
  AND U5605 ( .A(n4060), .B(n4061), .Z(n4058) );
  XNOR U5606 ( .A(x[1545]), .B(n4059), .Z(n4061) );
  XOR U5607 ( .A(n4062), .B(n4063), .Z(n4059) );
  AND U5608 ( .A(n4064), .B(n4065), .Z(n4062) );
  XNOR U5609 ( .A(x[1544]), .B(n4063), .Z(n4065) );
  XOR U5610 ( .A(n4066), .B(n4067), .Z(n4063) );
  AND U5611 ( .A(n4068), .B(n4069), .Z(n4066) );
  XNOR U5612 ( .A(x[1543]), .B(n4067), .Z(n4069) );
  XOR U5613 ( .A(n4070), .B(n4071), .Z(n4067) );
  AND U5614 ( .A(n4072), .B(n4073), .Z(n4070) );
  XNOR U5615 ( .A(x[1542]), .B(n4071), .Z(n4073) );
  XOR U5616 ( .A(n4074), .B(n4075), .Z(n4071) );
  AND U5617 ( .A(n4076), .B(n4077), .Z(n4074) );
  XNOR U5618 ( .A(x[1541]), .B(n4075), .Z(n4077) );
  XOR U5619 ( .A(n4078), .B(n4079), .Z(n4075) );
  AND U5620 ( .A(n4080), .B(n4081), .Z(n4078) );
  XNOR U5621 ( .A(x[1540]), .B(n4079), .Z(n4081) );
  XOR U5622 ( .A(n4082), .B(n4083), .Z(n4079) );
  AND U5623 ( .A(n4084), .B(n4085), .Z(n4082) );
  XNOR U5624 ( .A(x[1539]), .B(n4083), .Z(n4085) );
  XOR U5625 ( .A(n4086), .B(n4087), .Z(n4083) );
  AND U5626 ( .A(n4088), .B(n4089), .Z(n4086) );
  XNOR U5627 ( .A(x[1538]), .B(n4087), .Z(n4089) );
  XOR U5628 ( .A(n4090), .B(n4091), .Z(n4087) );
  AND U5629 ( .A(n4092), .B(n4093), .Z(n4090) );
  XNOR U5630 ( .A(x[1537]), .B(n4091), .Z(n4093) );
  XOR U5631 ( .A(n4094), .B(n4095), .Z(n4091) );
  AND U5632 ( .A(n4096), .B(n4097), .Z(n4094) );
  XNOR U5633 ( .A(x[1536]), .B(n4095), .Z(n4097) );
  XOR U5634 ( .A(n4098), .B(n4099), .Z(n4095) );
  AND U5635 ( .A(n4100), .B(n4101), .Z(n4098) );
  XNOR U5636 ( .A(x[1535]), .B(n4099), .Z(n4101) );
  XOR U5637 ( .A(n4102), .B(n4103), .Z(n4099) );
  AND U5638 ( .A(n4104), .B(n4105), .Z(n4102) );
  XNOR U5639 ( .A(x[1534]), .B(n4103), .Z(n4105) );
  XOR U5640 ( .A(n4106), .B(n4107), .Z(n4103) );
  AND U5641 ( .A(n4108), .B(n4109), .Z(n4106) );
  XNOR U5642 ( .A(x[1533]), .B(n4107), .Z(n4109) );
  XOR U5643 ( .A(n4110), .B(n4111), .Z(n4107) );
  AND U5644 ( .A(n4112), .B(n4113), .Z(n4110) );
  XNOR U5645 ( .A(x[1532]), .B(n4111), .Z(n4113) );
  XOR U5646 ( .A(n4114), .B(n4115), .Z(n4111) );
  AND U5647 ( .A(n4116), .B(n4117), .Z(n4114) );
  XNOR U5648 ( .A(x[1531]), .B(n4115), .Z(n4117) );
  XOR U5649 ( .A(n4118), .B(n4119), .Z(n4115) );
  AND U5650 ( .A(n4120), .B(n4121), .Z(n4118) );
  XNOR U5651 ( .A(x[1530]), .B(n4119), .Z(n4121) );
  XOR U5652 ( .A(n4122), .B(n4123), .Z(n4119) );
  AND U5653 ( .A(n4124), .B(n4125), .Z(n4122) );
  XNOR U5654 ( .A(x[1529]), .B(n4123), .Z(n4125) );
  XOR U5655 ( .A(n4126), .B(n4127), .Z(n4123) );
  AND U5656 ( .A(n4128), .B(n4129), .Z(n4126) );
  XNOR U5657 ( .A(x[1528]), .B(n4127), .Z(n4129) );
  XOR U5658 ( .A(n4130), .B(n4131), .Z(n4127) );
  AND U5659 ( .A(n4132), .B(n4133), .Z(n4130) );
  XNOR U5660 ( .A(x[1527]), .B(n4131), .Z(n4133) );
  XOR U5661 ( .A(n4134), .B(n4135), .Z(n4131) );
  AND U5662 ( .A(n4136), .B(n4137), .Z(n4134) );
  XNOR U5663 ( .A(x[1526]), .B(n4135), .Z(n4137) );
  XOR U5664 ( .A(n4138), .B(n4139), .Z(n4135) );
  AND U5665 ( .A(n4140), .B(n4141), .Z(n4138) );
  XNOR U5666 ( .A(x[1525]), .B(n4139), .Z(n4141) );
  XOR U5667 ( .A(n4142), .B(n4143), .Z(n4139) );
  AND U5668 ( .A(n4144), .B(n4145), .Z(n4142) );
  XNOR U5669 ( .A(x[1524]), .B(n4143), .Z(n4145) );
  XOR U5670 ( .A(n4146), .B(n4147), .Z(n4143) );
  AND U5671 ( .A(n4148), .B(n4149), .Z(n4146) );
  XNOR U5672 ( .A(x[1523]), .B(n4147), .Z(n4149) );
  XOR U5673 ( .A(n4150), .B(n4151), .Z(n4147) );
  AND U5674 ( .A(n4152), .B(n4153), .Z(n4150) );
  XNOR U5675 ( .A(x[1522]), .B(n4151), .Z(n4153) );
  XOR U5676 ( .A(n4154), .B(n4155), .Z(n4151) );
  AND U5677 ( .A(n4156), .B(n4157), .Z(n4154) );
  XNOR U5678 ( .A(x[1521]), .B(n4155), .Z(n4157) );
  XOR U5679 ( .A(n4158), .B(n4159), .Z(n4155) );
  AND U5680 ( .A(n4160), .B(n4161), .Z(n4158) );
  XNOR U5681 ( .A(x[1520]), .B(n4159), .Z(n4161) );
  XOR U5682 ( .A(n4162), .B(n4163), .Z(n4159) );
  AND U5683 ( .A(n4164), .B(n4165), .Z(n4162) );
  XNOR U5684 ( .A(x[1519]), .B(n4163), .Z(n4165) );
  XOR U5685 ( .A(n4166), .B(n4167), .Z(n4163) );
  AND U5686 ( .A(n4168), .B(n4169), .Z(n4166) );
  XNOR U5687 ( .A(x[1518]), .B(n4167), .Z(n4169) );
  XOR U5688 ( .A(n4170), .B(n4171), .Z(n4167) );
  AND U5689 ( .A(n4172), .B(n4173), .Z(n4170) );
  XNOR U5690 ( .A(x[1517]), .B(n4171), .Z(n4173) );
  XOR U5691 ( .A(n4174), .B(n4175), .Z(n4171) );
  AND U5692 ( .A(n4176), .B(n4177), .Z(n4174) );
  XNOR U5693 ( .A(x[1516]), .B(n4175), .Z(n4177) );
  XOR U5694 ( .A(n4178), .B(n4179), .Z(n4175) );
  AND U5695 ( .A(n4180), .B(n4181), .Z(n4178) );
  XNOR U5696 ( .A(x[1515]), .B(n4179), .Z(n4181) );
  XOR U5697 ( .A(n4182), .B(n4183), .Z(n4179) );
  AND U5698 ( .A(n4184), .B(n4185), .Z(n4182) );
  XNOR U5699 ( .A(x[1514]), .B(n4183), .Z(n4185) );
  XOR U5700 ( .A(n4186), .B(n4187), .Z(n4183) );
  AND U5701 ( .A(n4188), .B(n4189), .Z(n4186) );
  XNOR U5702 ( .A(x[1513]), .B(n4187), .Z(n4189) );
  XOR U5703 ( .A(n4190), .B(n4191), .Z(n4187) );
  AND U5704 ( .A(n4192), .B(n4193), .Z(n4190) );
  XNOR U5705 ( .A(x[1512]), .B(n4191), .Z(n4193) );
  XOR U5706 ( .A(n4194), .B(n4195), .Z(n4191) );
  AND U5707 ( .A(n4196), .B(n4197), .Z(n4194) );
  XNOR U5708 ( .A(x[1511]), .B(n4195), .Z(n4197) );
  XOR U5709 ( .A(n4198), .B(n4199), .Z(n4195) );
  AND U5710 ( .A(n4200), .B(n4201), .Z(n4198) );
  XNOR U5711 ( .A(x[1510]), .B(n4199), .Z(n4201) );
  XOR U5712 ( .A(n4202), .B(n4203), .Z(n4199) );
  AND U5713 ( .A(n4204), .B(n4205), .Z(n4202) );
  XNOR U5714 ( .A(x[1509]), .B(n4203), .Z(n4205) );
  XOR U5715 ( .A(n4206), .B(n4207), .Z(n4203) );
  AND U5716 ( .A(n4208), .B(n4209), .Z(n4206) );
  XNOR U5717 ( .A(x[1508]), .B(n4207), .Z(n4209) );
  XOR U5718 ( .A(n4210), .B(n4211), .Z(n4207) );
  AND U5719 ( .A(n4212), .B(n4213), .Z(n4210) );
  XNOR U5720 ( .A(x[1507]), .B(n4211), .Z(n4213) );
  XOR U5721 ( .A(n4214), .B(n4215), .Z(n4211) );
  AND U5722 ( .A(n4216), .B(n4217), .Z(n4214) );
  XNOR U5723 ( .A(x[1506]), .B(n4215), .Z(n4217) );
  XOR U5724 ( .A(n4218), .B(n4219), .Z(n4215) );
  AND U5725 ( .A(n4220), .B(n4221), .Z(n4218) );
  XNOR U5726 ( .A(x[1505]), .B(n4219), .Z(n4221) );
  XOR U5727 ( .A(n4222), .B(n4223), .Z(n4219) );
  AND U5728 ( .A(n4224), .B(n4225), .Z(n4222) );
  XNOR U5729 ( .A(x[1504]), .B(n4223), .Z(n4225) );
  XOR U5730 ( .A(n4226), .B(n4227), .Z(n4223) );
  AND U5731 ( .A(n4228), .B(n4229), .Z(n4226) );
  XNOR U5732 ( .A(x[1503]), .B(n4227), .Z(n4229) );
  XOR U5733 ( .A(n4230), .B(n4231), .Z(n4227) );
  AND U5734 ( .A(n4232), .B(n4233), .Z(n4230) );
  XNOR U5735 ( .A(x[1502]), .B(n4231), .Z(n4233) );
  XOR U5736 ( .A(n4234), .B(n4235), .Z(n4231) );
  AND U5737 ( .A(n4236), .B(n4237), .Z(n4234) );
  XNOR U5738 ( .A(x[1501]), .B(n4235), .Z(n4237) );
  XOR U5739 ( .A(n4238), .B(n4239), .Z(n4235) );
  AND U5740 ( .A(n4240), .B(n4241), .Z(n4238) );
  XNOR U5741 ( .A(x[1500]), .B(n4239), .Z(n4241) );
  XOR U5742 ( .A(n4242), .B(n4243), .Z(n4239) );
  AND U5743 ( .A(n4244), .B(n4245), .Z(n4242) );
  XNOR U5744 ( .A(x[1499]), .B(n4243), .Z(n4245) );
  XOR U5745 ( .A(n4246), .B(n4247), .Z(n4243) );
  AND U5746 ( .A(n4248), .B(n4249), .Z(n4246) );
  XNOR U5747 ( .A(x[1498]), .B(n4247), .Z(n4249) );
  XOR U5748 ( .A(n4250), .B(n4251), .Z(n4247) );
  AND U5749 ( .A(n4252), .B(n4253), .Z(n4250) );
  XNOR U5750 ( .A(x[1497]), .B(n4251), .Z(n4253) );
  XOR U5751 ( .A(n4254), .B(n4255), .Z(n4251) );
  AND U5752 ( .A(n4256), .B(n4257), .Z(n4254) );
  XNOR U5753 ( .A(x[1496]), .B(n4255), .Z(n4257) );
  XOR U5754 ( .A(n4258), .B(n4259), .Z(n4255) );
  AND U5755 ( .A(n4260), .B(n4261), .Z(n4258) );
  XNOR U5756 ( .A(x[1495]), .B(n4259), .Z(n4261) );
  XOR U5757 ( .A(n4262), .B(n4263), .Z(n4259) );
  AND U5758 ( .A(n4264), .B(n4265), .Z(n4262) );
  XNOR U5759 ( .A(x[1494]), .B(n4263), .Z(n4265) );
  XOR U5760 ( .A(n4266), .B(n4267), .Z(n4263) );
  AND U5761 ( .A(n4268), .B(n4269), .Z(n4266) );
  XNOR U5762 ( .A(x[1493]), .B(n4267), .Z(n4269) );
  XOR U5763 ( .A(n4270), .B(n4271), .Z(n4267) );
  AND U5764 ( .A(n4272), .B(n4273), .Z(n4270) );
  XNOR U5765 ( .A(x[1492]), .B(n4271), .Z(n4273) );
  XOR U5766 ( .A(n4274), .B(n4275), .Z(n4271) );
  AND U5767 ( .A(n4276), .B(n4277), .Z(n4274) );
  XNOR U5768 ( .A(x[1491]), .B(n4275), .Z(n4277) );
  XOR U5769 ( .A(n4278), .B(n4279), .Z(n4275) );
  AND U5770 ( .A(n4280), .B(n4281), .Z(n4278) );
  XNOR U5771 ( .A(x[1490]), .B(n4279), .Z(n4281) );
  XOR U5772 ( .A(n4282), .B(n4283), .Z(n4279) );
  AND U5773 ( .A(n4284), .B(n4285), .Z(n4282) );
  XNOR U5774 ( .A(x[1489]), .B(n4283), .Z(n4285) );
  XOR U5775 ( .A(n4286), .B(n4287), .Z(n4283) );
  AND U5776 ( .A(n4288), .B(n4289), .Z(n4286) );
  XNOR U5777 ( .A(x[1488]), .B(n4287), .Z(n4289) );
  XOR U5778 ( .A(n4290), .B(n4291), .Z(n4287) );
  AND U5779 ( .A(n4292), .B(n4293), .Z(n4290) );
  XNOR U5780 ( .A(x[1487]), .B(n4291), .Z(n4293) );
  XOR U5781 ( .A(n4294), .B(n4295), .Z(n4291) );
  AND U5782 ( .A(n4296), .B(n4297), .Z(n4294) );
  XNOR U5783 ( .A(x[1486]), .B(n4295), .Z(n4297) );
  XOR U5784 ( .A(n4298), .B(n4299), .Z(n4295) );
  AND U5785 ( .A(n4300), .B(n4301), .Z(n4298) );
  XNOR U5786 ( .A(x[1485]), .B(n4299), .Z(n4301) );
  XOR U5787 ( .A(n4302), .B(n4303), .Z(n4299) );
  AND U5788 ( .A(n4304), .B(n4305), .Z(n4302) );
  XNOR U5789 ( .A(x[1484]), .B(n4303), .Z(n4305) );
  XOR U5790 ( .A(n4306), .B(n4307), .Z(n4303) );
  AND U5791 ( .A(n4308), .B(n4309), .Z(n4306) );
  XNOR U5792 ( .A(x[1483]), .B(n4307), .Z(n4309) );
  XOR U5793 ( .A(n4310), .B(n4311), .Z(n4307) );
  AND U5794 ( .A(n4312), .B(n4313), .Z(n4310) );
  XNOR U5795 ( .A(x[1482]), .B(n4311), .Z(n4313) );
  XOR U5796 ( .A(n4314), .B(n4315), .Z(n4311) );
  AND U5797 ( .A(n4316), .B(n4317), .Z(n4314) );
  XNOR U5798 ( .A(x[1481]), .B(n4315), .Z(n4317) );
  XOR U5799 ( .A(n4318), .B(n4319), .Z(n4315) );
  AND U5800 ( .A(n4320), .B(n4321), .Z(n4318) );
  XNOR U5801 ( .A(x[1480]), .B(n4319), .Z(n4321) );
  XOR U5802 ( .A(n4322), .B(n4323), .Z(n4319) );
  AND U5803 ( .A(n4324), .B(n4325), .Z(n4322) );
  XNOR U5804 ( .A(x[1479]), .B(n4323), .Z(n4325) );
  XOR U5805 ( .A(n4326), .B(n4327), .Z(n4323) );
  AND U5806 ( .A(n4328), .B(n4329), .Z(n4326) );
  XNOR U5807 ( .A(x[1478]), .B(n4327), .Z(n4329) );
  XOR U5808 ( .A(n4330), .B(n4331), .Z(n4327) );
  AND U5809 ( .A(n4332), .B(n4333), .Z(n4330) );
  XNOR U5810 ( .A(x[1477]), .B(n4331), .Z(n4333) );
  XOR U5811 ( .A(n4334), .B(n4335), .Z(n4331) );
  AND U5812 ( .A(n4336), .B(n4337), .Z(n4334) );
  XNOR U5813 ( .A(x[1476]), .B(n4335), .Z(n4337) );
  XOR U5814 ( .A(n4338), .B(n4339), .Z(n4335) );
  AND U5815 ( .A(n4340), .B(n4341), .Z(n4338) );
  XNOR U5816 ( .A(x[1475]), .B(n4339), .Z(n4341) );
  XOR U5817 ( .A(n4342), .B(n4343), .Z(n4339) );
  AND U5818 ( .A(n4344), .B(n4345), .Z(n4342) );
  XNOR U5819 ( .A(x[1474]), .B(n4343), .Z(n4345) );
  XOR U5820 ( .A(n4346), .B(n4347), .Z(n4343) );
  AND U5821 ( .A(n4348), .B(n4349), .Z(n4346) );
  XNOR U5822 ( .A(x[1473]), .B(n4347), .Z(n4349) );
  XOR U5823 ( .A(n4350), .B(n4351), .Z(n4347) );
  AND U5824 ( .A(n4352), .B(n4353), .Z(n4350) );
  XNOR U5825 ( .A(x[1472]), .B(n4351), .Z(n4353) );
  XOR U5826 ( .A(n4354), .B(n4355), .Z(n4351) );
  AND U5827 ( .A(n4356), .B(n4357), .Z(n4354) );
  XNOR U5828 ( .A(x[1471]), .B(n4355), .Z(n4357) );
  XOR U5829 ( .A(n4358), .B(n4359), .Z(n4355) );
  AND U5830 ( .A(n4360), .B(n4361), .Z(n4358) );
  XNOR U5831 ( .A(x[1470]), .B(n4359), .Z(n4361) );
  XOR U5832 ( .A(n4362), .B(n4363), .Z(n4359) );
  AND U5833 ( .A(n4364), .B(n4365), .Z(n4362) );
  XNOR U5834 ( .A(x[1469]), .B(n4363), .Z(n4365) );
  XOR U5835 ( .A(n4366), .B(n4367), .Z(n4363) );
  AND U5836 ( .A(n4368), .B(n4369), .Z(n4366) );
  XNOR U5837 ( .A(x[1468]), .B(n4367), .Z(n4369) );
  XOR U5838 ( .A(n4370), .B(n4371), .Z(n4367) );
  AND U5839 ( .A(n4372), .B(n4373), .Z(n4370) );
  XNOR U5840 ( .A(x[1467]), .B(n4371), .Z(n4373) );
  XOR U5841 ( .A(n4374), .B(n4375), .Z(n4371) );
  AND U5842 ( .A(n4376), .B(n4377), .Z(n4374) );
  XNOR U5843 ( .A(x[1466]), .B(n4375), .Z(n4377) );
  XOR U5844 ( .A(n4378), .B(n4379), .Z(n4375) );
  AND U5845 ( .A(n4380), .B(n4381), .Z(n4378) );
  XNOR U5846 ( .A(x[1465]), .B(n4379), .Z(n4381) );
  XOR U5847 ( .A(n4382), .B(n4383), .Z(n4379) );
  AND U5848 ( .A(n4384), .B(n4385), .Z(n4382) );
  XNOR U5849 ( .A(x[1464]), .B(n4383), .Z(n4385) );
  XOR U5850 ( .A(n4386), .B(n4387), .Z(n4383) );
  AND U5851 ( .A(n4388), .B(n4389), .Z(n4386) );
  XNOR U5852 ( .A(x[1463]), .B(n4387), .Z(n4389) );
  XOR U5853 ( .A(n4390), .B(n4391), .Z(n4387) );
  AND U5854 ( .A(n4392), .B(n4393), .Z(n4390) );
  XNOR U5855 ( .A(x[1462]), .B(n4391), .Z(n4393) );
  XOR U5856 ( .A(n4394), .B(n4395), .Z(n4391) );
  AND U5857 ( .A(n4396), .B(n4397), .Z(n4394) );
  XNOR U5858 ( .A(x[1461]), .B(n4395), .Z(n4397) );
  XOR U5859 ( .A(n4398), .B(n4399), .Z(n4395) );
  AND U5860 ( .A(n4400), .B(n4401), .Z(n4398) );
  XNOR U5861 ( .A(x[1460]), .B(n4399), .Z(n4401) );
  XOR U5862 ( .A(n4402), .B(n4403), .Z(n4399) );
  AND U5863 ( .A(n4404), .B(n4405), .Z(n4402) );
  XNOR U5864 ( .A(x[1459]), .B(n4403), .Z(n4405) );
  XOR U5865 ( .A(n4406), .B(n4407), .Z(n4403) );
  AND U5866 ( .A(n4408), .B(n4409), .Z(n4406) );
  XNOR U5867 ( .A(x[1458]), .B(n4407), .Z(n4409) );
  XOR U5868 ( .A(n4410), .B(n4411), .Z(n4407) );
  AND U5869 ( .A(n4412), .B(n4413), .Z(n4410) );
  XNOR U5870 ( .A(x[1457]), .B(n4411), .Z(n4413) );
  XOR U5871 ( .A(n4414), .B(n4415), .Z(n4411) );
  AND U5872 ( .A(n4416), .B(n4417), .Z(n4414) );
  XNOR U5873 ( .A(x[1456]), .B(n4415), .Z(n4417) );
  XOR U5874 ( .A(n4418), .B(n4419), .Z(n4415) );
  AND U5875 ( .A(n4420), .B(n4421), .Z(n4418) );
  XNOR U5876 ( .A(x[1455]), .B(n4419), .Z(n4421) );
  XOR U5877 ( .A(n4422), .B(n4423), .Z(n4419) );
  AND U5878 ( .A(n4424), .B(n4425), .Z(n4422) );
  XNOR U5879 ( .A(x[1454]), .B(n4423), .Z(n4425) );
  XOR U5880 ( .A(n4426), .B(n4427), .Z(n4423) );
  AND U5881 ( .A(n4428), .B(n4429), .Z(n4426) );
  XNOR U5882 ( .A(x[1453]), .B(n4427), .Z(n4429) );
  XOR U5883 ( .A(n4430), .B(n4431), .Z(n4427) );
  AND U5884 ( .A(n4432), .B(n4433), .Z(n4430) );
  XNOR U5885 ( .A(x[1452]), .B(n4431), .Z(n4433) );
  XOR U5886 ( .A(n4434), .B(n4435), .Z(n4431) );
  AND U5887 ( .A(n4436), .B(n4437), .Z(n4434) );
  XNOR U5888 ( .A(x[1451]), .B(n4435), .Z(n4437) );
  XOR U5889 ( .A(n4438), .B(n4439), .Z(n4435) );
  AND U5890 ( .A(n4440), .B(n4441), .Z(n4438) );
  XNOR U5891 ( .A(x[1450]), .B(n4439), .Z(n4441) );
  XOR U5892 ( .A(n4442), .B(n4443), .Z(n4439) );
  AND U5893 ( .A(n4444), .B(n4445), .Z(n4442) );
  XNOR U5894 ( .A(x[1449]), .B(n4443), .Z(n4445) );
  XOR U5895 ( .A(n4446), .B(n4447), .Z(n4443) );
  AND U5896 ( .A(n4448), .B(n4449), .Z(n4446) );
  XNOR U5897 ( .A(x[1448]), .B(n4447), .Z(n4449) );
  XOR U5898 ( .A(n4450), .B(n4451), .Z(n4447) );
  AND U5899 ( .A(n4452), .B(n4453), .Z(n4450) );
  XNOR U5900 ( .A(x[1447]), .B(n4451), .Z(n4453) );
  XOR U5901 ( .A(n4454), .B(n4455), .Z(n4451) );
  AND U5902 ( .A(n4456), .B(n4457), .Z(n4454) );
  XNOR U5903 ( .A(x[1446]), .B(n4455), .Z(n4457) );
  XOR U5904 ( .A(n4458), .B(n4459), .Z(n4455) );
  AND U5905 ( .A(n4460), .B(n4461), .Z(n4458) );
  XNOR U5906 ( .A(x[1445]), .B(n4459), .Z(n4461) );
  XOR U5907 ( .A(n4462), .B(n4463), .Z(n4459) );
  AND U5908 ( .A(n4464), .B(n4465), .Z(n4462) );
  XNOR U5909 ( .A(x[1444]), .B(n4463), .Z(n4465) );
  XOR U5910 ( .A(n4466), .B(n4467), .Z(n4463) );
  AND U5911 ( .A(n4468), .B(n4469), .Z(n4466) );
  XNOR U5912 ( .A(x[1443]), .B(n4467), .Z(n4469) );
  XOR U5913 ( .A(n4470), .B(n4471), .Z(n4467) );
  AND U5914 ( .A(n4472), .B(n4473), .Z(n4470) );
  XNOR U5915 ( .A(x[1442]), .B(n4471), .Z(n4473) );
  XOR U5916 ( .A(n4474), .B(n4475), .Z(n4471) );
  AND U5917 ( .A(n4476), .B(n4477), .Z(n4474) );
  XNOR U5918 ( .A(x[1441]), .B(n4475), .Z(n4477) );
  XOR U5919 ( .A(n4478), .B(n4479), .Z(n4475) );
  AND U5920 ( .A(n4480), .B(n4481), .Z(n4478) );
  XNOR U5921 ( .A(x[1440]), .B(n4479), .Z(n4481) );
  XOR U5922 ( .A(n4482), .B(n4483), .Z(n4479) );
  AND U5923 ( .A(n4484), .B(n4485), .Z(n4482) );
  XNOR U5924 ( .A(x[1439]), .B(n4483), .Z(n4485) );
  XOR U5925 ( .A(n4486), .B(n4487), .Z(n4483) );
  AND U5926 ( .A(n4488), .B(n4489), .Z(n4486) );
  XNOR U5927 ( .A(x[1438]), .B(n4487), .Z(n4489) );
  XOR U5928 ( .A(n4490), .B(n4491), .Z(n4487) );
  AND U5929 ( .A(n4492), .B(n4493), .Z(n4490) );
  XNOR U5930 ( .A(x[1437]), .B(n4491), .Z(n4493) );
  XOR U5931 ( .A(n4494), .B(n4495), .Z(n4491) );
  AND U5932 ( .A(n4496), .B(n4497), .Z(n4494) );
  XNOR U5933 ( .A(x[1436]), .B(n4495), .Z(n4497) );
  XOR U5934 ( .A(n4498), .B(n4499), .Z(n4495) );
  AND U5935 ( .A(n4500), .B(n4501), .Z(n4498) );
  XNOR U5936 ( .A(x[1435]), .B(n4499), .Z(n4501) );
  XOR U5937 ( .A(n4502), .B(n4503), .Z(n4499) );
  AND U5938 ( .A(n4504), .B(n4505), .Z(n4502) );
  XNOR U5939 ( .A(x[1434]), .B(n4503), .Z(n4505) );
  XOR U5940 ( .A(n4506), .B(n4507), .Z(n4503) );
  AND U5941 ( .A(n4508), .B(n4509), .Z(n4506) );
  XNOR U5942 ( .A(x[1433]), .B(n4507), .Z(n4509) );
  XOR U5943 ( .A(n4510), .B(n4511), .Z(n4507) );
  AND U5944 ( .A(n4512), .B(n4513), .Z(n4510) );
  XNOR U5945 ( .A(x[1432]), .B(n4511), .Z(n4513) );
  XOR U5946 ( .A(n4514), .B(n4515), .Z(n4511) );
  AND U5947 ( .A(n4516), .B(n4517), .Z(n4514) );
  XNOR U5948 ( .A(x[1431]), .B(n4515), .Z(n4517) );
  XOR U5949 ( .A(n4518), .B(n4519), .Z(n4515) );
  AND U5950 ( .A(n4520), .B(n4521), .Z(n4518) );
  XNOR U5951 ( .A(x[1430]), .B(n4519), .Z(n4521) );
  XOR U5952 ( .A(n4522), .B(n4523), .Z(n4519) );
  AND U5953 ( .A(n4524), .B(n4525), .Z(n4522) );
  XNOR U5954 ( .A(x[1429]), .B(n4523), .Z(n4525) );
  XOR U5955 ( .A(n4526), .B(n4527), .Z(n4523) );
  AND U5956 ( .A(n4528), .B(n4529), .Z(n4526) );
  XNOR U5957 ( .A(x[1428]), .B(n4527), .Z(n4529) );
  XOR U5958 ( .A(n4530), .B(n4531), .Z(n4527) );
  AND U5959 ( .A(n4532), .B(n4533), .Z(n4530) );
  XNOR U5960 ( .A(x[1427]), .B(n4531), .Z(n4533) );
  XOR U5961 ( .A(n4534), .B(n4535), .Z(n4531) );
  AND U5962 ( .A(n4536), .B(n4537), .Z(n4534) );
  XNOR U5963 ( .A(x[1426]), .B(n4535), .Z(n4537) );
  XOR U5964 ( .A(n4538), .B(n4539), .Z(n4535) );
  AND U5965 ( .A(n4540), .B(n4541), .Z(n4538) );
  XNOR U5966 ( .A(x[1425]), .B(n4539), .Z(n4541) );
  XOR U5967 ( .A(n4542), .B(n4543), .Z(n4539) );
  AND U5968 ( .A(n4544), .B(n4545), .Z(n4542) );
  XNOR U5969 ( .A(x[1424]), .B(n4543), .Z(n4545) );
  XOR U5970 ( .A(n4546), .B(n4547), .Z(n4543) );
  AND U5971 ( .A(n4548), .B(n4549), .Z(n4546) );
  XNOR U5972 ( .A(x[1423]), .B(n4547), .Z(n4549) );
  XOR U5973 ( .A(n4550), .B(n4551), .Z(n4547) );
  AND U5974 ( .A(n4552), .B(n4553), .Z(n4550) );
  XNOR U5975 ( .A(x[1422]), .B(n4551), .Z(n4553) );
  XOR U5976 ( .A(n4554), .B(n4555), .Z(n4551) );
  AND U5977 ( .A(n4556), .B(n4557), .Z(n4554) );
  XNOR U5978 ( .A(x[1421]), .B(n4555), .Z(n4557) );
  XOR U5979 ( .A(n4558), .B(n4559), .Z(n4555) );
  AND U5980 ( .A(n4560), .B(n4561), .Z(n4558) );
  XNOR U5981 ( .A(x[1420]), .B(n4559), .Z(n4561) );
  XOR U5982 ( .A(n4562), .B(n4563), .Z(n4559) );
  AND U5983 ( .A(n4564), .B(n4565), .Z(n4562) );
  XNOR U5984 ( .A(x[1419]), .B(n4563), .Z(n4565) );
  XOR U5985 ( .A(n4566), .B(n4567), .Z(n4563) );
  AND U5986 ( .A(n4568), .B(n4569), .Z(n4566) );
  XNOR U5987 ( .A(x[1418]), .B(n4567), .Z(n4569) );
  XOR U5988 ( .A(n4570), .B(n4571), .Z(n4567) );
  AND U5989 ( .A(n4572), .B(n4573), .Z(n4570) );
  XNOR U5990 ( .A(x[1417]), .B(n4571), .Z(n4573) );
  XOR U5991 ( .A(n4574), .B(n4575), .Z(n4571) );
  AND U5992 ( .A(n4576), .B(n4577), .Z(n4574) );
  XNOR U5993 ( .A(x[1416]), .B(n4575), .Z(n4577) );
  XOR U5994 ( .A(n4578), .B(n4579), .Z(n4575) );
  AND U5995 ( .A(n4580), .B(n4581), .Z(n4578) );
  XNOR U5996 ( .A(x[1415]), .B(n4579), .Z(n4581) );
  XOR U5997 ( .A(n4582), .B(n4583), .Z(n4579) );
  AND U5998 ( .A(n4584), .B(n4585), .Z(n4582) );
  XNOR U5999 ( .A(x[1414]), .B(n4583), .Z(n4585) );
  XOR U6000 ( .A(n4586), .B(n4587), .Z(n4583) );
  AND U6001 ( .A(n4588), .B(n4589), .Z(n4586) );
  XNOR U6002 ( .A(x[1413]), .B(n4587), .Z(n4589) );
  XOR U6003 ( .A(n4590), .B(n4591), .Z(n4587) );
  AND U6004 ( .A(n4592), .B(n4593), .Z(n4590) );
  XNOR U6005 ( .A(x[1412]), .B(n4591), .Z(n4593) );
  XOR U6006 ( .A(n4594), .B(n4595), .Z(n4591) );
  AND U6007 ( .A(n4596), .B(n4597), .Z(n4594) );
  XNOR U6008 ( .A(x[1411]), .B(n4595), .Z(n4597) );
  XOR U6009 ( .A(n4598), .B(n4599), .Z(n4595) );
  AND U6010 ( .A(n4600), .B(n4601), .Z(n4598) );
  XNOR U6011 ( .A(x[1410]), .B(n4599), .Z(n4601) );
  XOR U6012 ( .A(n4602), .B(n4603), .Z(n4599) );
  AND U6013 ( .A(n4604), .B(n4605), .Z(n4602) );
  XNOR U6014 ( .A(x[1409]), .B(n4603), .Z(n4605) );
  XOR U6015 ( .A(n4606), .B(n4607), .Z(n4603) );
  AND U6016 ( .A(n4608), .B(n4609), .Z(n4606) );
  XNOR U6017 ( .A(x[1408]), .B(n4607), .Z(n4609) );
  XOR U6018 ( .A(n4610), .B(n4611), .Z(n4607) );
  AND U6019 ( .A(n4612), .B(n4613), .Z(n4610) );
  XNOR U6020 ( .A(x[1407]), .B(n4611), .Z(n4613) );
  XOR U6021 ( .A(n4614), .B(n4615), .Z(n4611) );
  AND U6022 ( .A(n4616), .B(n4617), .Z(n4614) );
  XNOR U6023 ( .A(x[1406]), .B(n4615), .Z(n4617) );
  XOR U6024 ( .A(n4618), .B(n4619), .Z(n4615) );
  AND U6025 ( .A(n4620), .B(n4621), .Z(n4618) );
  XNOR U6026 ( .A(x[1405]), .B(n4619), .Z(n4621) );
  XOR U6027 ( .A(n4622), .B(n4623), .Z(n4619) );
  AND U6028 ( .A(n4624), .B(n4625), .Z(n4622) );
  XNOR U6029 ( .A(x[1404]), .B(n4623), .Z(n4625) );
  XOR U6030 ( .A(n4626), .B(n4627), .Z(n4623) );
  AND U6031 ( .A(n4628), .B(n4629), .Z(n4626) );
  XNOR U6032 ( .A(x[1403]), .B(n4627), .Z(n4629) );
  XOR U6033 ( .A(n4630), .B(n4631), .Z(n4627) );
  AND U6034 ( .A(n4632), .B(n4633), .Z(n4630) );
  XNOR U6035 ( .A(x[1402]), .B(n4631), .Z(n4633) );
  XOR U6036 ( .A(n4634), .B(n4635), .Z(n4631) );
  AND U6037 ( .A(n4636), .B(n4637), .Z(n4634) );
  XNOR U6038 ( .A(x[1401]), .B(n4635), .Z(n4637) );
  XOR U6039 ( .A(n4638), .B(n4639), .Z(n4635) );
  AND U6040 ( .A(n4640), .B(n4641), .Z(n4638) );
  XNOR U6041 ( .A(x[1400]), .B(n4639), .Z(n4641) );
  XOR U6042 ( .A(n4642), .B(n4643), .Z(n4639) );
  AND U6043 ( .A(n4644), .B(n4645), .Z(n4642) );
  XNOR U6044 ( .A(x[1399]), .B(n4643), .Z(n4645) );
  XOR U6045 ( .A(n4646), .B(n4647), .Z(n4643) );
  AND U6046 ( .A(n4648), .B(n4649), .Z(n4646) );
  XNOR U6047 ( .A(x[1398]), .B(n4647), .Z(n4649) );
  XOR U6048 ( .A(n4650), .B(n4651), .Z(n4647) );
  AND U6049 ( .A(n4652), .B(n4653), .Z(n4650) );
  XNOR U6050 ( .A(x[1397]), .B(n4651), .Z(n4653) );
  XOR U6051 ( .A(n4654), .B(n4655), .Z(n4651) );
  AND U6052 ( .A(n4656), .B(n4657), .Z(n4654) );
  XNOR U6053 ( .A(x[1396]), .B(n4655), .Z(n4657) );
  XOR U6054 ( .A(n4658), .B(n4659), .Z(n4655) );
  AND U6055 ( .A(n4660), .B(n4661), .Z(n4658) );
  XNOR U6056 ( .A(x[1395]), .B(n4659), .Z(n4661) );
  XOR U6057 ( .A(n4662), .B(n4663), .Z(n4659) );
  AND U6058 ( .A(n4664), .B(n4665), .Z(n4662) );
  XNOR U6059 ( .A(x[1394]), .B(n4663), .Z(n4665) );
  XOR U6060 ( .A(n4666), .B(n4667), .Z(n4663) );
  AND U6061 ( .A(n4668), .B(n4669), .Z(n4666) );
  XNOR U6062 ( .A(x[1393]), .B(n4667), .Z(n4669) );
  XOR U6063 ( .A(n4670), .B(n4671), .Z(n4667) );
  AND U6064 ( .A(n4672), .B(n4673), .Z(n4670) );
  XNOR U6065 ( .A(x[1392]), .B(n4671), .Z(n4673) );
  XOR U6066 ( .A(n4674), .B(n4675), .Z(n4671) );
  AND U6067 ( .A(n4676), .B(n4677), .Z(n4674) );
  XNOR U6068 ( .A(x[1391]), .B(n4675), .Z(n4677) );
  XOR U6069 ( .A(n4678), .B(n4679), .Z(n4675) );
  AND U6070 ( .A(n4680), .B(n4681), .Z(n4678) );
  XNOR U6071 ( .A(x[1390]), .B(n4679), .Z(n4681) );
  XOR U6072 ( .A(n4682), .B(n4683), .Z(n4679) );
  AND U6073 ( .A(n4684), .B(n4685), .Z(n4682) );
  XNOR U6074 ( .A(x[1389]), .B(n4683), .Z(n4685) );
  XOR U6075 ( .A(n4686), .B(n4687), .Z(n4683) );
  AND U6076 ( .A(n4688), .B(n4689), .Z(n4686) );
  XNOR U6077 ( .A(x[1388]), .B(n4687), .Z(n4689) );
  XOR U6078 ( .A(n4690), .B(n4691), .Z(n4687) );
  AND U6079 ( .A(n4692), .B(n4693), .Z(n4690) );
  XNOR U6080 ( .A(x[1387]), .B(n4691), .Z(n4693) );
  XOR U6081 ( .A(n4694), .B(n4695), .Z(n4691) );
  AND U6082 ( .A(n4696), .B(n4697), .Z(n4694) );
  XNOR U6083 ( .A(x[1386]), .B(n4695), .Z(n4697) );
  XOR U6084 ( .A(n4698), .B(n4699), .Z(n4695) );
  AND U6085 ( .A(n4700), .B(n4701), .Z(n4698) );
  XNOR U6086 ( .A(x[1385]), .B(n4699), .Z(n4701) );
  XOR U6087 ( .A(n4702), .B(n4703), .Z(n4699) );
  AND U6088 ( .A(n4704), .B(n4705), .Z(n4702) );
  XNOR U6089 ( .A(x[1384]), .B(n4703), .Z(n4705) );
  XOR U6090 ( .A(n4706), .B(n4707), .Z(n4703) );
  AND U6091 ( .A(n4708), .B(n4709), .Z(n4706) );
  XNOR U6092 ( .A(x[1383]), .B(n4707), .Z(n4709) );
  XOR U6093 ( .A(n4710), .B(n4711), .Z(n4707) );
  AND U6094 ( .A(n4712), .B(n4713), .Z(n4710) );
  XNOR U6095 ( .A(x[1382]), .B(n4711), .Z(n4713) );
  XOR U6096 ( .A(n4714), .B(n4715), .Z(n4711) );
  AND U6097 ( .A(n4716), .B(n4717), .Z(n4714) );
  XNOR U6098 ( .A(x[1381]), .B(n4715), .Z(n4717) );
  XOR U6099 ( .A(n4718), .B(n4719), .Z(n4715) );
  AND U6100 ( .A(n4720), .B(n4721), .Z(n4718) );
  XNOR U6101 ( .A(x[1380]), .B(n4719), .Z(n4721) );
  XOR U6102 ( .A(n4722), .B(n4723), .Z(n4719) );
  AND U6103 ( .A(n4724), .B(n4725), .Z(n4722) );
  XNOR U6104 ( .A(x[1379]), .B(n4723), .Z(n4725) );
  XOR U6105 ( .A(n4726), .B(n4727), .Z(n4723) );
  AND U6106 ( .A(n4728), .B(n4729), .Z(n4726) );
  XNOR U6107 ( .A(x[1378]), .B(n4727), .Z(n4729) );
  XOR U6108 ( .A(n4730), .B(n4731), .Z(n4727) );
  AND U6109 ( .A(n4732), .B(n4733), .Z(n4730) );
  XNOR U6110 ( .A(x[1377]), .B(n4731), .Z(n4733) );
  XOR U6111 ( .A(n4734), .B(n4735), .Z(n4731) );
  AND U6112 ( .A(n4736), .B(n4737), .Z(n4734) );
  XNOR U6113 ( .A(x[1376]), .B(n4735), .Z(n4737) );
  XOR U6114 ( .A(n4738), .B(n4739), .Z(n4735) );
  AND U6115 ( .A(n4740), .B(n4741), .Z(n4738) );
  XNOR U6116 ( .A(x[1375]), .B(n4739), .Z(n4741) );
  XOR U6117 ( .A(n4742), .B(n4743), .Z(n4739) );
  AND U6118 ( .A(n4744), .B(n4745), .Z(n4742) );
  XNOR U6119 ( .A(x[1374]), .B(n4743), .Z(n4745) );
  XOR U6120 ( .A(n4746), .B(n4747), .Z(n4743) );
  AND U6121 ( .A(n4748), .B(n4749), .Z(n4746) );
  XNOR U6122 ( .A(x[1373]), .B(n4747), .Z(n4749) );
  XOR U6123 ( .A(n4750), .B(n4751), .Z(n4747) );
  AND U6124 ( .A(n4752), .B(n4753), .Z(n4750) );
  XNOR U6125 ( .A(x[1372]), .B(n4751), .Z(n4753) );
  XOR U6126 ( .A(n4754), .B(n4755), .Z(n4751) );
  AND U6127 ( .A(n4756), .B(n4757), .Z(n4754) );
  XNOR U6128 ( .A(x[1371]), .B(n4755), .Z(n4757) );
  XOR U6129 ( .A(n4758), .B(n4759), .Z(n4755) );
  AND U6130 ( .A(n4760), .B(n4761), .Z(n4758) );
  XNOR U6131 ( .A(x[1370]), .B(n4759), .Z(n4761) );
  XOR U6132 ( .A(n4762), .B(n4763), .Z(n4759) );
  AND U6133 ( .A(n4764), .B(n4765), .Z(n4762) );
  XNOR U6134 ( .A(x[1369]), .B(n4763), .Z(n4765) );
  XOR U6135 ( .A(n4766), .B(n4767), .Z(n4763) );
  AND U6136 ( .A(n4768), .B(n4769), .Z(n4766) );
  XNOR U6137 ( .A(x[1368]), .B(n4767), .Z(n4769) );
  XOR U6138 ( .A(n4770), .B(n4771), .Z(n4767) );
  AND U6139 ( .A(n4772), .B(n4773), .Z(n4770) );
  XNOR U6140 ( .A(x[1367]), .B(n4771), .Z(n4773) );
  XOR U6141 ( .A(n4774), .B(n4775), .Z(n4771) );
  AND U6142 ( .A(n4776), .B(n4777), .Z(n4774) );
  XNOR U6143 ( .A(x[1366]), .B(n4775), .Z(n4777) );
  XOR U6144 ( .A(n4778), .B(n4779), .Z(n4775) );
  AND U6145 ( .A(n4780), .B(n4781), .Z(n4778) );
  XNOR U6146 ( .A(x[1365]), .B(n4779), .Z(n4781) );
  XOR U6147 ( .A(n4782), .B(n4783), .Z(n4779) );
  AND U6148 ( .A(n4784), .B(n4785), .Z(n4782) );
  XNOR U6149 ( .A(x[1364]), .B(n4783), .Z(n4785) );
  XOR U6150 ( .A(n4786), .B(n4787), .Z(n4783) );
  AND U6151 ( .A(n4788), .B(n4789), .Z(n4786) );
  XNOR U6152 ( .A(x[1363]), .B(n4787), .Z(n4789) );
  XOR U6153 ( .A(n4790), .B(n4791), .Z(n4787) );
  AND U6154 ( .A(n4792), .B(n4793), .Z(n4790) );
  XNOR U6155 ( .A(x[1362]), .B(n4791), .Z(n4793) );
  XOR U6156 ( .A(n4794), .B(n4795), .Z(n4791) );
  AND U6157 ( .A(n4796), .B(n4797), .Z(n4794) );
  XNOR U6158 ( .A(x[1361]), .B(n4795), .Z(n4797) );
  XOR U6159 ( .A(n4798), .B(n4799), .Z(n4795) );
  AND U6160 ( .A(n4800), .B(n4801), .Z(n4798) );
  XNOR U6161 ( .A(x[1360]), .B(n4799), .Z(n4801) );
  XOR U6162 ( .A(n4802), .B(n4803), .Z(n4799) );
  AND U6163 ( .A(n4804), .B(n4805), .Z(n4802) );
  XNOR U6164 ( .A(x[1359]), .B(n4803), .Z(n4805) );
  XOR U6165 ( .A(n4806), .B(n4807), .Z(n4803) );
  AND U6166 ( .A(n4808), .B(n4809), .Z(n4806) );
  XNOR U6167 ( .A(x[1358]), .B(n4807), .Z(n4809) );
  XOR U6168 ( .A(n4810), .B(n4811), .Z(n4807) );
  AND U6169 ( .A(n4812), .B(n4813), .Z(n4810) );
  XNOR U6170 ( .A(x[1357]), .B(n4811), .Z(n4813) );
  XOR U6171 ( .A(n4814), .B(n4815), .Z(n4811) );
  AND U6172 ( .A(n4816), .B(n4817), .Z(n4814) );
  XNOR U6173 ( .A(x[1356]), .B(n4815), .Z(n4817) );
  XOR U6174 ( .A(n4818), .B(n4819), .Z(n4815) );
  AND U6175 ( .A(n4820), .B(n4821), .Z(n4818) );
  XNOR U6176 ( .A(x[1355]), .B(n4819), .Z(n4821) );
  XOR U6177 ( .A(n4822), .B(n4823), .Z(n4819) );
  AND U6178 ( .A(n4824), .B(n4825), .Z(n4822) );
  XNOR U6179 ( .A(x[1354]), .B(n4823), .Z(n4825) );
  XOR U6180 ( .A(n4826), .B(n4827), .Z(n4823) );
  AND U6181 ( .A(n4828), .B(n4829), .Z(n4826) );
  XNOR U6182 ( .A(x[1353]), .B(n4827), .Z(n4829) );
  XOR U6183 ( .A(n4830), .B(n4831), .Z(n4827) );
  AND U6184 ( .A(n4832), .B(n4833), .Z(n4830) );
  XNOR U6185 ( .A(x[1352]), .B(n4831), .Z(n4833) );
  XOR U6186 ( .A(n4834), .B(n4835), .Z(n4831) );
  AND U6187 ( .A(n4836), .B(n4837), .Z(n4834) );
  XNOR U6188 ( .A(x[1351]), .B(n4835), .Z(n4837) );
  XOR U6189 ( .A(n4838), .B(n4839), .Z(n4835) );
  AND U6190 ( .A(n4840), .B(n4841), .Z(n4838) );
  XNOR U6191 ( .A(x[1350]), .B(n4839), .Z(n4841) );
  XOR U6192 ( .A(n4842), .B(n4843), .Z(n4839) );
  AND U6193 ( .A(n4844), .B(n4845), .Z(n4842) );
  XNOR U6194 ( .A(x[1349]), .B(n4843), .Z(n4845) );
  XOR U6195 ( .A(n4846), .B(n4847), .Z(n4843) );
  AND U6196 ( .A(n4848), .B(n4849), .Z(n4846) );
  XNOR U6197 ( .A(x[1348]), .B(n4847), .Z(n4849) );
  XOR U6198 ( .A(n4850), .B(n4851), .Z(n4847) );
  AND U6199 ( .A(n4852), .B(n4853), .Z(n4850) );
  XNOR U6200 ( .A(x[1347]), .B(n4851), .Z(n4853) );
  XOR U6201 ( .A(n4854), .B(n4855), .Z(n4851) );
  AND U6202 ( .A(n4856), .B(n4857), .Z(n4854) );
  XNOR U6203 ( .A(x[1346]), .B(n4855), .Z(n4857) );
  XOR U6204 ( .A(n4858), .B(n4859), .Z(n4855) );
  AND U6205 ( .A(n4860), .B(n4861), .Z(n4858) );
  XNOR U6206 ( .A(x[1345]), .B(n4859), .Z(n4861) );
  XOR U6207 ( .A(n4862), .B(n4863), .Z(n4859) );
  AND U6208 ( .A(n4864), .B(n4865), .Z(n4862) );
  XNOR U6209 ( .A(x[1344]), .B(n4863), .Z(n4865) );
  XOR U6210 ( .A(n4866), .B(n4867), .Z(n4863) );
  AND U6211 ( .A(n4868), .B(n4869), .Z(n4866) );
  XNOR U6212 ( .A(x[1343]), .B(n4867), .Z(n4869) );
  XOR U6213 ( .A(n4870), .B(n4871), .Z(n4867) );
  AND U6214 ( .A(n4872), .B(n4873), .Z(n4870) );
  XNOR U6215 ( .A(x[1342]), .B(n4871), .Z(n4873) );
  XOR U6216 ( .A(n4874), .B(n4875), .Z(n4871) );
  AND U6217 ( .A(n4876), .B(n4877), .Z(n4874) );
  XNOR U6218 ( .A(x[1341]), .B(n4875), .Z(n4877) );
  XOR U6219 ( .A(n4878), .B(n4879), .Z(n4875) );
  AND U6220 ( .A(n4880), .B(n4881), .Z(n4878) );
  XNOR U6221 ( .A(x[1340]), .B(n4879), .Z(n4881) );
  XOR U6222 ( .A(n4882), .B(n4883), .Z(n4879) );
  AND U6223 ( .A(n4884), .B(n4885), .Z(n4882) );
  XNOR U6224 ( .A(x[1339]), .B(n4883), .Z(n4885) );
  XOR U6225 ( .A(n4886), .B(n4887), .Z(n4883) );
  AND U6226 ( .A(n4888), .B(n4889), .Z(n4886) );
  XNOR U6227 ( .A(x[1338]), .B(n4887), .Z(n4889) );
  XOR U6228 ( .A(n4890), .B(n4891), .Z(n4887) );
  AND U6229 ( .A(n4892), .B(n4893), .Z(n4890) );
  XNOR U6230 ( .A(x[1337]), .B(n4891), .Z(n4893) );
  XOR U6231 ( .A(n4894), .B(n4895), .Z(n4891) );
  AND U6232 ( .A(n4896), .B(n4897), .Z(n4894) );
  XNOR U6233 ( .A(x[1336]), .B(n4895), .Z(n4897) );
  XOR U6234 ( .A(n4898), .B(n4899), .Z(n4895) );
  AND U6235 ( .A(n4900), .B(n4901), .Z(n4898) );
  XNOR U6236 ( .A(x[1335]), .B(n4899), .Z(n4901) );
  XOR U6237 ( .A(n4902), .B(n4903), .Z(n4899) );
  AND U6238 ( .A(n4904), .B(n4905), .Z(n4902) );
  XNOR U6239 ( .A(x[1334]), .B(n4903), .Z(n4905) );
  XOR U6240 ( .A(n4906), .B(n4907), .Z(n4903) );
  AND U6241 ( .A(n4908), .B(n4909), .Z(n4906) );
  XNOR U6242 ( .A(x[1333]), .B(n4907), .Z(n4909) );
  XOR U6243 ( .A(n4910), .B(n4911), .Z(n4907) );
  AND U6244 ( .A(n4912), .B(n4913), .Z(n4910) );
  XNOR U6245 ( .A(x[1332]), .B(n4911), .Z(n4913) );
  XOR U6246 ( .A(n4914), .B(n4915), .Z(n4911) );
  AND U6247 ( .A(n4916), .B(n4917), .Z(n4914) );
  XNOR U6248 ( .A(x[1331]), .B(n4915), .Z(n4917) );
  XOR U6249 ( .A(n4918), .B(n4919), .Z(n4915) );
  AND U6250 ( .A(n4920), .B(n4921), .Z(n4918) );
  XNOR U6251 ( .A(x[1330]), .B(n4919), .Z(n4921) );
  XOR U6252 ( .A(n4922), .B(n4923), .Z(n4919) );
  AND U6253 ( .A(n4924), .B(n4925), .Z(n4922) );
  XNOR U6254 ( .A(x[1329]), .B(n4923), .Z(n4925) );
  XOR U6255 ( .A(n4926), .B(n4927), .Z(n4923) );
  AND U6256 ( .A(n4928), .B(n4929), .Z(n4926) );
  XNOR U6257 ( .A(x[1328]), .B(n4927), .Z(n4929) );
  XOR U6258 ( .A(n4930), .B(n4931), .Z(n4927) );
  AND U6259 ( .A(n4932), .B(n4933), .Z(n4930) );
  XNOR U6260 ( .A(x[1327]), .B(n4931), .Z(n4933) );
  XOR U6261 ( .A(n4934), .B(n4935), .Z(n4931) );
  AND U6262 ( .A(n4936), .B(n4937), .Z(n4934) );
  XNOR U6263 ( .A(x[1326]), .B(n4935), .Z(n4937) );
  XOR U6264 ( .A(n4938), .B(n4939), .Z(n4935) );
  AND U6265 ( .A(n4940), .B(n4941), .Z(n4938) );
  XNOR U6266 ( .A(x[1325]), .B(n4939), .Z(n4941) );
  XOR U6267 ( .A(n4942), .B(n4943), .Z(n4939) );
  AND U6268 ( .A(n4944), .B(n4945), .Z(n4942) );
  XNOR U6269 ( .A(x[1324]), .B(n4943), .Z(n4945) );
  XOR U6270 ( .A(n4946), .B(n4947), .Z(n4943) );
  AND U6271 ( .A(n4948), .B(n4949), .Z(n4946) );
  XNOR U6272 ( .A(x[1323]), .B(n4947), .Z(n4949) );
  XOR U6273 ( .A(n4950), .B(n4951), .Z(n4947) );
  AND U6274 ( .A(n4952), .B(n4953), .Z(n4950) );
  XNOR U6275 ( .A(x[1322]), .B(n4951), .Z(n4953) );
  XOR U6276 ( .A(n4954), .B(n4955), .Z(n4951) );
  AND U6277 ( .A(n4956), .B(n4957), .Z(n4954) );
  XNOR U6278 ( .A(x[1321]), .B(n4955), .Z(n4957) );
  XOR U6279 ( .A(n4958), .B(n4959), .Z(n4955) );
  AND U6280 ( .A(n4960), .B(n4961), .Z(n4958) );
  XNOR U6281 ( .A(x[1320]), .B(n4959), .Z(n4961) );
  XOR U6282 ( .A(n4962), .B(n4963), .Z(n4959) );
  AND U6283 ( .A(n4964), .B(n4965), .Z(n4962) );
  XNOR U6284 ( .A(x[1319]), .B(n4963), .Z(n4965) );
  XOR U6285 ( .A(n4966), .B(n4967), .Z(n4963) );
  AND U6286 ( .A(n4968), .B(n4969), .Z(n4966) );
  XNOR U6287 ( .A(x[1318]), .B(n4967), .Z(n4969) );
  XOR U6288 ( .A(n4970), .B(n4971), .Z(n4967) );
  AND U6289 ( .A(n4972), .B(n4973), .Z(n4970) );
  XNOR U6290 ( .A(x[1317]), .B(n4971), .Z(n4973) );
  XOR U6291 ( .A(n4974), .B(n4975), .Z(n4971) );
  AND U6292 ( .A(n4976), .B(n4977), .Z(n4974) );
  XNOR U6293 ( .A(x[1316]), .B(n4975), .Z(n4977) );
  XOR U6294 ( .A(n4978), .B(n4979), .Z(n4975) );
  AND U6295 ( .A(n4980), .B(n4981), .Z(n4978) );
  XNOR U6296 ( .A(x[1315]), .B(n4979), .Z(n4981) );
  XOR U6297 ( .A(n4982), .B(n4983), .Z(n4979) );
  AND U6298 ( .A(n4984), .B(n4985), .Z(n4982) );
  XNOR U6299 ( .A(x[1314]), .B(n4983), .Z(n4985) );
  XOR U6300 ( .A(n4986), .B(n4987), .Z(n4983) );
  AND U6301 ( .A(n4988), .B(n4989), .Z(n4986) );
  XNOR U6302 ( .A(x[1313]), .B(n4987), .Z(n4989) );
  XOR U6303 ( .A(n4990), .B(n4991), .Z(n4987) );
  AND U6304 ( .A(n4992), .B(n4993), .Z(n4990) );
  XNOR U6305 ( .A(x[1312]), .B(n4991), .Z(n4993) );
  XOR U6306 ( .A(n4994), .B(n4995), .Z(n4991) );
  AND U6307 ( .A(n4996), .B(n4997), .Z(n4994) );
  XNOR U6308 ( .A(x[1311]), .B(n4995), .Z(n4997) );
  XOR U6309 ( .A(n4998), .B(n4999), .Z(n4995) );
  AND U6310 ( .A(n5000), .B(n5001), .Z(n4998) );
  XNOR U6311 ( .A(x[1310]), .B(n4999), .Z(n5001) );
  XOR U6312 ( .A(n5002), .B(n5003), .Z(n4999) );
  AND U6313 ( .A(n5004), .B(n5005), .Z(n5002) );
  XNOR U6314 ( .A(x[1309]), .B(n5003), .Z(n5005) );
  XOR U6315 ( .A(n5006), .B(n5007), .Z(n5003) );
  AND U6316 ( .A(n5008), .B(n5009), .Z(n5006) );
  XNOR U6317 ( .A(x[1308]), .B(n5007), .Z(n5009) );
  XOR U6318 ( .A(n5010), .B(n5011), .Z(n5007) );
  AND U6319 ( .A(n5012), .B(n5013), .Z(n5010) );
  XNOR U6320 ( .A(x[1307]), .B(n5011), .Z(n5013) );
  XOR U6321 ( .A(n5014), .B(n5015), .Z(n5011) );
  AND U6322 ( .A(n5016), .B(n5017), .Z(n5014) );
  XNOR U6323 ( .A(x[1306]), .B(n5015), .Z(n5017) );
  XOR U6324 ( .A(n5018), .B(n5019), .Z(n5015) );
  AND U6325 ( .A(n5020), .B(n5021), .Z(n5018) );
  XNOR U6326 ( .A(x[1305]), .B(n5019), .Z(n5021) );
  XOR U6327 ( .A(n5022), .B(n5023), .Z(n5019) );
  AND U6328 ( .A(n5024), .B(n5025), .Z(n5022) );
  XNOR U6329 ( .A(x[1304]), .B(n5023), .Z(n5025) );
  XOR U6330 ( .A(n5026), .B(n5027), .Z(n5023) );
  AND U6331 ( .A(n5028), .B(n5029), .Z(n5026) );
  XNOR U6332 ( .A(x[1303]), .B(n5027), .Z(n5029) );
  XOR U6333 ( .A(n5030), .B(n5031), .Z(n5027) );
  AND U6334 ( .A(n5032), .B(n5033), .Z(n5030) );
  XNOR U6335 ( .A(x[1302]), .B(n5031), .Z(n5033) );
  XOR U6336 ( .A(n5034), .B(n5035), .Z(n5031) );
  AND U6337 ( .A(n5036), .B(n5037), .Z(n5034) );
  XNOR U6338 ( .A(x[1301]), .B(n5035), .Z(n5037) );
  XOR U6339 ( .A(n5038), .B(n5039), .Z(n5035) );
  AND U6340 ( .A(n5040), .B(n5041), .Z(n5038) );
  XNOR U6341 ( .A(x[1300]), .B(n5039), .Z(n5041) );
  XOR U6342 ( .A(n5042), .B(n5043), .Z(n5039) );
  AND U6343 ( .A(n5044), .B(n5045), .Z(n5042) );
  XNOR U6344 ( .A(x[1299]), .B(n5043), .Z(n5045) );
  XOR U6345 ( .A(n5046), .B(n5047), .Z(n5043) );
  AND U6346 ( .A(n5048), .B(n5049), .Z(n5046) );
  XNOR U6347 ( .A(x[1298]), .B(n5047), .Z(n5049) );
  XOR U6348 ( .A(n5050), .B(n5051), .Z(n5047) );
  AND U6349 ( .A(n5052), .B(n5053), .Z(n5050) );
  XNOR U6350 ( .A(x[1297]), .B(n5051), .Z(n5053) );
  XOR U6351 ( .A(n5054), .B(n5055), .Z(n5051) );
  AND U6352 ( .A(n5056), .B(n5057), .Z(n5054) );
  XNOR U6353 ( .A(x[1296]), .B(n5055), .Z(n5057) );
  XOR U6354 ( .A(n5058), .B(n5059), .Z(n5055) );
  AND U6355 ( .A(n5060), .B(n5061), .Z(n5058) );
  XNOR U6356 ( .A(x[1295]), .B(n5059), .Z(n5061) );
  XOR U6357 ( .A(n5062), .B(n5063), .Z(n5059) );
  AND U6358 ( .A(n5064), .B(n5065), .Z(n5062) );
  XNOR U6359 ( .A(x[1294]), .B(n5063), .Z(n5065) );
  XOR U6360 ( .A(n5066), .B(n5067), .Z(n5063) );
  AND U6361 ( .A(n5068), .B(n5069), .Z(n5066) );
  XNOR U6362 ( .A(x[1293]), .B(n5067), .Z(n5069) );
  XOR U6363 ( .A(n5070), .B(n5071), .Z(n5067) );
  AND U6364 ( .A(n5072), .B(n5073), .Z(n5070) );
  XNOR U6365 ( .A(x[1292]), .B(n5071), .Z(n5073) );
  XOR U6366 ( .A(n5074), .B(n5075), .Z(n5071) );
  AND U6367 ( .A(n5076), .B(n5077), .Z(n5074) );
  XNOR U6368 ( .A(x[1291]), .B(n5075), .Z(n5077) );
  XOR U6369 ( .A(n5078), .B(n5079), .Z(n5075) );
  AND U6370 ( .A(n5080), .B(n5081), .Z(n5078) );
  XNOR U6371 ( .A(x[1290]), .B(n5079), .Z(n5081) );
  XOR U6372 ( .A(n5082), .B(n5083), .Z(n5079) );
  AND U6373 ( .A(n5084), .B(n5085), .Z(n5082) );
  XNOR U6374 ( .A(x[1289]), .B(n5083), .Z(n5085) );
  XOR U6375 ( .A(n5086), .B(n5087), .Z(n5083) );
  AND U6376 ( .A(n5088), .B(n5089), .Z(n5086) );
  XNOR U6377 ( .A(x[1288]), .B(n5087), .Z(n5089) );
  XOR U6378 ( .A(n5090), .B(n5091), .Z(n5087) );
  AND U6379 ( .A(n5092), .B(n5093), .Z(n5090) );
  XNOR U6380 ( .A(x[1287]), .B(n5091), .Z(n5093) );
  XOR U6381 ( .A(n5094), .B(n5095), .Z(n5091) );
  AND U6382 ( .A(n5096), .B(n5097), .Z(n5094) );
  XNOR U6383 ( .A(x[1286]), .B(n5095), .Z(n5097) );
  XOR U6384 ( .A(n5098), .B(n5099), .Z(n5095) );
  AND U6385 ( .A(n5100), .B(n5101), .Z(n5098) );
  XNOR U6386 ( .A(x[1285]), .B(n5099), .Z(n5101) );
  XOR U6387 ( .A(n5102), .B(n5103), .Z(n5099) );
  AND U6388 ( .A(n5104), .B(n5105), .Z(n5102) );
  XNOR U6389 ( .A(x[1284]), .B(n5103), .Z(n5105) );
  XOR U6390 ( .A(n5106), .B(n5107), .Z(n5103) );
  AND U6391 ( .A(n5108), .B(n5109), .Z(n5106) );
  XNOR U6392 ( .A(x[1283]), .B(n5107), .Z(n5109) );
  XOR U6393 ( .A(n5110), .B(n5111), .Z(n5107) );
  AND U6394 ( .A(n5112), .B(n5113), .Z(n5110) );
  XNOR U6395 ( .A(x[1282]), .B(n5111), .Z(n5113) );
  XOR U6396 ( .A(n5114), .B(n5115), .Z(n5111) );
  AND U6397 ( .A(n5116), .B(n5117), .Z(n5114) );
  XNOR U6398 ( .A(x[1281]), .B(n5115), .Z(n5117) );
  XOR U6399 ( .A(n5118), .B(n5119), .Z(n5115) );
  AND U6400 ( .A(n5120), .B(n5121), .Z(n5118) );
  XNOR U6401 ( .A(x[1280]), .B(n5119), .Z(n5121) );
  XOR U6402 ( .A(n5122), .B(n5123), .Z(n5119) );
  AND U6403 ( .A(n5124), .B(n5125), .Z(n5122) );
  XNOR U6404 ( .A(x[1279]), .B(n5123), .Z(n5125) );
  XOR U6405 ( .A(n5126), .B(n5127), .Z(n5123) );
  AND U6406 ( .A(n5128), .B(n5129), .Z(n5126) );
  XNOR U6407 ( .A(x[1278]), .B(n5127), .Z(n5129) );
  XOR U6408 ( .A(n5130), .B(n5131), .Z(n5127) );
  AND U6409 ( .A(n5132), .B(n5133), .Z(n5130) );
  XNOR U6410 ( .A(x[1277]), .B(n5131), .Z(n5133) );
  XOR U6411 ( .A(n5134), .B(n5135), .Z(n5131) );
  AND U6412 ( .A(n5136), .B(n5137), .Z(n5134) );
  XNOR U6413 ( .A(x[1276]), .B(n5135), .Z(n5137) );
  XOR U6414 ( .A(n5138), .B(n5139), .Z(n5135) );
  AND U6415 ( .A(n5140), .B(n5141), .Z(n5138) );
  XNOR U6416 ( .A(x[1275]), .B(n5139), .Z(n5141) );
  XOR U6417 ( .A(n5142), .B(n5143), .Z(n5139) );
  AND U6418 ( .A(n5144), .B(n5145), .Z(n5142) );
  XNOR U6419 ( .A(x[1274]), .B(n5143), .Z(n5145) );
  XOR U6420 ( .A(n5146), .B(n5147), .Z(n5143) );
  AND U6421 ( .A(n5148), .B(n5149), .Z(n5146) );
  XNOR U6422 ( .A(x[1273]), .B(n5147), .Z(n5149) );
  XOR U6423 ( .A(n5150), .B(n5151), .Z(n5147) );
  AND U6424 ( .A(n5152), .B(n5153), .Z(n5150) );
  XNOR U6425 ( .A(x[1272]), .B(n5151), .Z(n5153) );
  XOR U6426 ( .A(n5154), .B(n5155), .Z(n5151) );
  AND U6427 ( .A(n5156), .B(n5157), .Z(n5154) );
  XNOR U6428 ( .A(x[1271]), .B(n5155), .Z(n5157) );
  XOR U6429 ( .A(n5158), .B(n5159), .Z(n5155) );
  AND U6430 ( .A(n5160), .B(n5161), .Z(n5158) );
  XNOR U6431 ( .A(x[1270]), .B(n5159), .Z(n5161) );
  XOR U6432 ( .A(n5162), .B(n5163), .Z(n5159) );
  AND U6433 ( .A(n5164), .B(n5165), .Z(n5162) );
  XNOR U6434 ( .A(x[1269]), .B(n5163), .Z(n5165) );
  XOR U6435 ( .A(n5166), .B(n5167), .Z(n5163) );
  AND U6436 ( .A(n5168), .B(n5169), .Z(n5166) );
  XNOR U6437 ( .A(x[1268]), .B(n5167), .Z(n5169) );
  XOR U6438 ( .A(n5170), .B(n5171), .Z(n5167) );
  AND U6439 ( .A(n5172), .B(n5173), .Z(n5170) );
  XNOR U6440 ( .A(x[1267]), .B(n5171), .Z(n5173) );
  XOR U6441 ( .A(n5174), .B(n5175), .Z(n5171) );
  AND U6442 ( .A(n5176), .B(n5177), .Z(n5174) );
  XNOR U6443 ( .A(x[1266]), .B(n5175), .Z(n5177) );
  XOR U6444 ( .A(n5178), .B(n5179), .Z(n5175) );
  AND U6445 ( .A(n5180), .B(n5181), .Z(n5178) );
  XNOR U6446 ( .A(x[1265]), .B(n5179), .Z(n5181) );
  XOR U6447 ( .A(n5182), .B(n5183), .Z(n5179) );
  AND U6448 ( .A(n5184), .B(n5185), .Z(n5182) );
  XNOR U6449 ( .A(x[1264]), .B(n5183), .Z(n5185) );
  XOR U6450 ( .A(n5186), .B(n5187), .Z(n5183) );
  AND U6451 ( .A(n5188), .B(n5189), .Z(n5186) );
  XNOR U6452 ( .A(x[1263]), .B(n5187), .Z(n5189) );
  XOR U6453 ( .A(n5190), .B(n5191), .Z(n5187) );
  AND U6454 ( .A(n5192), .B(n5193), .Z(n5190) );
  XNOR U6455 ( .A(x[1262]), .B(n5191), .Z(n5193) );
  XOR U6456 ( .A(n5194), .B(n5195), .Z(n5191) );
  AND U6457 ( .A(n5196), .B(n5197), .Z(n5194) );
  XNOR U6458 ( .A(x[1261]), .B(n5195), .Z(n5197) );
  XOR U6459 ( .A(n5198), .B(n5199), .Z(n5195) );
  AND U6460 ( .A(n5200), .B(n5201), .Z(n5198) );
  XNOR U6461 ( .A(x[1260]), .B(n5199), .Z(n5201) );
  XOR U6462 ( .A(n5202), .B(n5203), .Z(n5199) );
  AND U6463 ( .A(n5204), .B(n5205), .Z(n5202) );
  XNOR U6464 ( .A(x[1259]), .B(n5203), .Z(n5205) );
  XOR U6465 ( .A(n5206), .B(n5207), .Z(n5203) );
  AND U6466 ( .A(n5208), .B(n5209), .Z(n5206) );
  XNOR U6467 ( .A(x[1258]), .B(n5207), .Z(n5209) );
  XOR U6468 ( .A(n5210), .B(n5211), .Z(n5207) );
  AND U6469 ( .A(n5212), .B(n5213), .Z(n5210) );
  XNOR U6470 ( .A(x[1257]), .B(n5211), .Z(n5213) );
  XOR U6471 ( .A(n5214), .B(n5215), .Z(n5211) );
  AND U6472 ( .A(n5216), .B(n5217), .Z(n5214) );
  XNOR U6473 ( .A(x[1256]), .B(n5215), .Z(n5217) );
  XOR U6474 ( .A(n5218), .B(n5219), .Z(n5215) );
  AND U6475 ( .A(n5220), .B(n5221), .Z(n5218) );
  XNOR U6476 ( .A(x[1255]), .B(n5219), .Z(n5221) );
  XOR U6477 ( .A(n5222), .B(n5223), .Z(n5219) );
  AND U6478 ( .A(n5224), .B(n5225), .Z(n5222) );
  XNOR U6479 ( .A(x[1254]), .B(n5223), .Z(n5225) );
  XOR U6480 ( .A(n5226), .B(n5227), .Z(n5223) );
  AND U6481 ( .A(n5228), .B(n5229), .Z(n5226) );
  XNOR U6482 ( .A(x[1253]), .B(n5227), .Z(n5229) );
  XOR U6483 ( .A(n5230), .B(n5231), .Z(n5227) );
  AND U6484 ( .A(n5232), .B(n5233), .Z(n5230) );
  XNOR U6485 ( .A(x[1252]), .B(n5231), .Z(n5233) );
  XOR U6486 ( .A(n5234), .B(n5235), .Z(n5231) );
  AND U6487 ( .A(n5236), .B(n5237), .Z(n5234) );
  XNOR U6488 ( .A(x[1251]), .B(n5235), .Z(n5237) );
  XOR U6489 ( .A(n5238), .B(n5239), .Z(n5235) );
  AND U6490 ( .A(n5240), .B(n5241), .Z(n5238) );
  XNOR U6491 ( .A(x[1250]), .B(n5239), .Z(n5241) );
  XOR U6492 ( .A(n5242), .B(n5243), .Z(n5239) );
  AND U6493 ( .A(n5244), .B(n5245), .Z(n5242) );
  XNOR U6494 ( .A(x[1249]), .B(n5243), .Z(n5245) );
  XOR U6495 ( .A(n5246), .B(n5247), .Z(n5243) );
  AND U6496 ( .A(n5248), .B(n5249), .Z(n5246) );
  XNOR U6497 ( .A(x[1248]), .B(n5247), .Z(n5249) );
  XOR U6498 ( .A(n5250), .B(n5251), .Z(n5247) );
  AND U6499 ( .A(n5252), .B(n5253), .Z(n5250) );
  XNOR U6500 ( .A(x[1247]), .B(n5251), .Z(n5253) );
  XOR U6501 ( .A(n5254), .B(n5255), .Z(n5251) );
  AND U6502 ( .A(n5256), .B(n5257), .Z(n5254) );
  XNOR U6503 ( .A(x[1246]), .B(n5255), .Z(n5257) );
  XOR U6504 ( .A(n5258), .B(n5259), .Z(n5255) );
  AND U6505 ( .A(n5260), .B(n5261), .Z(n5258) );
  XNOR U6506 ( .A(x[1245]), .B(n5259), .Z(n5261) );
  XOR U6507 ( .A(n5262), .B(n5263), .Z(n5259) );
  AND U6508 ( .A(n5264), .B(n5265), .Z(n5262) );
  XNOR U6509 ( .A(x[1244]), .B(n5263), .Z(n5265) );
  XOR U6510 ( .A(n5266), .B(n5267), .Z(n5263) );
  AND U6511 ( .A(n5268), .B(n5269), .Z(n5266) );
  XNOR U6512 ( .A(x[1243]), .B(n5267), .Z(n5269) );
  XOR U6513 ( .A(n5270), .B(n5271), .Z(n5267) );
  AND U6514 ( .A(n5272), .B(n5273), .Z(n5270) );
  XNOR U6515 ( .A(x[1242]), .B(n5271), .Z(n5273) );
  XOR U6516 ( .A(n5274), .B(n5275), .Z(n5271) );
  AND U6517 ( .A(n5276), .B(n5277), .Z(n5274) );
  XNOR U6518 ( .A(x[1241]), .B(n5275), .Z(n5277) );
  XOR U6519 ( .A(n5278), .B(n5279), .Z(n5275) );
  AND U6520 ( .A(n5280), .B(n5281), .Z(n5278) );
  XNOR U6521 ( .A(x[1240]), .B(n5279), .Z(n5281) );
  XOR U6522 ( .A(n5282), .B(n5283), .Z(n5279) );
  AND U6523 ( .A(n5284), .B(n5285), .Z(n5282) );
  XNOR U6524 ( .A(x[1239]), .B(n5283), .Z(n5285) );
  XOR U6525 ( .A(n5286), .B(n5287), .Z(n5283) );
  AND U6526 ( .A(n5288), .B(n5289), .Z(n5286) );
  XNOR U6527 ( .A(x[1238]), .B(n5287), .Z(n5289) );
  XOR U6528 ( .A(n5290), .B(n5291), .Z(n5287) );
  AND U6529 ( .A(n5292), .B(n5293), .Z(n5290) );
  XNOR U6530 ( .A(x[1237]), .B(n5291), .Z(n5293) );
  XOR U6531 ( .A(n5294), .B(n5295), .Z(n5291) );
  AND U6532 ( .A(n5296), .B(n5297), .Z(n5294) );
  XNOR U6533 ( .A(x[1236]), .B(n5295), .Z(n5297) );
  XOR U6534 ( .A(n5298), .B(n5299), .Z(n5295) );
  AND U6535 ( .A(n5300), .B(n5301), .Z(n5298) );
  XNOR U6536 ( .A(x[1235]), .B(n5299), .Z(n5301) );
  XOR U6537 ( .A(n5302), .B(n5303), .Z(n5299) );
  AND U6538 ( .A(n5304), .B(n5305), .Z(n5302) );
  XNOR U6539 ( .A(x[1234]), .B(n5303), .Z(n5305) );
  XOR U6540 ( .A(n5306), .B(n5307), .Z(n5303) );
  AND U6541 ( .A(n5308), .B(n5309), .Z(n5306) );
  XNOR U6542 ( .A(x[1233]), .B(n5307), .Z(n5309) );
  XOR U6543 ( .A(n5310), .B(n5311), .Z(n5307) );
  AND U6544 ( .A(n5312), .B(n5313), .Z(n5310) );
  XNOR U6545 ( .A(x[1232]), .B(n5311), .Z(n5313) );
  XOR U6546 ( .A(n5314), .B(n5315), .Z(n5311) );
  AND U6547 ( .A(n5316), .B(n5317), .Z(n5314) );
  XNOR U6548 ( .A(x[1231]), .B(n5315), .Z(n5317) );
  XOR U6549 ( .A(n5318), .B(n5319), .Z(n5315) );
  AND U6550 ( .A(n5320), .B(n5321), .Z(n5318) );
  XNOR U6551 ( .A(x[1230]), .B(n5319), .Z(n5321) );
  XOR U6552 ( .A(n5322), .B(n5323), .Z(n5319) );
  AND U6553 ( .A(n5324), .B(n5325), .Z(n5322) );
  XNOR U6554 ( .A(x[1229]), .B(n5323), .Z(n5325) );
  XOR U6555 ( .A(n5326), .B(n5327), .Z(n5323) );
  AND U6556 ( .A(n5328), .B(n5329), .Z(n5326) );
  XNOR U6557 ( .A(x[1228]), .B(n5327), .Z(n5329) );
  XOR U6558 ( .A(n5330), .B(n5331), .Z(n5327) );
  AND U6559 ( .A(n5332), .B(n5333), .Z(n5330) );
  XNOR U6560 ( .A(x[1227]), .B(n5331), .Z(n5333) );
  XOR U6561 ( .A(n5334), .B(n5335), .Z(n5331) );
  AND U6562 ( .A(n5336), .B(n5337), .Z(n5334) );
  XNOR U6563 ( .A(x[1226]), .B(n5335), .Z(n5337) );
  XOR U6564 ( .A(n5338), .B(n5339), .Z(n5335) );
  AND U6565 ( .A(n5340), .B(n5341), .Z(n5338) );
  XNOR U6566 ( .A(x[1225]), .B(n5339), .Z(n5341) );
  XOR U6567 ( .A(n5342), .B(n5343), .Z(n5339) );
  AND U6568 ( .A(n5344), .B(n5345), .Z(n5342) );
  XNOR U6569 ( .A(x[1224]), .B(n5343), .Z(n5345) );
  XOR U6570 ( .A(n5346), .B(n5347), .Z(n5343) );
  AND U6571 ( .A(n5348), .B(n5349), .Z(n5346) );
  XNOR U6572 ( .A(x[1223]), .B(n5347), .Z(n5349) );
  XOR U6573 ( .A(n5350), .B(n5351), .Z(n5347) );
  AND U6574 ( .A(n5352), .B(n5353), .Z(n5350) );
  XNOR U6575 ( .A(x[1222]), .B(n5351), .Z(n5353) );
  XOR U6576 ( .A(n5354), .B(n5355), .Z(n5351) );
  AND U6577 ( .A(n5356), .B(n5357), .Z(n5354) );
  XNOR U6578 ( .A(x[1221]), .B(n5355), .Z(n5357) );
  XOR U6579 ( .A(n5358), .B(n5359), .Z(n5355) );
  AND U6580 ( .A(n5360), .B(n5361), .Z(n5358) );
  XNOR U6581 ( .A(x[1220]), .B(n5359), .Z(n5361) );
  XOR U6582 ( .A(n5362), .B(n5363), .Z(n5359) );
  AND U6583 ( .A(n5364), .B(n5365), .Z(n5362) );
  XNOR U6584 ( .A(x[1219]), .B(n5363), .Z(n5365) );
  XOR U6585 ( .A(n5366), .B(n5367), .Z(n5363) );
  AND U6586 ( .A(n5368), .B(n5369), .Z(n5366) );
  XNOR U6587 ( .A(x[1218]), .B(n5367), .Z(n5369) );
  XOR U6588 ( .A(n5370), .B(n5371), .Z(n5367) );
  AND U6589 ( .A(n5372), .B(n5373), .Z(n5370) );
  XNOR U6590 ( .A(x[1217]), .B(n5371), .Z(n5373) );
  XOR U6591 ( .A(n5374), .B(n5375), .Z(n5371) );
  AND U6592 ( .A(n5376), .B(n5377), .Z(n5374) );
  XNOR U6593 ( .A(x[1216]), .B(n5375), .Z(n5377) );
  XOR U6594 ( .A(n5378), .B(n5379), .Z(n5375) );
  AND U6595 ( .A(n5380), .B(n5381), .Z(n5378) );
  XNOR U6596 ( .A(x[1215]), .B(n5379), .Z(n5381) );
  XOR U6597 ( .A(n5382), .B(n5383), .Z(n5379) );
  AND U6598 ( .A(n5384), .B(n5385), .Z(n5382) );
  XNOR U6599 ( .A(x[1214]), .B(n5383), .Z(n5385) );
  XOR U6600 ( .A(n5386), .B(n5387), .Z(n5383) );
  AND U6601 ( .A(n5388), .B(n5389), .Z(n5386) );
  XNOR U6602 ( .A(x[1213]), .B(n5387), .Z(n5389) );
  XOR U6603 ( .A(n5390), .B(n5391), .Z(n5387) );
  AND U6604 ( .A(n5392), .B(n5393), .Z(n5390) );
  XNOR U6605 ( .A(x[1212]), .B(n5391), .Z(n5393) );
  XOR U6606 ( .A(n5394), .B(n5395), .Z(n5391) );
  AND U6607 ( .A(n5396), .B(n5397), .Z(n5394) );
  XNOR U6608 ( .A(x[1211]), .B(n5395), .Z(n5397) );
  XOR U6609 ( .A(n5398), .B(n5399), .Z(n5395) );
  AND U6610 ( .A(n5400), .B(n5401), .Z(n5398) );
  XNOR U6611 ( .A(x[1210]), .B(n5399), .Z(n5401) );
  XOR U6612 ( .A(n5402), .B(n5403), .Z(n5399) );
  AND U6613 ( .A(n5404), .B(n5405), .Z(n5402) );
  XNOR U6614 ( .A(x[1209]), .B(n5403), .Z(n5405) );
  XOR U6615 ( .A(n5406), .B(n5407), .Z(n5403) );
  AND U6616 ( .A(n5408), .B(n5409), .Z(n5406) );
  XNOR U6617 ( .A(x[1208]), .B(n5407), .Z(n5409) );
  XOR U6618 ( .A(n5410), .B(n5411), .Z(n5407) );
  AND U6619 ( .A(n5412), .B(n5413), .Z(n5410) );
  XNOR U6620 ( .A(x[1207]), .B(n5411), .Z(n5413) );
  XOR U6621 ( .A(n5414), .B(n5415), .Z(n5411) );
  AND U6622 ( .A(n5416), .B(n5417), .Z(n5414) );
  XNOR U6623 ( .A(x[1206]), .B(n5415), .Z(n5417) );
  XOR U6624 ( .A(n5418), .B(n5419), .Z(n5415) );
  AND U6625 ( .A(n5420), .B(n5421), .Z(n5418) );
  XNOR U6626 ( .A(x[1205]), .B(n5419), .Z(n5421) );
  XOR U6627 ( .A(n5422), .B(n5423), .Z(n5419) );
  AND U6628 ( .A(n5424), .B(n5425), .Z(n5422) );
  XNOR U6629 ( .A(x[1204]), .B(n5423), .Z(n5425) );
  XOR U6630 ( .A(n5426), .B(n5427), .Z(n5423) );
  AND U6631 ( .A(n5428), .B(n5429), .Z(n5426) );
  XNOR U6632 ( .A(x[1203]), .B(n5427), .Z(n5429) );
  XOR U6633 ( .A(n5430), .B(n5431), .Z(n5427) );
  AND U6634 ( .A(n5432), .B(n5433), .Z(n5430) );
  XNOR U6635 ( .A(x[1202]), .B(n5431), .Z(n5433) );
  XOR U6636 ( .A(n5434), .B(n5435), .Z(n5431) );
  AND U6637 ( .A(n5436), .B(n5437), .Z(n5434) );
  XNOR U6638 ( .A(x[1201]), .B(n5435), .Z(n5437) );
  XOR U6639 ( .A(n5438), .B(n5439), .Z(n5435) );
  AND U6640 ( .A(n5440), .B(n5441), .Z(n5438) );
  XNOR U6641 ( .A(x[1200]), .B(n5439), .Z(n5441) );
  XOR U6642 ( .A(n5442), .B(n5443), .Z(n5439) );
  AND U6643 ( .A(n5444), .B(n5445), .Z(n5442) );
  XNOR U6644 ( .A(x[1199]), .B(n5443), .Z(n5445) );
  XOR U6645 ( .A(n5446), .B(n5447), .Z(n5443) );
  AND U6646 ( .A(n5448), .B(n5449), .Z(n5446) );
  XNOR U6647 ( .A(x[1198]), .B(n5447), .Z(n5449) );
  XOR U6648 ( .A(n5450), .B(n5451), .Z(n5447) );
  AND U6649 ( .A(n5452), .B(n5453), .Z(n5450) );
  XNOR U6650 ( .A(x[1197]), .B(n5451), .Z(n5453) );
  XOR U6651 ( .A(n5454), .B(n5455), .Z(n5451) );
  AND U6652 ( .A(n5456), .B(n5457), .Z(n5454) );
  XNOR U6653 ( .A(x[1196]), .B(n5455), .Z(n5457) );
  XOR U6654 ( .A(n5458), .B(n5459), .Z(n5455) );
  AND U6655 ( .A(n5460), .B(n5461), .Z(n5458) );
  XNOR U6656 ( .A(x[1195]), .B(n5459), .Z(n5461) );
  XOR U6657 ( .A(n5462), .B(n5463), .Z(n5459) );
  AND U6658 ( .A(n5464), .B(n5465), .Z(n5462) );
  XNOR U6659 ( .A(x[1194]), .B(n5463), .Z(n5465) );
  XOR U6660 ( .A(n5466), .B(n5467), .Z(n5463) );
  AND U6661 ( .A(n5468), .B(n5469), .Z(n5466) );
  XNOR U6662 ( .A(x[1193]), .B(n5467), .Z(n5469) );
  XOR U6663 ( .A(n5470), .B(n5471), .Z(n5467) );
  AND U6664 ( .A(n5472), .B(n5473), .Z(n5470) );
  XNOR U6665 ( .A(x[1192]), .B(n5471), .Z(n5473) );
  XOR U6666 ( .A(n5474), .B(n5475), .Z(n5471) );
  AND U6667 ( .A(n5476), .B(n5477), .Z(n5474) );
  XNOR U6668 ( .A(x[1191]), .B(n5475), .Z(n5477) );
  XOR U6669 ( .A(n5478), .B(n5479), .Z(n5475) );
  AND U6670 ( .A(n5480), .B(n5481), .Z(n5478) );
  XNOR U6671 ( .A(x[1190]), .B(n5479), .Z(n5481) );
  XOR U6672 ( .A(n5482), .B(n5483), .Z(n5479) );
  AND U6673 ( .A(n5484), .B(n5485), .Z(n5482) );
  XNOR U6674 ( .A(x[1189]), .B(n5483), .Z(n5485) );
  XOR U6675 ( .A(n5486), .B(n5487), .Z(n5483) );
  AND U6676 ( .A(n5488), .B(n5489), .Z(n5486) );
  XNOR U6677 ( .A(x[1188]), .B(n5487), .Z(n5489) );
  XOR U6678 ( .A(n5490), .B(n5491), .Z(n5487) );
  AND U6679 ( .A(n5492), .B(n5493), .Z(n5490) );
  XNOR U6680 ( .A(x[1187]), .B(n5491), .Z(n5493) );
  XOR U6681 ( .A(n5494), .B(n5495), .Z(n5491) );
  AND U6682 ( .A(n5496), .B(n5497), .Z(n5494) );
  XNOR U6683 ( .A(x[1186]), .B(n5495), .Z(n5497) );
  XOR U6684 ( .A(n5498), .B(n5499), .Z(n5495) );
  AND U6685 ( .A(n5500), .B(n5501), .Z(n5498) );
  XNOR U6686 ( .A(x[1185]), .B(n5499), .Z(n5501) );
  XOR U6687 ( .A(n5502), .B(n5503), .Z(n5499) );
  AND U6688 ( .A(n5504), .B(n5505), .Z(n5502) );
  XNOR U6689 ( .A(x[1184]), .B(n5503), .Z(n5505) );
  XOR U6690 ( .A(n5506), .B(n5507), .Z(n5503) );
  AND U6691 ( .A(n5508), .B(n5509), .Z(n5506) );
  XNOR U6692 ( .A(x[1183]), .B(n5507), .Z(n5509) );
  XOR U6693 ( .A(n5510), .B(n5511), .Z(n5507) );
  AND U6694 ( .A(n5512), .B(n5513), .Z(n5510) );
  XNOR U6695 ( .A(x[1182]), .B(n5511), .Z(n5513) );
  XOR U6696 ( .A(n5514), .B(n5515), .Z(n5511) );
  AND U6697 ( .A(n5516), .B(n5517), .Z(n5514) );
  XNOR U6698 ( .A(x[1181]), .B(n5515), .Z(n5517) );
  XOR U6699 ( .A(n5518), .B(n5519), .Z(n5515) );
  AND U6700 ( .A(n5520), .B(n5521), .Z(n5518) );
  XNOR U6701 ( .A(x[1180]), .B(n5519), .Z(n5521) );
  XOR U6702 ( .A(n5522), .B(n5523), .Z(n5519) );
  AND U6703 ( .A(n5524), .B(n5525), .Z(n5522) );
  XNOR U6704 ( .A(x[1179]), .B(n5523), .Z(n5525) );
  XOR U6705 ( .A(n5526), .B(n5527), .Z(n5523) );
  AND U6706 ( .A(n5528), .B(n5529), .Z(n5526) );
  XNOR U6707 ( .A(x[1178]), .B(n5527), .Z(n5529) );
  XOR U6708 ( .A(n5530), .B(n5531), .Z(n5527) );
  AND U6709 ( .A(n5532), .B(n5533), .Z(n5530) );
  XNOR U6710 ( .A(x[1177]), .B(n5531), .Z(n5533) );
  XOR U6711 ( .A(n5534), .B(n5535), .Z(n5531) );
  AND U6712 ( .A(n5536), .B(n5537), .Z(n5534) );
  XNOR U6713 ( .A(x[1176]), .B(n5535), .Z(n5537) );
  XOR U6714 ( .A(n5538), .B(n5539), .Z(n5535) );
  AND U6715 ( .A(n5540), .B(n5541), .Z(n5538) );
  XNOR U6716 ( .A(x[1175]), .B(n5539), .Z(n5541) );
  XOR U6717 ( .A(n5542), .B(n5543), .Z(n5539) );
  AND U6718 ( .A(n5544), .B(n5545), .Z(n5542) );
  XNOR U6719 ( .A(x[1174]), .B(n5543), .Z(n5545) );
  XOR U6720 ( .A(n5546), .B(n5547), .Z(n5543) );
  AND U6721 ( .A(n5548), .B(n5549), .Z(n5546) );
  XNOR U6722 ( .A(x[1173]), .B(n5547), .Z(n5549) );
  XOR U6723 ( .A(n5550), .B(n5551), .Z(n5547) );
  AND U6724 ( .A(n5552), .B(n5553), .Z(n5550) );
  XNOR U6725 ( .A(x[1172]), .B(n5551), .Z(n5553) );
  XOR U6726 ( .A(n5554), .B(n5555), .Z(n5551) );
  AND U6727 ( .A(n5556), .B(n5557), .Z(n5554) );
  XNOR U6728 ( .A(x[1171]), .B(n5555), .Z(n5557) );
  XOR U6729 ( .A(n5558), .B(n5559), .Z(n5555) );
  AND U6730 ( .A(n5560), .B(n5561), .Z(n5558) );
  XNOR U6731 ( .A(x[1170]), .B(n5559), .Z(n5561) );
  XOR U6732 ( .A(n5562), .B(n5563), .Z(n5559) );
  AND U6733 ( .A(n5564), .B(n5565), .Z(n5562) );
  XNOR U6734 ( .A(x[1169]), .B(n5563), .Z(n5565) );
  XOR U6735 ( .A(n5566), .B(n5567), .Z(n5563) );
  AND U6736 ( .A(n5568), .B(n5569), .Z(n5566) );
  XNOR U6737 ( .A(x[1168]), .B(n5567), .Z(n5569) );
  XOR U6738 ( .A(n5570), .B(n5571), .Z(n5567) );
  AND U6739 ( .A(n5572), .B(n5573), .Z(n5570) );
  XNOR U6740 ( .A(x[1167]), .B(n5571), .Z(n5573) );
  XOR U6741 ( .A(n5574), .B(n5575), .Z(n5571) );
  AND U6742 ( .A(n5576), .B(n5577), .Z(n5574) );
  XNOR U6743 ( .A(x[1166]), .B(n5575), .Z(n5577) );
  XOR U6744 ( .A(n5578), .B(n5579), .Z(n5575) );
  AND U6745 ( .A(n5580), .B(n5581), .Z(n5578) );
  XNOR U6746 ( .A(x[1165]), .B(n5579), .Z(n5581) );
  XOR U6747 ( .A(n5582), .B(n5583), .Z(n5579) );
  AND U6748 ( .A(n5584), .B(n5585), .Z(n5582) );
  XNOR U6749 ( .A(x[1164]), .B(n5583), .Z(n5585) );
  XOR U6750 ( .A(n5586), .B(n5587), .Z(n5583) );
  AND U6751 ( .A(n5588), .B(n5589), .Z(n5586) );
  XNOR U6752 ( .A(x[1163]), .B(n5587), .Z(n5589) );
  XOR U6753 ( .A(n5590), .B(n5591), .Z(n5587) );
  AND U6754 ( .A(n5592), .B(n5593), .Z(n5590) );
  XNOR U6755 ( .A(x[1162]), .B(n5591), .Z(n5593) );
  XOR U6756 ( .A(n5594), .B(n5595), .Z(n5591) );
  AND U6757 ( .A(n5596), .B(n5597), .Z(n5594) );
  XNOR U6758 ( .A(x[1161]), .B(n5595), .Z(n5597) );
  XOR U6759 ( .A(n5598), .B(n5599), .Z(n5595) );
  AND U6760 ( .A(n5600), .B(n5601), .Z(n5598) );
  XNOR U6761 ( .A(x[1160]), .B(n5599), .Z(n5601) );
  XOR U6762 ( .A(n5602), .B(n5603), .Z(n5599) );
  AND U6763 ( .A(n5604), .B(n5605), .Z(n5602) );
  XNOR U6764 ( .A(x[1159]), .B(n5603), .Z(n5605) );
  XOR U6765 ( .A(n5606), .B(n5607), .Z(n5603) );
  AND U6766 ( .A(n5608), .B(n5609), .Z(n5606) );
  XNOR U6767 ( .A(x[1158]), .B(n5607), .Z(n5609) );
  XOR U6768 ( .A(n5610), .B(n5611), .Z(n5607) );
  AND U6769 ( .A(n5612), .B(n5613), .Z(n5610) );
  XNOR U6770 ( .A(x[1157]), .B(n5611), .Z(n5613) );
  XOR U6771 ( .A(n5614), .B(n5615), .Z(n5611) );
  AND U6772 ( .A(n5616), .B(n5617), .Z(n5614) );
  XNOR U6773 ( .A(x[1156]), .B(n5615), .Z(n5617) );
  XOR U6774 ( .A(n5618), .B(n5619), .Z(n5615) );
  AND U6775 ( .A(n5620), .B(n5621), .Z(n5618) );
  XNOR U6776 ( .A(x[1155]), .B(n5619), .Z(n5621) );
  XOR U6777 ( .A(n5622), .B(n5623), .Z(n5619) );
  AND U6778 ( .A(n5624), .B(n5625), .Z(n5622) );
  XNOR U6779 ( .A(x[1154]), .B(n5623), .Z(n5625) );
  XOR U6780 ( .A(n5626), .B(n5627), .Z(n5623) );
  AND U6781 ( .A(n5628), .B(n5629), .Z(n5626) );
  XNOR U6782 ( .A(x[1153]), .B(n5627), .Z(n5629) );
  XOR U6783 ( .A(n5630), .B(n5631), .Z(n5627) );
  AND U6784 ( .A(n5632), .B(n5633), .Z(n5630) );
  XNOR U6785 ( .A(x[1152]), .B(n5631), .Z(n5633) );
  XOR U6786 ( .A(n5634), .B(n5635), .Z(n5631) );
  AND U6787 ( .A(n5636), .B(n5637), .Z(n5634) );
  XNOR U6788 ( .A(x[1151]), .B(n5635), .Z(n5637) );
  XOR U6789 ( .A(n5638), .B(n5639), .Z(n5635) );
  AND U6790 ( .A(n5640), .B(n5641), .Z(n5638) );
  XNOR U6791 ( .A(x[1150]), .B(n5639), .Z(n5641) );
  XOR U6792 ( .A(n5642), .B(n5643), .Z(n5639) );
  AND U6793 ( .A(n5644), .B(n5645), .Z(n5642) );
  XNOR U6794 ( .A(x[1149]), .B(n5643), .Z(n5645) );
  XOR U6795 ( .A(n5646), .B(n5647), .Z(n5643) );
  AND U6796 ( .A(n5648), .B(n5649), .Z(n5646) );
  XNOR U6797 ( .A(x[1148]), .B(n5647), .Z(n5649) );
  XOR U6798 ( .A(n5650), .B(n5651), .Z(n5647) );
  AND U6799 ( .A(n5652), .B(n5653), .Z(n5650) );
  XNOR U6800 ( .A(x[1147]), .B(n5651), .Z(n5653) );
  XOR U6801 ( .A(n5654), .B(n5655), .Z(n5651) );
  AND U6802 ( .A(n5656), .B(n5657), .Z(n5654) );
  XNOR U6803 ( .A(x[1146]), .B(n5655), .Z(n5657) );
  XOR U6804 ( .A(n5658), .B(n5659), .Z(n5655) );
  AND U6805 ( .A(n5660), .B(n5661), .Z(n5658) );
  XNOR U6806 ( .A(x[1145]), .B(n5659), .Z(n5661) );
  XOR U6807 ( .A(n5662), .B(n5663), .Z(n5659) );
  AND U6808 ( .A(n5664), .B(n5665), .Z(n5662) );
  XNOR U6809 ( .A(x[1144]), .B(n5663), .Z(n5665) );
  XOR U6810 ( .A(n5666), .B(n5667), .Z(n5663) );
  AND U6811 ( .A(n5668), .B(n5669), .Z(n5666) );
  XNOR U6812 ( .A(x[1143]), .B(n5667), .Z(n5669) );
  XOR U6813 ( .A(n5670), .B(n5671), .Z(n5667) );
  AND U6814 ( .A(n5672), .B(n5673), .Z(n5670) );
  XNOR U6815 ( .A(x[1142]), .B(n5671), .Z(n5673) );
  XOR U6816 ( .A(n5674), .B(n5675), .Z(n5671) );
  AND U6817 ( .A(n5676), .B(n5677), .Z(n5674) );
  XNOR U6818 ( .A(x[1141]), .B(n5675), .Z(n5677) );
  XOR U6819 ( .A(n5678), .B(n5679), .Z(n5675) );
  AND U6820 ( .A(n5680), .B(n5681), .Z(n5678) );
  XNOR U6821 ( .A(x[1140]), .B(n5679), .Z(n5681) );
  XOR U6822 ( .A(n5682), .B(n5683), .Z(n5679) );
  AND U6823 ( .A(n5684), .B(n5685), .Z(n5682) );
  XNOR U6824 ( .A(x[1139]), .B(n5683), .Z(n5685) );
  XOR U6825 ( .A(n5686), .B(n5687), .Z(n5683) );
  AND U6826 ( .A(n5688), .B(n5689), .Z(n5686) );
  XNOR U6827 ( .A(x[1138]), .B(n5687), .Z(n5689) );
  XOR U6828 ( .A(n5690), .B(n5691), .Z(n5687) );
  AND U6829 ( .A(n5692), .B(n5693), .Z(n5690) );
  XNOR U6830 ( .A(x[1137]), .B(n5691), .Z(n5693) );
  XOR U6831 ( .A(n5694), .B(n5695), .Z(n5691) );
  AND U6832 ( .A(n5696), .B(n5697), .Z(n5694) );
  XNOR U6833 ( .A(x[1136]), .B(n5695), .Z(n5697) );
  XOR U6834 ( .A(n5698), .B(n5699), .Z(n5695) );
  AND U6835 ( .A(n5700), .B(n5701), .Z(n5698) );
  XNOR U6836 ( .A(x[1135]), .B(n5699), .Z(n5701) );
  XOR U6837 ( .A(n5702), .B(n5703), .Z(n5699) );
  AND U6838 ( .A(n5704), .B(n5705), .Z(n5702) );
  XNOR U6839 ( .A(x[1134]), .B(n5703), .Z(n5705) );
  XOR U6840 ( .A(n5706), .B(n5707), .Z(n5703) );
  AND U6841 ( .A(n5708), .B(n5709), .Z(n5706) );
  XNOR U6842 ( .A(x[1133]), .B(n5707), .Z(n5709) );
  XOR U6843 ( .A(n5710), .B(n5711), .Z(n5707) );
  AND U6844 ( .A(n5712), .B(n5713), .Z(n5710) );
  XNOR U6845 ( .A(x[1132]), .B(n5711), .Z(n5713) );
  XOR U6846 ( .A(n5714), .B(n5715), .Z(n5711) );
  AND U6847 ( .A(n5716), .B(n5717), .Z(n5714) );
  XNOR U6848 ( .A(x[1131]), .B(n5715), .Z(n5717) );
  XOR U6849 ( .A(n5718), .B(n5719), .Z(n5715) );
  AND U6850 ( .A(n5720), .B(n5721), .Z(n5718) );
  XNOR U6851 ( .A(x[1130]), .B(n5719), .Z(n5721) );
  XOR U6852 ( .A(n5722), .B(n5723), .Z(n5719) );
  AND U6853 ( .A(n5724), .B(n5725), .Z(n5722) );
  XNOR U6854 ( .A(x[1129]), .B(n5723), .Z(n5725) );
  XOR U6855 ( .A(n5726), .B(n5727), .Z(n5723) );
  AND U6856 ( .A(n5728), .B(n5729), .Z(n5726) );
  XNOR U6857 ( .A(x[1128]), .B(n5727), .Z(n5729) );
  XOR U6858 ( .A(n5730), .B(n5731), .Z(n5727) );
  AND U6859 ( .A(n5732), .B(n5733), .Z(n5730) );
  XNOR U6860 ( .A(x[1127]), .B(n5731), .Z(n5733) );
  XOR U6861 ( .A(n5734), .B(n5735), .Z(n5731) );
  AND U6862 ( .A(n5736), .B(n5737), .Z(n5734) );
  XNOR U6863 ( .A(x[1126]), .B(n5735), .Z(n5737) );
  XOR U6864 ( .A(n5738), .B(n5739), .Z(n5735) );
  AND U6865 ( .A(n5740), .B(n5741), .Z(n5738) );
  XNOR U6866 ( .A(x[1125]), .B(n5739), .Z(n5741) );
  XOR U6867 ( .A(n5742), .B(n5743), .Z(n5739) );
  AND U6868 ( .A(n5744), .B(n5745), .Z(n5742) );
  XNOR U6869 ( .A(x[1124]), .B(n5743), .Z(n5745) );
  XOR U6870 ( .A(n5746), .B(n5747), .Z(n5743) );
  AND U6871 ( .A(n5748), .B(n5749), .Z(n5746) );
  XNOR U6872 ( .A(x[1123]), .B(n5747), .Z(n5749) );
  XOR U6873 ( .A(n5750), .B(n5751), .Z(n5747) );
  AND U6874 ( .A(n5752), .B(n5753), .Z(n5750) );
  XNOR U6875 ( .A(x[1122]), .B(n5751), .Z(n5753) );
  XOR U6876 ( .A(n5754), .B(n5755), .Z(n5751) );
  AND U6877 ( .A(n5756), .B(n5757), .Z(n5754) );
  XNOR U6878 ( .A(x[1121]), .B(n5755), .Z(n5757) );
  XOR U6879 ( .A(n5758), .B(n5759), .Z(n5755) );
  AND U6880 ( .A(n5760), .B(n5761), .Z(n5758) );
  XNOR U6881 ( .A(x[1120]), .B(n5759), .Z(n5761) );
  XOR U6882 ( .A(n5762), .B(n5763), .Z(n5759) );
  AND U6883 ( .A(n5764), .B(n5765), .Z(n5762) );
  XNOR U6884 ( .A(x[1119]), .B(n5763), .Z(n5765) );
  XOR U6885 ( .A(n5766), .B(n5767), .Z(n5763) );
  AND U6886 ( .A(n5768), .B(n5769), .Z(n5766) );
  XNOR U6887 ( .A(x[1118]), .B(n5767), .Z(n5769) );
  XOR U6888 ( .A(n5770), .B(n5771), .Z(n5767) );
  AND U6889 ( .A(n5772), .B(n5773), .Z(n5770) );
  XNOR U6890 ( .A(x[1117]), .B(n5771), .Z(n5773) );
  XOR U6891 ( .A(n5774), .B(n5775), .Z(n5771) );
  AND U6892 ( .A(n5776), .B(n5777), .Z(n5774) );
  XNOR U6893 ( .A(x[1116]), .B(n5775), .Z(n5777) );
  XOR U6894 ( .A(n5778), .B(n5779), .Z(n5775) );
  AND U6895 ( .A(n5780), .B(n5781), .Z(n5778) );
  XNOR U6896 ( .A(x[1115]), .B(n5779), .Z(n5781) );
  XOR U6897 ( .A(n5782), .B(n5783), .Z(n5779) );
  AND U6898 ( .A(n5784), .B(n5785), .Z(n5782) );
  XNOR U6899 ( .A(x[1114]), .B(n5783), .Z(n5785) );
  XOR U6900 ( .A(n5786), .B(n5787), .Z(n5783) );
  AND U6901 ( .A(n5788), .B(n5789), .Z(n5786) );
  XNOR U6902 ( .A(x[1113]), .B(n5787), .Z(n5789) );
  XOR U6903 ( .A(n5790), .B(n5791), .Z(n5787) );
  AND U6904 ( .A(n5792), .B(n5793), .Z(n5790) );
  XNOR U6905 ( .A(x[1112]), .B(n5791), .Z(n5793) );
  XOR U6906 ( .A(n5794), .B(n5795), .Z(n5791) );
  AND U6907 ( .A(n5796), .B(n5797), .Z(n5794) );
  XNOR U6908 ( .A(x[1111]), .B(n5795), .Z(n5797) );
  XOR U6909 ( .A(n5798), .B(n5799), .Z(n5795) );
  AND U6910 ( .A(n5800), .B(n5801), .Z(n5798) );
  XNOR U6911 ( .A(x[1110]), .B(n5799), .Z(n5801) );
  XOR U6912 ( .A(n5802), .B(n5803), .Z(n5799) );
  AND U6913 ( .A(n5804), .B(n5805), .Z(n5802) );
  XNOR U6914 ( .A(x[1109]), .B(n5803), .Z(n5805) );
  XOR U6915 ( .A(n5806), .B(n5807), .Z(n5803) );
  AND U6916 ( .A(n5808), .B(n5809), .Z(n5806) );
  XNOR U6917 ( .A(x[1108]), .B(n5807), .Z(n5809) );
  XOR U6918 ( .A(n5810), .B(n5811), .Z(n5807) );
  AND U6919 ( .A(n5812), .B(n5813), .Z(n5810) );
  XNOR U6920 ( .A(x[1107]), .B(n5811), .Z(n5813) );
  XOR U6921 ( .A(n5814), .B(n5815), .Z(n5811) );
  AND U6922 ( .A(n5816), .B(n5817), .Z(n5814) );
  XNOR U6923 ( .A(x[1106]), .B(n5815), .Z(n5817) );
  XOR U6924 ( .A(n5818), .B(n5819), .Z(n5815) );
  AND U6925 ( .A(n5820), .B(n5821), .Z(n5818) );
  XNOR U6926 ( .A(x[1105]), .B(n5819), .Z(n5821) );
  XOR U6927 ( .A(n5822), .B(n5823), .Z(n5819) );
  AND U6928 ( .A(n5824), .B(n5825), .Z(n5822) );
  XNOR U6929 ( .A(x[1104]), .B(n5823), .Z(n5825) );
  XOR U6930 ( .A(n5826), .B(n5827), .Z(n5823) );
  AND U6931 ( .A(n5828), .B(n5829), .Z(n5826) );
  XNOR U6932 ( .A(x[1103]), .B(n5827), .Z(n5829) );
  XOR U6933 ( .A(n5830), .B(n5831), .Z(n5827) );
  AND U6934 ( .A(n5832), .B(n5833), .Z(n5830) );
  XNOR U6935 ( .A(x[1102]), .B(n5831), .Z(n5833) );
  XOR U6936 ( .A(n5834), .B(n5835), .Z(n5831) );
  AND U6937 ( .A(n5836), .B(n5837), .Z(n5834) );
  XNOR U6938 ( .A(x[1101]), .B(n5835), .Z(n5837) );
  XOR U6939 ( .A(n5838), .B(n5839), .Z(n5835) );
  AND U6940 ( .A(n5840), .B(n5841), .Z(n5838) );
  XNOR U6941 ( .A(x[1100]), .B(n5839), .Z(n5841) );
  XOR U6942 ( .A(n5842), .B(n5843), .Z(n5839) );
  AND U6943 ( .A(n5844), .B(n5845), .Z(n5842) );
  XNOR U6944 ( .A(x[1099]), .B(n5843), .Z(n5845) );
  XOR U6945 ( .A(n5846), .B(n5847), .Z(n5843) );
  AND U6946 ( .A(n5848), .B(n5849), .Z(n5846) );
  XNOR U6947 ( .A(x[1098]), .B(n5847), .Z(n5849) );
  XOR U6948 ( .A(n5850), .B(n5851), .Z(n5847) );
  AND U6949 ( .A(n5852), .B(n5853), .Z(n5850) );
  XNOR U6950 ( .A(x[1097]), .B(n5851), .Z(n5853) );
  XOR U6951 ( .A(n5854), .B(n5855), .Z(n5851) );
  AND U6952 ( .A(n5856), .B(n5857), .Z(n5854) );
  XNOR U6953 ( .A(x[1096]), .B(n5855), .Z(n5857) );
  XOR U6954 ( .A(n5858), .B(n5859), .Z(n5855) );
  AND U6955 ( .A(n5860), .B(n5861), .Z(n5858) );
  XNOR U6956 ( .A(x[1095]), .B(n5859), .Z(n5861) );
  XOR U6957 ( .A(n5862), .B(n5863), .Z(n5859) );
  AND U6958 ( .A(n5864), .B(n5865), .Z(n5862) );
  XNOR U6959 ( .A(x[1094]), .B(n5863), .Z(n5865) );
  XOR U6960 ( .A(n5866), .B(n5867), .Z(n5863) );
  AND U6961 ( .A(n5868), .B(n5869), .Z(n5866) );
  XNOR U6962 ( .A(x[1093]), .B(n5867), .Z(n5869) );
  XOR U6963 ( .A(n5870), .B(n5871), .Z(n5867) );
  AND U6964 ( .A(n5872), .B(n5873), .Z(n5870) );
  XNOR U6965 ( .A(x[1092]), .B(n5871), .Z(n5873) );
  XOR U6966 ( .A(n5874), .B(n5875), .Z(n5871) );
  AND U6967 ( .A(n5876), .B(n5877), .Z(n5874) );
  XNOR U6968 ( .A(x[1091]), .B(n5875), .Z(n5877) );
  XOR U6969 ( .A(n5878), .B(n5879), .Z(n5875) );
  AND U6970 ( .A(n5880), .B(n5881), .Z(n5878) );
  XNOR U6971 ( .A(x[1090]), .B(n5879), .Z(n5881) );
  XOR U6972 ( .A(n5882), .B(n5883), .Z(n5879) );
  AND U6973 ( .A(n5884), .B(n5885), .Z(n5882) );
  XNOR U6974 ( .A(x[1089]), .B(n5883), .Z(n5885) );
  XOR U6975 ( .A(n5886), .B(n5887), .Z(n5883) );
  AND U6976 ( .A(n5888), .B(n5889), .Z(n5886) );
  XNOR U6977 ( .A(x[1088]), .B(n5887), .Z(n5889) );
  XOR U6978 ( .A(n5890), .B(n5891), .Z(n5887) );
  AND U6979 ( .A(n5892), .B(n5893), .Z(n5890) );
  XNOR U6980 ( .A(x[1087]), .B(n5891), .Z(n5893) );
  XOR U6981 ( .A(n5894), .B(n5895), .Z(n5891) );
  AND U6982 ( .A(n5896), .B(n5897), .Z(n5894) );
  XNOR U6983 ( .A(x[1086]), .B(n5895), .Z(n5897) );
  XOR U6984 ( .A(n5898), .B(n5899), .Z(n5895) );
  AND U6985 ( .A(n5900), .B(n5901), .Z(n5898) );
  XNOR U6986 ( .A(x[1085]), .B(n5899), .Z(n5901) );
  XOR U6987 ( .A(n5902), .B(n5903), .Z(n5899) );
  AND U6988 ( .A(n5904), .B(n5905), .Z(n5902) );
  XNOR U6989 ( .A(x[1084]), .B(n5903), .Z(n5905) );
  XOR U6990 ( .A(n5906), .B(n5907), .Z(n5903) );
  AND U6991 ( .A(n5908), .B(n5909), .Z(n5906) );
  XNOR U6992 ( .A(x[1083]), .B(n5907), .Z(n5909) );
  XOR U6993 ( .A(n5910), .B(n5911), .Z(n5907) );
  AND U6994 ( .A(n5912), .B(n5913), .Z(n5910) );
  XNOR U6995 ( .A(x[1082]), .B(n5911), .Z(n5913) );
  XOR U6996 ( .A(n5914), .B(n5915), .Z(n5911) );
  AND U6997 ( .A(n5916), .B(n5917), .Z(n5914) );
  XNOR U6998 ( .A(x[1081]), .B(n5915), .Z(n5917) );
  XOR U6999 ( .A(n5918), .B(n5919), .Z(n5915) );
  AND U7000 ( .A(n5920), .B(n5921), .Z(n5918) );
  XNOR U7001 ( .A(x[1080]), .B(n5919), .Z(n5921) );
  XOR U7002 ( .A(n5922), .B(n5923), .Z(n5919) );
  AND U7003 ( .A(n5924), .B(n5925), .Z(n5922) );
  XNOR U7004 ( .A(x[1079]), .B(n5923), .Z(n5925) );
  XOR U7005 ( .A(n5926), .B(n5927), .Z(n5923) );
  AND U7006 ( .A(n5928), .B(n5929), .Z(n5926) );
  XNOR U7007 ( .A(x[1078]), .B(n5927), .Z(n5929) );
  XOR U7008 ( .A(n5930), .B(n5931), .Z(n5927) );
  AND U7009 ( .A(n5932), .B(n5933), .Z(n5930) );
  XNOR U7010 ( .A(x[1077]), .B(n5931), .Z(n5933) );
  XOR U7011 ( .A(n5934), .B(n5935), .Z(n5931) );
  AND U7012 ( .A(n5936), .B(n5937), .Z(n5934) );
  XNOR U7013 ( .A(x[1076]), .B(n5935), .Z(n5937) );
  XOR U7014 ( .A(n5938), .B(n5939), .Z(n5935) );
  AND U7015 ( .A(n5940), .B(n5941), .Z(n5938) );
  XNOR U7016 ( .A(x[1075]), .B(n5939), .Z(n5941) );
  XOR U7017 ( .A(n5942), .B(n5943), .Z(n5939) );
  AND U7018 ( .A(n5944), .B(n5945), .Z(n5942) );
  XNOR U7019 ( .A(x[1074]), .B(n5943), .Z(n5945) );
  XOR U7020 ( .A(n5946), .B(n5947), .Z(n5943) );
  AND U7021 ( .A(n5948), .B(n5949), .Z(n5946) );
  XNOR U7022 ( .A(x[1073]), .B(n5947), .Z(n5949) );
  XOR U7023 ( .A(n5950), .B(n5951), .Z(n5947) );
  AND U7024 ( .A(n5952), .B(n5953), .Z(n5950) );
  XNOR U7025 ( .A(x[1072]), .B(n5951), .Z(n5953) );
  XOR U7026 ( .A(n5954), .B(n5955), .Z(n5951) );
  AND U7027 ( .A(n5956), .B(n5957), .Z(n5954) );
  XNOR U7028 ( .A(x[1071]), .B(n5955), .Z(n5957) );
  XOR U7029 ( .A(n5958), .B(n5959), .Z(n5955) );
  AND U7030 ( .A(n5960), .B(n5961), .Z(n5958) );
  XNOR U7031 ( .A(x[1070]), .B(n5959), .Z(n5961) );
  XOR U7032 ( .A(n5962), .B(n5963), .Z(n5959) );
  AND U7033 ( .A(n5964), .B(n5965), .Z(n5962) );
  XNOR U7034 ( .A(x[1069]), .B(n5963), .Z(n5965) );
  XOR U7035 ( .A(n5966), .B(n5967), .Z(n5963) );
  AND U7036 ( .A(n5968), .B(n5969), .Z(n5966) );
  XNOR U7037 ( .A(x[1068]), .B(n5967), .Z(n5969) );
  XOR U7038 ( .A(n5970), .B(n5971), .Z(n5967) );
  AND U7039 ( .A(n5972), .B(n5973), .Z(n5970) );
  XNOR U7040 ( .A(x[1067]), .B(n5971), .Z(n5973) );
  XOR U7041 ( .A(n5974), .B(n5975), .Z(n5971) );
  AND U7042 ( .A(n5976), .B(n5977), .Z(n5974) );
  XNOR U7043 ( .A(x[1066]), .B(n5975), .Z(n5977) );
  XOR U7044 ( .A(n5978), .B(n5979), .Z(n5975) );
  AND U7045 ( .A(n5980), .B(n5981), .Z(n5978) );
  XNOR U7046 ( .A(x[1065]), .B(n5979), .Z(n5981) );
  XOR U7047 ( .A(n5982), .B(n5983), .Z(n5979) );
  AND U7048 ( .A(n5984), .B(n5985), .Z(n5982) );
  XNOR U7049 ( .A(x[1064]), .B(n5983), .Z(n5985) );
  XOR U7050 ( .A(n5986), .B(n5987), .Z(n5983) );
  AND U7051 ( .A(n5988), .B(n5989), .Z(n5986) );
  XNOR U7052 ( .A(x[1063]), .B(n5987), .Z(n5989) );
  XOR U7053 ( .A(n5990), .B(n5991), .Z(n5987) );
  AND U7054 ( .A(n5992), .B(n5993), .Z(n5990) );
  XNOR U7055 ( .A(x[1062]), .B(n5991), .Z(n5993) );
  XOR U7056 ( .A(n5994), .B(n5995), .Z(n5991) );
  AND U7057 ( .A(n5996), .B(n5997), .Z(n5994) );
  XNOR U7058 ( .A(x[1061]), .B(n5995), .Z(n5997) );
  XOR U7059 ( .A(n5998), .B(n5999), .Z(n5995) );
  AND U7060 ( .A(n6000), .B(n6001), .Z(n5998) );
  XNOR U7061 ( .A(x[1060]), .B(n5999), .Z(n6001) );
  XOR U7062 ( .A(n6002), .B(n6003), .Z(n5999) );
  AND U7063 ( .A(n6004), .B(n6005), .Z(n6002) );
  XNOR U7064 ( .A(x[1059]), .B(n6003), .Z(n6005) );
  XOR U7065 ( .A(n6006), .B(n6007), .Z(n6003) );
  AND U7066 ( .A(n6008), .B(n6009), .Z(n6006) );
  XNOR U7067 ( .A(x[1058]), .B(n6007), .Z(n6009) );
  XOR U7068 ( .A(n6010), .B(n6011), .Z(n6007) );
  AND U7069 ( .A(n6012), .B(n6013), .Z(n6010) );
  XNOR U7070 ( .A(x[1057]), .B(n6011), .Z(n6013) );
  XOR U7071 ( .A(n6014), .B(n6015), .Z(n6011) );
  AND U7072 ( .A(n6016), .B(n6017), .Z(n6014) );
  XNOR U7073 ( .A(x[1056]), .B(n6015), .Z(n6017) );
  XOR U7074 ( .A(n6018), .B(n6019), .Z(n6015) );
  AND U7075 ( .A(n6020), .B(n6021), .Z(n6018) );
  XNOR U7076 ( .A(x[1055]), .B(n6019), .Z(n6021) );
  XOR U7077 ( .A(n6022), .B(n6023), .Z(n6019) );
  AND U7078 ( .A(n6024), .B(n6025), .Z(n6022) );
  XNOR U7079 ( .A(x[1054]), .B(n6023), .Z(n6025) );
  XOR U7080 ( .A(n6026), .B(n6027), .Z(n6023) );
  AND U7081 ( .A(n6028), .B(n6029), .Z(n6026) );
  XNOR U7082 ( .A(x[1053]), .B(n6027), .Z(n6029) );
  XOR U7083 ( .A(n6030), .B(n6031), .Z(n6027) );
  AND U7084 ( .A(n6032), .B(n6033), .Z(n6030) );
  XNOR U7085 ( .A(x[1052]), .B(n6031), .Z(n6033) );
  XOR U7086 ( .A(n6034), .B(n6035), .Z(n6031) );
  AND U7087 ( .A(n6036), .B(n6037), .Z(n6034) );
  XNOR U7088 ( .A(x[1051]), .B(n6035), .Z(n6037) );
  XOR U7089 ( .A(n6038), .B(n6039), .Z(n6035) );
  AND U7090 ( .A(n6040), .B(n6041), .Z(n6038) );
  XNOR U7091 ( .A(x[1050]), .B(n6039), .Z(n6041) );
  XOR U7092 ( .A(n6042), .B(n6043), .Z(n6039) );
  AND U7093 ( .A(n6044), .B(n6045), .Z(n6042) );
  XNOR U7094 ( .A(x[1049]), .B(n6043), .Z(n6045) );
  XOR U7095 ( .A(n6046), .B(n6047), .Z(n6043) );
  AND U7096 ( .A(n6048), .B(n6049), .Z(n6046) );
  XNOR U7097 ( .A(x[1048]), .B(n6047), .Z(n6049) );
  XOR U7098 ( .A(n6050), .B(n6051), .Z(n6047) );
  AND U7099 ( .A(n6052), .B(n6053), .Z(n6050) );
  XNOR U7100 ( .A(x[1047]), .B(n6051), .Z(n6053) );
  XOR U7101 ( .A(n6054), .B(n6055), .Z(n6051) );
  AND U7102 ( .A(n6056), .B(n6057), .Z(n6054) );
  XNOR U7103 ( .A(x[1046]), .B(n6055), .Z(n6057) );
  XOR U7104 ( .A(n6058), .B(n6059), .Z(n6055) );
  AND U7105 ( .A(n6060), .B(n6061), .Z(n6058) );
  XNOR U7106 ( .A(x[1045]), .B(n6059), .Z(n6061) );
  XOR U7107 ( .A(n6062), .B(n6063), .Z(n6059) );
  AND U7108 ( .A(n6064), .B(n6065), .Z(n6062) );
  XNOR U7109 ( .A(x[1044]), .B(n6063), .Z(n6065) );
  XOR U7110 ( .A(n6066), .B(n6067), .Z(n6063) );
  AND U7111 ( .A(n6068), .B(n6069), .Z(n6066) );
  XNOR U7112 ( .A(x[1043]), .B(n6067), .Z(n6069) );
  XOR U7113 ( .A(n6070), .B(n6071), .Z(n6067) );
  AND U7114 ( .A(n6072), .B(n6073), .Z(n6070) );
  XNOR U7115 ( .A(x[1042]), .B(n6071), .Z(n6073) );
  XOR U7116 ( .A(n6074), .B(n6075), .Z(n6071) );
  AND U7117 ( .A(n6076), .B(n6077), .Z(n6074) );
  XNOR U7118 ( .A(x[1041]), .B(n6075), .Z(n6077) );
  XOR U7119 ( .A(n6078), .B(n6079), .Z(n6075) );
  AND U7120 ( .A(n6080), .B(n6081), .Z(n6078) );
  XNOR U7121 ( .A(x[1040]), .B(n6079), .Z(n6081) );
  XOR U7122 ( .A(n6082), .B(n6083), .Z(n6079) );
  AND U7123 ( .A(n6084), .B(n6085), .Z(n6082) );
  XNOR U7124 ( .A(x[1039]), .B(n6083), .Z(n6085) );
  XOR U7125 ( .A(n6086), .B(n6087), .Z(n6083) );
  AND U7126 ( .A(n6088), .B(n6089), .Z(n6086) );
  XNOR U7127 ( .A(x[1038]), .B(n6087), .Z(n6089) );
  XOR U7128 ( .A(n6090), .B(n6091), .Z(n6087) );
  AND U7129 ( .A(n6092), .B(n6093), .Z(n6090) );
  XNOR U7130 ( .A(x[1037]), .B(n6091), .Z(n6093) );
  XOR U7131 ( .A(n6094), .B(n6095), .Z(n6091) );
  AND U7132 ( .A(n6096), .B(n6097), .Z(n6094) );
  XNOR U7133 ( .A(x[1036]), .B(n6095), .Z(n6097) );
  XOR U7134 ( .A(n6098), .B(n6099), .Z(n6095) );
  AND U7135 ( .A(n6100), .B(n6101), .Z(n6098) );
  XNOR U7136 ( .A(x[1035]), .B(n6099), .Z(n6101) );
  XOR U7137 ( .A(n6102), .B(n6103), .Z(n6099) );
  AND U7138 ( .A(n6104), .B(n6105), .Z(n6102) );
  XNOR U7139 ( .A(x[1034]), .B(n6103), .Z(n6105) );
  XOR U7140 ( .A(n6106), .B(n6107), .Z(n6103) );
  AND U7141 ( .A(n6108), .B(n6109), .Z(n6106) );
  XNOR U7142 ( .A(x[1033]), .B(n6107), .Z(n6109) );
  XOR U7143 ( .A(n6110), .B(n6111), .Z(n6107) );
  AND U7144 ( .A(n6112), .B(n6113), .Z(n6110) );
  XNOR U7145 ( .A(x[1032]), .B(n6111), .Z(n6113) );
  XOR U7146 ( .A(n6114), .B(n6115), .Z(n6111) );
  AND U7147 ( .A(n6116), .B(n6117), .Z(n6114) );
  XNOR U7148 ( .A(x[1031]), .B(n6115), .Z(n6117) );
  XOR U7149 ( .A(n6118), .B(n6119), .Z(n6115) );
  AND U7150 ( .A(n6120), .B(n6121), .Z(n6118) );
  XNOR U7151 ( .A(x[1030]), .B(n6119), .Z(n6121) );
  XOR U7152 ( .A(n6122), .B(n6123), .Z(n6119) );
  AND U7153 ( .A(n6124), .B(n6125), .Z(n6122) );
  XNOR U7154 ( .A(x[1029]), .B(n6123), .Z(n6125) );
  XOR U7155 ( .A(n6126), .B(n6127), .Z(n6123) );
  AND U7156 ( .A(n6128), .B(n6129), .Z(n6126) );
  XNOR U7157 ( .A(x[1028]), .B(n6127), .Z(n6129) );
  XOR U7158 ( .A(n6130), .B(n6131), .Z(n6127) );
  AND U7159 ( .A(n6132), .B(n6133), .Z(n6130) );
  XNOR U7160 ( .A(x[1027]), .B(n6131), .Z(n6133) );
  XOR U7161 ( .A(n6134), .B(n6135), .Z(n6131) );
  AND U7162 ( .A(n6136), .B(n6137), .Z(n6134) );
  XNOR U7163 ( .A(x[1026]), .B(n6135), .Z(n6137) );
  XOR U7164 ( .A(n6138), .B(n6139), .Z(n6135) );
  AND U7165 ( .A(n6140), .B(n6141), .Z(n6138) );
  XNOR U7166 ( .A(x[1025]), .B(n6139), .Z(n6141) );
  XOR U7167 ( .A(n6142), .B(n6143), .Z(n6139) );
  AND U7168 ( .A(n6144), .B(n6145), .Z(n6142) );
  XNOR U7169 ( .A(x[1024]), .B(n6143), .Z(n6145) );
  XOR U7170 ( .A(n6146), .B(n6147), .Z(n6143) );
  AND U7171 ( .A(n6148), .B(n6149), .Z(n6146) );
  XNOR U7172 ( .A(x[1023]), .B(n6147), .Z(n6149) );
  XOR U7173 ( .A(n6150), .B(n6151), .Z(n6147) );
  AND U7174 ( .A(n6152), .B(n6153), .Z(n6150) );
  XNOR U7175 ( .A(x[1022]), .B(n6151), .Z(n6153) );
  XOR U7176 ( .A(n6154), .B(n6155), .Z(n6151) );
  AND U7177 ( .A(n6156), .B(n6157), .Z(n6154) );
  XNOR U7178 ( .A(x[1021]), .B(n6155), .Z(n6157) );
  XOR U7179 ( .A(n6158), .B(n6159), .Z(n6155) );
  AND U7180 ( .A(n6160), .B(n6161), .Z(n6158) );
  XNOR U7181 ( .A(x[1020]), .B(n6159), .Z(n6161) );
  XOR U7182 ( .A(n6162), .B(n6163), .Z(n6159) );
  AND U7183 ( .A(n6164), .B(n6165), .Z(n6162) );
  XNOR U7184 ( .A(x[1019]), .B(n6163), .Z(n6165) );
  XOR U7185 ( .A(n6166), .B(n6167), .Z(n6163) );
  AND U7186 ( .A(n6168), .B(n6169), .Z(n6166) );
  XNOR U7187 ( .A(x[1018]), .B(n6167), .Z(n6169) );
  XOR U7188 ( .A(n6170), .B(n6171), .Z(n6167) );
  AND U7189 ( .A(n6172), .B(n6173), .Z(n6170) );
  XNOR U7190 ( .A(x[1017]), .B(n6171), .Z(n6173) );
  XOR U7191 ( .A(n6174), .B(n6175), .Z(n6171) );
  AND U7192 ( .A(n6176), .B(n6177), .Z(n6174) );
  XNOR U7193 ( .A(x[1016]), .B(n6175), .Z(n6177) );
  XOR U7194 ( .A(n6178), .B(n6179), .Z(n6175) );
  AND U7195 ( .A(n6180), .B(n6181), .Z(n6178) );
  XNOR U7196 ( .A(x[1015]), .B(n6179), .Z(n6181) );
  XOR U7197 ( .A(n6182), .B(n6183), .Z(n6179) );
  AND U7198 ( .A(n6184), .B(n6185), .Z(n6182) );
  XNOR U7199 ( .A(x[1014]), .B(n6183), .Z(n6185) );
  XOR U7200 ( .A(n6186), .B(n6187), .Z(n6183) );
  AND U7201 ( .A(n6188), .B(n6189), .Z(n6186) );
  XNOR U7202 ( .A(x[1013]), .B(n6187), .Z(n6189) );
  XOR U7203 ( .A(n6190), .B(n6191), .Z(n6187) );
  AND U7204 ( .A(n6192), .B(n6193), .Z(n6190) );
  XNOR U7205 ( .A(x[1012]), .B(n6191), .Z(n6193) );
  XOR U7206 ( .A(n6194), .B(n6195), .Z(n6191) );
  AND U7207 ( .A(n6196), .B(n6197), .Z(n6194) );
  XNOR U7208 ( .A(x[1011]), .B(n6195), .Z(n6197) );
  XOR U7209 ( .A(n6198), .B(n6199), .Z(n6195) );
  AND U7210 ( .A(n6200), .B(n6201), .Z(n6198) );
  XNOR U7211 ( .A(x[1010]), .B(n6199), .Z(n6201) );
  XOR U7212 ( .A(n6202), .B(n6203), .Z(n6199) );
  AND U7213 ( .A(n6204), .B(n6205), .Z(n6202) );
  XNOR U7214 ( .A(x[1009]), .B(n6203), .Z(n6205) );
  XOR U7215 ( .A(n6206), .B(n6207), .Z(n6203) );
  AND U7216 ( .A(n6208), .B(n6209), .Z(n6206) );
  XNOR U7217 ( .A(x[1008]), .B(n6207), .Z(n6209) );
  XOR U7218 ( .A(n6210), .B(n6211), .Z(n6207) );
  AND U7219 ( .A(n6212), .B(n6213), .Z(n6210) );
  XNOR U7220 ( .A(x[1007]), .B(n6211), .Z(n6213) );
  XOR U7221 ( .A(n6214), .B(n6215), .Z(n6211) );
  AND U7222 ( .A(n6216), .B(n6217), .Z(n6214) );
  XNOR U7223 ( .A(x[1006]), .B(n6215), .Z(n6217) );
  XOR U7224 ( .A(n6218), .B(n6219), .Z(n6215) );
  AND U7225 ( .A(n6220), .B(n6221), .Z(n6218) );
  XNOR U7226 ( .A(x[1005]), .B(n6219), .Z(n6221) );
  XOR U7227 ( .A(n6222), .B(n6223), .Z(n6219) );
  AND U7228 ( .A(n6224), .B(n6225), .Z(n6222) );
  XNOR U7229 ( .A(x[1004]), .B(n6223), .Z(n6225) );
  XOR U7230 ( .A(n6226), .B(n6227), .Z(n6223) );
  AND U7231 ( .A(n6228), .B(n6229), .Z(n6226) );
  XNOR U7232 ( .A(x[1003]), .B(n6227), .Z(n6229) );
  XOR U7233 ( .A(n6230), .B(n6231), .Z(n6227) );
  AND U7234 ( .A(n6232), .B(n6233), .Z(n6230) );
  XNOR U7235 ( .A(x[1002]), .B(n6231), .Z(n6233) );
  XOR U7236 ( .A(n6234), .B(n6235), .Z(n6231) );
  AND U7237 ( .A(n6236), .B(n6237), .Z(n6234) );
  XNOR U7238 ( .A(x[1001]), .B(n6235), .Z(n6237) );
  XOR U7239 ( .A(n6238), .B(n6239), .Z(n6235) );
  AND U7240 ( .A(n6240), .B(n6241), .Z(n6238) );
  XNOR U7241 ( .A(x[1000]), .B(n6239), .Z(n6241) );
  XOR U7242 ( .A(n6242), .B(n6243), .Z(n6239) );
  AND U7243 ( .A(n6244), .B(n6245), .Z(n6242) );
  XNOR U7244 ( .A(x[999]), .B(n6243), .Z(n6245) );
  XOR U7245 ( .A(n6246), .B(n6247), .Z(n6243) );
  AND U7246 ( .A(n6248), .B(n6249), .Z(n6246) );
  XNOR U7247 ( .A(x[998]), .B(n6247), .Z(n6249) );
  XOR U7248 ( .A(n6250), .B(n6251), .Z(n6247) );
  AND U7249 ( .A(n6252), .B(n6253), .Z(n6250) );
  XNOR U7250 ( .A(x[997]), .B(n6251), .Z(n6253) );
  XOR U7251 ( .A(n6254), .B(n6255), .Z(n6251) );
  AND U7252 ( .A(n6256), .B(n6257), .Z(n6254) );
  XNOR U7253 ( .A(x[996]), .B(n6255), .Z(n6257) );
  XOR U7254 ( .A(n6258), .B(n6259), .Z(n6255) );
  AND U7255 ( .A(n6260), .B(n6261), .Z(n6258) );
  XNOR U7256 ( .A(x[995]), .B(n6259), .Z(n6261) );
  XOR U7257 ( .A(n6262), .B(n6263), .Z(n6259) );
  AND U7258 ( .A(n6264), .B(n6265), .Z(n6262) );
  XNOR U7259 ( .A(x[994]), .B(n6263), .Z(n6265) );
  XOR U7260 ( .A(n6266), .B(n6267), .Z(n6263) );
  AND U7261 ( .A(n6268), .B(n6269), .Z(n6266) );
  XNOR U7262 ( .A(x[993]), .B(n6267), .Z(n6269) );
  XOR U7263 ( .A(n6270), .B(n6271), .Z(n6267) );
  AND U7264 ( .A(n6272), .B(n6273), .Z(n6270) );
  XNOR U7265 ( .A(x[992]), .B(n6271), .Z(n6273) );
  XOR U7266 ( .A(n6274), .B(n6275), .Z(n6271) );
  AND U7267 ( .A(n6276), .B(n6277), .Z(n6274) );
  XNOR U7268 ( .A(x[991]), .B(n6275), .Z(n6277) );
  XOR U7269 ( .A(n6278), .B(n6279), .Z(n6275) );
  AND U7270 ( .A(n6280), .B(n6281), .Z(n6278) );
  XNOR U7271 ( .A(x[990]), .B(n6279), .Z(n6281) );
  XOR U7272 ( .A(n6282), .B(n6283), .Z(n6279) );
  AND U7273 ( .A(n6284), .B(n6285), .Z(n6282) );
  XNOR U7274 ( .A(x[989]), .B(n6283), .Z(n6285) );
  XOR U7275 ( .A(n6286), .B(n6287), .Z(n6283) );
  AND U7276 ( .A(n6288), .B(n6289), .Z(n6286) );
  XNOR U7277 ( .A(x[988]), .B(n6287), .Z(n6289) );
  XOR U7278 ( .A(n6290), .B(n6291), .Z(n6287) );
  AND U7279 ( .A(n6292), .B(n6293), .Z(n6290) );
  XNOR U7280 ( .A(x[987]), .B(n6291), .Z(n6293) );
  XOR U7281 ( .A(n6294), .B(n6295), .Z(n6291) );
  AND U7282 ( .A(n6296), .B(n6297), .Z(n6294) );
  XNOR U7283 ( .A(x[986]), .B(n6295), .Z(n6297) );
  XOR U7284 ( .A(n6298), .B(n6299), .Z(n6295) );
  AND U7285 ( .A(n6300), .B(n6301), .Z(n6298) );
  XNOR U7286 ( .A(x[985]), .B(n6299), .Z(n6301) );
  XOR U7287 ( .A(n6302), .B(n6303), .Z(n6299) );
  AND U7288 ( .A(n6304), .B(n6305), .Z(n6302) );
  XNOR U7289 ( .A(x[984]), .B(n6303), .Z(n6305) );
  XOR U7290 ( .A(n6306), .B(n6307), .Z(n6303) );
  AND U7291 ( .A(n6308), .B(n6309), .Z(n6306) );
  XNOR U7292 ( .A(x[983]), .B(n6307), .Z(n6309) );
  XOR U7293 ( .A(n6310), .B(n6311), .Z(n6307) );
  AND U7294 ( .A(n6312), .B(n6313), .Z(n6310) );
  XNOR U7295 ( .A(x[982]), .B(n6311), .Z(n6313) );
  XOR U7296 ( .A(n6314), .B(n6315), .Z(n6311) );
  AND U7297 ( .A(n6316), .B(n6317), .Z(n6314) );
  XNOR U7298 ( .A(x[981]), .B(n6315), .Z(n6317) );
  XOR U7299 ( .A(n6318), .B(n6319), .Z(n6315) );
  AND U7300 ( .A(n6320), .B(n6321), .Z(n6318) );
  XNOR U7301 ( .A(x[980]), .B(n6319), .Z(n6321) );
  XOR U7302 ( .A(n6322), .B(n6323), .Z(n6319) );
  AND U7303 ( .A(n6324), .B(n6325), .Z(n6322) );
  XNOR U7304 ( .A(x[979]), .B(n6323), .Z(n6325) );
  XOR U7305 ( .A(n6326), .B(n6327), .Z(n6323) );
  AND U7306 ( .A(n6328), .B(n6329), .Z(n6326) );
  XNOR U7307 ( .A(x[978]), .B(n6327), .Z(n6329) );
  XOR U7308 ( .A(n6330), .B(n6331), .Z(n6327) );
  AND U7309 ( .A(n6332), .B(n6333), .Z(n6330) );
  XNOR U7310 ( .A(x[977]), .B(n6331), .Z(n6333) );
  XOR U7311 ( .A(n6334), .B(n6335), .Z(n6331) );
  AND U7312 ( .A(n6336), .B(n6337), .Z(n6334) );
  XNOR U7313 ( .A(x[976]), .B(n6335), .Z(n6337) );
  XOR U7314 ( .A(n6338), .B(n6339), .Z(n6335) );
  AND U7315 ( .A(n6340), .B(n6341), .Z(n6338) );
  XNOR U7316 ( .A(x[975]), .B(n6339), .Z(n6341) );
  XOR U7317 ( .A(n6342), .B(n6343), .Z(n6339) );
  AND U7318 ( .A(n6344), .B(n6345), .Z(n6342) );
  XNOR U7319 ( .A(x[974]), .B(n6343), .Z(n6345) );
  XOR U7320 ( .A(n6346), .B(n6347), .Z(n6343) );
  AND U7321 ( .A(n6348), .B(n6349), .Z(n6346) );
  XNOR U7322 ( .A(x[973]), .B(n6347), .Z(n6349) );
  XOR U7323 ( .A(n6350), .B(n6351), .Z(n6347) );
  AND U7324 ( .A(n6352), .B(n6353), .Z(n6350) );
  XNOR U7325 ( .A(x[972]), .B(n6351), .Z(n6353) );
  XOR U7326 ( .A(n6354), .B(n6355), .Z(n6351) );
  AND U7327 ( .A(n6356), .B(n6357), .Z(n6354) );
  XNOR U7328 ( .A(x[971]), .B(n6355), .Z(n6357) );
  XOR U7329 ( .A(n6358), .B(n6359), .Z(n6355) );
  AND U7330 ( .A(n6360), .B(n6361), .Z(n6358) );
  XNOR U7331 ( .A(x[970]), .B(n6359), .Z(n6361) );
  XOR U7332 ( .A(n6362), .B(n6363), .Z(n6359) );
  AND U7333 ( .A(n6364), .B(n6365), .Z(n6362) );
  XNOR U7334 ( .A(x[969]), .B(n6363), .Z(n6365) );
  XOR U7335 ( .A(n6366), .B(n6367), .Z(n6363) );
  AND U7336 ( .A(n6368), .B(n6369), .Z(n6366) );
  XNOR U7337 ( .A(x[968]), .B(n6367), .Z(n6369) );
  XOR U7338 ( .A(n6370), .B(n6371), .Z(n6367) );
  AND U7339 ( .A(n6372), .B(n6373), .Z(n6370) );
  XNOR U7340 ( .A(x[967]), .B(n6371), .Z(n6373) );
  XOR U7341 ( .A(n6374), .B(n6375), .Z(n6371) );
  AND U7342 ( .A(n6376), .B(n6377), .Z(n6374) );
  XNOR U7343 ( .A(x[966]), .B(n6375), .Z(n6377) );
  XOR U7344 ( .A(n6378), .B(n6379), .Z(n6375) );
  AND U7345 ( .A(n6380), .B(n6381), .Z(n6378) );
  XNOR U7346 ( .A(x[965]), .B(n6379), .Z(n6381) );
  XOR U7347 ( .A(n6382), .B(n6383), .Z(n6379) );
  AND U7348 ( .A(n6384), .B(n6385), .Z(n6382) );
  XNOR U7349 ( .A(x[964]), .B(n6383), .Z(n6385) );
  XOR U7350 ( .A(n6386), .B(n6387), .Z(n6383) );
  AND U7351 ( .A(n6388), .B(n6389), .Z(n6386) );
  XNOR U7352 ( .A(x[963]), .B(n6387), .Z(n6389) );
  XOR U7353 ( .A(n6390), .B(n6391), .Z(n6387) );
  AND U7354 ( .A(n6392), .B(n6393), .Z(n6390) );
  XNOR U7355 ( .A(x[962]), .B(n6391), .Z(n6393) );
  XOR U7356 ( .A(n6394), .B(n6395), .Z(n6391) );
  AND U7357 ( .A(n6396), .B(n6397), .Z(n6394) );
  XNOR U7358 ( .A(x[961]), .B(n6395), .Z(n6397) );
  XOR U7359 ( .A(n6398), .B(n6399), .Z(n6395) );
  AND U7360 ( .A(n6400), .B(n6401), .Z(n6398) );
  XNOR U7361 ( .A(x[960]), .B(n6399), .Z(n6401) );
  XOR U7362 ( .A(n6402), .B(n6403), .Z(n6399) );
  AND U7363 ( .A(n6404), .B(n6405), .Z(n6402) );
  XNOR U7364 ( .A(x[959]), .B(n6403), .Z(n6405) );
  XOR U7365 ( .A(n6406), .B(n6407), .Z(n6403) );
  AND U7366 ( .A(n6408), .B(n6409), .Z(n6406) );
  XNOR U7367 ( .A(x[958]), .B(n6407), .Z(n6409) );
  XOR U7368 ( .A(n6410), .B(n6411), .Z(n6407) );
  AND U7369 ( .A(n6412), .B(n6413), .Z(n6410) );
  XNOR U7370 ( .A(x[957]), .B(n6411), .Z(n6413) );
  XOR U7371 ( .A(n6414), .B(n6415), .Z(n6411) );
  AND U7372 ( .A(n6416), .B(n6417), .Z(n6414) );
  XNOR U7373 ( .A(x[956]), .B(n6415), .Z(n6417) );
  XOR U7374 ( .A(n6418), .B(n6419), .Z(n6415) );
  AND U7375 ( .A(n6420), .B(n6421), .Z(n6418) );
  XNOR U7376 ( .A(x[955]), .B(n6419), .Z(n6421) );
  XOR U7377 ( .A(n6422), .B(n6423), .Z(n6419) );
  AND U7378 ( .A(n6424), .B(n6425), .Z(n6422) );
  XNOR U7379 ( .A(x[954]), .B(n6423), .Z(n6425) );
  XOR U7380 ( .A(n6426), .B(n6427), .Z(n6423) );
  AND U7381 ( .A(n6428), .B(n6429), .Z(n6426) );
  XNOR U7382 ( .A(x[953]), .B(n6427), .Z(n6429) );
  XOR U7383 ( .A(n6430), .B(n6431), .Z(n6427) );
  AND U7384 ( .A(n6432), .B(n6433), .Z(n6430) );
  XNOR U7385 ( .A(x[952]), .B(n6431), .Z(n6433) );
  XOR U7386 ( .A(n6434), .B(n6435), .Z(n6431) );
  AND U7387 ( .A(n6436), .B(n6437), .Z(n6434) );
  XNOR U7388 ( .A(x[951]), .B(n6435), .Z(n6437) );
  XOR U7389 ( .A(n6438), .B(n6439), .Z(n6435) );
  AND U7390 ( .A(n6440), .B(n6441), .Z(n6438) );
  XNOR U7391 ( .A(x[950]), .B(n6439), .Z(n6441) );
  XOR U7392 ( .A(n6442), .B(n6443), .Z(n6439) );
  AND U7393 ( .A(n6444), .B(n6445), .Z(n6442) );
  XNOR U7394 ( .A(x[949]), .B(n6443), .Z(n6445) );
  XOR U7395 ( .A(n6446), .B(n6447), .Z(n6443) );
  AND U7396 ( .A(n6448), .B(n6449), .Z(n6446) );
  XNOR U7397 ( .A(x[948]), .B(n6447), .Z(n6449) );
  XOR U7398 ( .A(n6450), .B(n6451), .Z(n6447) );
  AND U7399 ( .A(n6452), .B(n6453), .Z(n6450) );
  XNOR U7400 ( .A(x[947]), .B(n6451), .Z(n6453) );
  XOR U7401 ( .A(n6454), .B(n6455), .Z(n6451) );
  AND U7402 ( .A(n6456), .B(n6457), .Z(n6454) );
  XNOR U7403 ( .A(x[946]), .B(n6455), .Z(n6457) );
  XOR U7404 ( .A(n6458), .B(n6459), .Z(n6455) );
  AND U7405 ( .A(n6460), .B(n6461), .Z(n6458) );
  XNOR U7406 ( .A(x[945]), .B(n6459), .Z(n6461) );
  XOR U7407 ( .A(n6462), .B(n6463), .Z(n6459) );
  AND U7408 ( .A(n6464), .B(n6465), .Z(n6462) );
  XNOR U7409 ( .A(x[944]), .B(n6463), .Z(n6465) );
  XOR U7410 ( .A(n6466), .B(n6467), .Z(n6463) );
  AND U7411 ( .A(n6468), .B(n6469), .Z(n6466) );
  XNOR U7412 ( .A(x[943]), .B(n6467), .Z(n6469) );
  XOR U7413 ( .A(n6470), .B(n6471), .Z(n6467) );
  AND U7414 ( .A(n6472), .B(n6473), .Z(n6470) );
  XNOR U7415 ( .A(x[942]), .B(n6471), .Z(n6473) );
  XOR U7416 ( .A(n6474), .B(n6475), .Z(n6471) );
  AND U7417 ( .A(n6476), .B(n6477), .Z(n6474) );
  XNOR U7418 ( .A(x[941]), .B(n6475), .Z(n6477) );
  XOR U7419 ( .A(n6478), .B(n6479), .Z(n6475) );
  AND U7420 ( .A(n6480), .B(n6481), .Z(n6478) );
  XNOR U7421 ( .A(x[940]), .B(n6479), .Z(n6481) );
  XOR U7422 ( .A(n6482), .B(n6483), .Z(n6479) );
  AND U7423 ( .A(n6484), .B(n6485), .Z(n6482) );
  XNOR U7424 ( .A(x[939]), .B(n6483), .Z(n6485) );
  XOR U7425 ( .A(n6486), .B(n6487), .Z(n6483) );
  AND U7426 ( .A(n6488), .B(n6489), .Z(n6486) );
  XNOR U7427 ( .A(x[938]), .B(n6487), .Z(n6489) );
  XOR U7428 ( .A(n6490), .B(n6491), .Z(n6487) );
  AND U7429 ( .A(n6492), .B(n6493), .Z(n6490) );
  XNOR U7430 ( .A(x[937]), .B(n6491), .Z(n6493) );
  XOR U7431 ( .A(n6494), .B(n6495), .Z(n6491) );
  AND U7432 ( .A(n6496), .B(n6497), .Z(n6494) );
  XNOR U7433 ( .A(x[936]), .B(n6495), .Z(n6497) );
  XOR U7434 ( .A(n6498), .B(n6499), .Z(n6495) );
  AND U7435 ( .A(n6500), .B(n6501), .Z(n6498) );
  XNOR U7436 ( .A(x[935]), .B(n6499), .Z(n6501) );
  XOR U7437 ( .A(n6502), .B(n6503), .Z(n6499) );
  AND U7438 ( .A(n6504), .B(n6505), .Z(n6502) );
  XNOR U7439 ( .A(x[934]), .B(n6503), .Z(n6505) );
  XOR U7440 ( .A(n6506), .B(n6507), .Z(n6503) );
  AND U7441 ( .A(n6508), .B(n6509), .Z(n6506) );
  XNOR U7442 ( .A(x[933]), .B(n6507), .Z(n6509) );
  XOR U7443 ( .A(n6510), .B(n6511), .Z(n6507) );
  AND U7444 ( .A(n6512), .B(n6513), .Z(n6510) );
  XNOR U7445 ( .A(x[932]), .B(n6511), .Z(n6513) );
  XOR U7446 ( .A(n6514), .B(n6515), .Z(n6511) );
  AND U7447 ( .A(n6516), .B(n6517), .Z(n6514) );
  XNOR U7448 ( .A(x[931]), .B(n6515), .Z(n6517) );
  XOR U7449 ( .A(n6518), .B(n6519), .Z(n6515) );
  AND U7450 ( .A(n6520), .B(n6521), .Z(n6518) );
  XNOR U7451 ( .A(x[930]), .B(n6519), .Z(n6521) );
  XOR U7452 ( .A(n6522), .B(n6523), .Z(n6519) );
  AND U7453 ( .A(n6524), .B(n6525), .Z(n6522) );
  XNOR U7454 ( .A(x[929]), .B(n6523), .Z(n6525) );
  XOR U7455 ( .A(n6526), .B(n6527), .Z(n6523) );
  AND U7456 ( .A(n6528), .B(n6529), .Z(n6526) );
  XNOR U7457 ( .A(x[928]), .B(n6527), .Z(n6529) );
  XOR U7458 ( .A(n6530), .B(n6531), .Z(n6527) );
  AND U7459 ( .A(n6532), .B(n6533), .Z(n6530) );
  XNOR U7460 ( .A(x[927]), .B(n6531), .Z(n6533) );
  XOR U7461 ( .A(n6534), .B(n6535), .Z(n6531) );
  AND U7462 ( .A(n6536), .B(n6537), .Z(n6534) );
  XNOR U7463 ( .A(x[926]), .B(n6535), .Z(n6537) );
  XOR U7464 ( .A(n6538), .B(n6539), .Z(n6535) );
  AND U7465 ( .A(n6540), .B(n6541), .Z(n6538) );
  XNOR U7466 ( .A(x[925]), .B(n6539), .Z(n6541) );
  XOR U7467 ( .A(n6542), .B(n6543), .Z(n6539) );
  AND U7468 ( .A(n6544), .B(n6545), .Z(n6542) );
  XNOR U7469 ( .A(x[924]), .B(n6543), .Z(n6545) );
  XOR U7470 ( .A(n6546), .B(n6547), .Z(n6543) );
  AND U7471 ( .A(n6548), .B(n6549), .Z(n6546) );
  XNOR U7472 ( .A(x[923]), .B(n6547), .Z(n6549) );
  XOR U7473 ( .A(n6550), .B(n6551), .Z(n6547) );
  AND U7474 ( .A(n6552), .B(n6553), .Z(n6550) );
  XNOR U7475 ( .A(x[922]), .B(n6551), .Z(n6553) );
  XOR U7476 ( .A(n6554), .B(n6555), .Z(n6551) );
  AND U7477 ( .A(n6556), .B(n6557), .Z(n6554) );
  XNOR U7478 ( .A(x[921]), .B(n6555), .Z(n6557) );
  XOR U7479 ( .A(n6558), .B(n6559), .Z(n6555) );
  AND U7480 ( .A(n6560), .B(n6561), .Z(n6558) );
  XNOR U7481 ( .A(x[920]), .B(n6559), .Z(n6561) );
  XOR U7482 ( .A(n6562), .B(n6563), .Z(n6559) );
  AND U7483 ( .A(n6564), .B(n6565), .Z(n6562) );
  XNOR U7484 ( .A(x[919]), .B(n6563), .Z(n6565) );
  XOR U7485 ( .A(n6566), .B(n6567), .Z(n6563) );
  AND U7486 ( .A(n6568), .B(n6569), .Z(n6566) );
  XNOR U7487 ( .A(x[918]), .B(n6567), .Z(n6569) );
  XOR U7488 ( .A(n6570), .B(n6571), .Z(n6567) );
  AND U7489 ( .A(n6572), .B(n6573), .Z(n6570) );
  XNOR U7490 ( .A(x[917]), .B(n6571), .Z(n6573) );
  XOR U7491 ( .A(n6574), .B(n6575), .Z(n6571) );
  AND U7492 ( .A(n6576), .B(n6577), .Z(n6574) );
  XNOR U7493 ( .A(x[916]), .B(n6575), .Z(n6577) );
  XOR U7494 ( .A(n6578), .B(n6579), .Z(n6575) );
  AND U7495 ( .A(n6580), .B(n6581), .Z(n6578) );
  XNOR U7496 ( .A(x[915]), .B(n6579), .Z(n6581) );
  XOR U7497 ( .A(n6582), .B(n6583), .Z(n6579) );
  AND U7498 ( .A(n6584), .B(n6585), .Z(n6582) );
  XNOR U7499 ( .A(x[914]), .B(n6583), .Z(n6585) );
  XOR U7500 ( .A(n6586), .B(n6587), .Z(n6583) );
  AND U7501 ( .A(n6588), .B(n6589), .Z(n6586) );
  XNOR U7502 ( .A(x[913]), .B(n6587), .Z(n6589) );
  XOR U7503 ( .A(n6590), .B(n6591), .Z(n6587) );
  AND U7504 ( .A(n6592), .B(n6593), .Z(n6590) );
  XNOR U7505 ( .A(x[912]), .B(n6591), .Z(n6593) );
  XOR U7506 ( .A(n6594), .B(n6595), .Z(n6591) );
  AND U7507 ( .A(n6596), .B(n6597), .Z(n6594) );
  XNOR U7508 ( .A(x[911]), .B(n6595), .Z(n6597) );
  XOR U7509 ( .A(n6598), .B(n6599), .Z(n6595) );
  AND U7510 ( .A(n6600), .B(n6601), .Z(n6598) );
  XNOR U7511 ( .A(x[910]), .B(n6599), .Z(n6601) );
  XOR U7512 ( .A(n6602), .B(n6603), .Z(n6599) );
  AND U7513 ( .A(n6604), .B(n6605), .Z(n6602) );
  XNOR U7514 ( .A(x[909]), .B(n6603), .Z(n6605) );
  XOR U7515 ( .A(n6606), .B(n6607), .Z(n6603) );
  AND U7516 ( .A(n6608), .B(n6609), .Z(n6606) );
  XNOR U7517 ( .A(x[908]), .B(n6607), .Z(n6609) );
  XOR U7518 ( .A(n6610), .B(n6611), .Z(n6607) );
  AND U7519 ( .A(n6612), .B(n6613), .Z(n6610) );
  XNOR U7520 ( .A(x[907]), .B(n6611), .Z(n6613) );
  XOR U7521 ( .A(n6614), .B(n6615), .Z(n6611) );
  AND U7522 ( .A(n6616), .B(n6617), .Z(n6614) );
  XNOR U7523 ( .A(x[906]), .B(n6615), .Z(n6617) );
  XOR U7524 ( .A(n6618), .B(n6619), .Z(n6615) );
  AND U7525 ( .A(n6620), .B(n6621), .Z(n6618) );
  XNOR U7526 ( .A(x[905]), .B(n6619), .Z(n6621) );
  XOR U7527 ( .A(n6622), .B(n6623), .Z(n6619) );
  AND U7528 ( .A(n6624), .B(n6625), .Z(n6622) );
  XNOR U7529 ( .A(x[904]), .B(n6623), .Z(n6625) );
  XOR U7530 ( .A(n6626), .B(n6627), .Z(n6623) );
  AND U7531 ( .A(n6628), .B(n6629), .Z(n6626) );
  XNOR U7532 ( .A(x[903]), .B(n6627), .Z(n6629) );
  XOR U7533 ( .A(n6630), .B(n6631), .Z(n6627) );
  AND U7534 ( .A(n6632), .B(n6633), .Z(n6630) );
  XNOR U7535 ( .A(x[902]), .B(n6631), .Z(n6633) );
  XOR U7536 ( .A(n6634), .B(n6635), .Z(n6631) );
  AND U7537 ( .A(n6636), .B(n6637), .Z(n6634) );
  XNOR U7538 ( .A(x[901]), .B(n6635), .Z(n6637) );
  XOR U7539 ( .A(n6638), .B(n6639), .Z(n6635) );
  AND U7540 ( .A(n6640), .B(n6641), .Z(n6638) );
  XNOR U7541 ( .A(x[900]), .B(n6639), .Z(n6641) );
  XOR U7542 ( .A(n6642), .B(n6643), .Z(n6639) );
  AND U7543 ( .A(n6644), .B(n6645), .Z(n6642) );
  XNOR U7544 ( .A(x[899]), .B(n6643), .Z(n6645) );
  XOR U7545 ( .A(n6646), .B(n6647), .Z(n6643) );
  AND U7546 ( .A(n6648), .B(n6649), .Z(n6646) );
  XNOR U7547 ( .A(x[898]), .B(n6647), .Z(n6649) );
  XOR U7548 ( .A(n6650), .B(n6651), .Z(n6647) );
  AND U7549 ( .A(n6652), .B(n6653), .Z(n6650) );
  XNOR U7550 ( .A(x[897]), .B(n6651), .Z(n6653) );
  XOR U7551 ( .A(n6654), .B(n6655), .Z(n6651) );
  AND U7552 ( .A(n6656), .B(n6657), .Z(n6654) );
  XNOR U7553 ( .A(x[896]), .B(n6655), .Z(n6657) );
  XOR U7554 ( .A(n6658), .B(n6659), .Z(n6655) );
  AND U7555 ( .A(n6660), .B(n6661), .Z(n6658) );
  XNOR U7556 ( .A(x[895]), .B(n6659), .Z(n6661) );
  XOR U7557 ( .A(n6662), .B(n6663), .Z(n6659) );
  AND U7558 ( .A(n6664), .B(n6665), .Z(n6662) );
  XNOR U7559 ( .A(x[894]), .B(n6663), .Z(n6665) );
  XOR U7560 ( .A(n6666), .B(n6667), .Z(n6663) );
  AND U7561 ( .A(n6668), .B(n6669), .Z(n6666) );
  XNOR U7562 ( .A(x[893]), .B(n6667), .Z(n6669) );
  XOR U7563 ( .A(n6670), .B(n6671), .Z(n6667) );
  AND U7564 ( .A(n6672), .B(n6673), .Z(n6670) );
  XNOR U7565 ( .A(x[892]), .B(n6671), .Z(n6673) );
  XOR U7566 ( .A(n6674), .B(n6675), .Z(n6671) );
  AND U7567 ( .A(n6676), .B(n6677), .Z(n6674) );
  XNOR U7568 ( .A(x[891]), .B(n6675), .Z(n6677) );
  XOR U7569 ( .A(n6678), .B(n6679), .Z(n6675) );
  AND U7570 ( .A(n6680), .B(n6681), .Z(n6678) );
  XNOR U7571 ( .A(x[890]), .B(n6679), .Z(n6681) );
  XOR U7572 ( .A(n6682), .B(n6683), .Z(n6679) );
  AND U7573 ( .A(n6684), .B(n6685), .Z(n6682) );
  XNOR U7574 ( .A(x[889]), .B(n6683), .Z(n6685) );
  XOR U7575 ( .A(n6686), .B(n6687), .Z(n6683) );
  AND U7576 ( .A(n6688), .B(n6689), .Z(n6686) );
  XNOR U7577 ( .A(x[888]), .B(n6687), .Z(n6689) );
  XOR U7578 ( .A(n6690), .B(n6691), .Z(n6687) );
  AND U7579 ( .A(n6692), .B(n6693), .Z(n6690) );
  XNOR U7580 ( .A(x[887]), .B(n6691), .Z(n6693) );
  XOR U7581 ( .A(n6694), .B(n6695), .Z(n6691) );
  AND U7582 ( .A(n6696), .B(n6697), .Z(n6694) );
  XNOR U7583 ( .A(x[886]), .B(n6695), .Z(n6697) );
  XOR U7584 ( .A(n6698), .B(n6699), .Z(n6695) );
  AND U7585 ( .A(n6700), .B(n6701), .Z(n6698) );
  XNOR U7586 ( .A(x[885]), .B(n6699), .Z(n6701) );
  XOR U7587 ( .A(n6702), .B(n6703), .Z(n6699) );
  AND U7588 ( .A(n6704), .B(n6705), .Z(n6702) );
  XNOR U7589 ( .A(x[884]), .B(n6703), .Z(n6705) );
  XOR U7590 ( .A(n6706), .B(n6707), .Z(n6703) );
  AND U7591 ( .A(n6708), .B(n6709), .Z(n6706) );
  XNOR U7592 ( .A(x[883]), .B(n6707), .Z(n6709) );
  XOR U7593 ( .A(n6710), .B(n6711), .Z(n6707) );
  AND U7594 ( .A(n6712), .B(n6713), .Z(n6710) );
  XNOR U7595 ( .A(x[882]), .B(n6711), .Z(n6713) );
  XOR U7596 ( .A(n6714), .B(n6715), .Z(n6711) );
  AND U7597 ( .A(n6716), .B(n6717), .Z(n6714) );
  XNOR U7598 ( .A(x[881]), .B(n6715), .Z(n6717) );
  XOR U7599 ( .A(n6718), .B(n6719), .Z(n6715) );
  AND U7600 ( .A(n6720), .B(n6721), .Z(n6718) );
  XNOR U7601 ( .A(x[880]), .B(n6719), .Z(n6721) );
  XOR U7602 ( .A(n6722), .B(n6723), .Z(n6719) );
  AND U7603 ( .A(n6724), .B(n6725), .Z(n6722) );
  XNOR U7604 ( .A(x[879]), .B(n6723), .Z(n6725) );
  XOR U7605 ( .A(n6726), .B(n6727), .Z(n6723) );
  AND U7606 ( .A(n6728), .B(n6729), .Z(n6726) );
  XNOR U7607 ( .A(x[878]), .B(n6727), .Z(n6729) );
  XOR U7608 ( .A(n6730), .B(n6731), .Z(n6727) );
  AND U7609 ( .A(n6732), .B(n6733), .Z(n6730) );
  XNOR U7610 ( .A(x[877]), .B(n6731), .Z(n6733) );
  XOR U7611 ( .A(n6734), .B(n6735), .Z(n6731) );
  AND U7612 ( .A(n6736), .B(n6737), .Z(n6734) );
  XNOR U7613 ( .A(x[876]), .B(n6735), .Z(n6737) );
  XOR U7614 ( .A(n6738), .B(n6739), .Z(n6735) );
  AND U7615 ( .A(n6740), .B(n6741), .Z(n6738) );
  XNOR U7616 ( .A(x[875]), .B(n6739), .Z(n6741) );
  XOR U7617 ( .A(n6742), .B(n6743), .Z(n6739) );
  AND U7618 ( .A(n6744), .B(n6745), .Z(n6742) );
  XNOR U7619 ( .A(x[874]), .B(n6743), .Z(n6745) );
  XOR U7620 ( .A(n6746), .B(n6747), .Z(n6743) );
  AND U7621 ( .A(n6748), .B(n6749), .Z(n6746) );
  XNOR U7622 ( .A(x[873]), .B(n6747), .Z(n6749) );
  XOR U7623 ( .A(n6750), .B(n6751), .Z(n6747) );
  AND U7624 ( .A(n6752), .B(n6753), .Z(n6750) );
  XNOR U7625 ( .A(x[872]), .B(n6751), .Z(n6753) );
  XOR U7626 ( .A(n6754), .B(n6755), .Z(n6751) );
  AND U7627 ( .A(n6756), .B(n6757), .Z(n6754) );
  XNOR U7628 ( .A(x[871]), .B(n6755), .Z(n6757) );
  XOR U7629 ( .A(n6758), .B(n6759), .Z(n6755) );
  AND U7630 ( .A(n6760), .B(n6761), .Z(n6758) );
  XNOR U7631 ( .A(x[870]), .B(n6759), .Z(n6761) );
  XOR U7632 ( .A(n6762), .B(n6763), .Z(n6759) );
  AND U7633 ( .A(n6764), .B(n6765), .Z(n6762) );
  XNOR U7634 ( .A(x[869]), .B(n6763), .Z(n6765) );
  XOR U7635 ( .A(n6766), .B(n6767), .Z(n6763) );
  AND U7636 ( .A(n6768), .B(n6769), .Z(n6766) );
  XNOR U7637 ( .A(x[868]), .B(n6767), .Z(n6769) );
  XOR U7638 ( .A(n6770), .B(n6771), .Z(n6767) );
  AND U7639 ( .A(n6772), .B(n6773), .Z(n6770) );
  XNOR U7640 ( .A(x[867]), .B(n6771), .Z(n6773) );
  XOR U7641 ( .A(n6774), .B(n6775), .Z(n6771) );
  AND U7642 ( .A(n6776), .B(n6777), .Z(n6774) );
  XNOR U7643 ( .A(x[866]), .B(n6775), .Z(n6777) );
  XOR U7644 ( .A(n6778), .B(n6779), .Z(n6775) );
  AND U7645 ( .A(n6780), .B(n6781), .Z(n6778) );
  XNOR U7646 ( .A(x[865]), .B(n6779), .Z(n6781) );
  XOR U7647 ( .A(n6782), .B(n6783), .Z(n6779) );
  AND U7648 ( .A(n6784), .B(n6785), .Z(n6782) );
  XNOR U7649 ( .A(x[864]), .B(n6783), .Z(n6785) );
  XOR U7650 ( .A(n6786), .B(n6787), .Z(n6783) );
  AND U7651 ( .A(n6788), .B(n6789), .Z(n6786) );
  XNOR U7652 ( .A(x[863]), .B(n6787), .Z(n6789) );
  XOR U7653 ( .A(n6790), .B(n6791), .Z(n6787) );
  AND U7654 ( .A(n6792), .B(n6793), .Z(n6790) );
  XNOR U7655 ( .A(x[862]), .B(n6791), .Z(n6793) );
  XOR U7656 ( .A(n6794), .B(n6795), .Z(n6791) );
  AND U7657 ( .A(n6796), .B(n6797), .Z(n6794) );
  XNOR U7658 ( .A(x[861]), .B(n6795), .Z(n6797) );
  XOR U7659 ( .A(n6798), .B(n6799), .Z(n6795) );
  AND U7660 ( .A(n6800), .B(n6801), .Z(n6798) );
  XNOR U7661 ( .A(x[860]), .B(n6799), .Z(n6801) );
  XOR U7662 ( .A(n6802), .B(n6803), .Z(n6799) );
  AND U7663 ( .A(n6804), .B(n6805), .Z(n6802) );
  XNOR U7664 ( .A(x[859]), .B(n6803), .Z(n6805) );
  XOR U7665 ( .A(n6806), .B(n6807), .Z(n6803) );
  AND U7666 ( .A(n6808), .B(n6809), .Z(n6806) );
  XNOR U7667 ( .A(x[858]), .B(n6807), .Z(n6809) );
  XOR U7668 ( .A(n6810), .B(n6811), .Z(n6807) );
  AND U7669 ( .A(n6812), .B(n6813), .Z(n6810) );
  XNOR U7670 ( .A(x[857]), .B(n6811), .Z(n6813) );
  XOR U7671 ( .A(n6814), .B(n6815), .Z(n6811) );
  AND U7672 ( .A(n6816), .B(n6817), .Z(n6814) );
  XNOR U7673 ( .A(x[856]), .B(n6815), .Z(n6817) );
  XOR U7674 ( .A(n6818), .B(n6819), .Z(n6815) );
  AND U7675 ( .A(n6820), .B(n6821), .Z(n6818) );
  XNOR U7676 ( .A(x[855]), .B(n6819), .Z(n6821) );
  XOR U7677 ( .A(n6822), .B(n6823), .Z(n6819) );
  AND U7678 ( .A(n6824), .B(n6825), .Z(n6822) );
  XNOR U7679 ( .A(x[854]), .B(n6823), .Z(n6825) );
  XOR U7680 ( .A(n6826), .B(n6827), .Z(n6823) );
  AND U7681 ( .A(n6828), .B(n6829), .Z(n6826) );
  XNOR U7682 ( .A(x[853]), .B(n6827), .Z(n6829) );
  XOR U7683 ( .A(n6830), .B(n6831), .Z(n6827) );
  AND U7684 ( .A(n6832), .B(n6833), .Z(n6830) );
  XNOR U7685 ( .A(x[852]), .B(n6831), .Z(n6833) );
  XOR U7686 ( .A(n6834), .B(n6835), .Z(n6831) );
  AND U7687 ( .A(n6836), .B(n6837), .Z(n6834) );
  XNOR U7688 ( .A(x[851]), .B(n6835), .Z(n6837) );
  XOR U7689 ( .A(n6838), .B(n6839), .Z(n6835) );
  AND U7690 ( .A(n6840), .B(n6841), .Z(n6838) );
  XNOR U7691 ( .A(x[850]), .B(n6839), .Z(n6841) );
  XOR U7692 ( .A(n6842), .B(n6843), .Z(n6839) );
  AND U7693 ( .A(n6844), .B(n6845), .Z(n6842) );
  XNOR U7694 ( .A(x[849]), .B(n6843), .Z(n6845) );
  XOR U7695 ( .A(n6846), .B(n6847), .Z(n6843) );
  AND U7696 ( .A(n6848), .B(n6849), .Z(n6846) );
  XNOR U7697 ( .A(x[848]), .B(n6847), .Z(n6849) );
  XOR U7698 ( .A(n6850), .B(n6851), .Z(n6847) );
  AND U7699 ( .A(n6852), .B(n6853), .Z(n6850) );
  XNOR U7700 ( .A(x[847]), .B(n6851), .Z(n6853) );
  XOR U7701 ( .A(n6854), .B(n6855), .Z(n6851) );
  AND U7702 ( .A(n6856), .B(n6857), .Z(n6854) );
  XNOR U7703 ( .A(x[846]), .B(n6855), .Z(n6857) );
  XOR U7704 ( .A(n6858), .B(n6859), .Z(n6855) );
  AND U7705 ( .A(n6860), .B(n6861), .Z(n6858) );
  XNOR U7706 ( .A(x[845]), .B(n6859), .Z(n6861) );
  XOR U7707 ( .A(n6862), .B(n6863), .Z(n6859) );
  AND U7708 ( .A(n6864), .B(n6865), .Z(n6862) );
  XNOR U7709 ( .A(x[844]), .B(n6863), .Z(n6865) );
  XOR U7710 ( .A(n6866), .B(n6867), .Z(n6863) );
  AND U7711 ( .A(n6868), .B(n6869), .Z(n6866) );
  XNOR U7712 ( .A(x[843]), .B(n6867), .Z(n6869) );
  XOR U7713 ( .A(n6870), .B(n6871), .Z(n6867) );
  AND U7714 ( .A(n6872), .B(n6873), .Z(n6870) );
  XNOR U7715 ( .A(x[842]), .B(n6871), .Z(n6873) );
  XOR U7716 ( .A(n6874), .B(n6875), .Z(n6871) );
  AND U7717 ( .A(n6876), .B(n6877), .Z(n6874) );
  XNOR U7718 ( .A(x[841]), .B(n6875), .Z(n6877) );
  XOR U7719 ( .A(n6878), .B(n6879), .Z(n6875) );
  AND U7720 ( .A(n6880), .B(n6881), .Z(n6878) );
  XNOR U7721 ( .A(x[840]), .B(n6879), .Z(n6881) );
  XOR U7722 ( .A(n6882), .B(n6883), .Z(n6879) );
  AND U7723 ( .A(n6884), .B(n6885), .Z(n6882) );
  XNOR U7724 ( .A(x[839]), .B(n6883), .Z(n6885) );
  XOR U7725 ( .A(n6886), .B(n6887), .Z(n6883) );
  AND U7726 ( .A(n6888), .B(n6889), .Z(n6886) );
  XNOR U7727 ( .A(x[838]), .B(n6887), .Z(n6889) );
  XOR U7728 ( .A(n6890), .B(n6891), .Z(n6887) );
  AND U7729 ( .A(n6892), .B(n6893), .Z(n6890) );
  XNOR U7730 ( .A(x[837]), .B(n6891), .Z(n6893) );
  XOR U7731 ( .A(n6894), .B(n6895), .Z(n6891) );
  AND U7732 ( .A(n6896), .B(n6897), .Z(n6894) );
  XNOR U7733 ( .A(x[836]), .B(n6895), .Z(n6897) );
  XOR U7734 ( .A(n6898), .B(n6899), .Z(n6895) );
  AND U7735 ( .A(n6900), .B(n6901), .Z(n6898) );
  XNOR U7736 ( .A(x[835]), .B(n6899), .Z(n6901) );
  XOR U7737 ( .A(n6902), .B(n6903), .Z(n6899) );
  AND U7738 ( .A(n6904), .B(n6905), .Z(n6902) );
  XNOR U7739 ( .A(x[834]), .B(n6903), .Z(n6905) );
  XOR U7740 ( .A(n6906), .B(n6907), .Z(n6903) );
  AND U7741 ( .A(n6908), .B(n6909), .Z(n6906) );
  XNOR U7742 ( .A(x[833]), .B(n6907), .Z(n6909) );
  XOR U7743 ( .A(n6910), .B(n6911), .Z(n6907) );
  AND U7744 ( .A(n6912), .B(n6913), .Z(n6910) );
  XNOR U7745 ( .A(x[832]), .B(n6911), .Z(n6913) );
  XOR U7746 ( .A(n6914), .B(n6915), .Z(n6911) );
  AND U7747 ( .A(n6916), .B(n6917), .Z(n6914) );
  XNOR U7748 ( .A(x[831]), .B(n6915), .Z(n6917) );
  XOR U7749 ( .A(n6918), .B(n6919), .Z(n6915) );
  AND U7750 ( .A(n6920), .B(n6921), .Z(n6918) );
  XNOR U7751 ( .A(x[830]), .B(n6919), .Z(n6921) );
  XOR U7752 ( .A(n6922), .B(n6923), .Z(n6919) );
  AND U7753 ( .A(n6924), .B(n6925), .Z(n6922) );
  XNOR U7754 ( .A(x[829]), .B(n6923), .Z(n6925) );
  XOR U7755 ( .A(n6926), .B(n6927), .Z(n6923) );
  AND U7756 ( .A(n6928), .B(n6929), .Z(n6926) );
  XNOR U7757 ( .A(x[828]), .B(n6927), .Z(n6929) );
  XOR U7758 ( .A(n6930), .B(n6931), .Z(n6927) );
  AND U7759 ( .A(n6932), .B(n6933), .Z(n6930) );
  XNOR U7760 ( .A(x[827]), .B(n6931), .Z(n6933) );
  XOR U7761 ( .A(n6934), .B(n6935), .Z(n6931) );
  AND U7762 ( .A(n6936), .B(n6937), .Z(n6934) );
  XNOR U7763 ( .A(x[826]), .B(n6935), .Z(n6937) );
  XOR U7764 ( .A(n6938), .B(n6939), .Z(n6935) );
  AND U7765 ( .A(n6940), .B(n6941), .Z(n6938) );
  XNOR U7766 ( .A(x[825]), .B(n6939), .Z(n6941) );
  XOR U7767 ( .A(n6942), .B(n6943), .Z(n6939) );
  AND U7768 ( .A(n6944), .B(n6945), .Z(n6942) );
  XNOR U7769 ( .A(x[824]), .B(n6943), .Z(n6945) );
  XOR U7770 ( .A(n6946), .B(n6947), .Z(n6943) );
  AND U7771 ( .A(n6948), .B(n6949), .Z(n6946) );
  XNOR U7772 ( .A(x[823]), .B(n6947), .Z(n6949) );
  XOR U7773 ( .A(n6950), .B(n6951), .Z(n6947) );
  AND U7774 ( .A(n6952), .B(n6953), .Z(n6950) );
  XNOR U7775 ( .A(x[822]), .B(n6951), .Z(n6953) );
  XOR U7776 ( .A(n6954), .B(n6955), .Z(n6951) );
  AND U7777 ( .A(n6956), .B(n6957), .Z(n6954) );
  XNOR U7778 ( .A(x[821]), .B(n6955), .Z(n6957) );
  XOR U7779 ( .A(n6958), .B(n6959), .Z(n6955) );
  AND U7780 ( .A(n6960), .B(n6961), .Z(n6958) );
  XNOR U7781 ( .A(x[820]), .B(n6959), .Z(n6961) );
  XOR U7782 ( .A(n6962), .B(n6963), .Z(n6959) );
  AND U7783 ( .A(n6964), .B(n6965), .Z(n6962) );
  XNOR U7784 ( .A(x[819]), .B(n6963), .Z(n6965) );
  XOR U7785 ( .A(n6966), .B(n6967), .Z(n6963) );
  AND U7786 ( .A(n6968), .B(n6969), .Z(n6966) );
  XNOR U7787 ( .A(x[818]), .B(n6967), .Z(n6969) );
  XOR U7788 ( .A(n6970), .B(n6971), .Z(n6967) );
  AND U7789 ( .A(n6972), .B(n6973), .Z(n6970) );
  XNOR U7790 ( .A(x[817]), .B(n6971), .Z(n6973) );
  XOR U7791 ( .A(n6974), .B(n6975), .Z(n6971) );
  AND U7792 ( .A(n6976), .B(n6977), .Z(n6974) );
  XNOR U7793 ( .A(x[816]), .B(n6975), .Z(n6977) );
  XOR U7794 ( .A(n6978), .B(n6979), .Z(n6975) );
  AND U7795 ( .A(n6980), .B(n6981), .Z(n6978) );
  XNOR U7796 ( .A(x[815]), .B(n6979), .Z(n6981) );
  XOR U7797 ( .A(n6982), .B(n6983), .Z(n6979) );
  AND U7798 ( .A(n6984), .B(n6985), .Z(n6982) );
  XNOR U7799 ( .A(x[814]), .B(n6983), .Z(n6985) );
  XOR U7800 ( .A(n6986), .B(n6987), .Z(n6983) );
  AND U7801 ( .A(n6988), .B(n6989), .Z(n6986) );
  XNOR U7802 ( .A(x[813]), .B(n6987), .Z(n6989) );
  XOR U7803 ( .A(n6990), .B(n6991), .Z(n6987) );
  AND U7804 ( .A(n6992), .B(n6993), .Z(n6990) );
  XNOR U7805 ( .A(x[812]), .B(n6991), .Z(n6993) );
  XOR U7806 ( .A(n6994), .B(n6995), .Z(n6991) );
  AND U7807 ( .A(n6996), .B(n6997), .Z(n6994) );
  XNOR U7808 ( .A(x[811]), .B(n6995), .Z(n6997) );
  XOR U7809 ( .A(n6998), .B(n6999), .Z(n6995) );
  AND U7810 ( .A(n7000), .B(n7001), .Z(n6998) );
  XNOR U7811 ( .A(x[810]), .B(n6999), .Z(n7001) );
  XOR U7812 ( .A(n7002), .B(n7003), .Z(n6999) );
  AND U7813 ( .A(n7004), .B(n7005), .Z(n7002) );
  XNOR U7814 ( .A(x[809]), .B(n7003), .Z(n7005) );
  XOR U7815 ( .A(n7006), .B(n7007), .Z(n7003) );
  AND U7816 ( .A(n7008), .B(n7009), .Z(n7006) );
  XNOR U7817 ( .A(x[808]), .B(n7007), .Z(n7009) );
  XOR U7818 ( .A(n7010), .B(n7011), .Z(n7007) );
  AND U7819 ( .A(n7012), .B(n7013), .Z(n7010) );
  XNOR U7820 ( .A(x[807]), .B(n7011), .Z(n7013) );
  XOR U7821 ( .A(n7014), .B(n7015), .Z(n7011) );
  AND U7822 ( .A(n7016), .B(n7017), .Z(n7014) );
  XNOR U7823 ( .A(x[806]), .B(n7015), .Z(n7017) );
  XOR U7824 ( .A(n7018), .B(n7019), .Z(n7015) );
  AND U7825 ( .A(n7020), .B(n7021), .Z(n7018) );
  XNOR U7826 ( .A(x[805]), .B(n7019), .Z(n7021) );
  XOR U7827 ( .A(n7022), .B(n7023), .Z(n7019) );
  AND U7828 ( .A(n7024), .B(n7025), .Z(n7022) );
  XNOR U7829 ( .A(x[804]), .B(n7023), .Z(n7025) );
  XOR U7830 ( .A(n7026), .B(n7027), .Z(n7023) );
  AND U7831 ( .A(n7028), .B(n7029), .Z(n7026) );
  XNOR U7832 ( .A(x[803]), .B(n7027), .Z(n7029) );
  XOR U7833 ( .A(n7030), .B(n7031), .Z(n7027) );
  AND U7834 ( .A(n7032), .B(n7033), .Z(n7030) );
  XNOR U7835 ( .A(x[802]), .B(n7031), .Z(n7033) );
  XOR U7836 ( .A(n7034), .B(n7035), .Z(n7031) );
  AND U7837 ( .A(n7036), .B(n7037), .Z(n7034) );
  XNOR U7838 ( .A(x[801]), .B(n7035), .Z(n7037) );
  XOR U7839 ( .A(n7038), .B(n7039), .Z(n7035) );
  AND U7840 ( .A(n7040), .B(n7041), .Z(n7038) );
  XNOR U7841 ( .A(x[800]), .B(n7039), .Z(n7041) );
  XOR U7842 ( .A(n7042), .B(n7043), .Z(n7039) );
  AND U7843 ( .A(n7044), .B(n7045), .Z(n7042) );
  XNOR U7844 ( .A(x[799]), .B(n7043), .Z(n7045) );
  XOR U7845 ( .A(n7046), .B(n7047), .Z(n7043) );
  AND U7846 ( .A(n7048), .B(n7049), .Z(n7046) );
  XNOR U7847 ( .A(x[798]), .B(n7047), .Z(n7049) );
  XOR U7848 ( .A(n7050), .B(n7051), .Z(n7047) );
  AND U7849 ( .A(n7052), .B(n7053), .Z(n7050) );
  XNOR U7850 ( .A(x[797]), .B(n7051), .Z(n7053) );
  XOR U7851 ( .A(n7054), .B(n7055), .Z(n7051) );
  AND U7852 ( .A(n7056), .B(n7057), .Z(n7054) );
  XNOR U7853 ( .A(x[796]), .B(n7055), .Z(n7057) );
  XOR U7854 ( .A(n7058), .B(n7059), .Z(n7055) );
  AND U7855 ( .A(n7060), .B(n7061), .Z(n7058) );
  XNOR U7856 ( .A(x[795]), .B(n7059), .Z(n7061) );
  XOR U7857 ( .A(n7062), .B(n7063), .Z(n7059) );
  AND U7858 ( .A(n7064), .B(n7065), .Z(n7062) );
  XNOR U7859 ( .A(x[794]), .B(n7063), .Z(n7065) );
  XOR U7860 ( .A(n7066), .B(n7067), .Z(n7063) );
  AND U7861 ( .A(n7068), .B(n7069), .Z(n7066) );
  XNOR U7862 ( .A(x[793]), .B(n7067), .Z(n7069) );
  XOR U7863 ( .A(n7070), .B(n7071), .Z(n7067) );
  AND U7864 ( .A(n7072), .B(n7073), .Z(n7070) );
  XNOR U7865 ( .A(x[792]), .B(n7071), .Z(n7073) );
  XOR U7866 ( .A(n7074), .B(n7075), .Z(n7071) );
  AND U7867 ( .A(n7076), .B(n7077), .Z(n7074) );
  XNOR U7868 ( .A(x[791]), .B(n7075), .Z(n7077) );
  XOR U7869 ( .A(n7078), .B(n7079), .Z(n7075) );
  AND U7870 ( .A(n7080), .B(n7081), .Z(n7078) );
  XNOR U7871 ( .A(x[790]), .B(n7079), .Z(n7081) );
  XOR U7872 ( .A(n7082), .B(n7083), .Z(n7079) );
  AND U7873 ( .A(n7084), .B(n7085), .Z(n7082) );
  XNOR U7874 ( .A(x[789]), .B(n7083), .Z(n7085) );
  XOR U7875 ( .A(n7086), .B(n7087), .Z(n7083) );
  AND U7876 ( .A(n7088), .B(n7089), .Z(n7086) );
  XNOR U7877 ( .A(x[788]), .B(n7087), .Z(n7089) );
  XOR U7878 ( .A(n7090), .B(n7091), .Z(n7087) );
  AND U7879 ( .A(n7092), .B(n7093), .Z(n7090) );
  XNOR U7880 ( .A(x[787]), .B(n7091), .Z(n7093) );
  XOR U7881 ( .A(n7094), .B(n7095), .Z(n7091) );
  AND U7882 ( .A(n7096), .B(n7097), .Z(n7094) );
  XNOR U7883 ( .A(x[786]), .B(n7095), .Z(n7097) );
  XOR U7884 ( .A(n7098), .B(n7099), .Z(n7095) );
  AND U7885 ( .A(n7100), .B(n7101), .Z(n7098) );
  XNOR U7886 ( .A(x[785]), .B(n7099), .Z(n7101) );
  XOR U7887 ( .A(n7102), .B(n7103), .Z(n7099) );
  AND U7888 ( .A(n7104), .B(n7105), .Z(n7102) );
  XNOR U7889 ( .A(x[784]), .B(n7103), .Z(n7105) );
  XOR U7890 ( .A(n7106), .B(n7107), .Z(n7103) );
  AND U7891 ( .A(n7108), .B(n7109), .Z(n7106) );
  XNOR U7892 ( .A(x[783]), .B(n7107), .Z(n7109) );
  XOR U7893 ( .A(n7110), .B(n7111), .Z(n7107) );
  AND U7894 ( .A(n7112), .B(n7113), .Z(n7110) );
  XNOR U7895 ( .A(x[782]), .B(n7111), .Z(n7113) );
  XOR U7896 ( .A(n7114), .B(n7115), .Z(n7111) );
  AND U7897 ( .A(n7116), .B(n7117), .Z(n7114) );
  XNOR U7898 ( .A(x[781]), .B(n7115), .Z(n7117) );
  XOR U7899 ( .A(n7118), .B(n7119), .Z(n7115) );
  AND U7900 ( .A(n7120), .B(n7121), .Z(n7118) );
  XNOR U7901 ( .A(x[780]), .B(n7119), .Z(n7121) );
  XOR U7902 ( .A(n7122), .B(n7123), .Z(n7119) );
  AND U7903 ( .A(n7124), .B(n7125), .Z(n7122) );
  XNOR U7904 ( .A(x[779]), .B(n7123), .Z(n7125) );
  XOR U7905 ( .A(n7126), .B(n7127), .Z(n7123) );
  AND U7906 ( .A(n7128), .B(n7129), .Z(n7126) );
  XNOR U7907 ( .A(x[778]), .B(n7127), .Z(n7129) );
  XOR U7908 ( .A(n7130), .B(n7131), .Z(n7127) );
  AND U7909 ( .A(n7132), .B(n7133), .Z(n7130) );
  XNOR U7910 ( .A(x[777]), .B(n7131), .Z(n7133) );
  XOR U7911 ( .A(n7134), .B(n7135), .Z(n7131) );
  AND U7912 ( .A(n7136), .B(n7137), .Z(n7134) );
  XNOR U7913 ( .A(x[776]), .B(n7135), .Z(n7137) );
  XOR U7914 ( .A(n7138), .B(n7139), .Z(n7135) );
  AND U7915 ( .A(n7140), .B(n7141), .Z(n7138) );
  XNOR U7916 ( .A(x[775]), .B(n7139), .Z(n7141) );
  XOR U7917 ( .A(n7142), .B(n7143), .Z(n7139) );
  AND U7918 ( .A(n7144), .B(n7145), .Z(n7142) );
  XNOR U7919 ( .A(x[774]), .B(n7143), .Z(n7145) );
  XOR U7920 ( .A(n7146), .B(n7147), .Z(n7143) );
  AND U7921 ( .A(n7148), .B(n7149), .Z(n7146) );
  XNOR U7922 ( .A(x[773]), .B(n7147), .Z(n7149) );
  XOR U7923 ( .A(n7150), .B(n7151), .Z(n7147) );
  AND U7924 ( .A(n7152), .B(n7153), .Z(n7150) );
  XNOR U7925 ( .A(x[772]), .B(n7151), .Z(n7153) );
  XOR U7926 ( .A(n7154), .B(n7155), .Z(n7151) );
  AND U7927 ( .A(n7156), .B(n7157), .Z(n7154) );
  XNOR U7928 ( .A(x[771]), .B(n7155), .Z(n7157) );
  XOR U7929 ( .A(n7158), .B(n7159), .Z(n7155) );
  AND U7930 ( .A(n7160), .B(n7161), .Z(n7158) );
  XNOR U7931 ( .A(x[770]), .B(n7159), .Z(n7161) );
  XOR U7932 ( .A(n7162), .B(n7163), .Z(n7159) );
  AND U7933 ( .A(n7164), .B(n7165), .Z(n7162) );
  XNOR U7934 ( .A(x[769]), .B(n7163), .Z(n7165) );
  XOR U7935 ( .A(n7166), .B(n7167), .Z(n7163) );
  AND U7936 ( .A(n7168), .B(n7169), .Z(n7166) );
  XNOR U7937 ( .A(x[768]), .B(n7167), .Z(n7169) );
  XOR U7938 ( .A(n7170), .B(n7171), .Z(n7167) );
  AND U7939 ( .A(n7172), .B(n7173), .Z(n7170) );
  XNOR U7940 ( .A(x[767]), .B(n7171), .Z(n7173) );
  XOR U7941 ( .A(n7174), .B(n7175), .Z(n7171) );
  AND U7942 ( .A(n7176), .B(n7177), .Z(n7174) );
  XNOR U7943 ( .A(x[766]), .B(n7175), .Z(n7177) );
  XOR U7944 ( .A(n7178), .B(n7179), .Z(n7175) );
  AND U7945 ( .A(n7180), .B(n7181), .Z(n7178) );
  XNOR U7946 ( .A(x[765]), .B(n7179), .Z(n7181) );
  XOR U7947 ( .A(n7182), .B(n7183), .Z(n7179) );
  AND U7948 ( .A(n7184), .B(n7185), .Z(n7182) );
  XNOR U7949 ( .A(x[764]), .B(n7183), .Z(n7185) );
  XOR U7950 ( .A(n7186), .B(n7187), .Z(n7183) );
  AND U7951 ( .A(n7188), .B(n7189), .Z(n7186) );
  XNOR U7952 ( .A(x[763]), .B(n7187), .Z(n7189) );
  XOR U7953 ( .A(n7190), .B(n7191), .Z(n7187) );
  AND U7954 ( .A(n7192), .B(n7193), .Z(n7190) );
  XNOR U7955 ( .A(x[762]), .B(n7191), .Z(n7193) );
  XOR U7956 ( .A(n7194), .B(n7195), .Z(n7191) );
  AND U7957 ( .A(n7196), .B(n7197), .Z(n7194) );
  XNOR U7958 ( .A(x[761]), .B(n7195), .Z(n7197) );
  XOR U7959 ( .A(n7198), .B(n7199), .Z(n7195) );
  AND U7960 ( .A(n7200), .B(n7201), .Z(n7198) );
  XNOR U7961 ( .A(x[760]), .B(n7199), .Z(n7201) );
  XOR U7962 ( .A(n7202), .B(n7203), .Z(n7199) );
  AND U7963 ( .A(n7204), .B(n7205), .Z(n7202) );
  XNOR U7964 ( .A(x[759]), .B(n7203), .Z(n7205) );
  XOR U7965 ( .A(n7206), .B(n7207), .Z(n7203) );
  AND U7966 ( .A(n7208), .B(n7209), .Z(n7206) );
  XNOR U7967 ( .A(x[758]), .B(n7207), .Z(n7209) );
  XOR U7968 ( .A(n7210), .B(n7211), .Z(n7207) );
  AND U7969 ( .A(n7212), .B(n7213), .Z(n7210) );
  XNOR U7970 ( .A(x[757]), .B(n7211), .Z(n7213) );
  XOR U7971 ( .A(n7214), .B(n7215), .Z(n7211) );
  AND U7972 ( .A(n7216), .B(n7217), .Z(n7214) );
  XNOR U7973 ( .A(x[756]), .B(n7215), .Z(n7217) );
  XOR U7974 ( .A(n7218), .B(n7219), .Z(n7215) );
  AND U7975 ( .A(n7220), .B(n7221), .Z(n7218) );
  XNOR U7976 ( .A(x[755]), .B(n7219), .Z(n7221) );
  XOR U7977 ( .A(n7222), .B(n7223), .Z(n7219) );
  AND U7978 ( .A(n7224), .B(n7225), .Z(n7222) );
  XNOR U7979 ( .A(x[754]), .B(n7223), .Z(n7225) );
  XOR U7980 ( .A(n7226), .B(n7227), .Z(n7223) );
  AND U7981 ( .A(n7228), .B(n7229), .Z(n7226) );
  XNOR U7982 ( .A(x[753]), .B(n7227), .Z(n7229) );
  XOR U7983 ( .A(n7230), .B(n7231), .Z(n7227) );
  AND U7984 ( .A(n7232), .B(n7233), .Z(n7230) );
  XNOR U7985 ( .A(x[752]), .B(n7231), .Z(n7233) );
  XOR U7986 ( .A(n7234), .B(n7235), .Z(n7231) );
  AND U7987 ( .A(n7236), .B(n7237), .Z(n7234) );
  XNOR U7988 ( .A(x[751]), .B(n7235), .Z(n7237) );
  XOR U7989 ( .A(n7238), .B(n7239), .Z(n7235) );
  AND U7990 ( .A(n7240), .B(n7241), .Z(n7238) );
  XNOR U7991 ( .A(x[750]), .B(n7239), .Z(n7241) );
  XOR U7992 ( .A(n7242), .B(n7243), .Z(n7239) );
  AND U7993 ( .A(n7244), .B(n7245), .Z(n7242) );
  XNOR U7994 ( .A(x[749]), .B(n7243), .Z(n7245) );
  XOR U7995 ( .A(n7246), .B(n7247), .Z(n7243) );
  AND U7996 ( .A(n7248), .B(n7249), .Z(n7246) );
  XNOR U7997 ( .A(x[748]), .B(n7247), .Z(n7249) );
  XOR U7998 ( .A(n7250), .B(n7251), .Z(n7247) );
  AND U7999 ( .A(n7252), .B(n7253), .Z(n7250) );
  XNOR U8000 ( .A(x[747]), .B(n7251), .Z(n7253) );
  XOR U8001 ( .A(n7254), .B(n7255), .Z(n7251) );
  AND U8002 ( .A(n7256), .B(n7257), .Z(n7254) );
  XNOR U8003 ( .A(x[746]), .B(n7255), .Z(n7257) );
  XOR U8004 ( .A(n7258), .B(n7259), .Z(n7255) );
  AND U8005 ( .A(n7260), .B(n7261), .Z(n7258) );
  XNOR U8006 ( .A(x[745]), .B(n7259), .Z(n7261) );
  XOR U8007 ( .A(n7262), .B(n7263), .Z(n7259) );
  AND U8008 ( .A(n7264), .B(n7265), .Z(n7262) );
  XNOR U8009 ( .A(x[744]), .B(n7263), .Z(n7265) );
  XOR U8010 ( .A(n7266), .B(n7267), .Z(n7263) );
  AND U8011 ( .A(n7268), .B(n7269), .Z(n7266) );
  XNOR U8012 ( .A(x[743]), .B(n7267), .Z(n7269) );
  XOR U8013 ( .A(n7270), .B(n7271), .Z(n7267) );
  AND U8014 ( .A(n7272), .B(n7273), .Z(n7270) );
  XNOR U8015 ( .A(x[742]), .B(n7271), .Z(n7273) );
  XOR U8016 ( .A(n7274), .B(n7275), .Z(n7271) );
  AND U8017 ( .A(n7276), .B(n7277), .Z(n7274) );
  XNOR U8018 ( .A(x[741]), .B(n7275), .Z(n7277) );
  XOR U8019 ( .A(n7278), .B(n7279), .Z(n7275) );
  AND U8020 ( .A(n7280), .B(n7281), .Z(n7278) );
  XNOR U8021 ( .A(x[740]), .B(n7279), .Z(n7281) );
  XOR U8022 ( .A(n7282), .B(n7283), .Z(n7279) );
  AND U8023 ( .A(n7284), .B(n7285), .Z(n7282) );
  XNOR U8024 ( .A(x[739]), .B(n7283), .Z(n7285) );
  XOR U8025 ( .A(n7286), .B(n7287), .Z(n7283) );
  AND U8026 ( .A(n7288), .B(n7289), .Z(n7286) );
  XNOR U8027 ( .A(x[738]), .B(n7287), .Z(n7289) );
  XOR U8028 ( .A(n7290), .B(n7291), .Z(n7287) );
  AND U8029 ( .A(n7292), .B(n7293), .Z(n7290) );
  XNOR U8030 ( .A(x[737]), .B(n7291), .Z(n7293) );
  XOR U8031 ( .A(n7294), .B(n7295), .Z(n7291) );
  AND U8032 ( .A(n7296), .B(n7297), .Z(n7294) );
  XNOR U8033 ( .A(x[736]), .B(n7295), .Z(n7297) );
  XOR U8034 ( .A(n7298), .B(n7299), .Z(n7295) );
  AND U8035 ( .A(n7300), .B(n7301), .Z(n7298) );
  XNOR U8036 ( .A(x[735]), .B(n7299), .Z(n7301) );
  XOR U8037 ( .A(n7302), .B(n7303), .Z(n7299) );
  AND U8038 ( .A(n7304), .B(n7305), .Z(n7302) );
  XNOR U8039 ( .A(x[734]), .B(n7303), .Z(n7305) );
  XOR U8040 ( .A(n7306), .B(n7307), .Z(n7303) );
  AND U8041 ( .A(n7308), .B(n7309), .Z(n7306) );
  XNOR U8042 ( .A(x[733]), .B(n7307), .Z(n7309) );
  XOR U8043 ( .A(n7310), .B(n7311), .Z(n7307) );
  AND U8044 ( .A(n7312), .B(n7313), .Z(n7310) );
  XNOR U8045 ( .A(x[732]), .B(n7311), .Z(n7313) );
  XOR U8046 ( .A(n7314), .B(n7315), .Z(n7311) );
  AND U8047 ( .A(n7316), .B(n7317), .Z(n7314) );
  XNOR U8048 ( .A(x[731]), .B(n7315), .Z(n7317) );
  XOR U8049 ( .A(n7318), .B(n7319), .Z(n7315) );
  AND U8050 ( .A(n7320), .B(n7321), .Z(n7318) );
  XNOR U8051 ( .A(x[730]), .B(n7319), .Z(n7321) );
  XOR U8052 ( .A(n7322), .B(n7323), .Z(n7319) );
  AND U8053 ( .A(n7324), .B(n7325), .Z(n7322) );
  XNOR U8054 ( .A(x[729]), .B(n7323), .Z(n7325) );
  XOR U8055 ( .A(n7326), .B(n7327), .Z(n7323) );
  AND U8056 ( .A(n7328), .B(n7329), .Z(n7326) );
  XNOR U8057 ( .A(x[728]), .B(n7327), .Z(n7329) );
  XOR U8058 ( .A(n7330), .B(n7331), .Z(n7327) );
  AND U8059 ( .A(n7332), .B(n7333), .Z(n7330) );
  XNOR U8060 ( .A(x[727]), .B(n7331), .Z(n7333) );
  XOR U8061 ( .A(n7334), .B(n7335), .Z(n7331) );
  AND U8062 ( .A(n7336), .B(n7337), .Z(n7334) );
  XNOR U8063 ( .A(x[726]), .B(n7335), .Z(n7337) );
  XOR U8064 ( .A(n7338), .B(n7339), .Z(n7335) );
  AND U8065 ( .A(n7340), .B(n7341), .Z(n7338) );
  XNOR U8066 ( .A(x[725]), .B(n7339), .Z(n7341) );
  XOR U8067 ( .A(n7342), .B(n7343), .Z(n7339) );
  AND U8068 ( .A(n7344), .B(n7345), .Z(n7342) );
  XNOR U8069 ( .A(x[724]), .B(n7343), .Z(n7345) );
  XOR U8070 ( .A(n7346), .B(n7347), .Z(n7343) );
  AND U8071 ( .A(n7348), .B(n7349), .Z(n7346) );
  XNOR U8072 ( .A(x[723]), .B(n7347), .Z(n7349) );
  XOR U8073 ( .A(n7350), .B(n7351), .Z(n7347) );
  AND U8074 ( .A(n7352), .B(n7353), .Z(n7350) );
  XNOR U8075 ( .A(x[722]), .B(n7351), .Z(n7353) );
  XOR U8076 ( .A(n7354), .B(n7355), .Z(n7351) );
  AND U8077 ( .A(n7356), .B(n7357), .Z(n7354) );
  XNOR U8078 ( .A(x[721]), .B(n7355), .Z(n7357) );
  XOR U8079 ( .A(n7358), .B(n7359), .Z(n7355) );
  AND U8080 ( .A(n7360), .B(n7361), .Z(n7358) );
  XNOR U8081 ( .A(x[720]), .B(n7359), .Z(n7361) );
  XOR U8082 ( .A(n7362), .B(n7363), .Z(n7359) );
  AND U8083 ( .A(n7364), .B(n7365), .Z(n7362) );
  XNOR U8084 ( .A(x[719]), .B(n7363), .Z(n7365) );
  XOR U8085 ( .A(n7366), .B(n7367), .Z(n7363) );
  AND U8086 ( .A(n7368), .B(n7369), .Z(n7366) );
  XNOR U8087 ( .A(x[718]), .B(n7367), .Z(n7369) );
  XOR U8088 ( .A(n7370), .B(n7371), .Z(n7367) );
  AND U8089 ( .A(n7372), .B(n7373), .Z(n7370) );
  XNOR U8090 ( .A(x[717]), .B(n7371), .Z(n7373) );
  XOR U8091 ( .A(n7374), .B(n7375), .Z(n7371) );
  AND U8092 ( .A(n7376), .B(n7377), .Z(n7374) );
  XNOR U8093 ( .A(x[716]), .B(n7375), .Z(n7377) );
  XOR U8094 ( .A(n7378), .B(n7379), .Z(n7375) );
  AND U8095 ( .A(n7380), .B(n7381), .Z(n7378) );
  XNOR U8096 ( .A(x[715]), .B(n7379), .Z(n7381) );
  XOR U8097 ( .A(n7382), .B(n7383), .Z(n7379) );
  AND U8098 ( .A(n7384), .B(n7385), .Z(n7382) );
  XNOR U8099 ( .A(x[714]), .B(n7383), .Z(n7385) );
  XOR U8100 ( .A(n7386), .B(n7387), .Z(n7383) );
  AND U8101 ( .A(n7388), .B(n7389), .Z(n7386) );
  XNOR U8102 ( .A(x[713]), .B(n7387), .Z(n7389) );
  XOR U8103 ( .A(n7390), .B(n7391), .Z(n7387) );
  AND U8104 ( .A(n7392), .B(n7393), .Z(n7390) );
  XNOR U8105 ( .A(x[712]), .B(n7391), .Z(n7393) );
  XOR U8106 ( .A(n7394), .B(n7395), .Z(n7391) );
  AND U8107 ( .A(n7396), .B(n7397), .Z(n7394) );
  XNOR U8108 ( .A(x[711]), .B(n7395), .Z(n7397) );
  XOR U8109 ( .A(n7398), .B(n7399), .Z(n7395) );
  AND U8110 ( .A(n7400), .B(n7401), .Z(n7398) );
  XNOR U8111 ( .A(x[710]), .B(n7399), .Z(n7401) );
  XOR U8112 ( .A(n7402), .B(n7403), .Z(n7399) );
  AND U8113 ( .A(n7404), .B(n7405), .Z(n7402) );
  XNOR U8114 ( .A(x[709]), .B(n7403), .Z(n7405) );
  XOR U8115 ( .A(n7406), .B(n7407), .Z(n7403) );
  AND U8116 ( .A(n7408), .B(n7409), .Z(n7406) );
  XNOR U8117 ( .A(x[708]), .B(n7407), .Z(n7409) );
  XOR U8118 ( .A(n7410), .B(n7411), .Z(n7407) );
  AND U8119 ( .A(n7412), .B(n7413), .Z(n7410) );
  XNOR U8120 ( .A(x[707]), .B(n7411), .Z(n7413) );
  XOR U8121 ( .A(n7414), .B(n7415), .Z(n7411) );
  AND U8122 ( .A(n7416), .B(n7417), .Z(n7414) );
  XNOR U8123 ( .A(x[706]), .B(n7415), .Z(n7417) );
  XOR U8124 ( .A(n7418), .B(n7419), .Z(n7415) );
  AND U8125 ( .A(n7420), .B(n7421), .Z(n7418) );
  XNOR U8126 ( .A(x[705]), .B(n7419), .Z(n7421) );
  XOR U8127 ( .A(n7422), .B(n7423), .Z(n7419) );
  AND U8128 ( .A(n7424), .B(n7425), .Z(n7422) );
  XNOR U8129 ( .A(x[704]), .B(n7423), .Z(n7425) );
  XOR U8130 ( .A(n7426), .B(n7427), .Z(n7423) );
  AND U8131 ( .A(n7428), .B(n7429), .Z(n7426) );
  XNOR U8132 ( .A(x[703]), .B(n7427), .Z(n7429) );
  XOR U8133 ( .A(n7430), .B(n7431), .Z(n7427) );
  AND U8134 ( .A(n7432), .B(n7433), .Z(n7430) );
  XNOR U8135 ( .A(x[702]), .B(n7431), .Z(n7433) );
  XOR U8136 ( .A(n7434), .B(n7435), .Z(n7431) );
  AND U8137 ( .A(n7436), .B(n7437), .Z(n7434) );
  XNOR U8138 ( .A(x[701]), .B(n7435), .Z(n7437) );
  XOR U8139 ( .A(n7438), .B(n7439), .Z(n7435) );
  AND U8140 ( .A(n7440), .B(n7441), .Z(n7438) );
  XNOR U8141 ( .A(x[700]), .B(n7439), .Z(n7441) );
  XOR U8142 ( .A(n7442), .B(n7443), .Z(n7439) );
  AND U8143 ( .A(n7444), .B(n7445), .Z(n7442) );
  XNOR U8144 ( .A(x[699]), .B(n7443), .Z(n7445) );
  XOR U8145 ( .A(n7446), .B(n7447), .Z(n7443) );
  AND U8146 ( .A(n7448), .B(n7449), .Z(n7446) );
  XNOR U8147 ( .A(x[698]), .B(n7447), .Z(n7449) );
  XOR U8148 ( .A(n7450), .B(n7451), .Z(n7447) );
  AND U8149 ( .A(n7452), .B(n7453), .Z(n7450) );
  XNOR U8150 ( .A(x[697]), .B(n7451), .Z(n7453) );
  XOR U8151 ( .A(n7454), .B(n7455), .Z(n7451) );
  AND U8152 ( .A(n7456), .B(n7457), .Z(n7454) );
  XNOR U8153 ( .A(x[696]), .B(n7455), .Z(n7457) );
  XOR U8154 ( .A(n7458), .B(n7459), .Z(n7455) );
  AND U8155 ( .A(n7460), .B(n7461), .Z(n7458) );
  XNOR U8156 ( .A(x[695]), .B(n7459), .Z(n7461) );
  XOR U8157 ( .A(n7462), .B(n7463), .Z(n7459) );
  AND U8158 ( .A(n7464), .B(n7465), .Z(n7462) );
  XNOR U8159 ( .A(x[694]), .B(n7463), .Z(n7465) );
  XOR U8160 ( .A(n7466), .B(n7467), .Z(n7463) );
  AND U8161 ( .A(n7468), .B(n7469), .Z(n7466) );
  XNOR U8162 ( .A(x[693]), .B(n7467), .Z(n7469) );
  XOR U8163 ( .A(n7470), .B(n7471), .Z(n7467) );
  AND U8164 ( .A(n7472), .B(n7473), .Z(n7470) );
  XNOR U8165 ( .A(x[692]), .B(n7471), .Z(n7473) );
  XOR U8166 ( .A(n7474), .B(n7475), .Z(n7471) );
  AND U8167 ( .A(n7476), .B(n7477), .Z(n7474) );
  XNOR U8168 ( .A(x[691]), .B(n7475), .Z(n7477) );
  XOR U8169 ( .A(n7478), .B(n7479), .Z(n7475) );
  AND U8170 ( .A(n7480), .B(n7481), .Z(n7478) );
  XNOR U8171 ( .A(x[690]), .B(n7479), .Z(n7481) );
  XOR U8172 ( .A(n7482), .B(n7483), .Z(n7479) );
  AND U8173 ( .A(n7484), .B(n7485), .Z(n7482) );
  XNOR U8174 ( .A(x[689]), .B(n7483), .Z(n7485) );
  XOR U8175 ( .A(n7486), .B(n7487), .Z(n7483) );
  AND U8176 ( .A(n7488), .B(n7489), .Z(n7486) );
  XNOR U8177 ( .A(x[688]), .B(n7487), .Z(n7489) );
  XOR U8178 ( .A(n7490), .B(n7491), .Z(n7487) );
  AND U8179 ( .A(n7492), .B(n7493), .Z(n7490) );
  XNOR U8180 ( .A(x[687]), .B(n7491), .Z(n7493) );
  XOR U8181 ( .A(n7494), .B(n7495), .Z(n7491) );
  AND U8182 ( .A(n7496), .B(n7497), .Z(n7494) );
  XNOR U8183 ( .A(x[686]), .B(n7495), .Z(n7497) );
  XOR U8184 ( .A(n7498), .B(n7499), .Z(n7495) );
  AND U8185 ( .A(n7500), .B(n7501), .Z(n7498) );
  XNOR U8186 ( .A(x[685]), .B(n7499), .Z(n7501) );
  XOR U8187 ( .A(n7502), .B(n7503), .Z(n7499) );
  AND U8188 ( .A(n7504), .B(n7505), .Z(n7502) );
  XNOR U8189 ( .A(x[684]), .B(n7503), .Z(n7505) );
  XOR U8190 ( .A(n7506), .B(n7507), .Z(n7503) );
  AND U8191 ( .A(n7508), .B(n7509), .Z(n7506) );
  XNOR U8192 ( .A(x[683]), .B(n7507), .Z(n7509) );
  XOR U8193 ( .A(n7510), .B(n7511), .Z(n7507) );
  AND U8194 ( .A(n7512), .B(n7513), .Z(n7510) );
  XNOR U8195 ( .A(x[682]), .B(n7511), .Z(n7513) );
  XOR U8196 ( .A(n7514), .B(n7515), .Z(n7511) );
  AND U8197 ( .A(n7516), .B(n7517), .Z(n7514) );
  XNOR U8198 ( .A(x[681]), .B(n7515), .Z(n7517) );
  XOR U8199 ( .A(n7518), .B(n7519), .Z(n7515) );
  AND U8200 ( .A(n7520), .B(n7521), .Z(n7518) );
  XNOR U8201 ( .A(x[680]), .B(n7519), .Z(n7521) );
  XOR U8202 ( .A(n7522), .B(n7523), .Z(n7519) );
  AND U8203 ( .A(n7524), .B(n7525), .Z(n7522) );
  XNOR U8204 ( .A(x[679]), .B(n7523), .Z(n7525) );
  XOR U8205 ( .A(n7526), .B(n7527), .Z(n7523) );
  AND U8206 ( .A(n7528), .B(n7529), .Z(n7526) );
  XNOR U8207 ( .A(x[678]), .B(n7527), .Z(n7529) );
  XOR U8208 ( .A(n7530), .B(n7531), .Z(n7527) );
  AND U8209 ( .A(n7532), .B(n7533), .Z(n7530) );
  XNOR U8210 ( .A(x[677]), .B(n7531), .Z(n7533) );
  XOR U8211 ( .A(n7534), .B(n7535), .Z(n7531) );
  AND U8212 ( .A(n7536), .B(n7537), .Z(n7534) );
  XNOR U8213 ( .A(x[676]), .B(n7535), .Z(n7537) );
  XOR U8214 ( .A(n7538), .B(n7539), .Z(n7535) );
  AND U8215 ( .A(n7540), .B(n7541), .Z(n7538) );
  XNOR U8216 ( .A(x[675]), .B(n7539), .Z(n7541) );
  XOR U8217 ( .A(n7542), .B(n7543), .Z(n7539) );
  AND U8218 ( .A(n7544), .B(n7545), .Z(n7542) );
  XNOR U8219 ( .A(x[674]), .B(n7543), .Z(n7545) );
  XOR U8220 ( .A(n7546), .B(n7547), .Z(n7543) );
  AND U8221 ( .A(n7548), .B(n7549), .Z(n7546) );
  XNOR U8222 ( .A(x[673]), .B(n7547), .Z(n7549) );
  XOR U8223 ( .A(n7550), .B(n7551), .Z(n7547) );
  AND U8224 ( .A(n7552), .B(n7553), .Z(n7550) );
  XNOR U8225 ( .A(x[672]), .B(n7551), .Z(n7553) );
  XOR U8226 ( .A(n7554), .B(n7555), .Z(n7551) );
  AND U8227 ( .A(n7556), .B(n7557), .Z(n7554) );
  XNOR U8228 ( .A(x[671]), .B(n7555), .Z(n7557) );
  XOR U8229 ( .A(n7558), .B(n7559), .Z(n7555) );
  AND U8230 ( .A(n7560), .B(n7561), .Z(n7558) );
  XNOR U8231 ( .A(x[670]), .B(n7559), .Z(n7561) );
  XOR U8232 ( .A(n7562), .B(n7563), .Z(n7559) );
  AND U8233 ( .A(n7564), .B(n7565), .Z(n7562) );
  XNOR U8234 ( .A(x[669]), .B(n7563), .Z(n7565) );
  XOR U8235 ( .A(n7566), .B(n7567), .Z(n7563) );
  AND U8236 ( .A(n7568), .B(n7569), .Z(n7566) );
  XNOR U8237 ( .A(x[668]), .B(n7567), .Z(n7569) );
  XOR U8238 ( .A(n7570), .B(n7571), .Z(n7567) );
  AND U8239 ( .A(n7572), .B(n7573), .Z(n7570) );
  XNOR U8240 ( .A(x[667]), .B(n7571), .Z(n7573) );
  XOR U8241 ( .A(n7574), .B(n7575), .Z(n7571) );
  AND U8242 ( .A(n7576), .B(n7577), .Z(n7574) );
  XNOR U8243 ( .A(x[666]), .B(n7575), .Z(n7577) );
  XOR U8244 ( .A(n7578), .B(n7579), .Z(n7575) );
  AND U8245 ( .A(n7580), .B(n7581), .Z(n7578) );
  XNOR U8246 ( .A(x[665]), .B(n7579), .Z(n7581) );
  XOR U8247 ( .A(n7582), .B(n7583), .Z(n7579) );
  AND U8248 ( .A(n7584), .B(n7585), .Z(n7582) );
  XNOR U8249 ( .A(x[664]), .B(n7583), .Z(n7585) );
  XOR U8250 ( .A(n7586), .B(n7587), .Z(n7583) );
  AND U8251 ( .A(n7588), .B(n7589), .Z(n7586) );
  XNOR U8252 ( .A(x[663]), .B(n7587), .Z(n7589) );
  XOR U8253 ( .A(n7590), .B(n7591), .Z(n7587) );
  AND U8254 ( .A(n7592), .B(n7593), .Z(n7590) );
  XNOR U8255 ( .A(x[662]), .B(n7591), .Z(n7593) );
  XOR U8256 ( .A(n7594), .B(n7595), .Z(n7591) );
  AND U8257 ( .A(n7596), .B(n7597), .Z(n7594) );
  XNOR U8258 ( .A(x[661]), .B(n7595), .Z(n7597) );
  XOR U8259 ( .A(n7598), .B(n7599), .Z(n7595) );
  AND U8260 ( .A(n7600), .B(n7601), .Z(n7598) );
  XNOR U8261 ( .A(x[660]), .B(n7599), .Z(n7601) );
  XOR U8262 ( .A(n7602), .B(n7603), .Z(n7599) );
  AND U8263 ( .A(n7604), .B(n7605), .Z(n7602) );
  XNOR U8264 ( .A(x[659]), .B(n7603), .Z(n7605) );
  XOR U8265 ( .A(n7606), .B(n7607), .Z(n7603) );
  AND U8266 ( .A(n7608), .B(n7609), .Z(n7606) );
  XNOR U8267 ( .A(x[658]), .B(n7607), .Z(n7609) );
  XOR U8268 ( .A(n7610), .B(n7611), .Z(n7607) );
  AND U8269 ( .A(n7612), .B(n7613), .Z(n7610) );
  XNOR U8270 ( .A(x[657]), .B(n7611), .Z(n7613) );
  XOR U8271 ( .A(n7614), .B(n7615), .Z(n7611) );
  AND U8272 ( .A(n7616), .B(n7617), .Z(n7614) );
  XNOR U8273 ( .A(x[656]), .B(n7615), .Z(n7617) );
  XOR U8274 ( .A(n7618), .B(n7619), .Z(n7615) );
  AND U8275 ( .A(n7620), .B(n7621), .Z(n7618) );
  XNOR U8276 ( .A(x[655]), .B(n7619), .Z(n7621) );
  XOR U8277 ( .A(n7622), .B(n7623), .Z(n7619) );
  AND U8278 ( .A(n7624), .B(n7625), .Z(n7622) );
  XNOR U8279 ( .A(x[654]), .B(n7623), .Z(n7625) );
  XOR U8280 ( .A(n7626), .B(n7627), .Z(n7623) );
  AND U8281 ( .A(n7628), .B(n7629), .Z(n7626) );
  XNOR U8282 ( .A(x[653]), .B(n7627), .Z(n7629) );
  XOR U8283 ( .A(n7630), .B(n7631), .Z(n7627) );
  AND U8284 ( .A(n7632), .B(n7633), .Z(n7630) );
  XNOR U8285 ( .A(x[652]), .B(n7631), .Z(n7633) );
  XOR U8286 ( .A(n7634), .B(n7635), .Z(n7631) );
  AND U8287 ( .A(n7636), .B(n7637), .Z(n7634) );
  XNOR U8288 ( .A(x[651]), .B(n7635), .Z(n7637) );
  XOR U8289 ( .A(n7638), .B(n7639), .Z(n7635) );
  AND U8290 ( .A(n7640), .B(n7641), .Z(n7638) );
  XNOR U8291 ( .A(x[650]), .B(n7639), .Z(n7641) );
  XOR U8292 ( .A(n7642), .B(n7643), .Z(n7639) );
  AND U8293 ( .A(n7644), .B(n7645), .Z(n7642) );
  XNOR U8294 ( .A(x[649]), .B(n7643), .Z(n7645) );
  XOR U8295 ( .A(n7646), .B(n7647), .Z(n7643) );
  AND U8296 ( .A(n7648), .B(n7649), .Z(n7646) );
  XNOR U8297 ( .A(x[648]), .B(n7647), .Z(n7649) );
  XOR U8298 ( .A(n7650), .B(n7651), .Z(n7647) );
  AND U8299 ( .A(n7652), .B(n7653), .Z(n7650) );
  XNOR U8300 ( .A(x[647]), .B(n7651), .Z(n7653) );
  XOR U8301 ( .A(n7654), .B(n7655), .Z(n7651) );
  AND U8302 ( .A(n7656), .B(n7657), .Z(n7654) );
  XNOR U8303 ( .A(x[646]), .B(n7655), .Z(n7657) );
  XOR U8304 ( .A(n7658), .B(n7659), .Z(n7655) );
  AND U8305 ( .A(n7660), .B(n7661), .Z(n7658) );
  XNOR U8306 ( .A(x[645]), .B(n7659), .Z(n7661) );
  XOR U8307 ( .A(n7662), .B(n7663), .Z(n7659) );
  AND U8308 ( .A(n7664), .B(n7665), .Z(n7662) );
  XNOR U8309 ( .A(x[644]), .B(n7663), .Z(n7665) );
  XOR U8310 ( .A(n7666), .B(n7667), .Z(n7663) );
  AND U8311 ( .A(n7668), .B(n7669), .Z(n7666) );
  XNOR U8312 ( .A(x[643]), .B(n7667), .Z(n7669) );
  XOR U8313 ( .A(n7670), .B(n7671), .Z(n7667) );
  AND U8314 ( .A(n7672), .B(n7673), .Z(n7670) );
  XNOR U8315 ( .A(x[642]), .B(n7671), .Z(n7673) );
  XOR U8316 ( .A(n7674), .B(n7675), .Z(n7671) );
  AND U8317 ( .A(n7676), .B(n7677), .Z(n7674) );
  XNOR U8318 ( .A(x[641]), .B(n7675), .Z(n7677) );
  XOR U8319 ( .A(n7678), .B(n7679), .Z(n7675) );
  AND U8320 ( .A(n7680), .B(n7681), .Z(n7678) );
  XNOR U8321 ( .A(x[640]), .B(n7679), .Z(n7681) );
  XOR U8322 ( .A(n7682), .B(n7683), .Z(n7679) );
  AND U8323 ( .A(n7684), .B(n7685), .Z(n7682) );
  XNOR U8324 ( .A(x[639]), .B(n7683), .Z(n7685) );
  XOR U8325 ( .A(n7686), .B(n7687), .Z(n7683) );
  AND U8326 ( .A(n7688), .B(n7689), .Z(n7686) );
  XNOR U8327 ( .A(x[638]), .B(n7687), .Z(n7689) );
  XOR U8328 ( .A(n7690), .B(n7691), .Z(n7687) );
  AND U8329 ( .A(n7692), .B(n7693), .Z(n7690) );
  XNOR U8330 ( .A(x[637]), .B(n7691), .Z(n7693) );
  XOR U8331 ( .A(n7694), .B(n7695), .Z(n7691) );
  AND U8332 ( .A(n7696), .B(n7697), .Z(n7694) );
  XNOR U8333 ( .A(x[636]), .B(n7695), .Z(n7697) );
  XOR U8334 ( .A(n7698), .B(n7699), .Z(n7695) );
  AND U8335 ( .A(n7700), .B(n7701), .Z(n7698) );
  XNOR U8336 ( .A(x[635]), .B(n7699), .Z(n7701) );
  XOR U8337 ( .A(n7702), .B(n7703), .Z(n7699) );
  AND U8338 ( .A(n7704), .B(n7705), .Z(n7702) );
  XNOR U8339 ( .A(x[634]), .B(n7703), .Z(n7705) );
  XOR U8340 ( .A(n7706), .B(n7707), .Z(n7703) );
  AND U8341 ( .A(n7708), .B(n7709), .Z(n7706) );
  XNOR U8342 ( .A(x[633]), .B(n7707), .Z(n7709) );
  XOR U8343 ( .A(n7710), .B(n7711), .Z(n7707) );
  AND U8344 ( .A(n7712), .B(n7713), .Z(n7710) );
  XNOR U8345 ( .A(x[632]), .B(n7711), .Z(n7713) );
  XOR U8346 ( .A(n7714), .B(n7715), .Z(n7711) );
  AND U8347 ( .A(n7716), .B(n7717), .Z(n7714) );
  XNOR U8348 ( .A(x[631]), .B(n7715), .Z(n7717) );
  XOR U8349 ( .A(n7718), .B(n7719), .Z(n7715) );
  AND U8350 ( .A(n7720), .B(n7721), .Z(n7718) );
  XNOR U8351 ( .A(x[630]), .B(n7719), .Z(n7721) );
  XOR U8352 ( .A(n7722), .B(n7723), .Z(n7719) );
  AND U8353 ( .A(n7724), .B(n7725), .Z(n7722) );
  XNOR U8354 ( .A(x[629]), .B(n7723), .Z(n7725) );
  XOR U8355 ( .A(n7726), .B(n7727), .Z(n7723) );
  AND U8356 ( .A(n7728), .B(n7729), .Z(n7726) );
  XNOR U8357 ( .A(x[628]), .B(n7727), .Z(n7729) );
  XOR U8358 ( .A(n7730), .B(n7731), .Z(n7727) );
  AND U8359 ( .A(n7732), .B(n7733), .Z(n7730) );
  XNOR U8360 ( .A(x[627]), .B(n7731), .Z(n7733) );
  XOR U8361 ( .A(n7734), .B(n7735), .Z(n7731) );
  AND U8362 ( .A(n7736), .B(n7737), .Z(n7734) );
  XNOR U8363 ( .A(x[626]), .B(n7735), .Z(n7737) );
  XOR U8364 ( .A(n7738), .B(n7739), .Z(n7735) );
  AND U8365 ( .A(n7740), .B(n7741), .Z(n7738) );
  XNOR U8366 ( .A(x[625]), .B(n7739), .Z(n7741) );
  XOR U8367 ( .A(n7742), .B(n7743), .Z(n7739) );
  AND U8368 ( .A(n7744), .B(n7745), .Z(n7742) );
  XNOR U8369 ( .A(x[624]), .B(n7743), .Z(n7745) );
  XOR U8370 ( .A(n7746), .B(n7747), .Z(n7743) );
  AND U8371 ( .A(n7748), .B(n7749), .Z(n7746) );
  XNOR U8372 ( .A(x[623]), .B(n7747), .Z(n7749) );
  XOR U8373 ( .A(n7750), .B(n7751), .Z(n7747) );
  AND U8374 ( .A(n7752), .B(n7753), .Z(n7750) );
  XNOR U8375 ( .A(x[622]), .B(n7751), .Z(n7753) );
  XOR U8376 ( .A(n7754), .B(n7755), .Z(n7751) );
  AND U8377 ( .A(n7756), .B(n7757), .Z(n7754) );
  XNOR U8378 ( .A(x[621]), .B(n7755), .Z(n7757) );
  XOR U8379 ( .A(n7758), .B(n7759), .Z(n7755) );
  AND U8380 ( .A(n7760), .B(n7761), .Z(n7758) );
  XNOR U8381 ( .A(x[620]), .B(n7759), .Z(n7761) );
  XOR U8382 ( .A(n7762), .B(n7763), .Z(n7759) );
  AND U8383 ( .A(n7764), .B(n7765), .Z(n7762) );
  XNOR U8384 ( .A(x[619]), .B(n7763), .Z(n7765) );
  XOR U8385 ( .A(n7766), .B(n7767), .Z(n7763) );
  AND U8386 ( .A(n7768), .B(n7769), .Z(n7766) );
  XNOR U8387 ( .A(x[618]), .B(n7767), .Z(n7769) );
  XOR U8388 ( .A(n7770), .B(n7771), .Z(n7767) );
  AND U8389 ( .A(n7772), .B(n7773), .Z(n7770) );
  XNOR U8390 ( .A(x[617]), .B(n7771), .Z(n7773) );
  XOR U8391 ( .A(n7774), .B(n7775), .Z(n7771) );
  AND U8392 ( .A(n7776), .B(n7777), .Z(n7774) );
  XNOR U8393 ( .A(x[616]), .B(n7775), .Z(n7777) );
  XOR U8394 ( .A(n7778), .B(n7779), .Z(n7775) );
  AND U8395 ( .A(n7780), .B(n7781), .Z(n7778) );
  XNOR U8396 ( .A(x[615]), .B(n7779), .Z(n7781) );
  XOR U8397 ( .A(n7782), .B(n7783), .Z(n7779) );
  AND U8398 ( .A(n7784), .B(n7785), .Z(n7782) );
  XNOR U8399 ( .A(x[614]), .B(n7783), .Z(n7785) );
  XOR U8400 ( .A(n7786), .B(n7787), .Z(n7783) );
  AND U8401 ( .A(n7788), .B(n7789), .Z(n7786) );
  XNOR U8402 ( .A(x[613]), .B(n7787), .Z(n7789) );
  XOR U8403 ( .A(n7790), .B(n7791), .Z(n7787) );
  AND U8404 ( .A(n7792), .B(n7793), .Z(n7790) );
  XNOR U8405 ( .A(x[612]), .B(n7791), .Z(n7793) );
  XOR U8406 ( .A(n7794), .B(n7795), .Z(n7791) );
  AND U8407 ( .A(n7796), .B(n7797), .Z(n7794) );
  XNOR U8408 ( .A(x[611]), .B(n7795), .Z(n7797) );
  XOR U8409 ( .A(n7798), .B(n7799), .Z(n7795) );
  AND U8410 ( .A(n7800), .B(n7801), .Z(n7798) );
  XNOR U8411 ( .A(x[610]), .B(n7799), .Z(n7801) );
  XOR U8412 ( .A(n7802), .B(n7803), .Z(n7799) );
  AND U8413 ( .A(n7804), .B(n7805), .Z(n7802) );
  XNOR U8414 ( .A(x[609]), .B(n7803), .Z(n7805) );
  XOR U8415 ( .A(n7806), .B(n7807), .Z(n7803) );
  AND U8416 ( .A(n7808), .B(n7809), .Z(n7806) );
  XNOR U8417 ( .A(x[608]), .B(n7807), .Z(n7809) );
  XOR U8418 ( .A(n7810), .B(n7811), .Z(n7807) );
  AND U8419 ( .A(n7812), .B(n7813), .Z(n7810) );
  XNOR U8420 ( .A(x[607]), .B(n7811), .Z(n7813) );
  XOR U8421 ( .A(n7814), .B(n7815), .Z(n7811) );
  AND U8422 ( .A(n7816), .B(n7817), .Z(n7814) );
  XNOR U8423 ( .A(x[606]), .B(n7815), .Z(n7817) );
  XOR U8424 ( .A(n7818), .B(n7819), .Z(n7815) );
  AND U8425 ( .A(n7820), .B(n7821), .Z(n7818) );
  XNOR U8426 ( .A(x[605]), .B(n7819), .Z(n7821) );
  XOR U8427 ( .A(n7822), .B(n7823), .Z(n7819) );
  AND U8428 ( .A(n7824), .B(n7825), .Z(n7822) );
  XNOR U8429 ( .A(x[604]), .B(n7823), .Z(n7825) );
  XOR U8430 ( .A(n7826), .B(n7827), .Z(n7823) );
  AND U8431 ( .A(n7828), .B(n7829), .Z(n7826) );
  XNOR U8432 ( .A(x[603]), .B(n7827), .Z(n7829) );
  XOR U8433 ( .A(n7830), .B(n7831), .Z(n7827) );
  AND U8434 ( .A(n7832), .B(n7833), .Z(n7830) );
  XNOR U8435 ( .A(x[602]), .B(n7831), .Z(n7833) );
  XOR U8436 ( .A(n7834), .B(n7835), .Z(n7831) );
  AND U8437 ( .A(n7836), .B(n7837), .Z(n7834) );
  XNOR U8438 ( .A(x[601]), .B(n7835), .Z(n7837) );
  XOR U8439 ( .A(n7838), .B(n7839), .Z(n7835) );
  AND U8440 ( .A(n7840), .B(n7841), .Z(n7838) );
  XNOR U8441 ( .A(x[600]), .B(n7839), .Z(n7841) );
  XOR U8442 ( .A(n7842), .B(n7843), .Z(n7839) );
  AND U8443 ( .A(n7844), .B(n7845), .Z(n7842) );
  XNOR U8444 ( .A(x[599]), .B(n7843), .Z(n7845) );
  XOR U8445 ( .A(n7846), .B(n7847), .Z(n7843) );
  AND U8446 ( .A(n7848), .B(n7849), .Z(n7846) );
  XNOR U8447 ( .A(x[598]), .B(n7847), .Z(n7849) );
  XOR U8448 ( .A(n7850), .B(n7851), .Z(n7847) );
  AND U8449 ( .A(n7852), .B(n7853), .Z(n7850) );
  XNOR U8450 ( .A(x[597]), .B(n7851), .Z(n7853) );
  XOR U8451 ( .A(n7854), .B(n7855), .Z(n7851) );
  AND U8452 ( .A(n7856), .B(n7857), .Z(n7854) );
  XNOR U8453 ( .A(x[596]), .B(n7855), .Z(n7857) );
  XOR U8454 ( .A(n7858), .B(n7859), .Z(n7855) );
  AND U8455 ( .A(n7860), .B(n7861), .Z(n7858) );
  XNOR U8456 ( .A(x[595]), .B(n7859), .Z(n7861) );
  XOR U8457 ( .A(n7862), .B(n7863), .Z(n7859) );
  AND U8458 ( .A(n7864), .B(n7865), .Z(n7862) );
  XNOR U8459 ( .A(x[594]), .B(n7863), .Z(n7865) );
  XOR U8460 ( .A(n7866), .B(n7867), .Z(n7863) );
  AND U8461 ( .A(n7868), .B(n7869), .Z(n7866) );
  XNOR U8462 ( .A(x[593]), .B(n7867), .Z(n7869) );
  XOR U8463 ( .A(n7870), .B(n7871), .Z(n7867) );
  AND U8464 ( .A(n7872), .B(n7873), .Z(n7870) );
  XNOR U8465 ( .A(x[592]), .B(n7871), .Z(n7873) );
  XOR U8466 ( .A(n7874), .B(n7875), .Z(n7871) );
  AND U8467 ( .A(n7876), .B(n7877), .Z(n7874) );
  XNOR U8468 ( .A(x[591]), .B(n7875), .Z(n7877) );
  XOR U8469 ( .A(n7878), .B(n7879), .Z(n7875) );
  AND U8470 ( .A(n7880), .B(n7881), .Z(n7878) );
  XNOR U8471 ( .A(x[590]), .B(n7879), .Z(n7881) );
  XOR U8472 ( .A(n7882), .B(n7883), .Z(n7879) );
  AND U8473 ( .A(n7884), .B(n7885), .Z(n7882) );
  XNOR U8474 ( .A(x[589]), .B(n7883), .Z(n7885) );
  XOR U8475 ( .A(n7886), .B(n7887), .Z(n7883) );
  AND U8476 ( .A(n7888), .B(n7889), .Z(n7886) );
  XNOR U8477 ( .A(x[588]), .B(n7887), .Z(n7889) );
  XOR U8478 ( .A(n7890), .B(n7891), .Z(n7887) );
  AND U8479 ( .A(n7892), .B(n7893), .Z(n7890) );
  XNOR U8480 ( .A(x[587]), .B(n7891), .Z(n7893) );
  XOR U8481 ( .A(n7894), .B(n7895), .Z(n7891) );
  AND U8482 ( .A(n7896), .B(n7897), .Z(n7894) );
  XNOR U8483 ( .A(x[586]), .B(n7895), .Z(n7897) );
  XOR U8484 ( .A(n7898), .B(n7899), .Z(n7895) );
  AND U8485 ( .A(n7900), .B(n7901), .Z(n7898) );
  XNOR U8486 ( .A(x[585]), .B(n7899), .Z(n7901) );
  XOR U8487 ( .A(n7902), .B(n7903), .Z(n7899) );
  AND U8488 ( .A(n7904), .B(n7905), .Z(n7902) );
  XNOR U8489 ( .A(x[584]), .B(n7903), .Z(n7905) );
  XOR U8490 ( .A(n7906), .B(n7907), .Z(n7903) );
  AND U8491 ( .A(n7908), .B(n7909), .Z(n7906) );
  XNOR U8492 ( .A(x[583]), .B(n7907), .Z(n7909) );
  XOR U8493 ( .A(n7910), .B(n7911), .Z(n7907) );
  AND U8494 ( .A(n7912), .B(n7913), .Z(n7910) );
  XNOR U8495 ( .A(x[582]), .B(n7911), .Z(n7913) );
  XOR U8496 ( .A(n7914), .B(n7915), .Z(n7911) );
  AND U8497 ( .A(n7916), .B(n7917), .Z(n7914) );
  XNOR U8498 ( .A(x[581]), .B(n7915), .Z(n7917) );
  XOR U8499 ( .A(n7918), .B(n7919), .Z(n7915) );
  AND U8500 ( .A(n7920), .B(n7921), .Z(n7918) );
  XNOR U8501 ( .A(x[580]), .B(n7919), .Z(n7921) );
  XOR U8502 ( .A(n7922), .B(n7923), .Z(n7919) );
  AND U8503 ( .A(n7924), .B(n7925), .Z(n7922) );
  XNOR U8504 ( .A(x[579]), .B(n7923), .Z(n7925) );
  XOR U8505 ( .A(n7926), .B(n7927), .Z(n7923) );
  AND U8506 ( .A(n7928), .B(n7929), .Z(n7926) );
  XNOR U8507 ( .A(x[578]), .B(n7927), .Z(n7929) );
  XOR U8508 ( .A(n7930), .B(n7931), .Z(n7927) );
  AND U8509 ( .A(n7932), .B(n7933), .Z(n7930) );
  XNOR U8510 ( .A(x[577]), .B(n7931), .Z(n7933) );
  XOR U8511 ( .A(n7934), .B(n7935), .Z(n7931) );
  AND U8512 ( .A(n7936), .B(n7937), .Z(n7934) );
  XNOR U8513 ( .A(x[576]), .B(n7935), .Z(n7937) );
  XOR U8514 ( .A(n7938), .B(n7939), .Z(n7935) );
  AND U8515 ( .A(n7940), .B(n7941), .Z(n7938) );
  XNOR U8516 ( .A(x[575]), .B(n7939), .Z(n7941) );
  XOR U8517 ( .A(n7942), .B(n7943), .Z(n7939) );
  AND U8518 ( .A(n7944), .B(n7945), .Z(n7942) );
  XNOR U8519 ( .A(x[574]), .B(n7943), .Z(n7945) );
  XOR U8520 ( .A(n7946), .B(n7947), .Z(n7943) );
  AND U8521 ( .A(n7948), .B(n7949), .Z(n7946) );
  XNOR U8522 ( .A(x[573]), .B(n7947), .Z(n7949) );
  XOR U8523 ( .A(n7950), .B(n7951), .Z(n7947) );
  AND U8524 ( .A(n7952), .B(n7953), .Z(n7950) );
  XNOR U8525 ( .A(x[572]), .B(n7951), .Z(n7953) );
  XOR U8526 ( .A(n7954), .B(n7955), .Z(n7951) );
  AND U8527 ( .A(n7956), .B(n7957), .Z(n7954) );
  XNOR U8528 ( .A(x[571]), .B(n7955), .Z(n7957) );
  XOR U8529 ( .A(n7958), .B(n7959), .Z(n7955) );
  AND U8530 ( .A(n7960), .B(n7961), .Z(n7958) );
  XNOR U8531 ( .A(x[570]), .B(n7959), .Z(n7961) );
  XOR U8532 ( .A(n7962), .B(n7963), .Z(n7959) );
  AND U8533 ( .A(n7964), .B(n7965), .Z(n7962) );
  XNOR U8534 ( .A(x[569]), .B(n7963), .Z(n7965) );
  XOR U8535 ( .A(n7966), .B(n7967), .Z(n7963) );
  AND U8536 ( .A(n7968), .B(n7969), .Z(n7966) );
  XNOR U8537 ( .A(x[568]), .B(n7967), .Z(n7969) );
  XOR U8538 ( .A(n7970), .B(n7971), .Z(n7967) );
  AND U8539 ( .A(n7972), .B(n7973), .Z(n7970) );
  XNOR U8540 ( .A(x[567]), .B(n7971), .Z(n7973) );
  XOR U8541 ( .A(n7974), .B(n7975), .Z(n7971) );
  AND U8542 ( .A(n7976), .B(n7977), .Z(n7974) );
  XNOR U8543 ( .A(x[566]), .B(n7975), .Z(n7977) );
  XOR U8544 ( .A(n7978), .B(n7979), .Z(n7975) );
  AND U8545 ( .A(n7980), .B(n7981), .Z(n7978) );
  XNOR U8546 ( .A(x[565]), .B(n7979), .Z(n7981) );
  XOR U8547 ( .A(n7982), .B(n7983), .Z(n7979) );
  AND U8548 ( .A(n7984), .B(n7985), .Z(n7982) );
  XNOR U8549 ( .A(x[564]), .B(n7983), .Z(n7985) );
  XOR U8550 ( .A(n7986), .B(n7987), .Z(n7983) );
  AND U8551 ( .A(n7988), .B(n7989), .Z(n7986) );
  XNOR U8552 ( .A(x[563]), .B(n7987), .Z(n7989) );
  XOR U8553 ( .A(n7990), .B(n7991), .Z(n7987) );
  AND U8554 ( .A(n7992), .B(n7993), .Z(n7990) );
  XNOR U8555 ( .A(x[562]), .B(n7991), .Z(n7993) );
  XOR U8556 ( .A(n7994), .B(n7995), .Z(n7991) );
  AND U8557 ( .A(n7996), .B(n7997), .Z(n7994) );
  XNOR U8558 ( .A(x[561]), .B(n7995), .Z(n7997) );
  XOR U8559 ( .A(n7998), .B(n7999), .Z(n7995) );
  AND U8560 ( .A(n8000), .B(n8001), .Z(n7998) );
  XNOR U8561 ( .A(x[560]), .B(n7999), .Z(n8001) );
  XOR U8562 ( .A(n8002), .B(n8003), .Z(n7999) );
  AND U8563 ( .A(n8004), .B(n8005), .Z(n8002) );
  XNOR U8564 ( .A(x[559]), .B(n8003), .Z(n8005) );
  XOR U8565 ( .A(n8006), .B(n8007), .Z(n8003) );
  AND U8566 ( .A(n8008), .B(n8009), .Z(n8006) );
  XNOR U8567 ( .A(x[558]), .B(n8007), .Z(n8009) );
  XOR U8568 ( .A(n8010), .B(n8011), .Z(n8007) );
  AND U8569 ( .A(n8012), .B(n8013), .Z(n8010) );
  XNOR U8570 ( .A(x[557]), .B(n8011), .Z(n8013) );
  XOR U8571 ( .A(n8014), .B(n8015), .Z(n8011) );
  AND U8572 ( .A(n8016), .B(n8017), .Z(n8014) );
  XNOR U8573 ( .A(x[556]), .B(n8015), .Z(n8017) );
  XOR U8574 ( .A(n8018), .B(n8019), .Z(n8015) );
  AND U8575 ( .A(n8020), .B(n8021), .Z(n8018) );
  XNOR U8576 ( .A(x[555]), .B(n8019), .Z(n8021) );
  XOR U8577 ( .A(n8022), .B(n8023), .Z(n8019) );
  AND U8578 ( .A(n8024), .B(n8025), .Z(n8022) );
  XNOR U8579 ( .A(x[554]), .B(n8023), .Z(n8025) );
  XOR U8580 ( .A(n8026), .B(n8027), .Z(n8023) );
  AND U8581 ( .A(n8028), .B(n8029), .Z(n8026) );
  XNOR U8582 ( .A(x[553]), .B(n8027), .Z(n8029) );
  XOR U8583 ( .A(n8030), .B(n8031), .Z(n8027) );
  AND U8584 ( .A(n8032), .B(n8033), .Z(n8030) );
  XNOR U8585 ( .A(x[552]), .B(n8031), .Z(n8033) );
  XOR U8586 ( .A(n8034), .B(n8035), .Z(n8031) );
  AND U8587 ( .A(n8036), .B(n8037), .Z(n8034) );
  XNOR U8588 ( .A(x[551]), .B(n8035), .Z(n8037) );
  XOR U8589 ( .A(n8038), .B(n8039), .Z(n8035) );
  AND U8590 ( .A(n8040), .B(n8041), .Z(n8038) );
  XNOR U8591 ( .A(x[550]), .B(n8039), .Z(n8041) );
  XOR U8592 ( .A(n8042), .B(n8043), .Z(n8039) );
  AND U8593 ( .A(n8044), .B(n8045), .Z(n8042) );
  XNOR U8594 ( .A(x[549]), .B(n8043), .Z(n8045) );
  XOR U8595 ( .A(n8046), .B(n8047), .Z(n8043) );
  AND U8596 ( .A(n8048), .B(n8049), .Z(n8046) );
  XNOR U8597 ( .A(x[548]), .B(n8047), .Z(n8049) );
  XOR U8598 ( .A(n8050), .B(n8051), .Z(n8047) );
  AND U8599 ( .A(n8052), .B(n8053), .Z(n8050) );
  XNOR U8600 ( .A(x[547]), .B(n8051), .Z(n8053) );
  XOR U8601 ( .A(n8054), .B(n8055), .Z(n8051) );
  AND U8602 ( .A(n8056), .B(n8057), .Z(n8054) );
  XNOR U8603 ( .A(x[546]), .B(n8055), .Z(n8057) );
  XOR U8604 ( .A(n8058), .B(n8059), .Z(n8055) );
  AND U8605 ( .A(n8060), .B(n8061), .Z(n8058) );
  XNOR U8606 ( .A(x[545]), .B(n8059), .Z(n8061) );
  XOR U8607 ( .A(n8062), .B(n8063), .Z(n8059) );
  AND U8608 ( .A(n8064), .B(n8065), .Z(n8062) );
  XNOR U8609 ( .A(x[544]), .B(n8063), .Z(n8065) );
  XOR U8610 ( .A(n8066), .B(n8067), .Z(n8063) );
  AND U8611 ( .A(n8068), .B(n8069), .Z(n8066) );
  XNOR U8612 ( .A(x[543]), .B(n8067), .Z(n8069) );
  XOR U8613 ( .A(n8070), .B(n8071), .Z(n8067) );
  AND U8614 ( .A(n8072), .B(n8073), .Z(n8070) );
  XNOR U8615 ( .A(x[542]), .B(n8071), .Z(n8073) );
  XOR U8616 ( .A(n8074), .B(n8075), .Z(n8071) );
  AND U8617 ( .A(n8076), .B(n8077), .Z(n8074) );
  XNOR U8618 ( .A(x[541]), .B(n8075), .Z(n8077) );
  XOR U8619 ( .A(n8078), .B(n8079), .Z(n8075) );
  AND U8620 ( .A(n8080), .B(n8081), .Z(n8078) );
  XNOR U8621 ( .A(x[540]), .B(n8079), .Z(n8081) );
  XOR U8622 ( .A(n8082), .B(n8083), .Z(n8079) );
  AND U8623 ( .A(n8084), .B(n8085), .Z(n8082) );
  XNOR U8624 ( .A(x[539]), .B(n8083), .Z(n8085) );
  XOR U8625 ( .A(n8086), .B(n8087), .Z(n8083) );
  AND U8626 ( .A(n8088), .B(n8089), .Z(n8086) );
  XNOR U8627 ( .A(x[538]), .B(n8087), .Z(n8089) );
  XOR U8628 ( .A(n8090), .B(n8091), .Z(n8087) );
  AND U8629 ( .A(n8092), .B(n8093), .Z(n8090) );
  XNOR U8630 ( .A(x[537]), .B(n8091), .Z(n8093) );
  XOR U8631 ( .A(n8094), .B(n8095), .Z(n8091) );
  AND U8632 ( .A(n8096), .B(n8097), .Z(n8094) );
  XNOR U8633 ( .A(x[536]), .B(n8095), .Z(n8097) );
  XOR U8634 ( .A(n8098), .B(n8099), .Z(n8095) );
  AND U8635 ( .A(n8100), .B(n8101), .Z(n8098) );
  XNOR U8636 ( .A(x[535]), .B(n8099), .Z(n8101) );
  XOR U8637 ( .A(n8102), .B(n8103), .Z(n8099) );
  AND U8638 ( .A(n8104), .B(n8105), .Z(n8102) );
  XNOR U8639 ( .A(x[534]), .B(n8103), .Z(n8105) );
  XOR U8640 ( .A(n8106), .B(n8107), .Z(n8103) );
  AND U8641 ( .A(n8108), .B(n8109), .Z(n8106) );
  XNOR U8642 ( .A(x[533]), .B(n8107), .Z(n8109) );
  XOR U8643 ( .A(n8110), .B(n8111), .Z(n8107) );
  AND U8644 ( .A(n8112), .B(n8113), .Z(n8110) );
  XNOR U8645 ( .A(x[532]), .B(n8111), .Z(n8113) );
  XOR U8646 ( .A(n8114), .B(n8115), .Z(n8111) );
  AND U8647 ( .A(n8116), .B(n8117), .Z(n8114) );
  XNOR U8648 ( .A(x[531]), .B(n8115), .Z(n8117) );
  XOR U8649 ( .A(n8118), .B(n8119), .Z(n8115) );
  AND U8650 ( .A(n8120), .B(n8121), .Z(n8118) );
  XNOR U8651 ( .A(x[530]), .B(n8119), .Z(n8121) );
  XOR U8652 ( .A(n8122), .B(n8123), .Z(n8119) );
  AND U8653 ( .A(n8124), .B(n8125), .Z(n8122) );
  XNOR U8654 ( .A(x[529]), .B(n8123), .Z(n8125) );
  XOR U8655 ( .A(n8126), .B(n8127), .Z(n8123) );
  AND U8656 ( .A(n8128), .B(n8129), .Z(n8126) );
  XNOR U8657 ( .A(x[528]), .B(n8127), .Z(n8129) );
  XOR U8658 ( .A(n8130), .B(n8131), .Z(n8127) );
  AND U8659 ( .A(n8132), .B(n8133), .Z(n8130) );
  XNOR U8660 ( .A(x[527]), .B(n8131), .Z(n8133) );
  XOR U8661 ( .A(n8134), .B(n8135), .Z(n8131) );
  AND U8662 ( .A(n8136), .B(n8137), .Z(n8134) );
  XNOR U8663 ( .A(x[526]), .B(n8135), .Z(n8137) );
  XOR U8664 ( .A(n8138), .B(n8139), .Z(n8135) );
  AND U8665 ( .A(n8140), .B(n8141), .Z(n8138) );
  XNOR U8666 ( .A(x[525]), .B(n8139), .Z(n8141) );
  XOR U8667 ( .A(n8142), .B(n8143), .Z(n8139) );
  AND U8668 ( .A(n8144), .B(n8145), .Z(n8142) );
  XNOR U8669 ( .A(x[524]), .B(n8143), .Z(n8145) );
  XOR U8670 ( .A(n8146), .B(n8147), .Z(n8143) );
  AND U8671 ( .A(n8148), .B(n8149), .Z(n8146) );
  XNOR U8672 ( .A(x[523]), .B(n8147), .Z(n8149) );
  XOR U8673 ( .A(n8150), .B(n8151), .Z(n8147) );
  AND U8674 ( .A(n8152), .B(n8153), .Z(n8150) );
  XNOR U8675 ( .A(x[522]), .B(n8151), .Z(n8153) );
  XOR U8676 ( .A(n8154), .B(n8155), .Z(n8151) );
  AND U8677 ( .A(n8156), .B(n8157), .Z(n8154) );
  XNOR U8678 ( .A(x[521]), .B(n8155), .Z(n8157) );
  XOR U8679 ( .A(n8158), .B(n8159), .Z(n8155) );
  AND U8680 ( .A(n8160), .B(n8161), .Z(n8158) );
  XNOR U8681 ( .A(x[520]), .B(n8159), .Z(n8161) );
  XOR U8682 ( .A(n8162), .B(n8163), .Z(n8159) );
  AND U8683 ( .A(n8164), .B(n8165), .Z(n8162) );
  XNOR U8684 ( .A(x[519]), .B(n8163), .Z(n8165) );
  XOR U8685 ( .A(n8166), .B(n8167), .Z(n8163) );
  AND U8686 ( .A(n8168), .B(n8169), .Z(n8166) );
  XNOR U8687 ( .A(x[518]), .B(n8167), .Z(n8169) );
  XOR U8688 ( .A(n8170), .B(n8171), .Z(n8167) );
  AND U8689 ( .A(n8172), .B(n8173), .Z(n8170) );
  XNOR U8690 ( .A(x[517]), .B(n8171), .Z(n8173) );
  XOR U8691 ( .A(n8174), .B(n8175), .Z(n8171) );
  AND U8692 ( .A(n8176), .B(n8177), .Z(n8174) );
  XNOR U8693 ( .A(x[516]), .B(n8175), .Z(n8177) );
  XOR U8694 ( .A(n8178), .B(n8179), .Z(n8175) );
  AND U8695 ( .A(n8180), .B(n8181), .Z(n8178) );
  XNOR U8696 ( .A(x[515]), .B(n8179), .Z(n8181) );
  XOR U8697 ( .A(n8182), .B(n8183), .Z(n8179) );
  AND U8698 ( .A(n8184), .B(n8185), .Z(n8182) );
  XNOR U8699 ( .A(x[514]), .B(n8183), .Z(n8185) );
  XOR U8700 ( .A(n8186), .B(n8187), .Z(n8183) );
  AND U8701 ( .A(n8188), .B(n8189), .Z(n8186) );
  XNOR U8702 ( .A(x[513]), .B(n8187), .Z(n8189) );
  XOR U8703 ( .A(n8190), .B(n8191), .Z(n8187) );
  AND U8704 ( .A(n8192), .B(n8193), .Z(n8190) );
  XNOR U8705 ( .A(x[512]), .B(n8191), .Z(n8193) );
  XOR U8706 ( .A(n8194), .B(n8195), .Z(n8191) );
  AND U8707 ( .A(n8196), .B(n8197), .Z(n8194) );
  XNOR U8708 ( .A(x[511]), .B(n8195), .Z(n8197) );
  XOR U8709 ( .A(n8198), .B(n8199), .Z(n8195) );
  AND U8710 ( .A(n8200), .B(n8201), .Z(n8198) );
  XNOR U8711 ( .A(x[510]), .B(n8199), .Z(n8201) );
  XOR U8712 ( .A(n8202), .B(n8203), .Z(n8199) );
  AND U8713 ( .A(n8204), .B(n8205), .Z(n8202) );
  XNOR U8714 ( .A(x[509]), .B(n8203), .Z(n8205) );
  XOR U8715 ( .A(n8206), .B(n8207), .Z(n8203) );
  AND U8716 ( .A(n8208), .B(n8209), .Z(n8206) );
  XNOR U8717 ( .A(x[508]), .B(n8207), .Z(n8209) );
  XOR U8718 ( .A(n8210), .B(n8211), .Z(n8207) );
  AND U8719 ( .A(n8212), .B(n8213), .Z(n8210) );
  XNOR U8720 ( .A(x[507]), .B(n8211), .Z(n8213) );
  XOR U8721 ( .A(n8214), .B(n8215), .Z(n8211) );
  AND U8722 ( .A(n8216), .B(n8217), .Z(n8214) );
  XNOR U8723 ( .A(x[506]), .B(n8215), .Z(n8217) );
  XOR U8724 ( .A(n8218), .B(n8219), .Z(n8215) );
  AND U8725 ( .A(n8220), .B(n8221), .Z(n8218) );
  XNOR U8726 ( .A(x[505]), .B(n8219), .Z(n8221) );
  XOR U8727 ( .A(n8222), .B(n8223), .Z(n8219) );
  AND U8728 ( .A(n8224), .B(n8225), .Z(n8222) );
  XNOR U8729 ( .A(x[504]), .B(n8223), .Z(n8225) );
  XOR U8730 ( .A(n8226), .B(n8227), .Z(n8223) );
  AND U8731 ( .A(n8228), .B(n8229), .Z(n8226) );
  XNOR U8732 ( .A(x[503]), .B(n8227), .Z(n8229) );
  XOR U8733 ( .A(n8230), .B(n8231), .Z(n8227) );
  AND U8734 ( .A(n8232), .B(n8233), .Z(n8230) );
  XNOR U8735 ( .A(x[502]), .B(n8231), .Z(n8233) );
  XOR U8736 ( .A(n8234), .B(n8235), .Z(n8231) );
  AND U8737 ( .A(n8236), .B(n8237), .Z(n8234) );
  XNOR U8738 ( .A(x[501]), .B(n8235), .Z(n8237) );
  XOR U8739 ( .A(n8238), .B(n8239), .Z(n8235) );
  AND U8740 ( .A(n8240), .B(n8241), .Z(n8238) );
  XNOR U8741 ( .A(x[500]), .B(n8239), .Z(n8241) );
  XOR U8742 ( .A(n8242), .B(n8243), .Z(n8239) );
  AND U8743 ( .A(n8244), .B(n8245), .Z(n8242) );
  XNOR U8744 ( .A(x[499]), .B(n8243), .Z(n8245) );
  XOR U8745 ( .A(n8246), .B(n8247), .Z(n8243) );
  AND U8746 ( .A(n8248), .B(n8249), .Z(n8246) );
  XNOR U8747 ( .A(x[498]), .B(n8247), .Z(n8249) );
  XOR U8748 ( .A(n8250), .B(n8251), .Z(n8247) );
  AND U8749 ( .A(n8252), .B(n8253), .Z(n8250) );
  XNOR U8750 ( .A(x[497]), .B(n8251), .Z(n8253) );
  XOR U8751 ( .A(n8254), .B(n8255), .Z(n8251) );
  AND U8752 ( .A(n8256), .B(n8257), .Z(n8254) );
  XNOR U8753 ( .A(x[496]), .B(n8255), .Z(n8257) );
  XOR U8754 ( .A(n8258), .B(n8259), .Z(n8255) );
  AND U8755 ( .A(n8260), .B(n8261), .Z(n8258) );
  XNOR U8756 ( .A(x[495]), .B(n8259), .Z(n8261) );
  XOR U8757 ( .A(n8262), .B(n8263), .Z(n8259) );
  AND U8758 ( .A(n8264), .B(n8265), .Z(n8262) );
  XNOR U8759 ( .A(x[494]), .B(n8263), .Z(n8265) );
  XOR U8760 ( .A(n8266), .B(n8267), .Z(n8263) );
  AND U8761 ( .A(n8268), .B(n8269), .Z(n8266) );
  XNOR U8762 ( .A(x[493]), .B(n8267), .Z(n8269) );
  XOR U8763 ( .A(n8270), .B(n8271), .Z(n8267) );
  AND U8764 ( .A(n8272), .B(n8273), .Z(n8270) );
  XNOR U8765 ( .A(x[492]), .B(n8271), .Z(n8273) );
  XOR U8766 ( .A(n8274), .B(n8275), .Z(n8271) );
  AND U8767 ( .A(n8276), .B(n8277), .Z(n8274) );
  XNOR U8768 ( .A(x[491]), .B(n8275), .Z(n8277) );
  XOR U8769 ( .A(n8278), .B(n8279), .Z(n8275) );
  AND U8770 ( .A(n8280), .B(n8281), .Z(n8278) );
  XNOR U8771 ( .A(x[490]), .B(n8279), .Z(n8281) );
  XOR U8772 ( .A(n8282), .B(n8283), .Z(n8279) );
  AND U8773 ( .A(n8284), .B(n8285), .Z(n8282) );
  XNOR U8774 ( .A(x[489]), .B(n8283), .Z(n8285) );
  XOR U8775 ( .A(n8286), .B(n8287), .Z(n8283) );
  AND U8776 ( .A(n8288), .B(n8289), .Z(n8286) );
  XNOR U8777 ( .A(x[488]), .B(n8287), .Z(n8289) );
  XOR U8778 ( .A(n8290), .B(n8291), .Z(n8287) );
  AND U8779 ( .A(n8292), .B(n8293), .Z(n8290) );
  XNOR U8780 ( .A(x[487]), .B(n8291), .Z(n8293) );
  XOR U8781 ( .A(n8294), .B(n8295), .Z(n8291) );
  AND U8782 ( .A(n8296), .B(n8297), .Z(n8294) );
  XNOR U8783 ( .A(x[486]), .B(n8295), .Z(n8297) );
  XOR U8784 ( .A(n8298), .B(n8299), .Z(n8295) );
  AND U8785 ( .A(n8300), .B(n8301), .Z(n8298) );
  XNOR U8786 ( .A(x[485]), .B(n8299), .Z(n8301) );
  XOR U8787 ( .A(n8302), .B(n8303), .Z(n8299) );
  AND U8788 ( .A(n8304), .B(n8305), .Z(n8302) );
  XNOR U8789 ( .A(x[484]), .B(n8303), .Z(n8305) );
  XOR U8790 ( .A(n8306), .B(n8307), .Z(n8303) );
  AND U8791 ( .A(n8308), .B(n8309), .Z(n8306) );
  XNOR U8792 ( .A(x[483]), .B(n8307), .Z(n8309) );
  XOR U8793 ( .A(n8310), .B(n8311), .Z(n8307) );
  AND U8794 ( .A(n8312), .B(n8313), .Z(n8310) );
  XNOR U8795 ( .A(x[482]), .B(n8311), .Z(n8313) );
  XOR U8796 ( .A(n8314), .B(n8315), .Z(n8311) );
  AND U8797 ( .A(n8316), .B(n8317), .Z(n8314) );
  XNOR U8798 ( .A(x[481]), .B(n8315), .Z(n8317) );
  XOR U8799 ( .A(n8318), .B(n8319), .Z(n8315) );
  AND U8800 ( .A(n8320), .B(n8321), .Z(n8318) );
  XNOR U8801 ( .A(x[480]), .B(n8319), .Z(n8321) );
  XOR U8802 ( .A(n8322), .B(n8323), .Z(n8319) );
  AND U8803 ( .A(n8324), .B(n8325), .Z(n8322) );
  XNOR U8804 ( .A(x[479]), .B(n8323), .Z(n8325) );
  XOR U8805 ( .A(n8326), .B(n8327), .Z(n8323) );
  AND U8806 ( .A(n8328), .B(n8329), .Z(n8326) );
  XNOR U8807 ( .A(x[478]), .B(n8327), .Z(n8329) );
  XOR U8808 ( .A(n8330), .B(n8331), .Z(n8327) );
  AND U8809 ( .A(n8332), .B(n8333), .Z(n8330) );
  XNOR U8810 ( .A(x[477]), .B(n8331), .Z(n8333) );
  XOR U8811 ( .A(n8334), .B(n8335), .Z(n8331) );
  AND U8812 ( .A(n8336), .B(n8337), .Z(n8334) );
  XNOR U8813 ( .A(x[476]), .B(n8335), .Z(n8337) );
  XOR U8814 ( .A(n8338), .B(n8339), .Z(n8335) );
  AND U8815 ( .A(n8340), .B(n8341), .Z(n8338) );
  XNOR U8816 ( .A(x[475]), .B(n8339), .Z(n8341) );
  XOR U8817 ( .A(n8342), .B(n8343), .Z(n8339) );
  AND U8818 ( .A(n8344), .B(n8345), .Z(n8342) );
  XNOR U8819 ( .A(x[474]), .B(n8343), .Z(n8345) );
  XOR U8820 ( .A(n8346), .B(n8347), .Z(n8343) );
  AND U8821 ( .A(n8348), .B(n8349), .Z(n8346) );
  XNOR U8822 ( .A(x[473]), .B(n8347), .Z(n8349) );
  XOR U8823 ( .A(n8350), .B(n8351), .Z(n8347) );
  AND U8824 ( .A(n8352), .B(n8353), .Z(n8350) );
  XNOR U8825 ( .A(x[472]), .B(n8351), .Z(n8353) );
  XOR U8826 ( .A(n8354), .B(n8355), .Z(n8351) );
  AND U8827 ( .A(n8356), .B(n8357), .Z(n8354) );
  XNOR U8828 ( .A(x[471]), .B(n8355), .Z(n8357) );
  XOR U8829 ( .A(n8358), .B(n8359), .Z(n8355) );
  AND U8830 ( .A(n8360), .B(n8361), .Z(n8358) );
  XNOR U8831 ( .A(x[470]), .B(n8359), .Z(n8361) );
  XOR U8832 ( .A(n8362), .B(n8363), .Z(n8359) );
  AND U8833 ( .A(n8364), .B(n8365), .Z(n8362) );
  XNOR U8834 ( .A(x[469]), .B(n8363), .Z(n8365) );
  XOR U8835 ( .A(n8366), .B(n8367), .Z(n8363) );
  AND U8836 ( .A(n8368), .B(n8369), .Z(n8366) );
  XNOR U8837 ( .A(x[468]), .B(n8367), .Z(n8369) );
  XOR U8838 ( .A(n8370), .B(n8371), .Z(n8367) );
  AND U8839 ( .A(n8372), .B(n8373), .Z(n8370) );
  XNOR U8840 ( .A(x[467]), .B(n8371), .Z(n8373) );
  XOR U8841 ( .A(n8374), .B(n8375), .Z(n8371) );
  AND U8842 ( .A(n8376), .B(n8377), .Z(n8374) );
  XNOR U8843 ( .A(x[466]), .B(n8375), .Z(n8377) );
  XOR U8844 ( .A(n8378), .B(n8379), .Z(n8375) );
  AND U8845 ( .A(n8380), .B(n8381), .Z(n8378) );
  XNOR U8846 ( .A(x[465]), .B(n8379), .Z(n8381) );
  XOR U8847 ( .A(n8382), .B(n8383), .Z(n8379) );
  AND U8848 ( .A(n8384), .B(n8385), .Z(n8382) );
  XNOR U8849 ( .A(x[464]), .B(n8383), .Z(n8385) );
  XOR U8850 ( .A(n8386), .B(n8387), .Z(n8383) );
  AND U8851 ( .A(n8388), .B(n8389), .Z(n8386) );
  XNOR U8852 ( .A(x[463]), .B(n8387), .Z(n8389) );
  XOR U8853 ( .A(n8390), .B(n8391), .Z(n8387) );
  AND U8854 ( .A(n8392), .B(n8393), .Z(n8390) );
  XNOR U8855 ( .A(x[462]), .B(n8391), .Z(n8393) );
  XOR U8856 ( .A(n8394), .B(n8395), .Z(n8391) );
  AND U8857 ( .A(n8396), .B(n8397), .Z(n8394) );
  XNOR U8858 ( .A(x[461]), .B(n8395), .Z(n8397) );
  XOR U8859 ( .A(n8398), .B(n8399), .Z(n8395) );
  AND U8860 ( .A(n8400), .B(n8401), .Z(n8398) );
  XNOR U8861 ( .A(x[460]), .B(n8399), .Z(n8401) );
  XOR U8862 ( .A(n8402), .B(n8403), .Z(n8399) );
  AND U8863 ( .A(n8404), .B(n8405), .Z(n8402) );
  XNOR U8864 ( .A(x[459]), .B(n8403), .Z(n8405) );
  XOR U8865 ( .A(n8406), .B(n8407), .Z(n8403) );
  AND U8866 ( .A(n8408), .B(n8409), .Z(n8406) );
  XNOR U8867 ( .A(x[458]), .B(n8407), .Z(n8409) );
  XOR U8868 ( .A(n8410), .B(n8411), .Z(n8407) );
  AND U8869 ( .A(n8412), .B(n8413), .Z(n8410) );
  XNOR U8870 ( .A(x[457]), .B(n8411), .Z(n8413) );
  XOR U8871 ( .A(n8414), .B(n8415), .Z(n8411) );
  AND U8872 ( .A(n8416), .B(n8417), .Z(n8414) );
  XNOR U8873 ( .A(x[456]), .B(n8415), .Z(n8417) );
  XOR U8874 ( .A(n8418), .B(n8419), .Z(n8415) );
  AND U8875 ( .A(n8420), .B(n8421), .Z(n8418) );
  XNOR U8876 ( .A(x[455]), .B(n8419), .Z(n8421) );
  XOR U8877 ( .A(n8422), .B(n8423), .Z(n8419) );
  AND U8878 ( .A(n8424), .B(n8425), .Z(n8422) );
  XNOR U8879 ( .A(x[454]), .B(n8423), .Z(n8425) );
  XOR U8880 ( .A(n8426), .B(n8427), .Z(n8423) );
  AND U8881 ( .A(n8428), .B(n8429), .Z(n8426) );
  XNOR U8882 ( .A(x[453]), .B(n8427), .Z(n8429) );
  XOR U8883 ( .A(n8430), .B(n8431), .Z(n8427) );
  AND U8884 ( .A(n8432), .B(n8433), .Z(n8430) );
  XNOR U8885 ( .A(x[452]), .B(n8431), .Z(n8433) );
  XOR U8886 ( .A(n8434), .B(n8435), .Z(n8431) );
  AND U8887 ( .A(n8436), .B(n8437), .Z(n8434) );
  XNOR U8888 ( .A(x[451]), .B(n8435), .Z(n8437) );
  XOR U8889 ( .A(n8438), .B(n8439), .Z(n8435) );
  AND U8890 ( .A(n8440), .B(n8441), .Z(n8438) );
  XNOR U8891 ( .A(x[450]), .B(n8439), .Z(n8441) );
  XOR U8892 ( .A(n8442), .B(n8443), .Z(n8439) );
  AND U8893 ( .A(n8444), .B(n8445), .Z(n8442) );
  XNOR U8894 ( .A(x[449]), .B(n8443), .Z(n8445) );
  XOR U8895 ( .A(n8446), .B(n8447), .Z(n8443) );
  AND U8896 ( .A(n8448), .B(n8449), .Z(n8446) );
  XNOR U8897 ( .A(x[448]), .B(n8447), .Z(n8449) );
  XOR U8898 ( .A(n8450), .B(n8451), .Z(n8447) );
  AND U8899 ( .A(n8452), .B(n8453), .Z(n8450) );
  XNOR U8900 ( .A(x[447]), .B(n8451), .Z(n8453) );
  XOR U8901 ( .A(n8454), .B(n8455), .Z(n8451) );
  AND U8902 ( .A(n8456), .B(n8457), .Z(n8454) );
  XNOR U8903 ( .A(x[446]), .B(n8455), .Z(n8457) );
  XOR U8904 ( .A(n8458), .B(n8459), .Z(n8455) );
  AND U8905 ( .A(n8460), .B(n8461), .Z(n8458) );
  XNOR U8906 ( .A(x[445]), .B(n8459), .Z(n8461) );
  XOR U8907 ( .A(n8462), .B(n8463), .Z(n8459) );
  AND U8908 ( .A(n8464), .B(n8465), .Z(n8462) );
  XNOR U8909 ( .A(x[444]), .B(n8463), .Z(n8465) );
  XOR U8910 ( .A(n8466), .B(n8467), .Z(n8463) );
  AND U8911 ( .A(n8468), .B(n8469), .Z(n8466) );
  XNOR U8912 ( .A(x[443]), .B(n8467), .Z(n8469) );
  XOR U8913 ( .A(n8470), .B(n8471), .Z(n8467) );
  AND U8914 ( .A(n8472), .B(n8473), .Z(n8470) );
  XNOR U8915 ( .A(x[442]), .B(n8471), .Z(n8473) );
  XOR U8916 ( .A(n8474), .B(n8475), .Z(n8471) );
  AND U8917 ( .A(n8476), .B(n8477), .Z(n8474) );
  XNOR U8918 ( .A(x[441]), .B(n8475), .Z(n8477) );
  XOR U8919 ( .A(n8478), .B(n8479), .Z(n8475) );
  AND U8920 ( .A(n8480), .B(n8481), .Z(n8478) );
  XNOR U8921 ( .A(x[440]), .B(n8479), .Z(n8481) );
  XOR U8922 ( .A(n8482), .B(n8483), .Z(n8479) );
  AND U8923 ( .A(n8484), .B(n8485), .Z(n8482) );
  XNOR U8924 ( .A(x[439]), .B(n8483), .Z(n8485) );
  XOR U8925 ( .A(n8486), .B(n8487), .Z(n8483) );
  AND U8926 ( .A(n8488), .B(n8489), .Z(n8486) );
  XNOR U8927 ( .A(x[438]), .B(n8487), .Z(n8489) );
  XOR U8928 ( .A(n8490), .B(n8491), .Z(n8487) );
  AND U8929 ( .A(n8492), .B(n8493), .Z(n8490) );
  XNOR U8930 ( .A(x[437]), .B(n8491), .Z(n8493) );
  XOR U8931 ( .A(n8494), .B(n8495), .Z(n8491) );
  AND U8932 ( .A(n8496), .B(n8497), .Z(n8494) );
  XNOR U8933 ( .A(x[436]), .B(n8495), .Z(n8497) );
  XOR U8934 ( .A(n8498), .B(n8499), .Z(n8495) );
  AND U8935 ( .A(n8500), .B(n8501), .Z(n8498) );
  XNOR U8936 ( .A(x[435]), .B(n8499), .Z(n8501) );
  XOR U8937 ( .A(n8502), .B(n8503), .Z(n8499) );
  AND U8938 ( .A(n8504), .B(n8505), .Z(n8502) );
  XNOR U8939 ( .A(x[434]), .B(n8503), .Z(n8505) );
  XOR U8940 ( .A(n8506), .B(n8507), .Z(n8503) );
  AND U8941 ( .A(n8508), .B(n8509), .Z(n8506) );
  XNOR U8942 ( .A(x[433]), .B(n8507), .Z(n8509) );
  XOR U8943 ( .A(n8510), .B(n8511), .Z(n8507) );
  AND U8944 ( .A(n8512), .B(n8513), .Z(n8510) );
  XNOR U8945 ( .A(x[432]), .B(n8511), .Z(n8513) );
  XOR U8946 ( .A(n8514), .B(n8515), .Z(n8511) );
  AND U8947 ( .A(n8516), .B(n8517), .Z(n8514) );
  XNOR U8948 ( .A(x[431]), .B(n8515), .Z(n8517) );
  XOR U8949 ( .A(n8518), .B(n8519), .Z(n8515) );
  AND U8950 ( .A(n8520), .B(n8521), .Z(n8518) );
  XNOR U8951 ( .A(x[430]), .B(n8519), .Z(n8521) );
  XOR U8952 ( .A(n8522), .B(n8523), .Z(n8519) );
  AND U8953 ( .A(n8524), .B(n8525), .Z(n8522) );
  XNOR U8954 ( .A(x[429]), .B(n8523), .Z(n8525) );
  XOR U8955 ( .A(n8526), .B(n8527), .Z(n8523) );
  AND U8956 ( .A(n8528), .B(n8529), .Z(n8526) );
  XNOR U8957 ( .A(x[428]), .B(n8527), .Z(n8529) );
  XOR U8958 ( .A(n8530), .B(n8531), .Z(n8527) );
  AND U8959 ( .A(n8532), .B(n8533), .Z(n8530) );
  XNOR U8960 ( .A(x[427]), .B(n8531), .Z(n8533) );
  XOR U8961 ( .A(n8534), .B(n8535), .Z(n8531) );
  AND U8962 ( .A(n8536), .B(n8537), .Z(n8534) );
  XNOR U8963 ( .A(x[426]), .B(n8535), .Z(n8537) );
  XOR U8964 ( .A(n8538), .B(n8539), .Z(n8535) );
  AND U8965 ( .A(n8540), .B(n8541), .Z(n8538) );
  XNOR U8966 ( .A(x[425]), .B(n8539), .Z(n8541) );
  XOR U8967 ( .A(n8542), .B(n8543), .Z(n8539) );
  AND U8968 ( .A(n8544), .B(n8545), .Z(n8542) );
  XNOR U8969 ( .A(x[424]), .B(n8543), .Z(n8545) );
  XOR U8970 ( .A(n8546), .B(n8547), .Z(n8543) );
  AND U8971 ( .A(n8548), .B(n8549), .Z(n8546) );
  XNOR U8972 ( .A(x[423]), .B(n8547), .Z(n8549) );
  XOR U8973 ( .A(n8550), .B(n8551), .Z(n8547) );
  AND U8974 ( .A(n8552), .B(n8553), .Z(n8550) );
  XNOR U8975 ( .A(x[422]), .B(n8551), .Z(n8553) );
  XOR U8976 ( .A(n8554), .B(n8555), .Z(n8551) );
  AND U8977 ( .A(n8556), .B(n8557), .Z(n8554) );
  XNOR U8978 ( .A(x[421]), .B(n8555), .Z(n8557) );
  XOR U8979 ( .A(n8558), .B(n8559), .Z(n8555) );
  AND U8980 ( .A(n8560), .B(n8561), .Z(n8558) );
  XNOR U8981 ( .A(x[420]), .B(n8559), .Z(n8561) );
  XOR U8982 ( .A(n8562), .B(n8563), .Z(n8559) );
  AND U8983 ( .A(n8564), .B(n8565), .Z(n8562) );
  XNOR U8984 ( .A(x[419]), .B(n8563), .Z(n8565) );
  XOR U8985 ( .A(n8566), .B(n8567), .Z(n8563) );
  AND U8986 ( .A(n8568), .B(n8569), .Z(n8566) );
  XNOR U8987 ( .A(x[418]), .B(n8567), .Z(n8569) );
  XOR U8988 ( .A(n8570), .B(n8571), .Z(n8567) );
  AND U8989 ( .A(n8572), .B(n8573), .Z(n8570) );
  XNOR U8990 ( .A(x[417]), .B(n8571), .Z(n8573) );
  XOR U8991 ( .A(n8574), .B(n8575), .Z(n8571) );
  AND U8992 ( .A(n8576), .B(n8577), .Z(n8574) );
  XNOR U8993 ( .A(x[416]), .B(n8575), .Z(n8577) );
  XOR U8994 ( .A(n8578), .B(n8579), .Z(n8575) );
  AND U8995 ( .A(n8580), .B(n8581), .Z(n8578) );
  XNOR U8996 ( .A(x[415]), .B(n8579), .Z(n8581) );
  XOR U8997 ( .A(n8582), .B(n8583), .Z(n8579) );
  AND U8998 ( .A(n8584), .B(n8585), .Z(n8582) );
  XNOR U8999 ( .A(x[414]), .B(n8583), .Z(n8585) );
  XOR U9000 ( .A(n8586), .B(n8587), .Z(n8583) );
  AND U9001 ( .A(n8588), .B(n8589), .Z(n8586) );
  XNOR U9002 ( .A(x[413]), .B(n8587), .Z(n8589) );
  XOR U9003 ( .A(n8590), .B(n8591), .Z(n8587) );
  AND U9004 ( .A(n8592), .B(n8593), .Z(n8590) );
  XNOR U9005 ( .A(x[412]), .B(n8591), .Z(n8593) );
  XOR U9006 ( .A(n8594), .B(n8595), .Z(n8591) );
  AND U9007 ( .A(n8596), .B(n8597), .Z(n8594) );
  XNOR U9008 ( .A(x[411]), .B(n8595), .Z(n8597) );
  XOR U9009 ( .A(n8598), .B(n8599), .Z(n8595) );
  AND U9010 ( .A(n8600), .B(n8601), .Z(n8598) );
  XNOR U9011 ( .A(x[410]), .B(n8599), .Z(n8601) );
  XOR U9012 ( .A(n8602), .B(n8603), .Z(n8599) );
  AND U9013 ( .A(n8604), .B(n8605), .Z(n8602) );
  XNOR U9014 ( .A(x[409]), .B(n8603), .Z(n8605) );
  XOR U9015 ( .A(n8606), .B(n8607), .Z(n8603) );
  AND U9016 ( .A(n8608), .B(n8609), .Z(n8606) );
  XNOR U9017 ( .A(x[408]), .B(n8607), .Z(n8609) );
  XOR U9018 ( .A(n8610), .B(n8611), .Z(n8607) );
  AND U9019 ( .A(n8612), .B(n8613), .Z(n8610) );
  XNOR U9020 ( .A(x[407]), .B(n8611), .Z(n8613) );
  XOR U9021 ( .A(n8614), .B(n8615), .Z(n8611) );
  AND U9022 ( .A(n8616), .B(n8617), .Z(n8614) );
  XNOR U9023 ( .A(x[406]), .B(n8615), .Z(n8617) );
  XOR U9024 ( .A(n8618), .B(n8619), .Z(n8615) );
  AND U9025 ( .A(n8620), .B(n8621), .Z(n8618) );
  XNOR U9026 ( .A(x[405]), .B(n8619), .Z(n8621) );
  XOR U9027 ( .A(n8622), .B(n8623), .Z(n8619) );
  AND U9028 ( .A(n8624), .B(n8625), .Z(n8622) );
  XNOR U9029 ( .A(x[404]), .B(n8623), .Z(n8625) );
  XOR U9030 ( .A(n8626), .B(n8627), .Z(n8623) );
  AND U9031 ( .A(n8628), .B(n8629), .Z(n8626) );
  XNOR U9032 ( .A(x[403]), .B(n8627), .Z(n8629) );
  XOR U9033 ( .A(n8630), .B(n8631), .Z(n8627) );
  AND U9034 ( .A(n8632), .B(n8633), .Z(n8630) );
  XNOR U9035 ( .A(x[402]), .B(n8631), .Z(n8633) );
  XOR U9036 ( .A(n8634), .B(n8635), .Z(n8631) );
  AND U9037 ( .A(n8636), .B(n8637), .Z(n8634) );
  XNOR U9038 ( .A(x[401]), .B(n8635), .Z(n8637) );
  XOR U9039 ( .A(n8638), .B(n8639), .Z(n8635) );
  AND U9040 ( .A(n8640), .B(n8641), .Z(n8638) );
  XNOR U9041 ( .A(x[400]), .B(n8639), .Z(n8641) );
  XOR U9042 ( .A(n8642), .B(n8643), .Z(n8639) );
  AND U9043 ( .A(n8644), .B(n8645), .Z(n8642) );
  XNOR U9044 ( .A(x[399]), .B(n8643), .Z(n8645) );
  XOR U9045 ( .A(n8646), .B(n8647), .Z(n8643) );
  AND U9046 ( .A(n8648), .B(n8649), .Z(n8646) );
  XNOR U9047 ( .A(x[398]), .B(n8647), .Z(n8649) );
  XOR U9048 ( .A(n8650), .B(n8651), .Z(n8647) );
  AND U9049 ( .A(n8652), .B(n8653), .Z(n8650) );
  XNOR U9050 ( .A(x[397]), .B(n8651), .Z(n8653) );
  XOR U9051 ( .A(n8654), .B(n8655), .Z(n8651) );
  AND U9052 ( .A(n8656), .B(n8657), .Z(n8654) );
  XNOR U9053 ( .A(x[396]), .B(n8655), .Z(n8657) );
  XOR U9054 ( .A(n8658), .B(n8659), .Z(n8655) );
  AND U9055 ( .A(n8660), .B(n8661), .Z(n8658) );
  XNOR U9056 ( .A(x[395]), .B(n8659), .Z(n8661) );
  XOR U9057 ( .A(n8662), .B(n8663), .Z(n8659) );
  AND U9058 ( .A(n8664), .B(n8665), .Z(n8662) );
  XNOR U9059 ( .A(x[394]), .B(n8663), .Z(n8665) );
  XOR U9060 ( .A(n8666), .B(n8667), .Z(n8663) );
  AND U9061 ( .A(n8668), .B(n8669), .Z(n8666) );
  XNOR U9062 ( .A(x[393]), .B(n8667), .Z(n8669) );
  XOR U9063 ( .A(n8670), .B(n8671), .Z(n8667) );
  AND U9064 ( .A(n8672), .B(n8673), .Z(n8670) );
  XNOR U9065 ( .A(x[392]), .B(n8671), .Z(n8673) );
  XOR U9066 ( .A(n8674), .B(n8675), .Z(n8671) );
  AND U9067 ( .A(n8676), .B(n8677), .Z(n8674) );
  XNOR U9068 ( .A(x[391]), .B(n8675), .Z(n8677) );
  XOR U9069 ( .A(n8678), .B(n8679), .Z(n8675) );
  AND U9070 ( .A(n8680), .B(n8681), .Z(n8678) );
  XNOR U9071 ( .A(x[390]), .B(n8679), .Z(n8681) );
  XOR U9072 ( .A(n8682), .B(n8683), .Z(n8679) );
  AND U9073 ( .A(n8684), .B(n8685), .Z(n8682) );
  XNOR U9074 ( .A(x[389]), .B(n8683), .Z(n8685) );
  XOR U9075 ( .A(n8686), .B(n8687), .Z(n8683) );
  AND U9076 ( .A(n8688), .B(n8689), .Z(n8686) );
  XNOR U9077 ( .A(x[388]), .B(n8687), .Z(n8689) );
  XOR U9078 ( .A(n8690), .B(n8691), .Z(n8687) );
  AND U9079 ( .A(n8692), .B(n8693), .Z(n8690) );
  XNOR U9080 ( .A(x[387]), .B(n8691), .Z(n8693) );
  XOR U9081 ( .A(n8694), .B(n8695), .Z(n8691) );
  AND U9082 ( .A(n8696), .B(n8697), .Z(n8694) );
  XNOR U9083 ( .A(x[386]), .B(n8695), .Z(n8697) );
  XOR U9084 ( .A(n8698), .B(n8699), .Z(n8695) );
  AND U9085 ( .A(n8700), .B(n8701), .Z(n8698) );
  XNOR U9086 ( .A(x[385]), .B(n8699), .Z(n8701) );
  XOR U9087 ( .A(n8702), .B(n8703), .Z(n8699) );
  AND U9088 ( .A(n8704), .B(n8705), .Z(n8702) );
  XNOR U9089 ( .A(x[384]), .B(n8703), .Z(n8705) );
  XOR U9090 ( .A(n8706), .B(n8707), .Z(n8703) );
  AND U9091 ( .A(n8708), .B(n8709), .Z(n8706) );
  XNOR U9092 ( .A(x[383]), .B(n8707), .Z(n8709) );
  XOR U9093 ( .A(n8710), .B(n8711), .Z(n8707) );
  AND U9094 ( .A(n8712), .B(n8713), .Z(n8710) );
  XNOR U9095 ( .A(x[382]), .B(n8711), .Z(n8713) );
  XOR U9096 ( .A(n8714), .B(n8715), .Z(n8711) );
  AND U9097 ( .A(n8716), .B(n8717), .Z(n8714) );
  XNOR U9098 ( .A(x[381]), .B(n8715), .Z(n8717) );
  XOR U9099 ( .A(n8718), .B(n8719), .Z(n8715) );
  AND U9100 ( .A(n8720), .B(n8721), .Z(n8718) );
  XNOR U9101 ( .A(x[380]), .B(n8719), .Z(n8721) );
  XOR U9102 ( .A(n8722), .B(n8723), .Z(n8719) );
  AND U9103 ( .A(n8724), .B(n8725), .Z(n8722) );
  XNOR U9104 ( .A(x[379]), .B(n8723), .Z(n8725) );
  XOR U9105 ( .A(n8726), .B(n8727), .Z(n8723) );
  AND U9106 ( .A(n8728), .B(n8729), .Z(n8726) );
  XNOR U9107 ( .A(x[378]), .B(n8727), .Z(n8729) );
  XOR U9108 ( .A(n8730), .B(n8731), .Z(n8727) );
  AND U9109 ( .A(n8732), .B(n8733), .Z(n8730) );
  XNOR U9110 ( .A(x[377]), .B(n8731), .Z(n8733) );
  XOR U9111 ( .A(n8734), .B(n8735), .Z(n8731) );
  AND U9112 ( .A(n8736), .B(n8737), .Z(n8734) );
  XNOR U9113 ( .A(x[376]), .B(n8735), .Z(n8737) );
  XOR U9114 ( .A(n8738), .B(n8739), .Z(n8735) );
  AND U9115 ( .A(n8740), .B(n8741), .Z(n8738) );
  XNOR U9116 ( .A(x[375]), .B(n8739), .Z(n8741) );
  XOR U9117 ( .A(n8742), .B(n8743), .Z(n8739) );
  AND U9118 ( .A(n8744), .B(n8745), .Z(n8742) );
  XNOR U9119 ( .A(x[374]), .B(n8743), .Z(n8745) );
  XOR U9120 ( .A(n8746), .B(n8747), .Z(n8743) );
  AND U9121 ( .A(n8748), .B(n8749), .Z(n8746) );
  XNOR U9122 ( .A(x[373]), .B(n8747), .Z(n8749) );
  XOR U9123 ( .A(n8750), .B(n8751), .Z(n8747) );
  AND U9124 ( .A(n8752), .B(n8753), .Z(n8750) );
  XNOR U9125 ( .A(x[372]), .B(n8751), .Z(n8753) );
  XOR U9126 ( .A(n8754), .B(n8755), .Z(n8751) );
  AND U9127 ( .A(n8756), .B(n8757), .Z(n8754) );
  XNOR U9128 ( .A(x[371]), .B(n8755), .Z(n8757) );
  XOR U9129 ( .A(n8758), .B(n8759), .Z(n8755) );
  AND U9130 ( .A(n8760), .B(n8761), .Z(n8758) );
  XNOR U9131 ( .A(x[370]), .B(n8759), .Z(n8761) );
  XOR U9132 ( .A(n8762), .B(n8763), .Z(n8759) );
  AND U9133 ( .A(n8764), .B(n8765), .Z(n8762) );
  XNOR U9134 ( .A(x[369]), .B(n8763), .Z(n8765) );
  XOR U9135 ( .A(n8766), .B(n8767), .Z(n8763) );
  AND U9136 ( .A(n8768), .B(n8769), .Z(n8766) );
  XNOR U9137 ( .A(x[368]), .B(n8767), .Z(n8769) );
  XOR U9138 ( .A(n8770), .B(n8771), .Z(n8767) );
  AND U9139 ( .A(n8772), .B(n8773), .Z(n8770) );
  XNOR U9140 ( .A(x[367]), .B(n8771), .Z(n8773) );
  XOR U9141 ( .A(n8774), .B(n8775), .Z(n8771) );
  AND U9142 ( .A(n8776), .B(n8777), .Z(n8774) );
  XNOR U9143 ( .A(x[366]), .B(n8775), .Z(n8777) );
  XOR U9144 ( .A(n8778), .B(n8779), .Z(n8775) );
  AND U9145 ( .A(n8780), .B(n8781), .Z(n8778) );
  XNOR U9146 ( .A(x[365]), .B(n8779), .Z(n8781) );
  XOR U9147 ( .A(n8782), .B(n8783), .Z(n8779) );
  AND U9148 ( .A(n8784), .B(n8785), .Z(n8782) );
  XNOR U9149 ( .A(x[364]), .B(n8783), .Z(n8785) );
  XOR U9150 ( .A(n8786), .B(n8787), .Z(n8783) );
  AND U9151 ( .A(n8788), .B(n8789), .Z(n8786) );
  XNOR U9152 ( .A(x[363]), .B(n8787), .Z(n8789) );
  XOR U9153 ( .A(n8790), .B(n8791), .Z(n8787) );
  AND U9154 ( .A(n8792), .B(n8793), .Z(n8790) );
  XNOR U9155 ( .A(x[362]), .B(n8791), .Z(n8793) );
  XOR U9156 ( .A(n8794), .B(n8795), .Z(n8791) );
  AND U9157 ( .A(n8796), .B(n8797), .Z(n8794) );
  XNOR U9158 ( .A(x[361]), .B(n8795), .Z(n8797) );
  XOR U9159 ( .A(n8798), .B(n8799), .Z(n8795) );
  AND U9160 ( .A(n8800), .B(n8801), .Z(n8798) );
  XNOR U9161 ( .A(x[360]), .B(n8799), .Z(n8801) );
  XOR U9162 ( .A(n8802), .B(n8803), .Z(n8799) );
  AND U9163 ( .A(n8804), .B(n8805), .Z(n8802) );
  XNOR U9164 ( .A(x[359]), .B(n8803), .Z(n8805) );
  XOR U9165 ( .A(n8806), .B(n8807), .Z(n8803) );
  AND U9166 ( .A(n8808), .B(n8809), .Z(n8806) );
  XNOR U9167 ( .A(x[358]), .B(n8807), .Z(n8809) );
  XOR U9168 ( .A(n8810), .B(n8811), .Z(n8807) );
  AND U9169 ( .A(n8812), .B(n8813), .Z(n8810) );
  XNOR U9170 ( .A(x[357]), .B(n8811), .Z(n8813) );
  XOR U9171 ( .A(n8814), .B(n8815), .Z(n8811) );
  AND U9172 ( .A(n8816), .B(n8817), .Z(n8814) );
  XNOR U9173 ( .A(x[356]), .B(n8815), .Z(n8817) );
  XOR U9174 ( .A(n8818), .B(n8819), .Z(n8815) );
  AND U9175 ( .A(n8820), .B(n8821), .Z(n8818) );
  XNOR U9176 ( .A(x[355]), .B(n8819), .Z(n8821) );
  XOR U9177 ( .A(n8822), .B(n8823), .Z(n8819) );
  AND U9178 ( .A(n8824), .B(n8825), .Z(n8822) );
  XNOR U9179 ( .A(x[354]), .B(n8823), .Z(n8825) );
  XOR U9180 ( .A(n8826), .B(n8827), .Z(n8823) );
  AND U9181 ( .A(n8828), .B(n8829), .Z(n8826) );
  XNOR U9182 ( .A(x[353]), .B(n8827), .Z(n8829) );
  XOR U9183 ( .A(n8830), .B(n8831), .Z(n8827) );
  AND U9184 ( .A(n8832), .B(n8833), .Z(n8830) );
  XNOR U9185 ( .A(x[352]), .B(n8831), .Z(n8833) );
  XOR U9186 ( .A(n8834), .B(n8835), .Z(n8831) );
  AND U9187 ( .A(n8836), .B(n8837), .Z(n8834) );
  XNOR U9188 ( .A(x[351]), .B(n8835), .Z(n8837) );
  XOR U9189 ( .A(n8838), .B(n8839), .Z(n8835) );
  AND U9190 ( .A(n8840), .B(n8841), .Z(n8838) );
  XNOR U9191 ( .A(x[350]), .B(n8839), .Z(n8841) );
  XOR U9192 ( .A(n8842), .B(n8843), .Z(n8839) );
  AND U9193 ( .A(n8844), .B(n8845), .Z(n8842) );
  XNOR U9194 ( .A(x[349]), .B(n8843), .Z(n8845) );
  XOR U9195 ( .A(n8846), .B(n8847), .Z(n8843) );
  AND U9196 ( .A(n8848), .B(n8849), .Z(n8846) );
  XNOR U9197 ( .A(x[348]), .B(n8847), .Z(n8849) );
  XOR U9198 ( .A(n8850), .B(n8851), .Z(n8847) );
  AND U9199 ( .A(n8852), .B(n8853), .Z(n8850) );
  XNOR U9200 ( .A(x[347]), .B(n8851), .Z(n8853) );
  XOR U9201 ( .A(n8854), .B(n8855), .Z(n8851) );
  AND U9202 ( .A(n8856), .B(n8857), .Z(n8854) );
  XNOR U9203 ( .A(x[346]), .B(n8855), .Z(n8857) );
  XOR U9204 ( .A(n8858), .B(n8859), .Z(n8855) );
  AND U9205 ( .A(n8860), .B(n8861), .Z(n8858) );
  XNOR U9206 ( .A(x[345]), .B(n8859), .Z(n8861) );
  XOR U9207 ( .A(n8862), .B(n8863), .Z(n8859) );
  AND U9208 ( .A(n8864), .B(n8865), .Z(n8862) );
  XNOR U9209 ( .A(x[344]), .B(n8863), .Z(n8865) );
  XOR U9210 ( .A(n8866), .B(n8867), .Z(n8863) );
  AND U9211 ( .A(n8868), .B(n8869), .Z(n8866) );
  XNOR U9212 ( .A(x[343]), .B(n8867), .Z(n8869) );
  XOR U9213 ( .A(n8870), .B(n8871), .Z(n8867) );
  AND U9214 ( .A(n8872), .B(n8873), .Z(n8870) );
  XNOR U9215 ( .A(x[342]), .B(n8871), .Z(n8873) );
  XOR U9216 ( .A(n8874), .B(n8875), .Z(n8871) );
  AND U9217 ( .A(n8876), .B(n8877), .Z(n8874) );
  XNOR U9218 ( .A(x[341]), .B(n8875), .Z(n8877) );
  XOR U9219 ( .A(n8878), .B(n8879), .Z(n8875) );
  AND U9220 ( .A(n8880), .B(n8881), .Z(n8878) );
  XNOR U9221 ( .A(x[340]), .B(n8879), .Z(n8881) );
  XOR U9222 ( .A(n8882), .B(n8883), .Z(n8879) );
  AND U9223 ( .A(n8884), .B(n8885), .Z(n8882) );
  XNOR U9224 ( .A(x[339]), .B(n8883), .Z(n8885) );
  XOR U9225 ( .A(n8886), .B(n8887), .Z(n8883) );
  AND U9226 ( .A(n8888), .B(n8889), .Z(n8886) );
  XNOR U9227 ( .A(x[338]), .B(n8887), .Z(n8889) );
  XOR U9228 ( .A(n8890), .B(n8891), .Z(n8887) );
  AND U9229 ( .A(n8892), .B(n8893), .Z(n8890) );
  XNOR U9230 ( .A(x[337]), .B(n8891), .Z(n8893) );
  XOR U9231 ( .A(n8894), .B(n8895), .Z(n8891) );
  AND U9232 ( .A(n8896), .B(n8897), .Z(n8894) );
  XNOR U9233 ( .A(x[336]), .B(n8895), .Z(n8897) );
  XOR U9234 ( .A(n8898), .B(n8899), .Z(n8895) );
  AND U9235 ( .A(n8900), .B(n8901), .Z(n8898) );
  XNOR U9236 ( .A(x[335]), .B(n8899), .Z(n8901) );
  XOR U9237 ( .A(n8902), .B(n8903), .Z(n8899) );
  AND U9238 ( .A(n8904), .B(n8905), .Z(n8902) );
  XNOR U9239 ( .A(x[334]), .B(n8903), .Z(n8905) );
  XOR U9240 ( .A(n8906), .B(n8907), .Z(n8903) );
  AND U9241 ( .A(n8908), .B(n8909), .Z(n8906) );
  XNOR U9242 ( .A(x[333]), .B(n8907), .Z(n8909) );
  XOR U9243 ( .A(n8910), .B(n8911), .Z(n8907) );
  AND U9244 ( .A(n8912), .B(n8913), .Z(n8910) );
  XNOR U9245 ( .A(x[332]), .B(n8911), .Z(n8913) );
  XOR U9246 ( .A(n8914), .B(n8915), .Z(n8911) );
  AND U9247 ( .A(n8916), .B(n8917), .Z(n8914) );
  XNOR U9248 ( .A(x[331]), .B(n8915), .Z(n8917) );
  XOR U9249 ( .A(n8918), .B(n8919), .Z(n8915) );
  AND U9250 ( .A(n8920), .B(n8921), .Z(n8918) );
  XNOR U9251 ( .A(x[330]), .B(n8919), .Z(n8921) );
  XOR U9252 ( .A(n8922), .B(n8923), .Z(n8919) );
  AND U9253 ( .A(n8924), .B(n8925), .Z(n8922) );
  XNOR U9254 ( .A(x[329]), .B(n8923), .Z(n8925) );
  XOR U9255 ( .A(n8926), .B(n8927), .Z(n8923) );
  AND U9256 ( .A(n8928), .B(n8929), .Z(n8926) );
  XNOR U9257 ( .A(x[328]), .B(n8927), .Z(n8929) );
  XOR U9258 ( .A(n8930), .B(n8931), .Z(n8927) );
  AND U9259 ( .A(n8932), .B(n8933), .Z(n8930) );
  XNOR U9260 ( .A(x[327]), .B(n8931), .Z(n8933) );
  XOR U9261 ( .A(n8934), .B(n8935), .Z(n8931) );
  AND U9262 ( .A(n8936), .B(n8937), .Z(n8934) );
  XNOR U9263 ( .A(x[326]), .B(n8935), .Z(n8937) );
  XOR U9264 ( .A(n8938), .B(n8939), .Z(n8935) );
  AND U9265 ( .A(n8940), .B(n8941), .Z(n8938) );
  XNOR U9266 ( .A(x[325]), .B(n8939), .Z(n8941) );
  XOR U9267 ( .A(n8942), .B(n8943), .Z(n8939) );
  AND U9268 ( .A(n8944), .B(n8945), .Z(n8942) );
  XNOR U9269 ( .A(x[324]), .B(n8943), .Z(n8945) );
  XOR U9270 ( .A(n8946), .B(n8947), .Z(n8943) );
  AND U9271 ( .A(n8948), .B(n8949), .Z(n8946) );
  XNOR U9272 ( .A(x[323]), .B(n8947), .Z(n8949) );
  XOR U9273 ( .A(n8950), .B(n8951), .Z(n8947) );
  AND U9274 ( .A(n8952), .B(n8953), .Z(n8950) );
  XNOR U9275 ( .A(x[322]), .B(n8951), .Z(n8953) );
  XOR U9276 ( .A(n8954), .B(n8955), .Z(n8951) );
  AND U9277 ( .A(n8956), .B(n8957), .Z(n8954) );
  XNOR U9278 ( .A(x[321]), .B(n8955), .Z(n8957) );
  XOR U9279 ( .A(n8958), .B(n8959), .Z(n8955) );
  AND U9280 ( .A(n8960), .B(n8961), .Z(n8958) );
  XNOR U9281 ( .A(x[320]), .B(n8959), .Z(n8961) );
  XOR U9282 ( .A(n8962), .B(n8963), .Z(n8959) );
  AND U9283 ( .A(n8964), .B(n8965), .Z(n8962) );
  XNOR U9284 ( .A(x[319]), .B(n8963), .Z(n8965) );
  XOR U9285 ( .A(n8966), .B(n8967), .Z(n8963) );
  AND U9286 ( .A(n8968), .B(n8969), .Z(n8966) );
  XNOR U9287 ( .A(x[318]), .B(n8967), .Z(n8969) );
  XOR U9288 ( .A(n8970), .B(n8971), .Z(n8967) );
  AND U9289 ( .A(n8972), .B(n8973), .Z(n8970) );
  XNOR U9290 ( .A(x[317]), .B(n8971), .Z(n8973) );
  XOR U9291 ( .A(n8974), .B(n8975), .Z(n8971) );
  AND U9292 ( .A(n8976), .B(n8977), .Z(n8974) );
  XNOR U9293 ( .A(x[316]), .B(n8975), .Z(n8977) );
  XOR U9294 ( .A(n8978), .B(n8979), .Z(n8975) );
  AND U9295 ( .A(n8980), .B(n8981), .Z(n8978) );
  XNOR U9296 ( .A(x[315]), .B(n8979), .Z(n8981) );
  XOR U9297 ( .A(n8982), .B(n8983), .Z(n8979) );
  AND U9298 ( .A(n8984), .B(n8985), .Z(n8982) );
  XNOR U9299 ( .A(x[314]), .B(n8983), .Z(n8985) );
  XOR U9300 ( .A(n8986), .B(n8987), .Z(n8983) );
  AND U9301 ( .A(n8988), .B(n8989), .Z(n8986) );
  XNOR U9302 ( .A(x[313]), .B(n8987), .Z(n8989) );
  XOR U9303 ( .A(n8990), .B(n8991), .Z(n8987) );
  AND U9304 ( .A(n8992), .B(n8993), .Z(n8990) );
  XNOR U9305 ( .A(x[312]), .B(n8991), .Z(n8993) );
  XOR U9306 ( .A(n8994), .B(n8995), .Z(n8991) );
  AND U9307 ( .A(n8996), .B(n8997), .Z(n8994) );
  XNOR U9308 ( .A(x[311]), .B(n8995), .Z(n8997) );
  XOR U9309 ( .A(n8998), .B(n8999), .Z(n8995) );
  AND U9310 ( .A(n9000), .B(n9001), .Z(n8998) );
  XNOR U9311 ( .A(x[310]), .B(n8999), .Z(n9001) );
  XOR U9312 ( .A(n9002), .B(n9003), .Z(n8999) );
  AND U9313 ( .A(n9004), .B(n9005), .Z(n9002) );
  XNOR U9314 ( .A(x[309]), .B(n9003), .Z(n9005) );
  XOR U9315 ( .A(n9006), .B(n9007), .Z(n9003) );
  AND U9316 ( .A(n9008), .B(n9009), .Z(n9006) );
  XNOR U9317 ( .A(x[308]), .B(n9007), .Z(n9009) );
  XOR U9318 ( .A(n9010), .B(n9011), .Z(n9007) );
  AND U9319 ( .A(n9012), .B(n9013), .Z(n9010) );
  XNOR U9320 ( .A(x[307]), .B(n9011), .Z(n9013) );
  XOR U9321 ( .A(n9014), .B(n9015), .Z(n9011) );
  AND U9322 ( .A(n9016), .B(n9017), .Z(n9014) );
  XNOR U9323 ( .A(x[306]), .B(n9015), .Z(n9017) );
  XOR U9324 ( .A(n9018), .B(n9019), .Z(n9015) );
  AND U9325 ( .A(n9020), .B(n9021), .Z(n9018) );
  XNOR U9326 ( .A(x[305]), .B(n9019), .Z(n9021) );
  XOR U9327 ( .A(n9022), .B(n9023), .Z(n9019) );
  AND U9328 ( .A(n9024), .B(n9025), .Z(n9022) );
  XNOR U9329 ( .A(x[304]), .B(n9023), .Z(n9025) );
  XOR U9330 ( .A(n9026), .B(n9027), .Z(n9023) );
  AND U9331 ( .A(n9028), .B(n9029), .Z(n9026) );
  XNOR U9332 ( .A(x[303]), .B(n9027), .Z(n9029) );
  XOR U9333 ( .A(n9030), .B(n9031), .Z(n9027) );
  AND U9334 ( .A(n9032), .B(n9033), .Z(n9030) );
  XNOR U9335 ( .A(x[302]), .B(n9031), .Z(n9033) );
  XOR U9336 ( .A(n9034), .B(n9035), .Z(n9031) );
  AND U9337 ( .A(n9036), .B(n9037), .Z(n9034) );
  XNOR U9338 ( .A(x[301]), .B(n9035), .Z(n9037) );
  XOR U9339 ( .A(n9038), .B(n9039), .Z(n9035) );
  AND U9340 ( .A(n9040), .B(n9041), .Z(n9038) );
  XNOR U9341 ( .A(x[300]), .B(n9039), .Z(n9041) );
  XOR U9342 ( .A(n9042), .B(n9043), .Z(n9039) );
  AND U9343 ( .A(n9044), .B(n9045), .Z(n9042) );
  XNOR U9344 ( .A(x[299]), .B(n9043), .Z(n9045) );
  XOR U9345 ( .A(n9046), .B(n9047), .Z(n9043) );
  AND U9346 ( .A(n9048), .B(n9049), .Z(n9046) );
  XNOR U9347 ( .A(x[298]), .B(n9047), .Z(n9049) );
  XOR U9348 ( .A(n9050), .B(n9051), .Z(n9047) );
  AND U9349 ( .A(n9052), .B(n9053), .Z(n9050) );
  XNOR U9350 ( .A(x[297]), .B(n9051), .Z(n9053) );
  XOR U9351 ( .A(n9054), .B(n9055), .Z(n9051) );
  AND U9352 ( .A(n9056), .B(n9057), .Z(n9054) );
  XNOR U9353 ( .A(x[296]), .B(n9055), .Z(n9057) );
  XOR U9354 ( .A(n9058), .B(n9059), .Z(n9055) );
  AND U9355 ( .A(n9060), .B(n9061), .Z(n9058) );
  XNOR U9356 ( .A(x[295]), .B(n9059), .Z(n9061) );
  XOR U9357 ( .A(n9062), .B(n9063), .Z(n9059) );
  AND U9358 ( .A(n9064), .B(n9065), .Z(n9062) );
  XNOR U9359 ( .A(x[294]), .B(n9063), .Z(n9065) );
  XOR U9360 ( .A(n9066), .B(n9067), .Z(n9063) );
  AND U9361 ( .A(n9068), .B(n9069), .Z(n9066) );
  XNOR U9362 ( .A(x[293]), .B(n9067), .Z(n9069) );
  XOR U9363 ( .A(n9070), .B(n9071), .Z(n9067) );
  AND U9364 ( .A(n9072), .B(n9073), .Z(n9070) );
  XNOR U9365 ( .A(x[292]), .B(n9071), .Z(n9073) );
  XOR U9366 ( .A(n9074), .B(n9075), .Z(n9071) );
  AND U9367 ( .A(n9076), .B(n9077), .Z(n9074) );
  XNOR U9368 ( .A(x[291]), .B(n9075), .Z(n9077) );
  XOR U9369 ( .A(n9078), .B(n9079), .Z(n9075) );
  AND U9370 ( .A(n9080), .B(n9081), .Z(n9078) );
  XNOR U9371 ( .A(x[290]), .B(n9079), .Z(n9081) );
  XOR U9372 ( .A(n9082), .B(n9083), .Z(n9079) );
  AND U9373 ( .A(n9084), .B(n9085), .Z(n9082) );
  XNOR U9374 ( .A(x[289]), .B(n9083), .Z(n9085) );
  XOR U9375 ( .A(n9086), .B(n9087), .Z(n9083) );
  AND U9376 ( .A(n9088), .B(n9089), .Z(n9086) );
  XNOR U9377 ( .A(x[288]), .B(n9087), .Z(n9089) );
  XOR U9378 ( .A(n9090), .B(n9091), .Z(n9087) );
  AND U9379 ( .A(n9092), .B(n9093), .Z(n9090) );
  XNOR U9380 ( .A(x[287]), .B(n9091), .Z(n9093) );
  XOR U9381 ( .A(n9094), .B(n9095), .Z(n9091) );
  AND U9382 ( .A(n9096), .B(n9097), .Z(n9094) );
  XNOR U9383 ( .A(x[286]), .B(n9095), .Z(n9097) );
  XOR U9384 ( .A(n9098), .B(n9099), .Z(n9095) );
  AND U9385 ( .A(n9100), .B(n9101), .Z(n9098) );
  XNOR U9386 ( .A(x[285]), .B(n9099), .Z(n9101) );
  XOR U9387 ( .A(n9102), .B(n9103), .Z(n9099) );
  AND U9388 ( .A(n9104), .B(n9105), .Z(n9102) );
  XNOR U9389 ( .A(x[284]), .B(n9103), .Z(n9105) );
  XOR U9390 ( .A(n9106), .B(n9107), .Z(n9103) );
  AND U9391 ( .A(n9108), .B(n9109), .Z(n9106) );
  XNOR U9392 ( .A(x[283]), .B(n9107), .Z(n9109) );
  XOR U9393 ( .A(n9110), .B(n9111), .Z(n9107) );
  AND U9394 ( .A(n9112), .B(n9113), .Z(n9110) );
  XNOR U9395 ( .A(x[282]), .B(n9111), .Z(n9113) );
  XOR U9396 ( .A(n9114), .B(n9115), .Z(n9111) );
  AND U9397 ( .A(n9116), .B(n9117), .Z(n9114) );
  XNOR U9398 ( .A(x[281]), .B(n9115), .Z(n9117) );
  XOR U9399 ( .A(n9118), .B(n9119), .Z(n9115) );
  AND U9400 ( .A(n9120), .B(n9121), .Z(n9118) );
  XNOR U9401 ( .A(x[280]), .B(n9119), .Z(n9121) );
  XOR U9402 ( .A(n9122), .B(n9123), .Z(n9119) );
  AND U9403 ( .A(n9124), .B(n9125), .Z(n9122) );
  XNOR U9404 ( .A(x[279]), .B(n9123), .Z(n9125) );
  XOR U9405 ( .A(n9126), .B(n9127), .Z(n9123) );
  AND U9406 ( .A(n9128), .B(n9129), .Z(n9126) );
  XNOR U9407 ( .A(x[278]), .B(n9127), .Z(n9129) );
  XOR U9408 ( .A(n9130), .B(n9131), .Z(n9127) );
  AND U9409 ( .A(n9132), .B(n9133), .Z(n9130) );
  XNOR U9410 ( .A(x[277]), .B(n9131), .Z(n9133) );
  XOR U9411 ( .A(n9134), .B(n9135), .Z(n9131) );
  AND U9412 ( .A(n9136), .B(n9137), .Z(n9134) );
  XNOR U9413 ( .A(x[276]), .B(n9135), .Z(n9137) );
  XOR U9414 ( .A(n9138), .B(n9139), .Z(n9135) );
  AND U9415 ( .A(n9140), .B(n9141), .Z(n9138) );
  XNOR U9416 ( .A(x[275]), .B(n9139), .Z(n9141) );
  XOR U9417 ( .A(n9142), .B(n9143), .Z(n9139) );
  AND U9418 ( .A(n9144), .B(n9145), .Z(n9142) );
  XNOR U9419 ( .A(x[274]), .B(n9143), .Z(n9145) );
  XOR U9420 ( .A(n9146), .B(n9147), .Z(n9143) );
  AND U9421 ( .A(n9148), .B(n9149), .Z(n9146) );
  XNOR U9422 ( .A(x[273]), .B(n9147), .Z(n9149) );
  XOR U9423 ( .A(n9150), .B(n9151), .Z(n9147) );
  AND U9424 ( .A(n9152), .B(n9153), .Z(n9150) );
  XNOR U9425 ( .A(x[272]), .B(n9151), .Z(n9153) );
  XOR U9426 ( .A(n9154), .B(n9155), .Z(n9151) );
  AND U9427 ( .A(n9156), .B(n9157), .Z(n9154) );
  XNOR U9428 ( .A(x[271]), .B(n9155), .Z(n9157) );
  XOR U9429 ( .A(n9158), .B(n9159), .Z(n9155) );
  AND U9430 ( .A(n9160), .B(n9161), .Z(n9158) );
  XNOR U9431 ( .A(x[270]), .B(n9159), .Z(n9161) );
  XOR U9432 ( .A(n9162), .B(n9163), .Z(n9159) );
  AND U9433 ( .A(n9164), .B(n9165), .Z(n9162) );
  XNOR U9434 ( .A(x[269]), .B(n9163), .Z(n9165) );
  XOR U9435 ( .A(n9166), .B(n9167), .Z(n9163) );
  AND U9436 ( .A(n9168), .B(n9169), .Z(n9166) );
  XNOR U9437 ( .A(x[268]), .B(n9167), .Z(n9169) );
  XOR U9438 ( .A(n9170), .B(n9171), .Z(n9167) );
  AND U9439 ( .A(n9172), .B(n9173), .Z(n9170) );
  XNOR U9440 ( .A(x[267]), .B(n9171), .Z(n9173) );
  XOR U9441 ( .A(n9174), .B(n9175), .Z(n9171) );
  AND U9442 ( .A(n9176), .B(n9177), .Z(n9174) );
  XNOR U9443 ( .A(x[266]), .B(n9175), .Z(n9177) );
  XOR U9444 ( .A(n9178), .B(n9179), .Z(n9175) );
  AND U9445 ( .A(n9180), .B(n9181), .Z(n9178) );
  XNOR U9446 ( .A(x[265]), .B(n9179), .Z(n9181) );
  XOR U9447 ( .A(n9182), .B(n9183), .Z(n9179) );
  AND U9448 ( .A(n9184), .B(n9185), .Z(n9182) );
  XNOR U9449 ( .A(x[264]), .B(n9183), .Z(n9185) );
  XOR U9450 ( .A(n9186), .B(n9187), .Z(n9183) );
  AND U9451 ( .A(n9188), .B(n9189), .Z(n9186) );
  XNOR U9452 ( .A(x[263]), .B(n9187), .Z(n9189) );
  XOR U9453 ( .A(n9190), .B(n9191), .Z(n9187) );
  AND U9454 ( .A(n9192), .B(n9193), .Z(n9190) );
  XNOR U9455 ( .A(x[262]), .B(n9191), .Z(n9193) );
  XOR U9456 ( .A(n9194), .B(n9195), .Z(n9191) );
  AND U9457 ( .A(n9196), .B(n9197), .Z(n9194) );
  XNOR U9458 ( .A(x[261]), .B(n9195), .Z(n9197) );
  XOR U9459 ( .A(n9198), .B(n9199), .Z(n9195) );
  AND U9460 ( .A(n9200), .B(n9201), .Z(n9198) );
  XNOR U9461 ( .A(x[260]), .B(n9199), .Z(n9201) );
  XOR U9462 ( .A(n9202), .B(n9203), .Z(n9199) );
  AND U9463 ( .A(n9204), .B(n9205), .Z(n9202) );
  XNOR U9464 ( .A(x[259]), .B(n9203), .Z(n9205) );
  XOR U9465 ( .A(n9206), .B(n9207), .Z(n9203) );
  AND U9466 ( .A(n9208), .B(n9209), .Z(n9206) );
  XNOR U9467 ( .A(x[258]), .B(n9207), .Z(n9209) );
  XOR U9468 ( .A(n9210), .B(n9211), .Z(n9207) );
  AND U9469 ( .A(n9212), .B(n9213), .Z(n9210) );
  XNOR U9470 ( .A(x[257]), .B(n9211), .Z(n9213) );
  XOR U9471 ( .A(n9214), .B(n9215), .Z(n9211) );
  AND U9472 ( .A(n9216), .B(n9217), .Z(n9214) );
  XNOR U9473 ( .A(x[256]), .B(n9215), .Z(n9217) );
  XOR U9474 ( .A(n9218), .B(n9219), .Z(n9215) );
  AND U9475 ( .A(n9220), .B(n9221), .Z(n9218) );
  XNOR U9476 ( .A(x[255]), .B(n9219), .Z(n9221) );
  XOR U9477 ( .A(n9222), .B(n9223), .Z(n9219) );
  AND U9478 ( .A(n9224), .B(n9225), .Z(n9222) );
  XNOR U9479 ( .A(x[254]), .B(n9223), .Z(n9225) );
  XOR U9480 ( .A(n9226), .B(n9227), .Z(n9223) );
  AND U9481 ( .A(n9228), .B(n9229), .Z(n9226) );
  XNOR U9482 ( .A(x[253]), .B(n9227), .Z(n9229) );
  XOR U9483 ( .A(n9230), .B(n9231), .Z(n9227) );
  AND U9484 ( .A(n9232), .B(n9233), .Z(n9230) );
  XNOR U9485 ( .A(x[252]), .B(n9231), .Z(n9233) );
  XOR U9486 ( .A(n9234), .B(n9235), .Z(n9231) );
  AND U9487 ( .A(n9236), .B(n9237), .Z(n9234) );
  XNOR U9488 ( .A(x[251]), .B(n9235), .Z(n9237) );
  XOR U9489 ( .A(n9238), .B(n9239), .Z(n9235) );
  AND U9490 ( .A(n9240), .B(n9241), .Z(n9238) );
  XNOR U9491 ( .A(x[250]), .B(n9239), .Z(n9241) );
  XOR U9492 ( .A(n9242), .B(n9243), .Z(n9239) );
  AND U9493 ( .A(n9244), .B(n9245), .Z(n9242) );
  XNOR U9494 ( .A(x[249]), .B(n9243), .Z(n9245) );
  XOR U9495 ( .A(n9246), .B(n9247), .Z(n9243) );
  AND U9496 ( .A(n9248), .B(n9249), .Z(n9246) );
  XNOR U9497 ( .A(x[248]), .B(n9247), .Z(n9249) );
  XOR U9498 ( .A(n9250), .B(n9251), .Z(n9247) );
  AND U9499 ( .A(n9252), .B(n9253), .Z(n9250) );
  XNOR U9500 ( .A(x[247]), .B(n9251), .Z(n9253) );
  XOR U9501 ( .A(n9254), .B(n9255), .Z(n9251) );
  AND U9502 ( .A(n9256), .B(n9257), .Z(n9254) );
  XNOR U9503 ( .A(x[246]), .B(n9255), .Z(n9257) );
  XOR U9504 ( .A(n9258), .B(n9259), .Z(n9255) );
  AND U9505 ( .A(n9260), .B(n9261), .Z(n9258) );
  XNOR U9506 ( .A(x[245]), .B(n9259), .Z(n9261) );
  XOR U9507 ( .A(n9262), .B(n9263), .Z(n9259) );
  AND U9508 ( .A(n9264), .B(n9265), .Z(n9262) );
  XNOR U9509 ( .A(x[244]), .B(n9263), .Z(n9265) );
  XOR U9510 ( .A(n9266), .B(n9267), .Z(n9263) );
  AND U9511 ( .A(n9268), .B(n9269), .Z(n9266) );
  XNOR U9512 ( .A(x[243]), .B(n9267), .Z(n9269) );
  XOR U9513 ( .A(n9270), .B(n9271), .Z(n9267) );
  AND U9514 ( .A(n9272), .B(n9273), .Z(n9270) );
  XNOR U9515 ( .A(x[242]), .B(n9271), .Z(n9273) );
  XOR U9516 ( .A(n9274), .B(n9275), .Z(n9271) );
  AND U9517 ( .A(n9276), .B(n9277), .Z(n9274) );
  XNOR U9518 ( .A(x[241]), .B(n9275), .Z(n9277) );
  XOR U9519 ( .A(n9278), .B(n9279), .Z(n9275) );
  AND U9520 ( .A(n9280), .B(n9281), .Z(n9278) );
  XNOR U9521 ( .A(x[240]), .B(n9279), .Z(n9281) );
  XOR U9522 ( .A(n9282), .B(n9283), .Z(n9279) );
  AND U9523 ( .A(n9284), .B(n9285), .Z(n9282) );
  XNOR U9524 ( .A(x[239]), .B(n9283), .Z(n9285) );
  XOR U9525 ( .A(n9286), .B(n9287), .Z(n9283) );
  AND U9526 ( .A(n9288), .B(n9289), .Z(n9286) );
  XNOR U9527 ( .A(x[238]), .B(n9287), .Z(n9289) );
  XOR U9528 ( .A(n9290), .B(n9291), .Z(n9287) );
  AND U9529 ( .A(n9292), .B(n9293), .Z(n9290) );
  XNOR U9530 ( .A(x[237]), .B(n9291), .Z(n9293) );
  XOR U9531 ( .A(n9294), .B(n9295), .Z(n9291) );
  AND U9532 ( .A(n9296), .B(n9297), .Z(n9294) );
  XNOR U9533 ( .A(x[236]), .B(n9295), .Z(n9297) );
  XOR U9534 ( .A(n9298), .B(n9299), .Z(n9295) );
  AND U9535 ( .A(n9300), .B(n9301), .Z(n9298) );
  XNOR U9536 ( .A(x[235]), .B(n9299), .Z(n9301) );
  XOR U9537 ( .A(n9302), .B(n9303), .Z(n9299) );
  AND U9538 ( .A(n9304), .B(n9305), .Z(n9302) );
  XNOR U9539 ( .A(x[234]), .B(n9303), .Z(n9305) );
  XOR U9540 ( .A(n9306), .B(n9307), .Z(n9303) );
  AND U9541 ( .A(n9308), .B(n9309), .Z(n9306) );
  XNOR U9542 ( .A(x[233]), .B(n9307), .Z(n9309) );
  XOR U9543 ( .A(n9310), .B(n9311), .Z(n9307) );
  AND U9544 ( .A(n9312), .B(n9313), .Z(n9310) );
  XNOR U9545 ( .A(x[232]), .B(n9311), .Z(n9313) );
  XOR U9546 ( .A(n9314), .B(n9315), .Z(n9311) );
  AND U9547 ( .A(n9316), .B(n9317), .Z(n9314) );
  XNOR U9548 ( .A(x[231]), .B(n9315), .Z(n9317) );
  XOR U9549 ( .A(n9318), .B(n9319), .Z(n9315) );
  AND U9550 ( .A(n9320), .B(n9321), .Z(n9318) );
  XNOR U9551 ( .A(x[230]), .B(n9319), .Z(n9321) );
  XOR U9552 ( .A(n9322), .B(n9323), .Z(n9319) );
  AND U9553 ( .A(n9324), .B(n9325), .Z(n9322) );
  XNOR U9554 ( .A(x[229]), .B(n9323), .Z(n9325) );
  XOR U9555 ( .A(n9326), .B(n9327), .Z(n9323) );
  AND U9556 ( .A(n9328), .B(n9329), .Z(n9326) );
  XNOR U9557 ( .A(x[228]), .B(n9327), .Z(n9329) );
  XOR U9558 ( .A(n9330), .B(n9331), .Z(n9327) );
  AND U9559 ( .A(n9332), .B(n9333), .Z(n9330) );
  XNOR U9560 ( .A(x[227]), .B(n9331), .Z(n9333) );
  XOR U9561 ( .A(n9334), .B(n9335), .Z(n9331) );
  AND U9562 ( .A(n9336), .B(n9337), .Z(n9334) );
  XNOR U9563 ( .A(x[226]), .B(n9335), .Z(n9337) );
  XOR U9564 ( .A(n9338), .B(n9339), .Z(n9335) );
  AND U9565 ( .A(n9340), .B(n9341), .Z(n9338) );
  XNOR U9566 ( .A(x[225]), .B(n9339), .Z(n9341) );
  XOR U9567 ( .A(n9342), .B(n9343), .Z(n9339) );
  AND U9568 ( .A(n9344), .B(n9345), .Z(n9342) );
  XNOR U9569 ( .A(x[224]), .B(n9343), .Z(n9345) );
  XOR U9570 ( .A(n9346), .B(n9347), .Z(n9343) );
  AND U9571 ( .A(n9348), .B(n9349), .Z(n9346) );
  XNOR U9572 ( .A(x[223]), .B(n9347), .Z(n9349) );
  XOR U9573 ( .A(n9350), .B(n9351), .Z(n9347) );
  AND U9574 ( .A(n9352), .B(n9353), .Z(n9350) );
  XNOR U9575 ( .A(x[222]), .B(n9351), .Z(n9353) );
  XOR U9576 ( .A(n9354), .B(n9355), .Z(n9351) );
  AND U9577 ( .A(n9356), .B(n9357), .Z(n9354) );
  XNOR U9578 ( .A(x[221]), .B(n9355), .Z(n9357) );
  XOR U9579 ( .A(n9358), .B(n9359), .Z(n9355) );
  AND U9580 ( .A(n9360), .B(n9361), .Z(n9358) );
  XNOR U9581 ( .A(x[220]), .B(n9359), .Z(n9361) );
  XOR U9582 ( .A(n9362), .B(n9363), .Z(n9359) );
  AND U9583 ( .A(n9364), .B(n9365), .Z(n9362) );
  XNOR U9584 ( .A(x[219]), .B(n9363), .Z(n9365) );
  XOR U9585 ( .A(n9366), .B(n9367), .Z(n9363) );
  AND U9586 ( .A(n9368), .B(n9369), .Z(n9366) );
  XNOR U9587 ( .A(x[218]), .B(n9367), .Z(n9369) );
  XOR U9588 ( .A(n9370), .B(n9371), .Z(n9367) );
  AND U9589 ( .A(n9372), .B(n9373), .Z(n9370) );
  XNOR U9590 ( .A(x[217]), .B(n9371), .Z(n9373) );
  XOR U9591 ( .A(n9374), .B(n9375), .Z(n9371) );
  AND U9592 ( .A(n9376), .B(n9377), .Z(n9374) );
  XNOR U9593 ( .A(x[216]), .B(n9375), .Z(n9377) );
  XOR U9594 ( .A(n9378), .B(n9379), .Z(n9375) );
  AND U9595 ( .A(n9380), .B(n9381), .Z(n9378) );
  XNOR U9596 ( .A(x[215]), .B(n9379), .Z(n9381) );
  XOR U9597 ( .A(n9382), .B(n9383), .Z(n9379) );
  AND U9598 ( .A(n9384), .B(n9385), .Z(n9382) );
  XNOR U9599 ( .A(x[214]), .B(n9383), .Z(n9385) );
  XOR U9600 ( .A(n9386), .B(n9387), .Z(n9383) );
  AND U9601 ( .A(n9388), .B(n9389), .Z(n9386) );
  XNOR U9602 ( .A(x[213]), .B(n9387), .Z(n9389) );
  XOR U9603 ( .A(n9390), .B(n9391), .Z(n9387) );
  AND U9604 ( .A(n9392), .B(n9393), .Z(n9390) );
  XNOR U9605 ( .A(x[212]), .B(n9391), .Z(n9393) );
  XOR U9606 ( .A(n9394), .B(n9395), .Z(n9391) );
  AND U9607 ( .A(n9396), .B(n9397), .Z(n9394) );
  XNOR U9608 ( .A(x[211]), .B(n9395), .Z(n9397) );
  XOR U9609 ( .A(n9398), .B(n9399), .Z(n9395) );
  AND U9610 ( .A(n9400), .B(n9401), .Z(n9398) );
  XNOR U9611 ( .A(x[210]), .B(n9399), .Z(n9401) );
  XOR U9612 ( .A(n9402), .B(n9403), .Z(n9399) );
  AND U9613 ( .A(n9404), .B(n9405), .Z(n9402) );
  XNOR U9614 ( .A(x[209]), .B(n9403), .Z(n9405) );
  XOR U9615 ( .A(n9406), .B(n9407), .Z(n9403) );
  AND U9616 ( .A(n9408), .B(n9409), .Z(n9406) );
  XNOR U9617 ( .A(x[208]), .B(n9407), .Z(n9409) );
  XOR U9618 ( .A(n9410), .B(n9411), .Z(n9407) );
  AND U9619 ( .A(n9412), .B(n9413), .Z(n9410) );
  XNOR U9620 ( .A(x[207]), .B(n9411), .Z(n9413) );
  XOR U9621 ( .A(n9414), .B(n9415), .Z(n9411) );
  AND U9622 ( .A(n9416), .B(n9417), .Z(n9414) );
  XNOR U9623 ( .A(x[206]), .B(n9415), .Z(n9417) );
  XOR U9624 ( .A(n9418), .B(n9419), .Z(n9415) );
  AND U9625 ( .A(n9420), .B(n9421), .Z(n9418) );
  XNOR U9626 ( .A(x[205]), .B(n9419), .Z(n9421) );
  XOR U9627 ( .A(n9422), .B(n9423), .Z(n9419) );
  AND U9628 ( .A(n9424), .B(n9425), .Z(n9422) );
  XNOR U9629 ( .A(x[204]), .B(n9423), .Z(n9425) );
  XOR U9630 ( .A(n9426), .B(n9427), .Z(n9423) );
  AND U9631 ( .A(n9428), .B(n9429), .Z(n9426) );
  XNOR U9632 ( .A(x[203]), .B(n9427), .Z(n9429) );
  XOR U9633 ( .A(n9430), .B(n9431), .Z(n9427) );
  AND U9634 ( .A(n9432), .B(n9433), .Z(n9430) );
  XNOR U9635 ( .A(x[202]), .B(n9431), .Z(n9433) );
  XOR U9636 ( .A(n9434), .B(n9435), .Z(n9431) );
  AND U9637 ( .A(n9436), .B(n9437), .Z(n9434) );
  XNOR U9638 ( .A(x[201]), .B(n9435), .Z(n9437) );
  XOR U9639 ( .A(n9438), .B(n9439), .Z(n9435) );
  AND U9640 ( .A(n9440), .B(n9441), .Z(n9438) );
  XNOR U9641 ( .A(x[200]), .B(n9439), .Z(n9441) );
  XOR U9642 ( .A(n9442), .B(n9443), .Z(n9439) );
  AND U9643 ( .A(n9444), .B(n9445), .Z(n9442) );
  XNOR U9644 ( .A(x[199]), .B(n9443), .Z(n9445) );
  XOR U9645 ( .A(n9446), .B(n9447), .Z(n9443) );
  AND U9646 ( .A(n9448), .B(n9449), .Z(n9446) );
  XNOR U9647 ( .A(x[198]), .B(n9447), .Z(n9449) );
  XOR U9648 ( .A(n9450), .B(n9451), .Z(n9447) );
  AND U9649 ( .A(n9452), .B(n9453), .Z(n9450) );
  XNOR U9650 ( .A(x[197]), .B(n9451), .Z(n9453) );
  XOR U9651 ( .A(n9454), .B(n9455), .Z(n9451) );
  AND U9652 ( .A(n9456), .B(n9457), .Z(n9454) );
  XNOR U9653 ( .A(x[196]), .B(n9455), .Z(n9457) );
  XOR U9654 ( .A(n9458), .B(n9459), .Z(n9455) );
  AND U9655 ( .A(n9460), .B(n9461), .Z(n9458) );
  XNOR U9656 ( .A(x[195]), .B(n9459), .Z(n9461) );
  XOR U9657 ( .A(n9462), .B(n9463), .Z(n9459) );
  AND U9658 ( .A(n9464), .B(n9465), .Z(n9462) );
  XNOR U9659 ( .A(x[194]), .B(n9463), .Z(n9465) );
  XOR U9660 ( .A(n9466), .B(n9467), .Z(n9463) );
  AND U9661 ( .A(n9468), .B(n9469), .Z(n9466) );
  XNOR U9662 ( .A(x[193]), .B(n9467), .Z(n9469) );
  XOR U9663 ( .A(n9470), .B(n9471), .Z(n9467) );
  AND U9664 ( .A(n9472), .B(n9473), .Z(n9470) );
  XNOR U9665 ( .A(x[192]), .B(n9471), .Z(n9473) );
  XOR U9666 ( .A(n9474), .B(n9475), .Z(n9471) );
  AND U9667 ( .A(n9476), .B(n9477), .Z(n9474) );
  XNOR U9668 ( .A(x[191]), .B(n9475), .Z(n9477) );
  XOR U9669 ( .A(n9478), .B(n9479), .Z(n9475) );
  AND U9670 ( .A(n9480), .B(n9481), .Z(n9478) );
  XNOR U9671 ( .A(x[190]), .B(n9479), .Z(n9481) );
  XOR U9672 ( .A(n9482), .B(n9483), .Z(n9479) );
  AND U9673 ( .A(n9484), .B(n9485), .Z(n9482) );
  XNOR U9674 ( .A(x[189]), .B(n9483), .Z(n9485) );
  XOR U9675 ( .A(n9486), .B(n9487), .Z(n9483) );
  AND U9676 ( .A(n9488), .B(n9489), .Z(n9486) );
  XNOR U9677 ( .A(x[188]), .B(n9487), .Z(n9489) );
  XOR U9678 ( .A(n9490), .B(n9491), .Z(n9487) );
  AND U9679 ( .A(n9492), .B(n9493), .Z(n9490) );
  XNOR U9680 ( .A(x[187]), .B(n9491), .Z(n9493) );
  XOR U9681 ( .A(n9494), .B(n9495), .Z(n9491) );
  AND U9682 ( .A(n9496), .B(n9497), .Z(n9494) );
  XNOR U9683 ( .A(x[186]), .B(n9495), .Z(n9497) );
  XOR U9684 ( .A(n9498), .B(n9499), .Z(n9495) );
  AND U9685 ( .A(n9500), .B(n9501), .Z(n9498) );
  XNOR U9686 ( .A(x[185]), .B(n9499), .Z(n9501) );
  XOR U9687 ( .A(n9502), .B(n9503), .Z(n9499) );
  AND U9688 ( .A(n9504), .B(n9505), .Z(n9502) );
  XNOR U9689 ( .A(x[184]), .B(n9503), .Z(n9505) );
  XOR U9690 ( .A(n9506), .B(n9507), .Z(n9503) );
  AND U9691 ( .A(n9508), .B(n9509), .Z(n9506) );
  XNOR U9692 ( .A(x[183]), .B(n9507), .Z(n9509) );
  XOR U9693 ( .A(n9510), .B(n9511), .Z(n9507) );
  AND U9694 ( .A(n9512), .B(n9513), .Z(n9510) );
  XNOR U9695 ( .A(x[182]), .B(n9511), .Z(n9513) );
  XOR U9696 ( .A(n9514), .B(n9515), .Z(n9511) );
  AND U9697 ( .A(n9516), .B(n9517), .Z(n9514) );
  XNOR U9698 ( .A(x[181]), .B(n9515), .Z(n9517) );
  XOR U9699 ( .A(n9518), .B(n9519), .Z(n9515) );
  AND U9700 ( .A(n9520), .B(n9521), .Z(n9518) );
  XNOR U9701 ( .A(x[180]), .B(n9519), .Z(n9521) );
  XOR U9702 ( .A(n9522), .B(n9523), .Z(n9519) );
  AND U9703 ( .A(n9524), .B(n9525), .Z(n9522) );
  XNOR U9704 ( .A(x[179]), .B(n9523), .Z(n9525) );
  XOR U9705 ( .A(n9526), .B(n9527), .Z(n9523) );
  AND U9706 ( .A(n9528), .B(n9529), .Z(n9526) );
  XNOR U9707 ( .A(x[178]), .B(n9527), .Z(n9529) );
  XOR U9708 ( .A(n9530), .B(n9531), .Z(n9527) );
  AND U9709 ( .A(n9532), .B(n9533), .Z(n9530) );
  XNOR U9710 ( .A(x[177]), .B(n9531), .Z(n9533) );
  XOR U9711 ( .A(n9534), .B(n9535), .Z(n9531) );
  AND U9712 ( .A(n9536), .B(n9537), .Z(n9534) );
  XNOR U9713 ( .A(x[176]), .B(n9535), .Z(n9537) );
  XOR U9714 ( .A(n9538), .B(n9539), .Z(n9535) );
  AND U9715 ( .A(n9540), .B(n9541), .Z(n9538) );
  XNOR U9716 ( .A(x[175]), .B(n9539), .Z(n9541) );
  XOR U9717 ( .A(n9542), .B(n9543), .Z(n9539) );
  AND U9718 ( .A(n9544), .B(n9545), .Z(n9542) );
  XNOR U9719 ( .A(x[174]), .B(n9543), .Z(n9545) );
  XOR U9720 ( .A(n9546), .B(n9547), .Z(n9543) );
  AND U9721 ( .A(n9548), .B(n9549), .Z(n9546) );
  XNOR U9722 ( .A(x[173]), .B(n9547), .Z(n9549) );
  XOR U9723 ( .A(n9550), .B(n9551), .Z(n9547) );
  AND U9724 ( .A(n9552), .B(n9553), .Z(n9550) );
  XNOR U9725 ( .A(x[172]), .B(n9551), .Z(n9553) );
  XOR U9726 ( .A(n9554), .B(n9555), .Z(n9551) );
  AND U9727 ( .A(n9556), .B(n9557), .Z(n9554) );
  XNOR U9728 ( .A(x[171]), .B(n9555), .Z(n9557) );
  XOR U9729 ( .A(n9558), .B(n9559), .Z(n9555) );
  AND U9730 ( .A(n9560), .B(n9561), .Z(n9558) );
  XNOR U9731 ( .A(x[170]), .B(n9559), .Z(n9561) );
  XOR U9732 ( .A(n9562), .B(n9563), .Z(n9559) );
  AND U9733 ( .A(n9564), .B(n9565), .Z(n9562) );
  XNOR U9734 ( .A(x[169]), .B(n9563), .Z(n9565) );
  XOR U9735 ( .A(n9566), .B(n9567), .Z(n9563) );
  AND U9736 ( .A(n9568), .B(n9569), .Z(n9566) );
  XNOR U9737 ( .A(x[168]), .B(n9567), .Z(n9569) );
  XOR U9738 ( .A(n9570), .B(n9571), .Z(n9567) );
  AND U9739 ( .A(n9572), .B(n9573), .Z(n9570) );
  XNOR U9740 ( .A(x[167]), .B(n9571), .Z(n9573) );
  XOR U9741 ( .A(n9574), .B(n9575), .Z(n9571) );
  AND U9742 ( .A(n9576), .B(n9577), .Z(n9574) );
  XNOR U9743 ( .A(x[166]), .B(n9575), .Z(n9577) );
  XOR U9744 ( .A(n9578), .B(n9579), .Z(n9575) );
  AND U9745 ( .A(n9580), .B(n9581), .Z(n9578) );
  XNOR U9746 ( .A(x[165]), .B(n9579), .Z(n9581) );
  XOR U9747 ( .A(n9582), .B(n9583), .Z(n9579) );
  AND U9748 ( .A(n9584), .B(n9585), .Z(n9582) );
  XNOR U9749 ( .A(x[164]), .B(n9583), .Z(n9585) );
  XOR U9750 ( .A(n9586), .B(n9587), .Z(n9583) );
  AND U9751 ( .A(n9588), .B(n9589), .Z(n9586) );
  XNOR U9752 ( .A(x[163]), .B(n9587), .Z(n9589) );
  XOR U9753 ( .A(n9590), .B(n9591), .Z(n9587) );
  AND U9754 ( .A(n9592), .B(n9593), .Z(n9590) );
  XNOR U9755 ( .A(x[162]), .B(n9591), .Z(n9593) );
  XOR U9756 ( .A(n9594), .B(n9595), .Z(n9591) );
  AND U9757 ( .A(n9596), .B(n9597), .Z(n9594) );
  XNOR U9758 ( .A(x[161]), .B(n9595), .Z(n9597) );
  XOR U9759 ( .A(n9598), .B(n9599), .Z(n9595) );
  AND U9760 ( .A(n9600), .B(n9601), .Z(n9598) );
  XNOR U9761 ( .A(x[160]), .B(n9599), .Z(n9601) );
  XOR U9762 ( .A(n9602), .B(n9603), .Z(n9599) );
  AND U9763 ( .A(n9604), .B(n9605), .Z(n9602) );
  XNOR U9764 ( .A(x[159]), .B(n9603), .Z(n9605) );
  XOR U9765 ( .A(n9606), .B(n9607), .Z(n9603) );
  AND U9766 ( .A(n9608), .B(n9609), .Z(n9606) );
  XNOR U9767 ( .A(x[158]), .B(n9607), .Z(n9609) );
  XOR U9768 ( .A(n9610), .B(n9611), .Z(n9607) );
  AND U9769 ( .A(n9612), .B(n9613), .Z(n9610) );
  XNOR U9770 ( .A(x[157]), .B(n9611), .Z(n9613) );
  XOR U9771 ( .A(n9614), .B(n9615), .Z(n9611) );
  AND U9772 ( .A(n9616), .B(n9617), .Z(n9614) );
  XNOR U9773 ( .A(x[156]), .B(n9615), .Z(n9617) );
  XOR U9774 ( .A(n9618), .B(n9619), .Z(n9615) );
  AND U9775 ( .A(n9620), .B(n9621), .Z(n9618) );
  XNOR U9776 ( .A(x[155]), .B(n9619), .Z(n9621) );
  XOR U9777 ( .A(n9622), .B(n9623), .Z(n9619) );
  AND U9778 ( .A(n9624), .B(n9625), .Z(n9622) );
  XNOR U9779 ( .A(x[154]), .B(n9623), .Z(n9625) );
  XOR U9780 ( .A(n9626), .B(n9627), .Z(n9623) );
  AND U9781 ( .A(n9628), .B(n9629), .Z(n9626) );
  XNOR U9782 ( .A(x[153]), .B(n9627), .Z(n9629) );
  XOR U9783 ( .A(n9630), .B(n9631), .Z(n9627) );
  AND U9784 ( .A(n9632), .B(n9633), .Z(n9630) );
  XNOR U9785 ( .A(x[152]), .B(n9631), .Z(n9633) );
  XOR U9786 ( .A(n9634), .B(n9635), .Z(n9631) );
  AND U9787 ( .A(n9636), .B(n9637), .Z(n9634) );
  XNOR U9788 ( .A(x[151]), .B(n9635), .Z(n9637) );
  XOR U9789 ( .A(n9638), .B(n9639), .Z(n9635) );
  AND U9790 ( .A(n9640), .B(n9641), .Z(n9638) );
  XNOR U9791 ( .A(x[150]), .B(n9639), .Z(n9641) );
  XOR U9792 ( .A(n9642), .B(n9643), .Z(n9639) );
  AND U9793 ( .A(n9644), .B(n9645), .Z(n9642) );
  XNOR U9794 ( .A(x[149]), .B(n9643), .Z(n9645) );
  XOR U9795 ( .A(n9646), .B(n9647), .Z(n9643) );
  AND U9796 ( .A(n9648), .B(n9649), .Z(n9646) );
  XNOR U9797 ( .A(x[148]), .B(n9647), .Z(n9649) );
  XOR U9798 ( .A(n9650), .B(n9651), .Z(n9647) );
  AND U9799 ( .A(n9652), .B(n9653), .Z(n9650) );
  XNOR U9800 ( .A(x[147]), .B(n9651), .Z(n9653) );
  XOR U9801 ( .A(n9654), .B(n9655), .Z(n9651) );
  AND U9802 ( .A(n9656), .B(n9657), .Z(n9654) );
  XNOR U9803 ( .A(x[146]), .B(n9655), .Z(n9657) );
  XOR U9804 ( .A(n9658), .B(n9659), .Z(n9655) );
  AND U9805 ( .A(n9660), .B(n9661), .Z(n9658) );
  XNOR U9806 ( .A(x[145]), .B(n9659), .Z(n9661) );
  XOR U9807 ( .A(n9662), .B(n9663), .Z(n9659) );
  AND U9808 ( .A(n9664), .B(n9665), .Z(n9662) );
  XNOR U9809 ( .A(x[144]), .B(n9663), .Z(n9665) );
  XOR U9810 ( .A(n9666), .B(n9667), .Z(n9663) );
  AND U9811 ( .A(n9668), .B(n9669), .Z(n9666) );
  XNOR U9812 ( .A(x[143]), .B(n9667), .Z(n9669) );
  XOR U9813 ( .A(n9670), .B(n9671), .Z(n9667) );
  AND U9814 ( .A(n9672), .B(n9673), .Z(n9670) );
  XNOR U9815 ( .A(x[142]), .B(n9671), .Z(n9673) );
  XOR U9816 ( .A(n9674), .B(n9675), .Z(n9671) );
  AND U9817 ( .A(n9676), .B(n9677), .Z(n9674) );
  XNOR U9818 ( .A(x[141]), .B(n9675), .Z(n9677) );
  XOR U9819 ( .A(n9678), .B(n9679), .Z(n9675) );
  AND U9820 ( .A(n9680), .B(n9681), .Z(n9678) );
  XNOR U9821 ( .A(x[140]), .B(n9679), .Z(n9681) );
  XOR U9822 ( .A(n9682), .B(n9683), .Z(n9679) );
  AND U9823 ( .A(n9684), .B(n9685), .Z(n9682) );
  XNOR U9824 ( .A(x[139]), .B(n9683), .Z(n9685) );
  XOR U9825 ( .A(n9686), .B(n9687), .Z(n9683) );
  AND U9826 ( .A(n9688), .B(n9689), .Z(n9686) );
  XNOR U9827 ( .A(x[138]), .B(n9687), .Z(n9689) );
  XOR U9828 ( .A(n9690), .B(n9691), .Z(n9687) );
  AND U9829 ( .A(n9692), .B(n9693), .Z(n9690) );
  XNOR U9830 ( .A(x[137]), .B(n9691), .Z(n9693) );
  XOR U9831 ( .A(n9694), .B(n9695), .Z(n9691) );
  AND U9832 ( .A(n9696), .B(n9697), .Z(n9694) );
  XNOR U9833 ( .A(x[136]), .B(n9695), .Z(n9697) );
  XOR U9834 ( .A(n9698), .B(n9699), .Z(n9695) );
  AND U9835 ( .A(n9700), .B(n9701), .Z(n9698) );
  XNOR U9836 ( .A(x[135]), .B(n9699), .Z(n9701) );
  XOR U9837 ( .A(n9702), .B(n9703), .Z(n9699) );
  AND U9838 ( .A(n9704), .B(n9705), .Z(n9702) );
  XNOR U9839 ( .A(x[134]), .B(n9703), .Z(n9705) );
  XOR U9840 ( .A(n9706), .B(n9707), .Z(n9703) );
  AND U9841 ( .A(n9708), .B(n9709), .Z(n9706) );
  XNOR U9842 ( .A(x[133]), .B(n9707), .Z(n9709) );
  XOR U9843 ( .A(n9710), .B(n9711), .Z(n9707) );
  AND U9844 ( .A(n9712), .B(n9713), .Z(n9710) );
  XNOR U9845 ( .A(x[132]), .B(n9711), .Z(n9713) );
  XOR U9846 ( .A(n9714), .B(n9715), .Z(n9711) );
  AND U9847 ( .A(n9716), .B(n9717), .Z(n9714) );
  XNOR U9848 ( .A(x[131]), .B(n9715), .Z(n9717) );
  XOR U9849 ( .A(n9718), .B(n9719), .Z(n9715) );
  AND U9850 ( .A(n9720), .B(n9721), .Z(n9718) );
  XNOR U9851 ( .A(x[130]), .B(n9719), .Z(n9721) );
  XOR U9852 ( .A(n9722), .B(n9723), .Z(n9719) );
  AND U9853 ( .A(n9724), .B(n9725), .Z(n9722) );
  XNOR U9854 ( .A(x[129]), .B(n9723), .Z(n9725) );
  XOR U9855 ( .A(n9726), .B(n9727), .Z(n9723) );
  AND U9856 ( .A(n9728), .B(n9729), .Z(n9726) );
  XNOR U9857 ( .A(x[128]), .B(n9727), .Z(n9729) );
  XOR U9858 ( .A(n9730), .B(n9731), .Z(n9727) );
  AND U9859 ( .A(n9732), .B(n9733), .Z(n9730) );
  XNOR U9860 ( .A(x[127]), .B(n9731), .Z(n9733) );
  XOR U9861 ( .A(n9734), .B(n9735), .Z(n9731) );
  AND U9862 ( .A(n9736), .B(n9737), .Z(n9734) );
  XNOR U9863 ( .A(x[126]), .B(n9735), .Z(n9737) );
  XOR U9864 ( .A(n9738), .B(n9739), .Z(n9735) );
  AND U9865 ( .A(n9740), .B(n9741), .Z(n9738) );
  XNOR U9866 ( .A(x[125]), .B(n9739), .Z(n9741) );
  XOR U9867 ( .A(n9742), .B(n9743), .Z(n9739) );
  AND U9868 ( .A(n9744), .B(n9745), .Z(n9742) );
  XNOR U9869 ( .A(x[124]), .B(n9743), .Z(n9745) );
  XOR U9870 ( .A(n9746), .B(n9747), .Z(n9743) );
  AND U9871 ( .A(n9748), .B(n9749), .Z(n9746) );
  XNOR U9872 ( .A(x[123]), .B(n9747), .Z(n9749) );
  XOR U9873 ( .A(n9750), .B(n9751), .Z(n9747) );
  AND U9874 ( .A(n9752), .B(n9753), .Z(n9750) );
  XNOR U9875 ( .A(x[122]), .B(n9751), .Z(n9753) );
  XOR U9876 ( .A(n9754), .B(n9755), .Z(n9751) );
  AND U9877 ( .A(n9756), .B(n9757), .Z(n9754) );
  XNOR U9878 ( .A(x[121]), .B(n9755), .Z(n9757) );
  XOR U9879 ( .A(n9758), .B(n9759), .Z(n9755) );
  AND U9880 ( .A(n9760), .B(n9761), .Z(n9758) );
  XNOR U9881 ( .A(x[120]), .B(n9759), .Z(n9761) );
  XOR U9882 ( .A(n9762), .B(n9763), .Z(n9759) );
  AND U9883 ( .A(n9764), .B(n9765), .Z(n9762) );
  XNOR U9884 ( .A(x[119]), .B(n9763), .Z(n9765) );
  XOR U9885 ( .A(n9766), .B(n9767), .Z(n9763) );
  AND U9886 ( .A(n9768), .B(n9769), .Z(n9766) );
  XNOR U9887 ( .A(x[118]), .B(n9767), .Z(n9769) );
  XOR U9888 ( .A(n9770), .B(n9771), .Z(n9767) );
  AND U9889 ( .A(n9772), .B(n9773), .Z(n9770) );
  XNOR U9890 ( .A(x[117]), .B(n9771), .Z(n9773) );
  XOR U9891 ( .A(n9774), .B(n9775), .Z(n9771) );
  AND U9892 ( .A(n9776), .B(n9777), .Z(n9774) );
  XNOR U9893 ( .A(x[116]), .B(n9775), .Z(n9777) );
  XOR U9894 ( .A(n9778), .B(n9779), .Z(n9775) );
  AND U9895 ( .A(n9780), .B(n9781), .Z(n9778) );
  XNOR U9896 ( .A(x[115]), .B(n9779), .Z(n9781) );
  XOR U9897 ( .A(n9782), .B(n9783), .Z(n9779) );
  AND U9898 ( .A(n9784), .B(n9785), .Z(n9782) );
  XNOR U9899 ( .A(x[114]), .B(n9783), .Z(n9785) );
  XOR U9900 ( .A(n9786), .B(n9787), .Z(n9783) );
  AND U9901 ( .A(n9788), .B(n9789), .Z(n9786) );
  XNOR U9902 ( .A(x[113]), .B(n9787), .Z(n9789) );
  XOR U9903 ( .A(n9790), .B(n9791), .Z(n9787) );
  AND U9904 ( .A(n9792), .B(n9793), .Z(n9790) );
  XNOR U9905 ( .A(x[112]), .B(n9791), .Z(n9793) );
  XOR U9906 ( .A(n9794), .B(n9795), .Z(n9791) );
  AND U9907 ( .A(n9796), .B(n9797), .Z(n9794) );
  XNOR U9908 ( .A(x[111]), .B(n9795), .Z(n9797) );
  XOR U9909 ( .A(n9798), .B(n9799), .Z(n9795) );
  AND U9910 ( .A(n9800), .B(n9801), .Z(n9798) );
  XNOR U9911 ( .A(x[110]), .B(n9799), .Z(n9801) );
  XOR U9912 ( .A(n9802), .B(n9803), .Z(n9799) );
  AND U9913 ( .A(n9804), .B(n9805), .Z(n9802) );
  XNOR U9914 ( .A(x[109]), .B(n9803), .Z(n9805) );
  XOR U9915 ( .A(n9806), .B(n9807), .Z(n9803) );
  AND U9916 ( .A(n9808), .B(n9809), .Z(n9806) );
  XNOR U9917 ( .A(x[108]), .B(n9807), .Z(n9809) );
  XOR U9918 ( .A(n9810), .B(n9811), .Z(n9807) );
  AND U9919 ( .A(n9812), .B(n9813), .Z(n9810) );
  XNOR U9920 ( .A(x[107]), .B(n9811), .Z(n9813) );
  XOR U9921 ( .A(n9814), .B(n9815), .Z(n9811) );
  AND U9922 ( .A(n9816), .B(n9817), .Z(n9814) );
  XNOR U9923 ( .A(x[106]), .B(n9815), .Z(n9817) );
  XOR U9924 ( .A(n9818), .B(n9819), .Z(n9815) );
  AND U9925 ( .A(n9820), .B(n9821), .Z(n9818) );
  XNOR U9926 ( .A(x[105]), .B(n9819), .Z(n9821) );
  XOR U9927 ( .A(n9822), .B(n9823), .Z(n9819) );
  AND U9928 ( .A(n9824), .B(n9825), .Z(n9822) );
  XNOR U9929 ( .A(x[104]), .B(n9823), .Z(n9825) );
  XOR U9930 ( .A(n9826), .B(n9827), .Z(n9823) );
  AND U9931 ( .A(n9828), .B(n9829), .Z(n9826) );
  XNOR U9932 ( .A(x[103]), .B(n9827), .Z(n9829) );
  XOR U9933 ( .A(n9830), .B(n9831), .Z(n9827) );
  AND U9934 ( .A(n9832), .B(n9833), .Z(n9830) );
  XNOR U9935 ( .A(x[102]), .B(n9831), .Z(n9833) );
  XOR U9936 ( .A(n9834), .B(n9835), .Z(n9831) );
  AND U9937 ( .A(n9836), .B(n9837), .Z(n9834) );
  XNOR U9938 ( .A(x[101]), .B(n9835), .Z(n9837) );
  XOR U9939 ( .A(n9838), .B(n9839), .Z(n9835) );
  AND U9940 ( .A(n9840), .B(n9841), .Z(n9838) );
  XNOR U9941 ( .A(x[100]), .B(n9839), .Z(n9841) );
  XOR U9942 ( .A(n9842), .B(n9843), .Z(n9839) );
  AND U9943 ( .A(n9844), .B(n9845), .Z(n9842) );
  XNOR U9944 ( .A(x[99]), .B(n9843), .Z(n9845) );
  XOR U9945 ( .A(n9846), .B(n9847), .Z(n9843) );
  AND U9946 ( .A(n9848), .B(n9849), .Z(n9846) );
  XNOR U9947 ( .A(x[98]), .B(n9847), .Z(n9849) );
  XOR U9948 ( .A(n9850), .B(n9851), .Z(n9847) );
  AND U9949 ( .A(n9852), .B(n9853), .Z(n9850) );
  XNOR U9950 ( .A(x[97]), .B(n9851), .Z(n9853) );
  XOR U9951 ( .A(n9854), .B(n9855), .Z(n9851) );
  AND U9952 ( .A(n9856), .B(n9857), .Z(n9854) );
  XNOR U9953 ( .A(x[96]), .B(n9855), .Z(n9857) );
  XOR U9954 ( .A(n9858), .B(n9859), .Z(n9855) );
  AND U9955 ( .A(n9860), .B(n9861), .Z(n9858) );
  XNOR U9956 ( .A(x[95]), .B(n9859), .Z(n9861) );
  XOR U9957 ( .A(n9862), .B(n9863), .Z(n9859) );
  AND U9958 ( .A(n9864), .B(n9865), .Z(n9862) );
  XNOR U9959 ( .A(x[94]), .B(n9863), .Z(n9865) );
  XOR U9960 ( .A(n9866), .B(n9867), .Z(n9863) );
  AND U9961 ( .A(n9868), .B(n9869), .Z(n9866) );
  XNOR U9962 ( .A(x[93]), .B(n9867), .Z(n9869) );
  XOR U9963 ( .A(n9870), .B(n9871), .Z(n9867) );
  AND U9964 ( .A(n9872), .B(n9873), .Z(n9870) );
  XNOR U9965 ( .A(x[92]), .B(n9871), .Z(n9873) );
  XOR U9966 ( .A(n9874), .B(n9875), .Z(n9871) );
  AND U9967 ( .A(n9876), .B(n9877), .Z(n9874) );
  XNOR U9968 ( .A(x[91]), .B(n9875), .Z(n9877) );
  XOR U9969 ( .A(n9878), .B(n9879), .Z(n9875) );
  AND U9970 ( .A(n9880), .B(n9881), .Z(n9878) );
  XNOR U9971 ( .A(x[90]), .B(n9879), .Z(n9881) );
  XOR U9972 ( .A(n9882), .B(n9883), .Z(n9879) );
  AND U9973 ( .A(n9884), .B(n9885), .Z(n9882) );
  XNOR U9974 ( .A(x[89]), .B(n9883), .Z(n9885) );
  XOR U9975 ( .A(n9886), .B(n9887), .Z(n9883) );
  AND U9976 ( .A(n9888), .B(n9889), .Z(n9886) );
  XNOR U9977 ( .A(x[88]), .B(n9887), .Z(n9889) );
  XOR U9978 ( .A(n9890), .B(n9891), .Z(n9887) );
  AND U9979 ( .A(n9892), .B(n9893), .Z(n9890) );
  XNOR U9980 ( .A(x[87]), .B(n9891), .Z(n9893) );
  XOR U9981 ( .A(n9894), .B(n9895), .Z(n9891) );
  AND U9982 ( .A(n9896), .B(n9897), .Z(n9894) );
  XNOR U9983 ( .A(x[86]), .B(n9895), .Z(n9897) );
  XOR U9984 ( .A(n9898), .B(n9899), .Z(n9895) );
  AND U9985 ( .A(n9900), .B(n9901), .Z(n9898) );
  XNOR U9986 ( .A(x[85]), .B(n9899), .Z(n9901) );
  XOR U9987 ( .A(n9902), .B(n9903), .Z(n9899) );
  AND U9988 ( .A(n9904), .B(n9905), .Z(n9902) );
  XNOR U9989 ( .A(x[84]), .B(n9903), .Z(n9905) );
  XOR U9990 ( .A(n9906), .B(n9907), .Z(n9903) );
  AND U9991 ( .A(n9908), .B(n9909), .Z(n9906) );
  XNOR U9992 ( .A(x[83]), .B(n9907), .Z(n9909) );
  XOR U9993 ( .A(n9910), .B(n9911), .Z(n9907) );
  AND U9994 ( .A(n9912), .B(n9913), .Z(n9910) );
  XNOR U9995 ( .A(x[82]), .B(n9911), .Z(n9913) );
  XOR U9996 ( .A(n9914), .B(n9915), .Z(n9911) );
  AND U9997 ( .A(n9916), .B(n9917), .Z(n9914) );
  XNOR U9998 ( .A(x[81]), .B(n9915), .Z(n9917) );
  XOR U9999 ( .A(n9918), .B(n9919), .Z(n9915) );
  AND U10000 ( .A(n9920), .B(n9921), .Z(n9918) );
  XNOR U10001 ( .A(x[80]), .B(n9919), .Z(n9921) );
  XOR U10002 ( .A(n9922), .B(n9923), .Z(n9919) );
  AND U10003 ( .A(n9924), .B(n9925), .Z(n9922) );
  XNOR U10004 ( .A(x[79]), .B(n9923), .Z(n9925) );
  XOR U10005 ( .A(n9926), .B(n9927), .Z(n9923) );
  AND U10006 ( .A(n9928), .B(n9929), .Z(n9926) );
  XNOR U10007 ( .A(x[78]), .B(n9927), .Z(n9929) );
  XOR U10008 ( .A(n9930), .B(n9931), .Z(n9927) );
  AND U10009 ( .A(n9932), .B(n9933), .Z(n9930) );
  XNOR U10010 ( .A(x[77]), .B(n9931), .Z(n9933) );
  XOR U10011 ( .A(n9934), .B(n9935), .Z(n9931) );
  AND U10012 ( .A(n9936), .B(n9937), .Z(n9934) );
  XNOR U10013 ( .A(x[76]), .B(n9935), .Z(n9937) );
  XOR U10014 ( .A(n9938), .B(n9939), .Z(n9935) );
  AND U10015 ( .A(n9940), .B(n9941), .Z(n9938) );
  XNOR U10016 ( .A(x[75]), .B(n9939), .Z(n9941) );
  XOR U10017 ( .A(n9942), .B(n9943), .Z(n9939) );
  AND U10018 ( .A(n9944), .B(n9945), .Z(n9942) );
  XNOR U10019 ( .A(x[74]), .B(n9943), .Z(n9945) );
  XOR U10020 ( .A(n9946), .B(n9947), .Z(n9943) );
  AND U10021 ( .A(n9948), .B(n9949), .Z(n9946) );
  XNOR U10022 ( .A(x[73]), .B(n9947), .Z(n9949) );
  XOR U10023 ( .A(n9950), .B(n9951), .Z(n9947) );
  AND U10024 ( .A(n9952), .B(n9953), .Z(n9950) );
  XNOR U10025 ( .A(x[72]), .B(n9951), .Z(n9953) );
  XOR U10026 ( .A(n9954), .B(n9955), .Z(n9951) );
  AND U10027 ( .A(n9956), .B(n9957), .Z(n9954) );
  XNOR U10028 ( .A(x[71]), .B(n9955), .Z(n9957) );
  XOR U10029 ( .A(n9958), .B(n9959), .Z(n9955) );
  AND U10030 ( .A(n9960), .B(n9961), .Z(n9958) );
  XNOR U10031 ( .A(x[70]), .B(n9959), .Z(n9961) );
  XOR U10032 ( .A(n9962), .B(n9963), .Z(n9959) );
  AND U10033 ( .A(n9964), .B(n9965), .Z(n9962) );
  XNOR U10034 ( .A(x[69]), .B(n9963), .Z(n9965) );
  XOR U10035 ( .A(n9966), .B(n9967), .Z(n9963) );
  AND U10036 ( .A(n9968), .B(n9969), .Z(n9966) );
  XNOR U10037 ( .A(x[68]), .B(n9967), .Z(n9969) );
  XOR U10038 ( .A(n9970), .B(n9971), .Z(n9967) );
  AND U10039 ( .A(n9972), .B(n9973), .Z(n9970) );
  XNOR U10040 ( .A(x[67]), .B(n9971), .Z(n9973) );
  XOR U10041 ( .A(n9974), .B(n9975), .Z(n9971) );
  AND U10042 ( .A(n9976), .B(n9977), .Z(n9974) );
  XNOR U10043 ( .A(x[66]), .B(n9975), .Z(n9977) );
  XOR U10044 ( .A(n9978), .B(n9979), .Z(n9975) );
  AND U10045 ( .A(n9980), .B(n9981), .Z(n9978) );
  XNOR U10046 ( .A(x[65]), .B(n9979), .Z(n9981) );
  XOR U10047 ( .A(n9982), .B(n9983), .Z(n9979) );
  AND U10048 ( .A(n9984), .B(n9985), .Z(n9982) );
  XNOR U10049 ( .A(x[64]), .B(n9983), .Z(n9985) );
  XOR U10050 ( .A(n9986), .B(n9987), .Z(n9983) );
  AND U10051 ( .A(n9988), .B(n9989), .Z(n9986) );
  XNOR U10052 ( .A(x[63]), .B(n9987), .Z(n9989) );
  XOR U10053 ( .A(n9990), .B(n9991), .Z(n9987) );
  AND U10054 ( .A(n9992), .B(n9993), .Z(n9990) );
  XNOR U10055 ( .A(x[62]), .B(n9991), .Z(n9993) );
  XOR U10056 ( .A(n9994), .B(n9995), .Z(n9991) );
  AND U10057 ( .A(n9996), .B(n9997), .Z(n9994) );
  XNOR U10058 ( .A(x[61]), .B(n9995), .Z(n9997) );
  XOR U10059 ( .A(n9998), .B(n9999), .Z(n9995) );
  AND U10060 ( .A(n10000), .B(n10001), .Z(n9998) );
  XNOR U10061 ( .A(x[60]), .B(n9999), .Z(n10001) );
  XOR U10062 ( .A(n10002), .B(n10003), .Z(n9999) );
  AND U10063 ( .A(n10004), .B(n10005), .Z(n10002) );
  XNOR U10064 ( .A(x[59]), .B(n10003), .Z(n10005) );
  XOR U10065 ( .A(n10006), .B(n10007), .Z(n10003) );
  AND U10066 ( .A(n10008), .B(n10009), .Z(n10006) );
  XNOR U10067 ( .A(x[58]), .B(n10007), .Z(n10009) );
  XOR U10068 ( .A(n10010), .B(n10011), .Z(n10007) );
  AND U10069 ( .A(n10012), .B(n10013), .Z(n10010) );
  XNOR U10070 ( .A(x[57]), .B(n10011), .Z(n10013) );
  XOR U10071 ( .A(n10014), .B(n10015), .Z(n10011) );
  AND U10072 ( .A(n10016), .B(n10017), .Z(n10014) );
  XNOR U10073 ( .A(x[56]), .B(n10015), .Z(n10017) );
  XOR U10074 ( .A(n10018), .B(n10019), .Z(n10015) );
  AND U10075 ( .A(n10020), .B(n10021), .Z(n10018) );
  XNOR U10076 ( .A(x[55]), .B(n10019), .Z(n10021) );
  XOR U10077 ( .A(n10022), .B(n10023), .Z(n10019) );
  AND U10078 ( .A(n10024), .B(n10025), .Z(n10022) );
  XNOR U10079 ( .A(x[54]), .B(n10023), .Z(n10025) );
  XOR U10080 ( .A(n10026), .B(n10027), .Z(n10023) );
  AND U10081 ( .A(n10028), .B(n10029), .Z(n10026) );
  XNOR U10082 ( .A(x[53]), .B(n10027), .Z(n10029) );
  XOR U10083 ( .A(n10030), .B(n10031), .Z(n10027) );
  AND U10084 ( .A(n10032), .B(n10033), .Z(n10030) );
  XNOR U10085 ( .A(x[52]), .B(n10031), .Z(n10033) );
  XOR U10086 ( .A(n10034), .B(n10035), .Z(n10031) );
  AND U10087 ( .A(n10036), .B(n10037), .Z(n10034) );
  XNOR U10088 ( .A(x[51]), .B(n10035), .Z(n10037) );
  XOR U10089 ( .A(n10038), .B(n10039), .Z(n10035) );
  AND U10090 ( .A(n10040), .B(n10041), .Z(n10038) );
  XNOR U10091 ( .A(x[50]), .B(n10039), .Z(n10041) );
  XOR U10092 ( .A(n10042), .B(n10043), .Z(n10039) );
  AND U10093 ( .A(n10044), .B(n10045), .Z(n10042) );
  XNOR U10094 ( .A(x[49]), .B(n10043), .Z(n10045) );
  XOR U10095 ( .A(n10046), .B(n10047), .Z(n10043) );
  AND U10096 ( .A(n10048), .B(n10049), .Z(n10046) );
  XNOR U10097 ( .A(x[48]), .B(n10047), .Z(n10049) );
  XOR U10098 ( .A(n10050), .B(n10051), .Z(n10047) );
  AND U10099 ( .A(n10052), .B(n10053), .Z(n10050) );
  XNOR U10100 ( .A(x[47]), .B(n10051), .Z(n10053) );
  XOR U10101 ( .A(n10054), .B(n10055), .Z(n10051) );
  AND U10102 ( .A(n10056), .B(n10057), .Z(n10054) );
  XNOR U10103 ( .A(x[46]), .B(n10055), .Z(n10057) );
  XOR U10104 ( .A(n10058), .B(n10059), .Z(n10055) );
  AND U10105 ( .A(n10060), .B(n10061), .Z(n10058) );
  XNOR U10106 ( .A(x[45]), .B(n10059), .Z(n10061) );
  XOR U10107 ( .A(n10062), .B(n10063), .Z(n10059) );
  AND U10108 ( .A(n10064), .B(n10065), .Z(n10062) );
  XNOR U10109 ( .A(x[44]), .B(n10063), .Z(n10065) );
  XOR U10110 ( .A(n10066), .B(n10067), .Z(n10063) );
  AND U10111 ( .A(n10068), .B(n10069), .Z(n10066) );
  XNOR U10112 ( .A(x[43]), .B(n10067), .Z(n10069) );
  XOR U10113 ( .A(n10070), .B(n10071), .Z(n10067) );
  AND U10114 ( .A(n10072), .B(n10073), .Z(n10070) );
  XNOR U10115 ( .A(x[42]), .B(n10071), .Z(n10073) );
  XOR U10116 ( .A(n10074), .B(n10075), .Z(n10071) );
  AND U10117 ( .A(n10076), .B(n10077), .Z(n10074) );
  XNOR U10118 ( .A(x[41]), .B(n10075), .Z(n10077) );
  XOR U10119 ( .A(n10078), .B(n10079), .Z(n10075) );
  AND U10120 ( .A(n10080), .B(n10081), .Z(n10078) );
  XNOR U10121 ( .A(x[40]), .B(n10079), .Z(n10081) );
  XOR U10122 ( .A(n10082), .B(n10083), .Z(n10079) );
  AND U10123 ( .A(n10084), .B(n10085), .Z(n10082) );
  XNOR U10124 ( .A(x[39]), .B(n10083), .Z(n10085) );
  XOR U10125 ( .A(n10086), .B(n10087), .Z(n10083) );
  AND U10126 ( .A(n10088), .B(n10089), .Z(n10086) );
  XNOR U10127 ( .A(x[38]), .B(n10087), .Z(n10089) );
  XOR U10128 ( .A(n10090), .B(n10091), .Z(n10087) );
  AND U10129 ( .A(n10092), .B(n10093), .Z(n10090) );
  XNOR U10130 ( .A(x[37]), .B(n10091), .Z(n10093) );
  XOR U10131 ( .A(n10094), .B(n10095), .Z(n10091) );
  AND U10132 ( .A(n10096), .B(n10097), .Z(n10094) );
  XNOR U10133 ( .A(x[36]), .B(n10095), .Z(n10097) );
  XOR U10134 ( .A(n10098), .B(n10099), .Z(n10095) );
  AND U10135 ( .A(n10100), .B(n10101), .Z(n10098) );
  XNOR U10136 ( .A(x[35]), .B(n10099), .Z(n10101) );
  XOR U10137 ( .A(n10102), .B(n10103), .Z(n10099) );
  AND U10138 ( .A(n10104), .B(n10105), .Z(n10102) );
  XNOR U10139 ( .A(x[34]), .B(n10103), .Z(n10105) );
  XOR U10140 ( .A(n10106), .B(n10107), .Z(n10103) );
  AND U10141 ( .A(n10108), .B(n10109), .Z(n10106) );
  XNOR U10142 ( .A(x[33]), .B(n10107), .Z(n10109) );
  XOR U10143 ( .A(n10110), .B(n10111), .Z(n10107) );
  AND U10144 ( .A(n10112), .B(n10113), .Z(n10110) );
  XNOR U10145 ( .A(x[32]), .B(n10111), .Z(n10113) );
  XOR U10146 ( .A(n10114), .B(n10115), .Z(n10111) );
  AND U10147 ( .A(n10116), .B(n10117), .Z(n10114) );
  XNOR U10148 ( .A(x[31]), .B(n10115), .Z(n10117) );
  XOR U10149 ( .A(n10118), .B(n10119), .Z(n10115) );
  AND U10150 ( .A(n10120), .B(n10121), .Z(n10118) );
  XNOR U10151 ( .A(x[30]), .B(n10119), .Z(n10121) );
  XOR U10152 ( .A(n10122), .B(n10123), .Z(n10119) );
  AND U10153 ( .A(n10124), .B(n10125), .Z(n10122) );
  XNOR U10154 ( .A(x[29]), .B(n10123), .Z(n10125) );
  XOR U10155 ( .A(n10126), .B(n10127), .Z(n10123) );
  AND U10156 ( .A(n10128), .B(n10129), .Z(n10126) );
  XNOR U10157 ( .A(x[28]), .B(n10127), .Z(n10129) );
  XOR U10158 ( .A(n10130), .B(n10131), .Z(n10127) );
  AND U10159 ( .A(n10132), .B(n10133), .Z(n10130) );
  XNOR U10160 ( .A(x[27]), .B(n10131), .Z(n10133) );
  XOR U10161 ( .A(n10134), .B(n10135), .Z(n10131) );
  AND U10162 ( .A(n10136), .B(n10137), .Z(n10134) );
  XNOR U10163 ( .A(x[26]), .B(n10135), .Z(n10137) );
  XOR U10164 ( .A(n10138), .B(n10139), .Z(n10135) );
  AND U10165 ( .A(n10140), .B(n10141), .Z(n10138) );
  XNOR U10166 ( .A(x[25]), .B(n10139), .Z(n10141) );
  XOR U10167 ( .A(n10142), .B(n10143), .Z(n10139) );
  AND U10168 ( .A(n10144), .B(n10145), .Z(n10142) );
  XNOR U10169 ( .A(x[24]), .B(n10143), .Z(n10145) );
  XOR U10170 ( .A(n10146), .B(n10147), .Z(n10143) );
  AND U10171 ( .A(n10148), .B(n10149), .Z(n10146) );
  XNOR U10172 ( .A(x[23]), .B(n10147), .Z(n10149) );
  XOR U10173 ( .A(n10150), .B(n10151), .Z(n10147) );
  AND U10174 ( .A(n10152), .B(n10153), .Z(n10150) );
  XNOR U10175 ( .A(x[22]), .B(n10151), .Z(n10153) );
  XOR U10176 ( .A(n10154), .B(n10155), .Z(n10151) );
  AND U10177 ( .A(n10156), .B(n10157), .Z(n10154) );
  XNOR U10178 ( .A(x[21]), .B(n10155), .Z(n10157) );
  XOR U10179 ( .A(n10158), .B(n10159), .Z(n10155) );
  AND U10180 ( .A(n10160), .B(n10161), .Z(n10158) );
  XNOR U10181 ( .A(x[20]), .B(n10159), .Z(n10161) );
  XOR U10182 ( .A(n10162), .B(n10163), .Z(n10159) );
  AND U10183 ( .A(n10164), .B(n10165), .Z(n10162) );
  XNOR U10184 ( .A(x[19]), .B(n10163), .Z(n10165) );
  XOR U10185 ( .A(n10166), .B(n10167), .Z(n10163) );
  AND U10186 ( .A(n10168), .B(n10169), .Z(n10166) );
  XNOR U10187 ( .A(x[18]), .B(n10167), .Z(n10169) );
  XOR U10188 ( .A(n10170), .B(n10171), .Z(n10167) );
  AND U10189 ( .A(n10172), .B(n10173), .Z(n10170) );
  XNOR U10190 ( .A(x[17]), .B(n10171), .Z(n10173) );
  XOR U10191 ( .A(n10174), .B(n10175), .Z(n10171) );
  AND U10192 ( .A(n10176), .B(n10177), .Z(n10174) );
  XNOR U10193 ( .A(x[16]), .B(n10175), .Z(n10177) );
  XOR U10194 ( .A(n10178), .B(n10179), .Z(n10175) );
  AND U10195 ( .A(n10180), .B(n10181), .Z(n10178) );
  XNOR U10196 ( .A(x[15]), .B(n10179), .Z(n10181) );
  XOR U10197 ( .A(n10182), .B(n10183), .Z(n10179) );
  AND U10198 ( .A(n10184), .B(n10185), .Z(n10182) );
  XNOR U10199 ( .A(x[14]), .B(n10183), .Z(n10185) );
  XOR U10200 ( .A(n10186), .B(n10187), .Z(n10183) );
  AND U10201 ( .A(n10188), .B(n10189), .Z(n10186) );
  XNOR U10202 ( .A(x[13]), .B(n10187), .Z(n10189) );
  XOR U10203 ( .A(n10190), .B(n10191), .Z(n10187) );
  AND U10204 ( .A(n10192), .B(n10193), .Z(n10190) );
  XNOR U10205 ( .A(x[12]), .B(n10191), .Z(n10193) );
  XOR U10206 ( .A(n10194), .B(n10195), .Z(n10191) );
  AND U10207 ( .A(n10196), .B(n10197), .Z(n10194) );
  XNOR U10208 ( .A(x[11]), .B(n10195), .Z(n10197) );
  XOR U10209 ( .A(n10198), .B(n10199), .Z(n10195) );
  AND U10210 ( .A(n10200), .B(n10201), .Z(n10198) );
  XNOR U10211 ( .A(x[10]), .B(n10199), .Z(n10201) );
  XOR U10212 ( .A(n10202), .B(n10203), .Z(n10199) );
  AND U10213 ( .A(n10204), .B(n10205), .Z(n10202) );
  XNOR U10214 ( .A(x[9]), .B(n10203), .Z(n10205) );
  XOR U10215 ( .A(n10206), .B(n10207), .Z(n10203) );
  AND U10216 ( .A(n10208), .B(n10209), .Z(n10206) );
  XNOR U10217 ( .A(x[8]), .B(n10207), .Z(n10209) );
  XOR U10218 ( .A(n10210), .B(n10211), .Z(n10207) );
  AND U10219 ( .A(n10212), .B(n10213), .Z(n10210) );
  XNOR U10220 ( .A(x[7]), .B(n10211), .Z(n10213) );
  XOR U10221 ( .A(n10214), .B(n10215), .Z(n10211) );
  AND U10222 ( .A(n10216), .B(n10217), .Z(n10214) );
  XNOR U10223 ( .A(x[6]), .B(n10215), .Z(n10217) );
  XOR U10224 ( .A(n10218), .B(n10219), .Z(n10215) );
  AND U10225 ( .A(n10220), .B(n10221), .Z(n10218) );
  XNOR U10226 ( .A(x[5]), .B(n10219), .Z(n10221) );
  XOR U10227 ( .A(n10222), .B(n10223), .Z(n10219) );
  AND U10228 ( .A(n10224), .B(n10225), .Z(n10222) );
  XNOR U10229 ( .A(x[4]), .B(n10223), .Z(n10225) );
  XOR U10230 ( .A(n10226), .B(n10227), .Z(n10223) );
  AND U10231 ( .A(n10228), .B(n10229), .Z(n10226) );
  XNOR U10232 ( .A(x[3]), .B(n10227), .Z(n10229) );
  XOR U10233 ( .A(n10230), .B(n10231), .Z(n10227) );
  AND U10234 ( .A(n10232), .B(n10233), .Z(n10230) );
  XNOR U10235 ( .A(x[2]), .B(n10231), .Z(n10233) );
  XOR U10236 ( .A(n10234), .B(n10235), .Z(n10231) );
  AND U10237 ( .A(n10236), .B(n10237), .Z(n10234) );
  XNOR U10238 ( .A(x[1]), .B(n10235), .Z(n10237) );
  XOR U10239 ( .A(y[1]), .B(n10235), .Z(n10236) );
  XOR U10240 ( .A(ci), .B(n10238), .Z(n10235) );
  NANDN U10241 ( .A(n10239), .B(n10240), .Z(n10238) );
  XOR U10242 ( .A(x[0]), .B(ci), .Z(n10240) );
  XOR U10243 ( .A(y[0]), .B(ci), .Z(n10239) );
endmodule

