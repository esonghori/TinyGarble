
module sum_N16384_CC32 ( clk, rst, a, b, c );
  input [511:0] a;
  input [511:0] b;
  output [511:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        carry_on) );
  XOR U4 ( .A(n2), .B(n3), .Z(carry_on_d) );
  ANDN U5 ( .B(n4), .A(n5), .Z(n2) );
  XOR U6 ( .A(b[511]), .B(n3), .Z(n4) );
  XNOR U7 ( .A(b[9]), .B(n6), .Z(c[9]) );
  XNOR U8 ( .A(b[99]), .B(n7), .Z(c[99]) );
  XNOR U9 ( .A(b[98]), .B(n8), .Z(c[98]) );
  XNOR U10 ( .A(b[97]), .B(n9), .Z(c[97]) );
  XNOR U11 ( .A(b[96]), .B(n10), .Z(c[96]) );
  XNOR U12 ( .A(b[95]), .B(n11), .Z(c[95]) );
  XNOR U13 ( .A(b[94]), .B(n12), .Z(c[94]) );
  XNOR U14 ( .A(b[93]), .B(n13), .Z(c[93]) );
  XNOR U15 ( .A(b[92]), .B(n14), .Z(c[92]) );
  XNOR U16 ( .A(b[91]), .B(n15), .Z(c[91]) );
  XNOR U17 ( .A(b[90]), .B(n16), .Z(c[90]) );
  XNOR U18 ( .A(b[8]), .B(n17), .Z(c[8]) );
  XNOR U19 ( .A(b[89]), .B(n18), .Z(c[89]) );
  XNOR U20 ( .A(b[88]), .B(n19), .Z(c[88]) );
  XNOR U21 ( .A(b[87]), .B(n20), .Z(c[87]) );
  XNOR U22 ( .A(b[86]), .B(n21), .Z(c[86]) );
  XNOR U23 ( .A(b[85]), .B(n22), .Z(c[85]) );
  XNOR U24 ( .A(b[84]), .B(n23), .Z(c[84]) );
  XNOR U25 ( .A(b[83]), .B(n24), .Z(c[83]) );
  XNOR U26 ( .A(b[82]), .B(n25), .Z(c[82]) );
  XNOR U27 ( .A(b[81]), .B(n26), .Z(c[81]) );
  XNOR U28 ( .A(b[80]), .B(n27), .Z(c[80]) );
  XNOR U29 ( .A(b[7]), .B(n28), .Z(c[7]) );
  XNOR U30 ( .A(b[79]), .B(n29), .Z(c[79]) );
  XNOR U31 ( .A(b[78]), .B(n30), .Z(c[78]) );
  XNOR U32 ( .A(b[77]), .B(n31), .Z(c[77]) );
  XNOR U33 ( .A(b[76]), .B(n32), .Z(c[76]) );
  XNOR U34 ( .A(b[75]), .B(n33), .Z(c[75]) );
  XNOR U35 ( .A(b[74]), .B(n34), .Z(c[74]) );
  XNOR U36 ( .A(b[73]), .B(n35), .Z(c[73]) );
  XNOR U37 ( .A(b[72]), .B(n36), .Z(c[72]) );
  XNOR U38 ( .A(b[71]), .B(n37), .Z(c[71]) );
  XNOR U39 ( .A(b[70]), .B(n38), .Z(c[70]) );
  XNOR U40 ( .A(b[6]), .B(n39), .Z(c[6]) );
  XNOR U41 ( .A(b[69]), .B(n40), .Z(c[69]) );
  XNOR U42 ( .A(b[68]), .B(n41), .Z(c[68]) );
  XNOR U43 ( .A(b[67]), .B(n42), .Z(c[67]) );
  XNOR U44 ( .A(b[66]), .B(n43), .Z(c[66]) );
  XNOR U45 ( .A(b[65]), .B(n44), .Z(c[65]) );
  XNOR U46 ( .A(b[64]), .B(n45), .Z(c[64]) );
  XNOR U47 ( .A(b[63]), .B(n46), .Z(c[63]) );
  XNOR U48 ( .A(b[62]), .B(n47), .Z(c[62]) );
  XNOR U49 ( .A(b[61]), .B(n48), .Z(c[61]) );
  XNOR U50 ( .A(b[60]), .B(n49), .Z(c[60]) );
  XNOR U51 ( .A(b[5]), .B(n50), .Z(c[5]) );
  XNOR U52 ( .A(b[59]), .B(n51), .Z(c[59]) );
  XNOR U53 ( .A(b[58]), .B(n52), .Z(c[58]) );
  XNOR U54 ( .A(b[57]), .B(n53), .Z(c[57]) );
  XNOR U55 ( .A(b[56]), .B(n54), .Z(c[56]) );
  XNOR U56 ( .A(b[55]), .B(n55), .Z(c[55]) );
  XNOR U57 ( .A(b[54]), .B(n56), .Z(c[54]) );
  XNOR U58 ( .A(b[53]), .B(n57), .Z(c[53]) );
  XNOR U59 ( .A(b[52]), .B(n58), .Z(c[52]) );
  XNOR U60 ( .A(b[51]), .B(n59), .Z(c[51]) );
  XNOR U61 ( .A(b[511]), .B(n5), .Z(c[511]) );
  XNOR U62 ( .A(a[511]), .B(n3), .Z(n5) );
  XNOR U63 ( .A(n60), .B(n61), .Z(n3) );
  ANDN U64 ( .B(n62), .A(n63), .Z(n60) );
  XNOR U65 ( .A(b[510]), .B(n61), .Z(n62) );
  XNOR U66 ( .A(b[510]), .B(n63), .Z(c[510]) );
  XNOR U67 ( .A(a[510]), .B(n64), .Z(n63) );
  IV U68 ( .A(n61), .Z(n64) );
  XOR U69 ( .A(n65), .B(n66), .Z(n61) );
  ANDN U70 ( .B(n67), .A(n68), .Z(n65) );
  XNOR U71 ( .A(b[509]), .B(n66), .Z(n67) );
  XNOR U72 ( .A(b[50]), .B(n69), .Z(c[50]) );
  XNOR U73 ( .A(b[509]), .B(n68), .Z(c[509]) );
  XNOR U74 ( .A(a[509]), .B(n70), .Z(n68) );
  IV U75 ( .A(n66), .Z(n70) );
  XOR U76 ( .A(n71), .B(n72), .Z(n66) );
  ANDN U77 ( .B(n73), .A(n74), .Z(n71) );
  XNOR U78 ( .A(b[508]), .B(n72), .Z(n73) );
  XNOR U79 ( .A(b[508]), .B(n74), .Z(c[508]) );
  XNOR U80 ( .A(a[508]), .B(n75), .Z(n74) );
  IV U81 ( .A(n72), .Z(n75) );
  XOR U82 ( .A(n76), .B(n77), .Z(n72) );
  ANDN U83 ( .B(n78), .A(n79), .Z(n76) );
  XNOR U84 ( .A(b[507]), .B(n77), .Z(n78) );
  XNOR U85 ( .A(b[507]), .B(n79), .Z(c[507]) );
  XNOR U86 ( .A(a[507]), .B(n80), .Z(n79) );
  IV U87 ( .A(n77), .Z(n80) );
  XOR U88 ( .A(n81), .B(n82), .Z(n77) );
  ANDN U89 ( .B(n83), .A(n84), .Z(n81) );
  XNOR U90 ( .A(b[506]), .B(n82), .Z(n83) );
  XNOR U91 ( .A(b[506]), .B(n84), .Z(c[506]) );
  XNOR U92 ( .A(a[506]), .B(n85), .Z(n84) );
  IV U93 ( .A(n82), .Z(n85) );
  XOR U94 ( .A(n86), .B(n87), .Z(n82) );
  ANDN U95 ( .B(n88), .A(n89), .Z(n86) );
  XNOR U96 ( .A(b[505]), .B(n87), .Z(n88) );
  XNOR U97 ( .A(b[505]), .B(n89), .Z(c[505]) );
  XNOR U98 ( .A(a[505]), .B(n90), .Z(n89) );
  IV U99 ( .A(n87), .Z(n90) );
  XOR U100 ( .A(n91), .B(n92), .Z(n87) );
  ANDN U101 ( .B(n93), .A(n94), .Z(n91) );
  XNOR U102 ( .A(b[504]), .B(n92), .Z(n93) );
  XNOR U103 ( .A(b[504]), .B(n94), .Z(c[504]) );
  XNOR U104 ( .A(a[504]), .B(n95), .Z(n94) );
  IV U105 ( .A(n92), .Z(n95) );
  XOR U106 ( .A(n96), .B(n97), .Z(n92) );
  ANDN U107 ( .B(n98), .A(n99), .Z(n96) );
  XNOR U108 ( .A(b[503]), .B(n97), .Z(n98) );
  XNOR U109 ( .A(b[503]), .B(n99), .Z(c[503]) );
  XNOR U110 ( .A(a[503]), .B(n100), .Z(n99) );
  IV U111 ( .A(n97), .Z(n100) );
  XOR U112 ( .A(n101), .B(n102), .Z(n97) );
  ANDN U113 ( .B(n103), .A(n104), .Z(n101) );
  XNOR U114 ( .A(b[502]), .B(n102), .Z(n103) );
  XNOR U115 ( .A(b[502]), .B(n104), .Z(c[502]) );
  XNOR U116 ( .A(a[502]), .B(n105), .Z(n104) );
  IV U117 ( .A(n102), .Z(n105) );
  XOR U118 ( .A(n106), .B(n107), .Z(n102) );
  ANDN U119 ( .B(n108), .A(n109), .Z(n106) );
  XNOR U120 ( .A(b[501]), .B(n107), .Z(n108) );
  XNOR U121 ( .A(b[501]), .B(n109), .Z(c[501]) );
  XNOR U122 ( .A(a[501]), .B(n110), .Z(n109) );
  IV U123 ( .A(n107), .Z(n110) );
  XOR U124 ( .A(n111), .B(n112), .Z(n107) );
  ANDN U125 ( .B(n113), .A(n114), .Z(n111) );
  XNOR U126 ( .A(b[500]), .B(n112), .Z(n113) );
  XNOR U127 ( .A(b[500]), .B(n114), .Z(c[500]) );
  XNOR U128 ( .A(a[500]), .B(n115), .Z(n114) );
  IV U129 ( .A(n112), .Z(n115) );
  XOR U130 ( .A(n116), .B(n117), .Z(n112) );
  ANDN U131 ( .B(n118), .A(n119), .Z(n116) );
  XNOR U132 ( .A(b[499]), .B(n117), .Z(n118) );
  XNOR U133 ( .A(b[4]), .B(n120), .Z(c[4]) );
  XNOR U134 ( .A(b[49]), .B(n121), .Z(c[49]) );
  XNOR U135 ( .A(b[499]), .B(n119), .Z(c[499]) );
  XNOR U136 ( .A(a[499]), .B(n122), .Z(n119) );
  IV U137 ( .A(n117), .Z(n122) );
  XOR U138 ( .A(n123), .B(n124), .Z(n117) );
  ANDN U139 ( .B(n125), .A(n126), .Z(n123) );
  XNOR U140 ( .A(b[498]), .B(n124), .Z(n125) );
  XNOR U141 ( .A(b[498]), .B(n126), .Z(c[498]) );
  XNOR U142 ( .A(a[498]), .B(n127), .Z(n126) );
  IV U143 ( .A(n124), .Z(n127) );
  XOR U144 ( .A(n128), .B(n129), .Z(n124) );
  ANDN U145 ( .B(n130), .A(n131), .Z(n128) );
  XNOR U146 ( .A(b[497]), .B(n129), .Z(n130) );
  XNOR U147 ( .A(b[497]), .B(n131), .Z(c[497]) );
  XNOR U148 ( .A(a[497]), .B(n132), .Z(n131) );
  IV U149 ( .A(n129), .Z(n132) );
  XOR U150 ( .A(n133), .B(n134), .Z(n129) );
  ANDN U151 ( .B(n135), .A(n136), .Z(n133) );
  XNOR U152 ( .A(b[496]), .B(n134), .Z(n135) );
  XNOR U153 ( .A(b[496]), .B(n136), .Z(c[496]) );
  XNOR U154 ( .A(a[496]), .B(n137), .Z(n136) );
  IV U155 ( .A(n134), .Z(n137) );
  XOR U156 ( .A(n138), .B(n139), .Z(n134) );
  ANDN U157 ( .B(n140), .A(n141), .Z(n138) );
  XNOR U158 ( .A(b[495]), .B(n139), .Z(n140) );
  XNOR U159 ( .A(b[495]), .B(n141), .Z(c[495]) );
  XNOR U160 ( .A(a[495]), .B(n142), .Z(n141) );
  IV U161 ( .A(n139), .Z(n142) );
  XOR U162 ( .A(n143), .B(n144), .Z(n139) );
  ANDN U163 ( .B(n145), .A(n146), .Z(n143) );
  XNOR U164 ( .A(b[494]), .B(n144), .Z(n145) );
  XNOR U165 ( .A(b[494]), .B(n146), .Z(c[494]) );
  XNOR U166 ( .A(a[494]), .B(n147), .Z(n146) );
  IV U167 ( .A(n144), .Z(n147) );
  XOR U168 ( .A(n148), .B(n149), .Z(n144) );
  ANDN U169 ( .B(n150), .A(n151), .Z(n148) );
  XNOR U170 ( .A(b[493]), .B(n149), .Z(n150) );
  XNOR U171 ( .A(b[493]), .B(n151), .Z(c[493]) );
  XNOR U172 ( .A(a[493]), .B(n152), .Z(n151) );
  IV U173 ( .A(n149), .Z(n152) );
  XOR U174 ( .A(n153), .B(n154), .Z(n149) );
  ANDN U175 ( .B(n155), .A(n156), .Z(n153) );
  XNOR U176 ( .A(b[492]), .B(n154), .Z(n155) );
  XNOR U177 ( .A(b[492]), .B(n156), .Z(c[492]) );
  XNOR U178 ( .A(a[492]), .B(n157), .Z(n156) );
  IV U179 ( .A(n154), .Z(n157) );
  XOR U180 ( .A(n158), .B(n159), .Z(n154) );
  ANDN U181 ( .B(n160), .A(n161), .Z(n158) );
  XNOR U182 ( .A(b[491]), .B(n159), .Z(n160) );
  XNOR U183 ( .A(b[491]), .B(n161), .Z(c[491]) );
  XNOR U184 ( .A(a[491]), .B(n162), .Z(n161) );
  IV U185 ( .A(n159), .Z(n162) );
  XOR U186 ( .A(n163), .B(n164), .Z(n159) );
  ANDN U187 ( .B(n165), .A(n166), .Z(n163) );
  XNOR U188 ( .A(b[490]), .B(n164), .Z(n165) );
  XNOR U189 ( .A(b[490]), .B(n166), .Z(c[490]) );
  XNOR U190 ( .A(a[490]), .B(n167), .Z(n166) );
  IV U191 ( .A(n164), .Z(n167) );
  XOR U192 ( .A(n168), .B(n169), .Z(n164) );
  ANDN U193 ( .B(n170), .A(n171), .Z(n168) );
  XNOR U194 ( .A(b[489]), .B(n169), .Z(n170) );
  XNOR U195 ( .A(b[48]), .B(n172), .Z(c[48]) );
  XNOR U196 ( .A(b[489]), .B(n171), .Z(c[489]) );
  XNOR U197 ( .A(a[489]), .B(n173), .Z(n171) );
  IV U198 ( .A(n169), .Z(n173) );
  XOR U199 ( .A(n174), .B(n175), .Z(n169) );
  ANDN U200 ( .B(n176), .A(n177), .Z(n174) );
  XNOR U201 ( .A(b[488]), .B(n175), .Z(n176) );
  XNOR U202 ( .A(b[488]), .B(n177), .Z(c[488]) );
  XNOR U203 ( .A(a[488]), .B(n178), .Z(n177) );
  IV U204 ( .A(n175), .Z(n178) );
  XOR U205 ( .A(n179), .B(n180), .Z(n175) );
  ANDN U206 ( .B(n181), .A(n182), .Z(n179) );
  XNOR U207 ( .A(b[487]), .B(n180), .Z(n181) );
  XNOR U208 ( .A(b[487]), .B(n182), .Z(c[487]) );
  XNOR U209 ( .A(a[487]), .B(n183), .Z(n182) );
  IV U210 ( .A(n180), .Z(n183) );
  XOR U211 ( .A(n184), .B(n185), .Z(n180) );
  ANDN U212 ( .B(n186), .A(n187), .Z(n184) );
  XNOR U213 ( .A(b[486]), .B(n185), .Z(n186) );
  XNOR U214 ( .A(b[486]), .B(n187), .Z(c[486]) );
  XNOR U215 ( .A(a[486]), .B(n188), .Z(n187) );
  IV U216 ( .A(n185), .Z(n188) );
  XOR U217 ( .A(n189), .B(n190), .Z(n185) );
  ANDN U218 ( .B(n191), .A(n192), .Z(n189) );
  XNOR U219 ( .A(b[485]), .B(n190), .Z(n191) );
  XNOR U220 ( .A(b[485]), .B(n192), .Z(c[485]) );
  XNOR U221 ( .A(a[485]), .B(n193), .Z(n192) );
  IV U222 ( .A(n190), .Z(n193) );
  XOR U223 ( .A(n194), .B(n195), .Z(n190) );
  ANDN U224 ( .B(n196), .A(n197), .Z(n194) );
  XNOR U225 ( .A(b[484]), .B(n195), .Z(n196) );
  XNOR U226 ( .A(b[484]), .B(n197), .Z(c[484]) );
  XNOR U227 ( .A(a[484]), .B(n198), .Z(n197) );
  IV U228 ( .A(n195), .Z(n198) );
  XOR U229 ( .A(n199), .B(n200), .Z(n195) );
  ANDN U230 ( .B(n201), .A(n202), .Z(n199) );
  XNOR U231 ( .A(b[483]), .B(n200), .Z(n201) );
  XNOR U232 ( .A(b[483]), .B(n202), .Z(c[483]) );
  XNOR U233 ( .A(a[483]), .B(n203), .Z(n202) );
  IV U234 ( .A(n200), .Z(n203) );
  XOR U235 ( .A(n204), .B(n205), .Z(n200) );
  ANDN U236 ( .B(n206), .A(n207), .Z(n204) );
  XNOR U237 ( .A(b[482]), .B(n205), .Z(n206) );
  XNOR U238 ( .A(b[482]), .B(n207), .Z(c[482]) );
  XNOR U239 ( .A(a[482]), .B(n208), .Z(n207) );
  IV U240 ( .A(n205), .Z(n208) );
  XOR U241 ( .A(n209), .B(n210), .Z(n205) );
  ANDN U242 ( .B(n211), .A(n212), .Z(n209) );
  XNOR U243 ( .A(b[481]), .B(n210), .Z(n211) );
  XNOR U244 ( .A(b[481]), .B(n212), .Z(c[481]) );
  XNOR U245 ( .A(a[481]), .B(n213), .Z(n212) );
  IV U246 ( .A(n210), .Z(n213) );
  XOR U247 ( .A(n214), .B(n215), .Z(n210) );
  ANDN U248 ( .B(n216), .A(n217), .Z(n214) );
  XNOR U249 ( .A(b[480]), .B(n215), .Z(n216) );
  XNOR U250 ( .A(b[480]), .B(n217), .Z(c[480]) );
  XNOR U251 ( .A(a[480]), .B(n218), .Z(n217) );
  IV U252 ( .A(n215), .Z(n218) );
  XOR U253 ( .A(n219), .B(n220), .Z(n215) );
  ANDN U254 ( .B(n221), .A(n222), .Z(n219) );
  XNOR U255 ( .A(b[479]), .B(n220), .Z(n221) );
  XNOR U256 ( .A(b[47]), .B(n223), .Z(c[47]) );
  XNOR U257 ( .A(b[479]), .B(n222), .Z(c[479]) );
  XNOR U258 ( .A(a[479]), .B(n224), .Z(n222) );
  IV U259 ( .A(n220), .Z(n224) );
  XOR U260 ( .A(n225), .B(n226), .Z(n220) );
  ANDN U261 ( .B(n227), .A(n228), .Z(n225) );
  XNOR U262 ( .A(b[478]), .B(n226), .Z(n227) );
  XNOR U263 ( .A(b[478]), .B(n228), .Z(c[478]) );
  XNOR U264 ( .A(a[478]), .B(n229), .Z(n228) );
  IV U265 ( .A(n226), .Z(n229) );
  XOR U266 ( .A(n230), .B(n231), .Z(n226) );
  ANDN U267 ( .B(n232), .A(n233), .Z(n230) );
  XNOR U268 ( .A(b[477]), .B(n231), .Z(n232) );
  XNOR U269 ( .A(b[477]), .B(n233), .Z(c[477]) );
  XNOR U270 ( .A(a[477]), .B(n234), .Z(n233) );
  IV U271 ( .A(n231), .Z(n234) );
  XOR U272 ( .A(n235), .B(n236), .Z(n231) );
  ANDN U273 ( .B(n237), .A(n238), .Z(n235) );
  XNOR U274 ( .A(b[476]), .B(n236), .Z(n237) );
  XNOR U275 ( .A(b[476]), .B(n238), .Z(c[476]) );
  XNOR U276 ( .A(a[476]), .B(n239), .Z(n238) );
  IV U277 ( .A(n236), .Z(n239) );
  XOR U278 ( .A(n240), .B(n241), .Z(n236) );
  ANDN U279 ( .B(n242), .A(n243), .Z(n240) );
  XNOR U280 ( .A(b[475]), .B(n241), .Z(n242) );
  XNOR U281 ( .A(b[475]), .B(n243), .Z(c[475]) );
  XNOR U282 ( .A(a[475]), .B(n244), .Z(n243) );
  IV U283 ( .A(n241), .Z(n244) );
  XOR U284 ( .A(n245), .B(n246), .Z(n241) );
  ANDN U285 ( .B(n247), .A(n248), .Z(n245) );
  XNOR U286 ( .A(b[474]), .B(n246), .Z(n247) );
  XNOR U287 ( .A(b[474]), .B(n248), .Z(c[474]) );
  XNOR U288 ( .A(a[474]), .B(n249), .Z(n248) );
  IV U289 ( .A(n246), .Z(n249) );
  XOR U290 ( .A(n250), .B(n251), .Z(n246) );
  ANDN U291 ( .B(n252), .A(n253), .Z(n250) );
  XNOR U292 ( .A(b[473]), .B(n251), .Z(n252) );
  XNOR U293 ( .A(b[473]), .B(n253), .Z(c[473]) );
  XNOR U294 ( .A(a[473]), .B(n254), .Z(n253) );
  IV U295 ( .A(n251), .Z(n254) );
  XOR U296 ( .A(n255), .B(n256), .Z(n251) );
  ANDN U297 ( .B(n257), .A(n258), .Z(n255) );
  XNOR U298 ( .A(b[472]), .B(n256), .Z(n257) );
  XNOR U299 ( .A(b[472]), .B(n258), .Z(c[472]) );
  XNOR U300 ( .A(a[472]), .B(n259), .Z(n258) );
  IV U301 ( .A(n256), .Z(n259) );
  XOR U302 ( .A(n260), .B(n261), .Z(n256) );
  ANDN U303 ( .B(n262), .A(n263), .Z(n260) );
  XNOR U304 ( .A(b[471]), .B(n261), .Z(n262) );
  XNOR U305 ( .A(b[471]), .B(n263), .Z(c[471]) );
  XNOR U306 ( .A(a[471]), .B(n264), .Z(n263) );
  IV U307 ( .A(n261), .Z(n264) );
  XOR U308 ( .A(n265), .B(n266), .Z(n261) );
  ANDN U309 ( .B(n267), .A(n268), .Z(n265) );
  XNOR U310 ( .A(b[470]), .B(n266), .Z(n267) );
  XNOR U311 ( .A(b[470]), .B(n268), .Z(c[470]) );
  XNOR U312 ( .A(a[470]), .B(n269), .Z(n268) );
  IV U313 ( .A(n266), .Z(n269) );
  XOR U314 ( .A(n270), .B(n271), .Z(n266) );
  ANDN U315 ( .B(n272), .A(n273), .Z(n270) );
  XNOR U316 ( .A(b[469]), .B(n271), .Z(n272) );
  XNOR U317 ( .A(b[46]), .B(n274), .Z(c[46]) );
  XNOR U318 ( .A(b[469]), .B(n273), .Z(c[469]) );
  XNOR U319 ( .A(a[469]), .B(n275), .Z(n273) );
  IV U320 ( .A(n271), .Z(n275) );
  XOR U321 ( .A(n276), .B(n277), .Z(n271) );
  ANDN U322 ( .B(n278), .A(n279), .Z(n276) );
  XNOR U323 ( .A(b[468]), .B(n277), .Z(n278) );
  XNOR U324 ( .A(b[468]), .B(n279), .Z(c[468]) );
  XNOR U325 ( .A(a[468]), .B(n280), .Z(n279) );
  IV U326 ( .A(n277), .Z(n280) );
  XOR U327 ( .A(n281), .B(n282), .Z(n277) );
  ANDN U328 ( .B(n283), .A(n284), .Z(n281) );
  XNOR U329 ( .A(b[467]), .B(n282), .Z(n283) );
  XNOR U330 ( .A(b[467]), .B(n284), .Z(c[467]) );
  XNOR U331 ( .A(a[467]), .B(n285), .Z(n284) );
  IV U332 ( .A(n282), .Z(n285) );
  XOR U333 ( .A(n286), .B(n287), .Z(n282) );
  ANDN U334 ( .B(n288), .A(n289), .Z(n286) );
  XNOR U335 ( .A(b[466]), .B(n287), .Z(n288) );
  XNOR U336 ( .A(b[466]), .B(n289), .Z(c[466]) );
  XNOR U337 ( .A(a[466]), .B(n290), .Z(n289) );
  IV U338 ( .A(n287), .Z(n290) );
  XOR U339 ( .A(n291), .B(n292), .Z(n287) );
  ANDN U340 ( .B(n293), .A(n294), .Z(n291) );
  XNOR U341 ( .A(b[465]), .B(n292), .Z(n293) );
  XNOR U342 ( .A(b[465]), .B(n294), .Z(c[465]) );
  XNOR U343 ( .A(a[465]), .B(n295), .Z(n294) );
  IV U344 ( .A(n292), .Z(n295) );
  XOR U345 ( .A(n296), .B(n297), .Z(n292) );
  ANDN U346 ( .B(n298), .A(n299), .Z(n296) );
  XNOR U347 ( .A(b[464]), .B(n297), .Z(n298) );
  XNOR U348 ( .A(b[464]), .B(n299), .Z(c[464]) );
  XNOR U349 ( .A(a[464]), .B(n300), .Z(n299) );
  IV U350 ( .A(n297), .Z(n300) );
  XOR U351 ( .A(n301), .B(n302), .Z(n297) );
  ANDN U352 ( .B(n303), .A(n304), .Z(n301) );
  XNOR U353 ( .A(b[463]), .B(n302), .Z(n303) );
  XNOR U354 ( .A(b[463]), .B(n304), .Z(c[463]) );
  XNOR U355 ( .A(a[463]), .B(n305), .Z(n304) );
  IV U356 ( .A(n302), .Z(n305) );
  XOR U357 ( .A(n306), .B(n307), .Z(n302) );
  ANDN U358 ( .B(n308), .A(n309), .Z(n306) );
  XNOR U359 ( .A(b[462]), .B(n307), .Z(n308) );
  XNOR U360 ( .A(b[462]), .B(n309), .Z(c[462]) );
  XNOR U361 ( .A(a[462]), .B(n310), .Z(n309) );
  IV U362 ( .A(n307), .Z(n310) );
  XOR U363 ( .A(n311), .B(n312), .Z(n307) );
  ANDN U364 ( .B(n313), .A(n314), .Z(n311) );
  XNOR U365 ( .A(b[461]), .B(n312), .Z(n313) );
  XNOR U366 ( .A(b[461]), .B(n314), .Z(c[461]) );
  XNOR U367 ( .A(a[461]), .B(n315), .Z(n314) );
  IV U368 ( .A(n312), .Z(n315) );
  XOR U369 ( .A(n316), .B(n317), .Z(n312) );
  ANDN U370 ( .B(n318), .A(n319), .Z(n316) );
  XNOR U371 ( .A(b[460]), .B(n317), .Z(n318) );
  XNOR U372 ( .A(b[460]), .B(n319), .Z(c[460]) );
  XNOR U373 ( .A(a[460]), .B(n320), .Z(n319) );
  IV U374 ( .A(n317), .Z(n320) );
  XOR U375 ( .A(n321), .B(n322), .Z(n317) );
  ANDN U376 ( .B(n323), .A(n324), .Z(n321) );
  XNOR U377 ( .A(b[459]), .B(n322), .Z(n323) );
  XNOR U378 ( .A(b[45]), .B(n325), .Z(c[45]) );
  XNOR U379 ( .A(b[459]), .B(n324), .Z(c[459]) );
  XNOR U380 ( .A(a[459]), .B(n326), .Z(n324) );
  IV U381 ( .A(n322), .Z(n326) );
  XOR U382 ( .A(n327), .B(n328), .Z(n322) );
  ANDN U383 ( .B(n329), .A(n330), .Z(n327) );
  XNOR U384 ( .A(b[458]), .B(n328), .Z(n329) );
  XNOR U385 ( .A(b[458]), .B(n330), .Z(c[458]) );
  XNOR U386 ( .A(a[458]), .B(n331), .Z(n330) );
  IV U387 ( .A(n328), .Z(n331) );
  XOR U388 ( .A(n332), .B(n333), .Z(n328) );
  ANDN U389 ( .B(n334), .A(n335), .Z(n332) );
  XNOR U390 ( .A(b[457]), .B(n333), .Z(n334) );
  XNOR U391 ( .A(b[457]), .B(n335), .Z(c[457]) );
  XNOR U392 ( .A(a[457]), .B(n336), .Z(n335) );
  IV U393 ( .A(n333), .Z(n336) );
  XOR U394 ( .A(n337), .B(n338), .Z(n333) );
  ANDN U395 ( .B(n339), .A(n340), .Z(n337) );
  XNOR U396 ( .A(b[456]), .B(n338), .Z(n339) );
  XNOR U397 ( .A(b[456]), .B(n340), .Z(c[456]) );
  XNOR U398 ( .A(a[456]), .B(n341), .Z(n340) );
  IV U399 ( .A(n338), .Z(n341) );
  XOR U400 ( .A(n342), .B(n343), .Z(n338) );
  ANDN U401 ( .B(n344), .A(n345), .Z(n342) );
  XNOR U402 ( .A(b[455]), .B(n343), .Z(n344) );
  XNOR U403 ( .A(b[455]), .B(n345), .Z(c[455]) );
  XNOR U404 ( .A(a[455]), .B(n346), .Z(n345) );
  IV U405 ( .A(n343), .Z(n346) );
  XOR U406 ( .A(n347), .B(n348), .Z(n343) );
  ANDN U407 ( .B(n349), .A(n350), .Z(n347) );
  XNOR U408 ( .A(b[454]), .B(n348), .Z(n349) );
  XNOR U409 ( .A(b[454]), .B(n350), .Z(c[454]) );
  XNOR U410 ( .A(a[454]), .B(n351), .Z(n350) );
  IV U411 ( .A(n348), .Z(n351) );
  XOR U412 ( .A(n352), .B(n353), .Z(n348) );
  ANDN U413 ( .B(n354), .A(n355), .Z(n352) );
  XNOR U414 ( .A(b[453]), .B(n353), .Z(n354) );
  XNOR U415 ( .A(b[453]), .B(n355), .Z(c[453]) );
  XNOR U416 ( .A(a[453]), .B(n356), .Z(n355) );
  IV U417 ( .A(n353), .Z(n356) );
  XOR U418 ( .A(n357), .B(n358), .Z(n353) );
  ANDN U419 ( .B(n359), .A(n360), .Z(n357) );
  XNOR U420 ( .A(b[452]), .B(n358), .Z(n359) );
  XNOR U421 ( .A(b[452]), .B(n360), .Z(c[452]) );
  XNOR U422 ( .A(a[452]), .B(n361), .Z(n360) );
  IV U423 ( .A(n358), .Z(n361) );
  XOR U424 ( .A(n362), .B(n363), .Z(n358) );
  ANDN U425 ( .B(n364), .A(n365), .Z(n362) );
  XNOR U426 ( .A(b[451]), .B(n363), .Z(n364) );
  XNOR U427 ( .A(b[451]), .B(n365), .Z(c[451]) );
  XNOR U428 ( .A(a[451]), .B(n366), .Z(n365) );
  IV U429 ( .A(n363), .Z(n366) );
  XOR U430 ( .A(n367), .B(n368), .Z(n363) );
  ANDN U431 ( .B(n369), .A(n370), .Z(n367) );
  XNOR U432 ( .A(b[450]), .B(n368), .Z(n369) );
  XNOR U433 ( .A(b[450]), .B(n370), .Z(c[450]) );
  XNOR U434 ( .A(a[450]), .B(n371), .Z(n370) );
  IV U435 ( .A(n368), .Z(n371) );
  XOR U436 ( .A(n372), .B(n373), .Z(n368) );
  ANDN U437 ( .B(n374), .A(n375), .Z(n372) );
  XNOR U438 ( .A(b[449]), .B(n373), .Z(n374) );
  XNOR U439 ( .A(b[44]), .B(n376), .Z(c[44]) );
  XNOR U440 ( .A(b[449]), .B(n375), .Z(c[449]) );
  XNOR U441 ( .A(a[449]), .B(n377), .Z(n375) );
  IV U442 ( .A(n373), .Z(n377) );
  XOR U443 ( .A(n378), .B(n379), .Z(n373) );
  ANDN U444 ( .B(n380), .A(n381), .Z(n378) );
  XNOR U445 ( .A(b[448]), .B(n379), .Z(n380) );
  XNOR U446 ( .A(b[448]), .B(n381), .Z(c[448]) );
  XNOR U447 ( .A(a[448]), .B(n382), .Z(n381) );
  IV U448 ( .A(n379), .Z(n382) );
  XOR U449 ( .A(n383), .B(n384), .Z(n379) );
  ANDN U450 ( .B(n385), .A(n386), .Z(n383) );
  XNOR U451 ( .A(b[447]), .B(n384), .Z(n385) );
  XNOR U452 ( .A(b[447]), .B(n386), .Z(c[447]) );
  XNOR U453 ( .A(a[447]), .B(n387), .Z(n386) );
  IV U454 ( .A(n384), .Z(n387) );
  XOR U455 ( .A(n388), .B(n389), .Z(n384) );
  ANDN U456 ( .B(n390), .A(n391), .Z(n388) );
  XNOR U457 ( .A(b[446]), .B(n389), .Z(n390) );
  XNOR U458 ( .A(b[446]), .B(n391), .Z(c[446]) );
  XNOR U459 ( .A(a[446]), .B(n392), .Z(n391) );
  IV U460 ( .A(n389), .Z(n392) );
  XOR U461 ( .A(n393), .B(n394), .Z(n389) );
  ANDN U462 ( .B(n395), .A(n396), .Z(n393) );
  XNOR U463 ( .A(b[445]), .B(n394), .Z(n395) );
  XNOR U464 ( .A(b[445]), .B(n396), .Z(c[445]) );
  XNOR U465 ( .A(a[445]), .B(n397), .Z(n396) );
  IV U466 ( .A(n394), .Z(n397) );
  XOR U467 ( .A(n398), .B(n399), .Z(n394) );
  ANDN U468 ( .B(n400), .A(n401), .Z(n398) );
  XNOR U469 ( .A(b[444]), .B(n399), .Z(n400) );
  XNOR U470 ( .A(b[444]), .B(n401), .Z(c[444]) );
  XNOR U471 ( .A(a[444]), .B(n402), .Z(n401) );
  IV U472 ( .A(n399), .Z(n402) );
  XOR U473 ( .A(n403), .B(n404), .Z(n399) );
  ANDN U474 ( .B(n405), .A(n406), .Z(n403) );
  XNOR U475 ( .A(b[443]), .B(n404), .Z(n405) );
  XNOR U476 ( .A(b[443]), .B(n406), .Z(c[443]) );
  XNOR U477 ( .A(a[443]), .B(n407), .Z(n406) );
  IV U478 ( .A(n404), .Z(n407) );
  XOR U479 ( .A(n408), .B(n409), .Z(n404) );
  ANDN U480 ( .B(n410), .A(n411), .Z(n408) );
  XNOR U481 ( .A(b[442]), .B(n409), .Z(n410) );
  XNOR U482 ( .A(b[442]), .B(n411), .Z(c[442]) );
  XNOR U483 ( .A(a[442]), .B(n412), .Z(n411) );
  IV U484 ( .A(n409), .Z(n412) );
  XOR U485 ( .A(n413), .B(n414), .Z(n409) );
  ANDN U486 ( .B(n415), .A(n416), .Z(n413) );
  XNOR U487 ( .A(b[441]), .B(n414), .Z(n415) );
  XNOR U488 ( .A(b[441]), .B(n416), .Z(c[441]) );
  XNOR U489 ( .A(a[441]), .B(n417), .Z(n416) );
  IV U490 ( .A(n414), .Z(n417) );
  XOR U491 ( .A(n418), .B(n419), .Z(n414) );
  ANDN U492 ( .B(n420), .A(n421), .Z(n418) );
  XNOR U493 ( .A(b[440]), .B(n419), .Z(n420) );
  XNOR U494 ( .A(b[440]), .B(n421), .Z(c[440]) );
  XNOR U495 ( .A(a[440]), .B(n422), .Z(n421) );
  IV U496 ( .A(n419), .Z(n422) );
  XOR U497 ( .A(n423), .B(n424), .Z(n419) );
  ANDN U498 ( .B(n425), .A(n426), .Z(n423) );
  XNOR U499 ( .A(b[439]), .B(n424), .Z(n425) );
  XNOR U500 ( .A(b[43]), .B(n427), .Z(c[43]) );
  XNOR U501 ( .A(b[439]), .B(n426), .Z(c[439]) );
  XNOR U502 ( .A(a[439]), .B(n428), .Z(n426) );
  IV U503 ( .A(n424), .Z(n428) );
  XOR U504 ( .A(n429), .B(n430), .Z(n424) );
  ANDN U505 ( .B(n431), .A(n432), .Z(n429) );
  XNOR U506 ( .A(b[438]), .B(n430), .Z(n431) );
  XNOR U507 ( .A(b[438]), .B(n432), .Z(c[438]) );
  XNOR U508 ( .A(a[438]), .B(n433), .Z(n432) );
  IV U509 ( .A(n430), .Z(n433) );
  XOR U510 ( .A(n434), .B(n435), .Z(n430) );
  ANDN U511 ( .B(n436), .A(n437), .Z(n434) );
  XNOR U512 ( .A(b[437]), .B(n435), .Z(n436) );
  XNOR U513 ( .A(b[437]), .B(n437), .Z(c[437]) );
  XNOR U514 ( .A(a[437]), .B(n438), .Z(n437) );
  IV U515 ( .A(n435), .Z(n438) );
  XOR U516 ( .A(n439), .B(n440), .Z(n435) );
  ANDN U517 ( .B(n441), .A(n442), .Z(n439) );
  XNOR U518 ( .A(b[436]), .B(n440), .Z(n441) );
  XNOR U519 ( .A(b[436]), .B(n442), .Z(c[436]) );
  XNOR U520 ( .A(a[436]), .B(n443), .Z(n442) );
  IV U521 ( .A(n440), .Z(n443) );
  XOR U522 ( .A(n444), .B(n445), .Z(n440) );
  ANDN U523 ( .B(n446), .A(n447), .Z(n444) );
  XNOR U524 ( .A(b[435]), .B(n445), .Z(n446) );
  XNOR U525 ( .A(b[435]), .B(n447), .Z(c[435]) );
  XNOR U526 ( .A(a[435]), .B(n448), .Z(n447) );
  IV U527 ( .A(n445), .Z(n448) );
  XOR U528 ( .A(n449), .B(n450), .Z(n445) );
  ANDN U529 ( .B(n451), .A(n452), .Z(n449) );
  XNOR U530 ( .A(b[434]), .B(n450), .Z(n451) );
  XNOR U531 ( .A(b[434]), .B(n452), .Z(c[434]) );
  XNOR U532 ( .A(a[434]), .B(n453), .Z(n452) );
  IV U533 ( .A(n450), .Z(n453) );
  XOR U534 ( .A(n454), .B(n455), .Z(n450) );
  ANDN U535 ( .B(n456), .A(n457), .Z(n454) );
  XNOR U536 ( .A(b[433]), .B(n455), .Z(n456) );
  XNOR U537 ( .A(b[433]), .B(n457), .Z(c[433]) );
  XNOR U538 ( .A(a[433]), .B(n458), .Z(n457) );
  IV U539 ( .A(n455), .Z(n458) );
  XOR U540 ( .A(n459), .B(n460), .Z(n455) );
  ANDN U541 ( .B(n461), .A(n462), .Z(n459) );
  XNOR U542 ( .A(b[432]), .B(n460), .Z(n461) );
  XNOR U543 ( .A(b[432]), .B(n462), .Z(c[432]) );
  XNOR U544 ( .A(a[432]), .B(n463), .Z(n462) );
  IV U545 ( .A(n460), .Z(n463) );
  XOR U546 ( .A(n464), .B(n465), .Z(n460) );
  ANDN U547 ( .B(n466), .A(n467), .Z(n464) );
  XNOR U548 ( .A(b[431]), .B(n465), .Z(n466) );
  XNOR U549 ( .A(b[431]), .B(n467), .Z(c[431]) );
  XNOR U550 ( .A(a[431]), .B(n468), .Z(n467) );
  IV U551 ( .A(n465), .Z(n468) );
  XOR U552 ( .A(n469), .B(n470), .Z(n465) );
  ANDN U553 ( .B(n471), .A(n472), .Z(n469) );
  XNOR U554 ( .A(b[430]), .B(n470), .Z(n471) );
  XNOR U555 ( .A(b[430]), .B(n472), .Z(c[430]) );
  XNOR U556 ( .A(a[430]), .B(n473), .Z(n472) );
  IV U557 ( .A(n470), .Z(n473) );
  XOR U558 ( .A(n474), .B(n475), .Z(n470) );
  ANDN U559 ( .B(n476), .A(n477), .Z(n474) );
  XNOR U560 ( .A(b[429]), .B(n475), .Z(n476) );
  XNOR U561 ( .A(b[42]), .B(n478), .Z(c[42]) );
  XNOR U562 ( .A(b[429]), .B(n477), .Z(c[429]) );
  XNOR U563 ( .A(a[429]), .B(n479), .Z(n477) );
  IV U564 ( .A(n475), .Z(n479) );
  XOR U565 ( .A(n480), .B(n481), .Z(n475) );
  ANDN U566 ( .B(n482), .A(n483), .Z(n480) );
  XNOR U567 ( .A(b[428]), .B(n481), .Z(n482) );
  XNOR U568 ( .A(b[428]), .B(n483), .Z(c[428]) );
  XNOR U569 ( .A(a[428]), .B(n484), .Z(n483) );
  IV U570 ( .A(n481), .Z(n484) );
  XOR U571 ( .A(n485), .B(n486), .Z(n481) );
  ANDN U572 ( .B(n487), .A(n488), .Z(n485) );
  XNOR U573 ( .A(b[427]), .B(n486), .Z(n487) );
  XNOR U574 ( .A(b[427]), .B(n488), .Z(c[427]) );
  XNOR U575 ( .A(a[427]), .B(n489), .Z(n488) );
  IV U576 ( .A(n486), .Z(n489) );
  XOR U577 ( .A(n490), .B(n491), .Z(n486) );
  ANDN U578 ( .B(n492), .A(n493), .Z(n490) );
  XNOR U579 ( .A(b[426]), .B(n491), .Z(n492) );
  XNOR U580 ( .A(b[426]), .B(n493), .Z(c[426]) );
  XNOR U581 ( .A(a[426]), .B(n494), .Z(n493) );
  IV U582 ( .A(n491), .Z(n494) );
  XOR U583 ( .A(n495), .B(n496), .Z(n491) );
  ANDN U584 ( .B(n497), .A(n498), .Z(n495) );
  XNOR U585 ( .A(b[425]), .B(n496), .Z(n497) );
  XNOR U586 ( .A(b[425]), .B(n498), .Z(c[425]) );
  XNOR U587 ( .A(a[425]), .B(n499), .Z(n498) );
  IV U588 ( .A(n496), .Z(n499) );
  XOR U589 ( .A(n500), .B(n501), .Z(n496) );
  ANDN U590 ( .B(n502), .A(n503), .Z(n500) );
  XNOR U591 ( .A(b[424]), .B(n501), .Z(n502) );
  XNOR U592 ( .A(b[424]), .B(n503), .Z(c[424]) );
  XNOR U593 ( .A(a[424]), .B(n504), .Z(n503) );
  IV U594 ( .A(n501), .Z(n504) );
  XOR U595 ( .A(n505), .B(n506), .Z(n501) );
  ANDN U596 ( .B(n507), .A(n508), .Z(n505) );
  XNOR U597 ( .A(b[423]), .B(n506), .Z(n507) );
  XNOR U598 ( .A(b[423]), .B(n508), .Z(c[423]) );
  XNOR U599 ( .A(a[423]), .B(n509), .Z(n508) );
  IV U600 ( .A(n506), .Z(n509) );
  XOR U601 ( .A(n510), .B(n511), .Z(n506) );
  ANDN U602 ( .B(n512), .A(n513), .Z(n510) );
  XNOR U603 ( .A(b[422]), .B(n511), .Z(n512) );
  XNOR U604 ( .A(b[422]), .B(n513), .Z(c[422]) );
  XNOR U605 ( .A(a[422]), .B(n514), .Z(n513) );
  IV U606 ( .A(n511), .Z(n514) );
  XOR U607 ( .A(n515), .B(n516), .Z(n511) );
  ANDN U608 ( .B(n517), .A(n518), .Z(n515) );
  XNOR U609 ( .A(b[421]), .B(n516), .Z(n517) );
  XNOR U610 ( .A(b[421]), .B(n518), .Z(c[421]) );
  XNOR U611 ( .A(a[421]), .B(n519), .Z(n518) );
  IV U612 ( .A(n516), .Z(n519) );
  XOR U613 ( .A(n520), .B(n521), .Z(n516) );
  ANDN U614 ( .B(n522), .A(n523), .Z(n520) );
  XNOR U615 ( .A(b[420]), .B(n521), .Z(n522) );
  XNOR U616 ( .A(b[420]), .B(n523), .Z(c[420]) );
  XNOR U617 ( .A(a[420]), .B(n524), .Z(n523) );
  IV U618 ( .A(n521), .Z(n524) );
  XOR U619 ( .A(n525), .B(n526), .Z(n521) );
  ANDN U620 ( .B(n527), .A(n528), .Z(n525) );
  XNOR U621 ( .A(b[419]), .B(n526), .Z(n527) );
  XNOR U622 ( .A(b[41]), .B(n529), .Z(c[41]) );
  XNOR U623 ( .A(b[419]), .B(n528), .Z(c[419]) );
  XNOR U624 ( .A(a[419]), .B(n530), .Z(n528) );
  IV U625 ( .A(n526), .Z(n530) );
  XOR U626 ( .A(n531), .B(n532), .Z(n526) );
  ANDN U627 ( .B(n533), .A(n534), .Z(n531) );
  XNOR U628 ( .A(b[418]), .B(n532), .Z(n533) );
  XNOR U629 ( .A(b[418]), .B(n534), .Z(c[418]) );
  XNOR U630 ( .A(a[418]), .B(n535), .Z(n534) );
  IV U631 ( .A(n532), .Z(n535) );
  XOR U632 ( .A(n536), .B(n537), .Z(n532) );
  ANDN U633 ( .B(n538), .A(n539), .Z(n536) );
  XNOR U634 ( .A(b[417]), .B(n537), .Z(n538) );
  XNOR U635 ( .A(b[417]), .B(n539), .Z(c[417]) );
  XNOR U636 ( .A(a[417]), .B(n540), .Z(n539) );
  IV U637 ( .A(n537), .Z(n540) );
  XOR U638 ( .A(n541), .B(n542), .Z(n537) );
  ANDN U639 ( .B(n543), .A(n544), .Z(n541) );
  XNOR U640 ( .A(b[416]), .B(n542), .Z(n543) );
  XNOR U641 ( .A(b[416]), .B(n544), .Z(c[416]) );
  XNOR U642 ( .A(a[416]), .B(n545), .Z(n544) );
  IV U643 ( .A(n542), .Z(n545) );
  XOR U644 ( .A(n546), .B(n547), .Z(n542) );
  ANDN U645 ( .B(n548), .A(n549), .Z(n546) );
  XNOR U646 ( .A(b[415]), .B(n547), .Z(n548) );
  XNOR U647 ( .A(b[415]), .B(n549), .Z(c[415]) );
  XNOR U648 ( .A(a[415]), .B(n550), .Z(n549) );
  IV U649 ( .A(n547), .Z(n550) );
  XOR U650 ( .A(n551), .B(n552), .Z(n547) );
  ANDN U651 ( .B(n553), .A(n554), .Z(n551) );
  XNOR U652 ( .A(b[414]), .B(n552), .Z(n553) );
  XNOR U653 ( .A(b[414]), .B(n554), .Z(c[414]) );
  XNOR U654 ( .A(a[414]), .B(n555), .Z(n554) );
  IV U655 ( .A(n552), .Z(n555) );
  XOR U656 ( .A(n556), .B(n557), .Z(n552) );
  ANDN U657 ( .B(n558), .A(n559), .Z(n556) );
  XNOR U658 ( .A(b[413]), .B(n557), .Z(n558) );
  XNOR U659 ( .A(b[413]), .B(n559), .Z(c[413]) );
  XNOR U660 ( .A(a[413]), .B(n560), .Z(n559) );
  IV U661 ( .A(n557), .Z(n560) );
  XOR U662 ( .A(n561), .B(n562), .Z(n557) );
  ANDN U663 ( .B(n563), .A(n564), .Z(n561) );
  XNOR U664 ( .A(b[412]), .B(n562), .Z(n563) );
  XNOR U665 ( .A(b[412]), .B(n564), .Z(c[412]) );
  XNOR U666 ( .A(a[412]), .B(n565), .Z(n564) );
  IV U667 ( .A(n562), .Z(n565) );
  XOR U668 ( .A(n566), .B(n567), .Z(n562) );
  ANDN U669 ( .B(n568), .A(n569), .Z(n566) );
  XNOR U670 ( .A(b[411]), .B(n567), .Z(n568) );
  XNOR U671 ( .A(b[411]), .B(n569), .Z(c[411]) );
  XNOR U672 ( .A(a[411]), .B(n570), .Z(n569) );
  IV U673 ( .A(n567), .Z(n570) );
  XOR U674 ( .A(n571), .B(n572), .Z(n567) );
  ANDN U675 ( .B(n573), .A(n574), .Z(n571) );
  XNOR U676 ( .A(b[410]), .B(n572), .Z(n573) );
  XNOR U677 ( .A(b[410]), .B(n574), .Z(c[410]) );
  XNOR U678 ( .A(a[410]), .B(n575), .Z(n574) );
  IV U679 ( .A(n572), .Z(n575) );
  XOR U680 ( .A(n576), .B(n577), .Z(n572) );
  ANDN U681 ( .B(n578), .A(n579), .Z(n576) );
  XNOR U682 ( .A(b[409]), .B(n577), .Z(n578) );
  XNOR U683 ( .A(b[40]), .B(n580), .Z(c[40]) );
  XNOR U684 ( .A(b[409]), .B(n579), .Z(c[409]) );
  XNOR U685 ( .A(a[409]), .B(n581), .Z(n579) );
  IV U686 ( .A(n577), .Z(n581) );
  XOR U687 ( .A(n582), .B(n583), .Z(n577) );
  ANDN U688 ( .B(n584), .A(n585), .Z(n582) );
  XNOR U689 ( .A(b[408]), .B(n583), .Z(n584) );
  XNOR U690 ( .A(b[408]), .B(n585), .Z(c[408]) );
  XNOR U691 ( .A(a[408]), .B(n586), .Z(n585) );
  IV U692 ( .A(n583), .Z(n586) );
  XOR U693 ( .A(n587), .B(n588), .Z(n583) );
  ANDN U694 ( .B(n589), .A(n590), .Z(n587) );
  XNOR U695 ( .A(b[407]), .B(n588), .Z(n589) );
  XNOR U696 ( .A(b[407]), .B(n590), .Z(c[407]) );
  XNOR U697 ( .A(a[407]), .B(n591), .Z(n590) );
  IV U698 ( .A(n588), .Z(n591) );
  XOR U699 ( .A(n592), .B(n593), .Z(n588) );
  ANDN U700 ( .B(n594), .A(n595), .Z(n592) );
  XNOR U701 ( .A(b[406]), .B(n593), .Z(n594) );
  XNOR U702 ( .A(b[406]), .B(n595), .Z(c[406]) );
  XNOR U703 ( .A(a[406]), .B(n596), .Z(n595) );
  IV U704 ( .A(n593), .Z(n596) );
  XOR U705 ( .A(n597), .B(n598), .Z(n593) );
  ANDN U706 ( .B(n599), .A(n600), .Z(n597) );
  XNOR U707 ( .A(b[405]), .B(n598), .Z(n599) );
  XNOR U708 ( .A(b[405]), .B(n600), .Z(c[405]) );
  XNOR U709 ( .A(a[405]), .B(n601), .Z(n600) );
  IV U710 ( .A(n598), .Z(n601) );
  XOR U711 ( .A(n602), .B(n603), .Z(n598) );
  ANDN U712 ( .B(n604), .A(n605), .Z(n602) );
  XNOR U713 ( .A(b[404]), .B(n603), .Z(n604) );
  XNOR U714 ( .A(b[404]), .B(n605), .Z(c[404]) );
  XNOR U715 ( .A(a[404]), .B(n606), .Z(n605) );
  IV U716 ( .A(n603), .Z(n606) );
  XOR U717 ( .A(n607), .B(n608), .Z(n603) );
  ANDN U718 ( .B(n609), .A(n610), .Z(n607) );
  XNOR U719 ( .A(b[403]), .B(n608), .Z(n609) );
  XNOR U720 ( .A(b[403]), .B(n610), .Z(c[403]) );
  XNOR U721 ( .A(a[403]), .B(n611), .Z(n610) );
  IV U722 ( .A(n608), .Z(n611) );
  XOR U723 ( .A(n612), .B(n613), .Z(n608) );
  ANDN U724 ( .B(n614), .A(n615), .Z(n612) );
  XNOR U725 ( .A(b[402]), .B(n613), .Z(n614) );
  XNOR U726 ( .A(b[402]), .B(n615), .Z(c[402]) );
  XNOR U727 ( .A(a[402]), .B(n616), .Z(n615) );
  IV U728 ( .A(n613), .Z(n616) );
  XOR U729 ( .A(n617), .B(n618), .Z(n613) );
  ANDN U730 ( .B(n619), .A(n620), .Z(n617) );
  XNOR U731 ( .A(b[401]), .B(n618), .Z(n619) );
  XNOR U732 ( .A(b[401]), .B(n620), .Z(c[401]) );
  XNOR U733 ( .A(a[401]), .B(n621), .Z(n620) );
  IV U734 ( .A(n618), .Z(n621) );
  XOR U735 ( .A(n622), .B(n623), .Z(n618) );
  ANDN U736 ( .B(n624), .A(n625), .Z(n622) );
  XNOR U737 ( .A(b[400]), .B(n623), .Z(n624) );
  XNOR U738 ( .A(b[400]), .B(n625), .Z(c[400]) );
  XNOR U739 ( .A(a[400]), .B(n626), .Z(n625) );
  IV U740 ( .A(n623), .Z(n626) );
  XOR U741 ( .A(n627), .B(n628), .Z(n623) );
  ANDN U742 ( .B(n629), .A(n630), .Z(n627) );
  XNOR U743 ( .A(b[399]), .B(n628), .Z(n629) );
  XNOR U744 ( .A(b[3]), .B(n631), .Z(c[3]) );
  XNOR U745 ( .A(b[39]), .B(n632), .Z(c[39]) );
  XNOR U746 ( .A(b[399]), .B(n630), .Z(c[399]) );
  XNOR U747 ( .A(a[399]), .B(n633), .Z(n630) );
  IV U748 ( .A(n628), .Z(n633) );
  XOR U749 ( .A(n634), .B(n635), .Z(n628) );
  ANDN U750 ( .B(n636), .A(n637), .Z(n634) );
  XNOR U751 ( .A(b[398]), .B(n635), .Z(n636) );
  XNOR U752 ( .A(b[398]), .B(n637), .Z(c[398]) );
  XNOR U753 ( .A(a[398]), .B(n638), .Z(n637) );
  IV U754 ( .A(n635), .Z(n638) );
  XOR U755 ( .A(n639), .B(n640), .Z(n635) );
  ANDN U756 ( .B(n641), .A(n642), .Z(n639) );
  XNOR U757 ( .A(b[397]), .B(n640), .Z(n641) );
  XNOR U758 ( .A(b[397]), .B(n642), .Z(c[397]) );
  XNOR U759 ( .A(a[397]), .B(n643), .Z(n642) );
  IV U760 ( .A(n640), .Z(n643) );
  XOR U761 ( .A(n644), .B(n645), .Z(n640) );
  ANDN U762 ( .B(n646), .A(n647), .Z(n644) );
  XNOR U763 ( .A(b[396]), .B(n645), .Z(n646) );
  XNOR U764 ( .A(b[396]), .B(n647), .Z(c[396]) );
  XNOR U765 ( .A(a[396]), .B(n648), .Z(n647) );
  IV U766 ( .A(n645), .Z(n648) );
  XOR U767 ( .A(n649), .B(n650), .Z(n645) );
  ANDN U768 ( .B(n651), .A(n652), .Z(n649) );
  XNOR U769 ( .A(b[395]), .B(n650), .Z(n651) );
  XNOR U770 ( .A(b[395]), .B(n652), .Z(c[395]) );
  XNOR U771 ( .A(a[395]), .B(n653), .Z(n652) );
  IV U772 ( .A(n650), .Z(n653) );
  XOR U773 ( .A(n654), .B(n655), .Z(n650) );
  ANDN U774 ( .B(n656), .A(n657), .Z(n654) );
  XNOR U775 ( .A(b[394]), .B(n655), .Z(n656) );
  XNOR U776 ( .A(b[394]), .B(n657), .Z(c[394]) );
  XNOR U777 ( .A(a[394]), .B(n658), .Z(n657) );
  IV U778 ( .A(n655), .Z(n658) );
  XOR U779 ( .A(n659), .B(n660), .Z(n655) );
  ANDN U780 ( .B(n661), .A(n662), .Z(n659) );
  XNOR U781 ( .A(b[393]), .B(n660), .Z(n661) );
  XNOR U782 ( .A(b[393]), .B(n662), .Z(c[393]) );
  XNOR U783 ( .A(a[393]), .B(n663), .Z(n662) );
  IV U784 ( .A(n660), .Z(n663) );
  XOR U785 ( .A(n664), .B(n665), .Z(n660) );
  ANDN U786 ( .B(n666), .A(n667), .Z(n664) );
  XNOR U787 ( .A(b[392]), .B(n665), .Z(n666) );
  XNOR U788 ( .A(b[392]), .B(n667), .Z(c[392]) );
  XNOR U789 ( .A(a[392]), .B(n668), .Z(n667) );
  IV U790 ( .A(n665), .Z(n668) );
  XOR U791 ( .A(n669), .B(n670), .Z(n665) );
  ANDN U792 ( .B(n671), .A(n672), .Z(n669) );
  XNOR U793 ( .A(b[391]), .B(n670), .Z(n671) );
  XNOR U794 ( .A(b[391]), .B(n672), .Z(c[391]) );
  XNOR U795 ( .A(a[391]), .B(n673), .Z(n672) );
  IV U796 ( .A(n670), .Z(n673) );
  XOR U797 ( .A(n674), .B(n675), .Z(n670) );
  ANDN U798 ( .B(n676), .A(n677), .Z(n674) );
  XNOR U799 ( .A(b[390]), .B(n675), .Z(n676) );
  XNOR U800 ( .A(b[390]), .B(n677), .Z(c[390]) );
  XNOR U801 ( .A(a[390]), .B(n678), .Z(n677) );
  IV U802 ( .A(n675), .Z(n678) );
  XOR U803 ( .A(n679), .B(n680), .Z(n675) );
  ANDN U804 ( .B(n681), .A(n682), .Z(n679) );
  XNOR U805 ( .A(b[389]), .B(n680), .Z(n681) );
  XNOR U806 ( .A(b[38]), .B(n683), .Z(c[38]) );
  XNOR U807 ( .A(b[389]), .B(n682), .Z(c[389]) );
  XNOR U808 ( .A(a[389]), .B(n684), .Z(n682) );
  IV U809 ( .A(n680), .Z(n684) );
  XOR U810 ( .A(n685), .B(n686), .Z(n680) );
  ANDN U811 ( .B(n687), .A(n688), .Z(n685) );
  XNOR U812 ( .A(b[388]), .B(n686), .Z(n687) );
  XNOR U813 ( .A(b[388]), .B(n688), .Z(c[388]) );
  XNOR U814 ( .A(a[388]), .B(n689), .Z(n688) );
  IV U815 ( .A(n686), .Z(n689) );
  XOR U816 ( .A(n690), .B(n691), .Z(n686) );
  ANDN U817 ( .B(n692), .A(n693), .Z(n690) );
  XNOR U818 ( .A(b[387]), .B(n691), .Z(n692) );
  XNOR U819 ( .A(b[387]), .B(n693), .Z(c[387]) );
  XNOR U820 ( .A(a[387]), .B(n694), .Z(n693) );
  IV U821 ( .A(n691), .Z(n694) );
  XOR U822 ( .A(n695), .B(n696), .Z(n691) );
  ANDN U823 ( .B(n697), .A(n698), .Z(n695) );
  XNOR U824 ( .A(b[386]), .B(n696), .Z(n697) );
  XNOR U825 ( .A(b[386]), .B(n698), .Z(c[386]) );
  XNOR U826 ( .A(a[386]), .B(n699), .Z(n698) );
  IV U827 ( .A(n696), .Z(n699) );
  XOR U828 ( .A(n700), .B(n701), .Z(n696) );
  ANDN U829 ( .B(n702), .A(n703), .Z(n700) );
  XNOR U830 ( .A(b[385]), .B(n701), .Z(n702) );
  XNOR U831 ( .A(b[385]), .B(n703), .Z(c[385]) );
  XNOR U832 ( .A(a[385]), .B(n704), .Z(n703) );
  IV U833 ( .A(n701), .Z(n704) );
  XOR U834 ( .A(n705), .B(n706), .Z(n701) );
  ANDN U835 ( .B(n707), .A(n708), .Z(n705) );
  XNOR U836 ( .A(b[384]), .B(n706), .Z(n707) );
  XNOR U837 ( .A(b[384]), .B(n708), .Z(c[384]) );
  XNOR U838 ( .A(a[384]), .B(n709), .Z(n708) );
  IV U839 ( .A(n706), .Z(n709) );
  XOR U840 ( .A(n710), .B(n711), .Z(n706) );
  ANDN U841 ( .B(n712), .A(n713), .Z(n710) );
  XNOR U842 ( .A(b[383]), .B(n711), .Z(n712) );
  XNOR U843 ( .A(b[383]), .B(n713), .Z(c[383]) );
  XNOR U844 ( .A(a[383]), .B(n714), .Z(n713) );
  IV U845 ( .A(n711), .Z(n714) );
  XOR U846 ( .A(n715), .B(n716), .Z(n711) );
  ANDN U847 ( .B(n717), .A(n718), .Z(n715) );
  XNOR U848 ( .A(b[382]), .B(n716), .Z(n717) );
  XNOR U849 ( .A(b[382]), .B(n718), .Z(c[382]) );
  XNOR U850 ( .A(a[382]), .B(n719), .Z(n718) );
  IV U851 ( .A(n716), .Z(n719) );
  XOR U852 ( .A(n720), .B(n721), .Z(n716) );
  ANDN U853 ( .B(n722), .A(n723), .Z(n720) );
  XNOR U854 ( .A(b[381]), .B(n721), .Z(n722) );
  XNOR U855 ( .A(b[381]), .B(n723), .Z(c[381]) );
  XNOR U856 ( .A(a[381]), .B(n724), .Z(n723) );
  IV U857 ( .A(n721), .Z(n724) );
  XOR U858 ( .A(n725), .B(n726), .Z(n721) );
  ANDN U859 ( .B(n727), .A(n728), .Z(n725) );
  XNOR U860 ( .A(b[380]), .B(n726), .Z(n727) );
  XNOR U861 ( .A(b[380]), .B(n728), .Z(c[380]) );
  XNOR U862 ( .A(a[380]), .B(n729), .Z(n728) );
  IV U863 ( .A(n726), .Z(n729) );
  XOR U864 ( .A(n730), .B(n731), .Z(n726) );
  ANDN U865 ( .B(n732), .A(n733), .Z(n730) );
  XNOR U866 ( .A(b[379]), .B(n731), .Z(n732) );
  XNOR U867 ( .A(b[37]), .B(n734), .Z(c[37]) );
  XNOR U868 ( .A(b[379]), .B(n733), .Z(c[379]) );
  XNOR U869 ( .A(a[379]), .B(n735), .Z(n733) );
  IV U870 ( .A(n731), .Z(n735) );
  XOR U871 ( .A(n736), .B(n737), .Z(n731) );
  ANDN U872 ( .B(n738), .A(n739), .Z(n736) );
  XNOR U873 ( .A(b[378]), .B(n737), .Z(n738) );
  XNOR U874 ( .A(b[378]), .B(n739), .Z(c[378]) );
  XNOR U875 ( .A(a[378]), .B(n740), .Z(n739) );
  IV U876 ( .A(n737), .Z(n740) );
  XOR U877 ( .A(n741), .B(n742), .Z(n737) );
  ANDN U878 ( .B(n743), .A(n744), .Z(n741) );
  XNOR U879 ( .A(b[377]), .B(n742), .Z(n743) );
  XNOR U880 ( .A(b[377]), .B(n744), .Z(c[377]) );
  XNOR U881 ( .A(a[377]), .B(n745), .Z(n744) );
  IV U882 ( .A(n742), .Z(n745) );
  XOR U883 ( .A(n746), .B(n747), .Z(n742) );
  ANDN U884 ( .B(n748), .A(n749), .Z(n746) );
  XNOR U885 ( .A(b[376]), .B(n747), .Z(n748) );
  XNOR U886 ( .A(b[376]), .B(n749), .Z(c[376]) );
  XNOR U887 ( .A(a[376]), .B(n750), .Z(n749) );
  IV U888 ( .A(n747), .Z(n750) );
  XOR U889 ( .A(n751), .B(n752), .Z(n747) );
  ANDN U890 ( .B(n753), .A(n754), .Z(n751) );
  XNOR U891 ( .A(b[375]), .B(n752), .Z(n753) );
  XNOR U892 ( .A(b[375]), .B(n754), .Z(c[375]) );
  XNOR U893 ( .A(a[375]), .B(n755), .Z(n754) );
  IV U894 ( .A(n752), .Z(n755) );
  XOR U895 ( .A(n756), .B(n757), .Z(n752) );
  ANDN U896 ( .B(n758), .A(n759), .Z(n756) );
  XNOR U897 ( .A(b[374]), .B(n757), .Z(n758) );
  XNOR U898 ( .A(b[374]), .B(n759), .Z(c[374]) );
  XNOR U899 ( .A(a[374]), .B(n760), .Z(n759) );
  IV U900 ( .A(n757), .Z(n760) );
  XOR U901 ( .A(n761), .B(n762), .Z(n757) );
  ANDN U902 ( .B(n763), .A(n764), .Z(n761) );
  XNOR U903 ( .A(b[373]), .B(n762), .Z(n763) );
  XNOR U904 ( .A(b[373]), .B(n764), .Z(c[373]) );
  XNOR U905 ( .A(a[373]), .B(n765), .Z(n764) );
  IV U906 ( .A(n762), .Z(n765) );
  XOR U907 ( .A(n766), .B(n767), .Z(n762) );
  ANDN U908 ( .B(n768), .A(n769), .Z(n766) );
  XNOR U909 ( .A(b[372]), .B(n767), .Z(n768) );
  XNOR U910 ( .A(b[372]), .B(n769), .Z(c[372]) );
  XNOR U911 ( .A(a[372]), .B(n770), .Z(n769) );
  IV U912 ( .A(n767), .Z(n770) );
  XOR U913 ( .A(n771), .B(n772), .Z(n767) );
  ANDN U914 ( .B(n773), .A(n774), .Z(n771) );
  XNOR U915 ( .A(b[371]), .B(n772), .Z(n773) );
  XNOR U916 ( .A(b[371]), .B(n774), .Z(c[371]) );
  XNOR U917 ( .A(a[371]), .B(n775), .Z(n774) );
  IV U918 ( .A(n772), .Z(n775) );
  XOR U919 ( .A(n776), .B(n777), .Z(n772) );
  ANDN U920 ( .B(n778), .A(n779), .Z(n776) );
  XNOR U921 ( .A(b[370]), .B(n777), .Z(n778) );
  XNOR U922 ( .A(b[370]), .B(n779), .Z(c[370]) );
  XNOR U923 ( .A(a[370]), .B(n780), .Z(n779) );
  IV U924 ( .A(n777), .Z(n780) );
  XOR U925 ( .A(n781), .B(n782), .Z(n777) );
  ANDN U926 ( .B(n783), .A(n784), .Z(n781) );
  XNOR U927 ( .A(b[369]), .B(n782), .Z(n783) );
  XNOR U928 ( .A(b[36]), .B(n785), .Z(c[36]) );
  XNOR U929 ( .A(b[369]), .B(n784), .Z(c[369]) );
  XNOR U930 ( .A(a[369]), .B(n786), .Z(n784) );
  IV U931 ( .A(n782), .Z(n786) );
  XOR U932 ( .A(n787), .B(n788), .Z(n782) );
  ANDN U933 ( .B(n789), .A(n790), .Z(n787) );
  XNOR U934 ( .A(b[368]), .B(n788), .Z(n789) );
  XNOR U935 ( .A(b[368]), .B(n790), .Z(c[368]) );
  XNOR U936 ( .A(a[368]), .B(n791), .Z(n790) );
  IV U937 ( .A(n788), .Z(n791) );
  XOR U938 ( .A(n792), .B(n793), .Z(n788) );
  ANDN U939 ( .B(n794), .A(n795), .Z(n792) );
  XNOR U940 ( .A(b[367]), .B(n793), .Z(n794) );
  XNOR U941 ( .A(b[367]), .B(n795), .Z(c[367]) );
  XNOR U942 ( .A(a[367]), .B(n796), .Z(n795) );
  IV U943 ( .A(n793), .Z(n796) );
  XOR U944 ( .A(n797), .B(n798), .Z(n793) );
  ANDN U945 ( .B(n799), .A(n800), .Z(n797) );
  XNOR U946 ( .A(b[366]), .B(n798), .Z(n799) );
  XNOR U947 ( .A(b[366]), .B(n800), .Z(c[366]) );
  XNOR U948 ( .A(a[366]), .B(n801), .Z(n800) );
  IV U949 ( .A(n798), .Z(n801) );
  XOR U950 ( .A(n802), .B(n803), .Z(n798) );
  ANDN U951 ( .B(n804), .A(n805), .Z(n802) );
  XNOR U952 ( .A(b[365]), .B(n803), .Z(n804) );
  XNOR U953 ( .A(b[365]), .B(n805), .Z(c[365]) );
  XNOR U954 ( .A(a[365]), .B(n806), .Z(n805) );
  IV U955 ( .A(n803), .Z(n806) );
  XOR U956 ( .A(n807), .B(n808), .Z(n803) );
  ANDN U957 ( .B(n809), .A(n810), .Z(n807) );
  XNOR U958 ( .A(b[364]), .B(n808), .Z(n809) );
  XNOR U959 ( .A(b[364]), .B(n810), .Z(c[364]) );
  XNOR U960 ( .A(a[364]), .B(n811), .Z(n810) );
  IV U961 ( .A(n808), .Z(n811) );
  XOR U962 ( .A(n812), .B(n813), .Z(n808) );
  ANDN U963 ( .B(n814), .A(n815), .Z(n812) );
  XNOR U964 ( .A(b[363]), .B(n813), .Z(n814) );
  XNOR U965 ( .A(b[363]), .B(n815), .Z(c[363]) );
  XNOR U966 ( .A(a[363]), .B(n816), .Z(n815) );
  IV U967 ( .A(n813), .Z(n816) );
  XOR U968 ( .A(n817), .B(n818), .Z(n813) );
  ANDN U969 ( .B(n819), .A(n820), .Z(n817) );
  XNOR U970 ( .A(b[362]), .B(n818), .Z(n819) );
  XNOR U971 ( .A(b[362]), .B(n820), .Z(c[362]) );
  XNOR U972 ( .A(a[362]), .B(n821), .Z(n820) );
  IV U973 ( .A(n818), .Z(n821) );
  XOR U974 ( .A(n822), .B(n823), .Z(n818) );
  ANDN U975 ( .B(n824), .A(n825), .Z(n822) );
  XNOR U976 ( .A(b[361]), .B(n823), .Z(n824) );
  XNOR U977 ( .A(b[361]), .B(n825), .Z(c[361]) );
  XNOR U978 ( .A(a[361]), .B(n826), .Z(n825) );
  IV U979 ( .A(n823), .Z(n826) );
  XOR U980 ( .A(n827), .B(n828), .Z(n823) );
  ANDN U981 ( .B(n829), .A(n830), .Z(n827) );
  XNOR U982 ( .A(b[360]), .B(n828), .Z(n829) );
  XNOR U983 ( .A(b[360]), .B(n830), .Z(c[360]) );
  XNOR U984 ( .A(a[360]), .B(n831), .Z(n830) );
  IV U985 ( .A(n828), .Z(n831) );
  XOR U986 ( .A(n832), .B(n833), .Z(n828) );
  ANDN U987 ( .B(n834), .A(n835), .Z(n832) );
  XNOR U988 ( .A(b[359]), .B(n833), .Z(n834) );
  XNOR U989 ( .A(b[35]), .B(n836), .Z(c[35]) );
  XNOR U990 ( .A(b[359]), .B(n835), .Z(c[359]) );
  XNOR U991 ( .A(a[359]), .B(n837), .Z(n835) );
  IV U992 ( .A(n833), .Z(n837) );
  XOR U993 ( .A(n838), .B(n839), .Z(n833) );
  ANDN U994 ( .B(n840), .A(n841), .Z(n838) );
  XNOR U995 ( .A(b[358]), .B(n839), .Z(n840) );
  XNOR U996 ( .A(b[358]), .B(n841), .Z(c[358]) );
  XNOR U997 ( .A(a[358]), .B(n842), .Z(n841) );
  IV U998 ( .A(n839), .Z(n842) );
  XOR U999 ( .A(n843), .B(n844), .Z(n839) );
  ANDN U1000 ( .B(n845), .A(n846), .Z(n843) );
  XNOR U1001 ( .A(b[357]), .B(n844), .Z(n845) );
  XNOR U1002 ( .A(b[357]), .B(n846), .Z(c[357]) );
  XNOR U1003 ( .A(a[357]), .B(n847), .Z(n846) );
  IV U1004 ( .A(n844), .Z(n847) );
  XOR U1005 ( .A(n848), .B(n849), .Z(n844) );
  ANDN U1006 ( .B(n850), .A(n851), .Z(n848) );
  XNOR U1007 ( .A(b[356]), .B(n849), .Z(n850) );
  XNOR U1008 ( .A(b[356]), .B(n851), .Z(c[356]) );
  XNOR U1009 ( .A(a[356]), .B(n852), .Z(n851) );
  IV U1010 ( .A(n849), .Z(n852) );
  XOR U1011 ( .A(n853), .B(n854), .Z(n849) );
  ANDN U1012 ( .B(n855), .A(n856), .Z(n853) );
  XNOR U1013 ( .A(b[355]), .B(n854), .Z(n855) );
  XNOR U1014 ( .A(b[355]), .B(n856), .Z(c[355]) );
  XNOR U1015 ( .A(a[355]), .B(n857), .Z(n856) );
  IV U1016 ( .A(n854), .Z(n857) );
  XOR U1017 ( .A(n858), .B(n859), .Z(n854) );
  ANDN U1018 ( .B(n860), .A(n861), .Z(n858) );
  XNOR U1019 ( .A(b[354]), .B(n859), .Z(n860) );
  XNOR U1020 ( .A(b[354]), .B(n861), .Z(c[354]) );
  XNOR U1021 ( .A(a[354]), .B(n862), .Z(n861) );
  IV U1022 ( .A(n859), .Z(n862) );
  XOR U1023 ( .A(n863), .B(n864), .Z(n859) );
  ANDN U1024 ( .B(n865), .A(n866), .Z(n863) );
  XNOR U1025 ( .A(b[353]), .B(n864), .Z(n865) );
  XNOR U1026 ( .A(b[353]), .B(n866), .Z(c[353]) );
  XNOR U1027 ( .A(a[353]), .B(n867), .Z(n866) );
  IV U1028 ( .A(n864), .Z(n867) );
  XOR U1029 ( .A(n868), .B(n869), .Z(n864) );
  ANDN U1030 ( .B(n870), .A(n871), .Z(n868) );
  XNOR U1031 ( .A(b[352]), .B(n869), .Z(n870) );
  XNOR U1032 ( .A(b[352]), .B(n871), .Z(c[352]) );
  XNOR U1033 ( .A(a[352]), .B(n872), .Z(n871) );
  IV U1034 ( .A(n869), .Z(n872) );
  XOR U1035 ( .A(n873), .B(n874), .Z(n869) );
  ANDN U1036 ( .B(n875), .A(n876), .Z(n873) );
  XNOR U1037 ( .A(b[351]), .B(n874), .Z(n875) );
  XNOR U1038 ( .A(b[351]), .B(n876), .Z(c[351]) );
  XNOR U1039 ( .A(a[351]), .B(n877), .Z(n876) );
  IV U1040 ( .A(n874), .Z(n877) );
  XOR U1041 ( .A(n878), .B(n879), .Z(n874) );
  ANDN U1042 ( .B(n880), .A(n881), .Z(n878) );
  XNOR U1043 ( .A(b[350]), .B(n879), .Z(n880) );
  XNOR U1044 ( .A(b[350]), .B(n881), .Z(c[350]) );
  XNOR U1045 ( .A(a[350]), .B(n882), .Z(n881) );
  IV U1046 ( .A(n879), .Z(n882) );
  XOR U1047 ( .A(n883), .B(n884), .Z(n879) );
  ANDN U1048 ( .B(n885), .A(n886), .Z(n883) );
  XNOR U1049 ( .A(b[349]), .B(n884), .Z(n885) );
  XNOR U1050 ( .A(b[34]), .B(n887), .Z(c[34]) );
  XNOR U1051 ( .A(b[349]), .B(n886), .Z(c[349]) );
  XNOR U1052 ( .A(a[349]), .B(n888), .Z(n886) );
  IV U1053 ( .A(n884), .Z(n888) );
  XOR U1054 ( .A(n889), .B(n890), .Z(n884) );
  ANDN U1055 ( .B(n891), .A(n892), .Z(n889) );
  XNOR U1056 ( .A(b[348]), .B(n890), .Z(n891) );
  XNOR U1057 ( .A(b[348]), .B(n892), .Z(c[348]) );
  XNOR U1058 ( .A(a[348]), .B(n893), .Z(n892) );
  IV U1059 ( .A(n890), .Z(n893) );
  XOR U1060 ( .A(n894), .B(n895), .Z(n890) );
  ANDN U1061 ( .B(n896), .A(n897), .Z(n894) );
  XNOR U1062 ( .A(b[347]), .B(n895), .Z(n896) );
  XNOR U1063 ( .A(b[347]), .B(n897), .Z(c[347]) );
  XNOR U1064 ( .A(a[347]), .B(n898), .Z(n897) );
  IV U1065 ( .A(n895), .Z(n898) );
  XOR U1066 ( .A(n899), .B(n900), .Z(n895) );
  ANDN U1067 ( .B(n901), .A(n902), .Z(n899) );
  XNOR U1068 ( .A(b[346]), .B(n900), .Z(n901) );
  XNOR U1069 ( .A(b[346]), .B(n902), .Z(c[346]) );
  XNOR U1070 ( .A(a[346]), .B(n903), .Z(n902) );
  IV U1071 ( .A(n900), .Z(n903) );
  XOR U1072 ( .A(n904), .B(n905), .Z(n900) );
  ANDN U1073 ( .B(n906), .A(n907), .Z(n904) );
  XNOR U1074 ( .A(b[345]), .B(n905), .Z(n906) );
  XNOR U1075 ( .A(b[345]), .B(n907), .Z(c[345]) );
  XNOR U1076 ( .A(a[345]), .B(n908), .Z(n907) );
  IV U1077 ( .A(n905), .Z(n908) );
  XOR U1078 ( .A(n909), .B(n910), .Z(n905) );
  ANDN U1079 ( .B(n911), .A(n912), .Z(n909) );
  XNOR U1080 ( .A(b[344]), .B(n910), .Z(n911) );
  XNOR U1081 ( .A(b[344]), .B(n912), .Z(c[344]) );
  XNOR U1082 ( .A(a[344]), .B(n913), .Z(n912) );
  IV U1083 ( .A(n910), .Z(n913) );
  XOR U1084 ( .A(n914), .B(n915), .Z(n910) );
  ANDN U1085 ( .B(n916), .A(n917), .Z(n914) );
  XNOR U1086 ( .A(b[343]), .B(n915), .Z(n916) );
  XNOR U1087 ( .A(b[343]), .B(n917), .Z(c[343]) );
  XNOR U1088 ( .A(a[343]), .B(n918), .Z(n917) );
  IV U1089 ( .A(n915), .Z(n918) );
  XOR U1090 ( .A(n919), .B(n920), .Z(n915) );
  ANDN U1091 ( .B(n921), .A(n922), .Z(n919) );
  XNOR U1092 ( .A(b[342]), .B(n920), .Z(n921) );
  XNOR U1093 ( .A(b[342]), .B(n922), .Z(c[342]) );
  XNOR U1094 ( .A(a[342]), .B(n923), .Z(n922) );
  IV U1095 ( .A(n920), .Z(n923) );
  XOR U1096 ( .A(n924), .B(n925), .Z(n920) );
  ANDN U1097 ( .B(n926), .A(n927), .Z(n924) );
  XNOR U1098 ( .A(b[341]), .B(n925), .Z(n926) );
  XNOR U1099 ( .A(b[341]), .B(n927), .Z(c[341]) );
  XNOR U1100 ( .A(a[341]), .B(n928), .Z(n927) );
  IV U1101 ( .A(n925), .Z(n928) );
  XOR U1102 ( .A(n929), .B(n930), .Z(n925) );
  ANDN U1103 ( .B(n931), .A(n932), .Z(n929) );
  XNOR U1104 ( .A(b[340]), .B(n930), .Z(n931) );
  XNOR U1105 ( .A(b[340]), .B(n932), .Z(c[340]) );
  XNOR U1106 ( .A(a[340]), .B(n933), .Z(n932) );
  IV U1107 ( .A(n930), .Z(n933) );
  XOR U1108 ( .A(n934), .B(n935), .Z(n930) );
  ANDN U1109 ( .B(n936), .A(n937), .Z(n934) );
  XNOR U1110 ( .A(b[339]), .B(n935), .Z(n936) );
  XNOR U1111 ( .A(b[33]), .B(n938), .Z(c[33]) );
  XNOR U1112 ( .A(b[339]), .B(n937), .Z(c[339]) );
  XNOR U1113 ( .A(a[339]), .B(n939), .Z(n937) );
  IV U1114 ( .A(n935), .Z(n939) );
  XOR U1115 ( .A(n940), .B(n941), .Z(n935) );
  ANDN U1116 ( .B(n942), .A(n943), .Z(n940) );
  XNOR U1117 ( .A(b[338]), .B(n941), .Z(n942) );
  XNOR U1118 ( .A(b[338]), .B(n943), .Z(c[338]) );
  XNOR U1119 ( .A(a[338]), .B(n944), .Z(n943) );
  IV U1120 ( .A(n941), .Z(n944) );
  XOR U1121 ( .A(n945), .B(n946), .Z(n941) );
  ANDN U1122 ( .B(n947), .A(n948), .Z(n945) );
  XNOR U1123 ( .A(b[337]), .B(n946), .Z(n947) );
  XNOR U1124 ( .A(b[337]), .B(n948), .Z(c[337]) );
  XNOR U1125 ( .A(a[337]), .B(n949), .Z(n948) );
  IV U1126 ( .A(n946), .Z(n949) );
  XOR U1127 ( .A(n950), .B(n951), .Z(n946) );
  ANDN U1128 ( .B(n952), .A(n953), .Z(n950) );
  XNOR U1129 ( .A(b[336]), .B(n951), .Z(n952) );
  XNOR U1130 ( .A(b[336]), .B(n953), .Z(c[336]) );
  XNOR U1131 ( .A(a[336]), .B(n954), .Z(n953) );
  IV U1132 ( .A(n951), .Z(n954) );
  XOR U1133 ( .A(n955), .B(n956), .Z(n951) );
  ANDN U1134 ( .B(n957), .A(n958), .Z(n955) );
  XNOR U1135 ( .A(b[335]), .B(n956), .Z(n957) );
  XNOR U1136 ( .A(b[335]), .B(n958), .Z(c[335]) );
  XNOR U1137 ( .A(a[335]), .B(n959), .Z(n958) );
  IV U1138 ( .A(n956), .Z(n959) );
  XOR U1139 ( .A(n960), .B(n961), .Z(n956) );
  ANDN U1140 ( .B(n962), .A(n963), .Z(n960) );
  XNOR U1141 ( .A(b[334]), .B(n961), .Z(n962) );
  XNOR U1142 ( .A(b[334]), .B(n963), .Z(c[334]) );
  XNOR U1143 ( .A(a[334]), .B(n964), .Z(n963) );
  IV U1144 ( .A(n961), .Z(n964) );
  XOR U1145 ( .A(n965), .B(n966), .Z(n961) );
  ANDN U1146 ( .B(n967), .A(n968), .Z(n965) );
  XNOR U1147 ( .A(b[333]), .B(n966), .Z(n967) );
  XNOR U1148 ( .A(b[333]), .B(n968), .Z(c[333]) );
  XNOR U1149 ( .A(a[333]), .B(n969), .Z(n968) );
  IV U1150 ( .A(n966), .Z(n969) );
  XOR U1151 ( .A(n970), .B(n971), .Z(n966) );
  ANDN U1152 ( .B(n972), .A(n973), .Z(n970) );
  XNOR U1153 ( .A(b[332]), .B(n971), .Z(n972) );
  XNOR U1154 ( .A(b[332]), .B(n973), .Z(c[332]) );
  XNOR U1155 ( .A(a[332]), .B(n974), .Z(n973) );
  IV U1156 ( .A(n971), .Z(n974) );
  XOR U1157 ( .A(n975), .B(n976), .Z(n971) );
  ANDN U1158 ( .B(n977), .A(n978), .Z(n975) );
  XNOR U1159 ( .A(b[331]), .B(n976), .Z(n977) );
  XNOR U1160 ( .A(b[331]), .B(n978), .Z(c[331]) );
  XNOR U1161 ( .A(a[331]), .B(n979), .Z(n978) );
  IV U1162 ( .A(n976), .Z(n979) );
  XOR U1163 ( .A(n980), .B(n981), .Z(n976) );
  ANDN U1164 ( .B(n982), .A(n983), .Z(n980) );
  XNOR U1165 ( .A(b[330]), .B(n981), .Z(n982) );
  XNOR U1166 ( .A(b[330]), .B(n983), .Z(c[330]) );
  XNOR U1167 ( .A(a[330]), .B(n984), .Z(n983) );
  IV U1168 ( .A(n981), .Z(n984) );
  XOR U1169 ( .A(n985), .B(n986), .Z(n981) );
  ANDN U1170 ( .B(n987), .A(n988), .Z(n985) );
  XNOR U1171 ( .A(b[329]), .B(n986), .Z(n987) );
  XNOR U1172 ( .A(b[32]), .B(n989), .Z(c[32]) );
  XNOR U1173 ( .A(b[329]), .B(n988), .Z(c[329]) );
  XNOR U1174 ( .A(a[329]), .B(n990), .Z(n988) );
  IV U1175 ( .A(n986), .Z(n990) );
  XOR U1176 ( .A(n991), .B(n992), .Z(n986) );
  ANDN U1177 ( .B(n993), .A(n994), .Z(n991) );
  XNOR U1178 ( .A(b[328]), .B(n992), .Z(n993) );
  XNOR U1179 ( .A(b[328]), .B(n994), .Z(c[328]) );
  XNOR U1180 ( .A(a[328]), .B(n995), .Z(n994) );
  IV U1181 ( .A(n992), .Z(n995) );
  XOR U1182 ( .A(n996), .B(n997), .Z(n992) );
  ANDN U1183 ( .B(n998), .A(n999), .Z(n996) );
  XNOR U1184 ( .A(b[327]), .B(n997), .Z(n998) );
  XNOR U1185 ( .A(b[327]), .B(n999), .Z(c[327]) );
  XNOR U1186 ( .A(a[327]), .B(n1000), .Z(n999) );
  IV U1187 ( .A(n997), .Z(n1000) );
  XOR U1188 ( .A(n1001), .B(n1002), .Z(n997) );
  ANDN U1189 ( .B(n1003), .A(n1004), .Z(n1001) );
  XNOR U1190 ( .A(b[326]), .B(n1002), .Z(n1003) );
  XNOR U1191 ( .A(b[326]), .B(n1004), .Z(c[326]) );
  XNOR U1192 ( .A(a[326]), .B(n1005), .Z(n1004) );
  IV U1193 ( .A(n1002), .Z(n1005) );
  XOR U1194 ( .A(n1006), .B(n1007), .Z(n1002) );
  ANDN U1195 ( .B(n1008), .A(n1009), .Z(n1006) );
  XNOR U1196 ( .A(b[325]), .B(n1007), .Z(n1008) );
  XNOR U1197 ( .A(b[325]), .B(n1009), .Z(c[325]) );
  XNOR U1198 ( .A(a[325]), .B(n1010), .Z(n1009) );
  IV U1199 ( .A(n1007), .Z(n1010) );
  XOR U1200 ( .A(n1011), .B(n1012), .Z(n1007) );
  ANDN U1201 ( .B(n1013), .A(n1014), .Z(n1011) );
  XNOR U1202 ( .A(b[324]), .B(n1012), .Z(n1013) );
  XNOR U1203 ( .A(b[324]), .B(n1014), .Z(c[324]) );
  XNOR U1204 ( .A(a[324]), .B(n1015), .Z(n1014) );
  IV U1205 ( .A(n1012), .Z(n1015) );
  XOR U1206 ( .A(n1016), .B(n1017), .Z(n1012) );
  ANDN U1207 ( .B(n1018), .A(n1019), .Z(n1016) );
  XNOR U1208 ( .A(b[323]), .B(n1017), .Z(n1018) );
  XNOR U1209 ( .A(b[323]), .B(n1019), .Z(c[323]) );
  XNOR U1210 ( .A(a[323]), .B(n1020), .Z(n1019) );
  IV U1211 ( .A(n1017), .Z(n1020) );
  XOR U1212 ( .A(n1021), .B(n1022), .Z(n1017) );
  ANDN U1213 ( .B(n1023), .A(n1024), .Z(n1021) );
  XNOR U1214 ( .A(b[322]), .B(n1022), .Z(n1023) );
  XNOR U1215 ( .A(b[322]), .B(n1024), .Z(c[322]) );
  XNOR U1216 ( .A(a[322]), .B(n1025), .Z(n1024) );
  IV U1217 ( .A(n1022), .Z(n1025) );
  XOR U1218 ( .A(n1026), .B(n1027), .Z(n1022) );
  ANDN U1219 ( .B(n1028), .A(n1029), .Z(n1026) );
  XNOR U1220 ( .A(b[321]), .B(n1027), .Z(n1028) );
  XNOR U1221 ( .A(b[321]), .B(n1029), .Z(c[321]) );
  XNOR U1222 ( .A(a[321]), .B(n1030), .Z(n1029) );
  IV U1223 ( .A(n1027), .Z(n1030) );
  XOR U1224 ( .A(n1031), .B(n1032), .Z(n1027) );
  ANDN U1225 ( .B(n1033), .A(n1034), .Z(n1031) );
  XNOR U1226 ( .A(b[320]), .B(n1032), .Z(n1033) );
  XNOR U1227 ( .A(b[320]), .B(n1034), .Z(c[320]) );
  XNOR U1228 ( .A(a[320]), .B(n1035), .Z(n1034) );
  IV U1229 ( .A(n1032), .Z(n1035) );
  XOR U1230 ( .A(n1036), .B(n1037), .Z(n1032) );
  ANDN U1231 ( .B(n1038), .A(n1039), .Z(n1036) );
  XNOR U1232 ( .A(b[319]), .B(n1037), .Z(n1038) );
  XNOR U1233 ( .A(b[31]), .B(n1040), .Z(c[31]) );
  XNOR U1234 ( .A(b[319]), .B(n1039), .Z(c[319]) );
  XNOR U1235 ( .A(a[319]), .B(n1041), .Z(n1039) );
  IV U1236 ( .A(n1037), .Z(n1041) );
  XOR U1237 ( .A(n1042), .B(n1043), .Z(n1037) );
  ANDN U1238 ( .B(n1044), .A(n1045), .Z(n1042) );
  XNOR U1239 ( .A(b[318]), .B(n1043), .Z(n1044) );
  XNOR U1240 ( .A(b[318]), .B(n1045), .Z(c[318]) );
  XNOR U1241 ( .A(a[318]), .B(n1046), .Z(n1045) );
  IV U1242 ( .A(n1043), .Z(n1046) );
  XOR U1243 ( .A(n1047), .B(n1048), .Z(n1043) );
  ANDN U1244 ( .B(n1049), .A(n1050), .Z(n1047) );
  XNOR U1245 ( .A(b[317]), .B(n1048), .Z(n1049) );
  XNOR U1246 ( .A(b[317]), .B(n1050), .Z(c[317]) );
  XNOR U1247 ( .A(a[317]), .B(n1051), .Z(n1050) );
  IV U1248 ( .A(n1048), .Z(n1051) );
  XOR U1249 ( .A(n1052), .B(n1053), .Z(n1048) );
  ANDN U1250 ( .B(n1054), .A(n1055), .Z(n1052) );
  XNOR U1251 ( .A(b[316]), .B(n1053), .Z(n1054) );
  XNOR U1252 ( .A(b[316]), .B(n1055), .Z(c[316]) );
  XNOR U1253 ( .A(a[316]), .B(n1056), .Z(n1055) );
  IV U1254 ( .A(n1053), .Z(n1056) );
  XOR U1255 ( .A(n1057), .B(n1058), .Z(n1053) );
  ANDN U1256 ( .B(n1059), .A(n1060), .Z(n1057) );
  XNOR U1257 ( .A(b[315]), .B(n1058), .Z(n1059) );
  XNOR U1258 ( .A(b[315]), .B(n1060), .Z(c[315]) );
  XNOR U1259 ( .A(a[315]), .B(n1061), .Z(n1060) );
  IV U1260 ( .A(n1058), .Z(n1061) );
  XOR U1261 ( .A(n1062), .B(n1063), .Z(n1058) );
  ANDN U1262 ( .B(n1064), .A(n1065), .Z(n1062) );
  XNOR U1263 ( .A(b[314]), .B(n1063), .Z(n1064) );
  XNOR U1264 ( .A(b[314]), .B(n1065), .Z(c[314]) );
  XNOR U1265 ( .A(a[314]), .B(n1066), .Z(n1065) );
  IV U1266 ( .A(n1063), .Z(n1066) );
  XOR U1267 ( .A(n1067), .B(n1068), .Z(n1063) );
  ANDN U1268 ( .B(n1069), .A(n1070), .Z(n1067) );
  XNOR U1269 ( .A(b[313]), .B(n1068), .Z(n1069) );
  XNOR U1270 ( .A(b[313]), .B(n1070), .Z(c[313]) );
  XNOR U1271 ( .A(a[313]), .B(n1071), .Z(n1070) );
  IV U1272 ( .A(n1068), .Z(n1071) );
  XOR U1273 ( .A(n1072), .B(n1073), .Z(n1068) );
  ANDN U1274 ( .B(n1074), .A(n1075), .Z(n1072) );
  XNOR U1275 ( .A(b[312]), .B(n1073), .Z(n1074) );
  XNOR U1276 ( .A(b[312]), .B(n1075), .Z(c[312]) );
  XNOR U1277 ( .A(a[312]), .B(n1076), .Z(n1075) );
  IV U1278 ( .A(n1073), .Z(n1076) );
  XOR U1279 ( .A(n1077), .B(n1078), .Z(n1073) );
  ANDN U1280 ( .B(n1079), .A(n1080), .Z(n1077) );
  XNOR U1281 ( .A(b[311]), .B(n1078), .Z(n1079) );
  XNOR U1282 ( .A(b[311]), .B(n1080), .Z(c[311]) );
  XNOR U1283 ( .A(a[311]), .B(n1081), .Z(n1080) );
  IV U1284 ( .A(n1078), .Z(n1081) );
  XOR U1285 ( .A(n1082), .B(n1083), .Z(n1078) );
  ANDN U1286 ( .B(n1084), .A(n1085), .Z(n1082) );
  XNOR U1287 ( .A(b[310]), .B(n1083), .Z(n1084) );
  XNOR U1288 ( .A(b[310]), .B(n1085), .Z(c[310]) );
  XNOR U1289 ( .A(a[310]), .B(n1086), .Z(n1085) );
  IV U1290 ( .A(n1083), .Z(n1086) );
  XOR U1291 ( .A(n1087), .B(n1088), .Z(n1083) );
  ANDN U1292 ( .B(n1089), .A(n1090), .Z(n1087) );
  XNOR U1293 ( .A(b[309]), .B(n1088), .Z(n1089) );
  XNOR U1294 ( .A(b[30]), .B(n1091), .Z(c[30]) );
  XNOR U1295 ( .A(b[309]), .B(n1090), .Z(c[309]) );
  XNOR U1296 ( .A(a[309]), .B(n1092), .Z(n1090) );
  IV U1297 ( .A(n1088), .Z(n1092) );
  XOR U1298 ( .A(n1093), .B(n1094), .Z(n1088) );
  ANDN U1299 ( .B(n1095), .A(n1096), .Z(n1093) );
  XNOR U1300 ( .A(b[308]), .B(n1094), .Z(n1095) );
  XNOR U1301 ( .A(b[308]), .B(n1096), .Z(c[308]) );
  XNOR U1302 ( .A(a[308]), .B(n1097), .Z(n1096) );
  IV U1303 ( .A(n1094), .Z(n1097) );
  XOR U1304 ( .A(n1098), .B(n1099), .Z(n1094) );
  ANDN U1305 ( .B(n1100), .A(n1101), .Z(n1098) );
  XNOR U1306 ( .A(b[307]), .B(n1099), .Z(n1100) );
  XNOR U1307 ( .A(b[307]), .B(n1101), .Z(c[307]) );
  XNOR U1308 ( .A(a[307]), .B(n1102), .Z(n1101) );
  IV U1309 ( .A(n1099), .Z(n1102) );
  XOR U1310 ( .A(n1103), .B(n1104), .Z(n1099) );
  ANDN U1311 ( .B(n1105), .A(n1106), .Z(n1103) );
  XNOR U1312 ( .A(b[306]), .B(n1104), .Z(n1105) );
  XNOR U1313 ( .A(b[306]), .B(n1106), .Z(c[306]) );
  XNOR U1314 ( .A(a[306]), .B(n1107), .Z(n1106) );
  IV U1315 ( .A(n1104), .Z(n1107) );
  XOR U1316 ( .A(n1108), .B(n1109), .Z(n1104) );
  ANDN U1317 ( .B(n1110), .A(n1111), .Z(n1108) );
  XNOR U1318 ( .A(b[305]), .B(n1109), .Z(n1110) );
  XNOR U1319 ( .A(b[305]), .B(n1111), .Z(c[305]) );
  XNOR U1320 ( .A(a[305]), .B(n1112), .Z(n1111) );
  IV U1321 ( .A(n1109), .Z(n1112) );
  XOR U1322 ( .A(n1113), .B(n1114), .Z(n1109) );
  ANDN U1323 ( .B(n1115), .A(n1116), .Z(n1113) );
  XNOR U1324 ( .A(b[304]), .B(n1114), .Z(n1115) );
  XNOR U1325 ( .A(b[304]), .B(n1116), .Z(c[304]) );
  XNOR U1326 ( .A(a[304]), .B(n1117), .Z(n1116) );
  IV U1327 ( .A(n1114), .Z(n1117) );
  XOR U1328 ( .A(n1118), .B(n1119), .Z(n1114) );
  ANDN U1329 ( .B(n1120), .A(n1121), .Z(n1118) );
  XNOR U1330 ( .A(b[303]), .B(n1119), .Z(n1120) );
  XNOR U1331 ( .A(b[303]), .B(n1121), .Z(c[303]) );
  XNOR U1332 ( .A(a[303]), .B(n1122), .Z(n1121) );
  IV U1333 ( .A(n1119), .Z(n1122) );
  XOR U1334 ( .A(n1123), .B(n1124), .Z(n1119) );
  ANDN U1335 ( .B(n1125), .A(n1126), .Z(n1123) );
  XNOR U1336 ( .A(b[302]), .B(n1124), .Z(n1125) );
  XNOR U1337 ( .A(b[302]), .B(n1126), .Z(c[302]) );
  XNOR U1338 ( .A(a[302]), .B(n1127), .Z(n1126) );
  IV U1339 ( .A(n1124), .Z(n1127) );
  XOR U1340 ( .A(n1128), .B(n1129), .Z(n1124) );
  ANDN U1341 ( .B(n1130), .A(n1131), .Z(n1128) );
  XNOR U1342 ( .A(b[301]), .B(n1129), .Z(n1130) );
  XNOR U1343 ( .A(b[301]), .B(n1131), .Z(c[301]) );
  XNOR U1344 ( .A(a[301]), .B(n1132), .Z(n1131) );
  IV U1345 ( .A(n1129), .Z(n1132) );
  XOR U1346 ( .A(n1133), .B(n1134), .Z(n1129) );
  ANDN U1347 ( .B(n1135), .A(n1136), .Z(n1133) );
  XNOR U1348 ( .A(b[300]), .B(n1134), .Z(n1135) );
  XNOR U1349 ( .A(b[300]), .B(n1136), .Z(c[300]) );
  XNOR U1350 ( .A(a[300]), .B(n1137), .Z(n1136) );
  IV U1351 ( .A(n1134), .Z(n1137) );
  XOR U1352 ( .A(n1138), .B(n1139), .Z(n1134) );
  ANDN U1353 ( .B(n1140), .A(n1141), .Z(n1138) );
  XNOR U1354 ( .A(b[299]), .B(n1139), .Z(n1140) );
  XNOR U1355 ( .A(b[2]), .B(n1142), .Z(c[2]) );
  XNOR U1356 ( .A(b[29]), .B(n1143), .Z(c[29]) );
  XNOR U1357 ( .A(b[299]), .B(n1141), .Z(c[299]) );
  XNOR U1358 ( .A(a[299]), .B(n1144), .Z(n1141) );
  IV U1359 ( .A(n1139), .Z(n1144) );
  XOR U1360 ( .A(n1145), .B(n1146), .Z(n1139) );
  ANDN U1361 ( .B(n1147), .A(n1148), .Z(n1145) );
  XNOR U1362 ( .A(b[298]), .B(n1146), .Z(n1147) );
  XNOR U1363 ( .A(b[298]), .B(n1148), .Z(c[298]) );
  XNOR U1364 ( .A(a[298]), .B(n1149), .Z(n1148) );
  IV U1365 ( .A(n1146), .Z(n1149) );
  XOR U1366 ( .A(n1150), .B(n1151), .Z(n1146) );
  ANDN U1367 ( .B(n1152), .A(n1153), .Z(n1150) );
  XNOR U1368 ( .A(b[297]), .B(n1151), .Z(n1152) );
  XNOR U1369 ( .A(b[297]), .B(n1153), .Z(c[297]) );
  XNOR U1370 ( .A(a[297]), .B(n1154), .Z(n1153) );
  IV U1371 ( .A(n1151), .Z(n1154) );
  XOR U1372 ( .A(n1155), .B(n1156), .Z(n1151) );
  ANDN U1373 ( .B(n1157), .A(n1158), .Z(n1155) );
  XNOR U1374 ( .A(b[296]), .B(n1156), .Z(n1157) );
  XNOR U1375 ( .A(b[296]), .B(n1158), .Z(c[296]) );
  XNOR U1376 ( .A(a[296]), .B(n1159), .Z(n1158) );
  IV U1377 ( .A(n1156), .Z(n1159) );
  XOR U1378 ( .A(n1160), .B(n1161), .Z(n1156) );
  ANDN U1379 ( .B(n1162), .A(n1163), .Z(n1160) );
  XNOR U1380 ( .A(b[295]), .B(n1161), .Z(n1162) );
  XNOR U1381 ( .A(b[295]), .B(n1163), .Z(c[295]) );
  XNOR U1382 ( .A(a[295]), .B(n1164), .Z(n1163) );
  IV U1383 ( .A(n1161), .Z(n1164) );
  XOR U1384 ( .A(n1165), .B(n1166), .Z(n1161) );
  ANDN U1385 ( .B(n1167), .A(n1168), .Z(n1165) );
  XNOR U1386 ( .A(b[294]), .B(n1166), .Z(n1167) );
  XNOR U1387 ( .A(b[294]), .B(n1168), .Z(c[294]) );
  XNOR U1388 ( .A(a[294]), .B(n1169), .Z(n1168) );
  IV U1389 ( .A(n1166), .Z(n1169) );
  XOR U1390 ( .A(n1170), .B(n1171), .Z(n1166) );
  ANDN U1391 ( .B(n1172), .A(n1173), .Z(n1170) );
  XNOR U1392 ( .A(b[293]), .B(n1171), .Z(n1172) );
  XNOR U1393 ( .A(b[293]), .B(n1173), .Z(c[293]) );
  XNOR U1394 ( .A(a[293]), .B(n1174), .Z(n1173) );
  IV U1395 ( .A(n1171), .Z(n1174) );
  XOR U1396 ( .A(n1175), .B(n1176), .Z(n1171) );
  ANDN U1397 ( .B(n1177), .A(n1178), .Z(n1175) );
  XNOR U1398 ( .A(b[292]), .B(n1176), .Z(n1177) );
  XNOR U1399 ( .A(b[292]), .B(n1178), .Z(c[292]) );
  XNOR U1400 ( .A(a[292]), .B(n1179), .Z(n1178) );
  IV U1401 ( .A(n1176), .Z(n1179) );
  XOR U1402 ( .A(n1180), .B(n1181), .Z(n1176) );
  ANDN U1403 ( .B(n1182), .A(n1183), .Z(n1180) );
  XNOR U1404 ( .A(b[291]), .B(n1181), .Z(n1182) );
  XNOR U1405 ( .A(b[291]), .B(n1183), .Z(c[291]) );
  XNOR U1406 ( .A(a[291]), .B(n1184), .Z(n1183) );
  IV U1407 ( .A(n1181), .Z(n1184) );
  XOR U1408 ( .A(n1185), .B(n1186), .Z(n1181) );
  ANDN U1409 ( .B(n1187), .A(n1188), .Z(n1185) );
  XNOR U1410 ( .A(b[290]), .B(n1186), .Z(n1187) );
  XNOR U1411 ( .A(b[290]), .B(n1188), .Z(c[290]) );
  XNOR U1412 ( .A(a[290]), .B(n1189), .Z(n1188) );
  IV U1413 ( .A(n1186), .Z(n1189) );
  XOR U1414 ( .A(n1190), .B(n1191), .Z(n1186) );
  ANDN U1415 ( .B(n1192), .A(n1193), .Z(n1190) );
  XNOR U1416 ( .A(b[289]), .B(n1191), .Z(n1192) );
  XNOR U1417 ( .A(b[28]), .B(n1194), .Z(c[28]) );
  XNOR U1418 ( .A(b[289]), .B(n1193), .Z(c[289]) );
  XNOR U1419 ( .A(a[289]), .B(n1195), .Z(n1193) );
  IV U1420 ( .A(n1191), .Z(n1195) );
  XOR U1421 ( .A(n1196), .B(n1197), .Z(n1191) );
  ANDN U1422 ( .B(n1198), .A(n1199), .Z(n1196) );
  XNOR U1423 ( .A(b[288]), .B(n1197), .Z(n1198) );
  XNOR U1424 ( .A(b[288]), .B(n1199), .Z(c[288]) );
  XNOR U1425 ( .A(a[288]), .B(n1200), .Z(n1199) );
  IV U1426 ( .A(n1197), .Z(n1200) );
  XOR U1427 ( .A(n1201), .B(n1202), .Z(n1197) );
  ANDN U1428 ( .B(n1203), .A(n1204), .Z(n1201) );
  XNOR U1429 ( .A(b[287]), .B(n1202), .Z(n1203) );
  XNOR U1430 ( .A(b[287]), .B(n1204), .Z(c[287]) );
  XNOR U1431 ( .A(a[287]), .B(n1205), .Z(n1204) );
  IV U1432 ( .A(n1202), .Z(n1205) );
  XOR U1433 ( .A(n1206), .B(n1207), .Z(n1202) );
  ANDN U1434 ( .B(n1208), .A(n1209), .Z(n1206) );
  XNOR U1435 ( .A(b[286]), .B(n1207), .Z(n1208) );
  XNOR U1436 ( .A(b[286]), .B(n1209), .Z(c[286]) );
  XNOR U1437 ( .A(a[286]), .B(n1210), .Z(n1209) );
  IV U1438 ( .A(n1207), .Z(n1210) );
  XOR U1439 ( .A(n1211), .B(n1212), .Z(n1207) );
  ANDN U1440 ( .B(n1213), .A(n1214), .Z(n1211) );
  XNOR U1441 ( .A(b[285]), .B(n1212), .Z(n1213) );
  XNOR U1442 ( .A(b[285]), .B(n1214), .Z(c[285]) );
  XNOR U1443 ( .A(a[285]), .B(n1215), .Z(n1214) );
  IV U1444 ( .A(n1212), .Z(n1215) );
  XOR U1445 ( .A(n1216), .B(n1217), .Z(n1212) );
  ANDN U1446 ( .B(n1218), .A(n1219), .Z(n1216) );
  XNOR U1447 ( .A(b[284]), .B(n1217), .Z(n1218) );
  XNOR U1448 ( .A(b[284]), .B(n1219), .Z(c[284]) );
  XNOR U1449 ( .A(a[284]), .B(n1220), .Z(n1219) );
  IV U1450 ( .A(n1217), .Z(n1220) );
  XOR U1451 ( .A(n1221), .B(n1222), .Z(n1217) );
  ANDN U1452 ( .B(n1223), .A(n1224), .Z(n1221) );
  XNOR U1453 ( .A(b[283]), .B(n1222), .Z(n1223) );
  XNOR U1454 ( .A(b[283]), .B(n1224), .Z(c[283]) );
  XNOR U1455 ( .A(a[283]), .B(n1225), .Z(n1224) );
  IV U1456 ( .A(n1222), .Z(n1225) );
  XOR U1457 ( .A(n1226), .B(n1227), .Z(n1222) );
  ANDN U1458 ( .B(n1228), .A(n1229), .Z(n1226) );
  XNOR U1459 ( .A(b[282]), .B(n1227), .Z(n1228) );
  XNOR U1460 ( .A(b[282]), .B(n1229), .Z(c[282]) );
  XNOR U1461 ( .A(a[282]), .B(n1230), .Z(n1229) );
  IV U1462 ( .A(n1227), .Z(n1230) );
  XOR U1463 ( .A(n1231), .B(n1232), .Z(n1227) );
  ANDN U1464 ( .B(n1233), .A(n1234), .Z(n1231) );
  XNOR U1465 ( .A(b[281]), .B(n1232), .Z(n1233) );
  XNOR U1466 ( .A(b[281]), .B(n1234), .Z(c[281]) );
  XNOR U1467 ( .A(a[281]), .B(n1235), .Z(n1234) );
  IV U1468 ( .A(n1232), .Z(n1235) );
  XOR U1469 ( .A(n1236), .B(n1237), .Z(n1232) );
  ANDN U1470 ( .B(n1238), .A(n1239), .Z(n1236) );
  XNOR U1471 ( .A(b[280]), .B(n1237), .Z(n1238) );
  XNOR U1472 ( .A(b[280]), .B(n1239), .Z(c[280]) );
  XNOR U1473 ( .A(a[280]), .B(n1240), .Z(n1239) );
  IV U1474 ( .A(n1237), .Z(n1240) );
  XOR U1475 ( .A(n1241), .B(n1242), .Z(n1237) );
  ANDN U1476 ( .B(n1243), .A(n1244), .Z(n1241) );
  XNOR U1477 ( .A(b[279]), .B(n1242), .Z(n1243) );
  XNOR U1478 ( .A(b[27]), .B(n1245), .Z(c[27]) );
  XNOR U1479 ( .A(b[279]), .B(n1244), .Z(c[279]) );
  XNOR U1480 ( .A(a[279]), .B(n1246), .Z(n1244) );
  IV U1481 ( .A(n1242), .Z(n1246) );
  XOR U1482 ( .A(n1247), .B(n1248), .Z(n1242) );
  ANDN U1483 ( .B(n1249), .A(n1250), .Z(n1247) );
  XNOR U1484 ( .A(b[278]), .B(n1248), .Z(n1249) );
  XNOR U1485 ( .A(b[278]), .B(n1250), .Z(c[278]) );
  XNOR U1486 ( .A(a[278]), .B(n1251), .Z(n1250) );
  IV U1487 ( .A(n1248), .Z(n1251) );
  XOR U1488 ( .A(n1252), .B(n1253), .Z(n1248) );
  ANDN U1489 ( .B(n1254), .A(n1255), .Z(n1252) );
  XNOR U1490 ( .A(b[277]), .B(n1253), .Z(n1254) );
  XNOR U1491 ( .A(b[277]), .B(n1255), .Z(c[277]) );
  XNOR U1492 ( .A(a[277]), .B(n1256), .Z(n1255) );
  IV U1493 ( .A(n1253), .Z(n1256) );
  XOR U1494 ( .A(n1257), .B(n1258), .Z(n1253) );
  ANDN U1495 ( .B(n1259), .A(n1260), .Z(n1257) );
  XNOR U1496 ( .A(b[276]), .B(n1258), .Z(n1259) );
  XNOR U1497 ( .A(b[276]), .B(n1260), .Z(c[276]) );
  XNOR U1498 ( .A(a[276]), .B(n1261), .Z(n1260) );
  IV U1499 ( .A(n1258), .Z(n1261) );
  XOR U1500 ( .A(n1262), .B(n1263), .Z(n1258) );
  ANDN U1501 ( .B(n1264), .A(n1265), .Z(n1262) );
  XNOR U1502 ( .A(b[275]), .B(n1263), .Z(n1264) );
  XNOR U1503 ( .A(b[275]), .B(n1265), .Z(c[275]) );
  XNOR U1504 ( .A(a[275]), .B(n1266), .Z(n1265) );
  IV U1505 ( .A(n1263), .Z(n1266) );
  XOR U1506 ( .A(n1267), .B(n1268), .Z(n1263) );
  ANDN U1507 ( .B(n1269), .A(n1270), .Z(n1267) );
  XNOR U1508 ( .A(b[274]), .B(n1268), .Z(n1269) );
  XNOR U1509 ( .A(b[274]), .B(n1270), .Z(c[274]) );
  XNOR U1510 ( .A(a[274]), .B(n1271), .Z(n1270) );
  IV U1511 ( .A(n1268), .Z(n1271) );
  XOR U1512 ( .A(n1272), .B(n1273), .Z(n1268) );
  ANDN U1513 ( .B(n1274), .A(n1275), .Z(n1272) );
  XNOR U1514 ( .A(b[273]), .B(n1273), .Z(n1274) );
  XNOR U1515 ( .A(b[273]), .B(n1275), .Z(c[273]) );
  XNOR U1516 ( .A(a[273]), .B(n1276), .Z(n1275) );
  IV U1517 ( .A(n1273), .Z(n1276) );
  XOR U1518 ( .A(n1277), .B(n1278), .Z(n1273) );
  ANDN U1519 ( .B(n1279), .A(n1280), .Z(n1277) );
  XNOR U1520 ( .A(b[272]), .B(n1278), .Z(n1279) );
  XNOR U1521 ( .A(b[272]), .B(n1280), .Z(c[272]) );
  XNOR U1522 ( .A(a[272]), .B(n1281), .Z(n1280) );
  IV U1523 ( .A(n1278), .Z(n1281) );
  XOR U1524 ( .A(n1282), .B(n1283), .Z(n1278) );
  ANDN U1525 ( .B(n1284), .A(n1285), .Z(n1282) );
  XNOR U1526 ( .A(b[271]), .B(n1283), .Z(n1284) );
  XNOR U1527 ( .A(b[271]), .B(n1285), .Z(c[271]) );
  XNOR U1528 ( .A(a[271]), .B(n1286), .Z(n1285) );
  IV U1529 ( .A(n1283), .Z(n1286) );
  XOR U1530 ( .A(n1287), .B(n1288), .Z(n1283) );
  ANDN U1531 ( .B(n1289), .A(n1290), .Z(n1287) );
  XNOR U1532 ( .A(b[270]), .B(n1288), .Z(n1289) );
  XNOR U1533 ( .A(b[270]), .B(n1290), .Z(c[270]) );
  XNOR U1534 ( .A(a[270]), .B(n1291), .Z(n1290) );
  IV U1535 ( .A(n1288), .Z(n1291) );
  XOR U1536 ( .A(n1292), .B(n1293), .Z(n1288) );
  ANDN U1537 ( .B(n1294), .A(n1295), .Z(n1292) );
  XNOR U1538 ( .A(b[269]), .B(n1293), .Z(n1294) );
  XNOR U1539 ( .A(b[26]), .B(n1296), .Z(c[26]) );
  XNOR U1540 ( .A(b[269]), .B(n1295), .Z(c[269]) );
  XNOR U1541 ( .A(a[269]), .B(n1297), .Z(n1295) );
  IV U1542 ( .A(n1293), .Z(n1297) );
  XOR U1543 ( .A(n1298), .B(n1299), .Z(n1293) );
  ANDN U1544 ( .B(n1300), .A(n1301), .Z(n1298) );
  XNOR U1545 ( .A(b[268]), .B(n1299), .Z(n1300) );
  XNOR U1546 ( .A(b[268]), .B(n1301), .Z(c[268]) );
  XNOR U1547 ( .A(a[268]), .B(n1302), .Z(n1301) );
  IV U1548 ( .A(n1299), .Z(n1302) );
  XOR U1549 ( .A(n1303), .B(n1304), .Z(n1299) );
  ANDN U1550 ( .B(n1305), .A(n1306), .Z(n1303) );
  XNOR U1551 ( .A(b[267]), .B(n1304), .Z(n1305) );
  XNOR U1552 ( .A(b[267]), .B(n1306), .Z(c[267]) );
  XNOR U1553 ( .A(a[267]), .B(n1307), .Z(n1306) );
  IV U1554 ( .A(n1304), .Z(n1307) );
  XOR U1555 ( .A(n1308), .B(n1309), .Z(n1304) );
  ANDN U1556 ( .B(n1310), .A(n1311), .Z(n1308) );
  XNOR U1557 ( .A(b[266]), .B(n1309), .Z(n1310) );
  XNOR U1558 ( .A(b[266]), .B(n1311), .Z(c[266]) );
  XNOR U1559 ( .A(a[266]), .B(n1312), .Z(n1311) );
  IV U1560 ( .A(n1309), .Z(n1312) );
  XOR U1561 ( .A(n1313), .B(n1314), .Z(n1309) );
  ANDN U1562 ( .B(n1315), .A(n1316), .Z(n1313) );
  XNOR U1563 ( .A(b[265]), .B(n1314), .Z(n1315) );
  XNOR U1564 ( .A(b[265]), .B(n1316), .Z(c[265]) );
  XNOR U1565 ( .A(a[265]), .B(n1317), .Z(n1316) );
  IV U1566 ( .A(n1314), .Z(n1317) );
  XOR U1567 ( .A(n1318), .B(n1319), .Z(n1314) );
  ANDN U1568 ( .B(n1320), .A(n1321), .Z(n1318) );
  XNOR U1569 ( .A(b[264]), .B(n1319), .Z(n1320) );
  XNOR U1570 ( .A(b[264]), .B(n1321), .Z(c[264]) );
  XNOR U1571 ( .A(a[264]), .B(n1322), .Z(n1321) );
  IV U1572 ( .A(n1319), .Z(n1322) );
  XOR U1573 ( .A(n1323), .B(n1324), .Z(n1319) );
  ANDN U1574 ( .B(n1325), .A(n1326), .Z(n1323) );
  XNOR U1575 ( .A(b[263]), .B(n1324), .Z(n1325) );
  XNOR U1576 ( .A(b[263]), .B(n1326), .Z(c[263]) );
  XNOR U1577 ( .A(a[263]), .B(n1327), .Z(n1326) );
  IV U1578 ( .A(n1324), .Z(n1327) );
  XOR U1579 ( .A(n1328), .B(n1329), .Z(n1324) );
  ANDN U1580 ( .B(n1330), .A(n1331), .Z(n1328) );
  XNOR U1581 ( .A(b[262]), .B(n1329), .Z(n1330) );
  XNOR U1582 ( .A(b[262]), .B(n1331), .Z(c[262]) );
  XNOR U1583 ( .A(a[262]), .B(n1332), .Z(n1331) );
  IV U1584 ( .A(n1329), .Z(n1332) );
  XOR U1585 ( .A(n1333), .B(n1334), .Z(n1329) );
  ANDN U1586 ( .B(n1335), .A(n1336), .Z(n1333) );
  XNOR U1587 ( .A(b[261]), .B(n1334), .Z(n1335) );
  XNOR U1588 ( .A(b[261]), .B(n1336), .Z(c[261]) );
  XNOR U1589 ( .A(a[261]), .B(n1337), .Z(n1336) );
  IV U1590 ( .A(n1334), .Z(n1337) );
  XOR U1591 ( .A(n1338), .B(n1339), .Z(n1334) );
  ANDN U1592 ( .B(n1340), .A(n1341), .Z(n1338) );
  XNOR U1593 ( .A(b[260]), .B(n1339), .Z(n1340) );
  XNOR U1594 ( .A(b[260]), .B(n1341), .Z(c[260]) );
  XNOR U1595 ( .A(a[260]), .B(n1342), .Z(n1341) );
  IV U1596 ( .A(n1339), .Z(n1342) );
  XOR U1597 ( .A(n1343), .B(n1344), .Z(n1339) );
  ANDN U1598 ( .B(n1345), .A(n1346), .Z(n1343) );
  XNOR U1599 ( .A(b[259]), .B(n1344), .Z(n1345) );
  XNOR U1600 ( .A(b[25]), .B(n1347), .Z(c[25]) );
  XNOR U1601 ( .A(b[259]), .B(n1346), .Z(c[259]) );
  XNOR U1602 ( .A(a[259]), .B(n1348), .Z(n1346) );
  IV U1603 ( .A(n1344), .Z(n1348) );
  XOR U1604 ( .A(n1349), .B(n1350), .Z(n1344) );
  ANDN U1605 ( .B(n1351), .A(n1352), .Z(n1349) );
  XNOR U1606 ( .A(b[258]), .B(n1350), .Z(n1351) );
  XNOR U1607 ( .A(b[258]), .B(n1352), .Z(c[258]) );
  XNOR U1608 ( .A(a[258]), .B(n1353), .Z(n1352) );
  IV U1609 ( .A(n1350), .Z(n1353) );
  XOR U1610 ( .A(n1354), .B(n1355), .Z(n1350) );
  ANDN U1611 ( .B(n1356), .A(n1357), .Z(n1354) );
  XNOR U1612 ( .A(b[257]), .B(n1355), .Z(n1356) );
  XNOR U1613 ( .A(b[257]), .B(n1357), .Z(c[257]) );
  XNOR U1614 ( .A(a[257]), .B(n1358), .Z(n1357) );
  IV U1615 ( .A(n1355), .Z(n1358) );
  XOR U1616 ( .A(n1359), .B(n1360), .Z(n1355) );
  ANDN U1617 ( .B(n1361), .A(n1362), .Z(n1359) );
  XNOR U1618 ( .A(b[256]), .B(n1360), .Z(n1361) );
  XNOR U1619 ( .A(b[256]), .B(n1362), .Z(c[256]) );
  XNOR U1620 ( .A(a[256]), .B(n1363), .Z(n1362) );
  IV U1621 ( .A(n1360), .Z(n1363) );
  XOR U1622 ( .A(n1364), .B(n1365), .Z(n1360) );
  ANDN U1623 ( .B(n1366), .A(n1367), .Z(n1364) );
  XNOR U1624 ( .A(b[255]), .B(n1365), .Z(n1366) );
  XNOR U1625 ( .A(b[255]), .B(n1367), .Z(c[255]) );
  XNOR U1626 ( .A(a[255]), .B(n1368), .Z(n1367) );
  IV U1627 ( .A(n1365), .Z(n1368) );
  XOR U1628 ( .A(n1369), .B(n1370), .Z(n1365) );
  ANDN U1629 ( .B(n1371), .A(n1372), .Z(n1369) );
  XNOR U1630 ( .A(b[254]), .B(n1370), .Z(n1371) );
  XNOR U1631 ( .A(b[254]), .B(n1372), .Z(c[254]) );
  XNOR U1632 ( .A(a[254]), .B(n1373), .Z(n1372) );
  IV U1633 ( .A(n1370), .Z(n1373) );
  XOR U1634 ( .A(n1374), .B(n1375), .Z(n1370) );
  ANDN U1635 ( .B(n1376), .A(n1377), .Z(n1374) );
  XNOR U1636 ( .A(b[253]), .B(n1375), .Z(n1376) );
  XNOR U1637 ( .A(b[253]), .B(n1377), .Z(c[253]) );
  XNOR U1638 ( .A(a[253]), .B(n1378), .Z(n1377) );
  IV U1639 ( .A(n1375), .Z(n1378) );
  XOR U1640 ( .A(n1379), .B(n1380), .Z(n1375) );
  ANDN U1641 ( .B(n1381), .A(n1382), .Z(n1379) );
  XNOR U1642 ( .A(b[252]), .B(n1380), .Z(n1381) );
  XNOR U1643 ( .A(b[252]), .B(n1382), .Z(c[252]) );
  XNOR U1644 ( .A(a[252]), .B(n1383), .Z(n1382) );
  IV U1645 ( .A(n1380), .Z(n1383) );
  XOR U1646 ( .A(n1384), .B(n1385), .Z(n1380) );
  ANDN U1647 ( .B(n1386), .A(n1387), .Z(n1384) );
  XNOR U1648 ( .A(b[251]), .B(n1385), .Z(n1386) );
  XNOR U1649 ( .A(b[251]), .B(n1387), .Z(c[251]) );
  XNOR U1650 ( .A(a[251]), .B(n1388), .Z(n1387) );
  IV U1651 ( .A(n1385), .Z(n1388) );
  XOR U1652 ( .A(n1389), .B(n1390), .Z(n1385) );
  ANDN U1653 ( .B(n1391), .A(n1392), .Z(n1389) );
  XNOR U1654 ( .A(b[250]), .B(n1390), .Z(n1391) );
  XNOR U1655 ( .A(b[250]), .B(n1392), .Z(c[250]) );
  XNOR U1656 ( .A(a[250]), .B(n1393), .Z(n1392) );
  IV U1657 ( .A(n1390), .Z(n1393) );
  XOR U1658 ( .A(n1394), .B(n1395), .Z(n1390) );
  ANDN U1659 ( .B(n1396), .A(n1397), .Z(n1394) );
  XNOR U1660 ( .A(b[249]), .B(n1395), .Z(n1396) );
  XNOR U1661 ( .A(b[24]), .B(n1398), .Z(c[24]) );
  XNOR U1662 ( .A(b[249]), .B(n1397), .Z(c[249]) );
  XNOR U1663 ( .A(a[249]), .B(n1399), .Z(n1397) );
  IV U1664 ( .A(n1395), .Z(n1399) );
  XOR U1665 ( .A(n1400), .B(n1401), .Z(n1395) );
  ANDN U1666 ( .B(n1402), .A(n1403), .Z(n1400) );
  XNOR U1667 ( .A(b[248]), .B(n1401), .Z(n1402) );
  XNOR U1668 ( .A(b[248]), .B(n1403), .Z(c[248]) );
  XNOR U1669 ( .A(a[248]), .B(n1404), .Z(n1403) );
  IV U1670 ( .A(n1401), .Z(n1404) );
  XOR U1671 ( .A(n1405), .B(n1406), .Z(n1401) );
  ANDN U1672 ( .B(n1407), .A(n1408), .Z(n1405) );
  XNOR U1673 ( .A(b[247]), .B(n1406), .Z(n1407) );
  XNOR U1674 ( .A(b[247]), .B(n1408), .Z(c[247]) );
  XNOR U1675 ( .A(a[247]), .B(n1409), .Z(n1408) );
  IV U1676 ( .A(n1406), .Z(n1409) );
  XOR U1677 ( .A(n1410), .B(n1411), .Z(n1406) );
  ANDN U1678 ( .B(n1412), .A(n1413), .Z(n1410) );
  XNOR U1679 ( .A(b[246]), .B(n1411), .Z(n1412) );
  XNOR U1680 ( .A(b[246]), .B(n1413), .Z(c[246]) );
  XNOR U1681 ( .A(a[246]), .B(n1414), .Z(n1413) );
  IV U1682 ( .A(n1411), .Z(n1414) );
  XOR U1683 ( .A(n1415), .B(n1416), .Z(n1411) );
  ANDN U1684 ( .B(n1417), .A(n1418), .Z(n1415) );
  XNOR U1685 ( .A(b[245]), .B(n1416), .Z(n1417) );
  XNOR U1686 ( .A(b[245]), .B(n1418), .Z(c[245]) );
  XNOR U1687 ( .A(a[245]), .B(n1419), .Z(n1418) );
  IV U1688 ( .A(n1416), .Z(n1419) );
  XOR U1689 ( .A(n1420), .B(n1421), .Z(n1416) );
  ANDN U1690 ( .B(n1422), .A(n1423), .Z(n1420) );
  XNOR U1691 ( .A(b[244]), .B(n1421), .Z(n1422) );
  XNOR U1692 ( .A(b[244]), .B(n1423), .Z(c[244]) );
  XNOR U1693 ( .A(a[244]), .B(n1424), .Z(n1423) );
  IV U1694 ( .A(n1421), .Z(n1424) );
  XOR U1695 ( .A(n1425), .B(n1426), .Z(n1421) );
  ANDN U1696 ( .B(n1427), .A(n1428), .Z(n1425) );
  XNOR U1697 ( .A(b[243]), .B(n1426), .Z(n1427) );
  XNOR U1698 ( .A(b[243]), .B(n1428), .Z(c[243]) );
  XNOR U1699 ( .A(a[243]), .B(n1429), .Z(n1428) );
  IV U1700 ( .A(n1426), .Z(n1429) );
  XOR U1701 ( .A(n1430), .B(n1431), .Z(n1426) );
  ANDN U1702 ( .B(n1432), .A(n1433), .Z(n1430) );
  XNOR U1703 ( .A(b[242]), .B(n1431), .Z(n1432) );
  XNOR U1704 ( .A(b[242]), .B(n1433), .Z(c[242]) );
  XNOR U1705 ( .A(a[242]), .B(n1434), .Z(n1433) );
  IV U1706 ( .A(n1431), .Z(n1434) );
  XOR U1707 ( .A(n1435), .B(n1436), .Z(n1431) );
  ANDN U1708 ( .B(n1437), .A(n1438), .Z(n1435) );
  XNOR U1709 ( .A(b[241]), .B(n1436), .Z(n1437) );
  XNOR U1710 ( .A(b[241]), .B(n1438), .Z(c[241]) );
  XNOR U1711 ( .A(a[241]), .B(n1439), .Z(n1438) );
  IV U1712 ( .A(n1436), .Z(n1439) );
  XOR U1713 ( .A(n1440), .B(n1441), .Z(n1436) );
  ANDN U1714 ( .B(n1442), .A(n1443), .Z(n1440) );
  XNOR U1715 ( .A(b[240]), .B(n1441), .Z(n1442) );
  XNOR U1716 ( .A(b[240]), .B(n1443), .Z(c[240]) );
  XNOR U1717 ( .A(a[240]), .B(n1444), .Z(n1443) );
  IV U1718 ( .A(n1441), .Z(n1444) );
  XOR U1719 ( .A(n1445), .B(n1446), .Z(n1441) );
  ANDN U1720 ( .B(n1447), .A(n1448), .Z(n1445) );
  XNOR U1721 ( .A(b[239]), .B(n1446), .Z(n1447) );
  XNOR U1722 ( .A(b[23]), .B(n1449), .Z(c[23]) );
  XNOR U1723 ( .A(b[239]), .B(n1448), .Z(c[239]) );
  XNOR U1724 ( .A(a[239]), .B(n1450), .Z(n1448) );
  IV U1725 ( .A(n1446), .Z(n1450) );
  XOR U1726 ( .A(n1451), .B(n1452), .Z(n1446) );
  ANDN U1727 ( .B(n1453), .A(n1454), .Z(n1451) );
  XNOR U1728 ( .A(b[238]), .B(n1452), .Z(n1453) );
  XNOR U1729 ( .A(b[238]), .B(n1454), .Z(c[238]) );
  XNOR U1730 ( .A(a[238]), .B(n1455), .Z(n1454) );
  IV U1731 ( .A(n1452), .Z(n1455) );
  XOR U1732 ( .A(n1456), .B(n1457), .Z(n1452) );
  ANDN U1733 ( .B(n1458), .A(n1459), .Z(n1456) );
  XNOR U1734 ( .A(b[237]), .B(n1457), .Z(n1458) );
  XNOR U1735 ( .A(b[237]), .B(n1459), .Z(c[237]) );
  XNOR U1736 ( .A(a[237]), .B(n1460), .Z(n1459) );
  IV U1737 ( .A(n1457), .Z(n1460) );
  XOR U1738 ( .A(n1461), .B(n1462), .Z(n1457) );
  ANDN U1739 ( .B(n1463), .A(n1464), .Z(n1461) );
  XNOR U1740 ( .A(b[236]), .B(n1462), .Z(n1463) );
  XNOR U1741 ( .A(b[236]), .B(n1464), .Z(c[236]) );
  XNOR U1742 ( .A(a[236]), .B(n1465), .Z(n1464) );
  IV U1743 ( .A(n1462), .Z(n1465) );
  XOR U1744 ( .A(n1466), .B(n1467), .Z(n1462) );
  ANDN U1745 ( .B(n1468), .A(n1469), .Z(n1466) );
  XNOR U1746 ( .A(b[235]), .B(n1467), .Z(n1468) );
  XNOR U1747 ( .A(b[235]), .B(n1469), .Z(c[235]) );
  XNOR U1748 ( .A(a[235]), .B(n1470), .Z(n1469) );
  IV U1749 ( .A(n1467), .Z(n1470) );
  XOR U1750 ( .A(n1471), .B(n1472), .Z(n1467) );
  ANDN U1751 ( .B(n1473), .A(n1474), .Z(n1471) );
  XNOR U1752 ( .A(b[234]), .B(n1472), .Z(n1473) );
  XNOR U1753 ( .A(b[234]), .B(n1474), .Z(c[234]) );
  XNOR U1754 ( .A(a[234]), .B(n1475), .Z(n1474) );
  IV U1755 ( .A(n1472), .Z(n1475) );
  XOR U1756 ( .A(n1476), .B(n1477), .Z(n1472) );
  ANDN U1757 ( .B(n1478), .A(n1479), .Z(n1476) );
  XNOR U1758 ( .A(b[233]), .B(n1477), .Z(n1478) );
  XNOR U1759 ( .A(b[233]), .B(n1479), .Z(c[233]) );
  XNOR U1760 ( .A(a[233]), .B(n1480), .Z(n1479) );
  IV U1761 ( .A(n1477), .Z(n1480) );
  XOR U1762 ( .A(n1481), .B(n1482), .Z(n1477) );
  ANDN U1763 ( .B(n1483), .A(n1484), .Z(n1481) );
  XNOR U1764 ( .A(b[232]), .B(n1482), .Z(n1483) );
  XNOR U1765 ( .A(b[232]), .B(n1484), .Z(c[232]) );
  XNOR U1766 ( .A(a[232]), .B(n1485), .Z(n1484) );
  IV U1767 ( .A(n1482), .Z(n1485) );
  XOR U1768 ( .A(n1486), .B(n1487), .Z(n1482) );
  ANDN U1769 ( .B(n1488), .A(n1489), .Z(n1486) );
  XNOR U1770 ( .A(b[231]), .B(n1487), .Z(n1488) );
  XNOR U1771 ( .A(b[231]), .B(n1489), .Z(c[231]) );
  XNOR U1772 ( .A(a[231]), .B(n1490), .Z(n1489) );
  IV U1773 ( .A(n1487), .Z(n1490) );
  XOR U1774 ( .A(n1491), .B(n1492), .Z(n1487) );
  ANDN U1775 ( .B(n1493), .A(n1494), .Z(n1491) );
  XNOR U1776 ( .A(b[230]), .B(n1492), .Z(n1493) );
  XNOR U1777 ( .A(b[230]), .B(n1494), .Z(c[230]) );
  XNOR U1778 ( .A(a[230]), .B(n1495), .Z(n1494) );
  IV U1779 ( .A(n1492), .Z(n1495) );
  XOR U1780 ( .A(n1496), .B(n1497), .Z(n1492) );
  ANDN U1781 ( .B(n1498), .A(n1499), .Z(n1496) );
  XNOR U1782 ( .A(b[229]), .B(n1497), .Z(n1498) );
  XNOR U1783 ( .A(b[22]), .B(n1500), .Z(c[22]) );
  XNOR U1784 ( .A(b[229]), .B(n1499), .Z(c[229]) );
  XNOR U1785 ( .A(a[229]), .B(n1501), .Z(n1499) );
  IV U1786 ( .A(n1497), .Z(n1501) );
  XOR U1787 ( .A(n1502), .B(n1503), .Z(n1497) );
  ANDN U1788 ( .B(n1504), .A(n1505), .Z(n1502) );
  XNOR U1789 ( .A(b[228]), .B(n1503), .Z(n1504) );
  XNOR U1790 ( .A(b[228]), .B(n1505), .Z(c[228]) );
  XNOR U1791 ( .A(a[228]), .B(n1506), .Z(n1505) );
  IV U1792 ( .A(n1503), .Z(n1506) );
  XOR U1793 ( .A(n1507), .B(n1508), .Z(n1503) );
  ANDN U1794 ( .B(n1509), .A(n1510), .Z(n1507) );
  XNOR U1795 ( .A(b[227]), .B(n1508), .Z(n1509) );
  XNOR U1796 ( .A(b[227]), .B(n1510), .Z(c[227]) );
  XNOR U1797 ( .A(a[227]), .B(n1511), .Z(n1510) );
  IV U1798 ( .A(n1508), .Z(n1511) );
  XOR U1799 ( .A(n1512), .B(n1513), .Z(n1508) );
  ANDN U1800 ( .B(n1514), .A(n1515), .Z(n1512) );
  XNOR U1801 ( .A(b[226]), .B(n1513), .Z(n1514) );
  XNOR U1802 ( .A(b[226]), .B(n1515), .Z(c[226]) );
  XNOR U1803 ( .A(a[226]), .B(n1516), .Z(n1515) );
  IV U1804 ( .A(n1513), .Z(n1516) );
  XOR U1805 ( .A(n1517), .B(n1518), .Z(n1513) );
  ANDN U1806 ( .B(n1519), .A(n1520), .Z(n1517) );
  XNOR U1807 ( .A(b[225]), .B(n1518), .Z(n1519) );
  XNOR U1808 ( .A(b[225]), .B(n1520), .Z(c[225]) );
  XNOR U1809 ( .A(a[225]), .B(n1521), .Z(n1520) );
  IV U1810 ( .A(n1518), .Z(n1521) );
  XOR U1811 ( .A(n1522), .B(n1523), .Z(n1518) );
  ANDN U1812 ( .B(n1524), .A(n1525), .Z(n1522) );
  XNOR U1813 ( .A(b[224]), .B(n1523), .Z(n1524) );
  XNOR U1814 ( .A(b[224]), .B(n1525), .Z(c[224]) );
  XNOR U1815 ( .A(a[224]), .B(n1526), .Z(n1525) );
  IV U1816 ( .A(n1523), .Z(n1526) );
  XOR U1817 ( .A(n1527), .B(n1528), .Z(n1523) );
  ANDN U1818 ( .B(n1529), .A(n1530), .Z(n1527) );
  XNOR U1819 ( .A(b[223]), .B(n1528), .Z(n1529) );
  XNOR U1820 ( .A(b[223]), .B(n1530), .Z(c[223]) );
  XNOR U1821 ( .A(a[223]), .B(n1531), .Z(n1530) );
  IV U1822 ( .A(n1528), .Z(n1531) );
  XOR U1823 ( .A(n1532), .B(n1533), .Z(n1528) );
  ANDN U1824 ( .B(n1534), .A(n1535), .Z(n1532) );
  XNOR U1825 ( .A(b[222]), .B(n1533), .Z(n1534) );
  XNOR U1826 ( .A(b[222]), .B(n1535), .Z(c[222]) );
  XNOR U1827 ( .A(a[222]), .B(n1536), .Z(n1535) );
  IV U1828 ( .A(n1533), .Z(n1536) );
  XOR U1829 ( .A(n1537), .B(n1538), .Z(n1533) );
  ANDN U1830 ( .B(n1539), .A(n1540), .Z(n1537) );
  XNOR U1831 ( .A(b[221]), .B(n1538), .Z(n1539) );
  XNOR U1832 ( .A(b[221]), .B(n1540), .Z(c[221]) );
  XNOR U1833 ( .A(a[221]), .B(n1541), .Z(n1540) );
  IV U1834 ( .A(n1538), .Z(n1541) );
  XOR U1835 ( .A(n1542), .B(n1543), .Z(n1538) );
  ANDN U1836 ( .B(n1544), .A(n1545), .Z(n1542) );
  XNOR U1837 ( .A(b[220]), .B(n1543), .Z(n1544) );
  XNOR U1838 ( .A(b[220]), .B(n1545), .Z(c[220]) );
  XNOR U1839 ( .A(a[220]), .B(n1546), .Z(n1545) );
  IV U1840 ( .A(n1543), .Z(n1546) );
  XOR U1841 ( .A(n1547), .B(n1548), .Z(n1543) );
  ANDN U1842 ( .B(n1549), .A(n1550), .Z(n1547) );
  XNOR U1843 ( .A(b[219]), .B(n1548), .Z(n1549) );
  XNOR U1844 ( .A(b[21]), .B(n1551), .Z(c[21]) );
  XNOR U1845 ( .A(b[219]), .B(n1550), .Z(c[219]) );
  XNOR U1846 ( .A(a[219]), .B(n1552), .Z(n1550) );
  IV U1847 ( .A(n1548), .Z(n1552) );
  XOR U1848 ( .A(n1553), .B(n1554), .Z(n1548) );
  ANDN U1849 ( .B(n1555), .A(n1556), .Z(n1553) );
  XNOR U1850 ( .A(b[218]), .B(n1554), .Z(n1555) );
  XNOR U1851 ( .A(b[218]), .B(n1556), .Z(c[218]) );
  XNOR U1852 ( .A(a[218]), .B(n1557), .Z(n1556) );
  IV U1853 ( .A(n1554), .Z(n1557) );
  XOR U1854 ( .A(n1558), .B(n1559), .Z(n1554) );
  ANDN U1855 ( .B(n1560), .A(n1561), .Z(n1558) );
  XNOR U1856 ( .A(b[217]), .B(n1559), .Z(n1560) );
  XNOR U1857 ( .A(b[217]), .B(n1561), .Z(c[217]) );
  XNOR U1858 ( .A(a[217]), .B(n1562), .Z(n1561) );
  IV U1859 ( .A(n1559), .Z(n1562) );
  XOR U1860 ( .A(n1563), .B(n1564), .Z(n1559) );
  ANDN U1861 ( .B(n1565), .A(n1566), .Z(n1563) );
  XNOR U1862 ( .A(b[216]), .B(n1564), .Z(n1565) );
  XNOR U1863 ( .A(b[216]), .B(n1566), .Z(c[216]) );
  XNOR U1864 ( .A(a[216]), .B(n1567), .Z(n1566) );
  IV U1865 ( .A(n1564), .Z(n1567) );
  XOR U1866 ( .A(n1568), .B(n1569), .Z(n1564) );
  ANDN U1867 ( .B(n1570), .A(n1571), .Z(n1568) );
  XNOR U1868 ( .A(b[215]), .B(n1569), .Z(n1570) );
  XNOR U1869 ( .A(b[215]), .B(n1571), .Z(c[215]) );
  XNOR U1870 ( .A(a[215]), .B(n1572), .Z(n1571) );
  IV U1871 ( .A(n1569), .Z(n1572) );
  XOR U1872 ( .A(n1573), .B(n1574), .Z(n1569) );
  ANDN U1873 ( .B(n1575), .A(n1576), .Z(n1573) );
  XNOR U1874 ( .A(b[214]), .B(n1574), .Z(n1575) );
  XNOR U1875 ( .A(b[214]), .B(n1576), .Z(c[214]) );
  XNOR U1876 ( .A(a[214]), .B(n1577), .Z(n1576) );
  IV U1877 ( .A(n1574), .Z(n1577) );
  XOR U1878 ( .A(n1578), .B(n1579), .Z(n1574) );
  ANDN U1879 ( .B(n1580), .A(n1581), .Z(n1578) );
  XNOR U1880 ( .A(b[213]), .B(n1579), .Z(n1580) );
  XNOR U1881 ( .A(b[213]), .B(n1581), .Z(c[213]) );
  XNOR U1882 ( .A(a[213]), .B(n1582), .Z(n1581) );
  IV U1883 ( .A(n1579), .Z(n1582) );
  XOR U1884 ( .A(n1583), .B(n1584), .Z(n1579) );
  ANDN U1885 ( .B(n1585), .A(n1586), .Z(n1583) );
  XNOR U1886 ( .A(b[212]), .B(n1584), .Z(n1585) );
  XNOR U1887 ( .A(b[212]), .B(n1586), .Z(c[212]) );
  XNOR U1888 ( .A(a[212]), .B(n1587), .Z(n1586) );
  IV U1889 ( .A(n1584), .Z(n1587) );
  XOR U1890 ( .A(n1588), .B(n1589), .Z(n1584) );
  ANDN U1891 ( .B(n1590), .A(n1591), .Z(n1588) );
  XNOR U1892 ( .A(b[211]), .B(n1589), .Z(n1590) );
  XNOR U1893 ( .A(b[211]), .B(n1591), .Z(c[211]) );
  XNOR U1894 ( .A(a[211]), .B(n1592), .Z(n1591) );
  IV U1895 ( .A(n1589), .Z(n1592) );
  XOR U1896 ( .A(n1593), .B(n1594), .Z(n1589) );
  ANDN U1897 ( .B(n1595), .A(n1596), .Z(n1593) );
  XNOR U1898 ( .A(b[210]), .B(n1594), .Z(n1595) );
  XNOR U1899 ( .A(b[210]), .B(n1596), .Z(c[210]) );
  XNOR U1900 ( .A(a[210]), .B(n1597), .Z(n1596) );
  IV U1901 ( .A(n1594), .Z(n1597) );
  XOR U1902 ( .A(n1598), .B(n1599), .Z(n1594) );
  ANDN U1903 ( .B(n1600), .A(n1601), .Z(n1598) );
  XNOR U1904 ( .A(b[209]), .B(n1599), .Z(n1600) );
  XNOR U1905 ( .A(b[20]), .B(n1602), .Z(c[20]) );
  XNOR U1906 ( .A(b[209]), .B(n1601), .Z(c[209]) );
  XNOR U1907 ( .A(a[209]), .B(n1603), .Z(n1601) );
  IV U1908 ( .A(n1599), .Z(n1603) );
  XOR U1909 ( .A(n1604), .B(n1605), .Z(n1599) );
  ANDN U1910 ( .B(n1606), .A(n1607), .Z(n1604) );
  XNOR U1911 ( .A(b[208]), .B(n1605), .Z(n1606) );
  XNOR U1912 ( .A(b[208]), .B(n1607), .Z(c[208]) );
  XNOR U1913 ( .A(a[208]), .B(n1608), .Z(n1607) );
  IV U1914 ( .A(n1605), .Z(n1608) );
  XOR U1915 ( .A(n1609), .B(n1610), .Z(n1605) );
  ANDN U1916 ( .B(n1611), .A(n1612), .Z(n1609) );
  XNOR U1917 ( .A(b[207]), .B(n1610), .Z(n1611) );
  XNOR U1918 ( .A(b[207]), .B(n1612), .Z(c[207]) );
  XNOR U1919 ( .A(a[207]), .B(n1613), .Z(n1612) );
  IV U1920 ( .A(n1610), .Z(n1613) );
  XOR U1921 ( .A(n1614), .B(n1615), .Z(n1610) );
  ANDN U1922 ( .B(n1616), .A(n1617), .Z(n1614) );
  XNOR U1923 ( .A(b[206]), .B(n1615), .Z(n1616) );
  XNOR U1924 ( .A(b[206]), .B(n1617), .Z(c[206]) );
  XNOR U1925 ( .A(a[206]), .B(n1618), .Z(n1617) );
  IV U1926 ( .A(n1615), .Z(n1618) );
  XOR U1927 ( .A(n1619), .B(n1620), .Z(n1615) );
  ANDN U1928 ( .B(n1621), .A(n1622), .Z(n1619) );
  XNOR U1929 ( .A(b[205]), .B(n1620), .Z(n1621) );
  XNOR U1930 ( .A(b[205]), .B(n1622), .Z(c[205]) );
  XNOR U1931 ( .A(a[205]), .B(n1623), .Z(n1622) );
  IV U1932 ( .A(n1620), .Z(n1623) );
  XOR U1933 ( .A(n1624), .B(n1625), .Z(n1620) );
  ANDN U1934 ( .B(n1626), .A(n1627), .Z(n1624) );
  XNOR U1935 ( .A(b[204]), .B(n1625), .Z(n1626) );
  XNOR U1936 ( .A(b[204]), .B(n1627), .Z(c[204]) );
  XNOR U1937 ( .A(a[204]), .B(n1628), .Z(n1627) );
  IV U1938 ( .A(n1625), .Z(n1628) );
  XOR U1939 ( .A(n1629), .B(n1630), .Z(n1625) );
  ANDN U1940 ( .B(n1631), .A(n1632), .Z(n1629) );
  XNOR U1941 ( .A(b[203]), .B(n1630), .Z(n1631) );
  XNOR U1942 ( .A(b[203]), .B(n1632), .Z(c[203]) );
  XNOR U1943 ( .A(a[203]), .B(n1633), .Z(n1632) );
  IV U1944 ( .A(n1630), .Z(n1633) );
  XOR U1945 ( .A(n1634), .B(n1635), .Z(n1630) );
  ANDN U1946 ( .B(n1636), .A(n1637), .Z(n1634) );
  XNOR U1947 ( .A(b[202]), .B(n1635), .Z(n1636) );
  XNOR U1948 ( .A(b[202]), .B(n1637), .Z(c[202]) );
  XNOR U1949 ( .A(a[202]), .B(n1638), .Z(n1637) );
  IV U1950 ( .A(n1635), .Z(n1638) );
  XOR U1951 ( .A(n1639), .B(n1640), .Z(n1635) );
  ANDN U1952 ( .B(n1641), .A(n1642), .Z(n1639) );
  XNOR U1953 ( .A(b[201]), .B(n1640), .Z(n1641) );
  XNOR U1954 ( .A(b[201]), .B(n1642), .Z(c[201]) );
  XNOR U1955 ( .A(a[201]), .B(n1643), .Z(n1642) );
  IV U1956 ( .A(n1640), .Z(n1643) );
  XOR U1957 ( .A(n1644), .B(n1645), .Z(n1640) );
  ANDN U1958 ( .B(n1646), .A(n1647), .Z(n1644) );
  XNOR U1959 ( .A(b[200]), .B(n1645), .Z(n1646) );
  XNOR U1960 ( .A(b[200]), .B(n1647), .Z(c[200]) );
  XNOR U1961 ( .A(a[200]), .B(n1648), .Z(n1647) );
  IV U1962 ( .A(n1645), .Z(n1648) );
  XOR U1963 ( .A(n1649), .B(n1650), .Z(n1645) );
  ANDN U1964 ( .B(n1651), .A(n1652), .Z(n1649) );
  XNOR U1965 ( .A(b[199]), .B(n1650), .Z(n1651) );
  XNOR U1966 ( .A(b[1]), .B(n1653), .Z(c[1]) );
  XNOR U1967 ( .A(b[19]), .B(n1654), .Z(c[19]) );
  XNOR U1968 ( .A(b[199]), .B(n1652), .Z(c[199]) );
  XNOR U1969 ( .A(a[199]), .B(n1655), .Z(n1652) );
  IV U1970 ( .A(n1650), .Z(n1655) );
  XOR U1971 ( .A(n1656), .B(n1657), .Z(n1650) );
  ANDN U1972 ( .B(n1658), .A(n1659), .Z(n1656) );
  XNOR U1973 ( .A(b[198]), .B(n1657), .Z(n1658) );
  XNOR U1974 ( .A(b[198]), .B(n1659), .Z(c[198]) );
  XNOR U1975 ( .A(a[198]), .B(n1660), .Z(n1659) );
  IV U1976 ( .A(n1657), .Z(n1660) );
  XOR U1977 ( .A(n1661), .B(n1662), .Z(n1657) );
  ANDN U1978 ( .B(n1663), .A(n1664), .Z(n1661) );
  XNOR U1979 ( .A(b[197]), .B(n1662), .Z(n1663) );
  XNOR U1980 ( .A(b[197]), .B(n1664), .Z(c[197]) );
  XNOR U1981 ( .A(a[197]), .B(n1665), .Z(n1664) );
  IV U1982 ( .A(n1662), .Z(n1665) );
  XOR U1983 ( .A(n1666), .B(n1667), .Z(n1662) );
  ANDN U1984 ( .B(n1668), .A(n1669), .Z(n1666) );
  XNOR U1985 ( .A(b[196]), .B(n1667), .Z(n1668) );
  XNOR U1986 ( .A(b[196]), .B(n1669), .Z(c[196]) );
  XNOR U1987 ( .A(a[196]), .B(n1670), .Z(n1669) );
  IV U1988 ( .A(n1667), .Z(n1670) );
  XOR U1989 ( .A(n1671), .B(n1672), .Z(n1667) );
  ANDN U1990 ( .B(n1673), .A(n1674), .Z(n1671) );
  XNOR U1991 ( .A(b[195]), .B(n1672), .Z(n1673) );
  XNOR U1992 ( .A(b[195]), .B(n1674), .Z(c[195]) );
  XNOR U1993 ( .A(a[195]), .B(n1675), .Z(n1674) );
  IV U1994 ( .A(n1672), .Z(n1675) );
  XOR U1995 ( .A(n1676), .B(n1677), .Z(n1672) );
  ANDN U1996 ( .B(n1678), .A(n1679), .Z(n1676) );
  XNOR U1997 ( .A(b[194]), .B(n1677), .Z(n1678) );
  XNOR U1998 ( .A(b[194]), .B(n1679), .Z(c[194]) );
  XNOR U1999 ( .A(a[194]), .B(n1680), .Z(n1679) );
  IV U2000 ( .A(n1677), .Z(n1680) );
  XOR U2001 ( .A(n1681), .B(n1682), .Z(n1677) );
  ANDN U2002 ( .B(n1683), .A(n1684), .Z(n1681) );
  XNOR U2003 ( .A(b[193]), .B(n1682), .Z(n1683) );
  XNOR U2004 ( .A(b[193]), .B(n1684), .Z(c[193]) );
  XNOR U2005 ( .A(a[193]), .B(n1685), .Z(n1684) );
  IV U2006 ( .A(n1682), .Z(n1685) );
  XOR U2007 ( .A(n1686), .B(n1687), .Z(n1682) );
  ANDN U2008 ( .B(n1688), .A(n1689), .Z(n1686) );
  XNOR U2009 ( .A(b[192]), .B(n1687), .Z(n1688) );
  XNOR U2010 ( .A(b[192]), .B(n1689), .Z(c[192]) );
  XNOR U2011 ( .A(a[192]), .B(n1690), .Z(n1689) );
  IV U2012 ( .A(n1687), .Z(n1690) );
  XOR U2013 ( .A(n1691), .B(n1692), .Z(n1687) );
  ANDN U2014 ( .B(n1693), .A(n1694), .Z(n1691) );
  XNOR U2015 ( .A(b[191]), .B(n1692), .Z(n1693) );
  XNOR U2016 ( .A(b[191]), .B(n1694), .Z(c[191]) );
  XNOR U2017 ( .A(a[191]), .B(n1695), .Z(n1694) );
  IV U2018 ( .A(n1692), .Z(n1695) );
  XOR U2019 ( .A(n1696), .B(n1697), .Z(n1692) );
  ANDN U2020 ( .B(n1698), .A(n1699), .Z(n1696) );
  XNOR U2021 ( .A(b[190]), .B(n1697), .Z(n1698) );
  XNOR U2022 ( .A(b[190]), .B(n1699), .Z(c[190]) );
  XNOR U2023 ( .A(a[190]), .B(n1700), .Z(n1699) );
  IV U2024 ( .A(n1697), .Z(n1700) );
  XOR U2025 ( .A(n1701), .B(n1702), .Z(n1697) );
  ANDN U2026 ( .B(n1703), .A(n1704), .Z(n1701) );
  XNOR U2027 ( .A(b[189]), .B(n1702), .Z(n1703) );
  XNOR U2028 ( .A(b[18]), .B(n1705), .Z(c[18]) );
  XNOR U2029 ( .A(b[189]), .B(n1704), .Z(c[189]) );
  XNOR U2030 ( .A(a[189]), .B(n1706), .Z(n1704) );
  IV U2031 ( .A(n1702), .Z(n1706) );
  XOR U2032 ( .A(n1707), .B(n1708), .Z(n1702) );
  ANDN U2033 ( .B(n1709), .A(n1710), .Z(n1707) );
  XNOR U2034 ( .A(b[188]), .B(n1708), .Z(n1709) );
  XNOR U2035 ( .A(b[188]), .B(n1710), .Z(c[188]) );
  XNOR U2036 ( .A(a[188]), .B(n1711), .Z(n1710) );
  IV U2037 ( .A(n1708), .Z(n1711) );
  XOR U2038 ( .A(n1712), .B(n1713), .Z(n1708) );
  ANDN U2039 ( .B(n1714), .A(n1715), .Z(n1712) );
  XNOR U2040 ( .A(b[187]), .B(n1713), .Z(n1714) );
  XNOR U2041 ( .A(b[187]), .B(n1715), .Z(c[187]) );
  XNOR U2042 ( .A(a[187]), .B(n1716), .Z(n1715) );
  IV U2043 ( .A(n1713), .Z(n1716) );
  XOR U2044 ( .A(n1717), .B(n1718), .Z(n1713) );
  ANDN U2045 ( .B(n1719), .A(n1720), .Z(n1717) );
  XNOR U2046 ( .A(b[186]), .B(n1718), .Z(n1719) );
  XNOR U2047 ( .A(b[186]), .B(n1720), .Z(c[186]) );
  XNOR U2048 ( .A(a[186]), .B(n1721), .Z(n1720) );
  IV U2049 ( .A(n1718), .Z(n1721) );
  XOR U2050 ( .A(n1722), .B(n1723), .Z(n1718) );
  ANDN U2051 ( .B(n1724), .A(n1725), .Z(n1722) );
  XNOR U2052 ( .A(b[185]), .B(n1723), .Z(n1724) );
  XNOR U2053 ( .A(b[185]), .B(n1725), .Z(c[185]) );
  XNOR U2054 ( .A(a[185]), .B(n1726), .Z(n1725) );
  IV U2055 ( .A(n1723), .Z(n1726) );
  XOR U2056 ( .A(n1727), .B(n1728), .Z(n1723) );
  ANDN U2057 ( .B(n1729), .A(n1730), .Z(n1727) );
  XNOR U2058 ( .A(b[184]), .B(n1728), .Z(n1729) );
  XNOR U2059 ( .A(b[184]), .B(n1730), .Z(c[184]) );
  XNOR U2060 ( .A(a[184]), .B(n1731), .Z(n1730) );
  IV U2061 ( .A(n1728), .Z(n1731) );
  XOR U2062 ( .A(n1732), .B(n1733), .Z(n1728) );
  ANDN U2063 ( .B(n1734), .A(n1735), .Z(n1732) );
  XNOR U2064 ( .A(b[183]), .B(n1733), .Z(n1734) );
  XNOR U2065 ( .A(b[183]), .B(n1735), .Z(c[183]) );
  XNOR U2066 ( .A(a[183]), .B(n1736), .Z(n1735) );
  IV U2067 ( .A(n1733), .Z(n1736) );
  XOR U2068 ( .A(n1737), .B(n1738), .Z(n1733) );
  ANDN U2069 ( .B(n1739), .A(n1740), .Z(n1737) );
  XNOR U2070 ( .A(b[182]), .B(n1738), .Z(n1739) );
  XNOR U2071 ( .A(b[182]), .B(n1740), .Z(c[182]) );
  XNOR U2072 ( .A(a[182]), .B(n1741), .Z(n1740) );
  IV U2073 ( .A(n1738), .Z(n1741) );
  XOR U2074 ( .A(n1742), .B(n1743), .Z(n1738) );
  ANDN U2075 ( .B(n1744), .A(n1745), .Z(n1742) );
  XNOR U2076 ( .A(b[181]), .B(n1743), .Z(n1744) );
  XNOR U2077 ( .A(b[181]), .B(n1745), .Z(c[181]) );
  XNOR U2078 ( .A(a[181]), .B(n1746), .Z(n1745) );
  IV U2079 ( .A(n1743), .Z(n1746) );
  XOR U2080 ( .A(n1747), .B(n1748), .Z(n1743) );
  ANDN U2081 ( .B(n1749), .A(n1750), .Z(n1747) );
  XNOR U2082 ( .A(b[180]), .B(n1748), .Z(n1749) );
  XNOR U2083 ( .A(b[180]), .B(n1750), .Z(c[180]) );
  XNOR U2084 ( .A(a[180]), .B(n1751), .Z(n1750) );
  IV U2085 ( .A(n1748), .Z(n1751) );
  XOR U2086 ( .A(n1752), .B(n1753), .Z(n1748) );
  ANDN U2087 ( .B(n1754), .A(n1755), .Z(n1752) );
  XNOR U2088 ( .A(b[179]), .B(n1753), .Z(n1754) );
  XNOR U2089 ( .A(b[17]), .B(n1756), .Z(c[17]) );
  XNOR U2090 ( .A(b[179]), .B(n1755), .Z(c[179]) );
  XNOR U2091 ( .A(a[179]), .B(n1757), .Z(n1755) );
  IV U2092 ( .A(n1753), .Z(n1757) );
  XOR U2093 ( .A(n1758), .B(n1759), .Z(n1753) );
  ANDN U2094 ( .B(n1760), .A(n1761), .Z(n1758) );
  XNOR U2095 ( .A(b[178]), .B(n1759), .Z(n1760) );
  XNOR U2096 ( .A(b[178]), .B(n1761), .Z(c[178]) );
  XNOR U2097 ( .A(a[178]), .B(n1762), .Z(n1761) );
  IV U2098 ( .A(n1759), .Z(n1762) );
  XOR U2099 ( .A(n1763), .B(n1764), .Z(n1759) );
  ANDN U2100 ( .B(n1765), .A(n1766), .Z(n1763) );
  XNOR U2101 ( .A(b[177]), .B(n1764), .Z(n1765) );
  XNOR U2102 ( .A(b[177]), .B(n1766), .Z(c[177]) );
  XNOR U2103 ( .A(a[177]), .B(n1767), .Z(n1766) );
  IV U2104 ( .A(n1764), .Z(n1767) );
  XOR U2105 ( .A(n1768), .B(n1769), .Z(n1764) );
  ANDN U2106 ( .B(n1770), .A(n1771), .Z(n1768) );
  XNOR U2107 ( .A(b[176]), .B(n1769), .Z(n1770) );
  XNOR U2108 ( .A(b[176]), .B(n1771), .Z(c[176]) );
  XNOR U2109 ( .A(a[176]), .B(n1772), .Z(n1771) );
  IV U2110 ( .A(n1769), .Z(n1772) );
  XOR U2111 ( .A(n1773), .B(n1774), .Z(n1769) );
  ANDN U2112 ( .B(n1775), .A(n1776), .Z(n1773) );
  XNOR U2113 ( .A(b[175]), .B(n1774), .Z(n1775) );
  XNOR U2114 ( .A(b[175]), .B(n1776), .Z(c[175]) );
  XNOR U2115 ( .A(a[175]), .B(n1777), .Z(n1776) );
  IV U2116 ( .A(n1774), .Z(n1777) );
  XOR U2117 ( .A(n1778), .B(n1779), .Z(n1774) );
  ANDN U2118 ( .B(n1780), .A(n1781), .Z(n1778) );
  XNOR U2119 ( .A(b[174]), .B(n1779), .Z(n1780) );
  XNOR U2120 ( .A(b[174]), .B(n1781), .Z(c[174]) );
  XNOR U2121 ( .A(a[174]), .B(n1782), .Z(n1781) );
  IV U2122 ( .A(n1779), .Z(n1782) );
  XOR U2123 ( .A(n1783), .B(n1784), .Z(n1779) );
  ANDN U2124 ( .B(n1785), .A(n1786), .Z(n1783) );
  XNOR U2125 ( .A(b[173]), .B(n1784), .Z(n1785) );
  XNOR U2126 ( .A(b[173]), .B(n1786), .Z(c[173]) );
  XNOR U2127 ( .A(a[173]), .B(n1787), .Z(n1786) );
  IV U2128 ( .A(n1784), .Z(n1787) );
  XOR U2129 ( .A(n1788), .B(n1789), .Z(n1784) );
  ANDN U2130 ( .B(n1790), .A(n1791), .Z(n1788) );
  XNOR U2131 ( .A(b[172]), .B(n1789), .Z(n1790) );
  XNOR U2132 ( .A(b[172]), .B(n1791), .Z(c[172]) );
  XNOR U2133 ( .A(a[172]), .B(n1792), .Z(n1791) );
  IV U2134 ( .A(n1789), .Z(n1792) );
  XOR U2135 ( .A(n1793), .B(n1794), .Z(n1789) );
  ANDN U2136 ( .B(n1795), .A(n1796), .Z(n1793) );
  XNOR U2137 ( .A(b[171]), .B(n1794), .Z(n1795) );
  XNOR U2138 ( .A(b[171]), .B(n1796), .Z(c[171]) );
  XNOR U2139 ( .A(a[171]), .B(n1797), .Z(n1796) );
  IV U2140 ( .A(n1794), .Z(n1797) );
  XOR U2141 ( .A(n1798), .B(n1799), .Z(n1794) );
  ANDN U2142 ( .B(n1800), .A(n1801), .Z(n1798) );
  XNOR U2143 ( .A(b[170]), .B(n1799), .Z(n1800) );
  XNOR U2144 ( .A(b[170]), .B(n1801), .Z(c[170]) );
  XNOR U2145 ( .A(a[170]), .B(n1802), .Z(n1801) );
  IV U2146 ( .A(n1799), .Z(n1802) );
  XOR U2147 ( .A(n1803), .B(n1804), .Z(n1799) );
  ANDN U2148 ( .B(n1805), .A(n1806), .Z(n1803) );
  XNOR U2149 ( .A(b[169]), .B(n1804), .Z(n1805) );
  XNOR U2150 ( .A(b[16]), .B(n1807), .Z(c[16]) );
  XNOR U2151 ( .A(b[169]), .B(n1806), .Z(c[169]) );
  XNOR U2152 ( .A(a[169]), .B(n1808), .Z(n1806) );
  IV U2153 ( .A(n1804), .Z(n1808) );
  XOR U2154 ( .A(n1809), .B(n1810), .Z(n1804) );
  ANDN U2155 ( .B(n1811), .A(n1812), .Z(n1809) );
  XNOR U2156 ( .A(b[168]), .B(n1810), .Z(n1811) );
  XNOR U2157 ( .A(b[168]), .B(n1812), .Z(c[168]) );
  XNOR U2158 ( .A(a[168]), .B(n1813), .Z(n1812) );
  IV U2159 ( .A(n1810), .Z(n1813) );
  XOR U2160 ( .A(n1814), .B(n1815), .Z(n1810) );
  ANDN U2161 ( .B(n1816), .A(n1817), .Z(n1814) );
  XNOR U2162 ( .A(b[167]), .B(n1815), .Z(n1816) );
  XNOR U2163 ( .A(b[167]), .B(n1817), .Z(c[167]) );
  XNOR U2164 ( .A(a[167]), .B(n1818), .Z(n1817) );
  IV U2165 ( .A(n1815), .Z(n1818) );
  XOR U2166 ( .A(n1819), .B(n1820), .Z(n1815) );
  ANDN U2167 ( .B(n1821), .A(n1822), .Z(n1819) );
  XNOR U2168 ( .A(b[166]), .B(n1820), .Z(n1821) );
  XNOR U2169 ( .A(b[166]), .B(n1822), .Z(c[166]) );
  XNOR U2170 ( .A(a[166]), .B(n1823), .Z(n1822) );
  IV U2171 ( .A(n1820), .Z(n1823) );
  XOR U2172 ( .A(n1824), .B(n1825), .Z(n1820) );
  ANDN U2173 ( .B(n1826), .A(n1827), .Z(n1824) );
  XNOR U2174 ( .A(b[165]), .B(n1825), .Z(n1826) );
  XNOR U2175 ( .A(b[165]), .B(n1827), .Z(c[165]) );
  XNOR U2176 ( .A(a[165]), .B(n1828), .Z(n1827) );
  IV U2177 ( .A(n1825), .Z(n1828) );
  XOR U2178 ( .A(n1829), .B(n1830), .Z(n1825) );
  ANDN U2179 ( .B(n1831), .A(n1832), .Z(n1829) );
  XNOR U2180 ( .A(b[164]), .B(n1830), .Z(n1831) );
  XNOR U2181 ( .A(b[164]), .B(n1832), .Z(c[164]) );
  XNOR U2182 ( .A(a[164]), .B(n1833), .Z(n1832) );
  IV U2183 ( .A(n1830), .Z(n1833) );
  XOR U2184 ( .A(n1834), .B(n1835), .Z(n1830) );
  ANDN U2185 ( .B(n1836), .A(n1837), .Z(n1834) );
  XNOR U2186 ( .A(b[163]), .B(n1835), .Z(n1836) );
  XNOR U2187 ( .A(b[163]), .B(n1837), .Z(c[163]) );
  XNOR U2188 ( .A(a[163]), .B(n1838), .Z(n1837) );
  IV U2189 ( .A(n1835), .Z(n1838) );
  XOR U2190 ( .A(n1839), .B(n1840), .Z(n1835) );
  ANDN U2191 ( .B(n1841), .A(n1842), .Z(n1839) );
  XNOR U2192 ( .A(b[162]), .B(n1840), .Z(n1841) );
  XNOR U2193 ( .A(b[162]), .B(n1842), .Z(c[162]) );
  XNOR U2194 ( .A(a[162]), .B(n1843), .Z(n1842) );
  IV U2195 ( .A(n1840), .Z(n1843) );
  XOR U2196 ( .A(n1844), .B(n1845), .Z(n1840) );
  ANDN U2197 ( .B(n1846), .A(n1847), .Z(n1844) );
  XNOR U2198 ( .A(b[161]), .B(n1845), .Z(n1846) );
  XNOR U2199 ( .A(b[161]), .B(n1847), .Z(c[161]) );
  XNOR U2200 ( .A(a[161]), .B(n1848), .Z(n1847) );
  IV U2201 ( .A(n1845), .Z(n1848) );
  XOR U2202 ( .A(n1849), .B(n1850), .Z(n1845) );
  ANDN U2203 ( .B(n1851), .A(n1852), .Z(n1849) );
  XNOR U2204 ( .A(b[160]), .B(n1850), .Z(n1851) );
  XNOR U2205 ( .A(b[160]), .B(n1852), .Z(c[160]) );
  XNOR U2206 ( .A(a[160]), .B(n1853), .Z(n1852) );
  IV U2207 ( .A(n1850), .Z(n1853) );
  XOR U2208 ( .A(n1854), .B(n1855), .Z(n1850) );
  ANDN U2209 ( .B(n1856), .A(n1857), .Z(n1854) );
  XNOR U2210 ( .A(b[159]), .B(n1855), .Z(n1856) );
  XNOR U2211 ( .A(b[15]), .B(n1858), .Z(c[15]) );
  XNOR U2212 ( .A(b[159]), .B(n1857), .Z(c[159]) );
  XNOR U2213 ( .A(a[159]), .B(n1859), .Z(n1857) );
  IV U2214 ( .A(n1855), .Z(n1859) );
  XOR U2215 ( .A(n1860), .B(n1861), .Z(n1855) );
  ANDN U2216 ( .B(n1862), .A(n1863), .Z(n1860) );
  XNOR U2217 ( .A(b[158]), .B(n1861), .Z(n1862) );
  XNOR U2218 ( .A(b[158]), .B(n1863), .Z(c[158]) );
  XNOR U2219 ( .A(a[158]), .B(n1864), .Z(n1863) );
  IV U2220 ( .A(n1861), .Z(n1864) );
  XOR U2221 ( .A(n1865), .B(n1866), .Z(n1861) );
  ANDN U2222 ( .B(n1867), .A(n1868), .Z(n1865) );
  XNOR U2223 ( .A(b[157]), .B(n1866), .Z(n1867) );
  XNOR U2224 ( .A(b[157]), .B(n1868), .Z(c[157]) );
  XNOR U2225 ( .A(a[157]), .B(n1869), .Z(n1868) );
  IV U2226 ( .A(n1866), .Z(n1869) );
  XOR U2227 ( .A(n1870), .B(n1871), .Z(n1866) );
  ANDN U2228 ( .B(n1872), .A(n1873), .Z(n1870) );
  XNOR U2229 ( .A(b[156]), .B(n1871), .Z(n1872) );
  XNOR U2230 ( .A(b[156]), .B(n1873), .Z(c[156]) );
  XNOR U2231 ( .A(a[156]), .B(n1874), .Z(n1873) );
  IV U2232 ( .A(n1871), .Z(n1874) );
  XOR U2233 ( .A(n1875), .B(n1876), .Z(n1871) );
  ANDN U2234 ( .B(n1877), .A(n1878), .Z(n1875) );
  XNOR U2235 ( .A(b[155]), .B(n1876), .Z(n1877) );
  XNOR U2236 ( .A(b[155]), .B(n1878), .Z(c[155]) );
  XNOR U2237 ( .A(a[155]), .B(n1879), .Z(n1878) );
  IV U2238 ( .A(n1876), .Z(n1879) );
  XOR U2239 ( .A(n1880), .B(n1881), .Z(n1876) );
  ANDN U2240 ( .B(n1882), .A(n1883), .Z(n1880) );
  XNOR U2241 ( .A(b[154]), .B(n1881), .Z(n1882) );
  XNOR U2242 ( .A(b[154]), .B(n1883), .Z(c[154]) );
  XNOR U2243 ( .A(a[154]), .B(n1884), .Z(n1883) );
  IV U2244 ( .A(n1881), .Z(n1884) );
  XOR U2245 ( .A(n1885), .B(n1886), .Z(n1881) );
  ANDN U2246 ( .B(n1887), .A(n1888), .Z(n1885) );
  XNOR U2247 ( .A(b[153]), .B(n1886), .Z(n1887) );
  XNOR U2248 ( .A(b[153]), .B(n1888), .Z(c[153]) );
  XNOR U2249 ( .A(a[153]), .B(n1889), .Z(n1888) );
  IV U2250 ( .A(n1886), .Z(n1889) );
  XOR U2251 ( .A(n1890), .B(n1891), .Z(n1886) );
  ANDN U2252 ( .B(n1892), .A(n1893), .Z(n1890) );
  XNOR U2253 ( .A(b[152]), .B(n1891), .Z(n1892) );
  XNOR U2254 ( .A(b[152]), .B(n1893), .Z(c[152]) );
  XNOR U2255 ( .A(a[152]), .B(n1894), .Z(n1893) );
  IV U2256 ( .A(n1891), .Z(n1894) );
  XOR U2257 ( .A(n1895), .B(n1896), .Z(n1891) );
  ANDN U2258 ( .B(n1897), .A(n1898), .Z(n1895) );
  XNOR U2259 ( .A(b[151]), .B(n1896), .Z(n1897) );
  XNOR U2260 ( .A(b[151]), .B(n1898), .Z(c[151]) );
  XNOR U2261 ( .A(a[151]), .B(n1899), .Z(n1898) );
  IV U2262 ( .A(n1896), .Z(n1899) );
  XOR U2263 ( .A(n1900), .B(n1901), .Z(n1896) );
  ANDN U2264 ( .B(n1902), .A(n1903), .Z(n1900) );
  XNOR U2265 ( .A(b[150]), .B(n1901), .Z(n1902) );
  XNOR U2266 ( .A(b[150]), .B(n1903), .Z(c[150]) );
  XNOR U2267 ( .A(a[150]), .B(n1904), .Z(n1903) );
  IV U2268 ( .A(n1901), .Z(n1904) );
  XOR U2269 ( .A(n1905), .B(n1906), .Z(n1901) );
  ANDN U2270 ( .B(n1907), .A(n1908), .Z(n1905) );
  XNOR U2271 ( .A(b[149]), .B(n1906), .Z(n1907) );
  XNOR U2272 ( .A(b[14]), .B(n1909), .Z(c[14]) );
  XNOR U2273 ( .A(b[149]), .B(n1908), .Z(c[149]) );
  XNOR U2274 ( .A(a[149]), .B(n1910), .Z(n1908) );
  IV U2275 ( .A(n1906), .Z(n1910) );
  XOR U2276 ( .A(n1911), .B(n1912), .Z(n1906) );
  ANDN U2277 ( .B(n1913), .A(n1914), .Z(n1911) );
  XNOR U2278 ( .A(b[148]), .B(n1912), .Z(n1913) );
  XNOR U2279 ( .A(b[148]), .B(n1914), .Z(c[148]) );
  XNOR U2280 ( .A(a[148]), .B(n1915), .Z(n1914) );
  IV U2281 ( .A(n1912), .Z(n1915) );
  XOR U2282 ( .A(n1916), .B(n1917), .Z(n1912) );
  ANDN U2283 ( .B(n1918), .A(n1919), .Z(n1916) );
  XNOR U2284 ( .A(b[147]), .B(n1917), .Z(n1918) );
  XNOR U2285 ( .A(b[147]), .B(n1919), .Z(c[147]) );
  XNOR U2286 ( .A(a[147]), .B(n1920), .Z(n1919) );
  IV U2287 ( .A(n1917), .Z(n1920) );
  XOR U2288 ( .A(n1921), .B(n1922), .Z(n1917) );
  ANDN U2289 ( .B(n1923), .A(n1924), .Z(n1921) );
  XNOR U2290 ( .A(b[146]), .B(n1922), .Z(n1923) );
  XNOR U2291 ( .A(b[146]), .B(n1924), .Z(c[146]) );
  XNOR U2292 ( .A(a[146]), .B(n1925), .Z(n1924) );
  IV U2293 ( .A(n1922), .Z(n1925) );
  XOR U2294 ( .A(n1926), .B(n1927), .Z(n1922) );
  ANDN U2295 ( .B(n1928), .A(n1929), .Z(n1926) );
  XNOR U2296 ( .A(b[145]), .B(n1927), .Z(n1928) );
  XNOR U2297 ( .A(b[145]), .B(n1929), .Z(c[145]) );
  XNOR U2298 ( .A(a[145]), .B(n1930), .Z(n1929) );
  IV U2299 ( .A(n1927), .Z(n1930) );
  XOR U2300 ( .A(n1931), .B(n1932), .Z(n1927) );
  ANDN U2301 ( .B(n1933), .A(n1934), .Z(n1931) );
  XNOR U2302 ( .A(b[144]), .B(n1932), .Z(n1933) );
  XNOR U2303 ( .A(b[144]), .B(n1934), .Z(c[144]) );
  XNOR U2304 ( .A(a[144]), .B(n1935), .Z(n1934) );
  IV U2305 ( .A(n1932), .Z(n1935) );
  XOR U2306 ( .A(n1936), .B(n1937), .Z(n1932) );
  ANDN U2307 ( .B(n1938), .A(n1939), .Z(n1936) );
  XNOR U2308 ( .A(b[143]), .B(n1937), .Z(n1938) );
  XNOR U2309 ( .A(b[143]), .B(n1939), .Z(c[143]) );
  XNOR U2310 ( .A(a[143]), .B(n1940), .Z(n1939) );
  IV U2311 ( .A(n1937), .Z(n1940) );
  XOR U2312 ( .A(n1941), .B(n1942), .Z(n1937) );
  ANDN U2313 ( .B(n1943), .A(n1944), .Z(n1941) );
  XNOR U2314 ( .A(b[142]), .B(n1942), .Z(n1943) );
  XNOR U2315 ( .A(b[142]), .B(n1944), .Z(c[142]) );
  XNOR U2316 ( .A(a[142]), .B(n1945), .Z(n1944) );
  IV U2317 ( .A(n1942), .Z(n1945) );
  XOR U2318 ( .A(n1946), .B(n1947), .Z(n1942) );
  ANDN U2319 ( .B(n1948), .A(n1949), .Z(n1946) );
  XNOR U2320 ( .A(b[141]), .B(n1947), .Z(n1948) );
  XNOR U2321 ( .A(b[141]), .B(n1949), .Z(c[141]) );
  XNOR U2322 ( .A(a[141]), .B(n1950), .Z(n1949) );
  IV U2323 ( .A(n1947), .Z(n1950) );
  XOR U2324 ( .A(n1951), .B(n1952), .Z(n1947) );
  ANDN U2325 ( .B(n1953), .A(n1954), .Z(n1951) );
  XNOR U2326 ( .A(b[140]), .B(n1952), .Z(n1953) );
  XNOR U2327 ( .A(b[140]), .B(n1954), .Z(c[140]) );
  XNOR U2328 ( .A(a[140]), .B(n1955), .Z(n1954) );
  IV U2329 ( .A(n1952), .Z(n1955) );
  XOR U2330 ( .A(n1956), .B(n1957), .Z(n1952) );
  ANDN U2331 ( .B(n1958), .A(n1959), .Z(n1956) );
  XNOR U2332 ( .A(b[139]), .B(n1957), .Z(n1958) );
  XNOR U2333 ( .A(b[13]), .B(n1960), .Z(c[13]) );
  XNOR U2334 ( .A(b[139]), .B(n1959), .Z(c[139]) );
  XNOR U2335 ( .A(a[139]), .B(n1961), .Z(n1959) );
  IV U2336 ( .A(n1957), .Z(n1961) );
  XOR U2337 ( .A(n1962), .B(n1963), .Z(n1957) );
  ANDN U2338 ( .B(n1964), .A(n1965), .Z(n1962) );
  XNOR U2339 ( .A(b[138]), .B(n1963), .Z(n1964) );
  XNOR U2340 ( .A(b[138]), .B(n1965), .Z(c[138]) );
  XNOR U2341 ( .A(a[138]), .B(n1966), .Z(n1965) );
  IV U2342 ( .A(n1963), .Z(n1966) );
  XOR U2343 ( .A(n1967), .B(n1968), .Z(n1963) );
  ANDN U2344 ( .B(n1969), .A(n1970), .Z(n1967) );
  XNOR U2345 ( .A(b[137]), .B(n1968), .Z(n1969) );
  XNOR U2346 ( .A(b[137]), .B(n1970), .Z(c[137]) );
  XNOR U2347 ( .A(a[137]), .B(n1971), .Z(n1970) );
  IV U2348 ( .A(n1968), .Z(n1971) );
  XOR U2349 ( .A(n1972), .B(n1973), .Z(n1968) );
  ANDN U2350 ( .B(n1974), .A(n1975), .Z(n1972) );
  XNOR U2351 ( .A(b[136]), .B(n1973), .Z(n1974) );
  XNOR U2352 ( .A(b[136]), .B(n1975), .Z(c[136]) );
  XNOR U2353 ( .A(a[136]), .B(n1976), .Z(n1975) );
  IV U2354 ( .A(n1973), .Z(n1976) );
  XOR U2355 ( .A(n1977), .B(n1978), .Z(n1973) );
  ANDN U2356 ( .B(n1979), .A(n1980), .Z(n1977) );
  XNOR U2357 ( .A(b[135]), .B(n1978), .Z(n1979) );
  XNOR U2358 ( .A(b[135]), .B(n1980), .Z(c[135]) );
  XNOR U2359 ( .A(a[135]), .B(n1981), .Z(n1980) );
  IV U2360 ( .A(n1978), .Z(n1981) );
  XOR U2361 ( .A(n1982), .B(n1983), .Z(n1978) );
  ANDN U2362 ( .B(n1984), .A(n1985), .Z(n1982) );
  XNOR U2363 ( .A(b[134]), .B(n1983), .Z(n1984) );
  XNOR U2364 ( .A(b[134]), .B(n1985), .Z(c[134]) );
  XNOR U2365 ( .A(a[134]), .B(n1986), .Z(n1985) );
  IV U2366 ( .A(n1983), .Z(n1986) );
  XOR U2367 ( .A(n1987), .B(n1988), .Z(n1983) );
  ANDN U2368 ( .B(n1989), .A(n1990), .Z(n1987) );
  XNOR U2369 ( .A(b[133]), .B(n1988), .Z(n1989) );
  XNOR U2370 ( .A(b[133]), .B(n1990), .Z(c[133]) );
  XNOR U2371 ( .A(a[133]), .B(n1991), .Z(n1990) );
  IV U2372 ( .A(n1988), .Z(n1991) );
  XOR U2373 ( .A(n1992), .B(n1993), .Z(n1988) );
  ANDN U2374 ( .B(n1994), .A(n1995), .Z(n1992) );
  XNOR U2375 ( .A(b[132]), .B(n1993), .Z(n1994) );
  XNOR U2376 ( .A(b[132]), .B(n1995), .Z(c[132]) );
  XNOR U2377 ( .A(a[132]), .B(n1996), .Z(n1995) );
  IV U2378 ( .A(n1993), .Z(n1996) );
  XOR U2379 ( .A(n1997), .B(n1998), .Z(n1993) );
  ANDN U2380 ( .B(n1999), .A(n2000), .Z(n1997) );
  XNOR U2381 ( .A(b[131]), .B(n1998), .Z(n1999) );
  XNOR U2382 ( .A(b[131]), .B(n2000), .Z(c[131]) );
  XNOR U2383 ( .A(a[131]), .B(n2001), .Z(n2000) );
  IV U2384 ( .A(n1998), .Z(n2001) );
  XOR U2385 ( .A(n2002), .B(n2003), .Z(n1998) );
  ANDN U2386 ( .B(n2004), .A(n2005), .Z(n2002) );
  XNOR U2387 ( .A(b[130]), .B(n2003), .Z(n2004) );
  XNOR U2388 ( .A(b[130]), .B(n2005), .Z(c[130]) );
  XNOR U2389 ( .A(a[130]), .B(n2006), .Z(n2005) );
  IV U2390 ( .A(n2003), .Z(n2006) );
  XOR U2391 ( .A(n2007), .B(n2008), .Z(n2003) );
  ANDN U2392 ( .B(n2009), .A(n2010), .Z(n2007) );
  XNOR U2393 ( .A(b[129]), .B(n2008), .Z(n2009) );
  XNOR U2394 ( .A(b[12]), .B(n2011), .Z(c[12]) );
  XNOR U2395 ( .A(b[129]), .B(n2010), .Z(c[129]) );
  XNOR U2396 ( .A(a[129]), .B(n2012), .Z(n2010) );
  IV U2397 ( .A(n2008), .Z(n2012) );
  XOR U2398 ( .A(n2013), .B(n2014), .Z(n2008) );
  ANDN U2399 ( .B(n2015), .A(n2016), .Z(n2013) );
  XNOR U2400 ( .A(b[128]), .B(n2014), .Z(n2015) );
  XNOR U2401 ( .A(b[128]), .B(n2016), .Z(c[128]) );
  XNOR U2402 ( .A(a[128]), .B(n2017), .Z(n2016) );
  IV U2403 ( .A(n2014), .Z(n2017) );
  XOR U2404 ( .A(n2018), .B(n2019), .Z(n2014) );
  ANDN U2405 ( .B(n2020), .A(n2021), .Z(n2018) );
  XNOR U2406 ( .A(b[127]), .B(n2019), .Z(n2020) );
  XNOR U2407 ( .A(b[127]), .B(n2021), .Z(c[127]) );
  XNOR U2408 ( .A(a[127]), .B(n2022), .Z(n2021) );
  IV U2409 ( .A(n2019), .Z(n2022) );
  XOR U2410 ( .A(n2023), .B(n2024), .Z(n2019) );
  ANDN U2411 ( .B(n2025), .A(n2026), .Z(n2023) );
  XNOR U2412 ( .A(b[126]), .B(n2024), .Z(n2025) );
  XNOR U2413 ( .A(b[126]), .B(n2026), .Z(c[126]) );
  XNOR U2414 ( .A(a[126]), .B(n2027), .Z(n2026) );
  IV U2415 ( .A(n2024), .Z(n2027) );
  XOR U2416 ( .A(n2028), .B(n2029), .Z(n2024) );
  ANDN U2417 ( .B(n2030), .A(n2031), .Z(n2028) );
  XNOR U2418 ( .A(b[125]), .B(n2029), .Z(n2030) );
  XNOR U2419 ( .A(b[125]), .B(n2031), .Z(c[125]) );
  XNOR U2420 ( .A(a[125]), .B(n2032), .Z(n2031) );
  IV U2421 ( .A(n2029), .Z(n2032) );
  XOR U2422 ( .A(n2033), .B(n2034), .Z(n2029) );
  ANDN U2423 ( .B(n2035), .A(n2036), .Z(n2033) );
  XNOR U2424 ( .A(b[124]), .B(n2034), .Z(n2035) );
  XNOR U2425 ( .A(b[124]), .B(n2036), .Z(c[124]) );
  XNOR U2426 ( .A(a[124]), .B(n2037), .Z(n2036) );
  IV U2427 ( .A(n2034), .Z(n2037) );
  XOR U2428 ( .A(n2038), .B(n2039), .Z(n2034) );
  ANDN U2429 ( .B(n2040), .A(n2041), .Z(n2038) );
  XNOR U2430 ( .A(b[123]), .B(n2039), .Z(n2040) );
  XNOR U2431 ( .A(b[123]), .B(n2041), .Z(c[123]) );
  XNOR U2432 ( .A(a[123]), .B(n2042), .Z(n2041) );
  IV U2433 ( .A(n2039), .Z(n2042) );
  XOR U2434 ( .A(n2043), .B(n2044), .Z(n2039) );
  ANDN U2435 ( .B(n2045), .A(n2046), .Z(n2043) );
  XNOR U2436 ( .A(b[122]), .B(n2044), .Z(n2045) );
  XNOR U2437 ( .A(b[122]), .B(n2046), .Z(c[122]) );
  XNOR U2438 ( .A(a[122]), .B(n2047), .Z(n2046) );
  IV U2439 ( .A(n2044), .Z(n2047) );
  XOR U2440 ( .A(n2048), .B(n2049), .Z(n2044) );
  ANDN U2441 ( .B(n2050), .A(n2051), .Z(n2048) );
  XNOR U2442 ( .A(b[121]), .B(n2049), .Z(n2050) );
  XNOR U2443 ( .A(b[121]), .B(n2051), .Z(c[121]) );
  XNOR U2444 ( .A(a[121]), .B(n2052), .Z(n2051) );
  IV U2445 ( .A(n2049), .Z(n2052) );
  XOR U2446 ( .A(n2053), .B(n2054), .Z(n2049) );
  ANDN U2447 ( .B(n2055), .A(n2056), .Z(n2053) );
  XNOR U2448 ( .A(b[120]), .B(n2054), .Z(n2055) );
  XNOR U2449 ( .A(b[120]), .B(n2056), .Z(c[120]) );
  XNOR U2450 ( .A(a[120]), .B(n2057), .Z(n2056) );
  IV U2451 ( .A(n2054), .Z(n2057) );
  XOR U2452 ( .A(n2058), .B(n2059), .Z(n2054) );
  ANDN U2453 ( .B(n2060), .A(n2061), .Z(n2058) );
  XNOR U2454 ( .A(b[119]), .B(n2059), .Z(n2060) );
  XNOR U2455 ( .A(b[11]), .B(n2062), .Z(c[11]) );
  XNOR U2456 ( .A(b[119]), .B(n2061), .Z(c[119]) );
  XNOR U2457 ( .A(a[119]), .B(n2063), .Z(n2061) );
  IV U2458 ( .A(n2059), .Z(n2063) );
  XOR U2459 ( .A(n2064), .B(n2065), .Z(n2059) );
  ANDN U2460 ( .B(n2066), .A(n2067), .Z(n2064) );
  XNOR U2461 ( .A(b[118]), .B(n2065), .Z(n2066) );
  XNOR U2462 ( .A(b[118]), .B(n2067), .Z(c[118]) );
  XNOR U2463 ( .A(a[118]), .B(n2068), .Z(n2067) );
  IV U2464 ( .A(n2065), .Z(n2068) );
  XOR U2465 ( .A(n2069), .B(n2070), .Z(n2065) );
  ANDN U2466 ( .B(n2071), .A(n2072), .Z(n2069) );
  XNOR U2467 ( .A(b[117]), .B(n2070), .Z(n2071) );
  XNOR U2468 ( .A(b[117]), .B(n2072), .Z(c[117]) );
  XNOR U2469 ( .A(a[117]), .B(n2073), .Z(n2072) );
  IV U2470 ( .A(n2070), .Z(n2073) );
  XOR U2471 ( .A(n2074), .B(n2075), .Z(n2070) );
  ANDN U2472 ( .B(n2076), .A(n2077), .Z(n2074) );
  XNOR U2473 ( .A(b[116]), .B(n2075), .Z(n2076) );
  XNOR U2474 ( .A(b[116]), .B(n2077), .Z(c[116]) );
  XNOR U2475 ( .A(a[116]), .B(n2078), .Z(n2077) );
  IV U2476 ( .A(n2075), .Z(n2078) );
  XOR U2477 ( .A(n2079), .B(n2080), .Z(n2075) );
  ANDN U2478 ( .B(n2081), .A(n2082), .Z(n2079) );
  XNOR U2479 ( .A(b[115]), .B(n2080), .Z(n2081) );
  XNOR U2480 ( .A(b[115]), .B(n2082), .Z(c[115]) );
  XNOR U2481 ( .A(a[115]), .B(n2083), .Z(n2082) );
  IV U2482 ( .A(n2080), .Z(n2083) );
  XOR U2483 ( .A(n2084), .B(n2085), .Z(n2080) );
  ANDN U2484 ( .B(n2086), .A(n2087), .Z(n2084) );
  XNOR U2485 ( .A(b[114]), .B(n2085), .Z(n2086) );
  XNOR U2486 ( .A(b[114]), .B(n2087), .Z(c[114]) );
  XNOR U2487 ( .A(a[114]), .B(n2088), .Z(n2087) );
  IV U2488 ( .A(n2085), .Z(n2088) );
  XOR U2489 ( .A(n2089), .B(n2090), .Z(n2085) );
  ANDN U2490 ( .B(n2091), .A(n2092), .Z(n2089) );
  XNOR U2491 ( .A(b[113]), .B(n2090), .Z(n2091) );
  XNOR U2492 ( .A(b[113]), .B(n2092), .Z(c[113]) );
  XNOR U2493 ( .A(a[113]), .B(n2093), .Z(n2092) );
  IV U2494 ( .A(n2090), .Z(n2093) );
  XOR U2495 ( .A(n2094), .B(n2095), .Z(n2090) );
  ANDN U2496 ( .B(n2096), .A(n2097), .Z(n2094) );
  XNOR U2497 ( .A(b[112]), .B(n2095), .Z(n2096) );
  XNOR U2498 ( .A(b[112]), .B(n2097), .Z(c[112]) );
  XNOR U2499 ( .A(a[112]), .B(n2098), .Z(n2097) );
  IV U2500 ( .A(n2095), .Z(n2098) );
  XOR U2501 ( .A(n2099), .B(n2100), .Z(n2095) );
  ANDN U2502 ( .B(n2101), .A(n2102), .Z(n2099) );
  XNOR U2503 ( .A(b[111]), .B(n2100), .Z(n2101) );
  XNOR U2504 ( .A(b[111]), .B(n2102), .Z(c[111]) );
  XNOR U2505 ( .A(a[111]), .B(n2103), .Z(n2102) );
  IV U2506 ( .A(n2100), .Z(n2103) );
  XOR U2507 ( .A(n2104), .B(n2105), .Z(n2100) );
  ANDN U2508 ( .B(n2106), .A(n2107), .Z(n2104) );
  XNOR U2509 ( .A(b[110]), .B(n2105), .Z(n2106) );
  XNOR U2510 ( .A(b[110]), .B(n2107), .Z(c[110]) );
  XNOR U2511 ( .A(a[110]), .B(n2108), .Z(n2107) );
  IV U2512 ( .A(n2105), .Z(n2108) );
  XOR U2513 ( .A(n2109), .B(n2110), .Z(n2105) );
  ANDN U2514 ( .B(n2111), .A(n2112), .Z(n2109) );
  XNOR U2515 ( .A(b[109]), .B(n2110), .Z(n2111) );
  XNOR U2516 ( .A(b[10]), .B(n2113), .Z(c[10]) );
  XNOR U2517 ( .A(b[109]), .B(n2112), .Z(c[109]) );
  XNOR U2518 ( .A(a[109]), .B(n2114), .Z(n2112) );
  IV U2519 ( .A(n2110), .Z(n2114) );
  XOR U2520 ( .A(n2115), .B(n2116), .Z(n2110) );
  ANDN U2521 ( .B(n2117), .A(n2118), .Z(n2115) );
  XNOR U2522 ( .A(b[108]), .B(n2116), .Z(n2117) );
  XNOR U2523 ( .A(b[108]), .B(n2118), .Z(c[108]) );
  XNOR U2524 ( .A(a[108]), .B(n2119), .Z(n2118) );
  IV U2525 ( .A(n2116), .Z(n2119) );
  XOR U2526 ( .A(n2120), .B(n2121), .Z(n2116) );
  ANDN U2527 ( .B(n2122), .A(n2123), .Z(n2120) );
  XNOR U2528 ( .A(b[107]), .B(n2121), .Z(n2122) );
  XNOR U2529 ( .A(b[107]), .B(n2123), .Z(c[107]) );
  XNOR U2530 ( .A(a[107]), .B(n2124), .Z(n2123) );
  IV U2531 ( .A(n2121), .Z(n2124) );
  XOR U2532 ( .A(n2125), .B(n2126), .Z(n2121) );
  ANDN U2533 ( .B(n2127), .A(n2128), .Z(n2125) );
  XNOR U2534 ( .A(b[106]), .B(n2126), .Z(n2127) );
  XNOR U2535 ( .A(b[106]), .B(n2128), .Z(c[106]) );
  XNOR U2536 ( .A(a[106]), .B(n2129), .Z(n2128) );
  IV U2537 ( .A(n2126), .Z(n2129) );
  XOR U2538 ( .A(n2130), .B(n2131), .Z(n2126) );
  ANDN U2539 ( .B(n2132), .A(n2133), .Z(n2130) );
  XNOR U2540 ( .A(b[105]), .B(n2131), .Z(n2132) );
  XNOR U2541 ( .A(b[105]), .B(n2133), .Z(c[105]) );
  XNOR U2542 ( .A(a[105]), .B(n2134), .Z(n2133) );
  IV U2543 ( .A(n2131), .Z(n2134) );
  XOR U2544 ( .A(n2135), .B(n2136), .Z(n2131) );
  ANDN U2545 ( .B(n2137), .A(n2138), .Z(n2135) );
  XNOR U2546 ( .A(b[104]), .B(n2136), .Z(n2137) );
  XNOR U2547 ( .A(b[104]), .B(n2138), .Z(c[104]) );
  XNOR U2548 ( .A(a[104]), .B(n2139), .Z(n2138) );
  IV U2549 ( .A(n2136), .Z(n2139) );
  XOR U2550 ( .A(n2140), .B(n2141), .Z(n2136) );
  ANDN U2551 ( .B(n2142), .A(n2143), .Z(n2140) );
  XNOR U2552 ( .A(b[103]), .B(n2141), .Z(n2142) );
  XNOR U2553 ( .A(b[103]), .B(n2143), .Z(c[103]) );
  XNOR U2554 ( .A(a[103]), .B(n2144), .Z(n2143) );
  IV U2555 ( .A(n2141), .Z(n2144) );
  XOR U2556 ( .A(n2145), .B(n2146), .Z(n2141) );
  ANDN U2557 ( .B(n2147), .A(n2148), .Z(n2145) );
  XNOR U2558 ( .A(b[102]), .B(n2146), .Z(n2147) );
  XNOR U2559 ( .A(b[102]), .B(n2148), .Z(c[102]) );
  XNOR U2560 ( .A(a[102]), .B(n2149), .Z(n2148) );
  IV U2561 ( .A(n2146), .Z(n2149) );
  XOR U2562 ( .A(n2150), .B(n2151), .Z(n2146) );
  ANDN U2563 ( .B(n2152), .A(n2153), .Z(n2150) );
  XNOR U2564 ( .A(b[101]), .B(n2151), .Z(n2152) );
  XNOR U2565 ( .A(b[101]), .B(n2153), .Z(c[101]) );
  XNOR U2566 ( .A(a[101]), .B(n2154), .Z(n2153) );
  IV U2567 ( .A(n2151), .Z(n2154) );
  XOR U2568 ( .A(n2155), .B(n2156), .Z(n2151) );
  ANDN U2569 ( .B(n2157), .A(n2158), .Z(n2155) );
  XNOR U2570 ( .A(b[100]), .B(n2156), .Z(n2157) );
  XNOR U2571 ( .A(b[100]), .B(n2158), .Z(c[100]) );
  XNOR U2572 ( .A(a[100]), .B(n2159), .Z(n2158) );
  IV U2573 ( .A(n2156), .Z(n2159) );
  XOR U2574 ( .A(n2160), .B(n2161), .Z(n2156) );
  ANDN U2575 ( .B(n2162), .A(n7), .Z(n2160) );
  XNOR U2576 ( .A(a[99]), .B(n2163), .Z(n7) );
  IV U2577 ( .A(n2161), .Z(n2163) );
  XNOR U2578 ( .A(b[99]), .B(n2161), .Z(n2162) );
  XOR U2579 ( .A(n2164), .B(n2165), .Z(n2161) );
  ANDN U2580 ( .B(n2166), .A(n8), .Z(n2164) );
  XNOR U2581 ( .A(a[98]), .B(n2167), .Z(n8) );
  IV U2582 ( .A(n2165), .Z(n2167) );
  XNOR U2583 ( .A(b[98]), .B(n2165), .Z(n2166) );
  XOR U2584 ( .A(n2168), .B(n2169), .Z(n2165) );
  ANDN U2585 ( .B(n2170), .A(n9), .Z(n2168) );
  XNOR U2586 ( .A(a[97]), .B(n2171), .Z(n9) );
  IV U2587 ( .A(n2169), .Z(n2171) );
  XNOR U2588 ( .A(b[97]), .B(n2169), .Z(n2170) );
  XOR U2589 ( .A(n2172), .B(n2173), .Z(n2169) );
  ANDN U2590 ( .B(n2174), .A(n10), .Z(n2172) );
  XNOR U2591 ( .A(a[96]), .B(n2175), .Z(n10) );
  IV U2592 ( .A(n2173), .Z(n2175) );
  XNOR U2593 ( .A(b[96]), .B(n2173), .Z(n2174) );
  XOR U2594 ( .A(n2176), .B(n2177), .Z(n2173) );
  ANDN U2595 ( .B(n2178), .A(n11), .Z(n2176) );
  XNOR U2596 ( .A(a[95]), .B(n2179), .Z(n11) );
  IV U2597 ( .A(n2177), .Z(n2179) );
  XNOR U2598 ( .A(b[95]), .B(n2177), .Z(n2178) );
  XOR U2599 ( .A(n2180), .B(n2181), .Z(n2177) );
  ANDN U2600 ( .B(n2182), .A(n12), .Z(n2180) );
  XNOR U2601 ( .A(a[94]), .B(n2183), .Z(n12) );
  IV U2602 ( .A(n2181), .Z(n2183) );
  XNOR U2603 ( .A(b[94]), .B(n2181), .Z(n2182) );
  XOR U2604 ( .A(n2184), .B(n2185), .Z(n2181) );
  ANDN U2605 ( .B(n2186), .A(n13), .Z(n2184) );
  XNOR U2606 ( .A(a[93]), .B(n2187), .Z(n13) );
  IV U2607 ( .A(n2185), .Z(n2187) );
  XNOR U2608 ( .A(b[93]), .B(n2185), .Z(n2186) );
  XOR U2609 ( .A(n2188), .B(n2189), .Z(n2185) );
  ANDN U2610 ( .B(n2190), .A(n14), .Z(n2188) );
  XNOR U2611 ( .A(a[92]), .B(n2191), .Z(n14) );
  IV U2612 ( .A(n2189), .Z(n2191) );
  XNOR U2613 ( .A(b[92]), .B(n2189), .Z(n2190) );
  XOR U2614 ( .A(n2192), .B(n2193), .Z(n2189) );
  ANDN U2615 ( .B(n2194), .A(n15), .Z(n2192) );
  XNOR U2616 ( .A(a[91]), .B(n2195), .Z(n15) );
  IV U2617 ( .A(n2193), .Z(n2195) );
  XNOR U2618 ( .A(b[91]), .B(n2193), .Z(n2194) );
  XOR U2619 ( .A(n2196), .B(n2197), .Z(n2193) );
  ANDN U2620 ( .B(n2198), .A(n16), .Z(n2196) );
  XNOR U2621 ( .A(a[90]), .B(n2199), .Z(n16) );
  IV U2622 ( .A(n2197), .Z(n2199) );
  XNOR U2623 ( .A(b[90]), .B(n2197), .Z(n2198) );
  XOR U2624 ( .A(n2200), .B(n2201), .Z(n2197) );
  ANDN U2625 ( .B(n2202), .A(n18), .Z(n2200) );
  XNOR U2626 ( .A(a[89]), .B(n2203), .Z(n18) );
  IV U2627 ( .A(n2201), .Z(n2203) );
  XNOR U2628 ( .A(b[89]), .B(n2201), .Z(n2202) );
  XOR U2629 ( .A(n2204), .B(n2205), .Z(n2201) );
  ANDN U2630 ( .B(n2206), .A(n19), .Z(n2204) );
  XNOR U2631 ( .A(a[88]), .B(n2207), .Z(n19) );
  IV U2632 ( .A(n2205), .Z(n2207) );
  XNOR U2633 ( .A(b[88]), .B(n2205), .Z(n2206) );
  XOR U2634 ( .A(n2208), .B(n2209), .Z(n2205) );
  ANDN U2635 ( .B(n2210), .A(n20), .Z(n2208) );
  XNOR U2636 ( .A(a[87]), .B(n2211), .Z(n20) );
  IV U2637 ( .A(n2209), .Z(n2211) );
  XNOR U2638 ( .A(b[87]), .B(n2209), .Z(n2210) );
  XOR U2639 ( .A(n2212), .B(n2213), .Z(n2209) );
  ANDN U2640 ( .B(n2214), .A(n21), .Z(n2212) );
  XNOR U2641 ( .A(a[86]), .B(n2215), .Z(n21) );
  IV U2642 ( .A(n2213), .Z(n2215) );
  XNOR U2643 ( .A(b[86]), .B(n2213), .Z(n2214) );
  XOR U2644 ( .A(n2216), .B(n2217), .Z(n2213) );
  ANDN U2645 ( .B(n2218), .A(n22), .Z(n2216) );
  XNOR U2646 ( .A(a[85]), .B(n2219), .Z(n22) );
  IV U2647 ( .A(n2217), .Z(n2219) );
  XNOR U2648 ( .A(b[85]), .B(n2217), .Z(n2218) );
  XOR U2649 ( .A(n2220), .B(n2221), .Z(n2217) );
  ANDN U2650 ( .B(n2222), .A(n23), .Z(n2220) );
  XNOR U2651 ( .A(a[84]), .B(n2223), .Z(n23) );
  IV U2652 ( .A(n2221), .Z(n2223) );
  XNOR U2653 ( .A(b[84]), .B(n2221), .Z(n2222) );
  XOR U2654 ( .A(n2224), .B(n2225), .Z(n2221) );
  ANDN U2655 ( .B(n2226), .A(n24), .Z(n2224) );
  XNOR U2656 ( .A(a[83]), .B(n2227), .Z(n24) );
  IV U2657 ( .A(n2225), .Z(n2227) );
  XNOR U2658 ( .A(b[83]), .B(n2225), .Z(n2226) );
  XOR U2659 ( .A(n2228), .B(n2229), .Z(n2225) );
  ANDN U2660 ( .B(n2230), .A(n25), .Z(n2228) );
  XNOR U2661 ( .A(a[82]), .B(n2231), .Z(n25) );
  IV U2662 ( .A(n2229), .Z(n2231) );
  XNOR U2663 ( .A(b[82]), .B(n2229), .Z(n2230) );
  XOR U2664 ( .A(n2232), .B(n2233), .Z(n2229) );
  ANDN U2665 ( .B(n2234), .A(n26), .Z(n2232) );
  XNOR U2666 ( .A(a[81]), .B(n2235), .Z(n26) );
  IV U2667 ( .A(n2233), .Z(n2235) );
  XNOR U2668 ( .A(b[81]), .B(n2233), .Z(n2234) );
  XOR U2669 ( .A(n2236), .B(n2237), .Z(n2233) );
  ANDN U2670 ( .B(n2238), .A(n27), .Z(n2236) );
  XNOR U2671 ( .A(a[80]), .B(n2239), .Z(n27) );
  IV U2672 ( .A(n2237), .Z(n2239) );
  XNOR U2673 ( .A(b[80]), .B(n2237), .Z(n2238) );
  XOR U2674 ( .A(n2240), .B(n2241), .Z(n2237) );
  ANDN U2675 ( .B(n2242), .A(n29), .Z(n2240) );
  XNOR U2676 ( .A(a[79]), .B(n2243), .Z(n29) );
  IV U2677 ( .A(n2241), .Z(n2243) );
  XNOR U2678 ( .A(b[79]), .B(n2241), .Z(n2242) );
  XOR U2679 ( .A(n2244), .B(n2245), .Z(n2241) );
  ANDN U2680 ( .B(n2246), .A(n30), .Z(n2244) );
  XNOR U2681 ( .A(a[78]), .B(n2247), .Z(n30) );
  IV U2682 ( .A(n2245), .Z(n2247) );
  XNOR U2683 ( .A(b[78]), .B(n2245), .Z(n2246) );
  XOR U2684 ( .A(n2248), .B(n2249), .Z(n2245) );
  ANDN U2685 ( .B(n2250), .A(n31), .Z(n2248) );
  XNOR U2686 ( .A(a[77]), .B(n2251), .Z(n31) );
  IV U2687 ( .A(n2249), .Z(n2251) );
  XNOR U2688 ( .A(b[77]), .B(n2249), .Z(n2250) );
  XOR U2689 ( .A(n2252), .B(n2253), .Z(n2249) );
  ANDN U2690 ( .B(n2254), .A(n32), .Z(n2252) );
  XNOR U2691 ( .A(a[76]), .B(n2255), .Z(n32) );
  IV U2692 ( .A(n2253), .Z(n2255) );
  XNOR U2693 ( .A(b[76]), .B(n2253), .Z(n2254) );
  XOR U2694 ( .A(n2256), .B(n2257), .Z(n2253) );
  ANDN U2695 ( .B(n2258), .A(n33), .Z(n2256) );
  XNOR U2696 ( .A(a[75]), .B(n2259), .Z(n33) );
  IV U2697 ( .A(n2257), .Z(n2259) );
  XNOR U2698 ( .A(b[75]), .B(n2257), .Z(n2258) );
  XOR U2699 ( .A(n2260), .B(n2261), .Z(n2257) );
  ANDN U2700 ( .B(n2262), .A(n34), .Z(n2260) );
  XNOR U2701 ( .A(a[74]), .B(n2263), .Z(n34) );
  IV U2702 ( .A(n2261), .Z(n2263) );
  XNOR U2703 ( .A(b[74]), .B(n2261), .Z(n2262) );
  XOR U2704 ( .A(n2264), .B(n2265), .Z(n2261) );
  ANDN U2705 ( .B(n2266), .A(n35), .Z(n2264) );
  XNOR U2706 ( .A(a[73]), .B(n2267), .Z(n35) );
  IV U2707 ( .A(n2265), .Z(n2267) );
  XNOR U2708 ( .A(b[73]), .B(n2265), .Z(n2266) );
  XOR U2709 ( .A(n2268), .B(n2269), .Z(n2265) );
  ANDN U2710 ( .B(n2270), .A(n36), .Z(n2268) );
  XNOR U2711 ( .A(a[72]), .B(n2271), .Z(n36) );
  IV U2712 ( .A(n2269), .Z(n2271) );
  XNOR U2713 ( .A(b[72]), .B(n2269), .Z(n2270) );
  XOR U2714 ( .A(n2272), .B(n2273), .Z(n2269) );
  ANDN U2715 ( .B(n2274), .A(n37), .Z(n2272) );
  XNOR U2716 ( .A(a[71]), .B(n2275), .Z(n37) );
  IV U2717 ( .A(n2273), .Z(n2275) );
  XNOR U2718 ( .A(b[71]), .B(n2273), .Z(n2274) );
  XOR U2719 ( .A(n2276), .B(n2277), .Z(n2273) );
  ANDN U2720 ( .B(n2278), .A(n38), .Z(n2276) );
  XNOR U2721 ( .A(a[70]), .B(n2279), .Z(n38) );
  IV U2722 ( .A(n2277), .Z(n2279) );
  XNOR U2723 ( .A(b[70]), .B(n2277), .Z(n2278) );
  XOR U2724 ( .A(n2280), .B(n2281), .Z(n2277) );
  ANDN U2725 ( .B(n2282), .A(n40), .Z(n2280) );
  XNOR U2726 ( .A(a[69]), .B(n2283), .Z(n40) );
  IV U2727 ( .A(n2281), .Z(n2283) );
  XNOR U2728 ( .A(b[69]), .B(n2281), .Z(n2282) );
  XOR U2729 ( .A(n2284), .B(n2285), .Z(n2281) );
  ANDN U2730 ( .B(n2286), .A(n41), .Z(n2284) );
  XNOR U2731 ( .A(a[68]), .B(n2287), .Z(n41) );
  IV U2732 ( .A(n2285), .Z(n2287) );
  XNOR U2733 ( .A(b[68]), .B(n2285), .Z(n2286) );
  XOR U2734 ( .A(n2288), .B(n2289), .Z(n2285) );
  ANDN U2735 ( .B(n2290), .A(n42), .Z(n2288) );
  XNOR U2736 ( .A(a[67]), .B(n2291), .Z(n42) );
  IV U2737 ( .A(n2289), .Z(n2291) );
  XNOR U2738 ( .A(b[67]), .B(n2289), .Z(n2290) );
  XOR U2739 ( .A(n2292), .B(n2293), .Z(n2289) );
  ANDN U2740 ( .B(n2294), .A(n43), .Z(n2292) );
  XNOR U2741 ( .A(a[66]), .B(n2295), .Z(n43) );
  IV U2742 ( .A(n2293), .Z(n2295) );
  XNOR U2743 ( .A(b[66]), .B(n2293), .Z(n2294) );
  XOR U2744 ( .A(n2296), .B(n2297), .Z(n2293) );
  ANDN U2745 ( .B(n2298), .A(n44), .Z(n2296) );
  XNOR U2746 ( .A(a[65]), .B(n2299), .Z(n44) );
  IV U2747 ( .A(n2297), .Z(n2299) );
  XNOR U2748 ( .A(b[65]), .B(n2297), .Z(n2298) );
  XOR U2749 ( .A(n2300), .B(n2301), .Z(n2297) );
  ANDN U2750 ( .B(n2302), .A(n45), .Z(n2300) );
  XNOR U2751 ( .A(a[64]), .B(n2303), .Z(n45) );
  IV U2752 ( .A(n2301), .Z(n2303) );
  XNOR U2753 ( .A(b[64]), .B(n2301), .Z(n2302) );
  XOR U2754 ( .A(n2304), .B(n2305), .Z(n2301) );
  ANDN U2755 ( .B(n2306), .A(n46), .Z(n2304) );
  XNOR U2756 ( .A(a[63]), .B(n2307), .Z(n46) );
  IV U2757 ( .A(n2305), .Z(n2307) );
  XNOR U2758 ( .A(b[63]), .B(n2305), .Z(n2306) );
  XOR U2759 ( .A(n2308), .B(n2309), .Z(n2305) );
  ANDN U2760 ( .B(n2310), .A(n47), .Z(n2308) );
  XNOR U2761 ( .A(a[62]), .B(n2311), .Z(n47) );
  IV U2762 ( .A(n2309), .Z(n2311) );
  XNOR U2763 ( .A(b[62]), .B(n2309), .Z(n2310) );
  XOR U2764 ( .A(n2312), .B(n2313), .Z(n2309) );
  ANDN U2765 ( .B(n2314), .A(n48), .Z(n2312) );
  XNOR U2766 ( .A(a[61]), .B(n2315), .Z(n48) );
  IV U2767 ( .A(n2313), .Z(n2315) );
  XNOR U2768 ( .A(b[61]), .B(n2313), .Z(n2314) );
  XOR U2769 ( .A(n2316), .B(n2317), .Z(n2313) );
  ANDN U2770 ( .B(n2318), .A(n49), .Z(n2316) );
  XNOR U2771 ( .A(a[60]), .B(n2319), .Z(n49) );
  IV U2772 ( .A(n2317), .Z(n2319) );
  XNOR U2773 ( .A(b[60]), .B(n2317), .Z(n2318) );
  XOR U2774 ( .A(n2320), .B(n2321), .Z(n2317) );
  ANDN U2775 ( .B(n2322), .A(n51), .Z(n2320) );
  XNOR U2776 ( .A(a[59]), .B(n2323), .Z(n51) );
  IV U2777 ( .A(n2321), .Z(n2323) );
  XNOR U2778 ( .A(b[59]), .B(n2321), .Z(n2322) );
  XOR U2779 ( .A(n2324), .B(n2325), .Z(n2321) );
  ANDN U2780 ( .B(n2326), .A(n52), .Z(n2324) );
  XNOR U2781 ( .A(a[58]), .B(n2327), .Z(n52) );
  IV U2782 ( .A(n2325), .Z(n2327) );
  XNOR U2783 ( .A(b[58]), .B(n2325), .Z(n2326) );
  XOR U2784 ( .A(n2328), .B(n2329), .Z(n2325) );
  ANDN U2785 ( .B(n2330), .A(n53), .Z(n2328) );
  XNOR U2786 ( .A(a[57]), .B(n2331), .Z(n53) );
  IV U2787 ( .A(n2329), .Z(n2331) );
  XNOR U2788 ( .A(b[57]), .B(n2329), .Z(n2330) );
  XOR U2789 ( .A(n2332), .B(n2333), .Z(n2329) );
  ANDN U2790 ( .B(n2334), .A(n54), .Z(n2332) );
  XNOR U2791 ( .A(a[56]), .B(n2335), .Z(n54) );
  IV U2792 ( .A(n2333), .Z(n2335) );
  XNOR U2793 ( .A(b[56]), .B(n2333), .Z(n2334) );
  XOR U2794 ( .A(n2336), .B(n2337), .Z(n2333) );
  ANDN U2795 ( .B(n2338), .A(n55), .Z(n2336) );
  XNOR U2796 ( .A(a[55]), .B(n2339), .Z(n55) );
  IV U2797 ( .A(n2337), .Z(n2339) );
  XNOR U2798 ( .A(b[55]), .B(n2337), .Z(n2338) );
  XOR U2799 ( .A(n2340), .B(n2341), .Z(n2337) );
  ANDN U2800 ( .B(n2342), .A(n56), .Z(n2340) );
  XNOR U2801 ( .A(a[54]), .B(n2343), .Z(n56) );
  IV U2802 ( .A(n2341), .Z(n2343) );
  XNOR U2803 ( .A(b[54]), .B(n2341), .Z(n2342) );
  XOR U2804 ( .A(n2344), .B(n2345), .Z(n2341) );
  ANDN U2805 ( .B(n2346), .A(n57), .Z(n2344) );
  XNOR U2806 ( .A(a[53]), .B(n2347), .Z(n57) );
  IV U2807 ( .A(n2345), .Z(n2347) );
  XNOR U2808 ( .A(b[53]), .B(n2345), .Z(n2346) );
  XOR U2809 ( .A(n2348), .B(n2349), .Z(n2345) );
  ANDN U2810 ( .B(n2350), .A(n58), .Z(n2348) );
  XNOR U2811 ( .A(a[52]), .B(n2351), .Z(n58) );
  IV U2812 ( .A(n2349), .Z(n2351) );
  XNOR U2813 ( .A(b[52]), .B(n2349), .Z(n2350) );
  XOR U2814 ( .A(n2352), .B(n2353), .Z(n2349) );
  ANDN U2815 ( .B(n2354), .A(n59), .Z(n2352) );
  XNOR U2816 ( .A(a[51]), .B(n2355), .Z(n59) );
  IV U2817 ( .A(n2353), .Z(n2355) );
  XNOR U2818 ( .A(b[51]), .B(n2353), .Z(n2354) );
  XOR U2819 ( .A(n2356), .B(n2357), .Z(n2353) );
  ANDN U2820 ( .B(n2358), .A(n69), .Z(n2356) );
  XNOR U2821 ( .A(a[50]), .B(n2359), .Z(n69) );
  IV U2822 ( .A(n2357), .Z(n2359) );
  XNOR U2823 ( .A(b[50]), .B(n2357), .Z(n2358) );
  XOR U2824 ( .A(n2360), .B(n2361), .Z(n2357) );
  ANDN U2825 ( .B(n2362), .A(n121), .Z(n2360) );
  XNOR U2826 ( .A(a[49]), .B(n2363), .Z(n121) );
  IV U2827 ( .A(n2361), .Z(n2363) );
  XNOR U2828 ( .A(b[49]), .B(n2361), .Z(n2362) );
  XOR U2829 ( .A(n2364), .B(n2365), .Z(n2361) );
  ANDN U2830 ( .B(n2366), .A(n172), .Z(n2364) );
  XNOR U2831 ( .A(a[48]), .B(n2367), .Z(n172) );
  IV U2832 ( .A(n2365), .Z(n2367) );
  XNOR U2833 ( .A(b[48]), .B(n2365), .Z(n2366) );
  XOR U2834 ( .A(n2368), .B(n2369), .Z(n2365) );
  ANDN U2835 ( .B(n2370), .A(n223), .Z(n2368) );
  XNOR U2836 ( .A(a[47]), .B(n2371), .Z(n223) );
  IV U2837 ( .A(n2369), .Z(n2371) );
  XNOR U2838 ( .A(b[47]), .B(n2369), .Z(n2370) );
  XOR U2839 ( .A(n2372), .B(n2373), .Z(n2369) );
  ANDN U2840 ( .B(n2374), .A(n274), .Z(n2372) );
  XNOR U2841 ( .A(a[46]), .B(n2375), .Z(n274) );
  IV U2842 ( .A(n2373), .Z(n2375) );
  XNOR U2843 ( .A(b[46]), .B(n2373), .Z(n2374) );
  XOR U2844 ( .A(n2376), .B(n2377), .Z(n2373) );
  ANDN U2845 ( .B(n2378), .A(n325), .Z(n2376) );
  XNOR U2846 ( .A(a[45]), .B(n2379), .Z(n325) );
  IV U2847 ( .A(n2377), .Z(n2379) );
  XNOR U2848 ( .A(b[45]), .B(n2377), .Z(n2378) );
  XOR U2849 ( .A(n2380), .B(n2381), .Z(n2377) );
  ANDN U2850 ( .B(n2382), .A(n376), .Z(n2380) );
  XNOR U2851 ( .A(a[44]), .B(n2383), .Z(n376) );
  IV U2852 ( .A(n2381), .Z(n2383) );
  XNOR U2853 ( .A(b[44]), .B(n2381), .Z(n2382) );
  XOR U2854 ( .A(n2384), .B(n2385), .Z(n2381) );
  ANDN U2855 ( .B(n2386), .A(n427), .Z(n2384) );
  XNOR U2856 ( .A(a[43]), .B(n2387), .Z(n427) );
  IV U2857 ( .A(n2385), .Z(n2387) );
  XNOR U2858 ( .A(b[43]), .B(n2385), .Z(n2386) );
  XOR U2859 ( .A(n2388), .B(n2389), .Z(n2385) );
  ANDN U2860 ( .B(n2390), .A(n478), .Z(n2388) );
  XNOR U2861 ( .A(a[42]), .B(n2391), .Z(n478) );
  IV U2862 ( .A(n2389), .Z(n2391) );
  XNOR U2863 ( .A(b[42]), .B(n2389), .Z(n2390) );
  XOR U2864 ( .A(n2392), .B(n2393), .Z(n2389) );
  ANDN U2865 ( .B(n2394), .A(n529), .Z(n2392) );
  XNOR U2866 ( .A(a[41]), .B(n2395), .Z(n529) );
  IV U2867 ( .A(n2393), .Z(n2395) );
  XNOR U2868 ( .A(b[41]), .B(n2393), .Z(n2394) );
  XOR U2869 ( .A(n2396), .B(n2397), .Z(n2393) );
  ANDN U2870 ( .B(n2398), .A(n580), .Z(n2396) );
  XNOR U2871 ( .A(a[40]), .B(n2399), .Z(n580) );
  IV U2872 ( .A(n2397), .Z(n2399) );
  XNOR U2873 ( .A(b[40]), .B(n2397), .Z(n2398) );
  XOR U2874 ( .A(n2400), .B(n2401), .Z(n2397) );
  ANDN U2875 ( .B(n2402), .A(n632), .Z(n2400) );
  XNOR U2876 ( .A(a[39]), .B(n2403), .Z(n632) );
  IV U2877 ( .A(n2401), .Z(n2403) );
  XNOR U2878 ( .A(b[39]), .B(n2401), .Z(n2402) );
  XOR U2879 ( .A(n2404), .B(n2405), .Z(n2401) );
  ANDN U2880 ( .B(n2406), .A(n683), .Z(n2404) );
  XNOR U2881 ( .A(a[38]), .B(n2407), .Z(n683) );
  IV U2882 ( .A(n2405), .Z(n2407) );
  XNOR U2883 ( .A(b[38]), .B(n2405), .Z(n2406) );
  XOR U2884 ( .A(n2408), .B(n2409), .Z(n2405) );
  ANDN U2885 ( .B(n2410), .A(n734), .Z(n2408) );
  XNOR U2886 ( .A(a[37]), .B(n2411), .Z(n734) );
  IV U2887 ( .A(n2409), .Z(n2411) );
  XNOR U2888 ( .A(b[37]), .B(n2409), .Z(n2410) );
  XOR U2889 ( .A(n2412), .B(n2413), .Z(n2409) );
  ANDN U2890 ( .B(n2414), .A(n785), .Z(n2412) );
  XNOR U2891 ( .A(a[36]), .B(n2415), .Z(n785) );
  IV U2892 ( .A(n2413), .Z(n2415) );
  XNOR U2893 ( .A(b[36]), .B(n2413), .Z(n2414) );
  XOR U2894 ( .A(n2416), .B(n2417), .Z(n2413) );
  ANDN U2895 ( .B(n2418), .A(n836), .Z(n2416) );
  XNOR U2896 ( .A(a[35]), .B(n2419), .Z(n836) );
  IV U2897 ( .A(n2417), .Z(n2419) );
  XNOR U2898 ( .A(b[35]), .B(n2417), .Z(n2418) );
  XOR U2899 ( .A(n2420), .B(n2421), .Z(n2417) );
  ANDN U2900 ( .B(n2422), .A(n887), .Z(n2420) );
  XNOR U2901 ( .A(a[34]), .B(n2423), .Z(n887) );
  IV U2902 ( .A(n2421), .Z(n2423) );
  XNOR U2903 ( .A(b[34]), .B(n2421), .Z(n2422) );
  XOR U2904 ( .A(n2424), .B(n2425), .Z(n2421) );
  ANDN U2905 ( .B(n2426), .A(n938), .Z(n2424) );
  XNOR U2906 ( .A(a[33]), .B(n2427), .Z(n938) );
  IV U2907 ( .A(n2425), .Z(n2427) );
  XNOR U2908 ( .A(b[33]), .B(n2425), .Z(n2426) );
  XOR U2909 ( .A(n2428), .B(n2429), .Z(n2425) );
  ANDN U2910 ( .B(n2430), .A(n989), .Z(n2428) );
  XNOR U2911 ( .A(a[32]), .B(n2431), .Z(n989) );
  IV U2912 ( .A(n2429), .Z(n2431) );
  XNOR U2913 ( .A(b[32]), .B(n2429), .Z(n2430) );
  XOR U2914 ( .A(n2432), .B(n2433), .Z(n2429) );
  ANDN U2915 ( .B(n2434), .A(n1040), .Z(n2432) );
  XNOR U2916 ( .A(a[31]), .B(n2435), .Z(n1040) );
  IV U2917 ( .A(n2433), .Z(n2435) );
  XNOR U2918 ( .A(b[31]), .B(n2433), .Z(n2434) );
  XOR U2919 ( .A(n2436), .B(n2437), .Z(n2433) );
  ANDN U2920 ( .B(n2438), .A(n1091), .Z(n2436) );
  XNOR U2921 ( .A(a[30]), .B(n2439), .Z(n1091) );
  IV U2922 ( .A(n2437), .Z(n2439) );
  XNOR U2923 ( .A(b[30]), .B(n2437), .Z(n2438) );
  XOR U2924 ( .A(n2440), .B(n2441), .Z(n2437) );
  ANDN U2925 ( .B(n2442), .A(n1143), .Z(n2440) );
  XNOR U2926 ( .A(a[29]), .B(n2443), .Z(n1143) );
  IV U2927 ( .A(n2441), .Z(n2443) );
  XNOR U2928 ( .A(b[29]), .B(n2441), .Z(n2442) );
  XOR U2929 ( .A(n2444), .B(n2445), .Z(n2441) );
  ANDN U2930 ( .B(n2446), .A(n1194), .Z(n2444) );
  XNOR U2931 ( .A(a[28]), .B(n2447), .Z(n1194) );
  IV U2932 ( .A(n2445), .Z(n2447) );
  XNOR U2933 ( .A(b[28]), .B(n2445), .Z(n2446) );
  XOR U2934 ( .A(n2448), .B(n2449), .Z(n2445) );
  ANDN U2935 ( .B(n2450), .A(n1245), .Z(n2448) );
  XNOR U2936 ( .A(a[27]), .B(n2451), .Z(n1245) );
  IV U2937 ( .A(n2449), .Z(n2451) );
  XNOR U2938 ( .A(b[27]), .B(n2449), .Z(n2450) );
  XOR U2939 ( .A(n2452), .B(n2453), .Z(n2449) );
  ANDN U2940 ( .B(n2454), .A(n1296), .Z(n2452) );
  XNOR U2941 ( .A(a[26]), .B(n2455), .Z(n1296) );
  IV U2942 ( .A(n2453), .Z(n2455) );
  XNOR U2943 ( .A(b[26]), .B(n2453), .Z(n2454) );
  XOR U2944 ( .A(n2456), .B(n2457), .Z(n2453) );
  ANDN U2945 ( .B(n2458), .A(n1347), .Z(n2456) );
  XNOR U2946 ( .A(a[25]), .B(n2459), .Z(n1347) );
  IV U2947 ( .A(n2457), .Z(n2459) );
  XNOR U2948 ( .A(b[25]), .B(n2457), .Z(n2458) );
  XOR U2949 ( .A(n2460), .B(n2461), .Z(n2457) );
  ANDN U2950 ( .B(n2462), .A(n1398), .Z(n2460) );
  XNOR U2951 ( .A(a[24]), .B(n2463), .Z(n1398) );
  IV U2952 ( .A(n2461), .Z(n2463) );
  XNOR U2953 ( .A(b[24]), .B(n2461), .Z(n2462) );
  XOR U2954 ( .A(n2464), .B(n2465), .Z(n2461) );
  ANDN U2955 ( .B(n2466), .A(n1449), .Z(n2464) );
  XNOR U2956 ( .A(a[23]), .B(n2467), .Z(n1449) );
  IV U2957 ( .A(n2465), .Z(n2467) );
  XNOR U2958 ( .A(b[23]), .B(n2465), .Z(n2466) );
  XOR U2959 ( .A(n2468), .B(n2469), .Z(n2465) );
  ANDN U2960 ( .B(n2470), .A(n1500), .Z(n2468) );
  XNOR U2961 ( .A(a[22]), .B(n2471), .Z(n1500) );
  IV U2962 ( .A(n2469), .Z(n2471) );
  XNOR U2963 ( .A(b[22]), .B(n2469), .Z(n2470) );
  XOR U2964 ( .A(n2472), .B(n2473), .Z(n2469) );
  ANDN U2965 ( .B(n2474), .A(n1551), .Z(n2472) );
  XNOR U2966 ( .A(a[21]), .B(n2475), .Z(n1551) );
  IV U2967 ( .A(n2473), .Z(n2475) );
  XNOR U2968 ( .A(b[21]), .B(n2473), .Z(n2474) );
  XOR U2969 ( .A(n2476), .B(n2477), .Z(n2473) );
  ANDN U2970 ( .B(n2478), .A(n1602), .Z(n2476) );
  XNOR U2971 ( .A(a[20]), .B(n2479), .Z(n1602) );
  IV U2972 ( .A(n2477), .Z(n2479) );
  XNOR U2973 ( .A(b[20]), .B(n2477), .Z(n2478) );
  XOR U2974 ( .A(n2480), .B(n2481), .Z(n2477) );
  ANDN U2975 ( .B(n2482), .A(n1654), .Z(n2480) );
  XNOR U2976 ( .A(a[19]), .B(n2483), .Z(n1654) );
  IV U2977 ( .A(n2481), .Z(n2483) );
  XNOR U2978 ( .A(b[19]), .B(n2481), .Z(n2482) );
  XOR U2979 ( .A(n2484), .B(n2485), .Z(n2481) );
  ANDN U2980 ( .B(n2486), .A(n1705), .Z(n2484) );
  XNOR U2981 ( .A(a[18]), .B(n2487), .Z(n1705) );
  IV U2982 ( .A(n2485), .Z(n2487) );
  XNOR U2983 ( .A(b[18]), .B(n2485), .Z(n2486) );
  XOR U2984 ( .A(n2488), .B(n2489), .Z(n2485) );
  ANDN U2985 ( .B(n2490), .A(n1756), .Z(n2488) );
  XNOR U2986 ( .A(a[17]), .B(n2491), .Z(n1756) );
  IV U2987 ( .A(n2489), .Z(n2491) );
  XNOR U2988 ( .A(b[17]), .B(n2489), .Z(n2490) );
  XOR U2989 ( .A(n2492), .B(n2493), .Z(n2489) );
  ANDN U2990 ( .B(n2494), .A(n1807), .Z(n2492) );
  XNOR U2991 ( .A(a[16]), .B(n2495), .Z(n1807) );
  IV U2992 ( .A(n2493), .Z(n2495) );
  XNOR U2993 ( .A(b[16]), .B(n2493), .Z(n2494) );
  XOR U2994 ( .A(n2496), .B(n2497), .Z(n2493) );
  ANDN U2995 ( .B(n2498), .A(n1858), .Z(n2496) );
  XNOR U2996 ( .A(a[15]), .B(n2499), .Z(n1858) );
  IV U2997 ( .A(n2497), .Z(n2499) );
  XNOR U2998 ( .A(b[15]), .B(n2497), .Z(n2498) );
  XOR U2999 ( .A(n2500), .B(n2501), .Z(n2497) );
  ANDN U3000 ( .B(n2502), .A(n1909), .Z(n2500) );
  XNOR U3001 ( .A(a[14]), .B(n2503), .Z(n1909) );
  IV U3002 ( .A(n2501), .Z(n2503) );
  XNOR U3003 ( .A(b[14]), .B(n2501), .Z(n2502) );
  XOR U3004 ( .A(n2504), .B(n2505), .Z(n2501) );
  ANDN U3005 ( .B(n2506), .A(n1960), .Z(n2504) );
  XNOR U3006 ( .A(a[13]), .B(n2507), .Z(n1960) );
  IV U3007 ( .A(n2505), .Z(n2507) );
  XNOR U3008 ( .A(b[13]), .B(n2505), .Z(n2506) );
  XOR U3009 ( .A(n2508), .B(n2509), .Z(n2505) );
  ANDN U3010 ( .B(n2510), .A(n2011), .Z(n2508) );
  XNOR U3011 ( .A(a[12]), .B(n2511), .Z(n2011) );
  IV U3012 ( .A(n2509), .Z(n2511) );
  XNOR U3013 ( .A(b[12]), .B(n2509), .Z(n2510) );
  XOR U3014 ( .A(n2512), .B(n2513), .Z(n2509) );
  ANDN U3015 ( .B(n2514), .A(n2062), .Z(n2512) );
  XNOR U3016 ( .A(a[11]), .B(n2515), .Z(n2062) );
  IV U3017 ( .A(n2513), .Z(n2515) );
  XNOR U3018 ( .A(b[11]), .B(n2513), .Z(n2514) );
  XOR U3019 ( .A(n2516), .B(n2517), .Z(n2513) );
  ANDN U3020 ( .B(n2518), .A(n2113), .Z(n2516) );
  XNOR U3021 ( .A(a[10]), .B(n2519), .Z(n2113) );
  IV U3022 ( .A(n2517), .Z(n2519) );
  XNOR U3023 ( .A(b[10]), .B(n2517), .Z(n2518) );
  XOR U3024 ( .A(n2520), .B(n2521), .Z(n2517) );
  ANDN U3025 ( .B(n2522), .A(n6), .Z(n2520) );
  XNOR U3026 ( .A(a[9]), .B(n2523), .Z(n6) );
  IV U3027 ( .A(n2521), .Z(n2523) );
  XNOR U3028 ( .A(b[9]), .B(n2521), .Z(n2522) );
  XOR U3029 ( .A(n2524), .B(n2525), .Z(n2521) );
  ANDN U3030 ( .B(n2526), .A(n17), .Z(n2524) );
  XNOR U3031 ( .A(a[8]), .B(n2527), .Z(n17) );
  IV U3032 ( .A(n2525), .Z(n2527) );
  XNOR U3033 ( .A(b[8]), .B(n2525), .Z(n2526) );
  XOR U3034 ( .A(n2528), .B(n2529), .Z(n2525) );
  ANDN U3035 ( .B(n2530), .A(n28), .Z(n2528) );
  XNOR U3036 ( .A(a[7]), .B(n2531), .Z(n28) );
  IV U3037 ( .A(n2529), .Z(n2531) );
  XNOR U3038 ( .A(b[7]), .B(n2529), .Z(n2530) );
  XOR U3039 ( .A(n2532), .B(n2533), .Z(n2529) );
  ANDN U3040 ( .B(n2534), .A(n39), .Z(n2532) );
  XNOR U3041 ( .A(a[6]), .B(n2535), .Z(n39) );
  IV U3042 ( .A(n2533), .Z(n2535) );
  XNOR U3043 ( .A(b[6]), .B(n2533), .Z(n2534) );
  XOR U3044 ( .A(n2536), .B(n2537), .Z(n2533) );
  ANDN U3045 ( .B(n2538), .A(n50), .Z(n2536) );
  XNOR U3046 ( .A(a[5]), .B(n2539), .Z(n50) );
  IV U3047 ( .A(n2537), .Z(n2539) );
  XNOR U3048 ( .A(b[5]), .B(n2537), .Z(n2538) );
  XOR U3049 ( .A(n2540), .B(n2541), .Z(n2537) );
  ANDN U3050 ( .B(n2542), .A(n120), .Z(n2540) );
  XNOR U3051 ( .A(a[4]), .B(n2543), .Z(n120) );
  IV U3052 ( .A(n2541), .Z(n2543) );
  XNOR U3053 ( .A(b[4]), .B(n2541), .Z(n2542) );
  XOR U3054 ( .A(n2544), .B(n2545), .Z(n2541) );
  ANDN U3055 ( .B(n2546), .A(n631), .Z(n2544) );
  XNOR U3056 ( .A(a[3]), .B(n2547), .Z(n631) );
  IV U3057 ( .A(n2545), .Z(n2547) );
  XNOR U3058 ( .A(b[3]), .B(n2545), .Z(n2546) );
  XOR U3059 ( .A(n2548), .B(n2549), .Z(n2545) );
  ANDN U3060 ( .B(n2550), .A(n1142), .Z(n2548) );
  XNOR U3061 ( .A(a[2]), .B(n2551), .Z(n1142) );
  IV U3062 ( .A(n2549), .Z(n2551) );
  XNOR U3063 ( .A(b[2]), .B(n2549), .Z(n2550) );
  XOR U3064 ( .A(n2552), .B(n2553), .Z(n2549) );
  ANDN U3065 ( .B(n2554), .A(n1653), .Z(n2552) );
  XNOR U3066 ( .A(a[1]), .B(n2555), .Z(n1653) );
  IV U3067 ( .A(n2553), .Z(n2555) );
  XNOR U3068 ( .A(b[1]), .B(n2553), .Z(n2554) );
  XOR U3069 ( .A(carry_on), .B(n2556), .Z(n2553) );
  NANDN U3070 ( .A(n2557), .B(n2558), .Z(n2556) );
  XOR U3071 ( .A(carry_on), .B(b[0]), .Z(n2558) );
  XNOR U3072 ( .A(b[0]), .B(n2557), .Z(c[0]) );
  XNOR U3073 ( .A(a[0]), .B(carry_on), .Z(n2557) );
endmodule

