
module sha3_seq_CC6 ( clk, rst, in, out );
  input [575:0] in;
  output [1599:0] out;
  input clk, rst;
  wire   init, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,
         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,
         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,
         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,
         n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,
         n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,
         n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
         n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,
         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,
         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,
         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
         n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,
         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,
         n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,
         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,
         n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
         n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,
         n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,
         n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
         n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,
         n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,
         n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
         n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272,
         n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280,
         n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
         n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,
         n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,
         n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312,
         n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,
         n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,
         n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
         n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344,
         n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352,
         n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
         n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368,
         n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376,
         n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384,
         n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,
         n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400,
         n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
         n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416,
         n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,
         n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
         n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440,
         n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
         n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456,
         n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464,
         n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472,
         n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
         n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488,
         n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
         n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
         n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512,
         n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,
         n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528,
         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
         n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
         n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560,
         n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
         n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584,
         n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
         n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600,
         n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
         n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
         n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
         n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
         n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
         n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
         n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,
         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
         n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
         n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,
         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
         n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
         n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
         n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
         n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000,
         n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,
         n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016,
         n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
         n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032,
         n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040,
         n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048,
         n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
         n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064,
         n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072,
         n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080,
         n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088,
         n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096,
         n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104,
         n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112,
         n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
         n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
         n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136,
         n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144,
         n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
         n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160,
         n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
         n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,
         n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184,
         n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216,
         n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
         n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232,
         n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
         n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
         n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,
         n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,
         n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
         n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280,
         n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288,
         n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
         n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,
         n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
         n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320,
         n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328,
         n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,
         n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
         n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352,
         n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360,
         n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
         n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,
         n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
         n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
         n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
         n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
         n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
         n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424,
         n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432,
         n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
         n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
         n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,
         n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,
         n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
         n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
         n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496,
         n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
         n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
         n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
         n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
         n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536,
         n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544,
         n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,
         n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
         n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568,
         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
         n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,
         n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
         n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608,
         n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616,
         n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,
         n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
         n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
         n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,
         n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,
         n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664,
         n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,
         n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680,
         n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688,
         n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696,
         n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
         n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712,
         n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720,
         n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,
         n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736,
         n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
         n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752,
         n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,
         n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
         n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
         n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792,
         n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
         n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808,
         n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
         n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824,
         n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,
         n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840,
         n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
         n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856,
         n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864,
         n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872,
         n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880,
         n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,
         n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896,
         n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904,
         n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,
         n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920,
         n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928,
         n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936,
         n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944,
         n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952,
         n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960,
         n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968,
         n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976,
         n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984,
         n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992,
         n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000,
         n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008,
         n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016,
         n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024,
         n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032,
         n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040,
         n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048,
         n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056,
         n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064,
         n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072,
         n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080,
         n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088,
         n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096,
         n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104,
         n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112,
         n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120,
         n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128,
         n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136,
         n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144,
         n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152,
         n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160,
         n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168,
         n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176,
         n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184,
         n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192,
         n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200,
         n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208,
         n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216,
         n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224,
         n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232,
         n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240,
         n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248,
         n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256,
         n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264,
         n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272,
         n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280,
         n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288,
         n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296,
         n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304,
         n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312,
         n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320,
         n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328,
         n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336,
         n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344,
         n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352,
         n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360,
         n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368,
         n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376,
         n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384,
         n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392,
         n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400,
         n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408,
         n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416,
         n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424,
         n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432,
         n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440,
         n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448,
         n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456,
         n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464,
         n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472,
         n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480,
         n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488,
         n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496,
         n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504,
         n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512,
         n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520,
         n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528,
         n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536,
         n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544,
         n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552,
         n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560,
         n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568,
         n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576,
         n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584,
         n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592,
         n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600,
         n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608,
         n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616,
         n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624,
         n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632,
         n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640,
         n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648,
         n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656,
         n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664,
         n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672,
         n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680,
         n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688,
         n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696,
         n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704,
         n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712,
         n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720,
         n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728,
         n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736,
         n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744,
         n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752,
         n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760,
         n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768,
         n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776,
         n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784,
         n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792,
         n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800,
         n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808,
         n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816,
         n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824,
         n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832,
         n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840,
         n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848,
         n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856,
         n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864,
         n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872,
         n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880,
         n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888,
         n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896,
         n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904,
         n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912,
         n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920,
         n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928,
         n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936,
         n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944,
         n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952,
         n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960,
         n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968,
         n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976,
         n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984,
         n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992,
         n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000,
         n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008,
         n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016,
         n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024,
         n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032,
         n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040,
         n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048,
         n22049, n22050, n22051, n22052, n22053, n22054, n22055, n22056,
         n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064,
         n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072,
         n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080,
         n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088,
         n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096,
         n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104,
         n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112,
         n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120,
         n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128,
         n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136,
         n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144,
         n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152,
         n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160,
         n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168,
         n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176,
         n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184,
         n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192,
         n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200,
         n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208,
         n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216,
         n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224,
         n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232,
         n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240,
         n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248,
         n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256,
         n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264,
         n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272,
         n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280,
         n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288,
         n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296,
         n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304,
         n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312,
         n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320,
         n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328,
         n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336,
         n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344,
         n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352,
         n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360,
         n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368,
         n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376,
         n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384,
         n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392,
         n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400,
         n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408,
         n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416,
         n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424,
         n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432,
         n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440,
         n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448,
         n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456,
         n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464,
         n22465, n22466, n22467, n22468, n22469, n22470, n22471, n22472,
         n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480,
         n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488,
         n22489, n22490, n22491, n22492, n22493, n22494, n22495, n22496,
         n22497, n22498, n22499, n22500, n22501, n22502, n22503, n22504,
         n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512,
         n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520,
         n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528,
         n22529, n22530, n22531, n22532, n22533, n22534, n22535, n22536,
         n22537, n22538, n22539, n22540, n22541, n22542, n22543, n22544,
         n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552,
         n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560,
         n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568,
         n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576,
         n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584,
         n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592,
         n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600,
         n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608,
         n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616,
         n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624,
         n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632,
         n22633, n22634, n22635, n22636, n22637, n22638, n22639, n22640,
         n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648,
         n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656,
         n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664,
         n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672,
         n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680,
         n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688,
         n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696,
         n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704,
         n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712,
         n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720,
         n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728,
         n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736,
         n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744,
         n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752,
         n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760,
         n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768,
         n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776,
         n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784,
         n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792,
         n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800,
         n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808,
         n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816,
         n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824,
         n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832,
         n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840,
         n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848,
         n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856,
         n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864,
         n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872,
         n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880,
         n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888,
         n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22896,
         n22897, n22898, n22899, n22900, n22901, n22902, n22903, n22904,
         n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912,
         n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920,
         n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928,
         n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936,
         n22937, n22938, n22939, n22940, n22941, n22942, n22943, n22944,
         n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952,
         n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960,
         n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968,
         n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976,
         n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984,
         n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992,
         n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000,
         n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008,
         n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016,
         n23017, n23018, n23019, n23020, n23021, n23022, n23023, n23024,
         n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032,
         n23033, n23034, n23035, n23036, n23037, n23038, n23039, n23040,
         n23041, n23042, n23043, n23044, n23045, n23046, n23047, n23048,
         n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056,
         n23057, n23058, n23059, n23060, n23061, n23062, n23063, n23064,
         n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072,
         n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080,
         n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088,
         n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096,
         n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104,
         n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112,
         n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23120,
         n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128,
         n23129, n23130, n23131, n23132, n23133, n23134, n23135, n23136,
         n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144,
         n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152,
         n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160,
         n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168,
         n23169, n23170, n23171, n23172, n23173, n23174, n23175, n23176,
         n23177, n23178, n23179, n23180, n23181, n23182, n23183, n23184,
         n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192,
         n23193, n23194, n23195, n23196, n23197, n23198, n23199, n23200,
         n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208,
         n23209, n23210, n23211, n23212, n23213, n23214, n23215, n23216,
         n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224,
         n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232,
         n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240,
         n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248,
         n23249, n23250, n23251, n23252, n23253, n23254, n23255, n23256,
         n23257, n23258, n23259, n23260, n23261, n23262, n23263, n23264,
         n23265, n23266, n23267, n23268, n23269, n23270, n23271, n23272,
         n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280,
         n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288,
         n23289, n23290, n23291, n23292, n23293, n23294, n23295, n23296,
         n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304,
         n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23312,
         n23313, n23314, n23315, n23316, n23317, n23318, n23319, n23320,
         n23321, n23322, n23323, n23324, n23325, n23326, n23327, n23328,
         n23329, n23330, n23331, n23332, n23333, n23334, n23335, n23336,
         n23337, n23338, n23339, n23340, n23341, n23342, n23343, n23344,
         n23345, n23346, n23347, n23348, n23349, n23350, n23351, n23352,
         n23353, n23354, n23355, n23356, n23357, n23358, n23359, n23360,
         n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368,
         n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376,
         n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384,
         n23385, n23386, n23387, n23388, n23389, n23390, n23391, n23392,
         n23393, n23394, n23395, n23396, n23397, n23398, n23399, n23400,
         n23401, n23402, n23403, n23404, n23405, n23406, n23407, n23408,
         n23409, n23410, n23411, n23412, n23413, n23414, n23415, n23416,
         n23417, n23418, n23419, n23420, n23421, n23422, n23423, n23424,
         n23425, n23426, n23427, n23428, n23429, n23430, n23431, n23432,
         n23433, n23434, n23435, n23436, n23437, n23438, n23439, n23440,
         n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448,
         n23449, n23450, n23451, n23452, n23453, n23454, n23455, n23456,
         n23457, n23458, n23459, n23460, n23461, n23462, n23463, n23464,
         n23465, n23466, n23467, n23468, n23469, n23470, n23471, n23472,
         n23473, n23474, n23475, n23476, n23477, n23478, n23479, n23480,
         n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488,
         n23489, n23490, n23491, n23492, n23493, n23494, n23495, n23496,
         n23497, n23498, n23499, n23500, n23501, n23502, n23503, n23504,
         n23505, n23506, n23507, n23508, n23509, n23510, n23511, n23512,
         n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520,
         n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528,
         n23529, n23530, n23531, n23532, n23533, n23534, n23535, n23536,
         n23537, n23538, n23539, n23540, n23541, n23542, n23543, n23544,
         n23545, n23546, n23547, n23548, n23549, n23550, n23551, n23552,
         n23553, n23554, n23555, n23556, n23557, n23558, n23559, n23560,
         n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568,
         n23569, n23570, n23571, n23572, n23573, n23574, n23575, n23576,
         n23577, n23578, n23579, n23580, n23581, n23582, n23583, n23584,
         n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592,
         n23593, n23594, n23595, n23596, n23597, n23598, n23599, n23600,
         n23601, n23602, n23603, n23604, n23605, n23606, n23607, n23608,
         n23609, n23610, n23611, n23612, n23613, n23614, n23615, n23616,
         n23617, n23618, n23619, n23620, n23621, n23622, n23623, n23624,
         n23625, n23626, n23627, n23628, n23629, n23630, n23631, n23632,
         n23633, n23634, n23635, n23636, n23637, n23638, n23639, n23640,
         n23641, n23642, n23643, n23644, n23645, n23646, n23647, n23648,
         n23649, n23650, n23651, n23652, n23653, n23654, n23655, n23656,
         n23657, n23658, n23659, n23660, n23661, n23662, n23663, n23664,
         n23665, n23666, n23667, n23668, n23669, n23670, n23671, n23672,
         n23673, n23674, n23675, n23676, n23677, n23678, n23679, n23680,
         n23681, n23682, n23683, n23684, n23685, n23686, n23687, n23688,
         n23689, n23690, n23691, n23692, n23693, n23694, n23695, n23696,
         n23697, n23698, n23699, n23700, n23701, n23702, n23703, n23704,
         n23705, n23706, n23707, n23708, n23709, n23710, n23711, n23712,
         n23713, n23714, n23715, n23716, n23717, n23718, n23719, n23720,
         n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728,
         n23729, n23730, n23731, n23732, n23733, n23734, n23735, n23736,
         n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744,
         n23745, n23746, n23747, n23748, n23749, n23750, n23751, n23752,
         n23753, n23754, n23755, n23756, n23757, n23758, n23759, n23760,
         n23761, n23762, n23763, n23764, n23765, n23766, n23767, n23768,
         n23769, n23770, n23771, n23772, n23773, n23774, n23775, n23776,
         n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784,
         n23785, n23786, n23787, n23788, n23789, n23790, n23791, n23792,
         n23793, n23794, n23795, n23796, n23797, n23798, n23799, n23800,
         n23801, n23802, n23803, n23804, n23805, n23806, n23807, n23808,
         n23809, n23810, n23811, n23812, n23813, n23814, n23815, n23816,
         n23817, n23818, n23819, n23820, n23821, n23822, n23823, n23824,
         n23825, n23826, n23827, n23828, n23829, n23830, n23831, n23832,
         n23833, n23834, n23835, n23836, n23837, n23838, n23839, n23840,
         n23841, n23842, n23843, n23844, n23845, n23846, n23847, n23848,
         n23849, n23850, n23851, n23852, n23853, n23854, n23855, n23856,
         n23857, n23858, n23859, n23860, n23861, n23862, n23863, n23864,
         n23865, n23866, n23867, n23868, n23869, n23870, n23871, n23872,
         n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23880,
         n23881, n23882, n23883, n23884, n23885, n23886, n23887, n23888,
         n23889, n23890, n23891, n23892, n23893, n23894, n23895, n23896,
         n23897, n23898, n23899, n23900, n23901, n23902, n23903, n23904,
         n23905, n23906, n23907, n23908, n23909, n23910, n23911, n23912,
         n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920,
         n23921, n23922, n23923, n23924, n23925, n23926, n23927, n23928,
         n23929, n23930, n23931, n23932, n23933, n23934, n23935, n23936,
         n23937, n23938, n23939, n23940, n23941, n23942, n23943, n23944,
         n23945, n23946, n23947, n23948, n23949, n23950, n23951, n23952,
         n23953, n23954, n23955, n23956, n23957, n23958, n23959, n23960,
         n23961, n23962, n23963, n23964, n23965, n23966, n23967, n23968,
         n23969, n23970, n23971, n23972, n23973, n23974, n23975, n23976,
         n23977, n23978, n23979, n23980, n23981, n23982, n23983, n23984,
         n23985, n23986, n23987, n23988, n23989, n23990, n23991, n23992,
         n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000,
         n24001, n24002, n24003, n24004, n24005, n24006, n24007, n24008,
         n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016,
         n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024,
         n24025, n24026, n24027, n24028, n24029, n24030, n24031, n24032,
         n24033, n24034, n24035, n24036, n24037, n24038, n24039, n24040,
         n24041, n24042, n24043, n24044, n24045, n24046, n24047, n24048,
         n24049, n24050, n24051, n24052, n24053, n24054, n24055, n24056,
         n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064,
         n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072,
         n24073, n24074, n24075, n24076, n24077, n24078, n24079, n24080,
         n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088,
         n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096,
         n24097, n24098, n24099, n24100, n24101, n24102, n24103, n24104,
         n24105, n24106, n24107, n24108, n24109, n24110, n24111, n24112,
         n24113, n24114, n24115, n24116, n24117, n24118, n24119, n24120,
         n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128,
         n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136,
         n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144,
         n24145, n24146, n24147, n24148, n24149, n24150, n24151, n24152,
         n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160,
         n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168,
         n24169, n24170, n24171, n24172, n24173, n24174, n24175, n24176,
         n24177, n24178, n24179, n24180, n24181, n24182, n24183, n24184,
         n24185, n24186, n24187, n24188, n24189, n24190, n24191, n24192,
         n24193, n24194, n24195, n24196, n24197, n24198, n24199, n24200,
         n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208,
         n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24216,
         n24217, n24218, n24219, n24220, n24221, n24222, n24223, n24224,
         n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232,
         n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240,
         n24241, n24242, n24243, n24244, n24245, n24246, n24247, n24248,
         n24249, n24250, n24251, n24252, n24253, n24254, n24255, n24256,
         n24257, n24258, n24259, n24260, n24261, n24262, n24263, n24264,
         n24265, n24266, n24267, n24268, n24269, n24270, n24271, n24272,
         n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280,
         n24281, n24282, n24283, n24284, n24285, n24286, n24287, n24288,
         n24289, n24290, n24291, n24292, n24293, n24294, n24295, n24296,
         n24297, n24298, n24299, n24300, n24301, n24302, n24303, n24304,
         n24305, n24306, n24307, n24308, n24309, n24310, n24311, n24312,
         n24313, n24314, n24315, n24316, n24317, n24318, n24319, n24320,
         n24321, n24322, n24323, n24324, n24325, n24326, n24327, n24328,
         n24329, n24330, n24331, n24332, n24333, n24334, n24335, n24336,
         n24337, n24338, n24339, n24340, n24341, n24342, n24343, n24344,
         n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352,
         n24353, n24354, n24355, n24356, n24357, n24358, n24359, n24360,
         n24361, n24362, n24363, n24364, n24365, n24366, n24367, n24368,
         n24369, n24370, n24371, n24372, n24373, n24374, n24375, n24376,
         n24377, n24378, n24379, n24380, n24381, n24382, n24383, n24384,
         n24385, n24386, n24387, n24388, n24389, n24390, n24391, n24392,
         n24393, n24394, n24395, n24396, n24397, n24398, n24399, n24400,
         n24401, n24402, n24403, n24404, n24405, n24406, n24407, n24408,
         n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416,
         n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424,
         n24425, n24426, n24427, n24428, n24429, n24430, n24431, n24432,
         n24433, n24434, n24435, n24436, n24437, n24438, n24439, n24440,
         n24441, n24442, n24443, n24444, n24445, n24446, n24447, n24448,
         n24449, n24450, n24451, n24452, n24453, n24454, n24455, n24456,
         n24457, n24458, n24459, n24460, n24461, n24462, n24463, n24464,
         n24465, n24466, n24467, n24468, n24469, n24470, n24471, n24472,
         n24473, n24474, n24475, n24476, n24477, n24478, n24479, n24480,
         n24481, n24482, n24483, n24484, n24485, n24486, n24487, n24488,
         n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496,
         n24497, n24498, n24499, n24500, n24501, n24502, n24503, n24504,
         n24505, n24506, n24507, n24508, n24509, n24510, n24511, n24512,
         n24513, n24514, n24515, n24516, n24517, n24518, n24519, n24520,
         n24521, n24522, n24523, n24524, n24525, n24526, n24527, n24528,
         n24529, n24530, n24531, n24532, n24533, n24534, n24535, n24536,
         n24537, n24538, n24539, n24540, n24541, n24542, n24543, n24544,
         n24545, n24546, n24547, n24548, n24549, n24550, n24551, n24552,
         n24553, n24554, n24555, n24556, n24557, n24558, n24559, n24560,
         n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568,
         n24569, n24570, n24571, n24572, n24573, n24574, n24575, n24576,
         n24577, n24578, n24579, n24580, n24581, n24582, n24583, n24584,
         n24585, n24586, n24587, n24588, n24589, n24590, n24591, n24592,
         n24593, n24594, n24595, n24596, n24597, n24598, n24599, n24600,
         n24601, n24602, n24603, n24604, n24605, n24606, n24607, n24608,
         n24609, n24610, n24611, n24612, n24613, n24614, n24615, n24616,
         n24617, n24618, n24619, n24620, n24621, n24622, n24623, n24624,
         n24625, n24626, n24627, n24628, n24629, n24630, n24631, n24632,
         n24633, n24634, n24635, n24636, n24637, n24638, n24639, n24640,
         n24641, n24642, n24643, n24644, n24645, n24646, n24647, n24648,
         n24649, n24650, n24651, n24652, n24653, n24654, n24655, n24656,
         n24657, n24658, n24659, n24660, n24661, n24662, n24663, n24664,
         n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672,
         n24673, n24674, n24675, n24676, n24677, n24678, n24679, n24680,
         n24681, n24682, n24683, n24684, n24685, n24686, n24687, n24688,
         n24689, n24690, n24691, n24692, n24693, n24694, n24695, n24696,
         n24697, n24698, n24699, n24700, n24701, n24702, n24703, n24704,
         n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712,
         n24713, n24714, n24715, n24716, n24717, n24718, n24719, n24720,
         n24721, n24722, n24723, n24724, n24725, n24726, n24727, n24728,
         n24729, n24730, n24731, n24732, n24733, n24734, n24735, n24736,
         n24737, n24738, n24739, n24740, n24741, n24742, n24743, n24744,
         n24745, n24746, n24747, n24748, n24749, n24750, n24751, n24752,
         n24753, n24754, n24755, n24756, n24757, n24758, n24759, n24760,
         n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768,
         n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776,
         n24777, n24778, n24779, n24780, n24781, n24782, n24783, n24784,
         n24785, n24786, n24787, n24788, n24789, n24790, n24791, n24792,
         n24793, n24794, n24795, n24796, n24797, n24798, n24799, n24800,
         n24801, n24802, n24803, n24804, n24805, n24806, n24807, n24808,
         n24809, n24810, n24811, n24812, n24813, n24814, n24815, n24816,
         n24817, n24818, n24819, n24820, n24821, n24822, n24823, n24824,
         n24825, n24826, n24827, n24828, n24829, n24830, n24831, n24832,
         n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24840,
         n24841, n24842, n24843, n24844, n24845, n24846, n24847, n24848,
         n24849, n24850, n24851, n24852, n24853, n24854, n24855, n24856,
         n24857, n24858, n24859, n24860, n24861, n24862, n24863, n24864,
         n24865, n24866, n24867, n24868, n24869, n24870, n24871, n24872,
         n24873, n24874, n24875, n24876, n24877, n24878, n24879, n24880,
         n24881, n24882, n24883, n24884, n24885, n24886, n24887, n24888,
         n24889, n24890, n24891, n24892, n24893, n24894, n24895, n24896,
         n24897, n24898, n24899, n24900, n24901, n24902, n24903, n24904,
         n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912,
         n24913, n24914, n24915, n24916, n24917, n24918, n24919, n24920,
         n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928,
         n24929, n24930, n24931, n24932, n24933, n24934, n24935, n24936,
         n24937, n24938, n24939, n24940, n24941, n24942, n24943, n24944,
         n24945, n24946, n24947, n24948, n24949, n24950, n24951, n24952,
         n24953, n24954, n24955, n24956, n24957, n24958, n24959, n24960,
         n24961, n24962, n24963, n24964, n24965, n24966, n24967, n24968,
         n24969, n24970, n24971, n24972, n24973, n24974, n24975, n24976,
         n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984,
         n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992,
         n24993, n24994, n24995, n24996, n24997, n24998, n24999, n25000,
         n25001, n25002, n25003, n25004, n25005, n25006, n25007, n25008,
         n25009, n25010, n25011, n25012, n25013, n25014, n25015, n25016,
         n25017, n25018, n25019, n25020, n25021, n25022, n25023, n25024,
         n25025, n25026, n25027, n25028, n25029, n25030, n25031, n25032,
         n25033, n25034, n25035, n25036, n25037, n25038, n25039, n25040,
         n25041, n25042, n25043, n25044, n25045, n25046, n25047, n25048,
         n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056,
         n25057, n25058, n25059, n25060, n25061, n25062, n25063, n25064,
         n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072,
         n25073, n25074, n25075, n25076, n25077, n25078, n25079, n25080,
         n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088,
         n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096,
         n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104,
         n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112,
         n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120,
         n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128,
         n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136,
         n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144,
         n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152,
         n25153, n25154, n25155, n25156, n25157, n25158, n25159, n25160,
         n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168,
         n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176,
         n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184,
         n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192,
         n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200,
         n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208,
         n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216,
         n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224,
         n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232,
         n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240,
         n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248,
         n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256,
         n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264,
         n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272,
         n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280,
         n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288,
         n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296,
         n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304,
         n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312,
         n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320,
         n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25328,
         n25329, n25330, n25331, n25332, n25333, n25334, n25335, n25336,
         n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344,
         n25345, n25346, n25347, n25348, n25349, n25350, n25351, n25352,
         n25353, n25354, n25355, n25356, n25357, n25358, n25359, n25360,
         n25361, n25362, n25363, n25364, n25365, n25366, n25367, n25368,
         n25369, n25370, n25371, n25372, n25373, n25374, n25375, n25376,
         n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384,
         n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392,
         n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400,
         n25401, n25402, n25403, n25404, n25405, n25406, n25407, n25408,
         n25409, n25410, n25411, n25412, n25413, n25414, n25415, n25416,
         n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424,
         n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432,
         n25433, n25434, n25435, n25436, n25437, n25438, n25439, n25440,
         n25441, n25442, n25443, n25444, n25445, n25446, n25447, n25448,
         n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456,
         n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464,
         n25465, n25466, n25467, n25468, n25469, n25470, n25471, n25472,
         n25473, n25474, n25475, n25476, n25477, n25478, n25479, n25480,
         n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488,
         n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496,
         n25497, n25498, n25499, n25500, n25501, n25502, n25503, n25504,
         n25505, n25506, n25507, n25508, n25509, n25510, n25511, n25512,
         n25513, n25514, n25515, n25516, n25517, n25518, n25519, n25520,
         n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528,
         n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536,
         n25537, n25538, n25539, n25540, n25541, n25542, n25543, n25544,
         n25545, n25546, n25547, n25548, n25549, n25550, n25551, n25552,
         n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560,
         n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568,
         n25569, n25570, n25571, n25572, n25573, n25574, n25575, n25576,
         n25577, n25578, n25579, n25580, n25581, n25582, n25583, n25584,
         n25585, n25586, n25587, n25588, n25589, n25590, n25591, n25592,
         n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600,
         n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608,
         n25609, n25610, n25611, n25612, n25613, n25614, n25615, n25616,
         n25617, n25618, n25619, n25620, n25621, n25622, n25623, n25624,
         n25625, n25626, n25627, n25628, n25629, n25630, n25631, n25632,
         n25633, n25634, n25635, n25636, n25637, n25638, n25639, n25640,
         n25641, n25642, n25643, n25644, n25645, n25646, n25647, n25648,
         n25649, n25650, n25651, n25652, n25653, n25654, n25655, n25656,
         n25657, n25658, n25659, n25660, n25661, n25662, n25663, n25664,
         n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672,
         n25673, n25674, n25675, n25676, n25677, n25678, n25679, n25680,
         n25681, n25682, n25683, n25684, n25685, n25686, n25687, n25688,
         n25689, n25690, n25691, n25692, n25693, n25694, n25695, n25696,
         n25697, n25698, n25699, n25700, n25701, n25702, n25703, n25704,
         n25705, n25706, n25707, n25708, n25709, n25710, n25711, n25712,
         n25713, n25714, n25715, n25716, n25717, n25718, n25719, n25720,
         n25721, n25722, n25723, n25724, n25725, n25726, n25727, n25728,
         n25729, n25730, n25731, n25732, n25733, n25734, n25735, n25736,
         n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744,
         n25745, n25746, n25747, n25748, n25749, n25750, n25751, n25752,
         n25753, n25754, n25755, n25756, n25757, n25758, n25759, n25760,
         n25761, n25762, n25763, n25764, n25765, n25766, n25767, n25768,
         n25769, n25770, n25771, n25772, n25773, n25774, n25775, n25776,
         n25777, n25778, n25779, n25780, n25781, n25782, n25783, n25784,
         n25785, n25786, n25787, n25788, n25789, n25790, n25791, n25792,
         n25793, n25794, n25795, n25796, n25797, n25798, n25799, n25800,
         n25801, n25802, n25803, n25804, n25805, n25806, n25807, n25808,
         n25809, n25810, n25811, n25812, n25813, n25814, n25815, n25816,
         n25817, n25818, n25819, n25820, n25821, n25822, n25823, n25824,
         n25825, n25826, n25827, n25828, n25829, n25830, n25831, n25832,
         n25833, n25834, n25835, n25836, n25837, n25838, n25839, n25840,
         n25841, n25842, n25843, n25844, n25845, n25846, n25847, n25848,
         n25849, n25850, n25851, n25852, n25853, n25854, n25855, n25856,
         n25857, n25858, n25859, n25860, n25861, n25862, n25863, n25864,
         n25865, n25866, n25867, n25868, n25869, n25870, n25871, n25872,
         n25873, n25874, n25875, n25876, n25877, n25878, n25879, n25880,
         n25881, n25882, n25883, n25884, n25885, n25886, n25887, n25888,
         n25889, n25890, n25891, n25892, n25893, n25894, n25895, n25896,
         n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904,
         n25905, n25906, n25907, n25908, n25909, n25910, n25911, n25912,
         n25913, n25914, n25915, n25916, n25917, n25918, n25919, n25920,
         n25921, n25922, n25923, n25924, n25925, n25926, n25927, n25928,
         n25929, n25930, n25931, n25932, n25933, n25934, n25935, n25936,
         n25937, n25938, n25939, n25940, n25941, n25942, n25943, n25944,
         n25945, n25946, n25947, n25948, n25949, n25950, n25951, n25952,
         n25953, n25954, n25955, n25956, n25957, n25958, n25959, n25960,
         n25961, n25962, n25963, n25964, n25965, n25966, n25967, n25968,
         n25969, n25970, n25971, n25972, n25973, n25974, n25975, n25976,
         n25977, n25978, n25979, n25980, n25981, n25982, n25983, n25984,
         n25985, n25986, n25987, n25988, n25989, n25990, n25991, n25992,
         n25993, n25994, n25995, n25996, n25997, n25998, n25999, n26000,
         n26001, n26002, n26003, n26004, n26005, n26006, n26007, n26008,
         n26009, n26010, n26011, n26012, n26013, n26014, n26015, n26016,
         n26017, n26018, n26019, n26020, n26021, n26022, n26023, n26024,
         n26025, n26026, n26027, n26028, n26029, n26030, n26031, n26032,
         n26033, n26034, n26035, n26036, n26037, n26038, n26039, n26040,
         n26041, n26042, n26043, n26044, n26045, n26046, n26047, n26048,
         n26049, n26050, n26051, n26052, n26053, n26054, n26055, n26056,
         n26057, n26058, n26059, n26060, n26061, n26062, n26063, n26064,
         n26065, n26066, n26067, n26068, n26069, n26070, n26071, n26072,
         n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080,
         n26081, n26082, n26083, n26084, n26085, n26086, n26087, n26088,
         n26089, n26090, n26091, n26092, n26093, n26094, n26095, n26096,
         n26097, n26098, n26099, n26100, n26101, n26102, n26103, n26104,
         n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112,
         n26113, n26114, n26115, n26116, n26117, n26118, n26119, n26120,
         n26121, n26122, n26123, n26124, n26125, n26126, n26127, n26128,
         n26129, n26130, n26131, n26132, n26133, n26134, n26135, n26136,
         n26137, n26138, n26139, n26140, n26141, n26142, n26143, n26144,
         n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152,
         n26153, n26154, n26155, n26156, n26157, n26158, n26159, n26160,
         n26161, n26162, n26163, n26164, n26165, n26166, n26167, n26168,
         n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176,
         n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184,
         n26185, n26186, n26187, n26188, n26189, n26190, n26191, n26192,
         n26193, n26194, n26195, n26196, n26197, n26198, n26199, n26200,
         n26201, n26202, n26203, n26204, n26205, n26206, n26207, n26208,
         n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216,
         n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224,
         n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232,
         n26233, n26234, n26235, n26236, n26237, n26238, n26239, n26240,
         n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248,
         n26249, n26250, n26251, n26252, n26253, n26254, n26255, n26256,
         n26257, n26258, n26259, n26260, n26261, n26262, n26263, n26264,
         n26265, n26266, n26267, n26268, n26269, n26270, n26271, n26272,
         n26273, n26274, n26275, n26276, n26277, n26278, n26279, n26280,
         n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288,
         n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296,
         n26297, n26298, n26299, n26300, n26301, n26302, n26303, n26304,
         n26305, n26306, n26307, n26308, n26309, n26310, n26311, n26312,
         n26313, n26314, n26315, n26316, n26317, n26318, n26319, n26320,
         n26321, n26322, n26323, n26324, n26325, n26326, n26327, n26328,
         n26329, n26330, n26331, n26332, n26333, n26334, n26335, n26336,
         n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344,
         n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352,
         n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360,
         n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368,
         n26369, n26370, n26371, n26372, n26373, n26374, n26375, n26376,
         n26377, n26378, n26379, n26380, n26381, n26382, n26383, n26384,
         n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392,
         n26393, n26394, n26395, n26396, n26397, n26398, n26399, n26400,
         n26401, n26402, n26403, n26404, n26405, n26406, n26407, n26408,
         n26409, n26410, n26411, n26412, n26413, n26414, n26415, n26416,
         n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424,
         n26425, n26426, n26427, n26428, n26429, n26430, n26431, n26432,
         n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440,
         n26441, n26442, n26443, n26444, n26445, n26446, n26447, n26448,
         n26449, n26450, n26451, n26452, n26453, n26454, n26455, n26456,
         n26457, n26458, n26459, n26460, n26461, n26462, n26463, n26464,
         n26465, n26466, n26467, n26468, n26469, n26470, n26471, n26472,
         n26473, n26474, n26475, n26476, n26477, n26478, n26479, n26480,
         n26481, n26482, n26483, n26484, n26485, n26486, n26487, n26488,
         n26489, n26490, n26491, n26492, n26493, n26494, n26495, n26496,
         n26497, n26498, n26499, n26500, n26501, n26502, n26503, n26504,
         n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26512,
         n26513, n26514, n26515, n26516, n26517, n26518;
  wire   [5:0] rc_i;
  wire   [1599:0] round_reg;

  DFF init_reg ( .D(1'b1), .CLK(clk), .RST(rst), .I(1'b0), .Q(init) );
  DFF \rc_i_reg[0]  ( .D(n1032), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[0])
         );
  DFF \rc_i_reg[1]  ( .D(rc_i[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[1])
         );
  DFF \rc_i_reg[2]  ( .D(rc_i[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[2])
         );
  DFF \rc_i_reg[3]  ( .D(rc_i[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[3])
         );
  DFF \rc_i_reg[4]  ( .D(rc_i[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[4])
         );
  DFF \rc_i_reg[5]  ( .D(rc_i[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[5])
         );
  DFF \round_reg_reg[0]  ( .D(out[0]), .CLK(clk), .RST(rst), .I(in[0]), .Q(
        round_reg[0]) );
  DFF \round_reg_reg[1]  ( .D(out[1]), .CLK(clk), .RST(rst), .I(in[1]), .Q(
        round_reg[1]) );
  DFF \round_reg_reg[2]  ( .D(out[2]), .CLK(clk), .RST(rst), .I(in[2]), .Q(
        round_reg[2]) );
  DFF \round_reg_reg[3]  ( .D(out[3]), .CLK(clk), .RST(rst), .I(in[3]), .Q(
        round_reg[3]) );
  DFF \round_reg_reg[4]  ( .D(out[4]), .CLK(clk), .RST(rst), .I(in[4]), .Q(
        round_reg[4]) );
  DFF \round_reg_reg[5]  ( .D(out[5]), .CLK(clk), .RST(rst), .I(in[5]), .Q(
        round_reg[5]) );
  DFF \round_reg_reg[6]  ( .D(out[6]), .CLK(clk), .RST(rst), .I(in[6]), .Q(
        round_reg[6]) );
  DFF \round_reg_reg[7]  ( .D(out[7]), .CLK(clk), .RST(rst), .I(in[7]), .Q(
        round_reg[7]) );
  DFF \round_reg_reg[8]  ( .D(out[8]), .CLK(clk), .RST(rst), .I(in[8]), .Q(
        round_reg[8]) );
  DFF \round_reg_reg[9]  ( .D(out[9]), .CLK(clk), .RST(rst), .I(in[9]), .Q(
        round_reg[9]) );
  DFF \round_reg_reg[10]  ( .D(out[10]), .CLK(clk), .RST(rst), .I(in[10]), .Q(
        round_reg[10]) );
  DFF \round_reg_reg[11]  ( .D(out[11]), .CLK(clk), .RST(rst), .I(in[11]), .Q(
        round_reg[11]) );
  DFF \round_reg_reg[12]  ( .D(out[12]), .CLK(clk), .RST(rst), .I(in[12]), .Q(
        round_reg[12]) );
  DFF \round_reg_reg[13]  ( .D(out[13]), .CLK(clk), .RST(rst), .I(in[13]), .Q(
        round_reg[13]) );
  DFF \round_reg_reg[14]  ( .D(out[14]), .CLK(clk), .RST(rst), .I(in[14]), .Q(
        round_reg[14]) );
  DFF \round_reg_reg[15]  ( .D(out[15]), .CLK(clk), .RST(rst), .I(in[15]), .Q(
        round_reg[15]) );
  DFF \round_reg_reg[16]  ( .D(out[16]), .CLK(clk), .RST(rst), .I(in[16]), .Q(
        round_reg[16]) );
  DFF \round_reg_reg[17]  ( .D(out[17]), .CLK(clk), .RST(rst), .I(in[17]), .Q(
        round_reg[17]) );
  DFF \round_reg_reg[18]  ( .D(out[18]), .CLK(clk), .RST(rst), .I(in[18]), .Q(
        round_reg[18]) );
  DFF \round_reg_reg[19]  ( .D(out[19]), .CLK(clk), .RST(rst), .I(in[19]), .Q(
        round_reg[19]) );
  DFF \round_reg_reg[20]  ( .D(out[20]), .CLK(clk), .RST(rst), .I(in[20]), .Q(
        round_reg[20]) );
  DFF \round_reg_reg[21]  ( .D(out[21]), .CLK(clk), .RST(rst), .I(in[21]), .Q(
        round_reg[21]) );
  DFF \round_reg_reg[22]  ( .D(out[22]), .CLK(clk), .RST(rst), .I(in[22]), .Q(
        round_reg[22]) );
  DFF \round_reg_reg[23]  ( .D(out[23]), .CLK(clk), .RST(rst), .I(in[23]), .Q(
        round_reg[23]) );
  DFF \round_reg_reg[24]  ( .D(out[24]), .CLK(clk), .RST(rst), .I(in[24]), .Q(
        round_reg[24]) );
  DFF \round_reg_reg[25]  ( .D(out[25]), .CLK(clk), .RST(rst), .I(in[25]), .Q(
        round_reg[25]) );
  DFF \round_reg_reg[26]  ( .D(out[26]), .CLK(clk), .RST(rst), .I(in[26]), .Q(
        round_reg[26]) );
  DFF \round_reg_reg[27]  ( .D(out[27]), .CLK(clk), .RST(rst), .I(in[27]), .Q(
        round_reg[27]) );
  DFF \round_reg_reg[28]  ( .D(out[28]), .CLK(clk), .RST(rst), .I(in[28]), .Q(
        round_reg[28]) );
  DFF \round_reg_reg[29]  ( .D(out[29]), .CLK(clk), .RST(rst), .I(in[29]), .Q(
        round_reg[29]) );
  DFF \round_reg_reg[30]  ( .D(out[30]), .CLK(clk), .RST(rst), .I(in[30]), .Q(
        round_reg[30]) );
  DFF \round_reg_reg[31]  ( .D(out[31]), .CLK(clk), .RST(rst), .I(in[31]), .Q(
        round_reg[31]) );
  DFF \round_reg_reg[32]  ( .D(out[32]), .CLK(clk), .RST(rst), .I(in[32]), .Q(
        round_reg[32]) );
  DFF \round_reg_reg[33]  ( .D(out[33]), .CLK(clk), .RST(rst), .I(in[33]), .Q(
        round_reg[33]) );
  DFF \round_reg_reg[34]  ( .D(out[34]), .CLK(clk), .RST(rst), .I(in[34]), .Q(
        round_reg[34]) );
  DFF \round_reg_reg[35]  ( .D(out[35]), .CLK(clk), .RST(rst), .I(in[35]), .Q(
        round_reg[35]) );
  DFF \round_reg_reg[36]  ( .D(out[36]), .CLK(clk), .RST(rst), .I(in[36]), .Q(
        round_reg[36]) );
  DFF \round_reg_reg[37]  ( .D(out[37]), .CLK(clk), .RST(rst), .I(in[37]), .Q(
        round_reg[37]) );
  DFF \round_reg_reg[38]  ( .D(out[38]), .CLK(clk), .RST(rst), .I(in[38]), .Q(
        round_reg[38]) );
  DFF \round_reg_reg[39]  ( .D(out[39]), .CLK(clk), .RST(rst), .I(in[39]), .Q(
        round_reg[39]) );
  DFF \round_reg_reg[40]  ( .D(out[40]), .CLK(clk), .RST(rst), .I(in[40]), .Q(
        round_reg[40]) );
  DFF \round_reg_reg[41]  ( .D(out[41]), .CLK(clk), .RST(rst), .I(in[41]), .Q(
        round_reg[41]) );
  DFF \round_reg_reg[42]  ( .D(out[42]), .CLK(clk), .RST(rst), .I(in[42]), .Q(
        round_reg[42]) );
  DFF \round_reg_reg[43]  ( .D(out[43]), .CLK(clk), .RST(rst), .I(in[43]), .Q(
        round_reg[43]) );
  DFF \round_reg_reg[44]  ( .D(out[44]), .CLK(clk), .RST(rst), .I(in[44]), .Q(
        round_reg[44]) );
  DFF \round_reg_reg[45]  ( .D(out[45]), .CLK(clk), .RST(rst), .I(in[45]), .Q(
        round_reg[45]) );
  DFF \round_reg_reg[46]  ( .D(out[46]), .CLK(clk), .RST(rst), .I(in[46]), .Q(
        round_reg[46]) );
  DFF \round_reg_reg[47]  ( .D(out[47]), .CLK(clk), .RST(rst), .I(in[47]), .Q(
        round_reg[47]) );
  DFF \round_reg_reg[48]  ( .D(out[48]), .CLK(clk), .RST(rst), .I(in[48]), .Q(
        round_reg[48]) );
  DFF \round_reg_reg[49]  ( .D(out[49]), .CLK(clk), .RST(rst), .I(in[49]), .Q(
        round_reg[49]) );
  DFF \round_reg_reg[50]  ( .D(out[50]), .CLK(clk), .RST(rst), .I(in[50]), .Q(
        round_reg[50]) );
  DFF \round_reg_reg[51]  ( .D(out[51]), .CLK(clk), .RST(rst), .I(in[51]), .Q(
        round_reg[51]) );
  DFF \round_reg_reg[52]  ( .D(out[52]), .CLK(clk), .RST(rst), .I(in[52]), .Q(
        round_reg[52]) );
  DFF \round_reg_reg[53]  ( .D(out[53]), .CLK(clk), .RST(rst), .I(in[53]), .Q(
        round_reg[53]) );
  DFF \round_reg_reg[54]  ( .D(out[54]), .CLK(clk), .RST(rst), .I(in[54]), .Q(
        round_reg[54]) );
  DFF \round_reg_reg[55]  ( .D(out[55]), .CLK(clk), .RST(rst), .I(in[55]), .Q(
        round_reg[55]) );
  DFF \round_reg_reg[56]  ( .D(out[56]), .CLK(clk), .RST(rst), .I(in[56]), .Q(
        round_reg[56]) );
  DFF \round_reg_reg[57]  ( .D(out[57]), .CLK(clk), .RST(rst), .I(in[57]), .Q(
        round_reg[57]) );
  DFF \round_reg_reg[58]  ( .D(out[58]), .CLK(clk), .RST(rst), .I(in[58]), .Q(
        round_reg[58]) );
  DFF \round_reg_reg[59]  ( .D(out[59]), .CLK(clk), .RST(rst), .I(in[59]), .Q(
        round_reg[59]) );
  DFF \round_reg_reg[60]  ( .D(out[60]), .CLK(clk), .RST(rst), .I(in[60]), .Q(
        round_reg[60]) );
  DFF \round_reg_reg[61]  ( .D(out[61]), .CLK(clk), .RST(rst), .I(in[61]), .Q(
        round_reg[61]) );
  DFF \round_reg_reg[62]  ( .D(out[62]), .CLK(clk), .RST(rst), .I(in[62]), .Q(
        round_reg[62]) );
  DFF \round_reg_reg[63]  ( .D(out[63]), .CLK(clk), .RST(rst), .I(in[63]), .Q(
        round_reg[63]) );
  DFF \round_reg_reg[64]  ( .D(out[64]), .CLK(clk), .RST(rst), .I(in[64]), .Q(
        round_reg[64]) );
  DFF \round_reg_reg[65]  ( .D(out[65]), .CLK(clk), .RST(rst), .I(in[65]), .Q(
        round_reg[65]) );
  DFF \round_reg_reg[66]  ( .D(out[66]), .CLK(clk), .RST(rst), .I(in[66]), .Q(
        round_reg[66]) );
  DFF \round_reg_reg[67]  ( .D(out[67]), .CLK(clk), .RST(rst), .I(in[67]), .Q(
        round_reg[67]) );
  DFF \round_reg_reg[68]  ( .D(out[68]), .CLK(clk), .RST(rst), .I(in[68]), .Q(
        round_reg[68]) );
  DFF \round_reg_reg[69]  ( .D(out[69]), .CLK(clk), .RST(rst), .I(in[69]), .Q(
        round_reg[69]) );
  DFF \round_reg_reg[70]  ( .D(out[70]), .CLK(clk), .RST(rst), .I(in[70]), .Q(
        round_reg[70]) );
  DFF \round_reg_reg[71]  ( .D(out[71]), .CLK(clk), .RST(rst), .I(in[71]), .Q(
        round_reg[71]) );
  DFF \round_reg_reg[72]  ( .D(out[72]), .CLK(clk), .RST(rst), .I(in[72]), .Q(
        round_reg[72]) );
  DFF \round_reg_reg[73]  ( .D(out[73]), .CLK(clk), .RST(rst), .I(in[73]), .Q(
        round_reg[73]) );
  DFF \round_reg_reg[74]  ( .D(out[74]), .CLK(clk), .RST(rst), .I(in[74]), .Q(
        round_reg[74]) );
  DFF \round_reg_reg[75]  ( .D(out[75]), .CLK(clk), .RST(rst), .I(in[75]), .Q(
        round_reg[75]) );
  DFF \round_reg_reg[76]  ( .D(out[76]), .CLK(clk), .RST(rst), .I(in[76]), .Q(
        round_reg[76]) );
  DFF \round_reg_reg[77]  ( .D(out[77]), .CLK(clk), .RST(rst), .I(in[77]), .Q(
        round_reg[77]) );
  DFF \round_reg_reg[78]  ( .D(out[78]), .CLK(clk), .RST(rst), .I(in[78]), .Q(
        round_reg[78]) );
  DFF \round_reg_reg[79]  ( .D(out[79]), .CLK(clk), .RST(rst), .I(in[79]), .Q(
        round_reg[79]) );
  DFF \round_reg_reg[80]  ( .D(out[80]), .CLK(clk), .RST(rst), .I(in[80]), .Q(
        round_reg[80]) );
  DFF \round_reg_reg[81]  ( .D(out[81]), .CLK(clk), .RST(rst), .I(in[81]), .Q(
        round_reg[81]) );
  DFF \round_reg_reg[82]  ( .D(out[82]), .CLK(clk), .RST(rst), .I(in[82]), .Q(
        round_reg[82]) );
  DFF \round_reg_reg[83]  ( .D(out[83]), .CLK(clk), .RST(rst), .I(in[83]), .Q(
        round_reg[83]) );
  DFF \round_reg_reg[84]  ( .D(out[84]), .CLK(clk), .RST(rst), .I(in[84]), .Q(
        round_reg[84]) );
  DFF \round_reg_reg[85]  ( .D(out[85]), .CLK(clk), .RST(rst), .I(in[85]), .Q(
        round_reg[85]) );
  DFF \round_reg_reg[86]  ( .D(out[86]), .CLK(clk), .RST(rst), .I(in[86]), .Q(
        round_reg[86]) );
  DFF \round_reg_reg[87]  ( .D(out[87]), .CLK(clk), .RST(rst), .I(in[87]), .Q(
        round_reg[87]) );
  DFF \round_reg_reg[88]  ( .D(out[88]), .CLK(clk), .RST(rst), .I(in[88]), .Q(
        round_reg[88]) );
  DFF \round_reg_reg[89]  ( .D(out[89]), .CLK(clk), .RST(rst), .I(in[89]), .Q(
        round_reg[89]) );
  DFF \round_reg_reg[90]  ( .D(out[90]), .CLK(clk), .RST(rst), .I(in[90]), .Q(
        round_reg[90]) );
  DFF \round_reg_reg[91]  ( .D(out[91]), .CLK(clk), .RST(rst), .I(in[91]), .Q(
        round_reg[91]) );
  DFF \round_reg_reg[92]  ( .D(out[92]), .CLK(clk), .RST(rst), .I(in[92]), .Q(
        round_reg[92]) );
  DFF \round_reg_reg[93]  ( .D(out[93]), .CLK(clk), .RST(rst), .I(in[93]), .Q(
        round_reg[93]) );
  DFF \round_reg_reg[94]  ( .D(out[94]), .CLK(clk), .RST(rst), .I(in[94]), .Q(
        round_reg[94]) );
  DFF \round_reg_reg[95]  ( .D(out[95]), .CLK(clk), .RST(rst), .I(in[95]), .Q(
        round_reg[95]) );
  DFF \round_reg_reg[96]  ( .D(out[96]), .CLK(clk), .RST(rst), .I(in[96]), .Q(
        round_reg[96]) );
  DFF \round_reg_reg[97]  ( .D(out[97]), .CLK(clk), .RST(rst), .I(in[97]), .Q(
        round_reg[97]) );
  DFF \round_reg_reg[98]  ( .D(out[98]), .CLK(clk), .RST(rst), .I(in[98]), .Q(
        round_reg[98]) );
  DFF \round_reg_reg[99]  ( .D(out[99]), .CLK(clk), .RST(rst), .I(in[99]), .Q(
        round_reg[99]) );
  DFF \round_reg_reg[100]  ( .D(out[100]), .CLK(clk), .RST(rst), .I(in[100]), 
        .Q(round_reg[100]) );
  DFF \round_reg_reg[101]  ( .D(out[101]), .CLK(clk), .RST(rst), .I(in[101]), 
        .Q(round_reg[101]) );
  DFF \round_reg_reg[102]  ( .D(out[102]), .CLK(clk), .RST(rst), .I(in[102]), 
        .Q(round_reg[102]) );
  DFF \round_reg_reg[103]  ( .D(out[103]), .CLK(clk), .RST(rst), .I(in[103]), 
        .Q(round_reg[103]) );
  DFF \round_reg_reg[104]  ( .D(out[104]), .CLK(clk), .RST(rst), .I(in[104]), 
        .Q(round_reg[104]) );
  DFF \round_reg_reg[105]  ( .D(out[105]), .CLK(clk), .RST(rst), .I(in[105]), 
        .Q(round_reg[105]) );
  DFF \round_reg_reg[106]  ( .D(out[106]), .CLK(clk), .RST(rst), .I(in[106]), 
        .Q(round_reg[106]) );
  DFF \round_reg_reg[107]  ( .D(out[107]), .CLK(clk), .RST(rst), .I(in[107]), 
        .Q(round_reg[107]) );
  DFF \round_reg_reg[108]  ( .D(out[108]), .CLK(clk), .RST(rst), .I(in[108]), 
        .Q(round_reg[108]) );
  DFF \round_reg_reg[109]  ( .D(out[109]), .CLK(clk), .RST(rst), .I(in[109]), 
        .Q(round_reg[109]) );
  DFF \round_reg_reg[110]  ( .D(out[110]), .CLK(clk), .RST(rst), .I(in[110]), 
        .Q(round_reg[110]) );
  DFF \round_reg_reg[111]  ( .D(out[111]), .CLK(clk), .RST(rst), .I(in[111]), 
        .Q(round_reg[111]) );
  DFF \round_reg_reg[112]  ( .D(out[112]), .CLK(clk), .RST(rst), .I(in[112]), 
        .Q(round_reg[112]) );
  DFF \round_reg_reg[113]  ( .D(out[113]), .CLK(clk), .RST(rst), .I(in[113]), 
        .Q(round_reg[113]) );
  DFF \round_reg_reg[114]  ( .D(out[114]), .CLK(clk), .RST(rst), .I(in[114]), 
        .Q(round_reg[114]) );
  DFF \round_reg_reg[115]  ( .D(out[115]), .CLK(clk), .RST(rst), .I(in[115]), 
        .Q(round_reg[115]) );
  DFF \round_reg_reg[116]  ( .D(out[116]), .CLK(clk), .RST(rst), .I(in[116]), 
        .Q(round_reg[116]) );
  DFF \round_reg_reg[117]  ( .D(out[117]), .CLK(clk), .RST(rst), .I(in[117]), 
        .Q(round_reg[117]) );
  DFF \round_reg_reg[118]  ( .D(out[118]), .CLK(clk), .RST(rst), .I(in[118]), 
        .Q(round_reg[118]) );
  DFF \round_reg_reg[119]  ( .D(out[119]), .CLK(clk), .RST(rst), .I(in[119]), 
        .Q(round_reg[119]) );
  DFF \round_reg_reg[120]  ( .D(out[120]), .CLK(clk), .RST(rst), .I(in[120]), 
        .Q(round_reg[120]) );
  DFF \round_reg_reg[121]  ( .D(out[121]), .CLK(clk), .RST(rst), .I(in[121]), 
        .Q(round_reg[121]) );
  DFF \round_reg_reg[122]  ( .D(out[122]), .CLK(clk), .RST(rst), .I(in[122]), 
        .Q(round_reg[122]) );
  DFF \round_reg_reg[123]  ( .D(out[123]), .CLK(clk), .RST(rst), .I(in[123]), 
        .Q(round_reg[123]) );
  DFF \round_reg_reg[124]  ( .D(out[124]), .CLK(clk), .RST(rst), .I(in[124]), 
        .Q(round_reg[124]) );
  DFF \round_reg_reg[125]  ( .D(out[125]), .CLK(clk), .RST(rst), .I(in[125]), 
        .Q(round_reg[125]) );
  DFF \round_reg_reg[126]  ( .D(out[126]), .CLK(clk), .RST(rst), .I(in[126]), 
        .Q(round_reg[126]) );
  DFF \round_reg_reg[127]  ( .D(out[127]), .CLK(clk), .RST(rst), .I(in[127]), 
        .Q(round_reg[127]) );
  DFF \round_reg_reg[128]  ( .D(out[128]), .CLK(clk), .RST(rst), .I(in[128]), 
        .Q(round_reg[128]) );
  DFF \round_reg_reg[129]  ( .D(out[129]), .CLK(clk), .RST(rst), .I(in[129]), 
        .Q(round_reg[129]) );
  DFF \round_reg_reg[130]  ( .D(out[130]), .CLK(clk), .RST(rst), .I(in[130]), 
        .Q(round_reg[130]) );
  DFF \round_reg_reg[131]  ( .D(out[131]), .CLK(clk), .RST(rst), .I(in[131]), 
        .Q(round_reg[131]) );
  DFF \round_reg_reg[132]  ( .D(out[132]), .CLK(clk), .RST(rst), .I(in[132]), 
        .Q(round_reg[132]) );
  DFF \round_reg_reg[133]  ( .D(out[133]), .CLK(clk), .RST(rst), .I(in[133]), 
        .Q(round_reg[133]) );
  DFF \round_reg_reg[134]  ( .D(out[134]), .CLK(clk), .RST(rst), .I(in[134]), 
        .Q(round_reg[134]) );
  DFF \round_reg_reg[135]  ( .D(out[135]), .CLK(clk), .RST(rst), .I(in[135]), 
        .Q(round_reg[135]) );
  DFF \round_reg_reg[136]  ( .D(out[136]), .CLK(clk), .RST(rst), .I(in[136]), 
        .Q(round_reg[136]) );
  DFF \round_reg_reg[137]  ( .D(out[137]), .CLK(clk), .RST(rst), .I(in[137]), 
        .Q(round_reg[137]) );
  DFF \round_reg_reg[138]  ( .D(out[138]), .CLK(clk), .RST(rst), .I(in[138]), 
        .Q(round_reg[138]) );
  DFF \round_reg_reg[139]  ( .D(out[139]), .CLK(clk), .RST(rst), .I(in[139]), 
        .Q(round_reg[139]) );
  DFF \round_reg_reg[140]  ( .D(out[140]), .CLK(clk), .RST(rst), .I(in[140]), 
        .Q(round_reg[140]) );
  DFF \round_reg_reg[141]  ( .D(out[141]), .CLK(clk), .RST(rst), .I(in[141]), 
        .Q(round_reg[141]) );
  DFF \round_reg_reg[142]  ( .D(out[142]), .CLK(clk), .RST(rst), .I(in[142]), 
        .Q(round_reg[142]) );
  DFF \round_reg_reg[143]  ( .D(out[143]), .CLK(clk), .RST(rst), .I(in[143]), 
        .Q(round_reg[143]) );
  DFF \round_reg_reg[144]  ( .D(out[144]), .CLK(clk), .RST(rst), .I(in[144]), 
        .Q(round_reg[144]) );
  DFF \round_reg_reg[145]  ( .D(out[145]), .CLK(clk), .RST(rst), .I(in[145]), 
        .Q(round_reg[145]) );
  DFF \round_reg_reg[146]  ( .D(out[146]), .CLK(clk), .RST(rst), .I(in[146]), 
        .Q(round_reg[146]) );
  DFF \round_reg_reg[147]  ( .D(out[147]), .CLK(clk), .RST(rst), .I(in[147]), 
        .Q(round_reg[147]) );
  DFF \round_reg_reg[148]  ( .D(out[148]), .CLK(clk), .RST(rst), .I(in[148]), 
        .Q(round_reg[148]) );
  DFF \round_reg_reg[149]  ( .D(out[149]), .CLK(clk), .RST(rst), .I(in[149]), 
        .Q(round_reg[149]) );
  DFF \round_reg_reg[150]  ( .D(out[150]), .CLK(clk), .RST(rst), .I(in[150]), 
        .Q(round_reg[150]) );
  DFF \round_reg_reg[151]  ( .D(out[151]), .CLK(clk), .RST(rst), .I(in[151]), 
        .Q(round_reg[151]) );
  DFF \round_reg_reg[152]  ( .D(out[152]), .CLK(clk), .RST(rst), .I(in[152]), 
        .Q(round_reg[152]) );
  DFF \round_reg_reg[153]  ( .D(out[153]), .CLK(clk), .RST(rst), .I(in[153]), 
        .Q(round_reg[153]) );
  DFF \round_reg_reg[154]  ( .D(out[154]), .CLK(clk), .RST(rst), .I(in[154]), 
        .Q(round_reg[154]) );
  DFF \round_reg_reg[155]  ( .D(out[155]), .CLK(clk), .RST(rst), .I(in[155]), 
        .Q(round_reg[155]) );
  DFF \round_reg_reg[156]  ( .D(out[156]), .CLK(clk), .RST(rst), .I(in[156]), 
        .Q(round_reg[156]) );
  DFF \round_reg_reg[157]  ( .D(out[157]), .CLK(clk), .RST(rst), .I(in[157]), 
        .Q(round_reg[157]) );
  DFF \round_reg_reg[158]  ( .D(out[158]), .CLK(clk), .RST(rst), .I(in[158]), 
        .Q(round_reg[158]) );
  DFF \round_reg_reg[159]  ( .D(out[159]), .CLK(clk), .RST(rst), .I(in[159]), 
        .Q(round_reg[159]) );
  DFF \round_reg_reg[160]  ( .D(out[160]), .CLK(clk), .RST(rst), .I(in[160]), 
        .Q(round_reg[160]) );
  DFF \round_reg_reg[161]  ( .D(out[161]), .CLK(clk), .RST(rst), .I(in[161]), 
        .Q(round_reg[161]) );
  DFF \round_reg_reg[162]  ( .D(out[162]), .CLK(clk), .RST(rst), .I(in[162]), 
        .Q(round_reg[162]) );
  DFF \round_reg_reg[163]  ( .D(out[163]), .CLK(clk), .RST(rst), .I(in[163]), 
        .Q(round_reg[163]) );
  DFF \round_reg_reg[164]  ( .D(out[164]), .CLK(clk), .RST(rst), .I(in[164]), 
        .Q(round_reg[164]) );
  DFF \round_reg_reg[165]  ( .D(out[165]), .CLK(clk), .RST(rst), .I(in[165]), 
        .Q(round_reg[165]) );
  DFF \round_reg_reg[166]  ( .D(out[166]), .CLK(clk), .RST(rst), .I(in[166]), 
        .Q(round_reg[166]) );
  DFF \round_reg_reg[167]  ( .D(out[167]), .CLK(clk), .RST(rst), .I(in[167]), 
        .Q(round_reg[167]) );
  DFF \round_reg_reg[168]  ( .D(out[168]), .CLK(clk), .RST(rst), .I(in[168]), 
        .Q(round_reg[168]) );
  DFF \round_reg_reg[169]  ( .D(out[169]), .CLK(clk), .RST(rst), .I(in[169]), 
        .Q(round_reg[169]) );
  DFF \round_reg_reg[170]  ( .D(out[170]), .CLK(clk), .RST(rst), .I(in[170]), 
        .Q(round_reg[170]) );
  DFF \round_reg_reg[171]  ( .D(out[171]), .CLK(clk), .RST(rst), .I(in[171]), 
        .Q(round_reg[171]) );
  DFF \round_reg_reg[172]  ( .D(out[172]), .CLK(clk), .RST(rst), .I(in[172]), 
        .Q(round_reg[172]) );
  DFF \round_reg_reg[173]  ( .D(out[173]), .CLK(clk), .RST(rst), .I(in[173]), 
        .Q(round_reg[173]) );
  DFF \round_reg_reg[174]  ( .D(out[174]), .CLK(clk), .RST(rst), .I(in[174]), 
        .Q(round_reg[174]) );
  DFF \round_reg_reg[175]  ( .D(out[175]), .CLK(clk), .RST(rst), .I(in[175]), 
        .Q(round_reg[175]) );
  DFF \round_reg_reg[176]  ( .D(out[176]), .CLK(clk), .RST(rst), .I(in[176]), 
        .Q(round_reg[176]) );
  DFF \round_reg_reg[177]  ( .D(out[177]), .CLK(clk), .RST(rst), .I(in[177]), 
        .Q(round_reg[177]) );
  DFF \round_reg_reg[178]  ( .D(out[178]), .CLK(clk), .RST(rst), .I(in[178]), 
        .Q(round_reg[178]) );
  DFF \round_reg_reg[179]  ( .D(out[179]), .CLK(clk), .RST(rst), .I(in[179]), 
        .Q(round_reg[179]) );
  DFF \round_reg_reg[180]  ( .D(out[180]), .CLK(clk), .RST(rst), .I(in[180]), 
        .Q(round_reg[180]) );
  DFF \round_reg_reg[181]  ( .D(out[181]), .CLK(clk), .RST(rst), .I(in[181]), 
        .Q(round_reg[181]) );
  DFF \round_reg_reg[182]  ( .D(out[182]), .CLK(clk), .RST(rst), .I(in[182]), 
        .Q(round_reg[182]) );
  DFF \round_reg_reg[183]  ( .D(out[183]), .CLK(clk), .RST(rst), .I(in[183]), 
        .Q(round_reg[183]) );
  DFF \round_reg_reg[184]  ( .D(out[184]), .CLK(clk), .RST(rst), .I(in[184]), 
        .Q(round_reg[184]) );
  DFF \round_reg_reg[185]  ( .D(out[185]), .CLK(clk), .RST(rst), .I(in[185]), 
        .Q(round_reg[185]) );
  DFF \round_reg_reg[186]  ( .D(out[186]), .CLK(clk), .RST(rst), .I(in[186]), 
        .Q(round_reg[186]) );
  DFF \round_reg_reg[187]  ( .D(out[187]), .CLK(clk), .RST(rst), .I(in[187]), 
        .Q(round_reg[187]) );
  DFF \round_reg_reg[188]  ( .D(out[188]), .CLK(clk), .RST(rst), .I(in[188]), 
        .Q(round_reg[188]) );
  DFF \round_reg_reg[189]  ( .D(out[189]), .CLK(clk), .RST(rst), .I(in[189]), 
        .Q(round_reg[189]) );
  DFF \round_reg_reg[190]  ( .D(out[190]), .CLK(clk), .RST(rst), .I(in[190]), 
        .Q(round_reg[190]) );
  DFF \round_reg_reg[191]  ( .D(out[191]), .CLK(clk), .RST(rst), .I(in[191]), 
        .Q(round_reg[191]) );
  DFF \round_reg_reg[192]  ( .D(out[192]), .CLK(clk), .RST(rst), .I(in[192]), 
        .Q(round_reg[192]) );
  DFF \round_reg_reg[193]  ( .D(out[193]), .CLK(clk), .RST(rst), .I(in[193]), 
        .Q(round_reg[193]) );
  DFF \round_reg_reg[194]  ( .D(out[194]), .CLK(clk), .RST(rst), .I(in[194]), 
        .Q(round_reg[194]) );
  DFF \round_reg_reg[195]  ( .D(out[195]), .CLK(clk), .RST(rst), .I(in[195]), 
        .Q(round_reg[195]) );
  DFF \round_reg_reg[196]  ( .D(out[196]), .CLK(clk), .RST(rst), .I(in[196]), 
        .Q(round_reg[196]) );
  DFF \round_reg_reg[197]  ( .D(out[197]), .CLK(clk), .RST(rst), .I(in[197]), 
        .Q(round_reg[197]) );
  DFF \round_reg_reg[198]  ( .D(out[198]), .CLK(clk), .RST(rst), .I(in[198]), 
        .Q(round_reg[198]) );
  DFF \round_reg_reg[199]  ( .D(out[199]), .CLK(clk), .RST(rst), .I(in[199]), 
        .Q(round_reg[199]) );
  DFF \round_reg_reg[200]  ( .D(out[200]), .CLK(clk), .RST(rst), .I(in[200]), 
        .Q(round_reg[200]) );
  DFF \round_reg_reg[201]  ( .D(out[201]), .CLK(clk), .RST(rst), .I(in[201]), 
        .Q(round_reg[201]) );
  DFF \round_reg_reg[202]  ( .D(out[202]), .CLK(clk), .RST(rst), .I(in[202]), 
        .Q(round_reg[202]) );
  DFF \round_reg_reg[203]  ( .D(out[203]), .CLK(clk), .RST(rst), .I(in[203]), 
        .Q(round_reg[203]) );
  DFF \round_reg_reg[204]  ( .D(out[204]), .CLK(clk), .RST(rst), .I(in[204]), 
        .Q(round_reg[204]) );
  DFF \round_reg_reg[205]  ( .D(out[205]), .CLK(clk), .RST(rst), .I(in[205]), 
        .Q(round_reg[205]) );
  DFF \round_reg_reg[206]  ( .D(out[206]), .CLK(clk), .RST(rst), .I(in[206]), 
        .Q(round_reg[206]) );
  DFF \round_reg_reg[207]  ( .D(out[207]), .CLK(clk), .RST(rst), .I(in[207]), 
        .Q(round_reg[207]) );
  DFF \round_reg_reg[208]  ( .D(out[208]), .CLK(clk), .RST(rst), .I(in[208]), 
        .Q(round_reg[208]) );
  DFF \round_reg_reg[209]  ( .D(out[209]), .CLK(clk), .RST(rst), .I(in[209]), 
        .Q(round_reg[209]) );
  DFF \round_reg_reg[210]  ( .D(out[210]), .CLK(clk), .RST(rst), .I(in[210]), 
        .Q(round_reg[210]) );
  DFF \round_reg_reg[211]  ( .D(out[211]), .CLK(clk), .RST(rst), .I(in[211]), 
        .Q(round_reg[211]) );
  DFF \round_reg_reg[212]  ( .D(out[212]), .CLK(clk), .RST(rst), .I(in[212]), 
        .Q(round_reg[212]) );
  DFF \round_reg_reg[213]  ( .D(out[213]), .CLK(clk), .RST(rst), .I(in[213]), 
        .Q(round_reg[213]) );
  DFF \round_reg_reg[214]  ( .D(out[214]), .CLK(clk), .RST(rst), .I(in[214]), 
        .Q(round_reg[214]) );
  DFF \round_reg_reg[215]  ( .D(out[215]), .CLK(clk), .RST(rst), .I(in[215]), 
        .Q(round_reg[215]) );
  DFF \round_reg_reg[216]  ( .D(out[216]), .CLK(clk), .RST(rst), .I(in[216]), 
        .Q(round_reg[216]) );
  DFF \round_reg_reg[217]  ( .D(out[217]), .CLK(clk), .RST(rst), .I(in[217]), 
        .Q(round_reg[217]) );
  DFF \round_reg_reg[218]  ( .D(out[218]), .CLK(clk), .RST(rst), .I(in[218]), 
        .Q(round_reg[218]) );
  DFF \round_reg_reg[219]  ( .D(out[219]), .CLK(clk), .RST(rst), .I(in[219]), 
        .Q(round_reg[219]) );
  DFF \round_reg_reg[220]  ( .D(out[220]), .CLK(clk), .RST(rst), .I(in[220]), 
        .Q(round_reg[220]) );
  DFF \round_reg_reg[221]  ( .D(out[221]), .CLK(clk), .RST(rst), .I(in[221]), 
        .Q(round_reg[221]) );
  DFF \round_reg_reg[222]  ( .D(out[222]), .CLK(clk), .RST(rst), .I(in[222]), 
        .Q(round_reg[222]) );
  DFF \round_reg_reg[223]  ( .D(out[223]), .CLK(clk), .RST(rst), .I(in[223]), 
        .Q(round_reg[223]) );
  DFF \round_reg_reg[224]  ( .D(out[224]), .CLK(clk), .RST(rst), .I(in[224]), 
        .Q(round_reg[224]) );
  DFF \round_reg_reg[225]  ( .D(out[225]), .CLK(clk), .RST(rst), .I(in[225]), 
        .Q(round_reg[225]) );
  DFF \round_reg_reg[226]  ( .D(out[226]), .CLK(clk), .RST(rst), .I(in[226]), 
        .Q(round_reg[226]) );
  DFF \round_reg_reg[227]  ( .D(out[227]), .CLK(clk), .RST(rst), .I(in[227]), 
        .Q(round_reg[227]) );
  DFF \round_reg_reg[228]  ( .D(out[228]), .CLK(clk), .RST(rst), .I(in[228]), 
        .Q(round_reg[228]) );
  DFF \round_reg_reg[229]  ( .D(out[229]), .CLK(clk), .RST(rst), .I(in[229]), 
        .Q(round_reg[229]) );
  DFF \round_reg_reg[230]  ( .D(out[230]), .CLK(clk), .RST(rst), .I(in[230]), 
        .Q(round_reg[230]) );
  DFF \round_reg_reg[231]  ( .D(out[231]), .CLK(clk), .RST(rst), .I(in[231]), 
        .Q(round_reg[231]) );
  DFF \round_reg_reg[232]  ( .D(out[232]), .CLK(clk), .RST(rst), .I(in[232]), 
        .Q(round_reg[232]) );
  DFF \round_reg_reg[233]  ( .D(out[233]), .CLK(clk), .RST(rst), .I(in[233]), 
        .Q(round_reg[233]) );
  DFF \round_reg_reg[234]  ( .D(out[234]), .CLK(clk), .RST(rst), .I(in[234]), 
        .Q(round_reg[234]) );
  DFF \round_reg_reg[235]  ( .D(out[235]), .CLK(clk), .RST(rst), .I(in[235]), 
        .Q(round_reg[235]) );
  DFF \round_reg_reg[236]  ( .D(out[236]), .CLK(clk), .RST(rst), .I(in[236]), 
        .Q(round_reg[236]) );
  DFF \round_reg_reg[237]  ( .D(out[237]), .CLK(clk), .RST(rst), .I(in[237]), 
        .Q(round_reg[237]) );
  DFF \round_reg_reg[238]  ( .D(out[238]), .CLK(clk), .RST(rst), .I(in[238]), 
        .Q(round_reg[238]) );
  DFF \round_reg_reg[239]  ( .D(out[239]), .CLK(clk), .RST(rst), .I(in[239]), 
        .Q(round_reg[239]) );
  DFF \round_reg_reg[240]  ( .D(out[240]), .CLK(clk), .RST(rst), .I(in[240]), 
        .Q(round_reg[240]) );
  DFF \round_reg_reg[241]  ( .D(out[241]), .CLK(clk), .RST(rst), .I(in[241]), 
        .Q(round_reg[241]) );
  DFF \round_reg_reg[242]  ( .D(out[242]), .CLK(clk), .RST(rst), .I(in[242]), 
        .Q(round_reg[242]) );
  DFF \round_reg_reg[243]  ( .D(out[243]), .CLK(clk), .RST(rst), .I(in[243]), 
        .Q(round_reg[243]) );
  DFF \round_reg_reg[244]  ( .D(out[244]), .CLK(clk), .RST(rst), .I(in[244]), 
        .Q(round_reg[244]) );
  DFF \round_reg_reg[245]  ( .D(out[245]), .CLK(clk), .RST(rst), .I(in[245]), 
        .Q(round_reg[245]) );
  DFF \round_reg_reg[246]  ( .D(out[246]), .CLK(clk), .RST(rst), .I(in[246]), 
        .Q(round_reg[246]) );
  DFF \round_reg_reg[247]  ( .D(out[247]), .CLK(clk), .RST(rst), .I(in[247]), 
        .Q(round_reg[247]) );
  DFF \round_reg_reg[248]  ( .D(out[248]), .CLK(clk), .RST(rst), .I(in[248]), 
        .Q(round_reg[248]) );
  DFF \round_reg_reg[249]  ( .D(out[249]), .CLK(clk), .RST(rst), .I(in[249]), 
        .Q(round_reg[249]) );
  DFF \round_reg_reg[250]  ( .D(out[250]), .CLK(clk), .RST(rst), .I(in[250]), 
        .Q(round_reg[250]) );
  DFF \round_reg_reg[251]  ( .D(out[251]), .CLK(clk), .RST(rst), .I(in[251]), 
        .Q(round_reg[251]) );
  DFF \round_reg_reg[252]  ( .D(out[252]), .CLK(clk), .RST(rst), .I(in[252]), 
        .Q(round_reg[252]) );
  DFF \round_reg_reg[253]  ( .D(out[253]), .CLK(clk), .RST(rst), .I(in[253]), 
        .Q(round_reg[253]) );
  DFF \round_reg_reg[254]  ( .D(out[254]), .CLK(clk), .RST(rst), .I(in[254]), 
        .Q(round_reg[254]) );
  DFF \round_reg_reg[255]  ( .D(out[255]), .CLK(clk), .RST(rst), .I(in[255]), 
        .Q(round_reg[255]) );
  DFF \round_reg_reg[256]  ( .D(out[256]), .CLK(clk), .RST(rst), .I(in[256]), 
        .Q(round_reg[256]) );
  DFF \round_reg_reg[257]  ( .D(out[257]), .CLK(clk), .RST(rst), .I(in[257]), 
        .Q(round_reg[257]) );
  DFF \round_reg_reg[258]  ( .D(out[258]), .CLK(clk), .RST(rst), .I(in[258]), 
        .Q(round_reg[258]) );
  DFF \round_reg_reg[259]  ( .D(out[259]), .CLK(clk), .RST(rst), .I(in[259]), 
        .Q(round_reg[259]) );
  DFF \round_reg_reg[260]  ( .D(out[260]), .CLK(clk), .RST(rst), .I(in[260]), 
        .Q(round_reg[260]) );
  DFF \round_reg_reg[261]  ( .D(out[261]), .CLK(clk), .RST(rst), .I(in[261]), 
        .Q(round_reg[261]) );
  DFF \round_reg_reg[262]  ( .D(out[262]), .CLK(clk), .RST(rst), .I(in[262]), 
        .Q(round_reg[262]) );
  DFF \round_reg_reg[263]  ( .D(out[263]), .CLK(clk), .RST(rst), .I(in[263]), 
        .Q(round_reg[263]) );
  DFF \round_reg_reg[264]  ( .D(out[264]), .CLK(clk), .RST(rst), .I(in[264]), 
        .Q(round_reg[264]) );
  DFF \round_reg_reg[265]  ( .D(out[265]), .CLK(clk), .RST(rst), .I(in[265]), 
        .Q(round_reg[265]) );
  DFF \round_reg_reg[266]  ( .D(out[266]), .CLK(clk), .RST(rst), .I(in[266]), 
        .Q(round_reg[266]) );
  DFF \round_reg_reg[267]  ( .D(out[267]), .CLK(clk), .RST(rst), .I(in[267]), 
        .Q(round_reg[267]) );
  DFF \round_reg_reg[268]  ( .D(out[268]), .CLK(clk), .RST(rst), .I(in[268]), 
        .Q(round_reg[268]) );
  DFF \round_reg_reg[269]  ( .D(out[269]), .CLK(clk), .RST(rst), .I(in[269]), 
        .Q(round_reg[269]) );
  DFF \round_reg_reg[270]  ( .D(out[270]), .CLK(clk), .RST(rst), .I(in[270]), 
        .Q(round_reg[270]) );
  DFF \round_reg_reg[271]  ( .D(out[271]), .CLK(clk), .RST(rst), .I(in[271]), 
        .Q(round_reg[271]) );
  DFF \round_reg_reg[272]  ( .D(out[272]), .CLK(clk), .RST(rst), .I(in[272]), 
        .Q(round_reg[272]) );
  DFF \round_reg_reg[273]  ( .D(out[273]), .CLK(clk), .RST(rst), .I(in[273]), 
        .Q(round_reg[273]) );
  DFF \round_reg_reg[274]  ( .D(out[274]), .CLK(clk), .RST(rst), .I(in[274]), 
        .Q(round_reg[274]) );
  DFF \round_reg_reg[275]  ( .D(out[275]), .CLK(clk), .RST(rst), .I(in[275]), 
        .Q(round_reg[275]) );
  DFF \round_reg_reg[276]  ( .D(out[276]), .CLK(clk), .RST(rst), .I(in[276]), 
        .Q(round_reg[276]) );
  DFF \round_reg_reg[277]  ( .D(out[277]), .CLK(clk), .RST(rst), .I(in[277]), 
        .Q(round_reg[277]) );
  DFF \round_reg_reg[278]  ( .D(out[278]), .CLK(clk), .RST(rst), .I(in[278]), 
        .Q(round_reg[278]) );
  DFF \round_reg_reg[279]  ( .D(out[279]), .CLK(clk), .RST(rst), .I(in[279]), 
        .Q(round_reg[279]) );
  DFF \round_reg_reg[280]  ( .D(out[280]), .CLK(clk), .RST(rst), .I(in[280]), 
        .Q(round_reg[280]) );
  DFF \round_reg_reg[281]  ( .D(out[281]), .CLK(clk), .RST(rst), .I(in[281]), 
        .Q(round_reg[281]) );
  DFF \round_reg_reg[282]  ( .D(out[282]), .CLK(clk), .RST(rst), .I(in[282]), 
        .Q(round_reg[282]) );
  DFF \round_reg_reg[283]  ( .D(out[283]), .CLK(clk), .RST(rst), .I(in[283]), 
        .Q(round_reg[283]) );
  DFF \round_reg_reg[284]  ( .D(out[284]), .CLK(clk), .RST(rst), .I(in[284]), 
        .Q(round_reg[284]) );
  DFF \round_reg_reg[285]  ( .D(out[285]), .CLK(clk), .RST(rst), .I(in[285]), 
        .Q(round_reg[285]) );
  DFF \round_reg_reg[286]  ( .D(out[286]), .CLK(clk), .RST(rst), .I(in[286]), 
        .Q(round_reg[286]) );
  DFF \round_reg_reg[287]  ( .D(out[287]), .CLK(clk), .RST(rst), .I(in[287]), 
        .Q(round_reg[287]) );
  DFF \round_reg_reg[288]  ( .D(out[288]), .CLK(clk), .RST(rst), .I(in[288]), 
        .Q(round_reg[288]) );
  DFF \round_reg_reg[289]  ( .D(out[289]), .CLK(clk), .RST(rst), .I(in[289]), 
        .Q(round_reg[289]) );
  DFF \round_reg_reg[290]  ( .D(out[290]), .CLK(clk), .RST(rst), .I(in[290]), 
        .Q(round_reg[290]) );
  DFF \round_reg_reg[291]  ( .D(out[291]), .CLK(clk), .RST(rst), .I(in[291]), 
        .Q(round_reg[291]) );
  DFF \round_reg_reg[292]  ( .D(out[292]), .CLK(clk), .RST(rst), .I(in[292]), 
        .Q(round_reg[292]) );
  DFF \round_reg_reg[293]  ( .D(out[293]), .CLK(clk), .RST(rst), .I(in[293]), 
        .Q(round_reg[293]) );
  DFF \round_reg_reg[294]  ( .D(out[294]), .CLK(clk), .RST(rst), .I(in[294]), 
        .Q(round_reg[294]) );
  DFF \round_reg_reg[295]  ( .D(out[295]), .CLK(clk), .RST(rst), .I(in[295]), 
        .Q(round_reg[295]) );
  DFF \round_reg_reg[296]  ( .D(out[296]), .CLK(clk), .RST(rst), .I(in[296]), 
        .Q(round_reg[296]) );
  DFF \round_reg_reg[297]  ( .D(out[297]), .CLK(clk), .RST(rst), .I(in[297]), 
        .Q(round_reg[297]) );
  DFF \round_reg_reg[298]  ( .D(out[298]), .CLK(clk), .RST(rst), .I(in[298]), 
        .Q(round_reg[298]) );
  DFF \round_reg_reg[299]  ( .D(out[299]), .CLK(clk), .RST(rst), .I(in[299]), 
        .Q(round_reg[299]) );
  DFF \round_reg_reg[300]  ( .D(out[300]), .CLK(clk), .RST(rst), .I(in[300]), 
        .Q(round_reg[300]) );
  DFF \round_reg_reg[301]  ( .D(out[301]), .CLK(clk), .RST(rst), .I(in[301]), 
        .Q(round_reg[301]) );
  DFF \round_reg_reg[302]  ( .D(out[302]), .CLK(clk), .RST(rst), .I(in[302]), 
        .Q(round_reg[302]) );
  DFF \round_reg_reg[303]  ( .D(out[303]), .CLK(clk), .RST(rst), .I(in[303]), 
        .Q(round_reg[303]) );
  DFF \round_reg_reg[304]  ( .D(out[304]), .CLK(clk), .RST(rst), .I(in[304]), 
        .Q(round_reg[304]) );
  DFF \round_reg_reg[305]  ( .D(out[305]), .CLK(clk), .RST(rst), .I(in[305]), 
        .Q(round_reg[305]) );
  DFF \round_reg_reg[306]  ( .D(out[306]), .CLK(clk), .RST(rst), .I(in[306]), 
        .Q(round_reg[306]) );
  DFF \round_reg_reg[307]  ( .D(out[307]), .CLK(clk), .RST(rst), .I(in[307]), 
        .Q(round_reg[307]) );
  DFF \round_reg_reg[308]  ( .D(out[308]), .CLK(clk), .RST(rst), .I(in[308]), 
        .Q(round_reg[308]) );
  DFF \round_reg_reg[309]  ( .D(out[309]), .CLK(clk), .RST(rst), .I(in[309]), 
        .Q(round_reg[309]) );
  DFF \round_reg_reg[310]  ( .D(out[310]), .CLK(clk), .RST(rst), .I(in[310]), 
        .Q(round_reg[310]) );
  DFF \round_reg_reg[311]  ( .D(out[311]), .CLK(clk), .RST(rst), .I(in[311]), 
        .Q(round_reg[311]) );
  DFF \round_reg_reg[312]  ( .D(out[312]), .CLK(clk), .RST(rst), .I(in[312]), 
        .Q(round_reg[312]) );
  DFF \round_reg_reg[313]  ( .D(out[313]), .CLK(clk), .RST(rst), .I(in[313]), 
        .Q(round_reg[313]) );
  DFF \round_reg_reg[314]  ( .D(out[314]), .CLK(clk), .RST(rst), .I(in[314]), 
        .Q(round_reg[314]) );
  DFF \round_reg_reg[315]  ( .D(out[315]), .CLK(clk), .RST(rst), .I(in[315]), 
        .Q(round_reg[315]) );
  DFF \round_reg_reg[316]  ( .D(out[316]), .CLK(clk), .RST(rst), .I(in[316]), 
        .Q(round_reg[316]) );
  DFF \round_reg_reg[317]  ( .D(out[317]), .CLK(clk), .RST(rst), .I(in[317]), 
        .Q(round_reg[317]) );
  DFF \round_reg_reg[318]  ( .D(out[318]), .CLK(clk), .RST(rst), .I(in[318]), 
        .Q(round_reg[318]) );
  DFF \round_reg_reg[319]  ( .D(out[319]), .CLK(clk), .RST(rst), .I(in[319]), 
        .Q(round_reg[319]) );
  DFF \round_reg_reg[320]  ( .D(out[320]), .CLK(clk), .RST(rst), .I(in[320]), 
        .Q(round_reg[320]) );
  DFF \round_reg_reg[321]  ( .D(out[321]), .CLK(clk), .RST(rst), .I(in[321]), 
        .Q(round_reg[321]) );
  DFF \round_reg_reg[322]  ( .D(out[322]), .CLK(clk), .RST(rst), .I(in[322]), 
        .Q(round_reg[322]) );
  DFF \round_reg_reg[323]  ( .D(out[323]), .CLK(clk), .RST(rst), .I(in[323]), 
        .Q(round_reg[323]) );
  DFF \round_reg_reg[324]  ( .D(out[324]), .CLK(clk), .RST(rst), .I(in[324]), 
        .Q(round_reg[324]) );
  DFF \round_reg_reg[325]  ( .D(out[325]), .CLK(clk), .RST(rst), .I(in[325]), 
        .Q(round_reg[325]) );
  DFF \round_reg_reg[326]  ( .D(out[326]), .CLK(clk), .RST(rst), .I(in[326]), 
        .Q(round_reg[326]) );
  DFF \round_reg_reg[327]  ( .D(out[327]), .CLK(clk), .RST(rst), .I(in[327]), 
        .Q(round_reg[327]) );
  DFF \round_reg_reg[328]  ( .D(out[328]), .CLK(clk), .RST(rst), .I(in[328]), 
        .Q(round_reg[328]) );
  DFF \round_reg_reg[329]  ( .D(out[329]), .CLK(clk), .RST(rst), .I(in[329]), 
        .Q(round_reg[329]) );
  DFF \round_reg_reg[330]  ( .D(out[330]), .CLK(clk), .RST(rst), .I(in[330]), 
        .Q(round_reg[330]) );
  DFF \round_reg_reg[331]  ( .D(out[331]), .CLK(clk), .RST(rst), .I(in[331]), 
        .Q(round_reg[331]) );
  DFF \round_reg_reg[332]  ( .D(out[332]), .CLK(clk), .RST(rst), .I(in[332]), 
        .Q(round_reg[332]) );
  DFF \round_reg_reg[333]  ( .D(out[333]), .CLK(clk), .RST(rst), .I(in[333]), 
        .Q(round_reg[333]) );
  DFF \round_reg_reg[334]  ( .D(out[334]), .CLK(clk), .RST(rst), .I(in[334]), 
        .Q(round_reg[334]) );
  DFF \round_reg_reg[335]  ( .D(out[335]), .CLK(clk), .RST(rst), .I(in[335]), 
        .Q(round_reg[335]) );
  DFF \round_reg_reg[336]  ( .D(out[336]), .CLK(clk), .RST(rst), .I(in[336]), 
        .Q(round_reg[336]) );
  DFF \round_reg_reg[337]  ( .D(out[337]), .CLK(clk), .RST(rst), .I(in[337]), 
        .Q(round_reg[337]) );
  DFF \round_reg_reg[338]  ( .D(out[338]), .CLK(clk), .RST(rst), .I(in[338]), 
        .Q(round_reg[338]) );
  DFF \round_reg_reg[339]  ( .D(out[339]), .CLK(clk), .RST(rst), .I(in[339]), 
        .Q(round_reg[339]) );
  DFF \round_reg_reg[340]  ( .D(out[340]), .CLK(clk), .RST(rst), .I(in[340]), 
        .Q(round_reg[340]) );
  DFF \round_reg_reg[341]  ( .D(out[341]), .CLK(clk), .RST(rst), .I(in[341]), 
        .Q(round_reg[341]) );
  DFF \round_reg_reg[342]  ( .D(out[342]), .CLK(clk), .RST(rst), .I(in[342]), 
        .Q(round_reg[342]) );
  DFF \round_reg_reg[343]  ( .D(out[343]), .CLK(clk), .RST(rst), .I(in[343]), 
        .Q(round_reg[343]) );
  DFF \round_reg_reg[344]  ( .D(out[344]), .CLK(clk), .RST(rst), .I(in[344]), 
        .Q(round_reg[344]) );
  DFF \round_reg_reg[345]  ( .D(out[345]), .CLK(clk), .RST(rst), .I(in[345]), 
        .Q(round_reg[345]) );
  DFF \round_reg_reg[346]  ( .D(out[346]), .CLK(clk), .RST(rst), .I(in[346]), 
        .Q(round_reg[346]) );
  DFF \round_reg_reg[347]  ( .D(out[347]), .CLK(clk), .RST(rst), .I(in[347]), 
        .Q(round_reg[347]) );
  DFF \round_reg_reg[348]  ( .D(out[348]), .CLK(clk), .RST(rst), .I(in[348]), 
        .Q(round_reg[348]) );
  DFF \round_reg_reg[349]  ( .D(out[349]), .CLK(clk), .RST(rst), .I(in[349]), 
        .Q(round_reg[349]) );
  DFF \round_reg_reg[350]  ( .D(out[350]), .CLK(clk), .RST(rst), .I(in[350]), 
        .Q(round_reg[350]) );
  DFF \round_reg_reg[351]  ( .D(out[351]), .CLK(clk), .RST(rst), .I(in[351]), 
        .Q(round_reg[351]) );
  DFF \round_reg_reg[352]  ( .D(out[352]), .CLK(clk), .RST(rst), .I(in[352]), 
        .Q(round_reg[352]) );
  DFF \round_reg_reg[353]  ( .D(out[353]), .CLK(clk), .RST(rst), .I(in[353]), 
        .Q(round_reg[353]) );
  DFF \round_reg_reg[354]  ( .D(out[354]), .CLK(clk), .RST(rst), .I(in[354]), 
        .Q(round_reg[354]) );
  DFF \round_reg_reg[355]  ( .D(out[355]), .CLK(clk), .RST(rst), .I(in[355]), 
        .Q(round_reg[355]) );
  DFF \round_reg_reg[356]  ( .D(out[356]), .CLK(clk), .RST(rst), .I(in[356]), 
        .Q(round_reg[356]) );
  DFF \round_reg_reg[357]  ( .D(out[357]), .CLK(clk), .RST(rst), .I(in[357]), 
        .Q(round_reg[357]) );
  DFF \round_reg_reg[358]  ( .D(out[358]), .CLK(clk), .RST(rst), .I(in[358]), 
        .Q(round_reg[358]) );
  DFF \round_reg_reg[359]  ( .D(out[359]), .CLK(clk), .RST(rst), .I(in[359]), 
        .Q(round_reg[359]) );
  DFF \round_reg_reg[360]  ( .D(out[360]), .CLK(clk), .RST(rst), .I(in[360]), 
        .Q(round_reg[360]) );
  DFF \round_reg_reg[361]  ( .D(out[361]), .CLK(clk), .RST(rst), .I(in[361]), 
        .Q(round_reg[361]) );
  DFF \round_reg_reg[362]  ( .D(out[362]), .CLK(clk), .RST(rst), .I(in[362]), 
        .Q(round_reg[362]) );
  DFF \round_reg_reg[363]  ( .D(out[363]), .CLK(clk), .RST(rst), .I(in[363]), 
        .Q(round_reg[363]) );
  DFF \round_reg_reg[364]  ( .D(out[364]), .CLK(clk), .RST(rst), .I(in[364]), 
        .Q(round_reg[364]) );
  DFF \round_reg_reg[365]  ( .D(out[365]), .CLK(clk), .RST(rst), .I(in[365]), 
        .Q(round_reg[365]) );
  DFF \round_reg_reg[366]  ( .D(out[366]), .CLK(clk), .RST(rst), .I(in[366]), 
        .Q(round_reg[366]) );
  DFF \round_reg_reg[367]  ( .D(out[367]), .CLK(clk), .RST(rst), .I(in[367]), 
        .Q(round_reg[367]) );
  DFF \round_reg_reg[368]  ( .D(out[368]), .CLK(clk), .RST(rst), .I(in[368]), 
        .Q(round_reg[368]) );
  DFF \round_reg_reg[369]  ( .D(out[369]), .CLK(clk), .RST(rst), .I(in[369]), 
        .Q(round_reg[369]) );
  DFF \round_reg_reg[370]  ( .D(out[370]), .CLK(clk), .RST(rst), .I(in[370]), 
        .Q(round_reg[370]) );
  DFF \round_reg_reg[371]  ( .D(out[371]), .CLK(clk), .RST(rst), .I(in[371]), 
        .Q(round_reg[371]) );
  DFF \round_reg_reg[372]  ( .D(out[372]), .CLK(clk), .RST(rst), .I(in[372]), 
        .Q(round_reg[372]) );
  DFF \round_reg_reg[373]  ( .D(out[373]), .CLK(clk), .RST(rst), .I(in[373]), 
        .Q(round_reg[373]) );
  DFF \round_reg_reg[374]  ( .D(out[374]), .CLK(clk), .RST(rst), .I(in[374]), 
        .Q(round_reg[374]) );
  DFF \round_reg_reg[375]  ( .D(out[375]), .CLK(clk), .RST(rst), .I(in[375]), 
        .Q(round_reg[375]) );
  DFF \round_reg_reg[376]  ( .D(out[376]), .CLK(clk), .RST(rst), .I(in[376]), 
        .Q(round_reg[376]) );
  DFF \round_reg_reg[377]  ( .D(out[377]), .CLK(clk), .RST(rst), .I(in[377]), 
        .Q(round_reg[377]) );
  DFF \round_reg_reg[378]  ( .D(out[378]), .CLK(clk), .RST(rst), .I(in[378]), 
        .Q(round_reg[378]) );
  DFF \round_reg_reg[379]  ( .D(out[379]), .CLK(clk), .RST(rst), .I(in[379]), 
        .Q(round_reg[379]) );
  DFF \round_reg_reg[380]  ( .D(out[380]), .CLK(clk), .RST(rst), .I(in[380]), 
        .Q(round_reg[380]) );
  DFF \round_reg_reg[381]  ( .D(out[381]), .CLK(clk), .RST(rst), .I(in[381]), 
        .Q(round_reg[381]) );
  DFF \round_reg_reg[382]  ( .D(out[382]), .CLK(clk), .RST(rst), .I(in[382]), 
        .Q(round_reg[382]) );
  DFF \round_reg_reg[383]  ( .D(out[383]), .CLK(clk), .RST(rst), .I(in[383]), 
        .Q(round_reg[383]) );
  DFF \round_reg_reg[384]  ( .D(out[384]), .CLK(clk), .RST(rst), .I(in[384]), 
        .Q(round_reg[384]) );
  DFF \round_reg_reg[385]  ( .D(out[385]), .CLK(clk), .RST(rst), .I(in[385]), 
        .Q(round_reg[385]) );
  DFF \round_reg_reg[386]  ( .D(out[386]), .CLK(clk), .RST(rst), .I(in[386]), 
        .Q(round_reg[386]) );
  DFF \round_reg_reg[387]  ( .D(out[387]), .CLK(clk), .RST(rst), .I(in[387]), 
        .Q(round_reg[387]) );
  DFF \round_reg_reg[388]  ( .D(out[388]), .CLK(clk), .RST(rst), .I(in[388]), 
        .Q(round_reg[388]) );
  DFF \round_reg_reg[389]  ( .D(out[389]), .CLK(clk), .RST(rst), .I(in[389]), 
        .Q(round_reg[389]) );
  DFF \round_reg_reg[390]  ( .D(out[390]), .CLK(clk), .RST(rst), .I(in[390]), 
        .Q(round_reg[390]) );
  DFF \round_reg_reg[391]  ( .D(out[391]), .CLK(clk), .RST(rst), .I(in[391]), 
        .Q(round_reg[391]) );
  DFF \round_reg_reg[392]  ( .D(out[392]), .CLK(clk), .RST(rst), .I(in[392]), 
        .Q(round_reg[392]) );
  DFF \round_reg_reg[393]  ( .D(out[393]), .CLK(clk), .RST(rst), .I(in[393]), 
        .Q(round_reg[393]) );
  DFF \round_reg_reg[394]  ( .D(out[394]), .CLK(clk), .RST(rst), .I(in[394]), 
        .Q(round_reg[394]) );
  DFF \round_reg_reg[395]  ( .D(out[395]), .CLK(clk), .RST(rst), .I(in[395]), 
        .Q(round_reg[395]) );
  DFF \round_reg_reg[396]  ( .D(out[396]), .CLK(clk), .RST(rst), .I(in[396]), 
        .Q(round_reg[396]) );
  DFF \round_reg_reg[397]  ( .D(out[397]), .CLK(clk), .RST(rst), .I(in[397]), 
        .Q(round_reg[397]) );
  DFF \round_reg_reg[398]  ( .D(out[398]), .CLK(clk), .RST(rst), .I(in[398]), 
        .Q(round_reg[398]) );
  DFF \round_reg_reg[399]  ( .D(out[399]), .CLK(clk), .RST(rst), .I(in[399]), 
        .Q(round_reg[399]) );
  DFF \round_reg_reg[400]  ( .D(out[400]), .CLK(clk), .RST(rst), .I(in[400]), 
        .Q(round_reg[400]) );
  DFF \round_reg_reg[401]  ( .D(out[401]), .CLK(clk), .RST(rst), .I(in[401]), 
        .Q(round_reg[401]) );
  DFF \round_reg_reg[402]  ( .D(out[402]), .CLK(clk), .RST(rst), .I(in[402]), 
        .Q(round_reg[402]) );
  DFF \round_reg_reg[403]  ( .D(out[403]), .CLK(clk), .RST(rst), .I(in[403]), 
        .Q(round_reg[403]) );
  DFF \round_reg_reg[404]  ( .D(out[404]), .CLK(clk), .RST(rst), .I(in[404]), 
        .Q(round_reg[404]) );
  DFF \round_reg_reg[405]  ( .D(out[405]), .CLK(clk), .RST(rst), .I(in[405]), 
        .Q(round_reg[405]) );
  DFF \round_reg_reg[406]  ( .D(out[406]), .CLK(clk), .RST(rst), .I(in[406]), 
        .Q(round_reg[406]) );
  DFF \round_reg_reg[407]  ( .D(out[407]), .CLK(clk), .RST(rst), .I(in[407]), 
        .Q(round_reg[407]) );
  DFF \round_reg_reg[408]  ( .D(out[408]), .CLK(clk), .RST(rst), .I(in[408]), 
        .Q(round_reg[408]) );
  DFF \round_reg_reg[409]  ( .D(out[409]), .CLK(clk), .RST(rst), .I(in[409]), 
        .Q(round_reg[409]) );
  DFF \round_reg_reg[410]  ( .D(out[410]), .CLK(clk), .RST(rst), .I(in[410]), 
        .Q(round_reg[410]) );
  DFF \round_reg_reg[411]  ( .D(out[411]), .CLK(clk), .RST(rst), .I(in[411]), 
        .Q(round_reg[411]) );
  DFF \round_reg_reg[412]  ( .D(out[412]), .CLK(clk), .RST(rst), .I(in[412]), 
        .Q(round_reg[412]) );
  DFF \round_reg_reg[413]  ( .D(out[413]), .CLK(clk), .RST(rst), .I(in[413]), 
        .Q(round_reg[413]) );
  DFF \round_reg_reg[414]  ( .D(out[414]), .CLK(clk), .RST(rst), .I(in[414]), 
        .Q(round_reg[414]) );
  DFF \round_reg_reg[415]  ( .D(out[415]), .CLK(clk), .RST(rst), .I(in[415]), 
        .Q(round_reg[415]) );
  DFF \round_reg_reg[416]  ( .D(out[416]), .CLK(clk), .RST(rst), .I(in[416]), 
        .Q(round_reg[416]) );
  DFF \round_reg_reg[417]  ( .D(out[417]), .CLK(clk), .RST(rst), .I(in[417]), 
        .Q(round_reg[417]) );
  DFF \round_reg_reg[418]  ( .D(out[418]), .CLK(clk), .RST(rst), .I(in[418]), 
        .Q(round_reg[418]) );
  DFF \round_reg_reg[419]  ( .D(out[419]), .CLK(clk), .RST(rst), .I(in[419]), 
        .Q(round_reg[419]) );
  DFF \round_reg_reg[420]  ( .D(out[420]), .CLK(clk), .RST(rst), .I(in[420]), 
        .Q(round_reg[420]) );
  DFF \round_reg_reg[421]  ( .D(out[421]), .CLK(clk), .RST(rst), .I(in[421]), 
        .Q(round_reg[421]) );
  DFF \round_reg_reg[422]  ( .D(out[422]), .CLK(clk), .RST(rst), .I(in[422]), 
        .Q(round_reg[422]) );
  DFF \round_reg_reg[423]  ( .D(out[423]), .CLK(clk), .RST(rst), .I(in[423]), 
        .Q(round_reg[423]) );
  DFF \round_reg_reg[424]  ( .D(out[424]), .CLK(clk), .RST(rst), .I(in[424]), 
        .Q(round_reg[424]) );
  DFF \round_reg_reg[425]  ( .D(out[425]), .CLK(clk), .RST(rst), .I(in[425]), 
        .Q(round_reg[425]) );
  DFF \round_reg_reg[426]  ( .D(out[426]), .CLK(clk), .RST(rst), .I(in[426]), 
        .Q(round_reg[426]) );
  DFF \round_reg_reg[427]  ( .D(out[427]), .CLK(clk), .RST(rst), .I(in[427]), 
        .Q(round_reg[427]) );
  DFF \round_reg_reg[428]  ( .D(out[428]), .CLK(clk), .RST(rst), .I(in[428]), 
        .Q(round_reg[428]) );
  DFF \round_reg_reg[429]  ( .D(out[429]), .CLK(clk), .RST(rst), .I(in[429]), 
        .Q(round_reg[429]) );
  DFF \round_reg_reg[430]  ( .D(out[430]), .CLK(clk), .RST(rst), .I(in[430]), 
        .Q(round_reg[430]) );
  DFF \round_reg_reg[431]  ( .D(out[431]), .CLK(clk), .RST(rst), .I(in[431]), 
        .Q(round_reg[431]) );
  DFF \round_reg_reg[432]  ( .D(out[432]), .CLK(clk), .RST(rst), .I(in[432]), 
        .Q(round_reg[432]) );
  DFF \round_reg_reg[433]  ( .D(out[433]), .CLK(clk), .RST(rst), .I(in[433]), 
        .Q(round_reg[433]) );
  DFF \round_reg_reg[434]  ( .D(out[434]), .CLK(clk), .RST(rst), .I(in[434]), 
        .Q(round_reg[434]) );
  DFF \round_reg_reg[435]  ( .D(out[435]), .CLK(clk), .RST(rst), .I(in[435]), 
        .Q(round_reg[435]) );
  DFF \round_reg_reg[436]  ( .D(out[436]), .CLK(clk), .RST(rst), .I(in[436]), 
        .Q(round_reg[436]) );
  DFF \round_reg_reg[437]  ( .D(out[437]), .CLK(clk), .RST(rst), .I(in[437]), 
        .Q(round_reg[437]) );
  DFF \round_reg_reg[438]  ( .D(out[438]), .CLK(clk), .RST(rst), .I(in[438]), 
        .Q(round_reg[438]) );
  DFF \round_reg_reg[439]  ( .D(out[439]), .CLK(clk), .RST(rst), .I(in[439]), 
        .Q(round_reg[439]) );
  DFF \round_reg_reg[440]  ( .D(out[440]), .CLK(clk), .RST(rst), .I(in[440]), 
        .Q(round_reg[440]) );
  DFF \round_reg_reg[441]  ( .D(out[441]), .CLK(clk), .RST(rst), .I(in[441]), 
        .Q(round_reg[441]) );
  DFF \round_reg_reg[442]  ( .D(out[442]), .CLK(clk), .RST(rst), .I(in[442]), 
        .Q(round_reg[442]) );
  DFF \round_reg_reg[443]  ( .D(out[443]), .CLK(clk), .RST(rst), .I(in[443]), 
        .Q(round_reg[443]) );
  DFF \round_reg_reg[444]  ( .D(out[444]), .CLK(clk), .RST(rst), .I(in[444]), 
        .Q(round_reg[444]) );
  DFF \round_reg_reg[445]  ( .D(out[445]), .CLK(clk), .RST(rst), .I(in[445]), 
        .Q(round_reg[445]) );
  DFF \round_reg_reg[446]  ( .D(out[446]), .CLK(clk), .RST(rst), .I(in[446]), 
        .Q(round_reg[446]) );
  DFF \round_reg_reg[447]  ( .D(out[447]), .CLK(clk), .RST(rst), .I(in[447]), 
        .Q(round_reg[447]) );
  DFF \round_reg_reg[448]  ( .D(out[448]), .CLK(clk), .RST(rst), .I(in[448]), 
        .Q(round_reg[448]) );
  DFF \round_reg_reg[449]  ( .D(out[449]), .CLK(clk), .RST(rst), .I(in[449]), 
        .Q(round_reg[449]) );
  DFF \round_reg_reg[450]  ( .D(out[450]), .CLK(clk), .RST(rst), .I(in[450]), 
        .Q(round_reg[450]) );
  DFF \round_reg_reg[451]  ( .D(out[451]), .CLK(clk), .RST(rst), .I(in[451]), 
        .Q(round_reg[451]) );
  DFF \round_reg_reg[452]  ( .D(out[452]), .CLK(clk), .RST(rst), .I(in[452]), 
        .Q(round_reg[452]) );
  DFF \round_reg_reg[453]  ( .D(out[453]), .CLK(clk), .RST(rst), .I(in[453]), 
        .Q(round_reg[453]) );
  DFF \round_reg_reg[454]  ( .D(out[454]), .CLK(clk), .RST(rst), .I(in[454]), 
        .Q(round_reg[454]) );
  DFF \round_reg_reg[455]  ( .D(out[455]), .CLK(clk), .RST(rst), .I(in[455]), 
        .Q(round_reg[455]) );
  DFF \round_reg_reg[456]  ( .D(out[456]), .CLK(clk), .RST(rst), .I(in[456]), 
        .Q(round_reg[456]) );
  DFF \round_reg_reg[457]  ( .D(out[457]), .CLK(clk), .RST(rst), .I(in[457]), 
        .Q(round_reg[457]) );
  DFF \round_reg_reg[458]  ( .D(out[458]), .CLK(clk), .RST(rst), .I(in[458]), 
        .Q(round_reg[458]) );
  DFF \round_reg_reg[459]  ( .D(out[459]), .CLK(clk), .RST(rst), .I(in[459]), 
        .Q(round_reg[459]) );
  DFF \round_reg_reg[460]  ( .D(out[460]), .CLK(clk), .RST(rst), .I(in[460]), 
        .Q(round_reg[460]) );
  DFF \round_reg_reg[461]  ( .D(out[461]), .CLK(clk), .RST(rst), .I(in[461]), 
        .Q(round_reg[461]) );
  DFF \round_reg_reg[462]  ( .D(out[462]), .CLK(clk), .RST(rst), .I(in[462]), 
        .Q(round_reg[462]) );
  DFF \round_reg_reg[463]  ( .D(out[463]), .CLK(clk), .RST(rst), .I(in[463]), 
        .Q(round_reg[463]) );
  DFF \round_reg_reg[464]  ( .D(out[464]), .CLK(clk), .RST(rst), .I(in[464]), 
        .Q(round_reg[464]) );
  DFF \round_reg_reg[465]  ( .D(out[465]), .CLK(clk), .RST(rst), .I(in[465]), 
        .Q(round_reg[465]) );
  DFF \round_reg_reg[466]  ( .D(out[466]), .CLK(clk), .RST(rst), .I(in[466]), 
        .Q(round_reg[466]) );
  DFF \round_reg_reg[467]  ( .D(out[467]), .CLK(clk), .RST(rst), .I(in[467]), 
        .Q(round_reg[467]) );
  DFF \round_reg_reg[468]  ( .D(out[468]), .CLK(clk), .RST(rst), .I(in[468]), 
        .Q(round_reg[468]) );
  DFF \round_reg_reg[469]  ( .D(out[469]), .CLK(clk), .RST(rst), .I(in[469]), 
        .Q(round_reg[469]) );
  DFF \round_reg_reg[470]  ( .D(out[470]), .CLK(clk), .RST(rst), .I(in[470]), 
        .Q(round_reg[470]) );
  DFF \round_reg_reg[471]  ( .D(out[471]), .CLK(clk), .RST(rst), .I(in[471]), 
        .Q(round_reg[471]) );
  DFF \round_reg_reg[472]  ( .D(out[472]), .CLK(clk), .RST(rst), .I(in[472]), 
        .Q(round_reg[472]) );
  DFF \round_reg_reg[473]  ( .D(out[473]), .CLK(clk), .RST(rst), .I(in[473]), 
        .Q(round_reg[473]) );
  DFF \round_reg_reg[474]  ( .D(out[474]), .CLK(clk), .RST(rst), .I(in[474]), 
        .Q(round_reg[474]) );
  DFF \round_reg_reg[475]  ( .D(out[475]), .CLK(clk), .RST(rst), .I(in[475]), 
        .Q(round_reg[475]) );
  DFF \round_reg_reg[476]  ( .D(out[476]), .CLK(clk), .RST(rst), .I(in[476]), 
        .Q(round_reg[476]) );
  DFF \round_reg_reg[477]  ( .D(out[477]), .CLK(clk), .RST(rst), .I(in[477]), 
        .Q(round_reg[477]) );
  DFF \round_reg_reg[478]  ( .D(out[478]), .CLK(clk), .RST(rst), .I(in[478]), 
        .Q(round_reg[478]) );
  DFF \round_reg_reg[479]  ( .D(out[479]), .CLK(clk), .RST(rst), .I(in[479]), 
        .Q(round_reg[479]) );
  DFF \round_reg_reg[480]  ( .D(out[480]), .CLK(clk), .RST(rst), .I(in[480]), 
        .Q(round_reg[480]) );
  DFF \round_reg_reg[481]  ( .D(out[481]), .CLK(clk), .RST(rst), .I(in[481]), 
        .Q(round_reg[481]) );
  DFF \round_reg_reg[482]  ( .D(out[482]), .CLK(clk), .RST(rst), .I(in[482]), 
        .Q(round_reg[482]) );
  DFF \round_reg_reg[483]  ( .D(out[483]), .CLK(clk), .RST(rst), .I(in[483]), 
        .Q(round_reg[483]) );
  DFF \round_reg_reg[484]  ( .D(out[484]), .CLK(clk), .RST(rst), .I(in[484]), 
        .Q(round_reg[484]) );
  DFF \round_reg_reg[485]  ( .D(out[485]), .CLK(clk), .RST(rst), .I(in[485]), 
        .Q(round_reg[485]) );
  DFF \round_reg_reg[486]  ( .D(out[486]), .CLK(clk), .RST(rst), .I(in[486]), 
        .Q(round_reg[486]) );
  DFF \round_reg_reg[487]  ( .D(out[487]), .CLK(clk), .RST(rst), .I(in[487]), 
        .Q(round_reg[487]) );
  DFF \round_reg_reg[488]  ( .D(out[488]), .CLK(clk), .RST(rst), .I(in[488]), 
        .Q(round_reg[488]) );
  DFF \round_reg_reg[489]  ( .D(out[489]), .CLK(clk), .RST(rst), .I(in[489]), 
        .Q(round_reg[489]) );
  DFF \round_reg_reg[490]  ( .D(out[490]), .CLK(clk), .RST(rst), .I(in[490]), 
        .Q(round_reg[490]) );
  DFF \round_reg_reg[491]  ( .D(out[491]), .CLK(clk), .RST(rst), .I(in[491]), 
        .Q(round_reg[491]) );
  DFF \round_reg_reg[492]  ( .D(out[492]), .CLK(clk), .RST(rst), .I(in[492]), 
        .Q(round_reg[492]) );
  DFF \round_reg_reg[493]  ( .D(out[493]), .CLK(clk), .RST(rst), .I(in[493]), 
        .Q(round_reg[493]) );
  DFF \round_reg_reg[494]  ( .D(out[494]), .CLK(clk), .RST(rst), .I(in[494]), 
        .Q(round_reg[494]) );
  DFF \round_reg_reg[495]  ( .D(out[495]), .CLK(clk), .RST(rst), .I(in[495]), 
        .Q(round_reg[495]) );
  DFF \round_reg_reg[496]  ( .D(out[496]), .CLK(clk), .RST(rst), .I(in[496]), 
        .Q(round_reg[496]) );
  DFF \round_reg_reg[497]  ( .D(out[497]), .CLK(clk), .RST(rst), .I(in[497]), 
        .Q(round_reg[497]) );
  DFF \round_reg_reg[498]  ( .D(out[498]), .CLK(clk), .RST(rst), .I(in[498]), 
        .Q(round_reg[498]) );
  DFF \round_reg_reg[499]  ( .D(out[499]), .CLK(clk), .RST(rst), .I(in[499]), 
        .Q(round_reg[499]) );
  DFF \round_reg_reg[500]  ( .D(out[500]), .CLK(clk), .RST(rst), .I(in[500]), 
        .Q(round_reg[500]) );
  DFF \round_reg_reg[501]  ( .D(out[501]), .CLK(clk), .RST(rst), .I(in[501]), 
        .Q(round_reg[501]) );
  DFF \round_reg_reg[502]  ( .D(out[502]), .CLK(clk), .RST(rst), .I(in[502]), 
        .Q(round_reg[502]) );
  DFF \round_reg_reg[503]  ( .D(out[503]), .CLK(clk), .RST(rst), .I(in[503]), 
        .Q(round_reg[503]) );
  DFF \round_reg_reg[504]  ( .D(out[504]), .CLK(clk), .RST(rst), .I(in[504]), 
        .Q(round_reg[504]) );
  DFF \round_reg_reg[505]  ( .D(out[505]), .CLK(clk), .RST(rst), .I(in[505]), 
        .Q(round_reg[505]) );
  DFF \round_reg_reg[506]  ( .D(out[506]), .CLK(clk), .RST(rst), .I(in[506]), 
        .Q(round_reg[506]) );
  DFF \round_reg_reg[507]  ( .D(out[507]), .CLK(clk), .RST(rst), .I(in[507]), 
        .Q(round_reg[507]) );
  DFF \round_reg_reg[508]  ( .D(out[508]), .CLK(clk), .RST(rst), .I(in[508]), 
        .Q(round_reg[508]) );
  DFF \round_reg_reg[509]  ( .D(out[509]), .CLK(clk), .RST(rst), .I(in[509]), 
        .Q(round_reg[509]) );
  DFF \round_reg_reg[510]  ( .D(out[510]), .CLK(clk), .RST(rst), .I(in[510]), 
        .Q(round_reg[510]) );
  DFF \round_reg_reg[511]  ( .D(out[511]), .CLK(clk), .RST(rst), .I(in[511]), 
        .Q(round_reg[511]) );
  DFF \round_reg_reg[512]  ( .D(out[512]), .CLK(clk), .RST(rst), .I(in[512]), 
        .Q(round_reg[512]) );
  DFF \round_reg_reg[513]  ( .D(out[513]), .CLK(clk), .RST(rst), .I(in[513]), 
        .Q(round_reg[513]) );
  DFF \round_reg_reg[514]  ( .D(out[514]), .CLK(clk), .RST(rst), .I(in[514]), 
        .Q(round_reg[514]) );
  DFF \round_reg_reg[515]  ( .D(out[515]), .CLK(clk), .RST(rst), .I(in[515]), 
        .Q(round_reg[515]) );
  DFF \round_reg_reg[516]  ( .D(out[516]), .CLK(clk), .RST(rst), .I(in[516]), 
        .Q(round_reg[516]) );
  DFF \round_reg_reg[517]  ( .D(out[517]), .CLK(clk), .RST(rst), .I(in[517]), 
        .Q(round_reg[517]) );
  DFF \round_reg_reg[518]  ( .D(out[518]), .CLK(clk), .RST(rst), .I(in[518]), 
        .Q(round_reg[518]) );
  DFF \round_reg_reg[519]  ( .D(out[519]), .CLK(clk), .RST(rst), .I(in[519]), 
        .Q(round_reg[519]) );
  DFF \round_reg_reg[520]  ( .D(out[520]), .CLK(clk), .RST(rst), .I(in[520]), 
        .Q(round_reg[520]) );
  DFF \round_reg_reg[521]  ( .D(out[521]), .CLK(clk), .RST(rst), .I(in[521]), 
        .Q(round_reg[521]) );
  DFF \round_reg_reg[522]  ( .D(out[522]), .CLK(clk), .RST(rst), .I(in[522]), 
        .Q(round_reg[522]) );
  DFF \round_reg_reg[523]  ( .D(out[523]), .CLK(clk), .RST(rst), .I(in[523]), 
        .Q(round_reg[523]) );
  DFF \round_reg_reg[524]  ( .D(out[524]), .CLK(clk), .RST(rst), .I(in[524]), 
        .Q(round_reg[524]) );
  DFF \round_reg_reg[525]  ( .D(out[525]), .CLK(clk), .RST(rst), .I(in[525]), 
        .Q(round_reg[525]) );
  DFF \round_reg_reg[526]  ( .D(out[526]), .CLK(clk), .RST(rst), .I(in[526]), 
        .Q(round_reg[526]) );
  DFF \round_reg_reg[527]  ( .D(out[527]), .CLK(clk), .RST(rst), .I(in[527]), 
        .Q(round_reg[527]) );
  DFF \round_reg_reg[528]  ( .D(out[528]), .CLK(clk), .RST(rst), .I(in[528]), 
        .Q(round_reg[528]) );
  DFF \round_reg_reg[529]  ( .D(out[529]), .CLK(clk), .RST(rst), .I(in[529]), 
        .Q(round_reg[529]) );
  DFF \round_reg_reg[530]  ( .D(out[530]), .CLK(clk), .RST(rst), .I(in[530]), 
        .Q(round_reg[530]) );
  DFF \round_reg_reg[531]  ( .D(out[531]), .CLK(clk), .RST(rst), .I(in[531]), 
        .Q(round_reg[531]) );
  DFF \round_reg_reg[532]  ( .D(out[532]), .CLK(clk), .RST(rst), .I(in[532]), 
        .Q(round_reg[532]) );
  DFF \round_reg_reg[533]  ( .D(out[533]), .CLK(clk), .RST(rst), .I(in[533]), 
        .Q(round_reg[533]) );
  DFF \round_reg_reg[534]  ( .D(out[534]), .CLK(clk), .RST(rst), .I(in[534]), 
        .Q(round_reg[534]) );
  DFF \round_reg_reg[535]  ( .D(out[535]), .CLK(clk), .RST(rst), .I(in[535]), 
        .Q(round_reg[535]) );
  DFF \round_reg_reg[536]  ( .D(out[536]), .CLK(clk), .RST(rst), .I(in[536]), 
        .Q(round_reg[536]) );
  DFF \round_reg_reg[537]  ( .D(out[537]), .CLK(clk), .RST(rst), .I(in[537]), 
        .Q(round_reg[537]) );
  DFF \round_reg_reg[538]  ( .D(out[538]), .CLK(clk), .RST(rst), .I(in[538]), 
        .Q(round_reg[538]) );
  DFF \round_reg_reg[539]  ( .D(out[539]), .CLK(clk), .RST(rst), .I(in[539]), 
        .Q(round_reg[539]) );
  DFF \round_reg_reg[540]  ( .D(out[540]), .CLK(clk), .RST(rst), .I(in[540]), 
        .Q(round_reg[540]) );
  DFF \round_reg_reg[541]  ( .D(out[541]), .CLK(clk), .RST(rst), .I(in[541]), 
        .Q(round_reg[541]) );
  DFF \round_reg_reg[542]  ( .D(out[542]), .CLK(clk), .RST(rst), .I(in[542]), 
        .Q(round_reg[542]) );
  DFF \round_reg_reg[543]  ( .D(out[543]), .CLK(clk), .RST(rst), .I(in[543]), 
        .Q(round_reg[543]) );
  DFF \round_reg_reg[544]  ( .D(out[544]), .CLK(clk), .RST(rst), .I(in[544]), 
        .Q(round_reg[544]) );
  DFF \round_reg_reg[545]  ( .D(out[545]), .CLK(clk), .RST(rst), .I(in[545]), 
        .Q(round_reg[545]) );
  DFF \round_reg_reg[546]  ( .D(out[546]), .CLK(clk), .RST(rst), .I(in[546]), 
        .Q(round_reg[546]) );
  DFF \round_reg_reg[547]  ( .D(out[547]), .CLK(clk), .RST(rst), .I(in[547]), 
        .Q(round_reg[547]) );
  DFF \round_reg_reg[548]  ( .D(out[548]), .CLK(clk), .RST(rst), .I(in[548]), 
        .Q(round_reg[548]) );
  DFF \round_reg_reg[549]  ( .D(out[549]), .CLK(clk), .RST(rst), .I(in[549]), 
        .Q(round_reg[549]) );
  DFF \round_reg_reg[550]  ( .D(out[550]), .CLK(clk), .RST(rst), .I(in[550]), 
        .Q(round_reg[550]) );
  DFF \round_reg_reg[551]  ( .D(out[551]), .CLK(clk), .RST(rst), .I(in[551]), 
        .Q(round_reg[551]) );
  DFF \round_reg_reg[552]  ( .D(out[552]), .CLK(clk), .RST(rst), .I(in[552]), 
        .Q(round_reg[552]) );
  DFF \round_reg_reg[553]  ( .D(out[553]), .CLK(clk), .RST(rst), .I(in[553]), 
        .Q(round_reg[553]) );
  DFF \round_reg_reg[554]  ( .D(out[554]), .CLK(clk), .RST(rst), .I(in[554]), 
        .Q(round_reg[554]) );
  DFF \round_reg_reg[555]  ( .D(out[555]), .CLK(clk), .RST(rst), .I(in[555]), 
        .Q(round_reg[555]) );
  DFF \round_reg_reg[556]  ( .D(out[556]), .CLK(clk), .RST(rst), .I(in[556]), 
        .Q(round_reg[556]) );
  DFF \round_reg_reg[557]  ( .D(out[557]), .CLK(clk), .RST(rst), .I(in[557]), 
        .Q(round_reg[557]) );
  DFF \round_reg_reg[558]  ( .D(out[558]), .CLK(clk), .RST(rst), .I(in[558]), 
        .Q(round_reg[558]) );
  DFF \round_reg_reg[559]  ( .D(out[559]), .CLK(clk), .RST(rst), .I(in[559]), 
        .Q(round_reg[559]) );
  DFF \round_reg_reg[560]  ( .D(out[560]), .CLK(clk), .RST(rst), .I(in[560]), 
        .Q(round_reg[560]) );
  DFF \round_reg_reg[561]  ( .D(out[561]), .CLK(clk), .RST(rst), .I(in[561]), 
        .Q(round_reg[561]) );
  DFF \round_reg_reg[562]  ( .D(out[562]), .CLK(clk), .RST(rst), .I(in[562]), 
        .Q(round_reg[562]) );
  DFF \round_reg_reg[563]  ( .D(out[563]), .CLK(clk), .RST(rst), .I(in[563]), 
        .Q(round_reg[563]) );
  DFF \round_reg_reg[564]  ( .D(out[564]), .CLK(clk), .RST(rst), .I(in[564]), 
        .Q(round_reg[564]) );
  DFF \round_reg_reg[565]  ( .D(out[565]), .CLK(clk), .RST(rst), .I(in[565]), 
        .Q(round_reg[565]) );
  DFF \round_reg_reg[566]  ( .D(out[566]), .CLK(clk), .RST(rst), .I(in[566]), 
        .Q(round_reg[566]) );
  DFF \round_reg_reg[567]  ( .D(out[567]), .CLK(clk), .RST(rst), .I(in[567]), 
        .Q(round_reg[567]) );
  DFF \round_reg_reg[568]  ( .D(out[568]), .CLK(clk), .RST(rst), .I(in[568]), 
        .Q(round_reg[568]) );
  DFF \round_reg_reg[569]  ( .D(out[569]), .CLK(clk), .RST(rst), .I(in[569]), 
        .Q(round_reg[569]) );
  DFF \round_reg_reg[570]  ( .D(out[570]), .CLK(clk), .RST(rst), .I(in[570]), 
        .Q(round_reg[570]) );
  DFF \round_reg_reg[571]  ( .D(out[571]), .CLK(clk), .RST(rst), .I(in[571]), 
        .Q(round_reg[571]) );
  DFF \round_reg_reg[572]  ( .D(out[572]), .CLK(clk), .RST(rst), .I(in[572]), 
        .Q(round_reg[572]) );
  DFF \round_reg_reg[573]  ( .D(out[573]), .CLK(clk), .RST(rst), .I(in[573]), 
        .Q(round_reg[573]) );
  DFF \round_reg_reg[574]  ( .D(out[574]), .CLK(clk), .RST(rst), .I(in[574]), 
        .Q(round_reg[574]) );
  DFF \round_reg_reg[575]  ( .D(out[575]), .CLK(clk), .RST(rst), .I(in[575]), 
        .Q(round_reg[575]) );
  DFF \round_reg_reg[576]  ( .D(out[576]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[576]) );
  DFF \round_reg_reg[577]  ( .D(out[577]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[577]) );
  DFF \round_reg_reg[578]  ( .D(out[578]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[578]) );
  DFF \round_reg_reg[579]  ( .D(out[579]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[579]) );
  DFF \round_reg_reg[580]  ( .D(out[580]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[580]) );
  DFF \round_reg_reg[581]  ( .D(out[581]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[581]) );
  DFF \round_reg_reg[582]  ( .D(out[582]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[582]) );
  DFF \round_reg_reg[583]  ( .D(out[583]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[583]) );
  DFF \round_reg_reg[584]  ( .D(out[584]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[584]) );
  DFF \round_reg_reg[585]  ( .D(out[585]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[585]) );
  DFF \round_reg_reg[586]  ( .D(out[586]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[586]) );
  DFF \round_reg_reg[587]  ( .D(out[587]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[587]) );
  DFF \round_reg_reg[588]  ( .D(out[588]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[588]) );
  DFF \round_reg_reg[589]  ( .D(out[589]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[589]) );
  DFF \round_reg_reg[590]  ( .D(out[590]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[590]) );
  DFF \round_reg_reg[591]  ( .D(out[591]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[591]) );
  DFF \round_reg_reg[592]  ( .D(out[592]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[592]) );
  DFF \round_reg_reg[593]  ( .D(out[593]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[593]) );
  DFF \round_reg_reg[594]  ( .D(out[594]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[594]) );
  DFF \round_reg_reg[595]  ( .D(out[595]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[595]) );
  DFF \round_reg_reg[596]  ( .D(out[596]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[596]) );
  DFF \round_reg_reg[597]  ( .D(out[597]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[597]) );
  DFF \round_reg_reg[598]  ( .D(out[598]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[598]) );
  DFF \round_reg_reg[599]  ( .D(out[599]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[599]) );
  DFF \round_reg_reg[600]  ( .D(out[600]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[600]) );
  DFF \round_reg_reg[601]  ( .D(out[601]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[601]) );
  DFF \round_reg_reg[602]  ( .D(out[602]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[602]) );
  DFF \round_reg_reg[603]  ( .D(out[603]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[603]) );
  DFF \round_reg_reg[604]  ( .D(out[604]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[604]) );
  DFF \round_reg_reg[605]  ( .D(out[605]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[605]) );
  DFF \round_reg_reg[606]  ( .D(out[606]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[606]) );
  DFF \round_reg_reg[607]  ( .D(out[607]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[607]) );
  DFF \round_reg_reg[608]  ( .D(out[608]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[608]) );
  DFF \round_reg_reg[609]  ( .D(out[609]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[609]) );
  DFF \round_reg_reg[610]  ( .D(out[610]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[610]) );
  DFF \round_reg_reg[611]  ( .D(out[611]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[611]) );
  DFF \round_reg_reg[612]  ( .D(out[612]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[612]) );
  DFF \round_reg_reg[613]  ( .D(out[613]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[613]) );
  DFF \round_reg_reg[614]  ( .D(out[614]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[614]) );
  DFF \round_reg_reg[615]  ( .D(out[615]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[615]) );
  DFF \round_reg_reg[616]  ( .D(out[616]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[616]) );
  DFF \round_reg_reg[617]  ( .D(out[617]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[617]) );
  DFF \round_reg_reg[618]  ( .D(out[618]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[618]) );
  DFF \round_reg_reg[619]  ( .D(out[619]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[619]) );
  DFF \round_reg_reg[620]  ( .D(out[620]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[620]) );
  DFF \round_reg_reg[621]  ( .D(out[621]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[621]) );
  DFF \round_reg_reg[622]  ( .D(out[622]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[622]) );
  DFF \round_reg_reg[623]  ( .D(out[623]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[623]) );
  DFF \round_reg_reg[624]  ( .D(out[624]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[624]) );
  DFF \round_reg_reg[625]  ( .D(out[625]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[625]) );
  DFF \round_reg_reg[626]  ( .D(out[626]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[626]) );
  DFF \round_reg_reg[627]  ( .D(out[627]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[627]) );
  DFF \round_reg_reg[628]  ( .D(out[628]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[628]) );
  DFF \round_reg_reg[629]  ( .D(out[629]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[629]) );
  DFF \round_reg_reg[630]  ( .D(out[630]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[630]) );
  DFF \round_reg_reg[631]  ( .D(out[631]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[631]) );
  DFF \round_reg_reg[632]  ( .D(out[632]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[632]) );
  DFF \round_reg_reg[633]  ( .D(out[633]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[633]) );
  DFF \round_reg_reg[634]  ( .D(out[634]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[634]) );
  DFF \round_reg_reg[635]  ( .D(out[635]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[635]) );
  DFF \round_reg_reg[636]  ( .D(out[636]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[636]) );
  DFF \round_reg_reg[637]  ( .D(out[637]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[637]) );
  DFF \round_reg_reg[638]  ( .D(out[638]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[638]) );
  DFF \round_reg_reg[639]  ( .D(out[639]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[639]) );
  DFF \round_reg_reg[640]  ( .D(out[640]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[640]) );
  DFF \round_reg_reg[641]  ( .D(out[641]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[641]) );
  DFF \round_reg_reg[642]  ( .D(out[642]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[642]) );
  DFF \round_reg_reg[643]  ( .D(out[643]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[643]) );
  DFF \round_reg_reg[644]  ( .D(out[644]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[644]) );
  DFF \round_reg_reg[645]  ( .D(out[645]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[645]) );
  DFF \round_reg_reg[646]  ( .D(out[646]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[646]) );
  DFF \round_reg_reg[647]  ( .D(out[647]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[647]) );
  DFF \round_reg_reg[648]  ( .D(out[648]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[648]) );
  DFF \round_reg_reg[649]  ( .D(out[649]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[649]) );
  DFF \round_reg_reg[650]  ( .D(out[650]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[650]) );
  DFF \round_reg_reg[651]  ( .D(out[651]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[651]) );
  DFF \round_reg_reg[652]  ( .D(out[652]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[652]) );
  DFF \round_reg_reg[653]  ( .D(out[653]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[653]) );
  DFF \round_reg_reg[654]  ( .D(out[654]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[654]) );
  DFF \round_reg_reg[655]  ( .D(out[655]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[655]) );
  DFF \round_reg_reg[656]  ( .D(out[656]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[656]) );
  DFF \round_reg_reg[657]  ( .D(out[657]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[657]) );
  DFF \round_reg_reg[658]  ( .D(out[658]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[658]) );
  DFF \round_reg_reg[659]  ( .D(out[659]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[659]) );
  DFF \round_reg_reg[660]  ( .D(out[660]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[660]) );
  DFF \round_reg_reg[661]  ( .D(out[661]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[661]) );
  DFF \round_reg_reg[662]  ( .D(out[662]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[662]) );
  DFF \round_reg_reg[663]  ( .D(out[663]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[663]) );
  DFF \round_reg_reg[664]  ( .D(out[664]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[664]) );
  DFF \round_reg_reg[665]  ( .D(out[665]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[665]) );
  DFF \round_reg_reg[666]  ( .D(out[666]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[666]) );
  DFF \round_reg_reg[667]  ( .D(out[667]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[667]) );
  DFF \round_reg_reg[668]  ( .D(out[668]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[668]) );
  DFF \round_reg_reg[669]  ( .D(out[669]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[669]) );
  DFF \round_reg_reg[670]  ( .D(out[670]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[670]) );
  DFF \round_reg_reg[671]  ( .D(out[671]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[671]) );
  DFF \round_reg_reg[672]  ( .D(out[672]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[672]) );
  DFF \round_reg_reg[673]  ( .D(out[673]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[673]) );
  DFF \round_reg_reg[674]  ( .D(out[674]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[674]) );
  DFF \round_reg_reg[675]  ( .D(out[675]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[675]) );
  DFF \round_reg_reg[676]  ( .D(out[676]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[676]) );
  DFF \round_reg_reg[677]  ( .D(out[677]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[677]) );
  DFF \round_reg_reg[678]  ( .D(out[678]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[678]) );
  DFF \round_reg_reg[679]  ( .D(out[679]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[679]) );
  DFF \round_reg_reg[680]  ( .D(out[680]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[680]) );
  DFF \round_reg_reg[681]  ( .D(out[681]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[681]) );
  DFF \round_reg_reg[682]  ( .D(out[682]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[682]) );
  DFF \round_reg_reg[683]  ( .D(out[683]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[683]) );
  DFF \round_reg_reg[684]  ( .D(out[684]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[684]) );
  DFF \round_reg_reg[685]  ( .D(out[685]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[685]) );
  DFF \round_reg_reg[686]  ( .D(out[686]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[686]) );
  DFF \round_reg_reg[687]  ( .D(out[687]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[687]) );
  DFF \round_reg_reg[688]  ( .D(out[688]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[688]) );
  DFF \round_reg_reg[689]  ( .D(out[689]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[689]) );
  DFF \round_reg_reg[690]  ( .D(out[690]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[690]) );
  DFF \round_reg_reg[691]  ( .D(out[691]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[691]) );
  DFF \round_reg_reg[692]  ( .D(out[692]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[692]) );
  DFF \round_reg_reg[693]  ( .D(out[693]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[693]) );
  DFF \round_reg_reg[694]  ( .D(out[694]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[694]) );
  DFF \round_reg_reg[695]  ( .D(out[695]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[695]) );
  DFF \round_reg_reg[696]  ( .D(out[696]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[696]) );
  DFF \round_reg_reg[697]  ( .D(out[697]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[697]) );
  DFF \round_reg_reg[698]  ( .D(out[698]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[698]) );
  DFF \round_reg_reg[699]  ( .D(out[699]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[699]) );
  DFF \round_reg_reg[700]  ( .D(out[700]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[700]) );
  DFF \round_reg_reg[701]  ( .D(out[701]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[701]) );
  DFF \round_reg_reg[702]  ( .D(out[702]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[702]) );
  DFF \round_reg_reg[703]  ( .D(out[703]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[703]) );
  DFF \round_reg_reg[704]  ( .D(out[704]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[704]) );
  DFF \round_reg_reg[705]  ( .D(out[705]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[705]) );
  DFF \round_reg_reg[706]  ( .D(out[706]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[706]) );
  DFF \round_reg_reg[707]  ( .D(out[707]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[707]) );
  DFF \round_reg_reg[708]  ( .D(out[708]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[708]) );
  DFF \round_reg_reg[709]  ( .D(out[709]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[709]) );
  DFF \round_reg_reg[710]  ( .D(out[710]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[710]) );
  DFF \round_reg_reg[711]  ( .D(out[711]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[711]) );
  DFF \round_reg_reg[712]  ( .D(out[712]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[712]) );
  DFF \round_reg_reg[713]  ( .D(out[713]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[713]) );
  DFF \round_reg_reg[714]  ( .D(out[714]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[714]) );
  DFF \round_reg_reg[715]  ( .D(out[715]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[715]) );
  DFF \round_reg_reg[716]  ( .D(out[716]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[716]) );
  DFF \round_reg_reg[717]  ( .D(out[717]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[717]) );
  DFF \round_reg_reg[718]  ( .D(out[718]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[718]) );
  DFF \round_reg_reg[719]  ( .D(out[719]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[719]) );
  DFF \round_reg_reg[720]  ( .D(out[720]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[720]) );
  DFF \round_reg_reg[721]  ( .D(out[721]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[721]) );
  DFF \round_reg_reg[722]  ( .D(out[722]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[722]) );
  DFF \round_reg_reg[723]  ( .D(out[723]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[723]) );
  DFF \round_reg_reg[724]  ( .D(out[724]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[724]) );
  DFF \round_reg_reg[725]  ( .D(out[725]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[725]) );
  DFF \round_reg_reg[726]  ( .D(out[726]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[726]) );
  DFF \round_reg_reg[727]  ( .D(out[727]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[727]) );
  DFF \round_reg_reg[728]  ( .D(out[728]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[728]) );
  DFF \round_reg_reg[729]  ( .D(out[729]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[729]) );
  DFF \round_reg_reg[730]  ( .D(out[730]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[730]) );
  DFF \round_reg_reg[731]  ( .D(out[731]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[731]) );
  DFF \round_reg_reg[732]  ( .D(out[732]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[732]) );
  DFF \round_reg_reg[733]  ( .D(out[733]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[733]) );
  DFF \round_reg_reg[734]  ( .D(out[734]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[734]) );
  DFF \round_reg_reg[735]  ( .D(out[735]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[735]) );
  DFF \round_reg_reg[736]  ( .D(out[736]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[736]) );
  DFF \round_reg_reg[737]  ( .D(out[737]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[737]) );
  DFF \round_reg_reg[738]  ( .D(out[738]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[738]) );
  DFF \round_reg_reg[739]  ( .D(out[739]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[739]) );
  DFF \round_reg_reg[740]  ( .D(out[740]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[740]) );
  DFF \round_reg_reg[741]  ( .D(out[741]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[741]) );
  DFF \round_reg_reg[742]  ( .D(out[742]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[742]) );
  DFF \round_reg_reg[743]  ( .D(out[743]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[743]) );
  DFF \round_reg_reg[744]  ( .D(out[744]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[744]) );
  DFF \round_reg_reg[745]  ( .D(out[745]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[745]) );
  DFF \round_reg_reg[746]  ( .D(out[746]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[746]) );
  DFF \round_reg_reg[747]  ( .D(out[747]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[747]) );
  DFF \round_reg_reg[748]  ( .D(out[748]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[748]) );
  DFF \round_reg_reg[749]  ( .D(out[749]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[749]) );
  DFF \round_reg_reg[750]  ( .D(out[750]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[750]) );
  DFF \round_reg_reg[751]  ( .D(out[751]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[751]) );
  DFF \round_reg_reg[752]  ( .D(out[752]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[752]) );
  DFF \round_reg_reg[753]  ( .D(out[753]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[753]) );
  DFF \round_reg_reg[754]  ( .D(out[754]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[754]) );
  DFF \round_reg_reg[755]  ( .D(out[755]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[755]) );
  DFF \round_reg_reg[756]  ( .D(out[756]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[756]) );
  DFF \round_reg_reg[757]  ( .D(out[757]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[757]) );
  DFF \round_reg_reg[758]  ( .D(out[758]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[758]) );
  DFF \round_reg_reg[759]  ( .D(out[759]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[759]) );
  DFF \round_reg_reg[760]  ( .D(out[760]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[760]) );
  DFF \round_reg_reg[761]  ( .D(out[761]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[761]) );
  DFF \round_reg_reg[762]  ( .D(out[762]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[762]) );
  DFF \round_reg_reg[763]  ( .D(out[763]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[763]) );
  DFF \round_reg_reg[764]  ( .D(out[764]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[764]) );
  DFF \round_reg_reg[765]  ( .D(out[765]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[765]) );
  DFF \round_reg_reg[766]  ( .D(out[766]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[766]) );
  DFF \round_reg_reg[767]  ( .D(out[767]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[767]) );
  DFF \round_reg_reg[768]  ( .D(out[768]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[768]) );
  DFF \round_reg_reg[769]  ( .D(out[769]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[769]) );
  DFF \round_reg_reg[770]  ( .D(out[770]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[770]) );
  DFF \round_reg_reg[771]  ( .D(out[771]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[771]) );
  DFF \round_reg_reg[772]  ( .D(out[772]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[772]) );
  DFF \round_reg_reg[773]  ( .D(out[773]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[773]) );
  DFF \round_reg_reg[774]  ( .D(out[774]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[774]) );
  DFF \round_reg_reg[775]  ( .D(out[775]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[775]) );
  DFF \round_reg_reg[776]  ( .D(out[776]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[776]) );
  DFF \round_reg_reg[777]  ( .D(out[777]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[777]) );
  DFF \round_reg_reg[778]  ( .D(out[778]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[778]) );
  DFF \round_reg_reg[779]  ( .D(out[779]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[779]) );
  DFF \round_reg_reg[780]  ( .D(out[780]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[780]) );
  DFF \round_reg_reg[781]  ( .D(out[781]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[781]) );
  DFF \round_reg_reg[782]  ( .D(out[782]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[782]) );
  DFF \round_reg_reg[783]  ( .D(out[783]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[783]) );
  DFF \round_reg_reg[784]  ( .D(out[784]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[784]) );
  DFF \round_reg_reg[785]  ( .D(out[785]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[785]) );
  DFF \round_reg_reg[786]  ( .D(out[786]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[786]) );
  DFF \round_reg_reg[787]  ( .D(out[787]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[787]) );
  DFF \round_reg_reg[788]  ( .D(out[788]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[788]) );
  DFF \round_reg_reg[789]  ( .D(out[789]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[789]) );
  DFF \round_reg_reg[790]  ( .D(out[790]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[790]) );
  DFF \round_reg_reg[791]  ( .D(out[791]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[791]) );
  DFF \round_reg_reg[792]  ( .D(out[792]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[792]) );
  DFF \round_reg_reg[793]  ( .D(out[793]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[793]) );
  DFF \round_reg_reg[794]  ( .D(out[794]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[794]) );
  DFF \round_reg_reg[795]  ( .D(out[795]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[795]) );
  DFF \round_reg_reg[796]  ( .D(out[796]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[796]) );
  DFF \round_reg_reg[797]  ( .D(out[797]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[797]) );
  DFF \round_reg_reg[798]  ( .D(out[798]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[798]) );
  DFF \round_reg_reg[799]  ( .D(out[799]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[799]) );
  DFF \round_reg_reg[800]  ( .D(out[800]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[800]) );
  DFF \round_reg_reg[801]  ( .D(out[801]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[801]) );
  DFF \round_reg_reg[802]  ( .D(out[802]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[802]) );
  DFF \round_reg_reg[803]  ( .D(out[803]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[803]) );
  DFF \round_reg_reg[804]  ( .D(out[804]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[804]) );
  DFF \round_reg_reg[805]  ( .D(out[805]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[805]) );
  DFF \round_reg_reg[806]  ( .D(out[806]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[806]) );
  DFF \round_reg_reg[807]  ( .D(out[807]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[807]) );
  DFF \round_reg_reg[808]  ( .D(out[808]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[808]) );
  DFF \round_reg_reg[809]  ( .D(out[809]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[809]) );
  DFF \round_reg_reg[810]  ( .D(out[810]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[810]) );
  DFF \round_reg_reg[811]  ( .D(out[811]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[811]) );
  DFF \round_reg_reg[812]  ( .D(out[812]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[812]) );
  DFF \round_reg_reg[813]  ( .D(out[813]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[813]) );
  DFF \round_reg_reg[814]  ( .D(out[814]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[814]) );
  DFF \round_reg_reg[815]  ( .D(out[815]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[815]) );
  DFF \round_reg_reg[816]  ( .D(out[816]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[816]) );
  DFF \round_reg_reg[817]  ( .D(out[817]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[817]) );
  DFF \round_reg_reg[818]  ( .D(out[818]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[818]) );
  DFF \round_reg_reg[819]  ( .D(out[819]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[819]) );
  DFF \round_reg_reg[820]  ( .D(out[820]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[820]) );
  DFF \round_reg_reg[821]  ( .D(out[821]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[821]) );
  DFF \round_reg_reg[822]  ( .D(out[822]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[822]) );
  DFF \round_reg_reg[823]  ( .D(out[823]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[823]) );
  DFF \round_reg_reg[824]  ( .D(out[824]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[824]) );
  DFF \round_reg_reg[825]  ( .D(out[825]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[825]) );
  DFF \round_reg_reg[826]  ( .D(out[826]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[826]) );
  DFF \round_reg_reg[827]  ( .D(out[827]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[827]) );
  DFF \round_reg_reg[828]  ( .D(out[828]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[828]) );
  DFF \round_reg_reg[829]  ( .D(out[829]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[829]) );
  DFF \round_reg_reg[830]  ( .D(out[830]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[830]) );
  DFF \round_reg_reg[831]  ( .D(out[831]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[831]) );
  DFF \round_reg_reg[832]  ( .D(out[832]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[832]) );
  DFF \round_reg_reg[833]  ( .D(out[833]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[833]) );
  DFF \round_reg_reg[834]  ( .D(out[834]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[834]) );
  DFF \round_reg_reg[835]  ( .D(out[835]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[835]) );
  DFF \round_reg_reg[836]  ( .D(out[836]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[836]) );
  DFF \round_reg_reg[837]  ( .D(out[837]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[837]) );
  DFF \round_reg_reg[838]  ( .D(out[838]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[838]) );
  DFF \round_reg_reg[839]  ( .D(out[839]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[839]) );
  DFF \round_reg_reg[840]  ( .D(out[840]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[840]) );
  DFF \round_reg_reg[841]  ( .D(out[841]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[841]) );
  DFF \round_reg_reg[842]  ( .D(out[842]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[842]) );
  DFF \round_reg_reg[843]  ( .D(out[843]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[843]) );
  DFF \round_reg_reg[844]  ( .D(out[844]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[844]) );
  DFF \round_reg_reg[845]  ( .D(out[845]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[845]) );
  DFF \round_reg_reg[846]  ( .D(out[846]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[846]) );
  DFF \round_reg_reg[847]  ( .D(out[847]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[847]) );
  DFF \round_reg_reg[848]  ( .D(out[848]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[848]) );
  DFF \round_reg_reg[849]  ( .D(out[849]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[849]) );
  DFF \round_reg_reg[850]  ( .D(out[850]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[850]) );
  DFF \round_reg_reg[851]  ( .D(out[851]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[851]) );
  DFF \round_reg_reg[852]  ( .D(out[852]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[852]) );
  DFF \round_reg_reg[853]  ( .D(out[853]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[853]) );
  DFF \round_reg_reg[854]  ( .D(out[854]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[854]) );
  DFF \round_reg_reg[855]  ( .D(out[855]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[855]) );
  DFF \round_reg_reg[856]  ( .D(out[856]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[856]) );
  DFF \round_reg_reg[857]  ( .D(out[857]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[857]) );
  DFF \round_reg_reg[858]  ( .D(out[858]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[858]) );
  DFF \round_reg_reg[859]  ( .D(out[859]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[859]) );
  DFF \round_reg_reg[860]  ( .D(out[860]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[860]) );
  DFF \round_reg_reg[861]  ( .D(out[861]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[861]) );
  DFF \round_reg_reg[862]  ( .D(out[862]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[862]) );
  DFF \round_reg_reg[863]  ( .D(out[863]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[863]) );
  DFF \round_reg_reg[864]  ( .D(out[864]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[864]) );
  DFF \round_reg_reg[865]  ( .D(out[865]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[865]) );
  DFF \round_reg_reg[866]  ( .D(out[866]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[866]) );
  DFF \round_reg_reg[867]  ( .D(out[867]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[867]) );
  DFF \round_reg_reg[868]  ( .D(out[868]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[868]) );
  DFF \round_reg_reg[869]  ( .D(out[869]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[869]) );
  DFF \round_reg_reg[870]  ( .D(out[870]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[870]) );
  DFF \round_reg_reg[871]  ( .D(out[871]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[871]) );
  DFF \round_reg_reg[872]  ( .D(out[872]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[872]) );
  DFF \round_reg_reg[873]  ( .D(out[873]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[873]) );
  DFF \round_reg_reg[874]  ( .D(out[874]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[874]) );
  DFF \round_reg_reg[875]  ( .D(out[875]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[875]) );
  DFF \round_reg_reg[876]  ( .D(out[876]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[876]) );
  DFF \round_reg_reg[877]  ( .D(out[877]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[877]) );
  DFF \round_reg_reg[878]  ( .D(out[878]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[878]) );
  DFF \round_reg_reg[879]  ( .D(out[879]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[879]) );
  DFF \round_reg_reg[880]  ( .D(out[880]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[880]) );
  DFF \round_reg_reg[881]  ( .D(out[881]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[881]) );
  DFF \round_reg_reg[882]  ( .D(out[882]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[882]) );
  DFF \round_reg_reg[883]  ( .D(out[883]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[883]) );
  DFF \round_reg_reg[884]  ( .D(out[884]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[884]) );
  DFF \round_reg_reg[885]  ( .D(out[885]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[885]) );
  DFF \round_reg_reg[886]  ( .D(out[886]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[886]) );
  DFF \round_reg_reg[887]  ( .D(out[887]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[887]) );
  DFF \round_reg_reg[888]  ( .D(out[888]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[888]) );
  DFF \round_reg_reg[889]  ( .D(out[889]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[889]) );
  DFF \round_reg_reg[890]  ( .D(out[890]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[890]) );
  DFF \round_reg_reg[891]  ( .D(out[891]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[891]) );
  DFF \round_reg_reg[892]  ( .D(out[892]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[892]) );
  DFF \round_reg_reg[893]  ( .D(out[893]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[893]) );
  DFF \round_reg_reg[894]  ( .D(out[894]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[894]) );
  DFF \round_reg_reg[895]  ( .D(out[895]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[895]) );
  DFF \round_reg_reg[896]  ( .D(out[896]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[896]) );
  DFF \round_reg_reg[897]  ( .D(out[897]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[897]) );
  DFF \round_reg_reg[898]  ( .D(out[898]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[898]) );
  DFF \round_reg_reg[899]  ( .D(out[899]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[899]) );
  DFF \round_reg_reg[900]  ( .D(out[900]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[900]) );
  DFF \round_reg_reg[901]  ( .D(out[901]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[901]) );
  DFF \round_reg_reg[902]  ( .D(out[902]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[902]) );
  DFF \round_reg_reg[903]  ( .D(out[903]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[903]) );
  DFF \round_reg_reg[904]  ( .D(out[904]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[904]) );
  DFF \round_reg_reg[905]  ( .D(out[905]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[905]) );
  DFF \round_reg_reg[906]  ( .D(out[906]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[906]) );
  DFF \round_reg_reg[907]  ( .D(out[907]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[907]) );
  DFF \round_reg_reg[908]  ( .D(out[908]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[908]) );
  DFF \round_reg_reg[909]  ( .D(out[909]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[909]) );
  DFF \round_reg_reg[910]  ( .D(out[910]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[910]) );
  DFF \round_reg_reg[911]  ( .D(out[911]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[911]) );
  DFF \round_reg_reg[912]  ( .D(out[912]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[912]) );
  DFF \round_reg_reg[913]  ( .D(out[913]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[913]) );
  DFF \round_reg_reg[914]  ( .D(out[914]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[914]) );
  DFF \round_reg_reg[915]  ( .D(out[915]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[915]) );
  DFF \round_reg_reg[916]  ( .D(out[916]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[916]) );
  DFF \round_reg_reg[917]  ( .D(out[917]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[917]) );
  DFF \round_reg_reg[918]  ( .D(out[918]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[918]) );
  DFF \round_reg_reg[919]  ( .D(out[919]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[919]) );
  DFF \round_reg_reg[920]  ( .D(out[920]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[920]) );
  DFF \round_reg_reg[921]  ( .D(out[921]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[921]) );
  DFF \round_reg_reg[922]  ( .D(out[922]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[922]) );
  DFF \round_reg_reg[923]  ( .D(out[923]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[923]) );
  DFF \round_reg_reg[924]  ( .D(out[924]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[924]) );
  DFF \round_reg_reg[925]  ( .D(out[925]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[925]) );
  DFF \round_reg_reg[926]  ( .D(out[926]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[926]) );
  DFF \round_reg_reg[927]  ( .D(out[927]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[927]) );
  DFF \round_reg_reg[928]  ( .D(out[928]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[928]) );
  DFF \round_reg_reg[929]  ( .D(out[929]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[929]) );
  DFF \round_reg_reg[930]  ( .D(out[930]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[930]) );
  DFF \round_reg_reg[931]  ( .D(out[931]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[931]) );
  DFF \round_reg_reg[932]  ( .D(out[932]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[932]) );
  DFF \round_reg_reg[933]  ( .D(out[933]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[933]) );
  DFF \round_reg_reg[934]  ( .D(out[934]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[934]) );
  DFF \round_reg_reg[935]  ( .D(out[935]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[935]) );
  DFF \round_reg_reg[936]  ( .D(out[936]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[936]) );
  DFF \round_reg_reg[937]  ( .D(out[937]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[937]) );
  DFF \round_reg_reg[938]  ( .D(out[938]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[938]) );
  DFF \round_reg_reg[939]  ( .D(out[939]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[939]) );
  DFF \round_reg_reg[940]  ( .D(out[940]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[940]) );
  DFF \round_reg_reg[941]  ( .D(out[941]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[941]) );
  DFF \round_reg_reg[942]  ( .D(out[942]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[942]) );
  DFF \round_reg_reg[943]  ( .D(out[943]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[943]) );
  DFF \round_reg_reg[944]  ( .D(out[944]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[944]) );
  DFF \round_reg_reg[945]  ( .D(out[945]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[945]) );
  DFF \round_reg_reg[946]  ( .D(out[946]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[946]) );
  DFF \round_reg_reg[947]  ( .D(out[947]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[947]) );
  DFF \round_reg_reg[948]  ( .D(out[948]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[948]) );
  DFF \round_reg_reg[949]  ( .D(out[949]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[949]) );
  DFF \round_reg_reg[950]  ( .D(out[950]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[950]) );
  DFF \round_reg_reg[951]  ( .D(out[951]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[951]) );
  DFF \round_reg_reg[952]  ( .D(out[952]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[952]) );
  DFF \round_reg_reg[953]  ( .D(out[953]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[953]) );
  DFF \round_reg_reg[954]  ( .D(out[954]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[954]) );
  DFF \round_reg_reg[955]  ( .D(out[955]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[955]) );
  DFF \round_reg_reg[956]  ( .D(out[956]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[956]) );
  DFF \round_reg_reg[957]  ( .D(out[957]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[957]) );
  DFF \round_reg_reg[958]  ( .D(out[958]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[958]) );
  DFF \round_reg_reg[959]  ( .D(out[959]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[959]) );
  DFF \round_reg_reg[960]  ( .D(out[960]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[960]) );
  DFF \round_reg_reg[961]  ( .D(out[961]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[961]) );
  DFF \round_reg_reg[962]  ( .D(out[962]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[962]) );
  DFF \round_reg_reg[963]  ( .D(out[963]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[963]) );
  DFF \round_reg_reg[964]  ( .D(out[964]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[964]) );
  DFF \round_reg_reg[965]  ( .D(out[965]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[965]) );
  DFF \round_reg_reg[966]  ( .D(out[966]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[966]) );
  DFF \round_reg_reg[967]  ( .D(out[967]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[967]) );
  DFF \round_reg_reg[968]  ( .D(out[968]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[968]) );
  DFF \round_reg_reg[969]  ( .D(out[969]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[969]) );
  DFF \round_reg_reg[970]  ( .D(out[970]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[970]) );
  DFF \round_reg_reg[971]  ( .D(out[971]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[971]) );
  DFF \round_reg_reg[972]  ( .D(out[972]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[972]) );
  DFF \round_reg_reg[973]  ( .D(out[973]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[973]) );
  DFF \round_reg_reg[974]  ( .D(out[974]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[974]) );
  DFF \round_reg_reg[975]  ( .D(out[975]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[975]) );
  DFF \round_reg_reg[976]  ( .D(out[976]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[976]) );
  DFF \round_reg_reg[977]  ( .D(out[977]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[977]) );
  DFF \round_reg_reg[978]  ( .D(out[978]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[978]) );
  DFF \round_reg_reg[979]  ( .D(out[979]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[979]) );
  DFF \round_reg_reg[980]  ( .D(out[980]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[980]) );
  DFF \round_reg_reg[981]  ( .D(out[981]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[981]) );
  DFF \round_reg_reg[982]  ( .D(out[982]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[982]) );
  DFF \round_reg_reg[983]  ( .D(out[983]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[983]) );
  DFF \round_reg_reg[984]  ( .D(out[984]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[984]) );
  DFF \round_reg_reg[985]  ( .D(out[985]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[985]) );
  DFF \round_reg_reg[986]  ( .D(out[986]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[986]) );
  DFF \round_reg_reg[987]  ( .D(out[987]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[987]) );
  DFF \round_reg_reg[988]  ( .D(out[988]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[988]) );
  DFF \round_reg_reg[989]  ( .D(out[989]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[989]) );
  DFF \round_reg_reg[990]  ( .D(out[990]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[990]) );
  DFF \round_reg_reg[991]  ( .D(out[991]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[991]) );
  DFF \round_reg_reg[992]  ( .D(out[992]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[992]) );
  DFF \round_reg_reg[993]  ( .D(out[993]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[993]) );
  DFF \round_reg_reg[994]  ( .D(out[994]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[994]) );
  DFF \round_reg_reg[995]  ( .D(out[995]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[995]) );
  DFF \round_reg_reg[996]  ( .D(out[996]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[996]) );
  DFF \round_reg_reg[997]  ( .D(out[997]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[997]) );
  DFF \round_reg_reg[998]  ( .D(out[998]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[998]) );
  DFF \round_reg_reg[999]  ( .D(out[999]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[999]) );
  DFF \round_reg_reg[1000]  ( .D(out[1000]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1000]) );
  DFF \round_reg_reg[1001]  ( .D(out[1001]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1001]) );
  DFF \round_reg_reg[1002]  ( .D(out[1002]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1002]) );
  DFF \round_reg_reg[1003]  ( .D(out[1003]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1003]) );
  DFF \round_reg_reg[1004]  ( .D(out[1004]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1004]) );
  DFF \round_reg_reg[1005]  ( .D(out[1005]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1005]) );
  DFF \round_reg_reg[1006]  ( .D(out[1006]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1006]) );
  DFF \round_reg_reg[1007]  ( .D(out[1007]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1007]) );
  DFF \round_reg_reg[1008]  ( .D(out[1008]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1008]) );
  DFF \round_reg_reg[1009]  ( .D(out[1009]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1009]) );
  DFF \round_reg_reg[1010]  ( .D(out[1010]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1010]) );
  DFF \round_reg_reg[1011]  ( .D(out[1011]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1011]) );
  DFF \round_reg_reg[1012]  ( .D(out[1012]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1012]) );
  DFF \round_reg_reg[1013]  ( .D(out[1013]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1013]) );
  DFF \round_reg_reg[1014]  ( .D(out[1014]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1014]) );
  DFF \round_reg_reg[1015]  ( .D(out[1015]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1015]) );
  DFF \round_reg_reg[1016]  ( .D(out[1016]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1016]) );
  DFF \round_reg_reg[1017]  ( .D(out[1017]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1017]) );
  DFF \round_reg_reg[1018]  ( .D(out[1018]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1018]) );
  DFF \round_reg_reg[1019]  ( .D(out[1019]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1019]) );
  DFF \round_reg_reg[1020]  ( .D(out[1020]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1020]) );
  DFF \round_reg_reg[1021]  ( .D(out[1021]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1021]) );
  DFF \round_reg_reg[1022]  ( .D(out[1022]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1022]) );
  DFF \round_reg_reg[1023]  ( .D(out[1023]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1023]) );
  DFF \round_reg_reg[1024]  ( .D(out[1024]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1024]) );
  DFF \round_reg_reg[1025]  ( .D(out[1025]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1025]) );
  DFF \round_reg_reg[1026]  ( .D(out[1026]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1026]) );
  DFF \round_reg_reg[1027]  ( .D(out[1027]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1027]) );
  DFF \round_reg_reg[1028]  ( .D(out[1028]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1028]) );
  DFF \round_reg_reg[1029]  ( .D(out[1029]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1029]) );
  DFF \round_reg_reg[1030]  ( .D(out[1030]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1030]) );
  DFF \round_reg_reg[1031]  ( .D(out[1031]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1031]) );
  DFF \round_reg_reg[1032]  ( .D(out[1032]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1032]) );
  DFF \round_reg_reg[1033]  ( .D(out[1033]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1033]) );
  DFF \round_reg_reg[1034]  ( .D(out[1034]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1034]) );
  DFF \round_reg_reg[1035]  ( .D(out[1035]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1035]) );
  DFF \round_reg_reg[1036]  ( .D(out[1036]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1036]) );
  DFF \round_reg_reg[1037]  ( .D(out[1037]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1037]) );
  DFF \round_reg_reg[1038]  ( .D(out[1038]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1038]) );
  DFF \round_reg_reg[1039]  ( .D(out[1039]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1039]) );
  DFF \round_reg_reg[1040]  ( .D(out[1040]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1040]) );
  DFF \round_reg_reg[1041]  ( .D(out[1041]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1041]) );
  DFF \round_reg_reg[1042]  ( .D(out[1042]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1042]) );
  DFF \round_reg_reg[1043]  ( .D(out[1043]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1043]) );
  DFF \round_reg_reg[1044]  ( .D(out[1044]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1044]) );
  DFF \round_reg_reg[1045]  ( .D(out[1045]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1045]) );
  DFF \round_reg_reg[1046]  ( .D(out[1046]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1046]) );
  DFF \round_reg_reg[1047]  ( .D(out[1047]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1047]) );
  DFF \round_reg_reg[1048]  ( .D(out[1048]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1048]) );
  DFF \round_reg_reg[1049]  ( .D(out[1049]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1049]) );
  DFF \round_reg_reg[1050]  ( .D(out[1050]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1050]) );
  DFF \round_reg_reg[1051]  ( .D(out[1051]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1051]) );
  DFF \round_reg_reg[1052]  ( .D(out[1052]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1052]) );
  DFF \round_reg_reg[1053]  ( .D(out[1053]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1053]) );
  DFF \round_reg_reg[1054]  ( .D(out[1054]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1054]) );
  DFF \round_reg_reg[1055]  ( .D(out[1055]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1055]) );
  DFF \round_reg_reg[1056]  ( .D(out[1056]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1056]) );
  DFF \round_reg_reg[1057]  ( .D(out[1057]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1057]) );
  DFF \round_reg_reg[1058]  ( .D(out[1058]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1058]) );
  DFF \round_reg_reg[1059]  ( .D(out[1059]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1059]) );
  DFF \round_reg_reg[1060]  ( .D(out[1060]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1060]) );
  DFF \round_reg_reg[1061]  ( .D(out[1061]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1061]) );
  DFF \round_reg_reg[1062]  ( .D(out[1062]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1062]) );
  DFF \round_reg_reg[1063]  ( .D(out[1063]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1063]) );
  DFF \round_reg_reg[1064]  ( .D(out[1064]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1064]) );
  DFF \round_reg_reg[1065]  ( .D(out[1065]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1065]) );
  DFF \round_reg_reg[1066]  ( .D(out[1066]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1066]) );
  DFF \round_reg_reg[1067]  ( .D(out[1067]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1067]) );
  DFF \round_reg_reg[1068]  ( .D(out[1068]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1068]) );
  DFF \round_reg_reg[1069]  ( .D(out[1069]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1069]) );
  DFF \round_reg_reg[1070]  ( .D(out[1070]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1070]) );
  DFF \round_reg_reg[1071]  ( .D(out[1071]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1071]) );
  DFF \round_reg_reg[1072]  ( .D(out[1072]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1072]) );
  DFF \round_reg_reg[1073]  ( .D(out[1073]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1073]) );
  DFF \round_reg_reg[1074]  ( .D(out[1074]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1074]) );
  DFF \round_reg_reg[1075]  ( .D(out[1075]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1075]) );
  DFF \round_reg_reg[1076]  ( .D(out[1076]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1076]) );
  DFF \round_reg_reg[1077]  ( .D(out[1077]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1077]) );
  DFF \round_reg_reg[1078]  ( .D(out[1078]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1078]) );
  DFF \round_reg_reg[1079]  ( .D(out[1079]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1079]) );
  DFF \round_reg_reg[1080]  ( .D(out[1080]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1080]) );
  DFF \round_reg_reg[1081]  ( .D(out[1081]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1081]) );
  DFF \round_reg_reg[1082]  ( .D(out[1082]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1082]) );
  DFF \round_reg_reg[1083]  ( .D(out[1083]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1083]) );
  DFF \round_reg_reg[1084]  ( .D(out[1084]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1084]) );
  DFF \round_reg_reg[1085]  ( .D(out[1085]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1085]) );
  DFF \round_reg_reg[1086]  ( .D(out[1086]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1086]) );
  DFF \round_reg_reg[1087]  ( .D(out[1087]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1087]) );
  DFF \round_reg_reg[1088]  ( .D(out[1088]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1088]) );
  DFF \round_reg_reg[1089]  ( .D(out[1089]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1089]) );
  DFF \round_reg_reg[1090]  ( .D(out[1090]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1090]) );
  DFF \round_reg_reg[1091]  ( .D(out[1091]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1091]) );
  DFF \round_reg_reg[1092]  ( .D(out[1092]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1092]) );
  DFF \round_reg_reg[1093]  ( .D(out[1093]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1093]) );
  DFF \round_reg_reg[1094]  ( .D(out[1094]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1094]) );
  DFF \round_reg_reg[1095]  ( .D(out[1095]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1095]) );
  DFF \round_reg_reg[1096]  ( .D(out[1096]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1096]) );
  DFF \round_reg_reg[1097]  ( .D(out[1097]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1097]) );
  DFF \round_reg_reg[1098]  ( .D(out[1098]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1098]) );
  DFF \round_reg_reg[1099]  ( .D(out[1099]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1099]) );
  DFF \round_reg_reg[1100]  ( .D(out[1100]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1100]) );
  DFF \round_reg_reg[1101]  ( .D(out[1101]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1101]) );
  DFF \round_reg_reg[1102]  ( .D(out[1102]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1102]) );
  DFF \round_reg_reg[1103]  ( .D(out[1103]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1103]) );
  DFF \round_reg_reg[1104]  ( .D(out[1104]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1104]) );
  DFF \round_reg_reg[1105]  ( .D(out[1105]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1105]) );
  DFF \round_reg_reg[1106]  ( .D(out[1106]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1106]) );
  DFF \round_reg_reg[1107]  ( .D(out[1107]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1107]) );
  DFF \round_reg_reg[1108]  ( .D(out[1108]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1108]) );
  DFF \round_reg_reg[1109]  ( .D(out[1109]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1109]) );
  DFF \round_reg_reg[1110]  ( .D(out[1110]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1110]) );
  DFF \round_reg_reg[1111]  ( .D(out[1111]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1111]) );
  DFF \round_reg_reg[1112]  ( .D(out[1112]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1112]) );
  DFF \round_reg_reg[1113]  ( .D(out[1113]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1113]) );
  DFF \round_reg_reg[1114]  ( .D(out[1114]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1114]) );
  DFF \round_reg_reg[1115]  ( .D(out[1115]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1115]) );
  DFF \round_reg_reg[1116]  ( .D(out[1116]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1116]) );
  DFF \round_reg_reg[1117]  ( .D(out[1117]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1117]) );
  DFF \round_reg_reg[1118]  ( .D(out[1118]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1118]) );
  DFF \round_reg_reg[1119]  ( .D(out[1119]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1119]) );
  DFF \round_reg_reg[1120]  ( .D(out[1120]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1120]) );
  DFF \round_reg_reg[1121]  ( .D(out[1121]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1121]) );
  DFF \round_reg_reg[1122]  ( .D(out[1122]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1122]) );
  DFF \round_reg_reg[1123]  ( .D(out[1123]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1123]) );
  DFF \round_reg_reg[1124]  ( .D(out[1124]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1124]) );
  DFF \round_reg_reg[1125]  ( .D(out[1125]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1125]) );
  DFF \round_reg_reg[1126]  ( .D(out[1126]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1126]) );
  DFF \round_reg_reg[1127]  ( .D(out[1127]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1127]) );
  DFF \round_reg_reg[1128]  ( .D(out[1128]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1128]) );
  DFF \round_reg_reg[1129]  ( .D(out[1129]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1129]) );
  DFF \round_reg_reg[1130]  ( .D(out[1130]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1130]) );
  DFF \round_reg_reg[1131]  ( .D(out[1131]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1131]) );
  DFF \round_reg_reg[1132]  ( .D(out[1132]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1132]) );
  DFF \round_reg_reg[1133]  ( .D(out[1133]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1133]) );
  DFF \round_reg_reg[1134]  ( .D(out[1134]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1134]) );
  DFF \round_reg_reg[1135]  ( .D(out[1135]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1135]) );
  DFF \round_reg_reg[1136]  ( .D(out[1136]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1136]) );
  DFF \round_reg_reg[1137]  ( .D(out[1137]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1137]) );
  DFF \round_reg_reg[1138]  ( .D(out[1138]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1138]) );
  DFF \round_reg_reg[1139]  ( .D(out[1139]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1139]) );
  DFF \round_reg_reg[1140]  ( .D(out[1140]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1140]) );
  DFF \round_reg_reg[1141]  ( .D(out[1141]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1141]) );
  DFF \round_reg_reg[1142]  ( .D(out[1142]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1142]) );
  DFF \round_reg_reg[1143]  ( .D(out[1143]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1143]) );
  DFF \round_reg_reg[1144]  ( .D(out[1144]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1144]) );
  DFF \round_reg_reg[1145]  ( .D(out[1145]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1145]) );
  DFF \round_reg_reg[1146]  ( .D(out[1146]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1146]) );
  DFF \round_reg_reg[1147]  ( .D(out[1147]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1147]) );
  DFF \round_reg_reg[1148]  ( .D(out[1148]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1148]) );
  DFF \round_reg_reg[1149]  ( .D(out[1149]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1149]) );
  DFF \round_reg_reg[1150]  ( .D(out[1150]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1150]) );
  DFF \round_reg_reg[1151]  ( .D(out[1151]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1151]) );
  DFF \round_reg_reg[1152]  ( .D(out[1152]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1152]) );
  DFF \round_reg_reg[1153]  ( .D(out[1153]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1153]) );
  DFF \round_reg_reg[1154]  ( .D(out[1154]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1154]) );
  DFF \round_reg_reg[1155]  ( .D(out[1155]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1155]) );
  DFF \round_reg_reg[1156]  ( .D(out[1156]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1156]) );
  DFF \round_reg_reg[1157]  ( .D(out[1157]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1157]) );
  DFF \round_reg_reg[1158]  ( .D(out[1158]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1158]) );
  DFF \round_reg_reg[1159]  ( .D(out[1159]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1159]) );
  DFF \round_reg_reg[1160]  ( .D(out[1160]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1160]) );
  DFF \round_reg_reg[1161]  ( .D(out[1161]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1161]) );
  DFF \round_reg_reg[1162]  ( .D(out[1162]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1162]) );
  DFF \round_reg_reg[1163]  ( .D(out[1163]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1163]) );
  DFF \round_reg_reg[1164]  ( .D(out[1164]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1164]) );
  DFF \round_reg_reg[1165]  ( .D(out[1165]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1165]) );
  DFF \round_reg_reg[1166]  ( .D(out[1166]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1166]) );
  DFF \round_reg_reg[1167]  ( .D(out[1167]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1167]) );
  DFF \round_reg_reg[1168]  ( .D(out[1168]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1168]) );
  DFF \round_reg_reg[1169]  ( .D(out[1169]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1169]) );
  DFF \round_reg_reg[1170]  ( .D(out[1170]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1170]) );
  DFF \round_reg_reg[1171]  ( .D(out[1171]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1171]) );
  DFF \round_reg_reg[1172]  ( .D(out[1172]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1172]) );
  DFF \round_reg_reg[1173]  ( .D(out[1173]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1173]) );
  DFF \round_reg_reg[1174]  ( .D(out[1174]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1174]) );
  DFF \round_reg_reg[1175]  ( .D(out[1175]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1175]) );
  DFF \round_reg_reg[1176]  ( .D(out[1176]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1176]) );
  DFF \round_reg_reg[1177]  ( .D(out[1177]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1177]) );
  DFF \round_reg_reg[1178]  ( .D(out[1178]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1178]) );
  DFF \round_reg_reg[1179]  ( .D(out[1179]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1179]) );
  DFF \round_reg_reg[1180]  ( .D(out[1180]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1180]) );
  DFF \round_reg_reg[1181]  ( .D(out[1181]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1181]) );
  DFF \round_reg_reg[1182]  ( .D(out[1182]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1182]) );
  DFF \round_reg_reg[1183]  ( .D(out[1183]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1183]) );
  DFF \round_reg_reg[1184]  ( .D(out[1184]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1184]) );
  DFF \round_reg_reg[1185]  ( .D(out[1185]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1185]) );
  DFF \round_reg_reg[1186]  ( .D(out[1186]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1186]) );
  DFF \round_reg_reg[1187]  ( .D(out[1187]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1187]) );
  DFF \round_reg_reg[1188]  ( .D(out[1188]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1188]) );
  DFF \round_reg_reg[1189]  ( .D(out[1189]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1189]) );
  DFF \round_reg_reg[1190]  ( .D(out[1190]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1190]) );
  DFF \round_reg_reg[1191]  ( .D(out[1191]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1191]) );
  DFF \round_reg_reg[1192]  ( .D(out[1192]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1192]) );
  DFF \round_reg_reg[1193]  ( .D(out[1193]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1193]) );
  DFF \round_reg_reg[1194]  ( .D(out[1194]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1194]) );
  DFF \round_reg_reg[1195]  ( .D(out[1195]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1195]) );
  DFF \round_reg_reg[1196]  ( .D(out[1196]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1196]) );
  DFF \round_reg_reg[1197]  ( .D(out[1197]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1197]) );
  DFF \round_reg_reg[1198]  ( .D(out[1198]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1198]) );
  DFF \round_reg_reg[1199]  ( .D(out[1199]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1199]) );
  DFF \round_reg_reg[1200]  ( .D(out[1200]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1200]) );
  DFF \round_reg_reg[1201]  ( .D(out[1201]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1201]) );
  DFF \round_reg_reg[1202]  ( .D(out[1202]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1202]) );
  DFF \round_reg_reg[1203]  ( .D(out[1203]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1203]) );
  DFF \round_reg_reg[1204]  ( .D(out[1204]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1204]) );
  DFF \round_reg_reg[1205]  ( .D(out[1205]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1205]) );
  DFF \round_reg_reg[1206]  ( .D(out[1206]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1206]) );
  DFF \round_reg_reg[1207]  ( .D(out[1207]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1207]) );
  DFF \round_reg_reg[1208]  ( .D(out[1208]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1208]) );
  DFF \round_reg_reg[1209]  ( .D(out[1209]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1209]) );
  DFF \round_reg_reg[1210]  ( .D(out[1210]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1210]) );
  DFF \round_reg_reg[1211]  ( .D(out[1211]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1211]) );
  DFF \round_reg_reg[1212]  ( .D(out[1212]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1212]) );
  DFF \round_reg_reg[1213]  ( .D(out[1213]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1213]) );
  DFF \round_reg_reg[1214]  ( .D(out[1214]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1214]) );
  DFF \round_reg_reg[1215]  ( .D(out[1215]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1215]) );
  DFF \round_reg_reg[1216]  ( .D(out[1216]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1216]) );
  DFF \round_reg_reg[1217]  ( .D(out[1217]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1217]) );
  DFF \round_reg_reg[1218]  ( .D(out[1218]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1218]) );
  DFF \round_reg_reg[1219]  ( .D(out[1219]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1219]) );
  DFF \round_reg_reg[1220]  ( .D(out[1220]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1220]) );
  DFF \round_reg_reg[1221]  ( .D(out[1221]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1221]) );
  DFF \round_reg_reg[1222]  ( .D(out[1222]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1222]) );
  DFF \round_reg_reg[1223]  ( .D(out[1223]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1223]) );
  DFF \round_reg_reg[1224]  ( .D(out[1224]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1224]) );
  DFF \round_reg_reg[1225]  ( .D(out[1225]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1225]) );
  DFF \round_reg_reg[1226]  ( .D(out[1226]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1226]) );
  DFF \round_reg_reg[1227]  ( .D(out[1227]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1227]) );
  DFF \round_reg_reg[1228]  ( .D(out[1228]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1228]) );
  DFF \round_reg_reg[1229]  ( .D(out[1229]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1229]) );
  DFF \round_reg_reg[1230]  ( .D(out[1230]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1230]) );
  DFF \round_reg_reg[1231]  ( .D(out[1231]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1231]) );
  DFF \round_reg_reg[1232]  ( .D(out[1232]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1232]) );
  DFF \round_reg_reg[1233]  ( .D(out[1233]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1233]) );
  DFF \round_reg_reg[1234]  ( .D(out[1234]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1234]) );
  DFF \round_reg_reg[1235]  ( .D(out[1235]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1235]) );
  DFF \round_reg_reg[1236]  ( .D(out[1236]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1236]) );
  DFF \round_reg_reg[1237]  ( .D(out[1237]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1237]) );
  DFF \round_reg_reg[1238]  ( .D(out[1238]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1238]) );
  DFF \round_reg_reg[1239]  ( .D(out[1239]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1239]) );
  DFF \round_reg_reg[1240]  ( .D(out[1240]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1240]) );
  DFF \round_reg_reg[1241]  ( .D(out[1241]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1241]) );
  DFF \round_reg_reg[1242]  ( .D(out[1242]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1242]) );
  DFF \round_reg_reg[1243]  ( .D(out[1243]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1243]) );
  DFF \round_reg_reg[1244]  ( .D(out[1244]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1244]) );
  DFF \round_reg_reg[1245]  ( .D(out[1245]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1245]) );
  DFF \round_reg_reg[1246]  ( .D(out[1246]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1246]) );
  DFF \round_reg_reg[1247]  ( .D(out[1247]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1247]) );
  DFF \round_reg_reg[1248]  ( .D(out[1248]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1248]) );
  DFF \round_reg_reg[1249]  ( .D(out[1249]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1249]) );
  DFF \round_reg_reg[1250]  ( .D(out[1250]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1250]) );
  DFF \round_reg_reg[1251]  ( .D(out[1251]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1251]) );
  DFF \round_reg_reg[1252]  ( .D(out[1252]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1252]) );
  DFF \round_reg_reg[1253]  ( .D(out[1253]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1253]) );
  DFF \round_reg_reg[1254]  ( .D(out[1254]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1254]) );
  DFF \round_reg_reg[1255]  ( .D(out[1255]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1255]) );
  DFF \round_reg_reg[1256]  ( .D(out[1256]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1256]) );
  DFF \round_reg_reg[1257]  ( .D(out[1257]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1257]) );
  DFF \round_reg_reg[1258]  ( .D(out[1258]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1258]) );
  DFF \round_reg_reg[1259]  ( .D(out[1259]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1259]) );
  DFF \round_reg_reg[1260]  ( .D(out[1260]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1260]) );
  DFF \round_reg_reg[1261]  ( .D(out[1261]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1261]) );
  DFF \round_reg_reg[1262]  ( .D(out[1262]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1262]) );
  DFF \round_reg_reg[1263]  ( .D(out[1263]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1263]) );
  DFF \round_reg_reg[1264]  ( .D(out[1264]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1264]) );
  DFF \round_reg_reg[1265]  ( .D(out[1265]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1265]) );
  DFF \round_reg_reg[1266]  ( .D(out[1266]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1266]) );
  DFF \round_reg_reg[1267]  ( .D(out[1267]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1267]) );
  DFF \round_reg_reg[1268]  ( .D(out[1268]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1268]) );
  DFF \round_reg_reg[1269]  ( .D(out[1269]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1269]) );
  DFF \round_reg_reg[1270]  ( .D(out[1270]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1270]) );
  DFF \round_reg_reg[1271]  ( .D(out[1271]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1271]) );
  DFF \round_reg_reg[1272]  ( .D(out[1272]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1272]) );
  DFF \round_reg_reg[1273]  ( .D(out[1273]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1273]) );
  DFF \round_reg_reg[1274]  ( .D(out[1274]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1274]) );
  DFF \round_reg_reg[1275]  ( .D(out[1275]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1275]) );
  DFF \round_reg_reg[1276]  ( .D(out[1276]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1276]) );
  DFF \round_reg_reg[1277]  ( .D(out[1277]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1277]) );
  DFF \round_reg_reg[1278]  ( .D(out[1278]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1278]) );
  DFF \round_reg_reg[1279]  ( .D(out[1279]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1279]) );
  DFF \round_reg_reg[1280]  ( .D(out[1280]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1280]) );
  DFF \round_reg_reg[1281]  ( .D(out[1281]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1281]) );
  DFF \round_reg_reg[1282]  ( .D(out[1282]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1282]) );
  DFF \round_reg_reg[1283]  ( .D(out[1283]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1283]) );
  DFF \round_reg_reg[1284]  ( .D(out[1284]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1284]) );
  DFF \round_reg_reg[1285]  ( .D(out[1285]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1285]) );
  DFF \round_reg_reg[1286]  ( .D(out[1286]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1286]) );
  DFF \round_reg_reg[1287]  ( .D(out[1287]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1287]) );
  DFF \round_reg_reg[1288]  ( .D(out[1288]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1288]) );
  DFF \round_reg_reg[1289]  ( .D(out[1289]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1289]) );
  DFF \round_reg_reg[1290]  ( .D(out[1290]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1290]) );
  DFF \round_reg_reg[1291]  ( .D(out[1291]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1291]) );
  DFF \round_reg_reg[1292]  ( .D(out[1292]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1292]) );
  DFF \round_reg_reg[1293]  ( .D(out[1293]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1293]) );
  DFF \round_reg_reg[1294]  ( .D(out[1294]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1294]) );
  DFF \round_reg_reg[1295]  ( .D(out[1295]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1295]) );
  DFF \round_reg_reg[1296]  ( .D(out[1296]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1296]) );
  DFF \round_reg_reg[1297]  ( .D(out[1297]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1297]) );
  DFF \round_reg_reg[1298]  ( .D(out[1298]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1298]) );
  DFF \round_reg_reg[1299]  ( .D(out[1299]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1299]) );
  DFF \round_reg_reg[1300]  ( .D(out[1300]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1300]) );
  DFF \round_reg_reg[1301]  ( .D(out[1301]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1301]) );
  DFF \round_reg_reg[1302]  ( .D(out[1302]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1302]) );
  DFF \round_reg_reg[1303]  ( .D(out[1303]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1303]) );
  DFF \round_reg_reg[1304]  ( .D(out[1304]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1304]) );
  DFF \round_reg_reg[1305]  ( .D(out[1305]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1305]) );
  DFF \round_reg_reg[1306]  ( .D(out[1306]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1306]) );
  DFF \round_reg_reg[1307]  ( .D(out[1307]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1307]) );
  DFF \round_reg_reg[1308]  ( .D(out[1308]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1308]) );
  DFF \round_reg_reg[1309]  ( .D(out[1309]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1309]) );
  DFF \round_reg_reg[1310]  ( .D(out[1310]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1310]) );
  DFF \round_reg_reg[1311]  ( .D(out[1311]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1311]) );
  DFF \round_reg_reg[1312]  ( .D(out[1312]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1312]) );
  DFF \round_reg_reg[1313]  ( .D(out[1313]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1313]) );
  DFF \round_reg_reg[1314]  ( .D(out[1314]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1314]) );
  DFF \round_reg_reg[1315]  ( .D(out[1315]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1315]) );
  DFF \round_reg_reg[1316]  ( .D(out[1316]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1316]) );
  DFF \round_reg_reg[1317]  ( .D(out[1317]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1317]) );
  DFF \round_reg_reg[1318]  ( .D(out[1318]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1318]) );
  DFF \round_reg_reg[1319]  ( .D(out[1319]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1319]) );
  DFF \round_reg_reg[1320]  ( .D(out[1320]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1320]) );
  DFF \round_reg_reg[1321]  ( .D(out[1321]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1321]) );
  DFF \round_reg_reg[1322]  ( .D(out[1322]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1322]) );
  DFF \round_reg_reg[1323]  ( .D(out[1323]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1323]) );
  DFF \round_reg_reg[1324]  ( .D(out[1324]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1324]) );
  DFF \round_reg_reg[1325]  ( .D(out[1325]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1325]) );
  DFF \round_reg_reg[1326]  ( .D(out[1326]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1326]) );
  DFF \round_reg_reg[1327]  ( .D(out[1327]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1327]) );
  DFF \round_reg_reg[1328]  ( .D(out[1328]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1328]) );
  DFF \round_reg_reg[1329]  ( .D(out[1329]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1329]) );
  DFF \round_reg_reg[1330]  ( .D(out[1330]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1330]) );
  DFF \round_reg_reg[1331]  ( .D(out[1331]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1331]) );
  DFF \round_reg_reg[1332]  ( .D(out[1332]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1332]) );
  DFF \round_reg_reg[1333]  ( .D(out[1333]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1333]) );
  DFF \round_reg_reg[1334]  ( .D(out[1334]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1334]) );
  DFF \round_reg_reg[1335]  ( .D(out[1335]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1335]) );
  DFF \round_reg_reg[1336]  ( .D(out[1336]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1336]) );
  DFF \round_reg_reg[1337]  ( .D(out[1337]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1337]) );
  DFF \round_reg_reg[1338]  ( .D(out[1338]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1338]) );
  DFF \round_reg_reg[1339]  ( .D(out[1339]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1339]) );
  DFF \round_reg_reg[1340]  ( .D(out[1340]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1340]) );
  DFF \round_reg_reg[1341]  ( .D(out[1341]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1341]) );
  DFF \round_reg_reg[1342]  ( .D(out[1342]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1342]) );
  DFF \round_reg_reg[1343]  ( .D(out[1343]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1343]) );
  DFF \round_reg_reg[1344]  ( .D(out[1344]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1344]) );
  DFF \round_reg_reg[1345]  ( .D(out[1345]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1345]) );
  DFF \round_reg_reg[1346]  ( .D(out[1346]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1346]) );
  DFF \round_reg_reg[1347]  ( .D(out[1347]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1347]) );
  DFF \round_reg_reg[1348]  ( .D(out[1348]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1348]) );
  DFF \round_reg_reg[1349]  ( .D(out[1349]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1349]) );
  DFF \round_reg_reg[1350]  ( .D(out[1350]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1350]) );
  DFF \round_reg_reg[1351]  ( .D(out[1351]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1351]) );
  DFF \round_reg_reg[1352]  ( .D(out[1352]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1352]) );
  DFF \round_reg_reg[1353]  ( .D(out[1353]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1353]) );
  DFF \round_reg_reg[1354]  ( .D(out[1354]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1354]) );
  DFF \round_reg_reg[1355]  ( .D(out[1355]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1355]) );
  DFF \round_reg_reg[1356]  ( .D(out[1356]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1356]) );
  DFF \round_reg_reg[1357]  ( .D(out[1357]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1357]) );
  DFF \round_reg_reg[1358]  ( .D(out[1358]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1358]) );
  DFF \round_reg_reg[1359]  ( .D(out[1359]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1359]) );
  DFF \round_reg_reg[1360]  ( .D(out[1360]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1360]) );
  DFF \round_reg_reg[1361]  ( .D(out[1361]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1361]) );
  DFF \round_reg_reg[1362]  ( .D(out[1362]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1362]) );
  DFF \round_reg_reg[1363]  ( .D(out[1363]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1363]) );
  DFF \round_reg_reg[1364]  ( .D(out[1364]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1364]) );
  DFF \round_reg_reg[1365]  ( .D(out[1365]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1365]) );
  DFF \round_reg_reg[1366]  ( .D(out[1366]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1366]) );
  DFF \round_reg_reg[1367]  ( .D(out[1367]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1367]) );
  DFF \round_reg_reg[1368]  ( .D(out[1368]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1368]) );
  DFF \round_reg_reg[1369]  ( .D(out[1369]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1369]) );
  DFF \round_reg_reg[1370]  ( .D(out[1370]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1370]) );
  DFF \round_reg_reg[1371]  ( .D(out[1371]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1371]) );
  DFF \round_reg_reg[1372]  ( .D(out[1372]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1372]) );
  DFF \round_reg_reg[1373]  ( .D(out[1373]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1373]) );
  DFF \round_reg_reg[1374]  ( .D(out[1374]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1374]) );
  DFF \round_reg_reg[1375]  ( .D(out[1375]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1375]) );
  DFF \round_reg_reg[1376]  ( .D(out[1376]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1376]) );
  DFF \round_reg_reg[1377]  ( .D(out[1377]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1377]) );
  DFF \round_reg_reg[1378]  ( .D(out[1378]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1378]) );
  DFF \round_reg_reg[1379]  ( .D(out[1379]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1379]) );
  DFF \round_reg_reg[1380]  ( .D(out[1380]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1380]) );
  DFF \round_reg_reg[1381]  ( .D(out[1381]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1381]) );
  DFF \round_reg_reg[1382]  ( .D(out[1382]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1382]) );
  DFF \round_reg_reg[1383]  ( .D(out[1383]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1383]) );
  DFF \round_reg_reg[1384]  ( .D(out[1384]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1384]) );
  DFF \round_reg_reg[1385]  ( .D(out[1385]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1385]) );
  DFF \round_reg_reg[1386]  ( .D(out[1386]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1386]) );
  DFF \round_reg_reg[1387]  ( .D(out[1387]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1387]) );
  DFF \round_reg_reg[1388]  ( .D(out[1388]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1388]) );
  DFF \round_reg_reg[1389]  ( .D(out[1389]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1389]) );
  DFF \round_reg_reg[1390]  ( .D(out[1390]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1390]) );
  DFF \round_reg_reg[1391]  ( .D(out[1391]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1391]) );
  DFF \round_reg_reg[1392]  ( .D(out[1392]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1392]) );
  DFF \round_reg_reg[1393]  ( .D(out[1393]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1393]) );
  DFF \round_reg_reg[1394]  ( .D(out[1394]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1394]) );
  DFF \round_reg_reg[1395]  ( .D(out[1395]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1395]) );
  DFF \round_reg_reg[1396]  ( .D(out[1396]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1396]) );
  DFF \round_reg_reg[1397]  ( .D(out[1397]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1397]) );
  DFF \round_reg_reg[1398]  ( .D(out[1398]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1398]) );
  DFF \round_reg_reg[1399]  ( .D(out[1399]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1399]) );
  DFF \round_reg_reg[1400]  ( .D(out[1400]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1400]) );
  DFF \round_reg_reg[1401]  ( .D(out[1401]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1401]) );
  DFF \round_reg_reg[1402]  ( .D(out[1402]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1402]) );
  DFF \round_reg_reg[1403]  ( .D(out[1403]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1403]) );
  DFF \round_reg_reg[1404]  ( .D(out[1404]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1404]) );
  DFF \round_reg_reg[1405]  ( .D(out[1405]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1405]) );
  DFF \round_reg_reg[1406]  ( .D(out[1406]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1406]) );
  DFF \round_reg_reg[1407]  ( .D(out[1407]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1407]) );
  DFF \round_reg_reg[1408]  ( .D(out[1408]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1408]) );
  DFF \round_reg_reg[1409]  ( .D(out[1409]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1409]) );
  DFF \round_reg_reg[1410]  ( .D(out[1410]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1410]) );
  DFF \round_reg_reg[1411]  ( .D(out[1411]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1411]) );
  DFF \round_reg_reg[1412]  ( .D(out[1412]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1412]) );
  DFF \round_reg_reg[1413]  ( .D(out[1413]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1413]) );
  DFF \round_reg_reg[1414]  ( .D(out[1414]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1414]) );
  DFF \round_reg_reg[1415]  ( .D(out[1415]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1415]) );
  DFF \round_reg_reg[1416]  ( .D(out[1416]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1416]) );
  DFF \round_reg_reg[1417]  ( .D(out[1417]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1417]) );
  DFF \round_reg_reg[1418]  ( .D(out[1418]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1418]) );
  DFF \round_reg_reg[1419]  ( .D(out[1419]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1419]) );
  DFF \round_reg_reg[1420]  ( .D(out[1420]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1420]) );
  DFF \round_reg_reg[1421]  ( .D(out[1421]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1421]) );
  DFF \round_reg_reg[1422]  ( .D(out[1422]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1422]) );
  DFF \round_reg_reg[1423]  ( .D(out[1423]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1423]) );
  DFF \round_reg_reg[1424]  ( .D(out[1424]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1424]) );
  DFF \round_reg_reg[1425]  ( .D(out[1425]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1425]) );
  DFF \round_reg_reg[1426]  ( .D(out[1426]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1426]) );
  DFF \round_reg_reg[1427]  ( .D(out[1427]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1427]) );
  DFF \round_reg_reg[1428]  ( .D(out[1428]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1428]) );
  DFF \round_reg_reg[1429]  ( .D(out[1429]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1429]) );
  DFF \round_reg_reg[1430]  ( .D(out[1430]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1430]) );
  DFF \round_reg_reg[1431]  ( .D(out[1431]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1431]) );
  DFF \round_reg_reg[1432]  ( .D(out[1432]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1432]) );
  DFF \round_reg_reg[1433]  ( .D(out[1433]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1433]) );
  DFF \round_reg_reg[1434]  ( .D(out[1434]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1434]) );
  DFF \round_reg_reg[1435]  ( .D(out[1435]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1435]) );
  DFF \round_reg_reg[1436]  ( .D(out[1436]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1436]) );
  DFF \round_reg_reg[1437]  ( .D(out[1437]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1437]) );
  DFF \round_reg_reg[1438]  ( .D(out[1438]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1438]) );
  DFF \round_reg_reg[1439]  ( .D(out[1439]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1439]) );
  DFF \round_reg_reg[1440]  ( .D(out[1440]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1440]) );
  DFF \round_reg_reg[1441]  ( .D(out[1441]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1441]) );
  DFF \round_reg_reg[1442]  ( .D(out[1442]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1442]) );
  DFF \round_reg_reg[1443]  ( .D(out[1443]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1443]) );
  DFF \round_reg_reg[1444]  ( .D(out[1444]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1444]) );
  DFF \round_reg_reg[1445]  ( .D(out[1445]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1445]) );
  DFF \round_reg_reg[1446]  ( .D(out[1446]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1446]) );
  DFF \round_reg_reg[1447]  ( .D(out[1447]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1447]) );
  DFF \round_reg_reg[1448]  ( .D(out[1448]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1448]) );
  DFF \round_reg_reg[1449]  ( .D(out[1449]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1449]) );
  DFF \round_reg_reg[1450]  ( .D(out[1450]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1450]) );
  DFF \round_reg_reg[1451]  ( .D(out[1451]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1451]) );
  DFF \round_reg_reg[1452]  ( .D(out[1452]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1452]) );
  DFF \round_reg_reg[1453]  ( .D(out[1453]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1453]) );
  DFF \round_reg_reg[1454]  ( .D(out[1454]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1454]) );
  DFF \round_reg_reg[1455]  ( .D(out[1455]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1455]) );
  DFF \round_reg_reg[1456]  ( .D(out[1456]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1456]) );
  DFF \round_reg_reg[1457]  ( .D(out[1457]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1457]) );
  DFF \round_reg_reg[1458]  ( .D(out[1458]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1458]) );
  DFF \round_reg_reg[1459]  ( .D(out[1459]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1459]) );
  DFF \round_reg_reg[1460]  ( .D(out[1460]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1460]) );
  DFF \round_reg_reg[1461]  ( .D(out[1461]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1461]) );
  DFF \round_reg_reg[1462]  ( .D(out[1462]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1462]) );
  DFF \round_reg_reg[1463]  ( .D(out[1463]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1463]) );
  DFF \round_reg_reg[1464]  ( .D(out[1464]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1464]) );
  DFF \round_reg_reg[1465]  ( .D(out[1465]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1465]) );
  DFF \round_reg_reg[1466]  ( .D(out[1466]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1466]) );
  DFF \round_reg_reg[1467]  ( .D(out[1467]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1467]) );
  DFF \round_reg_reg[1468]  ( .D(out[1468]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1468]) );
  DFF \round_reg_reg[1469]  ( .D(out[1469]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1469]) );
  DFF \round_reg_reg[1470]  ( .D(out[1470]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1470]) );
  DFF \round_reg_reg[1471]  ( .D(out[1471]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1471]) );
  DFF \round_reg_reg[1472]  ( .D(out[1472]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1472]) );
  DFF \round_reg_reg[1473]  ( .D(out[1473]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1473]) );
  DFF \round_reg_reg[1474]  ( .D(out[1474]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1474]) );
  DFF \round_reg_reg[1475]  ( .D(out[1475]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1475]) );
  DFF \round_reg_reg[1476]  ( .D(out[1476]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1476]) );
  DFF \round_reg_reg[1477]  ( .D(out[1477]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1477]) );
  DFF \round_reg_reg[1478]  ( .D(out[1478]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1478]) );
  DFF \round_reg_reg[1479]  ( .D(out[1479]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1479]) );
  DFF \round_reg_reg[1480]  ( .D(out[1480]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1480]) );
  DFF \round_reg_reg[1481]  ( .D(out[1481]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1481]) );
  DFF \round_reg_reg[1482]  ( .D(out[1482]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1482]) );
  DFF \round_reg_reg[1483]  ( .D(out[1483]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1483]) );
  DFF \round_reg_reg[1484]  ( .D(out[1484]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1484]) );
  DFF \round_reg_reg[1485]  ( .D(out[1485]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1485]) );
  DFF \round_reg_reg[1486]  ( .D(out[1486]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1486]) );
  DFF \round_reg_reg[1487]  ( .D(out[1487]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1487]) );
  DFF \round_reg_reg[1488]  ( .D(out[1488]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1488]) );
  DFF \round_reg_reg[1489]  ( .D(out[1489]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1489]) );
  DFF \round_reg_reg[1490]  ( .D(out[1490]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1490]) );
  DFF \round_reg_reg[1491]  ( .D(out[1491]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1491]) );
  DFF \round_reg_reg[1492]  ( .D(out[1492]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1492]) );
  DFF \round_reg_reg[1493]  ( .D(out[1493]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1493]) );
  DFF \round_reg_reg[1494]  ( .D(out[1494]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1494]) );
  DFF \round_reg_reg[1495]  ( .D(out[1495]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1495]) );
  DFF \round_reg_reg[1496]  ( .D(out[1496]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1496]) );
  DFF \round_reg_reg[1497]  ( .D(out[1497]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1497]) );
  DFF \round_reg_reg[1498]  ( .D(out[1498]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1498]) );
  DFF \round_reg_reg[1499]  ( .D(out[1499]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1499]) );
  DFF \round_reg_reg[1500]  ( .D(out[1500]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1500]) );
  DFF \round_reg_reg[1501]  ( .D(out[1501]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1501]) );
  DFF \round_reg_reg[1502]  ( .D(out[1502]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1502]) );
  DFF \round_reg_reg[1503]  ( .D(out[1503]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1503]) );
  DFF \round_reg_reg[1504]  ( .D(out[1504]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1504]) );
  DFF \round_reg_reg[1505]  ( .D(out[1505]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1505]) );
  DFF \round_reg_reg[1506]  ( .D(out[1506]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1506]) );
  DFF \round_reg_reg[1507]  ( .D(out[1507]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1507]) );
  DFF \round_reg_reg[1508]  ( .D(out[1508]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1508]) );
  DFF \round_reg_reg[1509]  ( .D(out[1509]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1509]) );
  DFF \round_reg_reg[1510]  ( .D(out[1510]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1510]) );
  DFF \round_reg_reg[1511]  ( .D(out[1511]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1511]) );
  DFF \round_reg_reg[1512]  ( .D(out[1512]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1512]) );
  DFF \round_reg_reg[1513]  ( .D(out[1513]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1513]) );
  DFF \round_reg_reg[1514]  ( .D(out[1514]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1514]) );
  DFF \round_reg_reg[1515]  ( .D(out[1515]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1515]) );
  DFF \round_reg_reg[1516]  ( .D(out[1516]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1516]) );
  DFF \round_reg_reg[1517]  ( .D(out[1517]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1517]) );
  DFF \round_reg_reg[1518]  ( .D(out[1518]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1518]) );
  DFF \round_reg_reg[1519]  ( .D(out[1519]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1519]) );
  DFF \round_reg_reg[1520]  ( .D(out[1520]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1520]) );
  DFF \round_reg_reg[1521]  ( .D(out[1521]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1521]) );
  DFF \round_reg_reg[1522]  ( .D(out[1522]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1522]) );
  DFF \round_reg_reg[1523]  ( .D(out[1523]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1523]) );
  DFF \round_reg_reg[1524]  ( .D(out[1524]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1524]) );
  DFF \round_reg_reg[1525]  ( .D(out[1525]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1525]) );
  DFF \round_reg_reg[1526]  ( .D(out[1526]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1526]) );
  DFF \round_reg_reg[1527]  ( .D(out[1527]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1527]) );
  DFF \round_reg_reg[1528]  ( .D(out[1528]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1528]) );
  DFF \round_reg_reg[1529]  ( .D(out[1529]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1529]) );
  DFF \round_reg_reg[1530]  ( .D(out[1530]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1530]) );
  DFF \round_reg_reg[1531]  ( .D(out[1531]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1531]) );
  DFF \round_reg_reg[1532]  ( .D(out[1532]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1532]) );
  DFF \round_reg_reg[1533]  ( .D(out[1533]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1533]) );
  DFF \round_reg_reg[1534]  ( .D(out[1534]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1534]) );
  DFF \round_reg_reg[1535]  ( .D(out[1535]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1535]) );
  DFF \round_reg_reg[1536]  ( .D(out[1536]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1536]) );
  DFF \round_reg_reg[1537]  ( .D(out[1537]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1537]) );
  DFF \round_reg_reg[1538]  ( .D(out[1538]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1538]) );
  DFF \round_reg_reg[1539]  ( .D(out[1539]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1539]) );
  DFF \round_reg_reg[1540]  ( .D(out[1540]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1540]) );
  DFF \round_reg_reg[1541]  ( .D(out[1541]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1541]) );
  DFF \round_reg_reg[1542]  ( .D(out[1542]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1542]) );
  DFF \round_reg_reg[1543]  ( .D(out[1543]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1543]) );
  DFF \round_reg_reg[1544]  ( .D(out[1544]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1544]) );
  DFF \round_reg_reg[1545]  ( .D(out[1545]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1545]) );
  DFF \round_reg_reg[1546]  ( .D(out[1546]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1546]) );
  DFF \round_reg_reg[1547]  ( .D(out[1547]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1547]) );
  DFF \round_reg_reg[1548]  ( .D(out[1548]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1548]) );
  DFF \round_reg_reg[1549]  ( .D(out[1549]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1549]) );
  DFF \round_reg_reg[1550]  ( .D(out[1550]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1550]) );
  DFF \round_reg_reg[1551]  ( .D(out[1551]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1551]) );
  DFF \round_reg_reg[1552]  ( .D(out[1552]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1552]) );
  DFF \round_reg_reg[1553]  ( .D(out[1553]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1553]) );
  DFF \round_reg_reg[1554]  ( .D(out[1554]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1554]) );
  DFF \round_reg_reg[1555]  ( .D(out[1555]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1555]) );
  DFF \round_reg_reg[1556]  ( .D(out[1556]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1556]) );
  DFF \round_reg_reg[1557]  ( .D(out[1557]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1557]) );
  DFF \round_reg_reg[1558]  ( .D(out[1558]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1558]) );
  DFF \round_reg_reg[1559]  ( .D(out[1559]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1559]) );
  DFF \round_reg_reg[1560]  ( .D(out[1560]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1560]) );
  DFF \round_reg_reg[1561]  ( .D(out[1561]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1561]) );
  DFF \round_reg_reg[1562]  ( .D(out[1562]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1562]) );
  DFF \round_reg_reg[1563]  ( .D(out[1563]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1563]) );
  DFF \round_reg_reg[1564]  ( .D(out[1564]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1564]) );
  DFF \round_reg_reg[1565]  ( .D(out[1565]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1565]) );
  DFF \round_reg_reg[1566]  ( .D(out[1566]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1566]) );
  DFF \round_reg_reg[1567]  ( .D(out[1567]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1567]) );
  DFF \round_reg_reg[1568]  ( .D(out[1568]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1568]) );
  DFF \round_reg_reg[1569]  ( .D(out[1569]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1569]) );
  DFF \round_reg_reg[1570]  ( .D(out[1570]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1570]) );
  DFF \round_reg_reg[1571]  ( .D(out[1571]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1571]) );
  DFF \round_reg_reg[1572]  ( .D(out[1572]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1572]) );
  DFF \round_reg_reg[1573]  ( .D(out[1573]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1573]) );
  DFF \round_reg_reg[1574]  ( .D(out[1574]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1574]) );
  DFF \round_reg_reg[1575]  ( .D(out[1575]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1575]) );
  DFF \round_reg_reg[1576]  ( .D(out[1576]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1576]) );
  DFF \round_reg_reg[1577]  ( .D(out[1577]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1577]) );
  DFF \round_reg_reg[1578]  ( .D(out[1578]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1578]) );
  DFF \round_reg_reg[1579]  ( .D(out[1579]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1579]) );
  DFF \round_reg_reg[1580]  ( .D(out[1580]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1580]) );
  DFF \round_reg_reg[1581]  ( .D(out[1581]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1581]) );
  DFF \round_reg_reg[1582]  ( .D(out[1582]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1582]) );
  DFF \round_reg_reg[1583]  ( .D(out[1583]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1583]) );
  DFF \round_reg_reg[1584]  ( .D(out[1584]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1584]) );
  DFF \round_reg_reg[1585]  ( .D(out[1585]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1585]) );
  DFF \round_reg_reg[1586]  ( .D(out[1586]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1586]) );
  DFF \round_reg_reg[1587]  ( .D(out[1587]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1587]) );
  DFF \round_reg_reg[1588]  ( .D(out[1588]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1588]) );
  DFF \round_reg_reg[1589]  ( .D(out[1589]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1589]) );
  DFF \round_reg_reg[1590]  ( .D(out[1590]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1590]) );
  DFF \round_reg_reg[1591]  ( .D(out[1591]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1591]) );
  DFF \round_reg_reg[1592]  ( .D(out[1592]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1592]) );
  DFF \round_reg_reg[1593]  ( .D(out[1593]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1593]) );
  DFF \round_reg_reg[1594]  ( .D(out[1594]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1594]) );
  DFF \round_reg_reg[1595]  ( .D(out[1595]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1595]) );
  DFF \round_reg_reg[1596]  ( .D(out[1596]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1596]) );
  DFF \round_reg_reg[1597]  ( .D(out[1597]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1597]) );
  DFF \round_reg_reg[1598]  ( .D(out[1598]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1598]) );
  DFF \round_reg_reg[1599]  ( .D(out[1599]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1599]) );
  NOR U1035 ( .A(n21578), .B(n21576), .Z(n24768) );
  ANDN U1036 ( .B(n22194), .A(n22195), .Z(n22192) );
  ANDN U1037 ( .B(n21277), .A(n20815), .Z(n21276) );
  NOR U1038 ( .A(n22992), .B(n19766), .Z(n24574) );
  XNOR U1039 ( .A(n19790), .B(n26209), .Z(n15907) );
  ANDN U1040 ( .B(n20950), .A(n20952), .Z(n25158) );
  NOR U1041 ( .A(n21819), .B(n21818), .Z(n21816) );
  XNOR U1042 ( .A(n19457), .B(n18690), .Z(n14918) );
  XNOR U1043 ( .A(n23183), .B(n20310), .Z(n18121) );
  XOR U1044 ( .A(n13395), .B(n17748), .Z(n9768) );
  XOR U1045 ( .A(n6247), .B(n9439), .Z(n1738) );
  XOR U1046 ( .A(n26039), .B(n25251), .Z(n23621) );
  XNOR U1047 ( .A(n25161), .B(n25160), .Z(n21923) );
  XNOR U1048 ( .A(n25598), .B(n25777), .Z(n22372) );
  XNOR U1049 ( .A(n24817), .B(n25253), .Z(n23471) );
  XNOR U1050 ( .A(round_reg[305]), .B(n22962), .Z(n21590) );
  ANDN U1051 ( .B(n23898), .A(n20705), .Z(n23897) );
  NOR U1052 ( .A(n22661), .B(n22662), .Z(n24914) );
  ANDN U1053 ( .B(n19951), .A(n19949), .Z(n20623) );
  XNOR U1054 ( .A(n20580), .B(n20579), .Z(n16674) );
  ANDN U1055 ( .B(n21694), .A(n21695), .Z(n21692) );
  ANDN U1056 ( .B(n21853), .A(n24647), .Z(n24646) );
  NOR U1057 ( .A(n19675), .B(n19676), .Z(n20381) );
  NOR U1058 ( .A(n24177), .B(n22564), .Z(n24432) );
  ANDN U1059 ( .B(n22625), .A(n22758), .Z(n24713) );
  NOR U1060 ( .A(n21680), .B(n22967), .Z(n22965) );
  NOR U1061 ( .A(n19885), .B(n19887), .Z(n20572) );
  XOR U1062 ( .A(n24890), .B(n23183), .Z(n18789) );
  NOR U1063 ( .A(n23972), .B(n22246), .Z(n23971) );
  NOR U1064 ( .A(n22073), .B(n21689), .Z(n24579) );
  NOR U1065 ( .A(n24625), .B(n24624), .Z(n24623) );
  XNOR U1066 ( .A(n24869), .B(n23195), .Z(n18404) );
  XNOR U1067 ( .A(n21824), .B(n18912), .Z(n15591) );
  XOR U1068 ( .A(n18453), .B(n20135), .Z(n17483) );
  NOR U1069 ( .A(n13995), .B(n13996), .Z(n15897) );
  XNOR U1070 ( .A(n15771), .B(n15772), .Z(n11857) );
  ANDN U1071 ( .B(n14360), .A(n14361), .Z(n14358) );
  ANDN U1072 ( .B(n13147), .A(n13145), .Z(n17971) );
  ANDN U1073 ( .B(n14322), .A(n14323), .Z(n14320) );
  ANDN U1074 ( .B(n14745), .A(n14747), .Z(n16314) );
  ANDN U1075 ( .B(n14732), .A(n14733), .Z(n14730) );
  NOR U1076 ( .A(n16160), .B(n14677), .Z(n16661) );
  NOR U1077 ( .A(n15095), .B(n17161), .Z(n21279) );
  ANDN U1078 ( .B(n13678), .A(n13679), .Z(n13676) );
  NOR U1079 ( .A(n14068), .B(n14067), .Z(n14065) );
  NOR U1080 ( .A(n15073), .B(n15074), .Z(n18600) );
  XOR U1081 ( .A(n16127), .B(n16126), .Z(n10691) );
  XNOR U1082 ( .A(n12077), .B(n12076), .Z(n9784) );
  XNOR U1083 ( .A(n6273), .B(n6358), .Z(n5128) );
  ANDN U1084 ( .B(n9150), .A(n7927), .Z(n9235) );
  XNOR U1085 ( .A(n6172), .B(n8179), .Z(n1965) );
  XOR U1086 ( .A(n6163), .B(n8125), .Z(n1961) );
  ANDN U1087 ( .B(n4926), .A(n4732), .Z(n4923) );
  NOR U1088 ( .A(n4409), .B(n4866), .Z(n5089) );
  ANDN U1089 ( .B(n5615), .A(n6124), .Z(n6714) );
  XNOR U1090 ( .A(n25409), .B(n25031), .Z(n24906) );
  XNOR U1091 ( .A(n25119), .B(n25118), .Z(n23134) );
  XNOR U1092 ( .A(n24942), .B(n24941), .Z(n24727) );
  XNOR U1093 ( .A(n25127), .B(n25126), .Z(n23300) );
  XNOR U1094 ( .A(round_reg[189]), .B(n21609), .Z(n19925) );
  XOR U1095 ( .A(round_reg[169]), .B(n22372), .Z(n22328) );
  XNOR U1096 ( .A(round_reg[158]), .B(n21923), .Z(n20787) );
  XNOR U1097 ( .A(round_reg[754]), .B(n23197), .Z(n20653) );
  XOR U1098 ( .A(round_reg[835]), .B(n24697), .Z(n22875) );
  ANDN U1099 ( .B(n23707), .A(n21058), .Z(n23705) );
  NOR U1100 ( .A(n23716), .B(n21651), .Z(n24314) );
  XNOR U1101 ( .A(n22392), .B(n22393), .Z(n16759) );
  ANDN U1102 ( .B(n22447), .A(n23003), .Z(n23404) );
  ANDN U1103 ( .B(n23113), .A(n23112), .Z(n25500) );
  NOR U1104 ( .A(n20317), .B(n20458), .Z(n21308) );
  NOR U1105 ( .A(n20773), .B(n19830), .Z(n20772) );
  NOR U1106 ( .A(n20442), .B(n20441), .Z(n20439) );
  NOR U1107 ( .A(n20254), .B(n20253), .Z(n20251) );
  ANDN U1108 ( .B(n22035), .A(n19750), .Z(n22985) );
  XNOR U1109 ( .A(n19626), .B(n19625), .Z(n15597) );
  ANDN U1110 ( .B(n20511), .A(n20512), .Z(n20509) );
  ANDN U1111 ( .B(n22963), .A(n22075), .Z(n22961) );
  NOR U1112 ( .A(n21921), .B(n20543), .Z(n24537) );
  ANDN U1113 ( .B(n20906), .A(n20907), .Z(n20904) );
  NOR U1114 ( .A(n20299), .B(n20298), .Z(n20296) );
  XOR U1115 ( .A(n21574), .B(n20580), .Z(n17137) );
  NOR U1116 ( .A(n20390), .B(n20161), .Z(n22817) );
  NOR U1117 ( .A(n20222), .B(n21203), .Z(n21202) );
  NOR U1118 ( .A(n19807), .B(n19946), .Z(n21184) );
  ANDN U1119 ( .B(n20182), .A(n20702), .Z(n23985) );
  NOR U1120 ( .A(n20174), .B(n21232), .Z(n23903) );
  NOR U1121 ( .A(n21403), .B(n21404), .Z(n25371) );
  NOR U1122 ( .A(n22464), .B(n22465), .Z(n25947) );
  XNOR U1123 ( .A(n18749), .B(n18748), .Z(n15623) );
  NOR U1124 ( .A(n21969), .B(n22046), .Z(n24129) );
  ANDN U1125 ( .B(n23536), .A(n20880), .Z(n23535) );
  ANDN U1126 ( .B(n19753), .A(n20832), .Z(n24563) );
  XNOR U1127 ( .A(n19537), .B(n19536), .Z(n19291) );
  ANDN U1128 ( .B(n22546), .A(n22547), .Z(n22544) );
  XOR U1129 ( .A(n23331), .B(n23330), .Z(n16746) );
  XNOR U1130 ( .A(n19708), .B(n19707), .Z(n16543) );
  XOR U1131 ( .A(n17553), .B(n17552), .Z(n15465) );
  XOR U1132 ( .A(n15207), .B(n15208), .Z(n13106) );
  XNOR U1133 ( .A(n17220), .B(n19220), .Z(n14791) );
  XOR U1134 ( .A(n17192), .B(n18623), .Z(n16742) );
  XNOR U1135 ( .A(n15590), .B(n15591), .Z(n14417) );
  XOR U1136 ( .A(n20945), .B(n16476), .Z(n12378) );
  XNOR U1137 ( .A(n14918), .B(n18206), .Z(n15791) );
  ANDN U1138 ( .B(n15115), .A(n15113), .Z(n23922) );
  NOR U1139 ( .A(n17099), .B(n17100), .Z(n18050) );
  NOR U1140 ( .A(n12499), .B(n12500), .Z(n13565) );
  XNOR U1141 ( .A(n16636), .B(n15100), .Z(n10574) );
  ANDN U1142 ( .B(n12748), .A(n12749), .Z(n12746) );
  ANDN U1143 ( .B(n17756), .A(n17757), .Z(n17754) );
  NOR U1144 ( .A(n15215), .B(n14466), .Z(n17537) );
  ANDN U1145 ( .B(n14151), .A(n15758), .Z(n20201) );
  ANDN U1146 ( .B(n12903), .A(n14109), .Z(n16012) );
  NOR U1147 ( .A(n13825), .B(n14689), .Z(n18834) );
  NOR U1148 ( .A(n14190), .B(n14189), .Z(n14187) );
  NOR U1149 ( .A(n13633), .B(n13632), .Z(n13630) );
  NOR U1150 ( .A(n16359), .B(n15552), .Z(n16358) );
  NOR U1151 ( .A(n14441), .B(n16619), .Z(n16617) );
  ANDN U1152 ( .B(n15745), .A(n15746), .Z(n15743) );
  ANDN U1153 ( .B(n16439), .A(n16542), .Z(n19655) );
  NOR U1154 ( .A(n15692), .B(n14703), .Z(n15689) );
  ANDN U1155 ( .B(n11952), .A(n11951), .Z(n16301) );
  NOR U1156 ( .A(n16979), .B(n17008), .Z(n17005) );
  NOR U1157 ( .A(n13997), .B(n17955), .Z(n17975) );
  XNOR U1158 ( .A(n17298), .B(n17297), .Z(n10113) );
  XNOR U1159 ( .A(n10673), .B(n14031), .Z(n13115) );
  ANDN U1160 ( .B(n16662), .A(n14679), .Z(n25099) );
  NOR U1161 ( .A(n16388), .B(n16870), .Z(n17347) );
  ANDN U1162 ( .B(n15103), .A(n16630), .Z(n23508) );
  XNOR U1163 ( .A(n12682), .B(n11456), .Z(n11218) );
  ANDN U1164 ( .B(n8015), .A(n8013), .Z(n9055) );
  ANDN U1165 ( .B(n10508), .A(n10507), .Z(n11654) );
  ANDN U1166 ( .B(n10858), .A(n10857), .Z(n12292) );
  NOR U1167 ( .A(n6896), .B(n6895), .Z(n6894) );
  ANDN U1168 ( .B(n7622), .A(n7620), .Z(n11136) );
  ANDN U1169 ( .B(n6393), .A(n6394), .Z(n6391) );
  ANDN U1170 ( .B(n8697), .A(n12218), .Z(n12386) );
  XNOR U1171 ( .A(n10413), .B(n10414), .Z(n7528) );
  ANDN U1172 ( .B(n7733), .A(n10319), .Z(n10511) );
  NOR U1173 ( .A(n11225), .B(n11226), .Z(n12982) );
  NOR U1174 ( .A(n8341), .B(n9746), .Z(n9744) );
  NOR U1175 ( .A(n7850), .B(n7849), .Z(n8914) );
  NOR U1176 ( .A(n8712), .B(n8635), .Z(n8711) );
  XNOR U1177 ( .A(n7874), .B(n7875), .Z(n2445) );
  XOR U1178 ( .A(n6231), .B(n9029), .Z(n1720) );
  XOR U1179 ( .A(n6255), .B(n9649), .Z(n1747) );
  XNOR U1180 ( .A(n3826), .B(n2252), .Z(n2909) );
  XOR U1181 ( .A(n2477), .B(n4264), .Z(n1668) );
  ANDN U1182 ( .B(n4470), .A(n4471), .Z(n4468) );
  ANDN U1183 ( .B(n4547), .A(n4548), .Z(n4545) );
  ANDN U1184 ( .B(n4580), .A(n4581), .Z(n4578) );
  NOR U1185 ( .A(n4707), .B(n4442), .Z(n4706) );
  NOR U1186 ( .A(n4860), .B(n4682), .Z(n4857) );
  ANDN U1187 ( .B(n4919), .A(n4723), .Z(n4917) );
  ANDN U1188 ( .B(n4922), .A(n4730), .Z(n4920) );
  ANDN U1189 ( .B(n4629), .A(n5042), .Z(n5233) );
  ANDN U1190 ( .B(n5752), .A(n1196), .Z(n5751) );
  ANDN U1191 ( .B(n1055), .A(n1056), .Z(n1053) );
  ANDN U1192 ( .B(n1283), .A(n1284), .Z(n1281) );
  ANDN U1193 ( .B(n1320), .A(n1321), .Z(n1318) );
  ANDN U1194 ( .B(n1546), .A(n1287), .Z(n1545) );
  ANDN U1195 ( .B(n1561), .A(n1324), .Z(n1560) );
  NOR U1196 ( .A(n1704), .B(n1527), .Z(n1701) );
  XOR U1197 ( .A(n25306), .B(n25409), .Z(n24779) );
  XNOR U1198 ( .A(n25094), .B(n25093), .Z(n24996) );
  XOR U1199 ( .A(n25895), .B(n26215), .Z(n22230) );
  XNOR U1200 ( .A(n25207), .B(n25206), .Z(n23019) );
  XNOR U1201 ( .A(n25087), .B(n25195), .Z(n22272) );
  XNOR U1202 ( .A(n25287), .B(n25342), .Z(n25029) );
  XNOR U1203 ( .A(n25438), .B(n25696), .Z(n22649) );
  XNOR U1204 ( .A(n25843), .B(n25442), .Z(n23318) );
  XOR U1205 ( .A(n24735), .B(n24328), .Z(n23785) );
  XNOR U1206 ( .A(n25358), .B(n25330), .Z(n23016) );
  XNOR U1207 ( .A(n25440), .B(n25201), .Z(n23584) );
  XOR U1208 ( .A(round_reg[878]), .B(n23735), .Z(n22496) );
  XNOR U1209 ( .A(round_reg[250]), .B(n23249), .Z(n21817) );
  XOR U1210 ( .A(round_reg[409]), .B(n21760), .Z(n20216) );
  ANDN U1211 ( .B(n22847), .A(n20892), .Z(n24105) );
  NOR U1212 ( .A(n20535), .B(n21288), .Z(n21287) );
  NOR U1213 ( .A(n21045), .B(n20559), .Z(n24546) );
  ANDN U1214 ( .B(n21180), .A(n21178), .Z(n23513) );
  ANDN U1215 ( .B(n21740), .A(n21739), .Z(n24403) );
  ANDN U1216 ( .B(n19274), .A(n19275), .Z(n19272) );
  NOR U1217 ( .A(n19843), .B(n19844), .Z(n19924) );
  NOR U1218 ( .A(n21685), .B(n21684), .Z(n21682) );
  ANDN U1219 ( .B(n22500), .A(n24630), .Z(n24628) );
  XOR U1220 ( .A(n22355), .B(n21574), .Z(n17363) );
  NOR U1221 ( .A(n21533), .B(n23579), .Z(n24755) );
  ANDN U1222 ( .B(n20010), .A(n20008), .Z(n23620) );
  NOR U1223 ( .A(n20419), .B(n20144), .Z(n22815) );
  ANDN U1224 ( .B(n23710), .A(n23711), .Z(n23708) );
  NOR U1225 ( .A(n22300), .B(n22299), .Z(n22297) );
  NOR U1226 ( .A(n22125), .B(n22124), .Z(n22122) );
  NOR U1227 ( .A(n22674), .B(n22675), .Z(n24915) );
  XNOR U1228 ( .A(n20282), .B(n20281), .Z(n17389) );
  NOR U1229 ( .A(n21228), .B(n21227), .Z(n21226) );
  NOR U1230 ( .A(n21147), .B(n21148), .Z(n23530) );
  NOR U1231 ( .A(n22726), .B(n22727), .Z(n23071) );
  NOR U1232 ( .A(n20118), .B(n20117), .Z(n20116) );
  XNOR U1233 ( .A(n19528), .B(n18452), .Z(n17517) );
  XNOR U1234 ( .A(n19499), .B(n19498), .Z(n18824) );
  ANDN U1235 ( .B(n19510), .A(n21946), .Z(n23468) );
  ANDN U1236 ( .B(n20176), .A(n20700), .Z(n23990) );
  ANDN U1237 ( .B(n20815), .A(n20816), .Z(n20813) );
  XNOR U1238 ( .A(n25221), .B(n20520), .Z(n19342) );
  NOR U1239 ( .A(n24785), .B(n23821), .Z(n24786) );
  NOR U1240 ( .A(n20485), .B(n20484), .Z(n20482) );
  ANDN U1241 ( .B(n19468), .A(n19730), .Z(n19728) );
  ANDN U1242 ( .B(n22548), .A(n24428), .Z(n24434) );
  ANDN U1243 ( .B(n21337), .A(n21239), .Z(n23010) );
  NOR U1244 ( .A(n22329), .B(n22328), .Z(n22327) );
  XNOR U1245 ( .A(n21126), .B(n18329), .Z(n15615) );
  ANDN U1246 ( .B(n21153), .A(n22170), .Z(n25258) );
  XNOR U1247 ( .A(n19176), .B(n19175), .Z(n18904) );
  XOR U1248 ( .A(n19328), .B(n19327), .Z(n18473) );
  NOR U1249 ( .A(n21743), .B(n21744), .Z(n24032) );
  XNOR U1250 ( .A(n22586), .B(n22585), .Z(n18379) );
  XNOR U1251 ( .A(n19653), .B(n20444), .Z(n16934) );
  XOR U1252 ( .A(n20237), .B(n20236), .Z(n17469) );
  XNOR U1253 ( .A(n19718), .B(n18599), .Z(n18625) );
  ANDN U1254 ( .B(n19949), .A(n20624), .Z(n21187) );
  XNOR U1255 ( .A(n22653), .B(n18748), .Z(n19732) );
  NOR U1256 ( .A(n21400), .B(n21401), .Z(n25353) );
  XNOR U1257 ( .A(n20514), .B(n20463), .Z(n17472) );
  XNOR U1258 ( .A(n19637), .B(n19636), .Z(n16021) );
  NOR U1259 ( .A(n19828), .B(n20506), .Z(n20505) );
  XNOR U1260 ( .A(n22503), .B(n19906), .Z(n16465) );
  XNOR U1261 ( .A(n20011), .B(n19625), .Z(n17895) );
  XNOR U1262 ( .A(n18913), .B(n18912), .Z(n17458) );
  XNOR U1263 ( .A(n19307), .B(n17474), .Z(n14047) );
  XOR U1264 ( .A(n16054), .B(n16055), .Z(n15350) );
  XNOR U1265 ( .A(n17466), .B(n17467), .Z(n13664) );
  XOR U1266 ( .A(n22628), .B(n17439), .Z(n14790) );
  NOR U1267 ( .A(n17125), .B(n13495), .Z(n18184) );
  NOR U1268 ( .A(n14272), .B(n14273), .Z(n15624) );
  NOR U1269 ( .A(n17094), .B(n18664), .Z(n18661) );
  NOR U1270 ( .A(n14038), .B(n14037), .Z(n14035) );
  NOR U1271 ( .A(n13716), .B(n14559), .Z(n14558) );
  NOR U1272 ( .A(n15448), .B(n15449), .Z(n20394) );
  ANDN U1273 ( .B(n16718), .A(n15926), .Z(n17037) );
  ANDN U1274 ( .B(n13503), .A(n13504), .Z(n13501) );
  NOR U1275 ( .A(n13743), .B(n15847), .Z(n15845) );
  ANDN U1276 ( .B(n17649), .A(n15674), .Z(n18635) );
  NOR U1277 ( .A(n14574), .B(n15156), .Z(n24365) );
  ANDN U1278 ( .B(n13302), .A(n16158), .Z(n16166) );
  ANDN U1279 ( .B(n14769), .A(n14767), .Z(n16350) );
  ANDN U1280 ( .B(n12758), .A(n12757), .Z(n13461) );
  ANDN U1281 ( .B(n16810), .A(n14746), .Z(n18428) );
  ANDN U1282 ( .B(n11957), .A(n11956), .Z(n16295) );
  NOR U1283 ( .A(n13763), .B(n13762), .Z(n13760) );
  XNOR U1284 ( .A(n13512), .B(n13511), .Z(n9944) );
  XNOR U1285 ( .A(n16415), .B(n15530), .Z(n14429) );
  NOR U1286 ( .A(n14233), .B(n14232), .Z(n18893) );
  ANDN U1287 ( .B(n14475), .A(n15458), .Z(n16278) );
  ANDN U1288 ( .B(n15027), .A(n15028), .Z(n15025) );
  XNOR U1289 ( .A(n11525), .B(n13226), .Z(n10661) );
  ANDN U1290 ( .B(n15497), .A(n15498), .Z(n15495) );
  ANDN U1291 ( .B(n14577), .A(n16439), .Z(n16541) );
  XNOR U1292 ( .A(n18838), .B(n13834), .Z(n11697) );
  ANDN U1293 ( .B(n12301), .A(n12302), .Z(n12299) );
  ANDN U1294 ( .B(n15734), .A(n15735), .Z(n15732) );
  XNOR U1295 ( .A(n13376), .B(n12611), .Z(n10000) );
  NOR U1296 ( .A(n17769), .B(n17768), .Z(n17767) );
  XNOR U1297 ( .A(n17279), .B(n11965), .Z(n13071) );
  NOR U1298 ( .A(n14333), .B(n14332), .Z(n17409) );
  ANDN U1299 ( .B(n15250), .A(n12972), .Z(n15247) );
  NOR U1300 ( .A(n15111), .B(n15110), .Z(n15108) );
  NOR U1301 ( .A(n16566), .B(n16565), .Z(n16563) );
  XNOR U1302 ( .A(n11278), .B(n14546), .Z(n10830) );
  NOR U1303 ( .A(n12908), .B(n14117), .Z(n16007) );
  NOR U1304 ( .A(n13194), .B(n13195), .Z(n13573) );
  XNOR U1305 ( .A(n16629), .B(n15104), .Z(n11744) );
  ANDN U1306 ( .B(n15776), .A(n14862), .Z(n18540) );
  XNOR U1307 ( .A(n11943), .B(n11849), .Z(n12205) );
  XNOR U1308 ( .A(n11930), .B(n13878), .Z(n9168) );
  XNOR U1309 ( .A(n9537), .B(n11671), .Z(n10495) );
  XOR U1310 ( .A(n13936), .B(n12050), .Z(n8359) );
  XOR U1311 ( .A(n11923), .B(n9784), .Z(n7415) );
  XOR U1312 ( .A(n10919), .B(n10920), .Z(n9851) );
  XOR U1313 ( .A(n11057), .B(n10544), .Z(n7059) );
  ANDN U1314 ( .B(n8026), .A(n8027), .Z(n8025) );
  ANDN U1315 ( .B(n10749), .A(n10748), .Z(n12143) );
  ANDN U1316 ( .B(n7215), .A(n7216), .Z(n7213) );
  ANDN U1317 ( .B(n7647), .A(n7648), .Z(n7645) );
  ANDN U1318 ( .B(n8794), .A(n12615), .Z(n12839) );
  NOR U1319 ( .A(n9034), .B(n9033), .Z(n9031) );
  ANDN U1320 ( .B(n9225), .A(n9226), .Z(n9223) );
  NOR U1321 ( .A(n10639), .B(n7316), .Z(n10786) );
  ANDN U1322 ( .B(n11094), .A(n11095), .Z(n12708) );
  XNOR U1323 ( .A(n6295), .B(n6494), .Z(n5148) );
  ANDN U1324 ( .B(n7867), .A(n10615), .Z(n10760) );
  ANDN U1325 ( .B(n8434), .A(n8435), .Z(n8432) );
  NOR U1326 ( .A(n7025), .B(n6568), .Z(n9025) );
  ANDN U1327 ( .B(n7207), .A(n7206), .Z(n8294) );
  NOR U1328 ( .A(n7640), .B(n7638), .Z(n8723) );
  NOR U1329 ( .A(n8009), .B(n8011), .Z(n9057) );
  XNOR U1330 ( .A(n7440), .B(n6181), .Z(n2364) );
  ANDN U1331 ( .B(n8197), .A(n8198), .Z(n8195) );
  ANDN U1332 ( .B(n7033), .A(n7034), .Z(n7032) );
  NOR U1333 ( .A(n9725), .B(n9726), .Z(n11839) );
  ANDN U1334 ( .B(n8851), .A(n8934), .Z(n8933) );
  ANDN U1335 ( .B(n8782), .A(n10327), .Z(n10516) );
  NOR U1336 ( .A(n12022), .B(n8413), .Z(n12020) );
  XNOR U1337 ( .A(n6182), .B(n8289), .Z(n1664) );
  XNOR U1338 ( .A(n5942), .B(n5941), .Z(n3743) );
  ANDN U1339 ( .B(n7253), .A(n7254), .Z(n7251) );
  ANDN U1340 ( .B(n11221), .A(n11220), .Z(n12966) );
  ANDN U1341 ( .B(n6846), .A(n6848), .Z(n7583) );
  ANDN U1342 ( .B(n7716), .A(n7717), .Z(n7714) );
  XOR U1343 ( .A(n8969), .B(n8968), .Z(n2455) );
  XNOR U1344 ( .A(n2107), .B(n5850), .Z(n1056) );
  ANDN U1345 ( .B(n4366), .A(n4367), .Z(n4362) );
  ANDN U1346 ( .B(n4370), .A(n4371), .Z(n4368) );
  ANDN U1347 ( .B(n4598), .A(n4599), .Z(n4596) );
  ANDN U1348 ( .B(n4622), .A(n4623), .Z(n4620) );
  ANDN U1349 ( .B(n4930), .A(n4734), .Z(n4927) );
  ANDN U1350 ( .B(n5560), .A(n5561), .Z(n5558) );
  ANDN U1351 ( .B(n5568), .A(n5569), .Z(n5566) );
  ANDN U1352 ( .B(n5653), .A(n5654), .Z(n5651) );
  NOR U1353 ( .A(n5863), .B(n5674), .Z(n5859) );
  NOR U1354 ( .A(n6173), .B(n5826), .Z(n6169) );
  ANDN U1355 ( .B(n6178), .A(n5828), .Z(n6174) );
  NOR U1356 ( .A(n5883), .B(n1078), .Z(n6219) );
  ANDN U1357 ( .B(n1271), .A(n1272), .Z(n1269) );
  XNOR U1358 ( .A(n1293), .B(n1294), .Z(out[941]) );
  ANDN U1359 ( .B(n1360), .A(n1361), .Z(n1358) );
  ANDN U1360 ( .B(n1364), .A(n1365), .Z(n1362) );
  ANDN U1361 ( .B(n1463), .A(n1464), .Z(n1461) );
  ANDN U1362 ( .B(n1495), .A(n1496), .Z(n1493) );
  NOR U1363 ( .A(n1283), .B(n1735), .Z(n1539) );
  ANDN U1364 ( .B(n1556), .A(n1312), .Z(n1555) );
  ANDN U1365 ( .B(n1608), .A(n1408), .Z(n1607) );
  ANDN U1366 ( .B(n1632), .A(n1452), .Z(n1631) );
  ANDN U1367 ( .B(n1636), .A(n1460), .Z(n1635) );
  ANDN U1368 ( .B(n1657), .A(n1500), .Z(n1656) );
  ANDN U1369 ( .B(n1739), .A(n1546), .Z(n1736) );
  ANDN U1370 ( .B(n1704), .A(n1254), .Z(n1998) );
  NOR U1371 ( .A(n1708), .B(n1262), .Z(n2001) );
  NOR U1372 ( .A(n2832), .B(n2831), .Z(n2829) );
  ANDN U1373 ( .B(n3072), .A(n2873), .Z(n3071) );
  ANDN U1374 ( .B(n3286), .A(n2864), .Z(n3494) );
  NOR U1375 ( .A(n3911), .B(n3170), .Z(n3910) );
  ANDN U1376 ( .B(n4043), .A(n2224), .Z(n4041) );
  XOR U1377 ( .A(n25391), .B(n26066), .Z(n24285) );
  XOR U1378 ( .A(n24911), .B(n24933), .Z(n23991) );
  XNOR U1379 ( .A(n24929), .B(n24941), .Z(n24284) );
  XOR U1380 ( .A(n25045), .B(n26094), .Z(n25233) );
  XNOR U1381 ( .A(n24970), .B(n25976), .Z(n23464) );
  XNOR U1382 ( .A(n25378), .B(n25354), .Z(n21617) );
  XNOR U1383 ( .A(n25943), .B(n25998), .Z(n24305) );
  XNOR U1384 ( .A(n25317), .B(n24967), .Z(n24443) );
  XNOR U1385 ( .A(n26298), .B(n25744), .Z(n23865) );
  XNOR U1386 ( .A(n25185), .B(n25211), .Z(n24157) );
  XNOR U1387 ( .A(n24974), .B(n24973), .Z(n21306) );
  XNOR U1388 ( .A(n24822), .B(n24821), .Z(n22764) );
  XNOR U1389 ( .A(n25882), .B(n25904), .Z(n21763) );
  XOR U1390 ( .A(n24725), .B(n25027), .Z(n23011) );
  XNOR U1391 ( .A(n25818), .B(n25206), .Z(n22268) );
  XOR U1392 ( .A(round_reg[235]), .B(n22112), .Z(n19817) );
  XNOR U1393 ( .A(round_reg[1498]), .B(n23471), .Z(n21294) );
  XOR U1394 ( .A(round_reg[697]), .B(n23469), .Z(n20991) );
  XNOR U1395 ( .A(round_reg[436]), .B(n23289), .Z(n22666) );
  XOR U1396 ( .A(round_reg[1286]), .B(n23738), .Z(n21028) );
  XOR U1397 ( .A(round_reg[535]), .B(n24139), .Z(n20253) );
  XOR U1398 ( .A(round_reg[1333]), .B(n21313), .Z(n20744) );
  XOR U1399 ( .A(round_reg[1533]), .B(n23387), .Z(n22020) );
  ANDN U1400 ( .B(n19361), .A(n19362), .Z(n19359) );
  NOR U1401 ( .A(n22611), .B(n22609), .Z(n24641) );
  NOR U1402 ( .A(n21069), .B(n21070), .Z(n24696) );
  ANDN U1403 ( .B(n20367), .A(n20368), .Z(n24295) );
  ANDN U1404 ( .B(n23690), .A(n23691), .Z(n24073) );
  NOR U1405 ( .A(n20731), .B(n21761), .Z(n21759) );
  ANDN U1406 ( .B(n21119), .A(n21120), .Z(n21117) );
  NOR U1407 ( .A(n22529), .B(n24362), .Z(n26404) );
  XNOR U1408 ( .A(n19689), .B(n19688), .Z(n18505) );
  NOR U1409 ( .A(n22903), .B(n22902), .Z(n22901) );
  NOR U1410 ( .A(n22722), .B(n22723), .Z(n23076) );
  NOR U1411 ( .A(n22474), .B(n22475), .Z(n25980) );
  ANDN U1412 ( .B(n22411), .A(n22086), .Z(n24666) );
  ANDN U1413 ( .B(n21167), .A(n21165), .Z(n23516) );
  ANDN U1414 ( .B(n19804), .A(n19802), .Z(n24160) );
  ANDN U1415 ( .B(n19513), .A(n19512), .Z(n22454) );
  ANDN U1416 ( .B(n23165), .A(n21346), .Z(n23594) );
  NOR U1417 ( .A(n18841), .B(n18842), .Z(n20380) );
  ANDN U1418 ( .B(n19874), .A(n19872), .Z(n25752) );
  ANDN U1419 ( .B(n20305), .A(n20306), .Z(n25117) );
  ANDN U1420 ( .B(n22013), .A(n22012), .Z(n22639) );
  NOR U1421 ( .A(n23970), .B(n23969), .Z(n23968) );
  NOR U1422 ( .A(n20294), .B(n20293), .Z(n20291) );
  ANDN U1423 ( .B(n22181), .A(n22182), .Z(n22179) );
  XNOR U1424 ( .A(n19249), .B(n20568), .Z(n14951) );
  ANDN U1425 ( .B(n21297), .A(n20787), .Z(n21296) );
  ANDN U1426 ( .B(n21733), .A(n21732), .Z(n24394) );
  ANDN U1427 ( .B(n21359), .A(n21360), .Z(n21357) );
  ANDN U1428 ( .B(n23548), .A(n23724), .Z(n23723) );
  ANDN U1429 ( .B(n23772), .A(n24830), .Z(n24829) );
  ANDN U1430 ( .B(n21679), .A(n22064), .Z(n25142) );
  ANDN U1431 ( .B(n19763), .A(n19764), .Z(n19761) );
  XNOR U1432 ( .A(n23764), .B(n22168), .Z(n16348) );
  XNOR U1433 ( .A(n20943), .B(n20508), .Z(n20770) );
  XNOR U1434 ( .A(n22238), .B(n23627), .Z(n17876) );
  ANDN U1435 ( .B(n19807), .A(n19808), .Z(n19805) );
  ANDN U1436 ( .B(n20351), .A(n22009), .Z(n23875) );
  ANDN U1437 ( .B(n21254), .A(n23020), .Z(n23585) );
  XOR U1438 ( .A(n18285), .B(n18284), .Z(n13896) );
  ANDN U1439 ( .B(n20962), .A(n20963), .Z(n20960) );
  ANDN U1440 ( .B(n20899), .A(n20897), .Z(n24766) );
  XNOR U1441 ( .A(n20807), .B(n18885), .Z(n16041) );
  NOR U1442 ( .A(n24179), .B(n22560), .Z(n24435) );
  XNOR U1443 ( .A(n21795), .B(n21794), .Z(n18510) );
  XNOR U1444 ( .A(n20709), .B(n19560), .Z(n16062) );
  NOR U1445 ( .A(n22135), .B(n22134), .Z(n22132) );
  NOR U1446 ( .A(n21691), .B(n22960), .Z(n22958) );
  ANDN U1447 ( .B(n20917), .A(n20916), .Z(n22373) );
  NOR U1448 ( .A(n21302), .B(n20454), .Z(n21300) );
  NOR U1449 ( .A(n22744), .B(n23346), .Z(n24016) );
  ANDN U1450 ( .B(n21087), .A(n21525), .Z(n21524) );
  ANDN U1451 ( .B(n21002), .A(n23106), .Z(n25503) );
  XNOR U1452 ( .A(n21636), .B(n20828), .Z(n15647) );
  NOR U1453 ( .A(n20719), .B(n20720), .Z(n21715) );
  NOR U1454 ( .A(n21590), .B(n21591), .Z(n24895) );
  XNOR U1455 ( .A(n18908), .B(n18907), .Z(n15333) );
  XNOR U1456 ( .A(n20739), .B(n22786), .Z(n18193) );
  XNOR U1457 ( .A(n20610), .B(n21709), .Z(n17509) );
  XOR U1458 ( .A(n19283), .B(n18204), .Z(n14914) );
  NOR U1459 ( .A(n20649), .B(n23202), .Z(n23200) );
  NOR U1460 ( .A(n20653), .B(n20652), .Z(n20650) );
  XNOR U1461 ( .A(n18290), .B(n17197), .Z(n18237) );
  XNOR U1462 ( .A(n17563), .B(n17564), .Z(n15458) );
  XOR U1463 ( .A(n20959), .B(n18379), .Z(n14787) );
  XNOR U1464 ( .A(n18754), .B(n18434), .Z(n15180) );
  XOR U1465 ( .A(n20276), .B(n18707), .Z(n16843) );
  XNOR U1466 ( .A(n18273), .B(n17520), .Z(n14487) );
  XNOR U1467 ( .A(n19635), .B(n16021), .Z(n14660) );
  XOR U1468 ( .A(n17523), .B(n17458), .Z(n16719) );
  XOR U1469 ( .A(n17416), .B(n15132), .Z(n14340) );
  ANDN U1470 ( .B(n14864), .A(n15785), .Z(n15783) );
  NOR U1471 ( .A(n15665), .B(n18303), .Z(n18641) );
  XNOR U1472 ( .A(n12809), .B(n12810), .Z(n10358) );
  NOR U1473 ( .A(n15231), .B(n15230), .Z(n15228) );
  NOR U1474 ( .A(n15876), .B(n15878), .Z(n24889) );
  XNOR U1475 ( .A(n18823), .B(n13821), .Z(n11974) );
  ANDN U1476 ( .B(n13204), .A(n13205), .Z(n13202) );
  NOR U1477 ( .A(n12513), .B(n12514), .Z(n13578) );
  ANDN U1478 ( .B(n16507), .A(n14842), .Z(n18808) );
  ANDN U1479 ( .B(n13826), .A(n13824), .Z(n18567) );
  NOR U1480 ( .A(n12490), .B(n12491), .Z(n13567) );
  ANDN U1481 ( .B(n16317), .A(n14499), .Z(n20081) );
  NOR U1482 ( .A(n16123), .B(n13574), .Z(n16122) );
  ANDN U1483 ( .B(n13807), .A(n15190), .Z(n19373) );
  ANDN U1484 ( .B(n12772), .A(n12773), .Z(n12770) );
  NOR U1485 ( .A(n18061), .B(n17093), .Z(n19179) );
  ANDN U1486 ( .B(n17156), .A(n17177), .Z(n19621) );
  ANDN U1487 ( .B(n13691), .A(n14338), .Z(n14336) );
  ANDN U1488 ( .B(n13653), .A(n16089), .Z(n17607) );
  ANDN U1489 ( .B(n14426), .A(n14427), .Z(n14424) );
  NOR U1490 ( .A(n15412), .B(n13677), .Z(n15419) );
  ANDN U1491 ( .B(n13645), .A(n13646), .Z(n13643) );
  XNOR U1492 ( .A(n18311), .B(n13343), .Z(n13877) );
  NOR U1493 ( .A(n15618), .B(n14814), .Z(n15616) );
  NOR U1494 ( .A(n13440), .B(n16616), .Z(n16615) );
  ANDN U1495 ( .B(n13106), .A(n13107), .Z(n13104) );
  ANDN U1496 ( .B(n14927), .A(n15130), .Z(n15127) );
  NOR U1497 ( .A(n13927), .B(n13926), .Z(n13924) );
  ANDN U1498 ( .B(n14330), .A(n14329), .Z(n17396) );
  NOR U1499 ( .A(n14479), .B(n15462), .Z(n16275) );
  ANDN U1500 ( .B(n12749), .A(n12747), .Z(n13453) );
  ANDN U1501 ( .B(n17700), .A(n17310), .Z(n19772) );
  ANDN U1502 ( .B(n14359), .A(n14795), .Z(n14793) );
  XOR U1503 ( .A(n12986), .B(n12985), .Z(n9769) );
  ANDN U1504 ( .B(n13213), .A(n13214), .Z(n15836) );
  XNOR U1505 ( .A(n12162), .B(n12742), .Z(n11280) );
  XOR U1506 ( .A(n17662), .B(n14642), .Z(n9388) );
  NOR U1507 ( .A(n13636), .B(n13637), .Z(n14432) );
  ANDN U1508 ( .B(n17090), .A(n17091), .Z(n17088) );
  ANDN U1509 ( .B(n13450), .A(n15245), .Z(n17138) );
  XNOR U1510 ( .A(n14721), .B(n14722), .Z(n10771) );
  NOR U1511 ( .A(n14516), .B(n14517), .Z(n15995) );
  XOR U1512 ( .A(n14683), .B(n13905), .Z(n10373) );
  NOR U1513 ( .A(n13791), .B(n15195), .Z(n17375) );
  NOR U1514 ( .A(n14265), .B(n14264), .Z(n14262) );
  XOR U1515 ( .A(n13396), .B(n13395), .Z(n11684) );
  XNOR U1516 ( .A(n18138), .B(n15276), .Z(n12250) );
  XNOR U1517 ( .A(n19610), .B(n14090), .Z(n14080) );
  ANDN U1518 ( .B(n18619), .A(n15755), .Z(n20231) );
  XNOR U1519 ( .A(n15418), .B(n13939), .Z(n12640) );
  NOR U1520 ( .A(n13378), .B(n13118), .Z(n14902) );
  NOR U1521 ( .A(n13741), .B(n13742), .Z(n15790) );
  ANDN U1522 ( .B(n16578), .A(n16579), .Z(n16577) );
  NOR U1523 ( .A(n17286), .B(n16300), .Z(n17285) );
  XOR U1524 ( .A(n12584), .B(n12583), .Z(n10382) );
  NOR U1525 ( .A(n15177), .B(n15176), .Z(n15175) );
  NOR U1526 ( .A(n16373), .B(n16374), .Z(n17885) );
  XOR U1527 ( .A(n11790), .B(n11789), .Z(n9694) );
  NOR U1528 ( .A(n12904), .B(n12903), .Z(n12901) );
  XNOR U1529 ( .A(n11686), .B(n11685), .Z(n11500) );
  XOR U1530 ( .A(n10359), .B(n10818), .Z(n8092) );
  XOR U1531 ( .A(n12482), .B(n9187), .Z(n6401) );
  XNOR U1532 ( .A(n9526), .B(n11378), .Z(n7732) );
  NOR U1533 ( .A(n11492), .B(n11493), .Z(n14006) );
  NOR U1534 ( .A(n9852), .B(n9314), .Z(n9850) );
  ANDN U1535 ( .B(n6759), .A(n6760), .Z(n7348) );
  ANDN U1536 ( .B(n6876), .A(n6877), .Z(n7684) );
  ANDN U1537 ( .B(n8215), .A(n7109), .Z(n8213) );
  ANDN U1538 ( .B(n8337), .A(n8338), .Z(n8335) );
  XNOR U1539 ( .A(n8520), .B(n8521), .Z(n5546) );
  NOR U1540 ( .A(n7859), .B(n7858), .Z(n7856) );
  NOR U1541 ( .A(n6448), .B(n6447), .Z(n6445) );
  NOR U1542 ( .A(n6603), .B(n6602), .Z(n6600) );
  NOR U1543 ( .A(n11618), .B(n11617), .Z(n14625) );
  XNOR U1544 ( .A(n6291), .B(n6468), .Z(n4249) );
  NOR U1545 ( .A(n9753), .B(n8565), .Z(n9831) );
  ANDN U1546 ( .B(n7975), .A(n10740), .Z(n10866) );
  XNOR U1547 ( .A(n11672), .B(n7822), .Z(n1697) );
  ANDN U1548 ( .B(n10746), .A(n10745), .Z(n12157) );
  ANDN U1549 ( .B(n6595), .A(n6593), .Z(n7010) );
  XNOR U1550 ( .A(n12594), .B(n8865), .Z(n1927) );
  XNOR U1551 ( .A(n5987), .B(n5986), .Z(n1969) );
  XNOR U1552 ( .A(n5992), .B(n5991), .Z(n1972) );
  NOR U1553 ( .A(n10858), .B(n9032), .Z(n10856) );
  NOR U1554 ( .A(n6483), .B(n8882), .Z(n8881) );
  ANDN U1555 ( .B(n7963), .A(n7964), .Z(n7961) );
  NOR U1556 ( .A(n6902), .B(n6901), .Z(n6899) );
  ANDN U1557 ( .B(n7245), .A(n7155), .Z(n7244) );
  ANDN U1558 ( .B(n6997), .A(n6998), .Z(n6995) );
  ANDN U1559 ( .B(n7447), .A(n7526), .Z(n7525) );
  NOR U1560 ( .A(n8039), .B(n8038), .Z(n8037) );
  NOR U1561 ( .A(n7721), .B(n7720), .Z(n7718) );
  ANDN U1562 ( .B(n7870), .A(n7871), .Z(n7868) );
  NOR U1563 ( .A(n10738), .B(n7984), .Z(n10736) );
  ANDN U1564 ( .B(n6644), .A(n6643), .Z(n19538) );
  XNOR U1565 ( .A(n6158), .B(n8063), .Z(n1953) );
  XNOR U1566 ( .A(n6177), .B(n8233), .Z(n1660) );
  ANDN U1567 ( .B(n6831), .A(n6837), .Z(n7585) );
  NOR U1568 ( .A(n7404), .B(n7403), .Z(n7401) );
  ANDN U1569 ( .B(n7477), .A(n7478), .Z(n7475) );
  ANDN U1570 ( .B(n7559), .A(n7557), .Z(n8694) );
  ANDN U1571 ( .B(n7633), .A(n7634), .Z(n8728) );
  ANDN U1572 ( .B(n7844), .A(n7845), .Z(n8919) );
  ANDN U1573 ( .B(n7216), .A(n7214), .Z(n8296) );
  XNOR U1574 ( .A(n5997), .B(n5996), .Z(n4494) );
  NOR U1575 ( .A(n9979), .B(n7534), .Z(n9977) );
  ANDN U1576 ( .B(n9962), .A(n9961), .Z(n10419) );
  XOR U1577 ( .A(n6143), .B(n7836), .Z(n1939) );
  XOR U1578 ( .A(n6148), .B(n7945), .Z(n1943) );
  NOR U1579 ( .A(n9873), .B(n7434), .Z(n9959) );
  XOR U1580 ( .A(n6153), .B(n7996), .Z(n1947) );
  XNOR U1581 ( .A(n8842), .B(n8841), .Z(n3211) );
  XOR U1582 ( .A(n6239), .B(n9221), .Z(n1729) );
  XOR U1583 ( .A(n6243), .B(n9343), .Z(n1733) );
  XNOR U1584 ( .A(n6251), .B(n9541), .Z(n1742) );
  XNOR U1585 ( .A(n9498), .B(n6667), .Z(n5139) );
  ANDN U1586 ( .B(n7036), .A(n7037), .Z(n7035) );
  XOR U1587 ( .A(n2568), .B(n2569), .Z(n1902) );
  ANDN U1588 ( .B(n4390), .A(n4391), .Z(n4388) );
  ANDN U1589 ( .B(n4462), .A(n4463), .Z(n4460) );
  ANDN U1590 ( .B(n4474), .A(n4475), .Z(n4472) );
  NOR U1591 ( .A(n4512), .B(n4511), .Z(n4507) );
  ANDN U1592 ( .B(n4551), .A(n4552), .Z(n4549) );
  ANDN U1593 ( .B(n4555), .A(n4556), .Z(n4553) );
  ANDN U1594 ( .B(n4567), .A(n4568), .Z(n4565) );
  ANDN U1595 ( .B(n4585), .A(n4586), .Z(n4583) );
  ANDN U1596 ( .B(n4602), .A(n4603), .Z(n4600) );
  ANDN U1597 ( .B(n4630), .A(n4631), .Z(n4628) );
  ANDN U1598 ( .B(n4682), .A(n4399), .Z(n4681) );
  NOR U1599 ( .A(n4686), .B(n4410), .Z(n4685) );
  ANDN U1600 ( .B(n4690), .A(n4419), .Z(n4689) );
  ANDN U1601 ( .B(n4471), .A(n4721), .Z(n4720) );
  ANDN U1602 ( .B(n5028), .A(n4804), .Z(n5026) );
  NOR U1603 ( .A(n4950), .B(n4514), .Z(n5153) );
  ANDN U1604 ( .B(n4617), .A(n5031), .Z(n5219) );
  ANDN U1605 ( .B(n5666), .A(n1047), .Z(n5665) );
  ANDN U1606 ( .B(n5714), .A(n1132), .Z(n5713) );
  ANDN U1607 ( .B(n6109), .A(n5793), .Z(n6105) );
  NOR U1608 ( .A(n5848), .B(n1050), .Z(n6187) );
  NOR U1609 ( .A(n1208), .B(n1207), .Z(n1205) );
  ANDN U1610 ( .B(n1300), .A(n1301), .Z(n1298) );
  ANDN U1611 ( .B(n1352), .A(n1353), .Z(n1350) );
  ANDN U1612 ( .B(n1372), .A(n1373), .Z(n1370) );
  ANDN U1613 ( .B(n1376), .A(n1377), .Z(n1374) );
  XNOR U1614 ( .A(n1446), .B(n2156), .Z(out[907]) );
  ANDN U1615 ( .B(n1467), .A(n1468), .Z(n1465) );
  NOR U1616 ( .A(n1536), .B(n1275), .Z(n1535) );
  NOR U1617 ( .A(n1295), .B(n1749), .Z(n1549) );
  ANDN U1618 ( .B(n1603), .A(n1401), .Z(n1602) );
  NOR U1619 ( .A(n1826), .B(n1583), .Z(n1823) );
  ANDN U1620 ( .B(n1890), .A(n1620), .Z(n1887) );
  ANDN U1621 ( .B(n1966), .A(n1657), .Z(n1963) );
  NOR U1622 ( .A(n1250), .B(n1699), .Z(n1995) );
  XNOR U1623 ( .A(n2047), .B(n1777), .Z(out[744]) );
  NOR U1624 ( .A(n1945), .B(n1474), .Z(n2180) );
  NOR U1625 ( .A(n2840), .B(n2839), .Z(n2837) );
  ANDN U1626 ( .B(n3084), .A(n2889), .Z(n3083) );
  NOR U1627 ( .A(n3219), .B(n3020), .Z(n3217) );
  ANDN U1628 ( .B(n3238), .A(n3038), .Z(n3236) );
  NOR U1629 ( .A(n3292), .B(n3072), .Z(n3290) );
  NOR U1630 ( .A(n3152), .B(n2702), .Z(n3385) );
  NOR U1631 ( .A(n3174), .B(n2726), .Z(n3404) );
  ANDN U1632 ( .B(n2738), .A(n3183), .Z(n3411) );
  NOR U1633 ( .A(n2774), .B(n3212), .Z(n3434) );
  NOR U1634 ( .A(n2778), .B(n3216), .Z(n3436) );
  NOR U1635 ( .A(n2830), .B(n3259), .Z(n3472) );
  NOR U1636 ( .A(n3328), .B(n2912), .Z(n3527) );
  ANDN U1637 ( .B(n2932), .A(n3348), .Z(n3542) );
  NOR U1638 ( .A(n3894), .B(n2969), .Z(n3893) );
  NOR U1639 ( .A(n3478), .B(n3934), .Z(n3933) );
  ANDN U1640 ( .B(n4001), .A(n4002), .Z(n4000) );
  ANDN U1641 ( .B(n4019), .A(n4020), .Z(n4018) );
  ANDN U1642 ( .B(n4046), .A(n2846), .Z(n4044) );
  ANDN U1643 ( .B(n1516), .A(n3982), .Z(n4200) );
  NOR U1644 ( .A(n4043), .B(n2174), .Z(n4243) );
  NOR U1645 ( .A(n4100), .B(n3022), .Z(n4281) );
  NOR U1646 ( .A(n4117), .B(n3169), .Z(n4296) );
  ANDN U1647 ( .B(n2375), .A(n2376), .Z(n2373) );
  XNOR U1648 ( .A(n25141), .B(n25140), .Z(n24757) );
  XNOR U1649 ( .A(n26047), .B(n26046), .Z(n23121) );
  XOR U1650 ( .A(n25327), .B(n25113), .Z(n22831) );
  XNOR U1651 ( .A(n25468), .B(n25467), .Z(n22839) );
  XOR U1652 ( .A(n25486), .B(n25297), .Z(n21198) );
  XOR U1653 ( .A(n24549), .B(n25662), .Z(n24448) );
  XNOR U1654 ( .A(n25073), .B(n25393), .Z(n23241) );
  XNOR U1655 ( .A(n24881), .B(n25998), .Z(n22211) );
  XNOR U1656 ( .A(n25681), .B(n25680), .Z(n25133) );
  XOR U1657 ( .A(n25462), .B(n25461), .Z(n22635) );
  XNOR U1658 ( .A(n26094), .B(n25609), .Z(n24715) );
  XNOR U1659 ( .A(n25499), .B(n25230), .Z(n24171) );
  XNOR U1660 ( .A(n25660), .B(n24776), .Z(n22821) );
  XNOR U1661 ( .A(n25014), .B(n25013), .Z(n23599) );
  XNOR U1662 ( .A(n25144), .B(n25718), .Z(n24221) );
  XNOR U1663 ( .A(n24933), .B(n25653), .Z(n22371) );
  XNOR U1664 ( .A(n25336), .B(n25335), .Z(n21609) );
  XNOR U1665 ( .A(n24977), .B(n25126), .Z(n24183) );
  XOR U1666 ( .A(n25209), .B(n25768), .Z(n22432) );
  XNOR U1667 ( .A(n26007), .B(n25566), .Z(n23323) );
  XNOR U1668 ( .A(n25909), .B(n25092), .Z(n23777) );
  XNOR U1669 ( .A(n24510), .B(n24554), .Z(n22687) );
  XOR U1670 ( .A(n26066), .B(n24688), .Z(n23445) );
  XNOR U1671 ( .A(n24337), .B(n24336), .Z(n24219) );
  XNOR U1672 ( .A(n23829), .B(n24896), .Z(n22962) );
  XOR U1673 ( .A(n25899), .B(n26048), .Z(n24309) );
  XOR U1674 ( .A(n25535), .B(n24991), .Z(n25023) );
  XNOR U1675 ( .A(n25854), .B(n25466), .Z(n23295) );
  XNOR U1676 ( .A(n24665), .B(n25064), .Z(n23726) );
  XNOR U1677 ( .A(n25580), .B(n25932), .Z(n23904) );
  XOR U1678 ( .A(n24740), .B(n24739), .Z(n23130) );
  XOR U1679 ( .A(n25186), .B(n25185), .Z(n22822) );
  XOR U1680 ( .A(n25489), .B(n25091), .Z(n22278) );
  XOR U1681 ( .A(n24672), .B(n24671), .Z(n22221) );
  XNOR U1682 ( .A(n26175), .B(n25663), .Z(n21754) );
  XNOR U1683 ( .A(n25676), .B(n25460), .Z(n23595) );
  XNOR U1684 ( .A(n25274), .B(n25071), .Z(n24694) );
  XOR U1685 ( .A(n24566), .B(n24565), .Z(n21193) );
  XNOR U1686 ( .A(n24939), .B(n24938), .Z(n24872) );
  XOR U1687 ( .A(round_reg[1352]), .B(n24284), .Z(n21892) );
  XNOR U1688 ( .A(round_reg[1315]), .B(n23584), .Z(n22012) );
  XNOR U1689 ( .A(round_reg[71]), .B(n21316), .Z(n20602) );
  XOR U1690 ( .A(round_reg[804]), .B(n23482), .Z(n22801) );
  XOR U1691 ( .A(round_reg[1417]), .B(n23283), .Z(n21944) );
  XOR U1692 ( .A(round_reg[145]), .B(n22790), .Z(n23506) );
  XOR U1693 ( .A(round_reg[1182]), .B(n22751), .Z(n19104) );
  XNOR U1694 ( .A(round_reg[117]), .B(n23993), .Z(n19808) );
  XOR U1695 ( .A(round_reg[1569]), .B(n23745), .Z(n21024) );
  XOR U1696 ( .A(round_reg[814]), .B(n23908), .Z(n21648) );
  XOR U1697 ( .A(round_reg[848]), .B(n24229), .Z(n23573) );
  NOR U1698 ( .A(n20729), .B(n20730), .Z(n21722) );
  NOR U1699 ( .A(n22913), .B(n22912), .Z(n22911) );
  ANDN U1700 ( .B(n22290), .A(n22894), .Z(n22893) );
  NOR U1701 ( .A(n20358), .B(n23868), .Z(n23867) );
  ANDN U1702 ( .B(n20047), .A(n20045), .Z(n22443) );
  NOR U1703 ( .A(n22553), .B(n23633), .Z(n23632) );
  ANDN U1704 ( .B(n22162), .A(n23700), .Z(n23698) );
  ANDN U1705 ( .B(n22581), .A(n22460), .Z(n24590) );
  NOR U1706 ( .A(n23235), .B(n22487), .Z(n23233) );
  NOR U1707 ( .A(n23718), .B(n24039), .Z(n24310) );
  XNOR U1708 ( .A(n18856), .B(n18855), .Z(n17514) );
  ANDN U1709 ( .B(n21241), .A(n21328), .Z(n23589) );
  NOR U1710 ( .A(n22797), .B(n21666), .Z(n23281) );
  ANDN U1711 ( .B(n21585), .A(n21370), .Z(n24604) );
  XNOR U1712 ( .A(n20191), .B(n20190), .Z(n16471) );
  ANDN U1713 ( .B(n20419), .A(n22333), .Z(n22332) );
  ANDN U1714 ( .B(n22917), .A(n22918), .Z(n23498) );
  XNOR U1715 ( .A(n22453), .B(n22452), .Z(n19597) );
  NOR U1716 ( .A(n24603), .B(n24894), .Z(n24893) );
  NOR U1717 ( .A(n20264), .B(n20263), .Z(n20261) );
  ANDN U1718 ( .B(n20488), .A(n20489), .Z(n20486) );
  ANDN U1719 ( .B(n22190), .A(n22191), .Z(n22188) );
  XNOR U1720 ( .A(n19957), .B(n20194), .Z(n17154) );
  NOR U1721 ( .A(n19881), .B(n19883), .Z(n20575) );
  NOR U1722 ( .A(n20889), .B(n20887), .Z(n24765) );
  NOR U1723 ( .A(n19854), .B(n22226), .Z(n22224) );
  ANDN U1724 ( .B(n20656), .A(n20658), .Z(n24888) );
  XNOR U1725 ( .A(n18979), .B(n18978), .Z(n17360) );
  XNOR U1726 ( .A(n20688), .B(n20687), .Z(n17522) );
  XNOR U1727 ( .A(n21293), .B(n21052), .Z(n19982) );
  ANDN U1728 ( .B(n24263), .A(n21546), .Z(n24275) );
  XNOR U1729 ( .A(n21130), .B(n21129), .Z(n18832) );
  XNOR U1730 ( .A(n20604), .B(n20229), .Z(n18140) );
  XNOR U1731 ( .A(n24108), .B(n23191), .Z(n17928) );
  NOR U1732 ( .A(n22666), .B(n22667), .Z(n24916) );
  XNOR U1733 ( .A(n20703), .B(n19798), .Z(n17121) );
  XOR U1734 ( .A(n20940), .B(n23458), .Z(n16039) );
  NOR U1735 ( .A(n21631), .B(n20483), .Z(n22110) );
  XNOR U1736 ( .A(n20466), .B(n19632), .Z(n19423) );
  ANDN U1737 ( .B(n20009), .A(n20010), .Z(n20007) );
  XOR U1738 ( .A(n19322), .B(n19864), .Z(n18464) );
  NOR U1739 ( .A(n23173), .B(n23977), .Z(n24439) );
  XNOR U1740 ( .A(n21322), .B(n21321), .Z(n18180) );
  NOR U1741 ( .A(n21093), .B(n19965), .Z(n25472) );
  ANDN U1742 ( .B(n21115), .A(n21116), .Z(n21113) );
  ANDN U1743 ( .B(n21867), .A(n22619), .Z(n24645) );
  XNOR U1744 ( .A(n19344), .B(n19343), .Z(n16047) );
  XNOR U1745 ( .A(n21784), .B(n20579), .Z(n18399) );
  NOR U1746 ( .A(n23187), .B(n23186), .Z(n23184) );
  XNOR U1747 ( .A(n23128), .B(n18391), .Z(n16539) );
  NOR U1748 ( .A(n21975), .B(n23658), .Z(n24120) );
  ANDN U1749 ( .B(n21179), .A(n23929), .Z(n25296) );
  XNOR U1750 ( .A(n20327), .B(n20326), .Z(n20025) );
  XNOR U1751 ( .A(n21632), .B(n19961), .Z(n18109) );
  XNOR U1752 ( .A(n20085), .B(n22629), .Z(n17388) );
  NOR U1753 ( .A(n24173), .B(n22545), .Z(n24436) );
  XNOR U1754 ( .A(n18330), .B(n18329), .Z(n14948) );
  XNOR U1755 ( .A(n19769), .B(n19016), .Z(n17489) );
  XNOR U1756 ( .A(n22077), .B(n19902), .Z(n15208) );
  NOR U1757 ( .A(n20920), .B(n20921), .Z(n21705) );
  XNOR U1758 ( .A(n20030), .B(n20168), .Z(n18406) );
  XNOR U1759 ( .A(n22504), .B(n19327), .Z(n17951) );
  ANDN U1760 ( .B(n20891), .A(n22848), .Z(n22846) );
  XNOR U1761 ( .A(n20077), .B(n20076), .Z(n15851) );
  ANDN U1762 ( .B(n22493), .A(n22494), .Z(n22491) );
  XNOR U1763 ( .A(n21435), .B(n21434), .Z(n17560) );
  XNOR U1764 ( .A(n19744), .B(n19688), .Z(n15217) );
  XNOR U1765 ( .A(n19182), .B(n20444), .Z(n16343) );
  XOR U1766 ( .A(n21478), .B(n21477), .Z(n15252) );
  NOR U1767 ( .A(n20338), .B(n22020), .Z(n23878) );
  XNOR U1768 ( .A(n22382), .B(n22585), .Z(n19971) );
  XNOR U1769 ( .A(n17860), .B(n19686), .Z(n15896) );
  XOR U1770 ( .A(n18625), .B(n18624), .Z(n15753) );
  XOR U1771 ( .A(n15607), .B(n16762), .Z(n15017) );
  XOR U1772 ( .A(n20109), .B(n16751), .Z(n13119) );
  XNOR U1773 ( .A(n17244), .B(n17069), .Z(n13209) );
  XNOR U1774 ( .A(n19336), .B(n19337), .Z(n15193) );
  XNOR U1775 ( .A(n19714), .B(n16944), .Z(n14019) );
  XOR U1776 ( .A(n17251), .B(n16053), .Z(n13728) );
  XOR U1777 ( .A(n18044), .B(n18043), .Z(n15667) );
  XOR U1778 ( .A(n18747), .B(n15623), .Z(n15169) );
  XNOR U1779 ( .A(n17772), .B(n15525), .Z(n14074) );
  XNOR U1780 ( .A(n17944), .B(n17945), .Z(n16569) );
  NOR U1781 ( .A(n15179), .B(n13770), .Z(n18753) );
  XNOR U1782 ( .A(n19076), .B(n14995), .Z(n9923) );
  NOR U1783 ( .A(n18059), .B(n17089), .Z(n19177) );
  NOR U1784 ( .A(n13350), .B(n13351), .Z(n13872) );
  ANDN U1785 ( .B(n14307), .A(n14308), .Z(n19189) );
  ANDN U1786 ( .B(n15998), .A(n16096), .Z(n17622) );
  ANDN U1787 ( .B(n16886), .A(n17073), .Z(n20929) );
  ANDN U1788 ( .B(n13034), .A(n13035), .Z(n13032) );
  NOR U1789 ( .A(n16173), .B(n16172), .Z(n22142) );
  ANDN U1790 ( .B(n14897), .A(n15123), .Z(n15637) );
  NOR U1791 ( .A(n14864), .B(n14865), .Z(n19031) );
  NOR U1792 ( .A(n15381), .B(n14036), .Z(n18943) );
  NOR U1793 ( .A(n14720), .B(n16486), .Z(n23271) );
  NOR U1794 ( .A(n16590), .B(n15061), .Z(n17910) );
  NOR U1795 ( .A(n17701), .B(n17700), .Z(n17699) );
  XNOR U1796 ( .A(n18652), .B(n15669), .Z(n11557) );
  ANDN U1797 ( .B(n13629), .A(n13627), .Z(n14027) );
  ANDN U1798 ( .B(n14973), .A(n16604), .Z(n23611) );
  ANDN U1799 ( .B(n14791), .A(n14792), .Z(n14789) );
  XNOR U1800 ( .A(n13386), .B(n13385), .Z(n12832) );
  ANDN U1801 ( .B(n16189), .A(n16217), .Z(n17833) );
  XNOR U1802 ( .A(n17046), .B(n12805), .Z(n16442) );
  ANDN U1803 ( .B(n14616), .A(n13163), .Z(n17493) );
  NOR U1804 ( .A(n17653), .B(n15680), .Z(n17651) );
  NOR U1805 ( .A(n14501), .B(n16108), .Z(n16107) );
  ANDN U1806 ( .B(n14763), .A(n14764), .Z(n16346) );
  XNOR U1807 ( .A(n12785), .B(n11902), .Z(n11663) );
  ANDN U1808 ( .B(n16579), .A(n16407), .Z(n17935) );
  NOR U1809 ( .A(n13983), .B(n13982), .Z(n13980) );
  ANDN U1810 ( .B(n13519), .A(n13520), .Z(n13517) );
  ANDN U1811 ( .B(n13293), .A(n14671), .Z(n14669) );
  XOR U1812 ( .A(n12548), .B(n12547), .Z(n9894) );
  ANDN U1813 ( .B(n14767), .A(n15563), .Z(n15561) );
  XOR U1814 ( .A(n11754), .B(n11943), .Z(n9083) );
  ANDN U1815 ( .B(n13581), .A(n16114), .Z(n16113) );
  XOR U1816 ( .A(n12667), .B(n12666), .Z(n10692) );
  ANDN U1817 ( .B(n13173), .A(n15521), .Z(n15518) );
  XNOR U1818 ( .A(n18154), .B(n18155), .Z(n9662) );
  NOR U1819 ( .A(n15068), .B(n15067), .Z(n16583) );
  ANDN U1820 ( .B(n17883), .A(n16369), .Z(n18733) );
  ANDN U1821 ( .B(n14983), .A(n16149), .Z(n16147) );
  ANDN U1822 ( .B(n14752), .A(n16308), .Z(n16805) );
  XNOR U1823 ( .A(n14081), .B(n12319), .Z(n11875) );
  ANDN U1824 ( .B(n13141), .A(n13142), .Z(n17963) );
  XOR U1825 ( .A(n17460), .B(n12843), .Z(n9687) );
  ANDN U1826 ( .B(n18231), .A(n19792), .Z(n19786) );
  ANDN U1827 ( .B(n14347), .A(n13503), .Z(n18170) );
  ANDN U1828 ( .B(n13952), .A(n13953), .Z(n13950) );
  NOR U1829 ( .A(n11960), .B(n11961), .Z(n16299) );
  ANDN U1830 ( .B(n13665), .A(n13666), .Z(n13663) );
  ANDN U1831 ( .B(n15935), .A(n15934), .Z(n15932) );
  XNOR U1832 ( .A(n19232), .B(n15300), .Z(n11991) );
  ANDN U1833 ( .B(n15509), .A(n16428), .Z(n18921) );
  XNOR U1834 ( .A(n12578), .B(n12577), .Z(n11149) );
  XOR U1835 ( .A(n14009), .B(n13246), .Z(n11257) );
  ANDN U1836 ( .B(n16276), .A(n14481), .Z(n18281) );
  ANDN U1837 ( .B(n13233), .A(n13765), .Z(n13764) );
  NOR U1838 ( .A(n13203), .B(n13204), .Z(n15833) );
  ANDN U1839 ( .B(n14247), .A(n14246), .Z(n18902) );
  ANDN U1840 ( .B(n15725), .A(n13054), .Z(n15723) );
  ANDN U1841 ( .B(n14272), .A(n15625), .Z(n20794) );
  NOR U1842 ( .A(n15941), .B(n15942), .Z(n17022) );
  ANDN U1843 ( .B(n14798), .A(n14797), .Z(n21788) );
  XNOR U1844 ( .A(n15030), .B(n16211), .Z(n11837) );
  XNOR U1845 ( .A(n11075), .B(n12418), .Z(n12260) );
  XNOR U1846 ( .A(n12766), .B(n12765), .Z(n10557) );
  NOR U1847 ( .A(n15820), .B(n15819), .Z(n15818) );
  NOR U1848 ( .A(n13564), .B(n12486), .Z(n17448) );
  XNOR U1849 ( .A(n12687), .B(n11756), .Z(n9177) );
  ANDN U1850 ( .B(n15741), .A(n15742), .Z(n15740) );
  NOR U1851 ( .A(n14594), .B(n14022), .Z(n14593) );
  NOR U1852 ( .A(n18030), .B(n18671), .Z(n18669) );
  ANDN U1853 ( .B(n15150), .A(n14585), .Z(n16545) );
  NOR U1854 ( .A(n16856), .B(n17870), .Z(n17867) );
  XNOR U1855 ( .A(n15000), .B(n12714), .Z(n11309) );
  ANDN U1856 ( .B(n16537), .A(n15428), .Z(n24605) );
  XNOR U1857 ( .A(n10154), .B(n10153), .Z(n7807) );
  XOR U1858 ( .A(n11821), .B(n10679), .Z(n9834) );
  XOR U1859 ( .A(n16814), .B(n9505), .Z(n8548) );
  XNOR U1860 ( .A(n12205), .B(n13907), .Z(n8882) );
  ANDN U1861 ( .B(n7682), .A(n7756), .Z(n7755) );
  ANDN U1862 ( .B(n7822), .A(n10503), .Z(n10627) );
  XNOR U1863 ( .A(n10240), .B(n8585), .Z(n5064) );
  ANDN U1864 ( .B(n9746), .A(n9745), .Z(n11823) );
  NOR U1865 ( .A(n7258), .B(n7257), .Z(n7255) );
  ANDN U1866 ( .B(n7330), .A(n7331), .Z(n7328) );
  ANDN U1867 ( .B(n8263), .A(n8264), .Z(n11189) );
  NOR U1868 ( .A(n7670), .B(n7668), .Z(n11236) );
  ANDN U1869 ( .B(n10668), .A(n9733), .Z(n11861) );
  ANDN U1870 ( .B(n6788), .A(n6789), .Z(n7444) );
  NOR U1871 ( .A(n6781), .B(n6780), .Z(n6778) );
  NOR U1872 ( .A(n7060), .B(n8227), .Z(n11056) );
  XNOR U1873 ( .A(n6287), .B(n6438), .Z(n5142) );
  XNOR U1874 ( .A(n9933), .B(n9934), .Z(n7573) );
  ANDN U1875 ( .B(n8095), .A(n6991), .Z(n10829) );
  XNOR U1876 ( .A(n12214), .B(n8742), .Z(n8720) );
  ANDN U1877 ( .B(n7262), .A(n7261), .Z(n8369) );
  NOR U1878 ( .A(n8618), .B(n6392), .Z(n8616) );
  ANDN U1879 ( .B(n6401), .A(n6402), .Z(n12480) );
  NOR U1880 ( .A(n6681), .B(n6682), .Z(n7157) );
  ANDN U1881 ( .B(n6704), .A(n6703), .Z(n7227) );
  ANDN U1882 ( .B(n8176), .A(n8230), .Z(n8229) );
  ANDN U1883 ( .B(n8523), .A(n8647), .Z(n8646) );
  ANDN U1884 ( .B(n8936), .A(n8860), .Z(n8935) );
  NOR U1885 ( .A(n9048), .B(n8987), .Z(n9047) );
  ANDN U1886 ( .B(n6389), .A(n6390), .Z(n6387) );
  ANDN U1887 ( .B(n7828), .A(n7829), .Z(n7826) );
  ANDN U1888 ( .B(n6538), .A(n6539), .Z(n6536) );
  ANDN U1889 ( .B(n6653), .A(n6654), .Z(n6651) );
  ANDN U1890 ( .B(n6734), .A(n6735), .Z(n6732) );
  NOR U1891 ( .A(n7469), .B(n7351), .Z(n7468) );
  NOR U1892 ( .A(n8099), .B(n8162), .Z(n8161) );
  NOR U1893 ( .A(n9839), .B(n7389), .Z(n9837) );
  NOR U1894 ( .A(n10958), .B(n8116), .Z(n10956) );
  XNOR U1895 ( .A(n11480), .B(n11481), .Z(n3626) );
  NOR U1896 ( .A(n6687), .B(n6686), .Z(n6684) );
  ANDN U1897 ( .B(n6829), .A(n6830), .Z(n6827) );
  ANDN U1898 ( .B(n6890), .A(n6891), .Z(n6888) );
  ANDN U1899 ( .B(n9972), .A(n9973), .Z(n11124) );
  ANDN U1900 ( .B(n7198), .A(n7199), .Z(n7196) );
  ANDN U1901 ( .B(n7707), .A(n7708), .Z(n7705) );
  ANDN U1902 ( .B(n8001), .A(n8002), .Z(n7999) );
  ANDN U1903 ( .B(n7712), .A(n7710), .Z(n8791) );
  XNOR U1904 ( .A(n11633), .B(n11634), .Z(n3872) );
  XNOR U1905 ( .A(n9253), .B(n9254), .Z(n4905) );
  NOR U1906 ( .A(n11351), .B(n8274), .Z(n11349) );
  XNOR U1907 ( .A(n5982), .B(n5981), .Z(n4357) );
  NOR U1908 ( .A(n7344), .B(n7342), .Z(n8446) );
  ANDN U1909 ( .B(n7493), .A(n7494), .Z(n8627) );
  NOR U1910 ( .A(n7784), .B(n7783), .Z(n7781) );
  ANDN U1911 ( .B(n7859), .A(n7857), .Z(n8916) );
  ANDN U1912 ( .B(n8018), .A(n8017), .Z(n9059) );
  ANDN U1913 ( .B(n9471), .A(n9472), .Z(n9469) );
  NOR U1914 ( .A(n7978), .B(n10746), .Z(n10744) );
  ANDN U1915 ( .B(n6460), .A(n6461), .Z(n6458) );
  NOR U1916 ( .A(n6562), .B(n6561), .Z(n6559) );
  NOR U1917 ( .A(n6595), .B(n6594), .Z(n6592) );
  NOR U1918 ( .A(n6813), .B(n6812), .Z(n6810) );
  NOR U1919 ( .A(n7413), .B(n7412), .Z(n7410) );
  NOR U1920 ( .A(n7960), .B(n7959), .Z(n7957) );
  ANDN U1921 ( .B(n8781), .A(n8780), .Z(n11371) );
  NOR U1922 ( .A(n8032), .B(n8031), .Z(n8029) );
  NOR U1923 ( .A(n9135), .B(n9053), .Z(n9134) );
  ANDN U1924 ( .B(n7542), .A(n9969), .Z(n10411) );
  XOR U1925 ( .A(n6186), .B(n8560), .Z(n1672) );
  XNOR U1926 ( .A(n6190), .B(n9311), .Z(n1677) );
  ANDN U1927 ( .B(n8057), .A(n10844), .Z(n10982) );
  ANDN U1928 ( .B(n11358), .A(n10519), .Z(n11545) );
  ANDN U1929 ( .B(n11498), .A(n10632), .Z(n11679) );
  ANDN U1930 ( .B(n11934), .A(n10865), .Z(n12163) );
  NOR U1931 ( .A(n10978), .B(n12122), .Z(n12328) );
  NOR U1932 ( .A(n11086), .B(n12272), .Z(n12469) );
  XOR U1933 ( .A(n6235), .B(n9121), .Z(n1725) );
  ANDN U1934 ( .B(n12101), .A(n14464), .Z(n16754) );
  XNOR U1935 ( .A(n5411), .B(n2291), .Z(n4515) );
  XOR U1936 ( .A(n3709), .B(n2555), .Z(n2808) );
  XNOR U1937 ( .A(n4582), .B(n4577), .Z(out[1551]) );
  NOR U1938 ( .A(n4688), .B(n4414), .Z(n4687) );
  NOR U1939 ( .A(n4696), .B(n4430), .Z(n4695) );
  NOR U1940 ( .A(n4953), .B(n4747), .Z(n4951) );
  ANDN U1941 ( .B(n4956), .A(n4750), .Z(n4954) );
  ANDN U1942 ( .B(n5009), .A(n4794), .Z(n5006) );
  NOR U1943 ( .A(n4827), .B(n4360), .Z(n5061) );
  NOR U1944 ( .A(n4936), .B(n4498), .Z(n5146) );
  ANDN U1945 ( .B(n4530), .A(n4962), .Z(n5164) );
  NOR U1946 ( .A(n5005), .B(n4584), .Z(n5201) );
  NOR U1947 ( .A(n5037), .B(n4625), .Z(n5230) );
  ANDN U1948 ( .B(n5620), .A(n5621), .Z(n5618) );
  ANDN U1949 ( .B(n5657), .A(n5658), .Z(n5655) );
  ANDN U1950 ( .B(n5740), .A(n1175), .Z(n5739) );
  ANDN U1951 ( .B(n5650), .A(n5822), .Z(n5821) );
  NOR U1952 ( .A(n6018), .B(n5747), .Z(n6014) );
  NOR U1953 ( .A(n6074), .B(n5775), .Z(n6070) );
  NOR U1954 ( .A(n5833), .B(n1042), .Z(n6179) );
  NOR U1955 ( .A(n5903), .B(n1094), .Z(n6232) );
  NOR U1956 ( .A(n5918), .B(n1106), .Z(n6244) );
  NOR U1957 ( .A(n1292), .B(n1291), .Z(n1289) );
  ANDN U1958 ( .B(n1340), .A(n1341), .Z(n1338) );
  ANDN U1959 ( .B(n1412), .A(n1413), .Z(n1410) );
  NOR U1960 ( .A(n1300), .B(n1754), .Z(n1551) );
  NOR U1961 ( .A(n1320), .B(n1777), .Z(n1559) );
  ANDN U1962 ( .B(n1563), .A(n1329), .Z(n1562) );
  ANDN U1963 ( .B(n1599), .A(n1388), .Z(n1598) );
  ANDN U1964 ( .B(n1538), .A(n1730), .Z(n1727) );
  NOR U1965 ( .A(n1941), .B(n1646), .Z(n1938) );
  NOR U1966 ( .A(n1678), .B(n1230), .Z(n1976) );
  ANDN U1967 ( .B(n1323), .A(n1781), .Z(n2050) );
  NOR U1968 ( .A(n1439), .B(n1902), .Z(n2147) );
  NOR U1969 ( .A(n1914), .B(n2156), .Z(n2153) );
  NOR U1970 ( .A(n2780), .B(n2779), .Z(n2777) );
  ANDN U1971 ( .B(n2964), .A(n2691), .Z(n2963) );
  ANDN U1972 ( .B(n3016), .A(n2775), .Z(n3015) );
  ANDN U1973 ( .B(n3038), .A(n2811), .Z(n3037) );
  NOR U1974 ( .A(n3065), .B(n2861), .Z(n3064) );
  ANDN U1975 ( .B(n3223), .A(n3026), .Z(n3220) );
  NOR U1976 ( .A(n3249), .B(n3042), .Z(n3247) );
  ANDN U1977 ( .B(n3252), .A(n3044), .Z(n3250) );
  NOR U1978 ( .A(n3245), .B(n2814), .Z(n3462) );
  ANDN U1979 ( .B(n3270), .A(n2842), .Z(n3482) );
  ANDN U1980 ( .B(n3292), .A(n2872), .Z(n3499) );
  NOR U1981 ( .A(n3303), .B(n2884), .Z(n3513) );
  NOR U1982 ( .A(n2900), .B(n3313), .Z(n3521) );
  NOR U1983 ( .A(n2904), .B(n3321), .Z(n3523) );
  NOR U1984 ( .A(n3333), .B(n2916), .Z(n3529) );
  ANDN U1985 ( .B(n3904), .A(n3076), .Z(n3903) );
  ANDN U1986 ( .B(n3909), .A(n3129), .Z(n3908) );
  ANDN U1987 ( .B(n3280), .A(n3917), .Z(n3916) );
  NOR U1988 ( .A(n3919), .B(n3317), .Z(n3918) );
  ANDN U1989 ( .B(n3925), .A(n3966), .Z(n3964) );
  ANDN U1990 ( .B(n4037), .A(n1479), .Z(n4034) );
  XNOR U1991 ( .A(n4063), .B(n2597), .Z(out[256]) );
  ANDN U1992 ( .B(n4084), .A(n3890), .Z(n4082) );
  ANDN U1993 ( .B(n4090), .A(n3892), .Z(n4088) );
  NOR U1994 ( .A(n3957), .B(n1170), .Z(n4173) );
  NOR U1995 ( .A(n1908), .B(n4019), .Z(n4224) );
  NOR U1996 ( .A(n4049), .B(n4250), .Z(n4247) );
  ANDN U1997 ( .B(n2670), .A(n4068), .Z(n4258) );
  ANDN U1998 ( .B(n2758), .A(n4074), .Z(n4265) );
  NOR U1999 ( .A(n1518), .B(n1517), .Z(n1515) );
  NOR U2000 ( .A(n1567), .B(n1566), .Z(n1564) );
  NOR U2001 ( .A(n1640), .B(n1639), .Z(n1637) );
  NOR U2002 ( .A(n1669), .B(n1668), .Z(n1666) );
  ANDN U2003 ( .B(n1716), .A(n1717), .Z(n1714) );
  ANDN U2004 ( .B(n2027), .A(n2028), .Z(n2025) );
  ANDN U2005 ( .B(n2175), .A(n2176), .Z(n2173) );
  ANDN U2006 ( .B(n2227), .A(n2228), .Z(n2225) );
  ANDN U2007 ( .B(n2449), .A(n2450), .Z(n2447) );
  ANDN U2008 ( .B(n2969), .A(n2970), .Z(n2967) );
  ANDN U2009 ( .B(n3023), .A(n3024), .Z(n3021) );
  ANDN U2010 ( .B(n3049), .A(n3050), .Z(n3047) );
  ANDN U2011 ( .B(n3170), .A(n3171), .Z(n3168) );
  ANDN U2012 ( .B(n3359), .A(n3360), .Z(n3357) );
  ANDN U2013 ( .B(n3478), .A(n3479), .Z(n3476) );
  ANDN U2014 ( .B(n3573), .A(n3574), .Z(n3571) );
  ANDN U2015 ( .B(n3723), .A(n1084), .Z(n3722) );
  ANDN U2016 ( .B(n3775), .A(n1127), .Z(n3774) );
  ANDN U2017 ( .B(n3878), .A(n1215), .Z(n3877) );
  ANDN U2018 ( .B(n1035), .A(n1036), .Z(n1033) );
  NOR U2019 ( .A(n3508), .B(n2375), .Z(n3507) );
  XOR U2020 ( .A(n1033), .B(n1034), .Z(out[9]) );
  XNOR U2021 ( .A(n1037), .B(n1038), .Z(out[99]) );
  ANDN U2022 ( .B(n1039), .A(n1040), .Z(n1037) );
  XNOR U2023 ( .A(n1041), .B(n1042), .Z(out[999]) );
  AND U2024 ( .A(n1043), .B(n1044), .Z(n1041) );
  XNOR U2025 ( .A(n1045), .B(n1046), .Z(out[998]) );
  ANDN U2026 ( .B(n1047), .A(n1048), .Z(n1045) );
  XNOR U2027 ( .A(n1049), .B(n1050), .Z(out[997]) );
  ANDN U2028 ( .B(n1051), .A(n1052), .Z(n1049) );
  XNOR U2029 ( .A(n1053), .B(n1054), .Z(out[996]) );
  XNOR U2030 ( .A(n1057), .B(n1058), .Z(out[995]) );
  ANDN U2031 ( .B(n1059), .A(n1060), .Z(n1057) );
  XNOR U2032 ( .A(n1061), .B(n1062), .Z(out[994]) );
  AND U2033 ( .A(n1063), .B(n1064), .Z(n1061) );
  XNOR U2034 ( .A(n1065), .B(n1066), .Z(out[993]) );
  AND U2035 ( .A(n1067), .B(n1068), .Z(n1065) );
  XOR U2036 ( .A(n1069), .B(n1070), .Z(out[992]) );
  ANDN U2037 ( .B(n1071), .A(n1072), .Z(n1069) );
  XNOR U2038 ( .A(n1073), .B(n1074), .Z(out[991]) );
  AND U2039 ( .A(n1075), .B(n1076), .Z(n1073) );
  XNOR U2040 ( .A(n1077), .B(n1078), .Z(out[990]) );
  AND U2041 ( .A(n1079), .B(n1080), .Z(n1077) );
  XNOR U2042 ( .A(n1081), .B(n1082), .Z(out[98]) );
  AND U2043 ( .A(n1083), .B(n1084), .Z(n1081) );
  XNOR U2044 ( .A(n1085), .B(n1086), .Z(out[989]) );
  ANDN U2045 ( .B(n1087), .A(n1088), .Z(n1085) );
  XNOR U2046 ( .A(n1089), .B(n1090), .Z(out[988]) );
  ANDN U2047 ( .B(n1091), .A(n1092), .Z(n1089) );
  XNOR U2048 ( .A(n1093), .B(n1094), .Z(out[987]) );
  AND U2049 ( .A(n1095), .B(n1096), .Z(n1093) );
  XNOR U2050 ( .A(n1097), .B(n1098), .Z(out[986]) );
  NOR U2051 ( .A(n1099), .B(n1100), .Z(n1097) );
  XNOR U2052 ( .A(n1101), .B(n1102), .Z(out[985]) );
  ANDN U2053 ( .B(n1103), .A(n1104), .Z(n1101) );
  XNOR U2054 ( .A(n1105), .B(n1106), .Z(out[984]) );
  AND U2055 ( .A(n1107), .B(n1108), .Z(n1105) );
  XNOR U2056 ( .A(n1109), .B(n1110), .Z(out[983]) );
  AND U2057 ( .A(n1111), .B(n1112), .Z(n1109) );
  XNOR U2058 ( .A(n1113), .B(n1114), .Z(out[982]) );
  ANDN U2059 ( .B(n1115), .A(n1116), .Z(n1113) );
  XNOR U2060 ( .A(n1117), .B(n1118), .Z(out[981]) );
  NOR U2061 ( .A(n1119), .B(n1120), .Z(n1117) );
  XNOR U2062 ( .A(n1121), .B(n1122), .Z(out[980]) );
  AND U2063 ( .A(n1123), .B(n1124), .Z(n1121) );
  XOR U2064 ( .A(n1125), .B(n1126), .Z(out[97]) );
  ANDN U2065 ( .B(n1127), .A(n1128), .Z(n1125) );
  XNOR U2066 ( .A(n1129), .B(n1130), .Z(out[979]) );
  AND U2067 ( .A(n1131), .B(n1132), .Z(n1129) );
  XNOR U2068 ( .A(n1133), .B(n1134), .Z(out[978]) );
  NOR U2069 ( .A(n1135), .B(n1136), .Z(n1133) );
  XNOR U2070 ( .A(n1137), .B(n1138), .Z(out[977]) );
  ANDN U2071 ( .B(n1139), .A(n1140), .Z(n1137) );
  XNOR U2072 ( .A(n1141), .B(n1142), .Z(out[976]) );
  NOR U2073 ( .A(n1143), .B(n1144), .Z(n1141) );
  XNOR U2074 ( .A(n1145), .B(n1146), .Z(out[975]) );
  NOR U2075 ( .A(n1147), .B(n1148), .Z(n1145) );
  XNOR U2076 ( .A(n1149), .B(n1150), .Z(out[974]) );
  NOR U2077 ( .A(n1151), .B(n1152), .Z(n1149) );
  XNOR U2078 ( .A(n1153), .B(n1154), .Z(out[973]) );
  AND U2079 ( .A(n1155), .B(n1156), .Z(n1153) );
  XNOR U2080 ( .A(n1157), .B(n1158), .Z(out[972]) );
  AND U2081 ( .A(n1159), .B(n1160), .Z(n1157) );
  XNOR U2082 ( .A(n1161), .B(n1162), .Z(out[971]) );
  AND U2083 ( .A(n1163), .B(n1164), .Z(n1161) );
  XNOR U2084 ( .A(n1165), .B(n1166), .Z(out[970]) );
  AND U2085 ( .A(n1167), .B(n1168), .Z(n1165) );
  XNOR U2086 ( .A(n1169), .B(n1170), .Z(out[96]) );
  ANDN U2087 ( .B(n1171), .A(n1172), .Z(n1169) );
  XNOR U2088 ( .A(n1173), .B(n1174), .Z(out[969]) );
  ANDN U2089 ( .B(n1175), .A(n1176), .Z(n1173) );
  XNOR U2090 ( .A(n1177), .B(n1178), .Z(out[968]) );
  ANDN U2091 ( .B(n1179), .A(n1180), .Z(n1177) );
  XNOR U2092 ( .A(n1181), .B(n1182), .Z(out[967]) );
  AND U2093 ( .A(n1183), .B(n1184), .Z(n1181) );
  XNOR U2094 ( .A(n1185), .B(n1186), .Z(out[966]) );
  AND U2095 ( .A(n1187), .B(n1188), .Z(n1185) );
  XOR U2096 ( .A(n1189), .B(n1190), .Z(out[965]) );
  ANDN U2097 ( .B(n1191), .A(n1192), .Z(n1189) );
  XNOR U2098 ( .A(n1193), .B(n1194), .Z(out[964]) );
  AND U2099 ( .A(n1195), .B(n1196), .Z(n1193) );
  XNOR U2100 ( .A(n1197), .B(n1198), .Z(out[963]) );
  NOR U2101 ( .A(n1199), .B(n1200), .Z(n1197) );
  XOR U2102 ( .A(n1201), .B(n1202), .Z(out[962]) );
  ANDN U2103 ( .B(n1203), .A(n1204), .Z(n1201) );
  XNOR U2104 ( .A(n1205), .B(n1206), .Z(out[961]) );
  XNOR U2105 ( .A(n1209), .B(n1210), .Z(out[960]) );
  AND U2106 ( .A(n1211), .B(n1212), .Z(n1209) );
  XNOR U2107 ( .A(n1213), .B(n1214), .Z(out[95]) );
  ANDN U2108 ( .B(n1215), .A(n1216), .Z(n1213) );
  XNOR U2109 ( .A(n1217), .B(n1218), .Z(out[959]) );
  AND U2110 ( .A(n1219), .B(n1220), .Z(n1217) );
  XNOR U2111 ( .A(n1221), .B(n1222), .Z(out[958]) );
  AND U2112 ( .A(n1223), .B(n1224), .Z(n1221) );
  XNOR U2113 ( .A(n1225), .B(n1226), .Z(out[957]) );
  ANDN U2114 ( .B(n1227), .A(n1228), .Z(n1225) );
  XNOR U2115 ( .A(n1229), .B(n1230), .Z(out[956]) );
  ANDN U2116 ( .B(n1231), .A(n1232), .Z(n1229) );
  XNOR U2117 ( .A(n1233), .B(n1234), .Z(out[955]) );
  ANDN U2118 ( .B(n1235), .A(n1236), .Z(n1233) );
  XNOR U2119 ( .A(n1237), .B(n1238), .Z(out[954]) );
  AND U2120 ( .A(n1239), .B(n1240), .Z(n1237) );
  XNOR U2121 ( .A(n1241), .B(n1242), .Z(out[953]) );
  AND U2122 ( .A(n1243), .B(n1244), .Z(n1241) );
  XNOR U2123 ( .A(n1245), .B(n1246), .Z(out[952]) );
  AND U2124 ( .A(n1247), .B(n1248), .Z(n1245) );
  XNOR U2125 ( .A(n1249), .B(n1250), .Z(out[951]) );
  NOR U2126 ( .A(n1251), .B(n1252), .Z(n1249) );
  XNOR U2127 ( .A(n1253), .B(n1254), .Z(out[950]) );
  ANDN U2128 ( .B(n1255), .A(n1256), .Z(n1253) );
  XOR U2129 ( .A(n1257), .B(n1258), .Z(out[94]) );
  AND U2130 ( .A(n1259), .B(n1260), .Z(n1257) );
  XNOR U2131 ( .A(n1261), .B(n1262), .Z(out[949]) );
  ANDN U2132 ( .B(n1263), .A(n1264), .Z(n1261) );
  XNOR U2133 ( .A(n1265), .B(n1266), .Z(out[948]) );
  ANDN U2134 ( .B(n1267), .A(n1268), .Z(n1265) );
  XNOR U2135 ( .A(n1269), .B(n1270), .Z(out[947]) );
  XNOR U2136 ( .A(n1273), .B(n1274), .Z(out[946]) );
  AND U2137 ( .A(n1275), .B(n1276), .Z(n1273) );
  XNOR U2138 ( .A(n1277), .B(n1278), .Z(out[945]) );
  ANDN U2139 ( .B(n1279), .A(n1280), .Z(n1277) );
  XNOR U2140 ( .A(n1281), .B(n1282), .Z(out[944]) );
  XNOR U2141 ( .A(n1285), .B(n1286), .Z(out[943]) );
  ANDN U2142 ( .B(n1287), .A(n1288), .Z(n1285) );
  XOR U2143 ( .A(n1289), .B(n1290), .Z(out[942]) );
  AND U2144 ( .A(n1295), .B(n1296), .Z(n1293) );
  IV U2145 ( .A(n1297), .Z(n1296) );
  XNOR U2146 ( .A(n1298), .B(n1299), .Z(out[940]) );
  XNOR U2147 ( .A(n1302), .B(n1303), .Z(out[93]) );
  NOR U2148 ( .A(n1304), .B(n1305), .Z(n1302) );
  XOR U2149 ( .A(n1306), .B(n1307), .Z(out[939]) );
  ANDN U2150 ( .B(n1308), .A(n1309), .Z(n1306) );
  XOR U2151 ( .A(n1310), .B(n1311), .Z(out[938]) );
  ANDN U2152 ( .B(n1312), .A(n1313), .Z(n1310) );
  XOR U2153 ( .A(n1314), .B(n1315), .Z(out[937]) );
  NOR U2154 ( .A(n1316), .B(n1317), .Z(n1314) );
  XNOR U2155 ( .A(n1318), .B(n1319), .Z(out[936]) );
  XOR U2156 ( .A(n1322), .B(n1323), .Z(out[935]) );
  ANDN U2157 ( .B(n1324), .A(n1325), .Z(n1322) );
  XNOR U2158 ( .A(n1326), .B(n1327), .Z(out[934]) );
  AND U2159 ( .A(n1328), .B(n1329), .Z(n1326) );
  XNOR U2160 ( .A(n1330), .B(n1331), .Z(out[933]) );
  AND U2161 ( .A(n1332), .B(n1333), .Z(n1330) );
  XOR U2162 ( .A(n1334), .B(n1335), .Z(out[932]) );
  ANDN U2163 ( .B(n1336), .A(n1337), .Z(n1334) );
  XNOR U2164 ( .A(n1338), .B(n1339), .Z(out[931]) );
  XOR U2165 ( .A(n1342), .B(n1343), .Z(out[930]) );
  ANDN U2166 ( .B(n1344), .A(n1345), .Z(n1342) );
  XNOR U2167 ( .A(n1346), .B(n1347), .Z(out[92]) );
  AND U2168 ( .A(n1348), .B(n1349), .Z(n1346) );
  XNOR U2169 ( .A(n1350), .B(n1351), .Z(out[929]) );
  XNOR U2170 ( .A(n1354), .B(n1355), .Z(out[928]) );
  ANDN U2171 ( .B(n1356), .A(n1357), .Z(n1354) );
  XNOR U2172 ( .A(n1358), .B(n1359), .Z(out[927]) );
  XNOR U2173 ( .A(n1362), .B(n1363), .Z(out[926]) );
  XNOR U2174 ( .A(n1366), .B(n1367), .Z(out[925]) );
  ANDN U2175 ( .B(n1368), .A(n1369), .Z(n1366) );
  XNOR U2176 ( .A(n1370), .B(n1371), .Z(out[924]) );
  XNOR U2177 ( .A(n1374), .B(n1375), .Z(out[923]) );
  XNOR U2178 ( .A(n1378), .B(n1379), .Z(out[922]) );
  ANDN U2179 ( .B(n1380), .A(n1381), .Z(n1378) );
  XOR U2180 ( .A(n1382), .B(n1383), .Z(out[921]) );
  ANDN U2181 ( .B(n1384), .A(n1385), .Z(n1382) );
  XNOR U2182 ( .A(n1386), .B(n1387), .Z(out[920]) );
  ANDN U2183 ( .B(n1388), .A(n1389), .Z(n1386) );
  XNOR U2184 ( .A(n1390), .B(n1391), .Z(out[91]) );
  AND U2185 ( .A(n1392), .B(n1393), .Z(n1390) );
  XNOR U2186 ( .A(n1394), .B(n1395), .Z(out[919]) );
  AND U2187 ( .A(n1396), .B(n1397), .Z(n1394) );
  XOR U2188 ( .A(n1398), .B(n1399), .Z(out[918]) );
  AND U2189 ( .A(n1400), .B(n1401), .Z(n1398) );
  XNOR U2190 ( .A(n1402), .B(n1403), .Z(out[917]) );
  AND U2191 ( .A(n1404), .B(n1405), .Z(n1402) );
  XOR U2192 ( .A(n1406), .B(n1407), .Z(out[916]) );
  ANDN U2193 ( .B(n1408), .A(n1409), .Z(n1406) );
  XNOR U2194 ( .A(n1410), .B(n1411), .Z(out[915]) );
  XNOR U2195 ( .A(n1414), .B(n1415), .Z(out[914]) );
  ANDN U2196 ( .B(n1416), .A(n1417), .Z(n1414) );
  XOR U2197 ( .A(n1418), .B(n1419), .Z(out[913]) );
  ANDN U2198 ( .B(n1420), .A(n1421), .Z(n1418) );
  XNOR U2199 ( .A(n1422), .B(n1423), .Z(out[912]) );
  ANDN U2200 ( .B(n1424), .A(n1425), .Z(n1422) );
  XNOR U2201 ( .A(n1426), .B(n1427), .Z(out[911]) );
  ANDN U2202 ( .B(n1428), .A(n1429), .Z(n1426) );
  XNOR U2203 ( .A(n1430), .B(n1431), .Z(out[910]) );
  AND U2204 ( .A(n1432), .B(n1433), .Z(n1430) );
  XNOR U2205 ( .A(n1434), .B(n1435), .Z(out[90]) );
  ANDN U2206 ( .B(n1436), .A(n1437), .Z(n1434) );
  XNOR U2207 ( .A(n1438), .B(n1439), .Z(out[909]) );
  NOR U2208 ( .A(n1440), .B(n1441), .Z(n1438) );
  XNOR U2209 ( .A(n1442), .B(n1443), .Z(out[908]) );
  AND U2210 ( .A(n1444), .B(n1445), .Z(n1442) );
  NOR U2211 ( .A(n1447), .B(n1448), .Z(n1446) );
  XNOR U2212 ( .A(n1449), .B(n1450), .Z(out[906]) );
  AND U2213 ( .A(n1451), .B(n1452), .Z(n1449) );
  XNOR U2214 ( .A(n1453), .B(n1454), .Z(out[905]) );
  NOR U2215 ( .A(n1455), .B(n1456), .Z(n1453) );
  XNOR U2216 ( .A(n1457), .B(n1458), .Z(out[904]) );
  AND U2217 ( .A(n1459), .B(n1460), .Z(n1457) );
  XNOR U2218 ( .A(n1461), .B(n1462), .Z(out[903]) );
  XNOR U2219 ( .A(n1465), .B(n1466), .Z(out[902]) );
  XNOR U2220 ( .A(n1469), .B(n1470), .Z(out[901]) );
  AND U2221 ( .A(n1471), .B(n1472), .Z(n1469) );
  XNOR U2222 ( .A(n1473), .B(n1474), .Z(out[900]) );
  ANDN U2223 ( .B(n1475), .A(n1476), .Z(n1473) );
  XOR U2224 ( .A(n1477), .B(n1478), .Z(out[8]) );
  ANDN U2225 ( .B(n1479), .A(n1480), .Z(n1477) );
  XNOR U2226 ( .A(n1481), .B(n1482), .Z(out[89]) );
  AND U2227 ( .A(n1483), .B(n1484), .Z(n1481) );
  XNOR U2228 ( .A(n1485), .B(n1486), .Z(out[899]) );
  ANDN U2229 ( .B(n1487), .A(n1488), .Z(n1485) );
  XNOR U2230 ( .A(n1489), .B(n1490), .Z(out[898]) );
  AND U2231 ( .A(n1491), .B(n1492), .Z(n1489) );
  XNOR U2232 ( .A(n1493), .B(n1494), .Z(out[897]) );
  XNOR U2233 ( .A(n1497), .B(n1498), .Z(out[896]) );
  AND U2234 ( .A(n1499), .B(n1500), .Z(n1497) );
  XNOR U2235 ( .A(n1501), .B(n1219), .Z(out[895]) );
  AND U2236 ( .A(n1502), .B(n1503), .Z(n1501) );
  XNOR U2237 ( .A(n1504), .B(n1224), .Z(out[894]) );
  ANDN U2238 ( .B(n1505), .A(n1223), .Z(n1504) );
  XNOR U2239 ( .A(n1506), .B(n1227), .Z(out[893]) );
  AND U2240 ( .A(n1228), .B(n1507), .Z(n1506) );
  XNOR U2241 ( .A(n1508), .B(n1231), .Z(out[892]) );
  AND U2242 ( .A(n1232), .B(n1509), .Z(n1508) );
  XOR U2243 ( .A(n1510), .B(n1236), .Z(out[891]) );
  ANDN U2244 ( .B(n1511), .A(n1235), .Z(n1510) );
  XNOR U2245 ( .A(n1512), .B(n1239), .Z(out[890]) );
  AND U2246 ( .A(n1513), .B(n1514), .Z(n1512) );
  XOR U2247 ( .A(n1515), .B(n1516), .Z(out[88]) );
  XNOR U2248 ( .A(n1519), .B(n1243), .Z(out[889]) );
  AND U2249 ( .A(n1520), .B(n1521), .Z(n1519) );
  XNOR U2250 ( .A(n1522), .B(n1248), .Z(out[888]) );
  ANDN U2251 ( .B(n1523), .A(n1247), .Z(n1522) );
  XOR U2252 ( .A(n1524), .B(n1252), .Z(out[887]) );
  AND U2253 ( .A(n1251), .B(n1525), .Z(n1524) );
  XOR U2254 ( .A(n1526), .B(n1256), .Z(out[886]) );
  AND U2255 ( .A(n1527), .B(n1528), .Z(n1526) );
  XNOR U2256 ( .A(n1529), .B(n1263), .Z(out[885]) );
  AND U2257 ( .A(n1264), .B(n1530), .Z(n1529) );
  XNOR U2258 ( .A(n1531), .B(n1267), .Z(out[884]) );
  AND U2259 ( .A(n1268), .B(n1532), .Z(n1531) );
  XNOR U2260 ( .A(n1533), .B(n1271), .Z(out[883]) );
  AND U2261 ( .A(n1272), .B(n1534), .Z(n1533) );
  XNOR U2262 ( .A(n1535), .B(n1276), .Z(out[882]) );
  XNOR U2263 ( .A(n1537), .B(n1279), .Z(out[881]) );
  ANDN U2264 ( .B(n1280), .A(n1538), .Z(n1537) );
  XOR U2265 ( .A(n1539), .B(n1284), .Z(out[880]) );
  XOR U2266 ( .A(n1541), .B(n1542), .Z(out[87]) );
  NOR U2267 ( .A(n1543), .B(n1544), .Z(n1541) );
  XOR U2268 ( .A(n1545), .B(n1288), .Z(out[879]) );
  XOR U2269 ( .A(n1547), .B(n1291), .Z(out[878]) );
  AND U2270 ( .A(n1292), .B(n1548), .Z(n1547) );
  XOR U2271 ( .A(n1549), .B(n1297), .Z(out[877]) );
  XOR U2272 ( .A(n1551), .B(n1301), .Z(out[876]) );
  XOR U2273 ( .A(n1553), .B(n1309), .Z(out[875]) );
  ANDN U2274 ( .B(n1554), .A(n1308), .Z(n1553) );
  XOR U2275 ( .A(n1555), .B(n1313), .Z(out[874]) );
  XOR U2276 ( .A(n1557), .B(n1317), .Z(out[873]) );
  AND U2277 ( .A(n1316), .B(n1558), .Z(n1557) );
  XOR U2278 ( .A(n1559), .B(n1321), .Z(out[872]) );
  XOR U2279 ( .A(n1560), .B(n1325), .Z(out[871]) );
  XNOR U2280 ( .A(n1562), .B(n1328), .Z(out[870]) );
  XOR U2281 ( .A(n1564), .B(n1565), .Z(out[86]) );
  XNOR U2282 ( .A(n1568), .B(n1333), .Z(out[869]) );
  ANDN U2283 ( .B(n1569), .A(n1332), .Z(n1568) );
  XOR U2284 ( .A(n1570), .B(n1337), .Z(out[868]) );
  NOR U2285 ( .A(n1571), .B(n1336), .Z(n1570) );
  XOR U2286 ( .A(n1572), .B(n1341), .Z(out[867]) );
  ANDN U2287 ( .B(n1573), .A(n1340), .Z(n1572) );
  XOR U2288 ( .A(n1574), .B(n1345), .Z(out[866]) );
  ANDN U2289 ( .B(n1575), .A(n1344), .Z(n1574) );
  XOR U2290 ( .A(n1576), .B(n1353), .Z(out[865]) );
  ANDN U2291 ( .B(n1577), .A(n1352), .Z(n1576) );
  XOR U2292 ( .A(n1578), .B(n1357), .Z(out[864]) );
  NOR U2293 ( .A(n1356), .B(n1579), .Z(n1578) );
  XOR U2294 ( .A(n1580), .B(n1361), .Z(out[863]) );
  ANDN U2295 ( .B(n1581), .A(n1360), .Z(n1580) );
  XOR U2296 ( .A(n1582), .B(n1365), .Z(out[862]) );
  ANDN U2297 ( .B(n1583), .A(n1364), .Z(n1582) );
  XOR U2298 ( .A(n1584), .B(n1369), .Z(out[861]) );
  NOR U2299 ( .A(n1585), .B(n1368), .Z(n1584) );
  XOR U2300 ( .A(n1586), .B(n1373), .Z(out[860]) );
  ANDN U2301 ( .B(n1587), .A(n1372), .Z(n1586) );
  XNOR U2302 ( .A(n1588), .B(n1589), .Z(out[85]) );
  AND U2303 ( .A(n1590), .B(n1591), .Z(n1588) );
  XOR U2304 ( .A(n1592), .B(n1377), .Z(out[859]) );
  ANDN U2305 ( .B(n1593), .A(n1376), .Z(n1592) );
  XOR U2306 ( .A(n1594), .B(n1381), .Z(out[858]) );
  ANDN U2307 ( .B(n1595), .A(n1380), .Z(n1594) );
  XOR U2308 ( .A(n1596), .B(n1385), .Z(out[857]) );
  ANDN U2309 ( .B(n1597), .A(n1384), .Z(n1596) );
  XOR U2310 ( .A(n1598), .B(n1389), .Z(out[856]) );
  XNOR U2311 ( .A(n1600), .B(n1397), .Z(out[855]) );
  ANDN U2312 ( .B(n1601), .A(n1396), .Z(n1600) );
  XNOR U2313 ( .A(n1602), .B(n1400), .Z(out[854]) );
  XNOR U2314 ( .A(n1604), .B(n1404), .Z(out[853]) );
  AND U2315 ( .A(n1605), .B(n1606), .Z(n1604) );
  XOR U2316 ( .A(n1607), .B(n1409), .Z(out[852]) );
  XNOR U2317 ( .A(n1609), .B(n1412), .Z(out[851]) );
  AND U2318 ( .A(n1610), .B(n1413), .Z(n1609) );
  XNOR U2319 ( .A(n1611), .B(n1416), .Z(out[850]) );
  AND U2320 ( .A(n1417), .B(n1612), .Z(n1611) );
  XNOR U2321 ( .A(n1613), .B(n1614), .Z(out[84]) );
  NOR U2322 ( .A(n1615), .B(n1616), .Z(n1613) );
  XOR U2323 ( .A(n1617), .B(n1421), .Z(out[849]) );
  ANDN U2324 ( .B(n1618), .A(n1420), .Z(n1617) );
  XOR U2325 ( .A(n1619), .B(n1425), .Z(out[848]) );
  ANDN U2326 ( .B(n1620), .A(n1424), .Z(n1619) );
  XOR U2327 ( .A(n1621), .B(n1429), .Z(out[847]) );
  ANDN U2328 ( .B(n1622), .A(n1428), .Z(n1621) );
  XNOR U2329 ( .A(n1623), .B(n1433), .Z(out[846]) );
  NOR U2330 ( .A(n1624), .B(n1432), .Z(n1623) );
  XOR U2331 ( .A(n1625), .B(n1441), .Z(out[845]) );
  ANDN U2332 ( .B(n1440), .A(n1626), .Z(n1625) );
  XNOR U2333 ( .A(n1627), .B(n1445), .Z(out[844]) );
  NOR U2334 ( .A(n1628), .B(n1444), .Z(n1627) );
  XOR U2335 ( .A(n1629), .B(n1448), .Z(out[843]) );
  AND U2336 ( .A(n1447), .B(n1630), .Z(n1629) );
  XNOR U2337 ( .A(n1631), .B(n1451), .Z(out[842]) );
  XOR U2338 ( .A(n1633), .B(n1455), .Z(out[841]) );
  AND U2339 ( .A(n1456), .B(n1634), .Z(n1633) );
  XNOR U2340 ( .A(n1635), .B(n1459), .Z(out[840]) );
  XOR U2341 ( .A(n1637), .B(n1638), .Z(out[83]) );
  XNOR U2342 ( .A(n1641), .B(n1463), .Z(out[839]) );
  AND U2343 ( .A(n1642), .B(n1464), .Z(n1641) );
  XNOR U2344 ( .A(n1643), .B(n1467), .Z(out[838]) );
  AND U2345 ( .A(n1468), .B(n1644), .Z(n1643) );
  XNOR U2346 ( .A(n1645), .B(n1472), .Z(out[837]) );
  ANDN U2347 ( .B(n1646), .A(n1471), .Z(n1645) );
  XNOR U2348 ( .A(n1647), .B(n1475), .Z(out[836]) );
  AND U2349 ( .A(n1476), .B(n1648), .Z(n1647) );
  XNOR U2350 ( .A(n1649), .B(n1487), .Z(out[835]) );
  AND U2351 ( .A(n1488), .B(n1650), .Z(n1649) );
  XNOR U2352 ( .A(n1651), .B(n1491), .Z(out[834]) );
  AND U2353 ( .A(n1652), .B(n1653), .Z(n1651) );
  XNOR U2354 ( .A(n1654), .B(n1495), .Z(out[833]) );
  AND U2355 ( .A(n1655), .B(n1496), .Z(n1654) );
  XNOR U2356 ( .A(n1656), .B(n1499), .Z(out[832]) );
  XOR U2357 ( .A(n1658), .B(n1220), .Z(out[831]) );
  IV U2358 ( .A(n1503), .Z(n1220) );
  XOR U2359 ( .A(n1659), .B(n1660), .Z(n1503) );
  ANDN U2360 ( .B(n1661), .A(n1502), .Z(n1658) );
  XOR U2361 ( .A(n1662), .B(n1223), .Z(out[830]) );
  XOR U2362 ( .A(n1663), .B(n1664), .Z(n1223) );
  ANDN U2363 ( .B(n1665), .A(n1505), .Z(n1662) );
  XNOR U2364 ( .A(n1666), .B(n1667), .Z(out[82]) );
  XNOR U2365 ( .A(n1670), .B(n1228), .Z(out[829]) );
  XNOR U2366 ( .A(n1671), .B(n1672), .Z(n1228) );
  AND U2367 ( .A(n1673), .B(n1674), .Z(n1670) );
  XNOR U2368 ( .A(n1675), .B(n1232), .Z(out[828]) );
  XNOR U2369 ( .A(n1676), .B(n1677), .Z(n1232) );
  AND U2370 ( .A(n1678), .B(n1679), .Z(n1675) );
  XOR U2371 ( .A(n1680), .B(n1235), .Z(out[827]) );
  XOR U2372 ( .A(n1681), .B(n1682), .Z(n1235) );
  ANDN U2373 ( .B(n1683), .A(n1511), .Z(n1680) );
  XOR U2374 ( .A(n1684), .B(n1240), .Z(out[826]) );
  IV U2375 ( .A(n1514), .Z(n1240) );
  XNOR U2376 ( .A(n1685), .B(n1686), .Z(n1514) );
  ANDN U2377 ( .B(n1687), .A(n1513), .Z(n1684) );
  XOR U2378 ( .A(n1688), .B(n1244), .Z(out[825]) );
  IV U2379 ( .A(n1521), .Z(n1244) );
  XNOR U2380 ( .A(n1689), .B(n1690), .Z(n1521) );
  ANDN U2381 ( .B(n1691), .A(n1520), .Z(n1688) );
  XOR U2382 ( .A(n1692), .B(n1247), .Z(out[824]) );
  XOR U2383 ( .A(n1693), .B(n1694), .Z(n1247) );
  ANDN U2384 ( .B(n1695), .A(n1523), .Z(n1692) );
  XNOR U2385 ( .A(n1696), .B(n1251), .Z(out[823]) );
  XNOR U2386 ( .A(n1697), .B(n1698), .Z(n1251) );
  AND U2387 ( .A(n1699), .B(n1700), .Z(n1696) );
  XOR U2388 ( .A(n1701), .B(n1255), .Z(out[822]) );
  IV U2389 ( .A(n1528), .Z(n1255) );
  XNOR U2390 ( .A(n1702), .B(n1703), .Z(n1528) );
  XNOR U2391 ( .A(n1705), .B(n1264), .Z(out[821]) );
  XOR U2392 ( .A(n1706), .B(n1707), .Z(n1264) );
  ANDN U2393 ( .B(n1708), .A(n1530), .Z(n1705) );
  XNOR U2394 ( .A(n1709), .B(n1268), .Z(out[820]) );
  XOR U2395 ( .A(n1710), .B(n1711), .Z(n1268) );
  AND U2396 ( .A(n1712), .B(n1713), .Z(n1709) );
  XNOR U2397 ( .A(n1714), .B(n1715), .Z(out[81]) );
  XNOR U2398 ( .A(n1718), .B(n1272), .Z(out[819]) );
  XNOR U2399 ( .A(n1719), .B(n1720), .Z(n1272) );
  NOR U2400 ( .A(n1534), .B(n1721), .Z(n1718) );
  IV U2401 ( .A(n1722), .Z(n1534) );
  XOR U2402 ( .A(n1723), .B(n1275), .Z(out[818]) );
  XOR U2403 ( .A(n1724), .B(n1725), .Z(n1275) );
  AND U2404 ( .A(n1726), .B(n1536), .Z(n1723) );
  XNOR U2405 ( .A(n1727), .B(n1280), .Z(out[817]) );
  XNOR U2406 ( .A(n1728), .B(n1729), .Z(n1280) );
  XOR U2407 ( .A(n1731), .B(n1283), .Z(out[816]) );
  XNOR U2408 ( .A(n1732), .B(n1733), .Z(n1283) );
  AND U2409 ( .A(n1734), .B(n1735), .Z(n1731) );
  XOR U2410 ( .A(n1736), .B(n1287), .Z(out[815]) );
  XNOR U2411 ( .A(n1737), .B(n1738), .Z(n1287) );
  XNOR U2412 ( .A(n1740), .B(n1292), .Z(out[814]) );
  XOR U2413 ( .A(n1741), .B(n1742), .Z(n1292) );
  AND U2414 ( .A(n1743), .B(n1744), .Z(n1740) );
  XOR U2415 ( .A(n1745), .B(n1295), .Z(out[813]) );
  XNOR U2416 ( .A(n1746), .B(n1747), .Z(n1295) );
  AND U2417 ( .A(n1748), .B(n1749), .Z(n1745) );
  XOR U2418 ( .A(n1750), .B(n1300), .Z(out[812]) );
  XOR U2419 ( .A(n1751), .B(n1752), .Z(n1300) );
  AND U2420 ( .A(n1753), .B(n1754), .Z(n1750) );
  XOR U2421 ( .A(n1755), .B(n1308), .Z(out[811]) );
  XNOR U2422 ( .A(n1756), .B(n1757), .Z(n1308) );
  AND U2423 ( .A(n1758), .B(n1759), .Z(n1755) );
  XOR U2424 ( .A(n1760), .B(n1312), .Z(out[810]) );
  XOR U2425 ( .A(n1761), .B(n1762), .Z(n1312) );
  ANDN U2426 ( .B(n1763), .A(n1556), .Z(n1760) );
  XNOR U2427 ( .A(n1764), .B(n1765), .Z(out[80]) );
  ANDN U2428 ( .B(n1766), .A(n1767), .Z(n1764) );
  XNOR U2429 ( .A(n1768), .B(n1316), .Z(out[809]) );
  XNOR U2430 ( .A(n1769), .B(n1770), .Z(n1316) );
  AND U2431 ( .A(n1771), .B(n1772), .Z(n1768) );
  XOR U2432 ( .A(n1773), .B(n1320), .Z(out[808]) );
  XOR U2433 ( .A(n1774), .B(n1775), .Z(n1320) );
  AND U2434 ( .A(n1776), .B(n1777), .Z(n1773) );
  XOR U2435 ( .A(n1778), .B(n1324), .Z(out[807]) );
  XOR U2436 ( .A(n1779), .B(n1780), .Z(n1324) );
  ANDN U2437 ( .B(n1781), .A(n1561), .Z(n1778) );
  XOR U2438 ( .A(n1782), .B(n1329), .Z(out[806]) );
  XOR U2439 ( .A(n1783), .B(n1784), .Z(n1329) );
  ANDN U2440 ( .B(n1785), .A(n1563), .Z(n1782) );
  XOR U2441 ( .A(n1786), .B(n1332), .Z(out[805]) );
  XNOR U2442 ( .A(n1787), .B(n1788), .Z(n1332) );
  AND U2443 ( .A(n1789), .B(n1790), .Z(n1786) );
  XOR U2444 ( .A(n1791), .B(n1336), .Z(out[804]) );
  XNOR U2445 ( .A(n1792), .B(n1793), .Z(n1336) );
  AND U2446 ( .A(n1571), .B(n1794), .Z(n1791) );
  XOR U2447 ( .A(n1795), .B(n1340), .Z(out[803]) );
  XOR U2448 ( .A(n1796), .B(n1797), .Z(n1340) );
  ANDN U2449 ( .B(n1798), .A(n1573), .Z(n1795) );
  XOR U2450 ( .A(n1799), .B(n1344), .Z(out[802]) );
  XNOR U2451 ( .A(n1800), .B(n1801), .Z(n1344) );
  ANDN U2452 ( .B(n1802), .A(n1575), .Z(n1799) );
  XOR U2453 ( .A(n1803), .B(n1352), .Z(out[801]) );
  XNOR U2454 ( .A(n1804), .B(n1805), .Z(n1352) );
  ANDN U2455 ( .B(n1806), .A(n1577), .Z(n1803) );
  XOR U2456 ( .A(n1807), .B(n1356), .Z(out[800]) );
  XNOR U2457 ( .A(n1808), .B(n1809), .Z(n1356) );
  AND U2458 ( .A(n1579), .B(n1810), .Z(n1807) );
  XOR U2459 ( .A(n1811), .B(n1812), .Z(out[7]) );
  NOR U2460 ( .A(n1813), .B(n1814), .Z(n1811) );
  XOR U2461 ( .A(n1815), .B(n1816), .Z(out[79]) );
  NOR U2462 ( .A(n1817), .B(n1818), .Z(n1815) );
  XOR U2463 ( .A(n1819), .B(n1360), .Z(out[799]) );
  XOR U2464 ( .A(n1820), .B(n1821), .Z(n1360) );
  NOR U2465 ( .A(n1822), .B(n1581), .Z(n1819) );
  XOR U2466 ( .A(n1823), .B(n1364), .Z(out[798]) );
  XOR U2467 ( .A(n1824), .B(n1825), .Z(n1364) );
  XOR U2468 ( .A(n1827), .B(n1368), .Z(out[797]) );
  XOR U2469 ( .A(n1828), .B(n1829), .Z(n1368) );
  AND U2470 ( .A(n1585), .B(n1830), .Z(n1827) );
  XOR U2471 ( .A(n1831), .B(n1372), .Z(out[796]) );
  XOR U2472 ( .A(n1832), .B(n1833), .Z(n1372) );
  AND U2473 ( .A(n1834), .B(n1835), .Z(n1831) );
  XOR U2474 ( .A(n1836), .B(n1376), .Z(out[795]) );
  XOR U2475 ( .A(n1837), .B(n1838), .Z(n1376) );
  ANDN U2476 ( .B(n1839), .A(n1593), .Z(n1836) );
  XOR U2477 ( .A(n1840), .B(n1380), .Z(out[794]) );
  XOR U2478 ( .A(n1841), .B(n1842), .Z(n1380) );
  ANDN U2479 ( .B(n1843), .A(n1595), .Z(n1840) );
  XOR U2480 ( .A(n1844), .B(n1384), .Z(out[793]) );
  XOR U2481 ( .A(n1845), .B(n1846), .Z(n1384) );
  AND U2482 ( .A(n1847), .B(n1848), .Z(n1844) );
  XOR U2483 ( .A(n1849), .B(n1388), .Z(out[792]) );
  XOR U2484 ( .A(n1850), .B(n1851), .Z(n1388) );
  ANDN U2485 ( .B(n1852), .A(n1599), .Z(n1849) );
  XOR U2486 ( .A(n1853), .B(n1396), .Z(out[791]) );
  XNOR U2487 ( .A(n1854), .B(n1855), .Z(n1396) );
  NOR U2488 ( .A(n1856), .B(n1601), .Z(n1853) );
  XOR U2489 ( .A(n1857), .B(n1401), .Z(out[790]) );
  XOR U2490 ( .A(n1858), .B(n1859), .Z(n1401) );
  NOR U2491 ( .A(n1860), .B(n1603), .Z(n1857) );
  XNOR U2492 ( .A(n1861), .B(n1862), .Z(out[78]) );
  AND U2493 ( .A(n1863), .B(n1864), .Z(n1861) );
  XOR U2494 ( .A(n1865), .B(n1405), .Z(out[789]) );
  IV U2495 ( .A(n1606), .Z(n1405) );
  XOR U2496 ( .A(n1866), .B(n1867), .Z(n1606) );
  ANDN U2497 ( .B(n1868), .A(n1605), .Z(n1865) );
  XOR U2498 ( .A(n1869), .B(n1408), .Z(out[788]) );
  XOR U2499 ( .A(n1870), .B(n1871), .Z(n1408) );
  ANDN U2500 ( .B(n1872), .A(n1608), .Z(n1869) );
  XNOR U2501 ( .A(n1873), .B(n1413), .Z(out[787]) );
  XOR U2502 ( .A(n1874), .B(n1875), .Z(n1413) );
  ANDN U2503 ( .B(n1876), .A(n1610), .Z(n1873) );
  XNOR U2504 ( .A(n1877), .B(n1417), .Z(out[786]) );
  XNOR U2505 ( .A(n1878), .B(n1879), .Z(n1417) );
  AND U2506 ( .A(n1880), .B(n1881), .Z(n1877) );
  XOR U2507 ( .A(n1882), .B(n1420), .Z(out[785]) );
  XNOR U2508 ( .A(n1883), .B(n1884), .Z(n1420) );
  AND U2509 ( .A(n1885), .B(n1886), .Z(n1882) );
  XOR U2510 ( .A(n1887), .B(n1424), .Z(out[784]) );
  XNOR U2511 ( .A(n1888), .B(n1889), .Z(n1424) );
  XOR U2512 ( .A(n1891), .B(n1428), .Z(out[783]) );
  XNOR U2513 ( .A(n1892), .B(n1893), .Z(n1428) );
  NOR U2514 ( .A(n1894), .B(n1622), .Z(n1891) );
  XOR U2515 ( .A(n1895), .B(n1432), .Z(out[782]) );
  XNOR U2516 ( .A(n1896), .B(n1897), .Z(n1432) );
  ANDN U2517 ( .B(n1624), .A(n1898), .Z(n1895) );
  XNOR U2518 ( .A(n1899), .B(n1440), .Z(out[781]) );
  XNOR U2519 ( .A(n1900), .B(n1901), .Z(n1440) );
  AND U2520 ( .A(n1626), .B(n1902), .Z(n1899) );
  XOR U2521 ( .A(n1903), .B(n1444), .Z(out[780]) );
  XNOR U2522 ( .A(n1904), .B(n1905), .Z(n1444) );
  ANDN U2523 ( .B(n1628), .A(n1906), .Z(n1903) );
  XNOR U2524 ( .A(n1907), .B(n1908), .Z(out[77]) );
  NOR U2525 ( .A(n1909), .B(n1910), .Z(n1907) );
  XNOR U2526 ( .A(n1911), .B(n1447), .Z(out[779]) );
  XOR U2527 ( .A(n1912), .B(n1913), .Z(n1447) );
  AND U2528 ( .A(n1914), .B(n1915), .Z(n1911) );
  XOR U2529 ( .A(n1916), .B(n1452), .Z(out[778]) );
  XOR U2530 ( .A(n1917), .B(n1918), .Z(n1452) );
  ANDN U2531 ( .B(n1919), .A(n1632), .Z(n1916) );
  XNOR U2532 ( .A(n1920), .B(n1456), .Z(out[777]) );
  XNOR U2533 ( .A(n1921), .B(n1922), .Z(n1456) );
  AND U2534 ( .A(n1923), .B(n1924), .Z(n1920) );
  XOR U2535 ( .A(n1925), .B(n1460), .Z(out[776]) );
  XOR U2536 ( .A(n1926), .B(n1927), .Z(n1460) );
  NOR U2537 ( .A(n1928), .B(n1636), .Z(n1925) );
  XNOR U2538 ( .A(n1929), .B(n1464), .Z(out[775]) );
  XOR U2539 ( .A(n1930), .B(n1931), .Z(n1464) );
  ANDN U2540 ( .B(n1932), .A(n1642), .Z(n1929) );
  XNOR U2541 ( .A(n1933), .B(n1468), .Z(out[774]) );
  XOR U2542 ( .A(n1934), .B(n1935), .Z(n1468) );
  AND U2543 ( .A(n1936), .B(n1937), .Z(n1933) );
  XOR U2544 ( .A(n1938), .B(n1471), .Z(out[773]) );
  XOR U2545 ( .A(n1939), .B(n1940), .Z(n1471) );
  XNOR U2546 ( .A(n1942), .B(n1476), .Z(out[772]) );
  XOR U2547 ( .A(n1943), .B(n1944), .Z(n1476) );
  ANDN U2548 ( .B(n1945), .A(n1648), .Z(n1942) );
  XNOR U2549 ( .A(n1946), .B(n1488), .Z(out[771]) );
  XOR U2550 ( .A(n1947), .B(n1948), .Z(n1488) );
  AND U2551 ( .A(n1949), .B(n1950), .Z(n1946) );
  XOR U2552 ( .A(n1951), .B(n1492), .Z(out[770]) );
  IV U2553 ( .A(n1653), .Z(n1492) );
  XOR U2554 ( .A(n1952), .B(n1953), .Z(n1653) );
  ANDN U2555 ( .B(n1954), .A(n1652), .Z(n1951) );
  XNOR U2556 ( .A(n1955), .B(n1956), .Z(out[76]) );
  NOR U2557 ( .A(n1957), .B(n1958), .Z(n1955) );
  XNOR U2558 ( .A(n1959), .B(n1496), .Z(out[769]) );
  XNOR U2559 ( .A(n1960), .B(n1961), .Z(n1496) );
  NOR U2560 ( .A(n1962), .B(n1655), .Z(n1959) );
  XOR U2561 ( .A(n1963), .B(n1500), .Z(out[768]) );
  XOR U2562 ( .A(n1964), .B(n1965), .Z(n1500) );
  XOR U2563 ( .A(n1967), .B(n1502), .Z(out[767]) );
  XOR U2564 ( .A(n1968), .B(n1969), .Z(n1502) );
  NOR U2565 ( .A(n1218), .B(n1661), .Z(n1967) );
  XOR U2566 ( .A(n1970), .B(n1505), .Z(out[766]) );
  XOR U2567 ( .A(n1971), .B(n1972), .Z(n1505) );
  NOR U2568 ( .A(n1665), .B(n1222), .Z(n1970) );
  XOR U2569 ( .A(n1973), .B(n1507), .Z(out[765]) );
  IV U2570 ( .A(n1674), .Z(n1507) );
  XOR U2571 ( .A(n1974), .B(n1975), .Z(n1674) );
  NOR U2572 ( .A(n1226), .B(n1673), .Z(n1973) );
  XOR U2573 ( .A(n1976), .B(n1509), .Z(out[764]) );
  IV U2574 ( .A(n1679), .Z(n1509) );
  XNOR U2575 ( .A(n1977), .B(n1978), .Z(n1679) );
  XOR U2576 ( .A(n1979), .B(n1511), .Z(out[763]) );
  XOR U2577 ( .A(n1980), .B(n1981), .Z(n1511) );
  NOR U2578 ( .A(n1683), .B(n1234), .Z(n1979) );
  XOR U2579 ( .A(n1982), .B(n1513), .Z(out[762]) );
  XOR U2580 ( .A(n1983), .B(n1984), .Z(n1513) );
  NOR U2581 ( .A(n1687), .B(n1238), .Z(n1982) );
  XOR U2582 ( .A(n1985), .B(n1520), .Z(out[761]) );
  XOR U2583 ( .A(n1986), .B(n1987), .Z(n1520) );
  NOR U2584 ( .A(n1242), .B(n1691), .Z(n1985) );
  XOR U2585 ( .A(n1988), .B(n1523), .Z(out[760]) );
  XOR U2586 ( .A(n1989), .B(n1990), .Z(n1523) );
  NOR U2587 ( .A(n1695), .B(n1246), .Z(n1988) );
  XNOR U2588 ( .A(n1991), .B(n1992), .Z(out[75]) );
  NOR U2589 ( .A(n1993), .B(n1994), .Z(n1991) );
  XOR U2590 ( .A(n1995), .B(n1525), .Z(out[759]) );
  IV U2591 ( .A(n1700), .Z(n1525) );
  XOR U2592 ( .A(n1996), .B(n1997), .Z(n1700) );
  XOR U2593 ( .A(n1998), .B(n1527), .Z(out[758]) );
  XOR U2594 ( .A(n1999), .B(n2000), .Z(n1527) );
  XOR U2595 ( .A(n2001), .B(n1530), .Z(out[757]) );
  XOR U2596 ( .A(n2002), .B(n2003), .Z(n1530) );
  XOR U2597 ( .A(n2004), .B(n1532), .Z(out[756]) );
  IV U2598 ( .A(n1713), .Z(n1532) );
  XNOR U2599 ( .A(n2005), .B(n2006), .Z(n1713) );
  NOR U2600 ( .A(n1712), .B(n1266), .Z(n2004) );
  XNOR U2601 ( .A(n2007), .B(n1722), .Z(out[755]) );
  XOR U2602 ( .A(n2008), .B(n2009), .Z(n1722) );
  ANDN U2603 ( .B(n1721), .A(n1270), .Z(n2007) );
  XNOR U2604 ( .A(n2010), .B(n1536), .Z(out[754]) );
  XOR U2605 ( .A(n2011), .B(n2012), .Z(n1536) );
  NOR U2606 ( .A(n1726), .B(n1274), .Z(n2010) );
  XNOR U2607 ( .A(n2013), .B(n1538), .Z(out[753]) );
  XNOR U2608 ( .A(n2014), .B(n2015), .Z(n1538) );
  ANDN U2609 ( .B(n1730), .A(n1278), .Z(n2013) );
  XOR U2610 ( .A(n2016), .B(n1540), .Z(out[752]) );
  IV U2611 ( .A(n1735), .Z(n1540) );
  XOR U2612 ( .A(n2017), .B(n2018), .Z(n1735) );
  NOR U2613 ( .A(n1282), .B(n1734), .Z(n2016) );
  XOR U2614 ( .A(n2019), .B(n1546), .Z(out[751]) );
  XNOR U2615 ( .A(n2020), .B(n2021), .Z(n1546) );
  NOR U2616 ( .A(n1739), .B(n1286), .Z(n2019) );
  XOR U2617 ( .A(n2022), .B(n1548), .Z(out[750]) );
  IV U2618 ( .A(n1744), .Z(n1548) );
  XOR U2619 ( .A(n2023), .B(n2024), .Z(n1744) );
  ANDN U2620 ( .B(n1290), .A(n1743), .Z(n2022) );
  XNOR U2621 ( .A(n2025), .B(n2026), .Z(out[74]) );
  XOR U2622 ( .A(n2029), .B(n1550), .Z(out[749]) );
  IV U2623 ( .A(n1749), .Z(n1550) );
  XOR U2624 ( .A(n2030), .B(n2031), .Z(n1749) );
  NOR U2625 ( .A(n1294), .B(n1748), .Z(n2029) );
  XOR U2626 ( .A(n2032), .B(n1552), .Z(out[748]) );
  IV U2627 ( .A(n1754), .Z(n1552) );
  XOR U2628 ( .A(n2033), .B(n2034), .Z(n1754) );
  NOR U2629 ( .A(n1753), .B(n1299), .Z(n2032) );
  XOR U2630 ( .A(n2035), .B(n1554), .Z(out[747]) );
  IV U2631 ( .A(n1759), .Z(n1554) );
  XNOR U2632 ( .A(n2036), .B(n2037), .Z(n1759) );
  ANDN U2633 ( .B(n1307), .A(n1758), .Z(n2035) );
  IV U2634 ( .A(n2038), .Z(n1307) );
  XOR U2635 ( .A(n2039), .B(n1556), .Z(out[746]) );
  XOR U2636 ( .A(n2040), .B(n2041), .Z(n1556) );
  AND U2637 ( .A(n1311), .B(n2042), .Z(n2039) );
  IV U2638 ( .A(n2043), .Z(n1311) );
  XOR U2639 ( .A(n2044), .B(n1558), .Z(out[745]) );
  IV U2640 ( .A(n1772), .Z(n1558) );
  XOR U2641 ( .A(n2045), .B(n2046), .Z(n1772) );
  ANDN U2642 ( .B(n1315), .A(n1771), .Z(n2044) );
  XOR U2643 ( .A(n2048), .B(n2049), .Z(n1777) );
  NOR U2644 ( .A(n1319), .B(n1776), .Z(n2047) );
  XOR U2645 ( .A(n2050), .B(n1561), .Z(out[743]) );
  XOR U2646 ( .A(n2051), .B(n2052), .Z(n1561) );
  IV U2647 ( .A(n2053), .Z(n1323) );
  XOR U2648 ( .A(n2054), .B(n1563), .Z(out[742]) );
  XOR U2649 ( .A(n2055), .B(n2056), .Z(n1563) );
  NOR U2650 ( .A(n1327), .B(n1785), .Z(n2054) );
  XOR U2651 ( .A(n2057), .B(n1569), .Z(out[741]) );
  IV U2652 ( .A(n1790), .Z(n1569) );
  XOR U2653 ( .A(n2058), .B(n2059), .Z(n1790) );
  NOR U2654 ( .A(n1331), .B(n1789), .Z(n2057) );
  XNOR U2655 ( .A(n2060), .B(n1571), .Z(out[740]) );
  XNOR U2656 ( .A(n2061), .B(n2062), .Z(n1571) );
  AND U2657 ( .A(n1335), .B(n2063), .Z(n2060) );
  IV U2658 ( .A(n2064), .Z(n1335) );
  XNOR U2659 ( .A(n2065), .B(n2066), .Z(out[73]) );
  ANDN U2660 ( .B(n1036), .A(n1034), .Z(n2065) );
  XOR U2661 ( .A(n2067), .B(n1573), .Z(out[739]) );
  XNOR U2662 ( .A(n2068), .B(n2069), .Z(n1573) );
  NOR U2663 ( .A(n1798), .B(n1339), .Z(n2067) );
  XOR U2664 ( .A(n2070), .B(n1575), .Z(out[738]) );
  XNOR U2665 ( .A(n2071), .B(n2072), .Z(n1575) );
  ANDN U2666 ( .B(n1343), .A(n1802), .Z(n2070) );
  IV U2667 ( .A(n2073), .Z(n1343) );
  XOR U2668 ( .A(n2074), .B(n1577), .Z(out[737]) );
  XNOR U2669 ( .A(n2075), .B(n2076), .Z(n1577) );
  NOR U2670 ( .A(n1806), .B(n1351), .Z(n2074) );
  XNOR U2671 ( .A(n2077), .B(n1579), .Z(out[736]) );
  XNOR U2672 ( .A(n2078), .B(n2079), .Z(n1579) );
  NOR U2673 ( .A(n1355), .B(n1810), .Z(n2077) );
  XOR U2674 ( .A(n2080), .B(n1581), .Z(out[735]) );
  XNOR U2675 ( .A(n2081), .B(n2082), .Z(n1581) );
  ANDN U2676 ( .B(n1822), .A(n1359), .Z(n2080) );
  XOR U2677 ( .A(n2083), .B(n1583), .Z(out[734]) );
  XOR U2678 ( .A(n2084), .B(n2085), .Z(n1583) );
  ANDN U2679 ( .B(n1826), .A(n1363), .Z(n2083) );
  XNOR U2680 ( .A(n2086), .B(n1585), .Z(out[733]) );
  XNOR U2681 ( .A(n2087), .B(n2088), .Z(n1585) );
  ANDN U2682 ( .B(n2089), .A(n1830), .Z(n2086) );
  XOR U2683 ( .A(n2090), .B(n1587), .Z(out[732]) );
  IV U2684 ( .A(n1835), .Z(n1587) );
  XOR U2685 ( .A(n2091), .B(n2092), .Z(n1835) );
  NOR U2686 ( .A(n1834), .B(n1371), .Z(n2090) );
  XOR U2687 ( .A(n2093), .B(n1593), .Z(out[731]) );
  XOR U2688 ( .A(n2094), .B(n2095), .Z(n1593) );
  NOR U2689 ( .A(n1375), .B(n1839), .Z(n2093) );
  XOR U2690 ( .A(n2096), .B(n1595), .Z(out[730]) );
  XNOR U2691 ( .A(n2097), .B(n2098), .Z(n1595) );
  ANDN U2692 ( .B(n2099), .A(n1843), .Z(n2096) );
  XNOR U2693 ( .A(n2100), .B(n2101), .Z(out[72]) );
  AND U2694 ( .A(n1480), .B(n2102), .Z(n2100) );
  XOR U2695 ( .A(n2103), .B(n1597), .Z(out[729]) );
  IV U2696 ( .A(n1848), .Z(n1597) );
  XNOR U2697 ( .A(n2104), .B(n2105), .Z(n1848) );
  ANDN U2698 ( .B(n1383), .A(n1847), .Z(n2103) );
  XOR U2699 ( .A(n2106), .B(n1599), .Z(out[728]) );
  XOR U2700 ( .A(n2107), .B(n2108), .Z(n1599) );
  ANDN U2701 ( .B(n2109), .A(n1852), .Z(n2106) );
  XOR U2702 ( .A(n2110), .B(n1601), .Z(out[727]) );
  XNOR U2703 ( .A(n2111), .B(n2112), .Z(n1601) );
  ANDN U2704 ( .B(n1856), .A(n1395), .Z(n2110) );
  XOR U2705 ( .A(n2113), .B(n1603), .Z(out[726]) );
  XOR U2706 ( .A(n2114), .B(n2115), .Z(n1603) );
  AND U2707 ( .A(n1860), .B(n1399), .Z(n2113) );
  IV U2708 ( .A(n2116), .Z(n1399) );
  XOR U2709 ( .A(n2117), .B(n1605), .Z(out[725]) );
  XOR U2710 ( .A(n2118), .B(n2119), .Z(n1605) );
  ANDN U2711 ( .B(n2120), .A(n1403), .Z(n2117) );
  XOR U2712 ( .A(n2121), .B(n1608), .Z(out[724]) );
  XOR U2713 ( .A(n2122), .B(n2123), .Z(n1608) );
  ANDN U2714 ( .B(n1407), .A(n1872), .Z(n2121) );
  IV U2715 ( .A(n2124), .Z(n1407) );
  XOR U2716 ( .A(n2125), .B(n1610), .Z(out[723]) );
  XNOR U2717 ( .A(n2126), .B(n2127), .Z(n1610) );
  NOR U2718 ( .A(n1876), .B(n1411), .Z(n2125) );
  XOR U2719 ( .A(n2128), .B(n1612), .Z(out[722]) );
  IV U2720 ( .A(n1881), .Z(n1612) );
  XOR U2721 ( .A(n2129), .B(n2130), .Z(n1881) );
  NOR U2722 ( .A(n1880), .B(n1415), .Z(n2128) );
  XOR U2723 ( .A(n2131), .B(n1618), .Z(out[721]) );
  IV U2724 ( .A(n1886), .Z(n1618) );
  XNOR U2725 ( .A(n2132), .B(n2133), .Z(n1886) );
  ANDN U2726 ( .B(n1419), .A(n1885), .Z(n2131) );
  XOR U2727 ( .A(n2134), .B(n1620), .Z(out[720]) );
  XNOR U2728 ( .A(n2135), .B(n2136), .Z(n1620) );
  NOR U2729 ( .A(n1890), .B(n1423), .Z(n2134) );
  XNOR U2730 ( .A(n2137), .B(n2138), .Z(out[71]) );
  AND U2731 ( .A(n1814), .B(n2139), .Z(n2137) );
  XOR U2732 ( .A(n2140), .B(n1622), .Z(out[719]) );
  XOR U2733 ( .A(n2141), .B(n2142), .Z(n1622) );
  AND U2734 ( .A(n1894), .B(n2143), .Z(n2140) );
  XNOR U2735 ( .A(n2144), .B(n1624), .Z(out[718]) );
  XNOR U2736 ( .A(n2145), .B(n2146), .Z(n1624) );
  ANDN U2737 ( .B(n1898), .A(n1431), .Z(n2144) );
  XNOR U2738 ( .A(n2147), .B(n1626), .Z(out[717]) );
  XNOR U2739 ( .A(n2148), .B(n2149), .Z(n1626) );
  XNOR U2740 ( .A(n2150), .B(n1628), .Z(out[716]) );
  XOR U2741 ( .A(n2151), .B(n2152), .Z(n1628) );
  ANDN U2742 ( .B(n1906), .A(n1443), .Z(n2150) );
  XOR U2743 ( .A(n2153), .B(n1630), .Z(out[715]) );
  IV U2744 ( .A(n1915), .Z(n1630) );
  XOR U2745 ( .A(n2154), .B(n2155), .Z(n1915) );
  XOR U2746 ( .A(n2157), .B(n1632), .Z(out[714]) );
  XOR U2747 ( .A(n2158), .B(n2159), .Z(n1632) );
  ANDN U2748 ( .B(n2160), .A(n1450), .Z(n2157) );
  XOR U2749 ( .A(n2161), .B(n1634), .Z(out[713]) );
  IV U2750 ( .A(n1924), .Z(n1634) );
  XOR U2751 ( .A(n2162), .B(n2163), .Z(n1924) );
  NOR U2752 ( .A(n1454), .B(n1923), .Z(n2161) );
  XOR U2753 ( .A(n2164), .B(n1636), .Z(out[712]) );
  XOR U2754 ( .A(n2165), .B(n2166), .Z(n1636) );
  ANDN U2755 ( .B(n1928), .A(n1458), .Z(n2164) );
  XOR U2756 ( .A(n2167), .B(n1642), .Z(out[711]) );
  XOR U2757 ( .A(n2168), .B(n2169), .Z(n1642) );
  NOR U2758 ( .A(n1932), .B(n1462), .Z(n2167) );
  XOR U2759 ( .A(n2170), .B(n1644), .Z(out[710]) );
  IV U2760 ( .A(n1937), .Z(n1644) );
  XOR U2761 ( .A(n2171), .B(n2172), .Z(n1937) );
  NOR U2762 ( .A(n1936), .B(n1466), .Z(n2170) );
  XNOR U2763 ( .A(n2173), .B(n2174), .Z(out[70]) );
  XOR U2764 ( .A(n2177), .B(n1646), .Z(out[709]) );
  XNOR U2765 ( .A(n2178), .B(n2179), .Z(n1646) );
  ANDN U2766 ( .B(n1941), .A(n1470), .Z(n2177) );
  XOR U2767 ( .A(n2180), .B(n1648), .Z(out[708]) );
  XNOR U2768 ( .A(n2181), .B(n2182), .Z(n1648) );
  XOR U2769 ( .A(n2183), .B(n1650), .Z(out[707]) );
  IV U2770 ( .A(n1950), .Z(n1650) );
  XOR U2771 ( .A(n2184), .B(n2185), .Z(n1950) );
  NOR U2772 ( .A(n1486), .B(n1949), .Z(n2183) );
  XOR U2773 ( .A(n2186), .B(n1652), .Z(out[706]) );
  XOR U2774 ( .A(n2187), .B(n2188), .Z(n1652) );
  NOR U2775 ( .A(n1490), .B(n1954), .Z(n2186) );
  XOR U2776 ( .A(n2189), .B(n1655), .Z(out[705]) );
  XOR U2777 ( .A(n2190), .B(n2191), .Z(n1655) );
  ANDN U2778 ( .B(n1962), .A(n1494), .Z(n2189) );
  XOR U2779 ( .A(n2192), .B(n1657), .Z(out[704]) );
  XOR U2780 ( .A(n2193), .B(n2194), .Z(n1657) );
  NOR U2781 ( .A(n1966), .B(n1498), .Z(n2192) );
  XOR U2782 ( .A(n2195), .B(n1661), .Z(out[703]) );
  XOR U2783 ( .A(n2196), .B(n2197), .Z(n1661) );
  ANDN U2784 ( .B(n1218), .A(n1219), .Z(n2195) );
  XOR U2785 ( .A(n2198), .B(n2199), .Z(n1219) );
  XNOR U2786 ( .A(n2200), .B(n2201), .Z(n1218) );
  XOR U2787 ( .A(n2202), .B(n1665), .Z(out[702]) );
  XNOR U2788 ( .A(n2203), .B(n2204), .Z(n1665) );
  ANDN U2789 ( .B(n1222), .A(n1224), .Z(n2202) );
  XNOR U2790 ( .A(n2205), .B(n2206), .Z(n1224) );
  XNOR U2791 ( .A(n2207), .B(n2208), .Z(n1222) );
  XOR U2792 ( .A(n2209), .B(n1673), .Z(out[701]) );
  XOR U2793 ( .A(n2210), .B(n2211), .Z(n1673) );
  ANDN U2794 ( .B(n1226), .A(n1227), .Z(n2209) );
  XNOR U2795 ( .A(n2212), .B(n2213), .Z(n1227) );
  XNOR U2796 ( .A(n2214), .B(n2215), .Z(n1226) );
  XOR U2797 ( .A(n2216), .B(n1678), .Z(out[700]) );
  XOR U2798 ( .A(n2217), .B(n2218), .Z(n1678) );
  ANDN U2799 ( .B(n1230), .A(n1231), .Z(n2216) );
  XNOR U2800 ( .A(n2219), .B(n2220), .Z(n1231) );
  XNOR U2801 ( .A(n2221), .B(n2222), .Z(n1230) );
  XOR U2802 ( .A(n2223), .B(n2176), .Z(out[6]) );
  ANDN U2803 ( .B(n2224), .A(n2175), .Z(n2223) );
  XNOR U2804 ( .A(n2225), .B(n2226), .Z(out[69]) );
  XOR U2805 ( .A(n2229), .B(n1683), .Z(out[699]) );
  XOR U2806 ( .A(n2230), .B(n2231), .Z(n1683) );
  AND U2807 ( .A(n1236), .B(n1234), .Z(n2229) );
  XNOR U2808 ( .A(n2232), .B(n2233), .Z(n1234) );
  XNOR U2809 ( .A(n2234), .B(n2235), .Z(n1236) );
  XOR U2810 ( .A(n2236), .B(n1687), .Z(out[698]) );
  XNOR U2811 ( .A(n2237), .B(n2238), .Z(n1687) );
  ANDN U2812 ( .B(n1238), .A(n1239), .Z(n2236) );
  XOR U2813 ( .A(n2239), .B(n2240), .Z(n1239) );
  XNOR U2814 ( .A(n2241), .B(n2242), .Z(n1238) );
  XOR U2815 ( .A(n2243), .B(n1691), .Z(out[697]) );
  XNOR U2816 ( .A(n2244), .B(n2245), .Z(n1691) );
  ANDN U2817 ( .B(n1242), .A(n1243), .Z(n2243) );
  XOR U2818 ( .A(n2246), .B(n2247), .Z(n1243) );
  XOR U2819 ( .A(n2248), .B(n2249), .Z(n1242) );
  XOR U2820 ( .A(n2250), .B(n1695), .Z(out[696]) );
  XOR U2821 ( .A(n2251), .B(n2252), .Z(n1695) );
  ANDN U2822 ( .B(n1246), .A(n1248), .Z(n2250) );
  XNOR U2823 ( .A(n2253), .B(n2254), .Z(n1248) );
  XOR U2824 ( .A(n2255), .B(n2256), .Z(n1246) );
  XOR U2825 ( .A(n2257), .B(n1699), .Z(out[695]) );
  XNOR U2826 ( .A(n2258), .B(n2259), .Z(n1699) );
  AND U2827 ( .A(n1252), .B(n1250), .Z(n2257) );
  XOR U2828 ( .A(n2260), .B(n2261), .Z(n1250) );
  XNOR U2829 ( .A(n2262), .B(n2263), .Z(n1252) );
  XNOR U2830 ( .A(n2264), .B(n1704), .Z(out[694]) );
  XOR U2831 ( .A(n2265), .B(n2266), .Z(n1704) );
  AND U2832 ( .A(n1256), .B(n1254), .Z(n2264) );
  XOR U2833 ( .A(n2267), .B(n2268), .Z(n1254) );
  XNOR U2834 ( .A(n2269), .B(n2270), .Z(n1256) );
  XOR U2835 ( .A(n2271), .B(n1708), .Z(out[693]) );
  XOR U2836 ( .A(n2272), .B(n2273), .Z(n1708) );
  ANDN U2837 ( .B(n1262), .A(n1263), .Z(n2271) );
  XNOR U2838 ( .A(n2274), .B(n2275), .Z(n1263) );
  XNOR U2839 ( .A(n2276), .B(n2277), .Z(n1262) );
  XOR U2840 ( .A(n2278), .B(n1712), .Z(out[692]) );
  XOR U2841 ( .A(n2279), .B(n2280), .Z(n1712) );
  ANDN U2842 ( .B(n1266), .A(n1267), .Z(n2278) );
  XOR U2843 ( .A(n2281), .B(n2282), .Z(n1267) );
  XOR U2844 ( .A(n2283), .B(n2284), .Z(n1266) );
  XNOR U2845 ( .A(n2285), .B(n1721), .Z(out[691]) );
  XNOR U2846 ( .A(n2286), .B(n2287), .Z(n1721) );
  ANDN U2847 ( .B(n1270), .A(n1271), .Z(n2285) );
  XOR U2848 ( .A(n2288), .B(n2289), .Z(n1271) );
  XOR U2849 ( .A(n2290), .B(n2291), .Z(n1270) );
  XOR U2850 ( .A(n2292), .B(n1726), .Z(out[690]) );
  XNOR U2851 ( .A(n2293), .B(n2294), .Z(n1726) );
  ANDN U2852 ( .B(n1274), .A(n1276), .Z(n2292) );
  XNOR U2853 ( .A(n2295), .B(n2296), .Z(n1276) );
  XOR U2854 ( .A(n2297), .B(n2298), .Z(n1274) );
  XOR U2855 ( .A(n2299), .B(n2300), .Z(out[68]) );
  AND U2856 ( .A(n2301), .B(n2302), .Z(n2299) );
  XNOR U2857 ( .A(n2303), .B(n1730), .Z(out[689]) );
  XOR U2858 ( .A(n2304), .B(n2305), .Z(n1730) );
  ANDN U2859 ( .B(n1278), .A(n1279), .Z(n2303) );
  XNOR U2860 ( .A(n2306), .B(n2307), .Z(n1279) );
  XOR U2861 ( .A(n2308), .B(n2309), .Z(n1278) );
  XOR U2862 ( .A(n2310), .B(n1734), .Z(out[688]) );
  XNOR U2863 ( .A(n2311), .B(n2312), .Z(n1734) );
  AND U2864 ( .A(n1282), .B(n1284), .Z(n2310) );
  XOR U2865 ( .A(n2313), .B(n2314), .Z(n1284) );
  XOR U2866 ( .A(n2315), .B(n2316), .Z(n1282) );
  XOR U2867 ( .A(n2317), .B(n1739), .Z(out[687]) );
  XOR U2868 ( .A(n2318), .B(n2319), .Z(n1739) );
  AND U2869 ( .A(n1286), .B(n1288), .Z(n2317) );
  XOR U2870 ( .A(n2320), .B(n2321), .Z(n1288) );
  XNOR U2871 ( .A(n2322), .B(n2323), .Z(n1286) );
  XOR U2872 ( .A(n2324), .B(n1743), .Z(out[686]) );
  XNOR U2873 ( .A(n2325), .B(n2326), .Z(n1743) );
  ANDN U2874 ( .B(n1291), .A(n1290), .Z(n2324) );
  XOR U2875 ( .A(n2327), .B(n2328), .Z(n1290) );
  XNOR U2876 ( .A(n2329), .B(n2330), .Z(n1291) );
  XOR U2877 ( .A(n2331), .B(n1748), .Z(out[685]) );
  XNOR U2878 ( .A(n2332), .B(n2333), .Z(n1748) );
  AND U2879 ( .A(n1297), .B(n1294), .Z(n2331) );
  XOR U2880 ( .A(n2334), .B(n2335), .Z(n1294) );
  XOR U2881 ( .A(n2336), .B(n2337), .Z(n1297) );
  XOR U2882 ( .A(n2338), .B(n1753), .Z(out[684]) );
  XNOR U2883 ( .A(n2339), .B(n2340), .Z(n1753) );
  AND U2884 ( .A(n1299), .B(n1301), .Z(n2338) );
  XOR U2885 ( .A(n2341), .B(n2342), .Z(n1301) );
  XOR U2886 ( .A(n2343), .B(n2344), .Z(n1299) );
  XOR U2887 ( .A(n2345), .B(n1758), .Z(out[683]) );
  XNOR U2888 ( .A(n2346), .B(n2347), .Z(n1758) );
  AND U2889 ( .A(n1309), .B(n2038), .Z(n2345) );
  XNOR U2890 ( .A(n2348), .B(n2349), .Z(n2038) );
  XOR U2891 ( .A(n2350), .B(n2351), .Z(n1309) );
  XOR U2892 ( .A(n2352), .B(n1763), .Z(out[682]) );
  IV U2893 ( .A(n2042), .Z(n1763) );
  XOR U2894 ( .A(n2353), .B(n2354), .Z(n2042) );
  AND U2895 ( .A(n1313), .B(n2043), .Z(n2352) );
  XNOR U2896 ( .A(n2355), .B(n2356), .Z(n2043) );
  XNOR U2897 ( .A(n2357), .B(n2358), .Z(n1313) );
  XOR U2898 ( .A(n2359), .B(n1771), .Z(out[681]) );
  XNOR U2899 ( .A(n2360), .B(n2361), .Z(n1771) );
  ANDN U2900 ( .B(n1317), .A(n1315), .Z(n2359) );
  XNOR U2901 ( .A(n2362), .B(n2363), .Z(n1315) );
  XNOR U2902 ( .A(n2364), .B(n2365), .Z(n1317) );
  XOR U2903 ( .A(n2366), .B(n1776), .Z(out[680]) );
  XOR U2904 ( .A(n2367), .B(n2368), .Z(n1776) );
  AND U2905 ( .A(n1319), .B(n1321), .Z(n2366) );
  XOR U2906 ( .A(n2369), .B(n2370), .Z(n1321) );
  XNOR U2907 ( .A(n2371), .B(n2372), .Z(n1319) );
  XNOR U2908 ( .A(n2373), .B(n2374), .Z(out[67]) );
  XOR U2909 ( .A(n2377), .B(n1781), .Z(out[679]) );
  XOR U2910 ( .A(n2378), .B(n2379), .Z(n1781) );
  AND U2911 ( .A(n1325), .B(n2053), .Z(n2377) );
  XNOR U2912 ( .A(n2380), .B(n2381), .Z(n2053) );
  XNOR U2913 ( .A(n2382), .B(n2383), .Z(n1325) );
  XOR U2914 ( .A(n2384), .B(n1785), .Z(out[678]) );
  XNOR U2915 ( .A(n2385), .B(n2386), .Z(n1785) );
  ANDN U2916 ( .B(n1327), .A(n1328), .Z(n2384) );
  XOR U2917 ( .A(n2387), .B(n2388), .Z(n1328) );
  XNOR U2918 ( .A(n2389), .B(n2390), .Z(n1327) );
  XOR U2919 ( .A(n2391), .B(n1789), .Z(out[677]) );
  XNOR U2920 ( .A(n2392), .B(n2393), .Z(n1789) );
  ANDN U2921 ( .B(n1331), .A(n1333), .Z(n2391) );
  XOR U2922 ( .A(n2394), .B(n2395), .Z(n1333) );
  XNOR U2923 ( .A(n2396), .B(n2397), .Z(n1331) );
  XOR U2924 ( .A(n2398), .B(n1794), .Z(out[676]) );
  IV U2925 ( .A(n2063), .Z(n1794) );
  XNOR U2926 ( .A(n2399), .B(n2400), .Z(n2063) );
  AND U2927 ( .A(n1337), .B(n2064), .Z(n2398) );
  XNOR U2928 ( .A(n2401), .B(n2402), .Z(n2064) );
  XNOR U2929 ( .A(n2403), .B(n2404), .Z(n1337) );
  XOR U2930 ( .A(n2405), .B(n1798), .Z(out[675]) );
  XNOR U2931 ( .A(n2406), .B(n2407), .Z(n1798) );
  AND U2932 ( .A(n1339), .B(n1341), .Z(n2405) );
  XOR U2933 ( .A(n2408), .B(n2409), .Z(n1341) );
  XNOR U2934 ( .A(n2410), .B(n2411), .Z(n1339) );
  XOR U2935 ( .A(n2412), .B(n1802), .Z(out[674]) );
  XNOR U2936 ( .A(n2413), .B(n2414), .Z(n1802) );
  AND U2937 ( .A(n1345), .B(n2073), .Z(n2412) );
  XOR U2938 ( .A(n2415), .B(n2416), .Z(n2073) );
  XNOR U2939 ( .A(n2417), .B(n2418), .Z(n1345) );
  XOR U2940 ( .A(n2419), .B(n1806), .Z(out[673]) );
  XNOR U2941 ( .A(n2420), .B(n2421), .Z(n1806) );
  AND U2942 ( .A(n1351), .B(n1353), .Z(n2419) );
  XOR U2943 ( .A(n2422), .B(n2423), .Z(n1353) );
  XNOR U2944 ( .A(n2424), .B(n2425), .Z(n1351) );
  XOR U2945 ( .A(n2426), .B(n1810), .Z(out[672]) );
  XNOR U2946 ( .A(n2427), .B(n2428), .Z(n1810) );
  AND U2947 ( .A(n1357), .B(n1355), .Z(n2426) );
  XNOR U2948 ( .A(n2429), .B(n2430), .Z(n1355) );
  XNOR U2949 ( .A(n2431), .B(n2432), .Z(n1357) );
  XNOR U2950 ( .A(n2433), .B(n1822), .Z(out[671]) );
  XNOR U2951 ( .A(n2434), .B(n2435), .Z(n1822) );
  AND U2952 ( .A(n1359), .B(n1361), .Z(n2433) );
  XOR U2953 ( .A(n2436), .B(n2437), .Z(n1361) );
  XNOR U2954 ( .A(n2438), .B(n2439), .Z(n1359) );
  XNOR U2955 ( .A(n2440), .B(n1826), .Z(out[670]) );
  XOR U2956 ( .A(n2441), .B(n2442), .Z(n1826) );
  AND U2957 ( .A(n1363), .B(n1365), .Z(n2440) );
  XNOR U2958 ( .A(n2443), .B(n2444), .Z(n1365) );
  XNOR U2959 ( .A(n2445), .B(n2446), .Z(n1363) );
  XNOR U2960 ( .A(n2447), .B(n2448), .Z(out[66]) );
  XOR U2961 ( .A(n2451), .B(n1830), .Z(out[669]) );
  XOR U2962 ( .A(n2452), .B(n2453), .Z(n1830) );
  AND U2963 ( .A(n1369), .B(n1367), .Z(n2451) );
  IV U2964 ( .A(n2089), .Z(n1367) );
  XNOR U2965 ( .A(n2454), .B(n2455), .Z(n2089) );
  XOR U2966 ( .A(n2456), .B(n2457), .Z(n1369) );
  XOR U2967 ( .A(n2458), .B(n1834), .Z(out[668]) );
  XNOR U2968 ( .A(n2459), .B(n2460), .Z(n1834) );
  AND U2969 ( .A(n1371), .B(n1373), .Z(n2458) );
  XOR U2970 ( .A(n2461), .B(n2462), .Z(n1373) );
  XNOR U2971 ( .A(n2463), .B(n2464), .Z(n1371) );
  XOR U2972 ( .A(n2465), .B(n1839), .Z(out[667]) );
  XOR U2973 ( .A(n2466), .B(n2467), .Z(n1839) );
  AND U2974 ( .A(n1375), .B(n1377), .Z(n2465) );
  XNOR U2975 ( .A(n2468), .B(n2469), .Z(n1377) );
  XNOR U2976 ( .A(n2470), .B(n2471), .Z(n1375) );
  XOR U2977 ( .A(n2472), .B(n1843), .Z(out[666]) );
  XNOR U2978 ( .A(n2473), .B(n2474), .Z(n1843) );
  AND U2979 ( .A(n1381), .B(n1379), .Z(n2472) );
  IV U2980 ( .A(n2099), .Z(n1379) );
  XNOR U2981 ( .A(n2475), .B(n2476), .Z(n2099) );
  XNOR U2982 ( .A(n2477), .B(n2478), .Z(n1381) );
  XOR U2983 ( .A(n2479), .B(n1847), .Z(out[665]) );
  XOR U2984 ( .A(n2480), .B(n2481), .Z(n1847) );
  ANDN U2985 ( .B(n1385), .A(n1383), .Z(n2479) );
  XNOR U2986 ( .A(n2482), .B(n2483), .Z(n1383) );
  XOR U2987 ( .A(n2484), .B(n2485), .Z(n1385) );
  XOR U2988 ( .A(n2486), .B(n1852), .Z(out[664]) );
  XOR U2989 ( .A(n2487), .B(n2488), .Z(n1852) );
  AND U2990 ( .A(n1389), .B(n1387), .Z(n2486) );
  IV U2991 ( .A(n2109), .Z(n1387) );
  XNOR U2992 ( .A(n2489), .B(n2490), .Z(n2109) );
  XOR U2993 ( .A(n2491), .B(n2492), .Z(n1389) );
  XNOR U2994 ( .A(n2493), .B(n1856), .Z(out[663]) );
  XOR U2995 ( .A(n2494), .B(n2495), .Z(n1856) );
  ANDN U2996 ( .B(n1395), .A(n1397), .Z(n2493) );
  XOR U2997 ( .A(n2496), .B(n2497), .Z(n1397) );
  XNOR U2998 ( .A(n2498), .B(n2499), .Z(n1395) );
  XNOR U2999 ( .A(n2500), .B(n1860), .Z(out[662]) );
  XNOR U3000 ( .A(n2501), .B(n2502), .Z(n1860) );
  ANDN U3001 ( .B(n2116), .A(n1400), .Z(n2500) );
  XOR U3002 ( .A(n2503), .B(n2504), .Z(n1400) );
  XOR U3003 ( .A(n2505), .B(n2506), .Z(n2116) );
  XOR U3004 ( .A(n2507), .B(n1868), .Z(out[661]) );
  IV U3005 ( .A(n2120), .Z(n1868) );
  XOR U3006 ( .A(n2508), .B(n2509), .Z(n2120) );
  ANDN U3007 ( .B(n1403), .A(n1404), .Z(n2507) );
  XOR U3008 ( .A(n2510), .B(n2511), .Z(n1404) );
  XOR U3009 ( .A(n2512), .B(n2513), .Z(n1403) );
  XOR U3010 ( .A(n2514), .B(n1872), .Z(out[660]) );
  XOR U3011 ( .A(n2515), .B(n2516), .Z(n1872) );
  AND U3012 ( .A(n1409), .B(n2124), .Z(n2514) );
  XNOR U3013 ( .A(n2517), .B(n2518), .Z(n2124) );
  XOR U3014 ( .A(n2519), .B(n2520), .Z(n1409) );
  XNOR U3015 ( .A(n2521), .B(n2522), .Z(out[65]) );
  AND U3016 ( .A(n2523), .B(n2524), .Z(n2521) );
  XOR U3017 ( .A(n2525), .B(n1876), .Z(out[659]) );
  XOR U3018 ( .A(n2526), .B(n2527), .Z(n1876) );
  ANDN U3019 ( .B(n1411), .A(n1412), .Z(n2525) );
  XNOR U3020 ( .A(n2528), .B(n2529), .Z(n1412) );
  XNOR U3021 ( .A(n2530), .B(n2531), .Z(n1411) );
  XOR U3022 ( .A(n2532), .B(n1880), .Z(out[658]) );
  XNOR U3023 ( .A(n2533), .B(n2534), .Z(n1880) );
  ANDN U3024 ( .B(n1415), .A(n1416), .Z(n2532) );
  XNOR U3025 ( .A(n2535), .B(n2536), .Z(n1416) );
  XNOR U3026 ( .A(n2537), .B(n2538), .Z(n1415) );
  XOR U3027 ( .A(n2539), .B(n1885), .Z(out[657]) );
  XNOR U3028 ( .A(n2540), .B(n2541), .Z(n1885) );
  ANDN U3029 ( .B(n1421), .A(n1419), .Z(n2539) );
  XNOR U3030 ( .A(n2542), .B(n2543), .Z(n1419) );
  XNOR U3031 ( .A(n2544), .B(n2545), .Z(n1421) );
  XOR U3032 ( .A(n2546), .B(n1890), .Z(out[656]) );
  XOR U3033 ( .A(n2547), .B(n2548), .Z(n1890) );
  AND U3034 ( .A(n1425), .B(n1423), .Z(n2546) );
  XNOR U3035 ( .A(n2549), .B(n2550), .Z(n1423) );
  XNOR U3036 ( .A(n2551), .B(n2552), .Z(n1425) );
  XNOR U3037 ( .A(n2553), .B(n1894), .Z(out[655]) );
  XNOR U3038 ( .A(n2554), .B(n2555), .Z(n1894) );
  AND U3039 ( .A(n1429), .B(n1427), .Z(n2553) );
  IV U3040 ( .A(n2143), .Z(n1427) );
  XOR U3041 ( .A(n2556), .B(n2557), .Z(n2143) );
  XNOR U3042 ( .A(n2558), .B(n2559), .Z(n1429) );
  XNOR U3043 ( .A(n2560), .B(n1898), .Z(out[654]) );
  XOR U3044 ( .A(n2561), .B(n2562), .Z(n1898) );
  ANDN U3045 ( .B(n1431), .A(n1433), .Z(n2560) );
  XOR U3046 ( .A(n2563), .B(n2564), .Z(n1433) );
  XNOR U3047 ( .A(n2565), .B(n2566), .Z(n1431) );
  XOR U3048 ( .A(n2567), .B(n1902), .Z(out[653]) );
  AND U3049 ( .A(n1441), .B(n1439), .Z(n2567) );
  XOR U3050 ( .A(n2570), .B(n2571), .Z(n1439) );
  XOR U3051 ( .A(n2572), .B(n2573), .Z(n1441) );
  XNOR U3052 ( .A(n2574), .B(n1906), .Z(out[652]) );
  XNOR U3053 ( .A(n2575), .B(n2576), .Z(n1906) );
  ANDN U3054 ( .B(n1443), .A(n1445), .Z(n2574) );
  XNOR U3055 ( .A(n2577), .B(n2578), .Z(n1445) );
  XNOR U3056 ( .A(n2579), .B(n2580), .Z(n1443) );
  XOR U3057 ( .A(n2581), .B(n1914), .Z(out[651]) );
  XOR U3058 ( .A(n2582), .B(n2583), .Z(n1914) );
  AND U3059 ( .A(n1448), .B(n2156), .Z(n2581) );
  XOR U3060 ( .A(n2584), .B(n2585), .Z(n2156) );
  XNOR U3061 ( .A(n2586), .B(n2587), .Z(n1448) );
  XOR U3062 ( .A(n2588), .B(n1919), .Z(out[650]) );
  IV U3063 ( .A(n2160), .Z(n1919) );
  XOR U3064 ( .A(n2589), .B(n2590), .Z(n2160) );
  ANDN U3065 ( .B(n1450), .A(n1451), .Z(n2588) );
  XNOR U3066 ( .A(n2591), .B(n2592), .Z(n1451) );
  XOR U3067 ( .A(n2593), .B(n2594), .Z(n1450) );
  XNOR U3068 ( .A(n2595), .B(n2596), .Z(out[64]) );
  NOR U3069 ( .A(n2597), .B(n2598), .Z(n2595) );
  XOR U3070 ( .A(n2599), .B(n1923), .Z(out[649]) );
  XOR U3071 ( .A(n2600), .B(n2601), .Z(n1923) );
  AND U3072 ( .A(n1455), .B(n1454), .Z(n2599) );
  XOR U3073 ( .A(n2602), .B(n2603), .Z(n1454) );
  XNOR U3074 ( .A(n2604), .B(n2605), .Z(n1455) );
  XNOR U3075 ( .A(n2606), .B(n1928), .Z(out[648]) );
  XNOR U3076 ( .A(n2607), .B(n2608), .Z(n1928) );
  ANDN U3077 ( .B(n1458), .A(n1459), .Z(n2606) );
  XNOR U3078 ( .A(n2609), .B(n2610), .Z(n1459) );
  XOR U3079 ( .A(n2611), .B(n2612), .Z(n1458) );
  XOR U3080 ( .A(n2613), .B(n1932), .Z(out[647]) );
  XOR U3081 ( .A(n2614), .B(n2615), .Z(n1932) );
  ANDN U3082 ( .B(n1462), .A(n1463), .Z(n2613) );
  XOR U3083 ( .A(n2616), .B(n2617), .Z(n1463) );
  XNOR U3084 ( .A(n2618), .B(n2619), .Z(n1462) );
  XOR U3085 ( .A(n2620), .B(n1936), .Z(out[646]) );
  XOR U3086 ( .A(n2621), .B(n2622), .Z(n1936) );
  ANDN U3087 ( .B(n1466), .A(n1467), .Z(n2620) );
  XOR U3088 ( .A(n2623), .B(n2624), .Z(n1467) );
  XNOR U3089 ( .A(n2625), .B(n2626), .Z(n1466) );
  XNOR U3090 ( .A(n2627), .B(n1941), .Z(out[645]) );
  XOR U3091 ( .A(n2628), .B(n2629), .Z(n1941) );
  ANDN U3092 ( .B(n1470), .A(n1472), .Z(n2627) );
  XOR U3093 ( .A(n2630), .B(n2631), .Z(n1472) );
  XNOR U3094 ( .A(n2632), .B(n2633), .Z(n1470) );
  XOR U3095 ( .A(n2634), .B(n1945), .Z(out[644]) );
  XOR U3096 ( .A(n2635), .B(n2636), .Z(n1945) );
  ANDN U3097 ( .B(n1474), .A(n1475), .Z(n2634) );
  XOR U3098 ( .A(n2637), .B(n2638), .Z(n1475) );
  XNOR U3099 ( .A(n2639), .B(n2640), .Z(n1474) );
  XOR U3100 ( .A(n2641), .B(n1949), .Z(out[643]) );
  XNOR U3101 ( .A(n2642), .B(n2643), .Z(n1949) );
  ANDN U3102 ( .B(n1486), .A(n1487), .Z(n2641) );
  XNOR U3103 ( .A(n2644), .B(n2645), .Z(n1487) );
  XNOR U3104 ( .A(n2646), .B(n2647), .Z(n1486) );
  XOR U3105 ( .A(n2648), .B(n1954), .Z(out[642]) );
  XOR U3106 ( .A(n2649), .B(n2650), .Z(n1954) );
  ANDN U3107 ( .B(n1490), .A(n1491), .Z(n2648) );
  XOR U3108 ( .A(n2651), .B(n2652), .Z(n1491) );
  XOR U3109 ( .A(n2653), .B(n2654), .Z(n1490) );
  XNOR U3110 ( .A(n2655), .B(n1962), .Z(out[641]) );
  XOR U3111 ( .A(n2656), .B(n2657), .Z(n1962) );
  ANDN U3112 ( .B(n1494), .A(n1495), .Z(n2655) );
  XOR U3113 ( .A(n2658), .B(n2659), .Z(n1495) );
  XNOR U3114 ( .A(n2660), .B(n2661), .Z(n1494) );
  XOR U3115 ( .A(n2662), .B(n1966), .Z(out[640]) );
  XNOR U3116 ( .A(n2663), .B(n2664), .Z(n1966) );
  ANDN U3117 ( .B(n1498), .A(n1499), .Z(n2662) );
  XOR U3118 ( .A(n2665), .B(n2666), .Z(n1499) );
  XNOR U3119 ( .A(n2667), .B(n2668), .Z(n1498) );
  XOR U3120 ( .A(n2669), .B(n2670), .Z(out[63]) );
  AND U3121 ( .A(n2671), .B(n2672), .Z(n2669) );
  XNOR U3122 ( .A(n2673), .B(n2674), .Z(out[639]) );
  AND U3123 ( .A(n2675), .B(n2676), .Z(n2673) );
  XOR U3124 ( .A(n2677), .B(n2678), .Z(out[638]) );
  AND U3125 ( .A(n2679), .B(n2680), .Z(n2677) );
  XOR U3126 ( .A(n2681), .B(n2682), .Z(out[637]) );
  NOR U3127 ( .A(n2683), .B(n2684), .Z(n2681) );
  XNOR U3128 ( .A(n2685), .B(n2686), .Z(out[636]) );
  ANDN U3129 ( .B(n2687), .A(n2688), .Z(n2685) );
  XOR U3130 ( .A(n2689), .B(n2690), .Z(out[635]) );
  ANDN U3131 ( .B(n2691), .A(n2692), .Z(n2689) );
  XNOR U3132 ( .A(n2693), .B(n2694), .Z(out[634]) );
  ANDN U3133 ( .B(n2695), .A(n2696), .Z(n2693) );
  XNOR U3134 ( .A(n2697), .B(n2698), .Z(out[633]) );
  AND U3135 ( .A(n2699), .B(n2700), .Z(n2697) );
  XNOR U3136 ( .A(n2701), .B(n2702), .Z(out[632]) );
  AND U3137 ( .A(n2703), .B(n2704), .Z(n2701) );
  XOR U3138 ( .A(n2705), .B(n2706), .Z(out[631]) );
  ANDN U3139 ( .B(n2707), .A(n2708), .Z(n2705) );
  XNOR U3140 ( .A(n2709), .B(n2710), .Z(out[630]) );
  ANDN U3141 ( .B(n2711), .A(n2712), .Z(n2709) );
  XNOR U3142 ( .A(n2713), .B(n2714), .Z(out[62]) );
  AND U3143 ( .A(n2715), .B(n2716), .Z(n2713) );
  XNOR U3144 ( .A(n2717), .B(n2718), .Z(out[629]) );
  AND U3145 ( .A(n2719), .B(n2720), .Z(n2717) );
  XNOR U3146 ( .A(n2721), .B(n2722), .Z(out[628]) );
  ANDN U3147 ( .B(n2723), .A(n2724), .Z(n2721) );
  XNOR U3148 ( .A(n2725), .B(n2726), .Z(out[627]) );
  AND U3149 ( .A(n2727), .B(n2728), .Z(n2725) );
  XOR U3150 ( .A(n2729), .B(n2730), .Z(out[626]) );
  ANDN U3151 ( .B(n2731), .A(n2732), .Z(n2729) );
  XNOR U3152 ( .A(n2733), .B(n2734), .Z(out[625]) );
  AND U3153 ( .A(n2735), .B(n2736), .Z(n2733) );
  XOR U3154 ( .A(n2737), .B(n2738), .Z(out[624]) );
  ANDN U3155 ( .B(n2739), .A(n2740), .Z(n2737) );
  XNOR U3156 ( .A(n2741), .B(n2742), .Z(out[623]) );
  AND U3157 ( .A(n2743), .B(n2744), .Z(n2741) );
  XNOR U3158 ( .A(n2745), .B(n2746), .Z(out[622]) );
  AND U3159 ( .A(n2747), .B(n2748), .Z(n2745) );
  XNOR U3160 ( .A(n2749), .B(n2750), .Z(out[621]) );
  ANDN U3161 ( .B(n2751), .A(n2752), .Z(n2749) );
  XNOR U3162 ( .A(n2753), .B(n2754), .Z(out[620]) );
  NOR U3163 ( .A(n2755), .B(n2756), .Z(n2753) );
  XOR U3164 ( .A(n2757), .B(n2758), .Z(out[61]) );
  AND U3165 ( .A(n2759), .B(n2760), .Z(n2757) );
  XNOR U3166 ( .A(n2761), .B(n2762), .Z(out[619]) );
  AND U3167 ( .A(n2763), .B(n2764), .Z(n2761) );
  XNOR U3168 ( .A(n2765), .B(n2766), .Z(out[618]) );
  AND U3169 ( .A(n2767), .B(n2768), .Z(n2765) );
  XNOR U3170 ( .A(n2769), .B(n2770), .Z(out[617]) );
  AND U3171 ( .A(n2771), .B(n2772), .Z(n2769) );
  XNOR U3172 ( .A(n2773), .B(n2774), .Z(out[616]) );
  ANDN U3173 ( .B(n2775), .A(n2776), .Z(n2773) );
  XNOR U3174 ( .A(n2777), .B(n2778), .Z(out[615]) );
  XOR U3175 ( .A(n2781), .B(n2782), .Z(out[614]) );
  NOR U3176 ( .A(n2783), .B(n2784), .Z(n2781) );
  XNOR U3177 ( .A(n2785), .B(n2786), .Z(out[613]) );
  ANDN U3178 ( .B(n2787), .A(n2788), .Z(n2785) );
  XOR U3179 ( .A(n2789), .B(n2790), .Z(out[612]) );
  AND U3180 ( .A(n2791), .B(n2792), .Z(n2789) );
  XNOR U3181 ( .A(n2793), .B(n2794), .Z(out[611]) );
  AND U3182 ( .A(n2795), .B(n2796), .Z(n2793) );
  XNOR U3183 ( .A(n2797), .B(n2798), .Z(out[610]) );
  AND U3184 ( .A(n2799), .B(n2800), .Z(n2797) );
  XOR U3185 ( .A(n2801), .B(n2802), .Z(out[60]) );
  ANDN U3186 ( .B(n2803), .A(n2804), .Z(n2801) );
  XOR U3187 ( .A(n2805), .B(n2806), .Z(out[609]) );
  NOR U3188 ( .A(n2807), .B(n2808), .Z(n2805) );
  XOR U3189 ( .A(n2809), .B(n2810), .Z(out[608]) );
  ANDN U3190 ( .B(n2811), .A(n2812), .Z(n2809) );
  XNOR U3191 ( .A(n2813), .B(n2814), .Z(out[607]) );
  AND U3192 ( .A(n2815), .B(n2816), .Z(n2813) );
  XNOR U3193 ( .A(n2817), .B(n2818), .Z(out[606]) );
  AND U3194 ( .A(n2819), .B(n2820), .Z(n2817) );
  XNOR U3195 ( .A(n2821), .B(n2822), .Z(out[605]) );
  ANDN U3196 ( .B(n2823), .A(n2824), .Z(n2821) );
  XNOR U3197 ( .A(n2825), .B(n2826), .Z(out[604]) );
  NOR U3198 ( .A(n2827), .B(n2828), .Z(n2825) );
  XNOR U3199 ( .A(n2829), .B(n2830), .Z(out[603]) );
  XNOR U3200 ( .A(n2833), .B(n2834), .Z(out[602]) );
  NOR U3201 ( .A(n2835), .B(n2836), .Z(n2833) );
  XOR U3202 ( .A(n2837), .B(n2838), .Z(out[601]) );
  XNOR U3203 ( .A(n2841), .B(n2842), .Z(out[600]) );
  NOR U3204 ( .A(n2843), .B(n2844), .Z(n2841) );
  XOR U3205 ( .A(n2845), .B(n2228), .Z(out[5]) );
  ANDN U3206 ( .B(n2846), .A(n2227), .Z(n2845) );
  XNOR U3207 ( .A(n2847), .B(n2848), .Z(out[59]) );
  ANDN U3208 ( .B(n2849), .A(n2850), .Z(n2847) );
  XNOR U3209 ( .A(n2851), .B(n2852), .Z(out[599]) );
  NOR U3210 ( .A(n2853), .B(n2854), .Z(n2851) );
  XOR U3211 ( .A(n2855), .B(n2856), .Z(out[598]) );
  ANDN U3212 ( .B(n2857), .A(n2858), .Z(n2855) );
  XNOR U3213 ( .A(n2859), .B(n2860), .Z(out[597]) );
  AND U3214 ( .A(n2861), .B(n2862), .Z(n2859) );
  XNOR U3215 ( .A(n2863), .B(n2864), .Z(out[596]) );
  ANDN U3216 ( .B(n2865), .A(n2866), .Z(n2863) );
  XNOR U3217 ( .A(n2867), .B(n2868), .Z(out[595]) );
  NOR U3218 ( .A(n2869), .B(n2870), .Z(n2867) );
  XNOR U3219 ( .A(n2871), .B(n2872), .Z(out[594]) );
  ANDN U3220 ( .B(n2873), .A(n2874), .Z(n2871) );
  XOR U3221 ( .A(n2875), .B(n2876), .Z(out[593]) );
  ANDN U3222 ( .B(n2877), .A(n2878), .Z(n2875) );
  XNOR U3223 ( .A(n2879), .B(n2880), .Z(out[592]) );
  ANDN U3224 ( .B(n2881), .A(n2882), .Z(n2879) );
  XNOR U3225 ( .A(n2883), .B(n2884), .Z(out[591]) );
  AND U3226 ( .A(n2885), .B(n2886), .Z(n2883) );
  XOR U3227 ( .A(n2887), .B(n2888), .Z(out[590]) );
  ANDN U3228 ( .B(n2889), .A(n2890), .Z(n2887) );
  XOR U3229 ( .A(n2891), .B(n2892), .Z(out[58]) );
  AND U3230 ( .A(n2893), .B(n2894), .Z(n2891) );
  XNOR U3231 ( .A(n2895), .B(n2896), .Z(out[589]) );
  NOR U3232 ( .A(n2897), .B(n2898), .Z(n2895) );
  XNOR U3233 ( .A(n2899), .B(n2900), .Z(out[588]) );
  NOR U3234 ( .A(n2901), .B(n2902), .Z(n2899) );
  XNOR U3235 ( .A(n2903), .B(n2904), .Z(out[587]) );
  ANDN U3236 ( .B(n2905), .A(n2906), .Z(n2903) );
  XNOR U3237 ( .A(n2907), .B(n2908), .Z(out[586]) );
  ANDN U3238 ( .B(n2909), .A(n2910), .Z(n2907) );
  XNOR U3239 ( .A(n2911), .B(n2912), .Z(out[585]) );
  ANDN U3240 ( .B(n2913), .A(n2914), .Z(n2911) );
  XNOR U3241 ( .A(n2915), .B(n2916), .Z(out[584]) );
  ANDN U3242 ( .B(n2917), .A(n2918), .Z(n2915) );
  XNOR U3243 ( .A(n2919), .B(n2920), .Z(out[583]) );
  ANDN U3244 ( .B(n2921), .A(n2922), .Z(n2919) );
  XNOR U3245 ( .A(n2923), .B(n2924), .Z(out[582]) );
  ANDN U3246 ( .B(n2925), .A(n2926), .Z(n2923) );
  XNOR U3247 ( .A(n2927), .B(n2928), .Z(out[581]) );
  AND U3248 ( .A(n2929), .B(n2930), .Z(n2927) );
  XOR U3249 ( .A(n2931), .B(n2932), .Z(out[580]) );
  ANDN U3250 ( .B(n2933), .A(n2934), .Z(n2931) );
  XOR U3251 ( .A(n2935), .B(n2936), .Z(out[57]) );
  ANDN U3252 ( .B(n2937), .A(n2938), .Z(n2935) );
  XNOR U3253 ( .A(n2939), .B(n2940), .Z(out[579]) );
  ANDN U3254 ( .B(n2941), .A(n2942), .Z(n2939) );
  XNOR U3255 ( .A(n2943), .B(n2944), .Z(out[578]) );
  AND U3256 ( .A(n2945), .B(n2946), .Z(n2943) );
  XOR U3257 ( .A(n2947), .B(n2948), .Z(out[577]) );
  AND U3258 ( .A(n2949), .B(n2950), .Z(n2947) );
  XNOR U3259 ( .A(n2951), .B(n2952), .Z(out[576]) );
  ANDN U3260 ( .B(n2953), .A(n2954), .Z(n2951) );
  XNOR U3261 ( .A(n2955), .B(n2676), .Z(out[575]) );
  ANDN U3262 ( .B(n2956), .A(n2675), .Z(n2955) );
  XNOR U3263 ( .A(n2957), .B(n2680), .Z(out[574]) );
  ANDN U3264 ( .B(n2958), .A(n2679), .Z(n2957) );
  XOR U3265 ( .A(n2959), .B(n2684), .Z(out[573]) );
  ANDN U3266 ( .B(n2683), .A(n2960), .Z(n2959) );
  XNOR U3267 ( .A(n2961), .B(n2687), .Z(out[572]) );
  AND U3268 ( .A(n2688), .B(n2962), .Z(n2961) );
  XOR U3269 ( .A(n2963), .B(n2692), .Z(out[571]) );
  XNOR U3270 ( .A(n2965), .B(n2695), .Z(out[570]) );
  AND U3271 ( .A(n2696), .B(n2966), .Z(n2965) );
  XNOR U3272 ( .A(n2967), .B(n2968), .Z(out[56]) );
  XNOR U3273 ( .A(n2971), .B(n2700), .Z(out[569]) );
  ANDN U3274 ( .B(n2972), .A(n2699), .Z(n2971) );
  XNOR U3275 ( .A(n2973), .B(n2704), .Z(out[568]) );
  ANDN U3276 ( .B(n2974), .A(n2703), .Z(n2973) );
  XOR U3277 ( .A(n2975), .B(n2708), .Z(out[567]) );
  AND U3278 ( .A(n2976), .B(n2977), .Z(n2975) );
  XNOR U3279 ( .A(n2978), .B(n2711), .Z(out[566]) );
  AND U3280 ( .A(n2712), .B(n2979), .Z(n2978) );
  XNOR U3281 ( .A(n2980), .B(n2720), .Z(out[565]) );
  ANDN U3282 ( .B(n2981), .A(n2719), .Z(n2980) );
  XNOR U3283 ( .A(n2982), .B(n2723), .Z(out[564]) );
  AND U3284 ( .A(n2724), .B(n2983), .Z(n2982) );
  XNOR U3285 ( .A(n2984), .B(n2727), .Z(out[563]) );
  AND U3286 ( .A(n2985), .B(n2986), .Z(n2984) );
  XNOR U3287 ( .A(n2987), .B(n2731), .Z(out[562]) );
  AND U3288 ( .A(n2732), .B(n2988), .Z(n2987) );
  XNOR U3289 ( .A(n2989), .B(n2736), .Z(out[561]) );
  ANDN U3290 ( .B(n2990), .A(n2735), .Z(n2989) );
  XOR U3291 ( .A(n2991), .B(n2740), .Z(out[560]) );
  AND U3292 ( .A(n2992), .B(n2993), .Z(n2991) );
  XNOR U3293 ( .A(n2994), .B(n2995), .Z(out[55]) );
  AND U3294 ( .A(n2996), .B(n2997), .Z(n2994) );
  XNOR U3295 ( .A(n2998), .B(n2743), .Z(out[559]) );
  AND U3296 ( .A(n2999), .B(n3000), .Z(n2998) );
  XNOR U3297 ( .A(n3001), .B(n2748), .Z(out[558]) );
  ANDN U3298 ( .B(n3002), .A(n2747), .Z(n3001) );
  XOR U3299 ( .A(n3003), .B(n2752), .Z(out[557]) );
  AND U3300 ( .A(n3004), .B(n3005), .Z(n3003) );
  XOR U3301 ( .A(n3006), .B(n2756), .Z(out[556]) );
  AND U3302 ( .A(n2755), .B(n3007), .Z(n3006) );
  XNOR U3303 ( .A(n3008), .B(n2764), .Z(out[555]) );
  ANDN U3304 ( .B(n3009), .A(n2763), .Z(n3008) );
  XNOR U3305 ( .A(n3010), .B(n2767), .Z(out[554]) );
  AND U3306 ( .A(n3011), .B(n3012), .Z(n3010) );
  XNOR U3307 ( .A(n3013), .B(n2772), .Z(out[553]) );
  ANDN U3308 ( .B(n3014), .A(n2771), .Z(n3013) );
  XOR U3309 ( .A(n3015), .B(n2776), .Z(out[552]) );
  XOR U3310 ( .A(n3017), .B(n2779), .Z(out[551]) );
  AND U3311 ( .A(n3018), .B(n2780), .Z(n3017) );
  XOR U3312 ( .A(n3019), .B(n2784), .Z(out[550]) );
  AND U3313 ( .A(n2783), .B(n3020), .Z(n3019) );
  XNOR U3314 ( .A(n3021), .B(n3022), .Z(out[54]) );
  XOR U3315 ( .A(n3025), .B(n2788), .Z(out[549]) );
  AND U3316 ( .A(n3026), .B(n3027), .Z(n3025) );
  XNOR U3317 ( .A(n3028), .B(n2792), .Z(out[548]) );
  ANDN U3318 ( .B(n3029), .A(n2791), .Z(n3028) );
  XNOR U3319 ( .A(n3030), .B(n2796), .Z(out[547]) );
  ANDN U3320 ( .B(n3031), .A(n2795), .Z(n3030) );
  XNOR U3321 ( .A(n3032), .B(n2799), .Z(out[546]) );
  AND U3322 ( .A(n3033), .B(n3034), .Z(n3032) );
  XOR U3323 ( .A(n3035), .B(n2808), .Z(out[545]) );
  AND U3324 ( .A(n2807), .B(n3036), .Z(n3035) );
  XOR U3325 ( .A(n3037), .B(n2812), .Z(out[544]) );
  XNOR U3326 ( .A(n3039), .B(n2816), .Z(out[543]) );
  ANDN U3327 ( .B(n3040), .A(n2815), .Z(n3039) );
  XNOR U3328 ( .A(n3041), .B(n2820), .Z(out[542]) );
  ANDN U3329 ( .B(n3042), .A(n2819), .Z(n3041) );
  XNOR U3330 ( .A(n3043), .B(n2823), .Z(out[541]) );
  AND U3331 ( .A(n2824), .B(n3044), .Z(n3043) );
  XOR U3332 ( .A(n3045), .B(n2827), .Z(out[540]) );
  AND U3333 ( .A(n2828), .B(n3046), .Z(n3045) );
  XNOR U3334 ( .A(n3047), .B(n3048), .Z(out[53]) );
  XOR U3335 ( .A(n3051), .B(n2831), .Z(out[539]) );
  AND U3336 ( .A(n3052), .B(n2832), .Z(n3051) );
  XOR U3337 ( .A(n3053), .B(n2836), .Z(out[538]) );
  AND U3338 ( .A(n2835), .B(n3054), .Z(n3053) );
  XOR U3339 ( .A(n3055), .B(n2839), .Z(out[537]) );
  AND U3340 ( .A(n2840), .B(n3056), .Z(n3055) );
  XOR U3341 ( .A(n3057), .B(n2844), .Z(out[536]) );
  ANDN U3342 ( .B(n2843), .A(n3058), .Z(n3057) );
  XOR U3343 ( .A(n3059), .B(n2854), .Z(out[535]) );
  ANDN U3344 ( .B(n2853), .A(n3060), .Z(n3059) );
  XOR U3345 ( .A(n3061), .B(n2858), .Z(out[534]) );
  AND U3346 ( .A(n3062), .B(n3063), .Z(n3061) );
  XNOR U3347 ( .A(n3064), .B(n2862), .Z(out[533]) );
  XOR U3348 ( .A(n3066), .B(n2866), .Z(out[532]) );
  AND U3349 ( .A(n3067), .B(n3068), .Z(n3066) );
  XOR U3350 ( .A(n3069), .B(n2870), .Z(out[531]) );
  AND U3351 ( .A(n2869), .B(n3070), .Z(n3069) );
  XOR U3352 ( .A(n3071), .B(n2874), .Z(out[530]) );
  XNOR U3353 ( .A(n3073), .B(n3074), .Z(out[52]) );
  AND U3354 ( .A(n3075), .B(n3076), .Z(n3073) );
  XOR U3355 ( .A(n3077), .B(n2878), .Z(out[529]) );
  ANDN U3356 ( .B(n3078), .A(n2877), .Z(n3077) );
  XNOR U3357 ( .A(n3079), .B(n2881), .Z(out[528]) );
  ANDN U3358 ( .B(n2882), .A(n3080), .Z(n3079) );
  XNOR U3359 ( .A(n3081), .B(n2886), .Z(out[527]) );
  NOR U3360 ( .A(n3082), .B(n2885), .Z(n3081) );
  XOR U3361 ( .A(n3083), .B(n2890), .Z(out[526]) );
  XOR U3362 ( .A(n3085), .B(n2898), .Z(out[525]) );
  ANDN U3363 ( .B(n2897), .A(n3086), .Z(n3085) );
  XOR U3364 ( .A(n3087), .B(n2902), .Z(out[524]) );
  AND U3365 ( .A(n2901), .B(n3088), .Z(n3087) );
  XOR U3366 ( .A(n3089), .B(n2906), .Z(out[523]) );
  AND U3367 ( .A(n3090), .B(n3091), .Z(n3089) );
  XNOR U3368 ( .A(n3092), .B(n2909), .Z(out[522]) );
  ANDN U3369 ( .B(n2910), .A(n3093), .Z(n3092) );
  XNOR U3370 ( .A(n3094), .B(n2913), .Z(out[521]) );
  AND U3371 ( .A(n2914), .B(n3095), .Z(n3094) );
  XOR U3372 ( .A(n3096), .B(n2918), .Z(out[520]) );
  ANDN U3373 ( .B(n3097), .A(n2917), .Z(n3096) );
  XNOR U3374 ( .A(n3098), .B(n3099), .Z(out[51]) );
  AND U3375 ( .A(n3100), .B(n3101), .Z(n3098) );
  XOR U3376 ( .A(n3102), .B(n2922), .Z(out[519]) );
  NOR U3377 ( .A(n3103), .B(n2921), .Z(n3102) );
  XOR U3378 ( .A(n3104), .B(n2926), .Z(out[518]) );
  NOR U3379 ( .A(n3105), .B(n2925), .Z(n3104) );
  XNOR U3380 ( .A(n3106), .B(n2930), .Z(out[517]) );
  ANDN U3381 ( .B(n3107), .A(n2929), .Z(n3106) );
  XOR U3382 ( .A(n3108), .B(n2934), .Z(out[516]) );
  ANDN U3383 ( .B(n3109), .A(n2933), .Z(n3108) );
  XNOR U3384 ( .A(n3110), .B(n2941), .Z(out[515]) );
  ANDN U3385 ( .B(n2942), .A(n3111), .Z(n3110) );
  XNOR U3386 ( .A(n3112), .B(n2946), .Z(out[514]) );
  ANDN U3387 ( .B(n3113), .A(n2945), .Z(n3112) );
  XNOR U3388 ( .A(n3114), .B(n2950), .Z(out[513]) );
  NOR U3389 ( .A(n3115), .B(n2949), .Z(n3114) );
  XNOR U3390 ( .A(n3116), .B(n2953), .Z(out[512]) );
  ANDN U3391 ( .B(n2954), .A(n3117), .Z(n3116) );
  XOR U3392 ( .A(n3118), .B(n2675), .Z(out[511]) );
  XOR U3393 ( .A(n3119), .B(n2268), .Z(n2675) );
  AND U3394 ( .A(n3120), .B(n3121), .Z(n3118) );
  XOR U3395 ( .A(n3122), .B(n2679), .Z(out[510]) );
  XOR U3396 ( .A(n3123), .B(n2277), .Z(n2679) );
  AND U3397 ( .A(n3124), .B(n3125), .Z(n3122) );
  XNOR U3398 ( .A(n3126), .B(n3127), .Z(out[50]) );
  AND U3399 ( .A(n3128), .B(n3129), .Z(n3126) );
  XNOR U3400 ( .A(n3130), .B(n2683), .Z(out[509]) );
  XNOR U3401 ( .A(n3131), .B(n3132), .Z(n2683) );
  AND U3402 ( .A(n2960), .B(n3133), .Z(n3130) );
  XNOR U3403 ( .A(n3134), .B(n2688), .Z(out[508]) );
  XNOR U3404 ( .A(n3135), .B(n2291), .Z(n2688) );
  AND U3405 ( .A(n3136), .B(n3137), .Z(n3134) );
  XOR U3406 ( .A(n3138), .B(n2691), .Z(out[507]) );
  XOR U3407 ( .A(n3139), .B(n3140), .Z(n2691) );
  NOR U3408 ( .A(n2964), .B(n3141), .Z(n3138) );
  XNOR U3409 ( .A(n3142), .B(n2696), .Z(out[506]) );
  XNOR U3410 ( .A(n3143), .B(n3144), .Z(n2696) );
  AND U3411 ( .A(n3145), .B(n3146), .Z(n3142) );
  XOR U3412 ( .A(n3147), .B(n2699), .Z(out[505]) );
  XOR U3413 ( .A(n3148), .B(n2316), .Z(n2699) );
  ANDN U3414 ( .B(n3149), .A(n2972), .Z(n3147) );
  XOR U3415 ( .A(n3150), .B(n2703), .Z(out[504]) );
  XNOR U3416 ( .A(n3151), .B(n2323), .Z(n2703) );
  ANDN U3417 ( .B(n3152), .A(n2974), .Z(n3150) );
  XOR U3418 ( .A(n3153), .B(n2707), .Z(out[503]) );
  IV U3419 ( .A(n2977), .Z(n2707) );
  XOR U3420 ( .A(n3154), .B(n2328), .Z(n2977) );
  ANDN U3421 ( .B(n3155), .A(n2976), .Z(n3153) );
  XNOR U3422 ( .A(n3156), .B(n2712), .Z(out[502]) );
  XOR U3423 ( .A(n3157), .B(n2335), .Z(n2712) );
  ANDN U3424 ( .B(n3158), .A(n2979), .Z(n3156) );
  XOR U3425 ( .A(n3159), .B(n2719), .Z(out[501]) );
  XNOR U3426 ( .A(n3160), .B(n3161), .Z(n2719) );
  ANDN U3427 ( .B(n3162), .A(n2981), .Z(n3159) );
  XNOR U3428 ( .A(n3163), .B(n2724), .Z(out[500]) );
  XNOR U3429 ( .A(n3164), .B(n2349), .Z(n2724) );
  ANDN U3430 ( .B(n3165), .A(n2983), .Z(n3163) );
  XNOR U3431 ( .A(n3166), .B(n2302), .Z(out[4]) );
  ANDN U3432 ( .B(n3167), .A(n2301), .Z(n3166) );
  XNOR U3433 ( .A(n3168), .B(n3169), .Z(out[49]) );
  XOR U3434 ( .A(n3172), .B(n2728), .Z(out[499]) );
  IV U3435 ( .A(n2986), .Z(n2728) );
  XNOR U3436 ( .A(n3173), .B(n2356), .Z(n2986) );
  ANDN U3437 ( .B(n3174), .A(n2985), .Z(n3172) );
  XNOR U3438 ( .A(n3175), .B(n2732), .Z(out[498]) );
  XOR U3439 ( .A(n3176), .B(n2363), .Z(n2732) );
  ANDN U3440 ( .B(n3177), .A(n2988), .Z(n3175) );
  XOR U3441 ( .A(n3178), .B(n2735), .Z(out[497]) );
  XNOR U3442 ( .A(n3179), .B(n2372), .Z(n2735) );
  ANDN U3443 ( .B(n3180), .A(n2990), .Z(n3178) );
  XOR U3444 ( .A(n3181), .B(n2739), .Z(out[496]) );
  IV U3445 ( .A(n2993), .Z(n2739) );
  XNOR U3446 ( .A(n3182), .B(n2381), .Z(n2993) );
  ANDN U3447 ( .B(n3183), .A(n2992), .Z(n3181) );
  XOR U3448 ( .A(n3184), .B(n2744), .Z(out[495]) );
  IV U3449 ( .A(n3000), .Z(n2744) );
  XNOR U3450 ( .A(n3185), .B(n2390), .Z(n3000) );
  ANDN U3451 ( .B(n3186), .A(n2999), .Z(n3184) );
  XOR U3452 ( .A(n3187), .B(n2747), .Z(out[494]) );
  XNOR U3453 ( .A(n3188), .B(n2397), .Z(n2747) );
  NOR U3454 ( .A(n3189), .B(n3002), .Z(n3187) );
  XOR U3455 ( .A(n3190), .B(n2751), .Z(out[493]) );
  IV U3456 ( .A(n3005), .Z(n2751) );
  XNOR U3457 ( .A(n3191), .B(n2402), .Z(n3005) );
  NOR U3458 ( .A(n3192), .B(n3004), .Z(n3190) );
  XNOR U3459 ( .A(n3193), .B(n2755), .Z(out[492]) );
  XOR U3460 ( .A(n3194), .B(n2411), .Z(n2755) );
  ANDN U3461 ( .B(n3195), .A(n3007), .Z(n3193) );
  XOR U3462 ( .A(n3196), .B(n2763), .Z(out[491]) );
  XNOR U3463 ( .A(n2415), .B(n3197), .Z(n2763) );
  ANDN U3464 ( .B(n3198), .A(n3009), .Z(n3196) );
  XOR U3465 ( .A(n3199), .B(n2768), .Z(out[490]) );
  IV U3466 ( .A(n3012), .Z(n2768) );
  XNOR U3467 ( .A(n2424), .B(n3200), .Z(n3012) );
  ANDN U3468 ( .B(n3201), .A(n3011), .Z(n3199) );
  XNOR U3469 ( .A(n3202), .B(n3203), .Z(out[48]) );
  AND U3470 ( .A(n3204), .B(n3205), .Z(n3202) );
  XOR U3471 ( .A(n3206), .B(n2771), .Z(out[489]) );
  XNOR U3472 ( .A(n3207), .B(n2430), .Z(n2771) );
  ANDN U3473 ( .B(n3208), .A(n3014), .Z(n3206) );
  XOR U3474 ( .A(n3209), .B(n2775), .Z(out[488]) );
  XOR U3475 ( .A(n3210), .B(n3211), .Z(n2775) );
  ANDN U3476 ( .B(n3212), .A(n3016), .Z(n3209) );
  XNOR U3477 ( .A(n3213), .B(n2780), .Z(out[487]) );
  XOR U3478 ( .A(n3214), .B(n3215), .Z(n2780) );
  ANDN U3479 ( .B(n3216), .A(n3018), .Z(n3213) );
  XNOR U3480 ( .A(n3217), .B(n2783), .Z(out[486]) );
  XOR U3481 ( .A(n3218), .B(n2455), .Z(n2783) );
  XOR U3482 ( .A(n3220), .B(n2787), .Z(out[485]) );
  IV U3483 ( .A(n3027), .Z(n2787) );
  XOR U3484 ( .A(n3221), .B(n3222), .Z(n3027) );
  XOR U3485 ( .A(n3224), .B(n2791), .Z(out[484]) );
  XNOR U3486 ( .A(n3225), .B(n2471), .Z(n2791) );
  NOR U3487 ( .A(n3226), .B(n3029), .Z(n3224) );
  XOR U3488 ( .A(n3227), .B(n2795), .Z(out[483]) );
  XNOR U3489 ( .A(n3228), .B(n2476), .Z(n2795) );
  NOR U3490 ( .A(n3229), .B(n3031), .Z(n3227) );
  XOR U3491 ( .A(n3230), .B(n2800), .Z(out[482]) );
  IV U3492 ( .A(n3034), .Z(n2800) );
  XNOR U3493 ( .A(n3231), .B(n2483), .Z(n3034) );
  ANDN U3494 ( .B(n3232), .A(n3033), .Z(n3230) );
  XNOR U3495 ( .A(n3233), .B(n2807), .Z(out[481]) );
  XOR U3496 ( .A(n3234), .B(n2490), .Z(n2807) );
  ANDN U3497 ( .B(n3235), .A(n3036), .Z(n3233) );
  XOR U3498 ( .A(n3236), .B(n2811), .Z(out[480]) );
  XOR U3499 ( .A(n3237), .B(n2499), .Z(n2811) );
  XNOR U3500 ( .A(n3239), .B(n3240), .Z(out[47]) );
  ANDN U3501 ( .B(n3241), .A(n3242), .Z(n3239) );
  XOR U3502 ( .A(n3243), .B(n2815), .Z(out[479]) );
  XNOR U3503 ( .A(n3244), .B(n2506), .Z(n2815) );
  AND U3504 ( .A(n3245), .B(n3246), .Z(n3243) );
  XOR U3505 ( .A(n3247), .B(n2819), .Z(out[478]) );
  XNOR U3506 ( .A(n3248), .B(n2513), .Z(n2819) );
  XNOR U3507 ( .A(n3250), .B(n2824), .Z(out[477]) );
  XNOR U3508 ( .A(n3251), .B(n2518), .Z(n2824) );
  XNOR U3509 ( .A(n3253), .B(n2828), .Z(out[476]) );
  XNOR U3510 ( .A(n3254), .B(n2531), .Z(n2828) );
  ANDN U3511 ( .B(n3255), .A(n3046), .Z(n3253) );
  XNOR U3512 ( .A(n3256), .B(n2832), .Z(out[475]) );
  XOR U3513 ( .A(n3257), .B(n3258), .Z(n2832) );
  ANDN U3514 ( .B(n3259), .A(n3052), .Z(n3256) );
  XNOR U3515 ( .A(n3260), .B(n2835), .Z(out[474]) );
  XOR U3516 ( .A(n3261), .B(n2543), .Z(n2835) );
  NOR U3517 ( .A(n3262), .B(n3054), .Z(n3260) );
  XNOR U3518 ( .A(n3263), .B(n2840), .Z(out[473]) );
  XOR U3519 ( .A(n3264), .B(n3265), .Z(n2840) );
  AND U3520 ( .A(n3266), .B(n3267), .Z(n3263) );
  XNOR U3521 ( .A(n3268), .B(n2843), .Z(out[472]) );
  XNOR U3522 ( .A(n3269), .B(n2557), .Z(n2843) );
  ANDN U3523 ( .B(n3058), .A(n3270), .Z(n3268) );
  XNOR U3524 ( .A(n3271), .B(n2853), .Z(out[471]) );
  XNOR U3525 ( .A(n3272), .B(n2566), .Z(n2853) );
  ANDN U3526 ( .B(n3060), .A(n3273), .Z(n3271) );
  XOR U3527 ( .A(n3274), .B(n2857), .Z(out[470]) );
  IV U3528 ( .A(n3063), .Z(n2857) );
  XOR U3529 ( .A(n3275), .B(n2571), .Z(n3063) );
  ANDN U3530 ( .B(n3276), .A(n3062), .Z(n3274) );
  XNOR U3531 ( .A(n3277), .B(n3278), .Z(out[46]) );
  ANDN U3532 ( .B(n3279), .A(n3280), .Z(n3277) );
  XOR U3533 ( .A(n3281), .B(n2861), .Z(out[469]) );
  XNOR U3534 ( .A(n3282), .B(n2580), .Z(n2861) );
  AND U3535 ( .A(n3283), .B(n3065), .Z(n3281) );
  XOR U3536 ( .A(n3284), .B(n2865), .Z(out[468]) );
  IV U3537 ( .A(n3068), .Z(n2865) );
  XOR U3538 ( .A(n3285), .B(n2585), .Z(n3068) );
  NOR U3539 ( .A(n3286), .B(n3067), .Z(n3284) );
  XNOR U3540 ( .A(n3287), .B(n2869), .Z(out[467]) );
  XNOR U3541 ( .A(n3288), .B(n2594), .Z(n2869) );
  ANDN U3542 ( .B(n3289), .A(n3070), .Z(n3287) );
  XOR U3543 ( .A(n3290), .B(n2873), .Z(out[466]) );
  XOR U3544 ( .A(n3291), .B(n2603), .Z(n2873) );
  XOR U3545 ( .A(n3293), .B(n2877), .Z(out[465]) );
  XOR U3546 ( .A(n2611), .B(n3294), .Z(n2877) );
  ANDN U3547 ( .B(n3295), .A(n3078), .Z(n3293) );
  XNOR U3548 ( .A(n3296), .B(n2882), .Z(out[464]) );
  XNOR U3549 ( .A(n3297), .B(n3298), .Z(n2882) );
  AND U3550 ( .A(n3080), .B(n3299), .Z(n3296) );
  XOR U3551 ( .A(n3300), .B(n2885), .Z(out[463]) );
  XNOR U3552 ( .A(n3301), .B(n3302), .Z(n2885) );
  AND U3553 ( .A(n3082), .B(n3303), .Z(n3300) );
  XOR U3554 ( .A(n3304), .B(n2889), .Z(out[462]) );
  XOR U3555 ( .A(n3305), .B(n3306), .Z(n2889) );
  ANDN U3556 ( .B(n3307), .A(n3084), .Z(n3304) );
  XNOR U3557 ( .A(n3308), .B(n2897), .Z(out[461]) );
  XNOR U3558 ( .A(n3309), .B(n2640), .Z(n2897) );
  AND U3559 ( .A(n3086), .B(n3310), .Z(n3308) );
  XNOR U3560 ( .A(n3311), .B(n2901), .Z(out[460]) );
  XNOR U3561 ( .A(n3312), .B(n2647), .Z(n2901) );
  AND U3562 ( .A(n3313), .B(n3314), .Z(n3311) );
  XNOR U3563 ( .A(n3315), .B(n3316), .Z(out[45]) );
  AND U3564 ( .A(n3317), .B(n3318), .Z(n3315) );
  XOR U3565 ( .A(n3319), .B(n2905), .Z(out[459]) );
  IV U3566 ( .A(n3091), .Z(n2905) );
  XOR U3567 ( .A(n3320), .B(n2654), .Z(n3091) );
  ANDN U3568 ( .B(n3321), .A(n3090), .Z(n3319) );
  XNOR U3569 ( .A(n3322), .B(n2910), .Z(out[458]) );
  XNOR U3570 ( .A(n3323), .B(n3324), .Z(n2910) );
  AND U3571 ( .A(n3093), .B(n3325), .Z(n3322) );
  XNOR U3572 ( .A(n3326), .B(n2914), .Z(out[457]) );
  XNOR U3573 ( .A(n3327), .B(n2668), .Z(n2914) );
  AND U3574 ( .A(n3328), .B(n3329), .Z(n3326) );
  XOR U3575 ( .A(n3330), .B(n2917), .Z(out[456]) );
  XNOR U3576 ( .A(n3331), .B(n3332), .Z(n2917) );
  AND U3577 ( .A(n3333), .B(n3334), .Z(n3330) );
  XOR U3578 ( .A(n3335), .B(n2921), .Z(out[455]) );
  XNOR U3579 ( .A(n2207), .B(n3336), .Z(n2921) );
  AND U3580 ( .A(n3103), .B(n3337), .Z(n3335) );
  XOR U3581 ( .A(n3338), .B(n2925), .Z(out[454]) );
  XOR U3582 ( .A(n3339), .B(n3340), .Z(n2925) );
  AND U3583 ( .A(n3105), .B(n3341), .Z(n3338) );
  XOR U3584 ( .A(n3342), .B(n2929), .Z(out[453]) );
  XOR U3585 ( .A(n3343), .B(n3344), .Z(n2929) );
  ANDN U3586 ( .B(n3345), .A(n3107), .Z(n3342) );
  XOR U3587 ( .A(n3346), .B(n2933), .Z(out[452]) );
  XNOR U3588 ( .A(n2232), .B(n3347), .Z(n2933) );
  AND U3589 ( .A(n3348), .B(n3349), .Z(n3346) );
  XNOR U3590 ( .A(n3350), .B(n2942), .Z(out[451]) );
  XNOR U3591 ( .A(n3351), .B(n2242), .Z(n2942) );
  AND U3592 ( .A(n3111), .B(n3352), .Z(n3350) );
  XOR U3593 ( .A(n3353), .B(n2945), .Z(out[450]) );
  XNOR U3594 ( .A(n3354), .B(n2249), .Z(n2945) );
  AND U3595 ( .A(n3355), .B(n3356), .Z(n3353) );
  XNOR U3596 ( .A(n3357), .B(n3358), .Z(out[44]) );
  XOR U3597 ( .A(n3361), .B(n2949), .Z(out[449]) );
  XOR U3598 ( .A(n3362), .B(n3363), .Z(n2949) );
  AND U3599 ( .A(n3115), .B(n3364), .Z(n3361) );
  XNOR U3600 ( .A(n3365), .B(n2954), .Z(out[448]) );
  XNOR U3601 ( .A(n3366), .B(n3367), .Z(n2954) );
  AND U3602 ( .A(n3117), .B(n3368), .Z(n3365) );
  XOR U3603 ( .A(n3369), .B(n2956), .Z(out[447]) );
  IV U3604 ( .A(n3121), .Z(n2956) );
  XNOR U3605 ( .A(n3370), .B(n2270), .Z(n3121) );
  NOR U3606 ( .A(n2674), .B(n3120), .Z(n3369) );
  XOR U3607 ( .A(n3371), .B(n2958), .Z(out[446]) );
  IV U3608 ( .A(n3125), .Z(n2958) );
  XNOR U3609 ( .A(n3372), .B(n2275), .Z(n3125) );
  ANDN U3610 ( .B(n2678), .A(n3124), .Z(n3371) );
  XNOR U3611 ( .A(n3373), .B(n2960), .Z(out[445]) );
  XOR U3612 ( .A(n3374), .B(n2282), .Z(n2960) );
  ANDN U3613 ( .B(n2682), .A(n3133), .Z(n3373) );
  XOR U3614 ( .A(n3375), .B(n2962), .Z(out[444]) );
  IV U3615 ( .A(n3137), .Z(n2962) );
  XNOR U3616 ( .A(n3376), .B(n2289), .Z(n3137) );
  NOR U3617 ( .A(n2686), .B(n3136), .Z(n3375) );
  XOR U3618 ( .A(n3377), .B(n2964), .Z(out[443]) );
  XOR U3619 ( .A(n3378), .B(n2296), .Z(n2964) );
  AND U3620 ( .A(n3141), .B(n2690), .Z(n3377) );
  XOR U3621 ( .A(n3379), .B(n2966), .Z(out[442]) );
  IV U3622 ( .A(n3146), .Z(n2966) );
  XNOR U3623 ( .A(n3380), .B(n2307), .Z(n3146) );
  NOR U3624 ( .A(n3145), .B(n2694), .Z(n3379) );
  XOR U3625 ( .A(n3381), .B(n2972), .Z(out[441]) );
  XNOR U3626 ( .A(n3382), .B(n3383), .Z(n2972) );
  ANDN U3627 ( .B(n3384), .A(n2698), .Z(n3381) );
  XOR U3628 ( .A(n3385), .B(n2974), .Z(out[440]) );
  XOR U3629 ( .A(n2320), .B(n3386), .Z(n2974) );
  XOR U3630 ( .A(n3387), .B(n3388), .Z(out[43]) );
  ANDN U3631 ( .B(n3389), .A(n3390), .Z(n3387) );
  XOR U3632 ( .A(n3391), .B(n2976), .Z(out[439]) );
  XOR U3633 ( .A(n3392), .B(n3393), .Z(n2976) );
  ANDN U3634 ( .B(n2706), .A(n3155), .Z(n3391) );
  XOR U3635 ( .A(n3394), .B(n2979), .Z(out[438]) );
  XNOR U3636 ( .A(n3395), .B(n3396), .Z(n2979) );
  NOR U3637 ( .A(n2710), .B(n3158), .Z(n3394) );
  XOR U3638 ( .A(n3397), .B(n2981), .Z(out[437]) );
  XNOR U3639 ( .A(n3398), .B(n3399), .Z(n2981) );
  NOR U3640 ( .A(n2718), .B(n3162), .Z(n3397) );
  XOR U3641 ( .A(n3400), .B(n2983), .Z(out[436]) );
  XNOR U3642 ( .A(n3401), .B(n3402), .Z(n2983) );
  ANDN U3643 ( .B(n3403), .A(n2722), .Z(n3400) );
  XOR U3644 ( .A(n3404), .B(n2985), .Z(out[435]) );
  XNOR U3645 ( .A(n2357), .B(n3405), .Z(n2985) );
  XOR U3646 ( .A(n3406), .B(n2988), .Z(out[434]) );
  XOR U3647 ( .A(n3407), .B(n3408), .Z(n2988) );
  ANDN U3648 ( .B(n2730), .A(n3177), .Z(n3406) );
  XOR U3649 ( .A(n3409), .B(n2990), .Z(out[433]) );
  XOR U3650 ( .A(n2369), .B(n3410), .Z(n2990) );
  NOR U3651 ( .A(n2734), .B(n3180), .Z(n3409) );
  XOR U3652 ( .A(n3411), .B(n2992), .Z(out[432]) );
  XNOR U3653 ( .A(n3412), .B(n3413), .Z(n2992) );
  XOR U3654 ( .A(n3414), .B(n2999), .Z(out[431]) );
  XOR U3655 ( .A(n3415), .B(n2388), .Z(n2999) );
  NOR U3656 ( .A(n2742), .B(n3186), .Z(n3414) );
  XOR U3657 ( .A(n3416), .B(n3002), .Z(out[430]) );
  XNOR U3658 ( .A(n3417), .B(n2395), .Z(n3002) );
  ANDN U3659 ( .B(n3189), .A(n2746), .Z(n3416) );
  XOR U3660 ( .A(n3418), .B(n3419), .Z(out[42]) );
  ANDN U3661 ( .B(n3420), .A(n3421), .Z(n3418) );
  XOR U3662 ( .A(n3422), .B(n3004), .Z(out[429]) );
  XNOR U3663 ( .A(n2403), .B(n3423), .Z(n3004) );
  AND U3664 ( .A(n3192), .B(n3424), .Z(n3422) );
  XOR U3665 ( .A(n3425), .B(n3007), .Z(out[428]) );
  XOR U3666 ( .A(n2408), .B(n3426), .Z(n3007) );
  ANDN U3667 ( .B(n3427), .A(n3195), .Z(n3425) );
  XOR U3668 ( .A(n3428), .B(n3009), .Z(out[427]) );
  XNOR U3669 ( .A(n2417), .B(n3429), .Z(n3009) );
  NOR U3670 ( .A(n3198), .B(n2762), .Z(n3428) );
  XOR U3671 ( .A(n3430), .B(n3011), .Z(out[426]) );
  XOR U3672 ( .A(n2422), .B(n3431), .Z(n3011) );
  NOR U3673 ( .A(n3201), .B(n2766), .Z(n3430) );
  XOR U3674 ( .A(n3432), .B(n3014), .Z(out[425]) );
  XNOR U3675 ( .A(n2431), .B(n3433), .Z(n3014) );
  NOR U3676 ( .A(n2770), .B(n3208), .Z(n3432) );
  XOR U3677 ( .A(n3434), .B(n3016), .Z(out[424]) );
  XOR U3678 ( .A(n2436), .B(n3435), .Z(n3016) );
  XOR U3679 ( .A(n3436), .B(n3018), .Z(out[423]) );
  XNOR U3680 ( .A(n2443), .B(n3437), .Z(n3018) );
  XOR U3681 ( .A(n3438), .B(n3020), .Z(out[422]) );
  XOR U3682 ( .A(n2456), .B(n3439), .Z(n3020) );
  AND U3683 ( .A(n3219), .B(n2782), .Z(n3438) );
  IV U3684 ( .A(n3440), .Z(n2782) );
  XOR U3685 ( .A(n3441), .B(n3026), .Z(out[421]) );
  XOR U3686 ( .A(n2461), .B(n3442), .Z(n3026) );
  ANDN U3687 ( .B(n3443), .A(n3223), .Z(n3441) );
  XOR U3688 ( .A(n3444), .B(n3029), .Z(out[420]) );
  XNOR U3689 ( .A(n2468), .B(n3445), .Z(n3029) );
  AND U3690 ( .A(n3226), .B(n2790), .Z(n3444) );
  IV U3691 ( .A(n3446), .Z(n2790) );
  XNOR U3692 ( .A(n3447), .B(n3448), .Z(out[41]) );
  AND U3693 ( .A(n3449), .B(n3450), .Z(n3447) );
  XOR U3694 ( .A(n3451), .B(n3031), .Z(out[419]) );
  XNOR U3695 ( .A(n2477), .B(n3452), .Z(n3031) );
  ANDN U3696 ( .B(n3229), .A(n2794), .Z(n3451) );
  XOR U3697 ( .A(n3453), .B(n3033), .Z(out[418]) );
  XOR U3698 ( .A(n2484), .B(n3454), .Z(n3033) );
  ANDN U3699 ( .B(n3455), .A(n2798), .Z(n3453) );
  XOR U3700 ( .A(n3456), .B(n3036), .Z(out[417]) );
  XOR U3701 ( .A(n3457), .B(n2492), .Z(n3036) );
  ANDN U3702 ( .B(n2806), .A(n3235), .Z(n3456) );
  IV U3703 ( .A(n3458), .Z(n2806) );
  XOR U3704 ( .A(n3459), .B(n3038), .Z(out[416]) );
  XOR U3705 ( .A(n2496), .B(n3460), .Z(n3038) );
  ANDN U3706 ( .B(n2810), .A(n3238), .Z(n3459) );
  IV U3707 ( .A(n3461), .Z(n2810) );
  XOR U3708 ( .A(n3462), .B(n3040), .Z(out[415]) );
  IV U3709 ( .A(n3246), .Z(n3040) );
  XOR U3710 ( .A(n2503), .B(n3463), .Z(n3246) );
  XOR U3711 ( .A(n3464), .B(n3042), .Z(out[414]) );
  XOR U3712 ( .A(n3465), .B(n3466), .Z(n3042) );
  ANDN U3713 ( .B(n3249), .A(n2818), .Z(n3464) );
  XOR U3714 ( .A(n3467), .B(n3044), .Z(out[413]) );
  XOR U3715 ( .A(n3468), .B(n3469), .Z(n3044) );
  NOR U3716 ( .A(n2822), .B(n3252), .Z(n3467) );
  XOR U3717 ( .A(n3470), .B(n3046), .Z(out[412]) );
  XOR U3718 ( .A(n2528), .B(n3471), .Z(n3046) );
  NOR U3719 ( .A(n3255), .B(n2826), .Z(n3470) );
  XOR U3720 ( .A(n3472), .B(n3052), .Z(out[411]) );
  XNOR U3721 ( .A(n2535), .B(n3473), .Z(n3052) );
  XOR U3722 ( .A(n3474), .B(n3054), .Z(out[410]) );
  XNOR U3723 ( .A(n2544), .B(n3475), .Z(n3054) );
  ANDN U3724 ( .B(n3262), .A(n2834), .Z(n3474) );
  XNOR U3725 ( .A(n3476), .B(n3477), .Z(out[40]) );
  XOR U3726 ( .A(n3480), .B(n3056), .Z(out[409]) );
  IV U3727 ( .A(n3267), .Z(n3056) );
  XOR U3728 ( .A(n3481), .B(n2552), .Z(n3267) );
  ANDN U3729 ( .B(n2838), .A(n3266), .Z(n3480) );
  XNOR U3730 ( .A(n3482), .B(n3058), .Z(out[408]) );
  XNOR U3731 ( .A(n3483), .B(n3484), .Z(n3058) );
  XNOR U3732 ( .A(n3485), .B(n3060), .Z(out[407]) );
  XNOR U3733 ( .A(n3486), .B(n3487), .Z(n3060) );
  AND U3734 ( .A(n3273), .B(n3488), .Z(n3485) );
  XOR U3735 ( .A(n3489), .B(n3062), .Z(out[406]) );
  XOR U3736 ( .A(n3490), .B(n2573), .Z(n3062) );
  ANDN U3737 ( .B(n2856), .A(n3276), .Z(n3489) );
  IV U3738 ( .A(n3491), .Z(n2856) );
  XNOR U3739 ( .A(n3492), .B(n3065), .Z(out[405]) );
  XOR U3740 ( .A(n3493), .B(n2578), .Z(n3065) );
  NOR U3741 ( .A(n2860), .B(n3283), .Z(n3492) );
  XOR U3742 ( .A(n3494), .B(n3067), .Z(out[404]) );
  XOR U3743 ( .A(n3495), .B(n3496), .Z(n3067) );
  XOR U3744 ( .A(n3497), .B(n3070), .Z(out[403]) );
  XOR U3745 ( .A(n3498), .B(n2592), .Z(n3070) );
  NOR U3746 ( .A(n2868), .B(n3289), .Z(n3497) );
  XOR U3747 ( .A(n3499), .B(n3072), .Z(out[402]) );
  XNOR U3748 ( .A(n3500), .B(n3501), .Z(n3072) );
  XOR U3749 ( .A(n3502), .B(n3078), .Z(out[401]) );
  XOR U3750 ( .A(n3503), .B(n2610), .Z(n3078) );
  ANDN U3751 ( .B(n2876), .A(n3295), .Z(n3502) );
  IV U3752 ( .A(n3504), .Z(n2876) );
  XNOR U3753 ( .A(n3505), .B(n3080), .Z(out[400]) );
  XOR U3754 ( .A(n3506), .B(n2617), .Z(n3080) );
  NOR U3755 ( .A(n2880), .B(n3299), .Z(n3505) );
  XOR U3756 ( .A(n3507), .B(n2376), .Z(out[3]) );
  XOR U3757 ( .A(n3509), .B(n3510), .Z(out[39]) );
  ANDN U3758 ( .B(n3511), .A(n3512), .Z(n3509) );
  XNOR U3759 ( .A(n3513), .B(n3082), .Z(out[399]) );
  XOR U3760 ( .A(n3514), .B(n2624), .Z(n3082) );
  XOR U3761 ( .A(n3515), .B(n3084), .Z(out[398]) );
  XNOR U3762 ( .A(n3516), .B(n2631), .Z(n3084) );
  ANDN U3763 ( .B(n2888), .A(n3307), .Z(n3515) );
  IV U3764 ( .A(n3517), .Z(n2888) );
  XNOR U3765 ( .A(n3518), .B(n3086), .Z(out[397]) );
  XOR U3766 ( .A(n3519), .B(n2638), .Z(n3086) );
  ANDN U3767 ( .B(n3520), .A(n3310), .Z(n3518) );
  XOR U3768 ( .A(n3521), .B(n3088), .Z(out[396]) );
  IV U3769 ( .A(n3314), .Z(n3088) );
  XNOR U3770 ( .A(n3522), .B(n2645), .Z(n3314) );
  XOR U3771 ( .A(n3523), .B(n3090), .Z(out[395]) );
  XNOR U3772 ( .A(n3524), .B(n2652), .Z(n3090) );
  XNOR U3773 ( .A(n3525), .B(n3093), .Z(out[394]) );
  XOR U3774 ( .A(n3526), .B(n2659), .Z(n3093) );
  NOR U3775 ( .A(n3325), .B(n2908), .Z(n3525) );
  XOR U3776 ( .A(n3527), .B(n3095), .Z(out[393]) );
  IV U3777 ( .A(n3329), .Z(n3095) );
  XOR U3778 ( .A(n3528), .B(n2666), .Z(n3329) );
  XOR U3779 ( .A(n3529), .B(n3097), .Z(out[392]) );
  IV U3780 ( .A(n3334), .Z(n3097) );
  XOR U3781 ( .A(n3530), .B(n2199), .Z(n3334) );
  XNOR U3782 ( .A(n3531), .B(n3103), .Z(out[391]) );
  XNOR U3783 ( .A(n3532), .B(n2206), .Z(n3103) );
  ANDN U3784 ( .B(n3533), .A(n3337), .Z(n3531) );
  XNOR U3785 ( .A(n3534), .B(n3105), .Z(out[390]) );
  XNOR U3786 ( .A(n3535), .B(n2213), .Z(n3105) );
  NOR U3787 ( .A(n2924), .B(n3341), .Z(n3534) );
  XOR U3788 ( .A(n3536), .B(n3537), .Z(out[38]) );
  ANDN U3789 ( .B(n3538), .A(n3539), .Z(n3536) );
  XOR U3790 ( .A(n3540), .B(n3107), .Z(out[389]) );
  XOR U3791 ( .A(n3541), .B(n2220), .Z(n3107) );
  NOR U3792 ( .A(n2928), .B(n3345), .Z(n3540) );
  XOR U3793 ( .A(n3542), .B(n3109), .Z(out[388]) );
  IV U3794 ( .A(n3349), .Z(n3109) );
  XOR U3795 ( .A(n3543), .B(n2235), .Z(n3349) );
  XNOR U3796 ( .A(n3544), .B(n3111), .Z(out[387]) );
  XOR U3797 ( .A(n3545), .B(n2240), .Z(n3111) );
  NOR U3798 ( .A(n2940), .B(n3352), .Z(n3544) );
  XOR U3799 ( .A(n3546), .B(n3113), .Z(out[386]) );
  IV U3800 ( .A(n3356), .Z(n3113) );
  XOR U3801 ( .A(n3547), .B(n2247), .Z(n3356) );
  NOR U3802 ( .A(n3355), .B(n2944), .Z(n3546) );
  XNOR U3803 ( .A(n3548), .B(n3115), .Z(out[385]) );
  XOR U3804 ( .A(n3549), .B(n2254), .Z(n3115) );
  ANDN U3805 ( .B(n2948), .A(n3364), .Z(n3548) );
  XNOR U3806 ( .A(n3550), .B(n3117), .Z(out[384]) );
  XOR U3807 ( .A(n3551), .B(n2263), .Z(n3117) );
  NOR U3808 ( .A(n2952), .B(n3368), .Z(n3550) );
  XOR U3809 ( .A(n3552), .B(n3120), .Z(out[383]) );
  XNOR U3810 ( .A(n1808), .B(n3553), .Z(n3120) );
  ANDN U3811 ( .B(n2674), .A(n2676), .Z(n3552) );
  XOR U3812 ( .A(n3554), .B(n2333), .Z(n2676) );
  XOR U3813 ( .A(n3555), .B(n2034), .Z(n2674) );
  XOR U3814 ( .A(n3556), .B(n3124), .Z(out[382]) );
  XOR U3815 ( .A(n1820), .B(n3557), .Z(n3124) );
  NOR U3816 ( .A(n2680), .B(n2678), .Z(n3556) );
  XOR U3817 ( .A(n3558), .B(n2037), .Z(n2678) );
  XOR U3818 ( .A(n3559), .B(n2340), .Z(n2680) );
  XOR U3819 ( .A(n3560), .B(n3133), .Z(out[381]) );
  XNOR U3820 ( .A(n3561), .B(n3562), .Z(n3133) );
  ANDN U3821 ( .B(n2684), .A(n2682), .Z(n3560) );
  XOR U3822 ( .A(n3563), .B(n2041), .Z(n2682) );
  XOR U3823 ( .A(n3564), .B(n3565), .Z(n2684) );
  XOR U3824 ( .A(n3566), .B(n3136), .Z(out[380]) );
  XNOR U3825 ( .A(n3567), .B(n3568), .Z(n3136) );
  ANDN U3826 ( .B(n2686), .A(n2687), .Z(n3566) );
  XOR U3827 ( .A(n3569), .B(n2354), .Z(n2687) );
  XOR U3828 ( .A(n3570), .B(n2046), .Z(n2686) );
  XOR U3829 ( .A(n3571), .B(n3572), .Z(out[37]) );
  XNOR U3830 ( .A(n3575), .B(n3141), .Z(out[379]) );
  XNOR U3831 ( .A(n1832), .B(n3576), .Z(n3141) );
  ANDN U3832 ( .B(n2692), .A(n2690), .Z(n3575) );
  XOR U3833 ( .A(n3577), .B(n2049), .Z(n2690) );
  XOR U3834 ( .A(n3578), .B(n3579), .Z(n2692) );
  XOR U3835 ( .A(n3580), .B(n3145), .Z(out[378]) );
  XOR U3836 ( .A(n1837), .B(n3581), .Z(n3145) );
  ANDN U3837 ( .B(n2694), .A(n2695), .Z(n3580) );
  XNOR U3838 ( .A(n3582), .B(n2368), .Z(n2695) );
  XNOR U3839 ( .A(n3583), .B(n2052), .Z(n2694) );
  XOR U3840 ( .A(n3584), .B(n3149), .Z(out[377]) );
  IV U3841 ( .A(n3384), .Z(n3149) );
  XOR U3842 ( .A(n3585), .B(n3586), .Z(n3384) );
  ANDN U3843 ( .B(n2698), .A(n2700), .Z(n3584) );
  XNOR U3844 ( .A(n3587), .B(n2379), .Z(n2700) );
  IV U3845 ( .A(n3588), .Z(n2379) );
  XOR U3846 ( .A(n3589), .B(n2056), .Z(n2698) );
  XOR U3847 ( .A(n3590), .B(n3152), .Z(out[376]) );
  XOR U3848 ( .A(n1845), .B(n3591), .Z(n3152) );
  ANDN U3849 ( .B(n2702), .A(n2704), .Z(n3590) );
  XOR U3850 ( .A(n3592), .B(n2386), .Z(n2704) );
  XOR U3851 ( .A(n3593), .B(n2059), .Z(n2702) );
  XOR U3852 ( .A(n3594), .B(n3155), .Z(out[375]) );
  XOR U3853 ( .A(n1850), .B(n3595), .Z(n3155) );
  ANDN U3854 ( .B(n2708), .A(n2706), .Z(n3594) );
  XOR U3855 ( .A(n3596), .B(n2062), .Z(n2706) );
  XNOR U3856 ( .A(n3597), .B(n3598), .Z(n2708) );
  XOR U3857 ( .A(n3599), .B(n3158), .Z(out[374]) );
  XNOR U3858 ( .A(n1854), .B(n3600), .Z(n3158) );
  ANDN U3859 ( .B(n2710), .A(n2711), .Z(n3599) );
  XOR U3860 ( .A(n3601), .B(n2400), .Z(n2711) );
  XOR U3861 ( .A(n3602), .B(n2069), .Z(n2710) );
  XOR U3862 ( .A(n3603), .B(n3162), .Z(out[373]) );
  XOR U3863 ( .A(n1858), .B(n3604), .Z(n3162) );
  ANDN U3864 ( .B(n2718), .A(n2720), .Z(n3603) );
  XOR U3865 ( .A(n3605), .B(n2407), .Z(n2720) );
  XOR U3866 ( .A(n3606), .B(n2072), .Z(n2718) );
  XOR U3867 ( .A(n3607), .B(n3165), .Z(out[372]) );
  IV U3868 ( .A(n3403), .Z(n3165) );
  XOR U3869 ( .A(n1866), .B(n3608), .Z(n3403) );
  ANDN U3870 ( .B(n2722), .A(n2723), .Z(n3607) );
  XOR U3871 ( .A(n3609), .B(n2414), .Z(n2723) );
  XOR U3872 ( .A(n3610), .B(n2076), .Z(n2722) );
  XOR U3873 ( .A(n3611), .B(n3174), .Z(out[371]) );
  XOR U3874 ( .A(n1870), .B(n3612), .Z(n3174) );
  ANDN U3875 ( .B(n2726), .A(n2727), .Z(n3611) );
  XNOR U3876 ( .A(n3613), .B(n2421), .Z(n2727) );
  XOR U3877 ( .A(n3614), .B(n2079), .Z(n2726) );
  XOR U3878 ( .A(n3615), .B(n3177), .Z(out[370]) );
  XNOR U3879 ( .A(n1874), .B(n3616), .Z(n3177) );
  NOR U3880 ( .A(n2731), .B(n2730), .Z(n3615) );
  XOR U3881 ( .A(n3617), .B(n2082), .Z(n2730) );
  XOR U3882 ( .A(n3618), .B(n2428), .Z(n2731) );
  XOR U3883 ( .A(n3619), .B(n3620), .Z(out[36]) );
  ANDN U3884 ( .B(n3621), .A(n3622), .Z(n3619) );
  XOR U3885 ( .A(n3623), .B(n3180), .Z(out[369]) );
  XNOR U3886 ( .A(n1878), .B(n3624), .Z(n3180) );
  ANDN U3887 ( .B(n2734), .A(n2736), .Z(n3623) );
  XNOR U3888 ( .A(n3625), .B(n2435), .Z(n2736) );
  XNOR U3889 ( .A(n3626), .B(n2085), .Z(n2734) );
  XOR U3890 ( .A(n3627), .B(n3183), .Z(out[368]) );
  XOR U3891 ( .A(n3628), .B(n3629), .Z(n3183) );
  ANDN U3892 ( .B(n2740), .A(n2738), .Z(n3627) );
  XOR U3893 ( .A(n3630), .B(n2088), .Z(n2738) );
  XOR U3894 ( .A(n3631), .B(n3632), .Z(n2740) );
  XOR U3895 ( .A(n3633), .B(n3186), .Z(out[367]) );
  XNOR U3896 ( .A(n3634), .B(n3635), .Z(n3186) );
  ANDN U3897 ( .B(n2742), .A(n2743), .Z(n3633) );
  XNOR U3898 ( .A(n3636), .B(n2453), .Z(n2743) );
  XOR U3899 ( .A(n3637), .B(n2092), .Z(n2742) );
  XNOR U3900 ( .A(n3638), .B(n3189), .Z(out[366]) );
  XNOR U3901 ( .A(n3639), .B(n3640), .Z(n3189) );
  ANDN U3902 ( .B(n2746), .A(n2748), .Z(n3638) );
  XOR U3903 ( .A(n3641), .B(n3642), .Z(n2748) );
  XNOR U3904 ( .A(n2094), .B(n3643), .Z(n2746) );
  XNOR U3905 ( .A(n3644), .B(n3192), .Z(out[365]) );
  XOR U3906 ( .A(n1896), .B(n3645), .Z(n3192) );
  AND U3907 ( .A(n2752), .B(n2750), .Z(n3644) );
  IV U3908 ( .A(n3424), .Z(n2750) );
  XOR U3909 ( .A(n3646), .B(n3647), .Z(n3424) );
  XNOR U3910 ( .A(n3648), .B(n3649), .Z(n2752) );
  XOR U3911 ( .A(n3650), .B(n3195), .Z(out[364]) );
  XOR U3912 ( .A(n1900), .B(n3651), .Z(n3195) );
  AND U3913 ( .A(n2756), .B(n2754), .Z(n3650) );
  IV U3914 ( .A(n3427), .Z(n2754) );
  XNOR U3915 ( .A(n3652), .B(n2105), .Z(n3427) );
  XNOR U3916 ( .A(n3653), .B(n2474), .Z(n2756) );
  IV U3917 ( .A(n3654), .Z(n2474) );
  XOR U3918 ( .A(n3655), .B(n3198), .Z(out[363]) );
  XOR U3919 ( .A(n3656), .B(n3657), .Z(n3198) );
  ANDN U3920 ( .B(n2762), .A(n2764), .Z(n3655) );
  XNOR U3921 ( .A(n3658), .B(n2481), .Z(n2764) );
  XNOR U3922 ( .A(n2107), .B(n3659), .Z(n2762) );
  XOR U3923 ( .A(n3660), .B(n3201), .Z(out[362]) );
  XNOR U3924 ( .A(n1912), .B(n3661), .Z(n3201) );
  ANDN U3925 ( .B(n2766), .A(n2767), .Z(n3660) );
  XOR U3926 ( .A(n3662), .B(n3663), .Z(n2767) );
  XNOR U3927 ( .A(n3664), .B(n3665), .Z(n2766) );
  XOR U3928 ( .A(n3666), .B(n3208), .Z(out[361]) );
  XOR U3929 ( .A(n1917), .B(n3667), .Z(n3208) );
  ANDN U3930 ( .B(n2770), .A(n2772), .Z(n3666) );
  XOR U3931 ( .A(n3668), .B(n2495), .Z(n2772) );
  XNOR U3932 ( .A(n2114), .B(n3669), .Z(n2770) );
  XOR U3933 ( .A(n3670), .B(n3212), .Z(out[360]) );
  XOR U3934 ( .A(n1921), .B(n3671), .Z(n3212) );
  AND U3935 ( .A(n2776), .B(n2774), .Z(n3670) );
  XOR U3936 ( .A(n3672), .B(n3673), .Z(n2774) );
  XOR U3937 ( .A(n3674), .B(n2502), .Z(n2776) );
  XOR U3938 ( .A(n3675), .B(n1040), .Z(out[35]) );
  ANDN U3939 ( .B(n3676), .A(n1039), .Z(n3675) );
  XOR U3940 ( .A(n3677), .B(n3216), .Z(out[359]) );
  XOR U3941 ( .A(n1926), .B(n3678), .Z(n3216) );
  AND U3942 ( .A(n2779), .B(n2778), .Z(n3677) );
  XOR U3943 ( .A(n3679), .B(n3680), .Z(n2778) );
  XNOR U3944 ( .A(n3681), .B(n3682), .Z(n2779) );
  XNOR U3945 ( .A(n3683), .B(n3219), .Z(out[358]) );
  XOR U3946 ( .A(n1930), .B(n3684), .Z(n3219) );
  AND U3947 ( .A(n2784), .B(n3440), .Z(n3683) );
  XOR U3948 ( .A(n2126), .B(n3685), .Z(n3440) );
  XNOR U3949 ( .A(n3686), .B(n3687), .Z(n2784) );
  XOR U3950 ( .A(n3688), .B(n3223), .Z(out[357]) );
  XOR U3951 ( .A(n3689), .B(n3690), .Z(n3223) );
  AND U3952 ( .A(n2788), .B(n2786), .Z(n3688) );
  IV U3953 ( .A(n3443), .Z(n2786) );
  XOR U3954 ( .A(n3691), .B(n2130), .Z(n3443) );
  XNOR U3955 ( .A(n3692), .B(n3693), .Z(n2788) );
  XNOR U3956 ( .A(n3694), .B(n3226), .Z(out[356]) );
  XNOR U3957 ( .A(n1939), .B(n3695), .Z(n3226) );
  ANDN U3958 ( .B(n3446), .A(n2792), .Z(n3694) );
  XOR U3959 ( .A(n3696), .B(n2534), .Z(n2792) );
  XNOR U3960 ( .A(n3697), .B(n2133), .Z(n3446) );
  XNOR U3961 ( .A(n3698), .B(n3229), .Z(out[355]) );
  XOR U3962 ( .A(n1943), .B(n3699), .Z(n3229) );
  ANDN U3963 ( .B(n2794), .A(n2796), .Z(n3698) );
  XOR U3964 ( .A(n3700), .B(n2541), .Z(n2796) );
  XNOR U3965 ( .A(n3701), .B(n2136), .Z(n2794) );
  XOR U3966 ( .A(n3702), .B(n3232), .Z(out[354]) );
  IV U3967 ( .A(n3455), .Z(n3232) );
  XOR U3968 ( .A(n1947), .B(n3703), .Z(n3455) );
  ANDN U3969 ( .B(n2798), .A(n2799), .Z(n3702) );
  XNOR U3970 ( .A(n3704), .B(n2548), .Z(n2799) );
  XNOR U3971 ( .A(n3705), .B(n2142), .Z(n2798) );
  XOR U3972 ( .A(n3706), .B(n3235), .Z(out[353]) );
  XNOR U3973 ( .A(n3707), .B(n1953), .Z(n3235) );
  AND U3974 ( .A(n2808), .B(n3458), .Z(n3706) );
  XNOR U3975 ( .A(n3708), .B(n2146), .Z(n3458) );
  XOR U3976 ( .A(n3710), .B(n3238), .Z(out[352]) );
  XOR U3977 ( .A(n3711), .B(n1961), .Z(n3238) );
  AND U3978 ( .A(n2812), .B(n3461), .Z(n3710) );
  XNOR U3979 ( .A(n3712), .B(n2149), .Z(n3461) );
  XNOR U3980 ( .A(n3713), .B(n2562), .Z(n2812) );
  XOR U3981 ( .A(n3714), .B(n3245), .Z(out[351]) );
  XOR U3982 ( .A(n3715), .B(n1965), .Z(n3245) );
  ANDN U3983 ( .B(n2814), .A(n2816), .Z(n3714) );
  XNOR U3984 ( .A(n3716), .B(n2569), .Z(n2816) );
  XOR U3985 ( .A(n3717), .B(n2152), .Z(n2814) );
  XNOR U3986 ( .A(n3718), .B(n3249), .Z(out[350]) );
  XOR U3987 ( .A(n3719), .B(n1660), .Z(n3249) );
  ANDN U3988 ( .B(n2818), .A(n2820), .Z(n3718) );
  XNOR U3989 ( .A(n2575), .B(n3720), .Z(n2820) );
  XOR U3990 ( .A(n3721), .B(n2155), .Z(n2818) );
  XNOR U3991 ( .A(n3722), .B(n1083), .Z(out[34]) );
  XOR U3992 ( .A(n3724), .B(n3252), .Z(out[349]) );
  XOR U3993 ( .A(n3725), .B(n1664), .Z(n3252) );
  ANDN U3994 ( .B(n2822), .A(n2823), .Z(n3724) );
  XNOR U3995 ( .A(n2582), .B(n3726), .Z(n2823) );
  XOR U3996 ( .A(n3727), .B(n3728), .Z(n2822) );
  XOR U3997 ( .A(n3729), .B(n3255), .Z(out[348]) );
  XOR U3998 ( .A(n3730), .B(n1672), .Z(n3255) );
  AND U3999 ( .A(n2827), .B(n2826), .Z(n3729) );
  XOR U4000 ( .A(n3731), .B(n2163), .Z(n2826) );
  XNOR U4001 ( .A(n2589), .B(n3732), .Z(n2827) );
  XOR U4002 ( .A(n3733), .B(n3259), .Z(out[347]) );
  XNOR U4003 ( .A(n3734), .B(n3735), .Z(n3259) );
  AND U4004 ( .A(n2831), .B(n2830), .Z(n3733) );
  XOR U4005 ( .A(n3736), .B(n3737), .Z(n2830) );
  XOR U4006 ( .A(n3738), .B(n2601), .Z(n2831) );
  XNOR U4007 ( .A(n3739), .B(n3262), .Z(out[346]) );
  XNOR U4008 ( .A(n3740), .B(n1682), .Z(n3262) );
  AND U4009 ( .A(n2834), .B(n2836), .Z(n3739) );
  XOR U4010 ( .A(n3741), .B(n2608), .Z(n2836) );
  XNOR U4011 ( .A(n3742), .B(n3743), .Z(n2834) );
  XOR U4012 ( .A(n3744), .B(n3266), .Z(out[345]) );
  XOR U4013 ( .A(n3745), .B(n1686), .Z(n3266) );
  ANDN U4014 ( .B(n2839), .A(n2838), .Z(n3744) );
  XNOR U4015 ( .A(n3746), .B(n2172), .Z(n2838) );
  XNOR U4016 ( .A(n3747), .B(n2615), .Z(n2839) );
  XNOR U4017 ( .A(n3748), .B(n3270), .Z(out[344]) );
  XNOR U4018 ( .A(n3749), .B(n1690), .Z(n3270) );
  AND U4019 ( .A(n2844), .B(n2842), .Z(n3748) );
  XOR U4020 ( .A(n3750), .B(n3751), .Z(n2842) );
  XOR U4021 ( .A(n3752), .B(n2622), .Z(n2844) );
  XNOR U4022 ( .A(n3753), .B(n3273), .Z(out[343]) );
  XNOR U4023 ( .A(n3754), .B(n1694), .Z(n3273) );
  AND U4024 ( .A(n2854), .B(n2852), .Z(n3753) );
  IV U4025 ( .A(n3488), .Z(n2852) );
  XOR U4026 ( .A(n3755), .B(n3756), .Z(n3488) );
  XNOR U4027 ( .A(n3757), .B(n3758), .Z(n2854) );
  XOR U4028 ( .A(n3759), .B(n3276), .Z(out[342]) );
  XOR U4029 ( .A(n3760), .B(n1698), .Z(n3276) );
  AND U4030 ( .A(n2858), .B(n3491), .Z(n3759) );
  XOR U4031 ( .A(n3761), .B(n2185), .Z(n3491) );
  XNOR U4032 ( .A(n3762), .B(n3763), .Z(n2858) );
  XOR U4033 ( .A(n3764), .B(n3283), .Z(out[341]) );
  XNOR U4034 ( .A(n3765), .B(n1703), .Z(n3283) );
  ANDN U4035 ( .B(n2860), .A(n2862), .Z(n3764) );
  XOR U4036 ( .A(n3766), .B(n2643), .Z(n2862) );
  XNOR U4037 ( .A(n3767), .B(n2188), .Z(n2860) );
  XNOR U4038 ( .A(n3768), .B(n3286), .Z(out[340]) );
  XOR U4039 ( .A(n3769), .B(n1707), .Z(n3286) );
  AND U4040 ( .A(n2866), .B(n2864), .Z(n3768) );
  XOR U4041 ( .A(n3770), .B(n3771), .Z(n2864) );
  XNOR U4042 ( .A(n3772), .B(n3773), .Z(n2866) );
  XOR U4043 ( .A(n3774), .B(n1128), .Z(out[33]) );
  XOR U4044 ( .A(n3776), .B(n3289), .Z(out[339]) );
  XNOR U4045 ( .A(n3777), .B(n1711), .Z(n3289) );
  AND U4046 ( .A(n2868), .B(n2870), .Z(n3776) );
  XNOR U4047 ( .A(n3778), .B(n2657), .Z(n2870) );
  XNOR U4048 ( .A(n3779), .B(n2194), .Z(n2868) );
  XNOR U4049 ( .A(n3780), .B(n3292), .Z(out[338]) );
  XNOR U4050 ( .A(n3781), .B(n1720), .Z(n3292) );
  AND U4051 ( .A(n2874), .B(n2872), .Z(n3780) );
  XOR U4052 ( .A(n3782), .B(n3783), .Z(n2872) );
  XNOR U4053 ( .A(n3784), .B(n2664), .Z(n2874) );
  XOR U4054 ( .A(n3785), .B(n3295), .Z(out[337]) );
  XNOR U4055 ( .A(n3786), .B(n1725), .Z(n3295) );
  AND U4056 ( .A(n2878), .B(n3504), .Z(n3785) );
  XOR U4057 ( .A(n3787), .B(n3788), .Z(n3504) );
  XOR U4058 ( .A(n3789), .B(n2197), .Z(n2878) );
  XOR U4059 ( .A(n3790), .B(n3299), .Z(out[336]) );
  XOR U4060 ( .A(n3791), .B(n1729), .Z(n3299) );
  ANDN U4061 ( .B(n2880), .A(n2881), .Z(n3790) );
  XNOR U4062 ( .A(n3792), .B(n3793), .Z(n2881) );
  XNOR U4063 ( .A(n3794), .B(n1975), .Z(n2880) );
  XOR U4064 ( .A(n3795), .B(n3303), .Z(out[335]) );
  XNOR U4065 ( .A(n3796), .B(n1733), .Z(n3303) );
  ANDN U4066 ( .B(n2884), .A(n2886), .Z(n3795) );
  XOR U4067 ( .A(n3797), .B(n2211), .Z(n2886) );
  XNOR U4068 ( .A(n3798), .B(n1978), .Z(n2884) );
  XOR U4069 ( .A(n3799), .B(n3307), .Z(out[334]) );
  XOR U4070 ( .A(n3800), .B(n1738), .Z(n3307) );
  AND U4071 ( .A(n2890), .B(n3517), .Z(n3799) );
  XNOR U4072 ( .A(n3801), .B(n1981), .Z(n3517) );
  XNOR U4073 ( .A(n3802), .B(n3803), .Z(n2890) );
  XOR U4074 ( .A(n3804), .B(n3310), .Z(out[333]) );
  XOR U4075 ( .A(n3805), .B(n3806), .Z(n3310) );
  AND U4076 ( .A(n2898), .B(n2896), .Z(n3804) );
  IV U4077 ( .A(n3520), .Z(n2896) );
  XNOR U4078 ( .A(n3807), .B(n1984), .Z(n3520) );
  XNOR U4079 ( .A(n3808), .B(n3809), .Z(n2898) );
  XOR U4080 ( .A(n3810), .B(n3313), .Z(out[332]) );
  XNOR U4081 ( .A(n3811), .B(n1747), .Z(n3313) );
  AND U4082 ( .A(n2902), .B(n2900), .Z(n3810) );
  XOR U4083 ( .A(n3812), .B(n3813), .Z(n2900) );
  XNOR U4084 ( .A(n3814), .B(n3815), .Z(n2902) );
  XOR U4085 ( .A(n3816), .B(n3321), .Z(out[331]) );
  XNOR U4086 ( .A(n3817), .B(n3818), .Z(n3321) );
  AND U4087 ( .A(n2906), .B(n2904), .Z(n3816) );
  XOR U4088 ( .A(n3819), .B(n3820), .Z(n2904) );
  XNOR U4089 ( .A(n3821), .B(n3822), .Z(n2906) );
  XOR U4090 ( .A(n3823), .B(n3325), .Z(out[330]) );
  XOR U4091 ( .A(n3824), .B(n3825), .Z(n3325) );
  ANDN U4092 ( .B(n2908), .A(n2909), .Z(n3823) );
  XOR U4093 ( .A(n3827), .B(n1997), .Z(n2908) );
  XNOR U4094 ( .A(n3828), .B(n1171), .Z(out[32]) );
  ANDN U4095 ( .B(n1172), .A(n3829), .Z(n3828) );
  XOR U4096 ( .A(n3830), .B(n3328), .Z(out[329]) );
  XOR U4097 ( .A(n3831), .B(n1762), .Z(n3328) );
  ANDN U4098 ( .B(n2912), .A(n2913), .Z(n3830) );
  XOR U4099 ( .A(n3832), .B(n2259), .Z(n2913) );
  XNOR U4100 ( .A(n3833), .B(n2000), .Z(n2912) );
  XOR U4101 ( .A(n3834), .B(n3333), .Z(out[328]) );
  XOR U4102 ( .A(n3835), .B(n1770), .Z(n3333) );
  AND U4103 ( .A(n2918), .B(n2916), .Z(n3834) );
  XOR U4104 ( .A(n3836), .B(n3837), .Z(n2916) );
  XOR U4105 ( .A(n3838), .B(n3839), .Z(n2918) );
  XOR U4106 ( .A(n3840), .B(n3337), .Z(out[327]) );
  XNOR U4107 ( .A(n3841), .B(n3842), .Z(n3337) );
  AND U4108 ( .A(n2922), .B(n2920), .Z(n3840) );
  IV U4109 ( .A(n3533), .Z(n2920) );
  XNOR U4110 ( .A(n3843), .B(n2006), .Z(n3533) );
  XNOR U4111 ( .A(n3844), .B(n3845), .Z(n2922) );
  XOR U4112 ( .A(n3846), .B(n3341), .Z(out[326]) );
  XOR U4113 ( .A(n3847), .B(n1780), .Z(n3341) );
  AND U4114 ( .A(n2924), .B(n2926), .Z(n3846) );
  XNOR U4115 ( .A(n3848), .B(n3849), .Z(n2926) );
  XNOR U4116 ( .A(n3850), .B(n2009), .Z(n2924) );
  XOR U4117 ( .A(n3851), .B(n3345), .Z(out[325]) );
  XNOR U4118 ( .A(n3852), .B(n1784), .Z(n3345) );
  ANDN U4119 ( .B(n2928), .A(n2930), .Z(n3851) );
  XNOR U4120 ( .A(n3853), .B(n2287), .Z(n2930) );
  XNOR U4121 ( .A(n3854), .B(n2012), .Z(n2928) );
  XOR U4122 ( .A(n3855), .B(n3348), .Z(out[324]) );
  XOR U4123 ( .A(n3856), .B(n1788), .Z(n3348) );
  ANDN U4124 ( .B(n2934), .A(n2932), .Z(n3855) );
  XOR U4125 ( .A(n3857), .B(n2015), .Z(n2932) );
  XNOR U4126 ( .A(n3858), .B(n2294), .Z(n2934) );
  XOR U4127 ( .A(n3859), .B(n3352), .Z(out[323]) );
  XNOR U4128 ( .A(n3860), .B(n3861), .Z(n3352) );
  ANDN U4129 ( .B(n2940), .A(n2941), .Z(n3859) );
  XOR U4130 ( .A(n3862), .B(n2305), .Z(n2941) );
  XOR U4131 ( .A(n3863), .B(n2018), .Z(n2940) );
  XOR U4132 ( .A(n3864), .B(n3355), .Z(out[322]) );
  XOR U4133 ( .A(n3865), .B(n1797), .Z(n3355) );
  ANDN U4134 ( .B(n2944), .A(n2946), .Z(n3864) );
  XOR U4135 ( .A(n3866), .B(n2312), .Z(n2946) );
  XOR U4136 ( .A(n3867), .B(n2021), .Z(n2944) );
  XOR U4137 ( .A(n3868), .B(n3364), .Z(out[321]) );
  XOR U4138 ( .A(n3869), .B(n3870), .Z(n3364) );
  NOR U4139 ( .A(n2950), .B(n2948), .Z(n3868) );
  XOR U4140 ( .A(n3871), .B(n2024), .Z(n2948) );
  XNOR U4141 ( .A(n3872), .B(n2319), .Z(n2950) );
  XOR U4142 ( .A(n3873), .B(n3368), .Z(out[320]) );
  XNOR U4143 ( .A(n1804), .B(n3874), .Z(n3368) );
  ANDN U4144 ( .B(n2952), .A(n2953), .Z(n3873) );
  XNOR U4145 ( .A(n3875), .B(n2326), .Z(n2953) );
  XOR U4146 ( .A(n3876), .B(n2031), .Z(n2952) );
  XOR U4147 ( .A(n3877), .B(n1216), .Z(out[31]) );
  XNOR U4148 ( .A(n3879), .B(n2672), .Z(out[319]) );
  ANDN U4149 ( .B(n3880), .A(n2671), .Z(n3879) );
  XNOR U4150 ( .A(n3881), .B(n2716), .Z(out[318]) );
  ANDN U4151 ( .B(n3882), .A(n2715), .Z(n3881) );
  XNOR U4152 ( .A(n3883), .B(n2760), .Z(out[317]) );
  ANDN U4153 ( .B(n3884), .A(n2759), .Z(n3883) );
  XOR U4154 ( .A(n3885), .B(n2804), .Z(out[316]) );
  ANDN U4155 ( .B(n3886), .A(n2803), .Z(n3885) );
  XNOR U4156 ( .A(n3887), .B(n2849), .Z(out[315]) );
  ANDN U4157 ( .B(n2850), .A(n3888), .Z(n3887) );
  XNOR U4158 ( .A(n3889), .B(n2894), .Z(out[314]) );
  ANDN U4159 ( .B(n3890), .A(n2893), .Z(n3889) );
  XOR U4160 ( .A(n3891), .B(n2938), .Z(out[313]) );
  ANDN U4161 ( .B(n3892), .A(n2937), .Z(n3891) );
  XOR U4162 ( .A(n3893), .B(n2970), .Z(out[312]) );
  XNOR U4163 ( .A(n3895), .B(n2997), .Z(out[311]) );
  NOR U4164 ( .A(n3896), .B(n2996), .Z(n3895) );
  XOR U4165 ( .A(n3897), .B(n3024), .Z(out[310]) );
  ANDN U4166 ( .B(n3898), .A(n3023), .Z(n3897) );
  XNOR U4167 ( .A(n3899), .B(n1260), .Z(out[30]) );
  ANDN U4168 ( .B(n3900), .A(n1259), .Z(n3899) );
  XOR U4169 ( .A(n3901), .B(n3050), .Z(out[309]) );
  ANDN U4170 ( .B(n3902), .A(n3049), .Z(n3901) );
  XNOR U4171 ( .A(n3903), .B(n3075), .Z(out[308]) );
  XNOR U4172 ( .A(n3905), .B(n3100), .Z(out[307]) );
  AND U4173 ( .A(n3906), .B(n3907), .Z(n3905) );
  XNOR U4174 ( .A(n3908), .B(n3128), .Z(out[306]) );
  XOR U4175 ( .A(n3910), .B(n3171), .Z(out[305]) );
  XNOR U4176 ( .A(n3912), .B(n3205), .Z(out[304]) );
  ANDN U4177 ( .B(n3913), .A(n3204), .Z(n3912) );
  XNOR U4178 ( .A(n3914), .B(n3241), .Z(out[303]) );
  AND U4179 ( .A(n3242), .B(n3915), .Z(n3914) );
  XNOR U4180 ( .A(n3916), .B(n3279), .Z(out[302]) );
  XNOR U4181 ( .A(n3918), .B(n3318), .Z(out[301]) );
  XNOR U4182 ( .A(n3920), .B(n3359), .Z(out[300]) );
  AND U4183 ( .A(n3921), .B(n3360), .Z(n3920) );
  XOR U4184 ( .A(n3922), .B(n2450), .Z(out[2]) );
  ANDN U4185 ( .B(n3923), .A(n2449), .Z(n3922) );
  XOR U4186 ( .A(n3924), .B(n1305), .Z(out[29]) );
  ANDN U4187 ( .B(n1304), .A(n3925), .Z(n3924) );
  XOR U4188 ( .A(n3926), .B(n3390), .Z(out[299]) );
  ANDN U4189 ( .B(n3927), .A(n3389), .Z(n3926) );
  XNOR U4190 ( .A(n3928), .B(n3420), .Z(out[298]) );
  AND U4191 ( .A(n3421), .B(n3929), .Z(n3928) );
  XNOR U4192 ( .A(n3930), .B(n3449), .Z(out[297]) );
  AND U4193 ( .A(n3931), .B(n3932), .Z(n3930) );
  XOR U4194 ( .A(n3933), .B(n3479), .Z(out[296]) );
  XOR U4195 ( .A(n3935), .B(n3512), .Z(out[295]) );
  NOR U4196 ( .A(n3936), .B(n3511), .Z(n3935) );
  XOR U4197 ( .A(n3937), .B(n3539), .Z(out[294]) );
  NOR U4198 ( .A(n3938), .B(n3538), .Z(n3937) );
  XOR U4199 ( .A(n3939), .B(n3574), .Z(out[293]) );
  ANDN U4200 ( .B(n3940), .A(n3573), .Z(n3939) );
  XOR U4201 ( .A(n3941), .B(n3622), .Z(out[292]) );
  NOR U4202 ( .A(n3942), .B(n3621), .Z(n3941) );
  XOR U4203 ( .A(n3943), .B(n1039), .Z(out[291]) );
  XNOR U4204 ( .A(n3401), .B(n3944), .Z(n1039) );
  IV U4205 ( .A(n2350), .Z(n3401) );
  ANDN U4206 ( .B(n3945), .A(n3676), .Z(n3943) );
  XOR U4207 ( .A(n3946), .B(n1084), .Z(out[290]) );
  XOR U4208 ( .A(n3947), .B(n3948), .Z(n1084) );
  ANDN U4209 ( .B(n3949), .A(n3723), .Z(n3946) );
  XNOR U4210 ( .A(n3950), .B(n1349), .Z(out[28]) );
  ANDN U4211 ( .B(n3951), .A(n1348), .Z(n3950) );
  XOR U4212 ( .A(n3952), .B(n1127), .Z(out[289]) );
  XOR U4213 ( .A(n3407), .B(n3953), .Z(n1127) );
  ANDN U4214 ( .B(n3954), .A(n3775), .Z(n3952) );
  XNOR U4215 ( .A(n3955), .B(n1172), .Z(out[288]) );
  XNOR U4216 ( .A(n2369), .B(n3956), .Z(n1172) );
  AND U4217 ( .A(n3829), .B(n3957), .Z(n3955) );
  XOR U4218 ( .A(n3958), .B(n1215), .Z(out[287]) );
  XOR U4219 ( .A(n3412), .B(n3959), .Z(n1215) );
  ANDN U4220 ( .B(n3960), .A(n3878), .Z(n3958) );
  XOR U4221 ( .A(n3961), .B(n1259), .Z(out[286]) );
  XOR U4222 ( .A(n3962), .B(n2388), .Z(n1259) );
  NOR U4223 ( .A(n3963), .B(n3900), .Z(n3961) );
  XNOR U4224 ( .A(n3964), .B(n1304), .Z(out[285]) );
  XOR U4225 ( .A(n3965), .B(n2395), .Z(n1304) );
  XOR U4226 ( .A(n3967), .B(n1348), .Z(out[284]) );
  XNOR U4227 ( .A(n2403), .B(n3968), .Z(n1348) );
  AND U4228 ( .A(n3969), .B(n3970), .Z(n3967) );
  XOR U4229 ( .A(n3971), .B(n1392), .Z(out[283]) );
  AND U4230 ( .A(n3972), .B(n3973), .Z(n3971) );
  XNOR U4231 ( .A(n3974), .B(n1437), .Z(out[282]) );
  AND U4232 ( .A(n3975), .B(n3976), .Z(n3974) );
  XOR U4233 ( .A(n3977), .B(n1483), .Z(out[281]) );
  ANDN U4234 ( .B(n3978), .A(n3979), .Z(n3977) );
  XNOR U4235 ( .A(n3980), .B(n1518), .Z(out[280]) );
  AND U4236 ( .A(n3981), .B(n3982), .Z(n3980) );
  XNOR U4237 ( .A(n3983), .B(n1393), .Z(out[27]) );
  NOR U4238 ( .A(n1392), .B(n3972), .Z(n3983) );
  XOR U4239 ( .A(n2408), .B(n3984), .Z(n1392) );
  XNOR U4240 ( .A(n3985), .B(n1543), .Z(out[279]) );
  AND U4241 ( .A(n3986), .B(n3987), .Z(n3985) );
  XNOR U4242 ( .A(n3988), .B(n1567), .Z(out[278]) );
  AND U4243 ( .A(n3989), .B(n3990), .Z(n3988) );
  XOR U4244 ( .A(n3991), .B(n1590), .Z(out[277]) );
  ANDN U4245 ( .B(n3992), .A(n3993), .Z(n3991) );
  XNOR U4246 ( .A(n3994), .B(n1616), .Z(out[276]) );
  ANDN U4247 ( .B(n3995), .A(n3996), .Z(n3994) );
  XNOR U4248 ( .A(n3997), .B(n1640), .Z(out[275]) );
  ANDN U4249 ( .B(n3998), .A(n3999), .Z(n3997) );
  XNOR U4250 ( .A(n4000), .B(n1668), .Z(out[274]) );
  XNOR U4251 ( .A(n4003), .B(n1717), .Z(out[273]) );
  ANDN U4252 ( .B(n4004), .A(n4005), .Z(n4003) );
  XNOR U4253 ( .A(n4006), .B(n1767), .Z(out[272]) );
  AND U4254 ( .A(n4007), .B(n4008), .Z(n4006) );
  XNOR U4255 ( .A(n4009), .B(n1818), .Z(out[271]) );
  AND U4256 ( .A(n4010), .B(n4011), .Z(n4009) );
  XOR U4257 ( .A(n4012), .B(n1863), .Z(out[270]) );
  AND U4258 ( .A(n4013), .B(n4014), .Z(n4012) );
  XNOR U4259 ( .A(n4015), .B(n1436), .Z(out[26]) );
  ANDN U4260 ( .B(n1437), .A(n3975), .Z(n4015) );
  XNOR U4261 ( .A(n4016), .B(n4017), .Z(n1437) );
  XNOR U4262 ( .A(n4018), .B(n1909), .Z(out[269]) );
  XNOR U4263 ( .A(n4021), .B(n1958), .Z(out[268]) );
  ANDN U4264 ( .B(n4022), .A(n4023), .Z(n4021) );
  XNOR U4265 ( .A(n4024), .B(n1993), .Z(out[267]) );
  AND U4266 ( .A(n4025), .B(n4026), .Z(n4024) );
  XOR U4267 ( .A(n4027), .B(n2027), .Z(out[266]) );
  ANDN U4268 ( .B(n4028), .A(n4029), .Z(n4027) );
  XOR U4269 ( .A(n4030), .B(n1036), .Z(out[265]) );
  XOR U4270 ( .A(n4031), .B(n4032), .Z(n1036) );
  ANDN U4271 ( .B(n4033), .A(n1035), .Z(n4030) );
  XOR U4272 ( .A(n4034), .B(n1480), .Z(out[264]) );
  XOR U4273 ( .A(n4035), .B(n4036), .Z(n1480) );
  XOR U4274 ( .A(n4038), .B(n1814), .Z(out[263]) );
  XOR U4275 ( .A(n4039), .B(n3484), .Z(n1814) );
  AND U4276 ( .A(n1813), .B(n4040), .Z(n4038) );
  XOR U4277 ( .A(n4041), .B(n2175), .Z(out[262]) );
  XOR U4278 ( .A(n4042), .B(n3487), .Z(n2175) );
  XOR U4279 ( .A(n4044), .B(n2227), .Z(out[261]) );
  XOR U4280 ( .A(n4045), .B(n2573), .Z(n2227) );
  XOR U4281 ( .A(n4047), .B(n2301), .Z(out[260]) );
  XNOR U4282 ( .A(n4048), .B(n2578), .Z(n2301) );
  AND U4283 ( .A(n4049), .B(n4050), .Z(n4047) );
  XNOR U4284 ( .A(n4051), .B(n1484), .Z(out[25]) );
  ANDN U4285 ( .B(n3979), .A(n1483), .Z(n4051) );
  XOR U4286 ( .A(n2422), .B(n4052), .Z(n1483) );
  IV U4287 ( .A(n4053), .Z(n2422) );
  XOR U4288 ( .A(n4054), .B(n2375), .Z(out[259]) );
  XOR U4289 ( .A(n4055), .B(n3496), .Z(n2375) );
  AND U4290 ( .A(n4056), .B(n3508), .Z(n4054) );
  XOR U4291 ( .A(n4057), .B(n2449), .Z(out[258]) );
  XOR U4292 ( .A(n4058), .B(n2592), .Z(n2449) );
  ANDN U4293 ( .B(n4059), .A(n3923), .Z(n4057) );
  XOR U4294 ( .A(n4060), .B(n2523), .Z(out[257]) );
  AND U4295 ( .A(n4061), .B(n4062), .Z(n4060) );
  ANDN U4296 ( .B(n4064), .A(n4065), .Z(n4063) );
  XOR U4297 ( .A(n4066), .B(n2671), .Z(out[255]) );
  XNOR U4298 ( .A(n1804), .B(n4067), .Z(n2671) );
  ANDN U4299 ( .B(n4068), .A(n3880), .Z(n4066) );
  XOR U4300 ( .A(n4069), .B(n2715), .Z(out[254]) );
  XNOR U4301 ( .A(n1808), .B(n4070), .Z(n2715) );
  ANDN U4302 ( .B(n4071), .A(n3882), .Z(n4069) );
  XOR U4303 ( .A(n4072), .B(n2759), .Z(out[253]) );
  XOR U4304 ( .A(n1820), .B(n4073), .Z(n2759) );
  ANDN U4305 ( .B(n4074), .A(n3884), .Z(n4072) );
  XOR U4306 ( .A(n4075), .B(n2803), .Z(out[252]) );
  XOR U4307 ( .A(n1824), .B(n4076), .Z(n2803) );
  AND U4308 ( .A(n4077), .B(n4078), .Z(n4075) );
  XNOR U4309 ( .A(n4079), .B(n2850), .Z(out[251]) );
  XNOR U4310 ( .A(n1828), .B(n4080), .Z(n2850) );
  AND U4311 ( .A(n3888), .B(n4081), .Z(n4079) );
  XOR U4312 ( .A(n4082), .B(n2893), .Z(out[250]) );
  XOR U4313 ( .A(n1832), .B(n4083), .Z(n2893) );
  XOR U4314 ( .A(n4085), .B(n1517), .Z(out[24]) );
  ANDN U4315 ( .B(n1518), .A(n3981), .Z(n4085) );
  XOR U4316 ( .A(n2431), .B(n4086), .Z(n1518) );
  IV U4317 ( .A(n4087), .Z(n2431) );
  XOR U4318 ( .A(n4088), .B(n2937), .Z(out[249]) );
  XOR U4319 ( .A(n1837), .B(n4089), .Z(n2937) );
  XOR U4320 ( .A(n4091), .B(n2969), .Z(out[248]) );
  XOR U4321 ( .A(n1841), .B(n4092), .Z(n2969) );
  AND U4322 ( .A(n4093), .B(n3894), .Z(n4091) );
  XOR U4323 ( .A(n4094), .B(n2996), .Z(out[247]) );
  XOR U4324 ( .A(n1845), .B(n4095), .Z(n2996) );
  ANDN U4325 ( .B(n3896), .A(n4096), .Z(n4094) );
  XOR U4326 ( .A(n4097), .B(n3023), .Z(out[246]) );
  XNOR U4327 ( .A(n4098), .B(n4099), .Z(n3023) );
  ANDN U4328 ( .B(n4100), .A(n3898), .Z(n4097) );
  XOR U4329 ( .A(n4101), .B(n3049), .Z(out[245]) );
  XOR U4330 ( .A(n4102), .B(n4103), .Z(n3049) );
  ANDN U4331 ( .B(n4104), .A(n3902), .Z(n4101) );
  XOR U4332 ( .A(n4105), .B(n3076), .Z(out[244]) );
  XOR U4333 ( .A(n1858), .B(n4106), .Z(n3076) );
  NOR U4334 ( .A(n4107), .B(n3904), .Z(n4105) );
  XOR U4335 ( .A(n4108), .B(n3101), .Z(out[243]) );
  IV U4336 ( .A(n3907), .Z(n3101) );
  XOR U4337 ( .A(n1866), .B(n4109), .Z(n3907) );
  ANDN U4338 ( .B(n4110), .A(n3906), .Z(n4108) );
  XOR U4339 ( .A(n4111), .B(n3129), .Z(out[242]) );
  XOR U4340 ( .A(n1870), .B(n4112), .Z(n3129) );
  ANDN U4341 ( .B(n4113), .A(n3909), .Z(n4111) );
  XOR U4342 ( .A(n4114), .B(n3170), .Z(out[241]) );
  XOR U4343 ( .A(n4115), .B(n4116), .Z(n3170) );
  AND U4344 ( .A(n3911), .B(n4117), .Z(n4114) );
  XOR U4345 ( .A(n4118), .B(n3204), .Z(out[240]) );
  XOR U4346 ( .A(n1878), .B(n4119), .Z(n3204) );
  ANDN U4347 ( .B(n4120), .A(n3913), .Z(n4118) );
  XOR U4348 ( .A(n4121), .B(n1544), .Z(out[23]) );
  AND U4349 ( .A(n1543), .B(n4122), .Z(n4121) );
  XNOR U4350 ( .A(n2436), .B(n4123), .Z(n1543) );
  XNOR U4351 ( .A(n4124), .B(n3242), .Z(out[239]) );
  XNOR U4352 ( .A(n3628), .B(n4125), .Z(n3242) );
  ANDN U4353 ( .B(n4126), .A(n3915), .Z(n4124) );
  XNOR U4354 ( .A(n4127), .B(n3280), .Z(out[238]) );
  XNOR U4355 ( .A(n1888), .B(n4128), .Z(n3280) );
  AND U4356 ( .A(n4129), .B(n3917), .Z(n4127) );
  XOR U4357 ( .A(n4130), .B(n3317), .Z(out[237]) );
  XNOR U4358 ( .A(n1892), .B(n4131), .Z(n3317) );
  AND U4359 ( .A(n3919), .B(n4132), .Z(n4130) );
  XNOR U4360 ( .A(n4133), .B(n3360), .Z(out[236]) );
  XOR U4361 ( .A(n1896), .B(n4134), .Z(n3360) );
  ANDN U4362 ( .B(n4135), .A(n3921), .Z(n4133) );
  XOR U4363 ( .A(n4136), .B(n3389), .Z(out[235]) );
  XOR U4364 ( .A(n1900), .B(n4137), .Z(n3389) );
  AND U4365 ( .A(n4138), .B(n4139), .Z(n4136) );
  XNOR U4366 ( .A(n4140), .B(n3421), .Z(out[234]) );
  XNOR U4367 ( .A(n3656), .B(n4141), .Z(n3421) );
  NOR U4368 ( .A(n3929), .B(n4142), .Z(n4140) );
  IV U4369 ( .A(n4143), .Z(n3929) );
  XOR U4370 ( .A(n4144), .B(n3450), .Z(out[233]) );
  IV U4371 ( .A(n3932), .Z(n3450) );
  XOR U4372 ( .A(n1912), .B(n4145), .Z(n3932) );
  ANDN U4373 ( .B(n4146), .A(n3931), .Z(n4144) );
  XOR U4374 ( .A(n4147), .B(n3478), .Z(out[232]) );
  XOR U4375 ( .A(n1917), .B(n4148), .Z(n3478) );
  AND U4376 ( .A(n4149), .B(n3934), .Z(n4147) );
  XOR U4377 ( .A(n4150), .B(n3511), .Z(out[231]) );
  XOR U4378 ( .A(n1921), .B(n4151), .Z(n3511) );
  ANDN U4379 ( .B(n3936), .A(n4152), .Z(n4150) );
  XOR U4380 ( .A(n4153), .B(n3538), .Z(out[230]) );
  XNOR U4381 ( .A(n4154), .B(n4155), .Z(n3538) );
  AND U4382 ( .A(n3938), .B(n4156), .Z(n4153) );
  XOR U4383 ( .A(n4157), .B(n1566), .Z(out[22]) );
  AND U4384 ( .A(n1567), .B(n4158), .Z(n4157) );
  XOR U4385 ( .A(n2443), .B(n4159), .Z(n1567) );
  XOR U4386 ( .A(n4160), .B(n3573), .Z(out[229]) );
  XNOR U4387 ( .A(n1930), .B(n4161), .Z(n3573) );
  ANDN U4388 ( .B(n4162), .A(n3940), .Z(n4160) );
  XOR U4389 ( .A(n4163), .B(n3621), .Z(out[228]) );
  XNOR U4390 ( .A(n1934), .B(n4164), .Z(n3621) );
  ANDN U4391 ( .B(n3942), .A(n4165), .Z(n4163) );
  XOR U4392 ( .A(n4166), .B(n3676), .Z(out[227]) );
  XOR U4393 ( .A(n1939), .B(n4167), .Z(n3676) );
  NOR U4394 ( .A(n1038), .B(n3945), .Z(n4166) );
  XOR U4395 ( .A(n4168), .B(n3723), .Z(out[226]) );
  XNOR U4396 ( .A(n1943), .B(n4169), .Z(n3723) );
  ANDN U4397 ( .B(n4170), .A(n1082), .Z(n4168) );
  XOR U4398 ( .A(n4171), .B(n3775), .Z(out[225]) );
  XNOR U4399 ( .A(n1947), .B(n4172), .Z(n3775) );
  ANDN U4400 ( .B(n1126), .A(n3954), .Z(n4171) );
  XNOR U4401 ( .A(n4173), .B(n3829), .Z(out[224]) );
  XNOR U4402 ( .A(n4174), .B(n4175), .Z(n3829) );
  XOR U4403 ( .A(n4176), .B(n3878), .Z(out[223]) );
  XOR U4404 ( .A(n4177), .B(n1961), .Z(n3878) );
  ANDN U4405 ( .B(n4178), .A(n3960), .Z(n4176) );
  XOR U4406 ( .A(n4179), .B(n3900), .Z(out[222]) );
  XNOR U4407 ( .A(n4180), .B(n4181), .Z(n3900) );
  AND U4408 ( .A(n3963), .B(n1258), .Z(n4179) );
  IV U4409 ( .A(n4182), .Z(n1258) );
  XNOR U4410 ( .A(n4183), .B(n3925), .Z(out[221]) );
  XNOR U4411 ( .A(n4184), .B(n4185), .Z(n3925) );
  AND U4412 ( .A(n3966), .B(n4186), .Z(n4183) );
  XOR U4413 ( .A(n4187), .B(n3951), .Z(out[220]) );
  IV U4414 ( .A(n3970), .Z(n3951) );
  XOR U4415 ( .A(n4188), .B(n4189), .Z(n3970) );
  NOR U4416 ( .A(n3969), .B(n1347), .Z(n4187) );
  XNOR U4417 ( .A(n4190), .B(n1591), .Z(out[21]) );
  ANDN U4418 ( .B(n3993), .A(n1590), .Z(n4190) );
  XNOR U4419 ( .A(n4191), .B(n4192), .Z(n1590) );
  XNOR U4420 ( .A(n4193), .B(n3972), .Z(out[219]) );
  XNOR U4421 ( .A(n4194), .B(n1672), .Z(n3972) );
  NOR U4422 ( .A(n3973), .B(n1391), .Z(n4193) );
  XNOR U4423 ( .A(n4195), .B(n3975), .Z(out[218]) );
  XNOR U4424 ( .A(n4196), .B(n1677), .Z(n3975) );
  ANDN U4425 ( .B(n4197), .A(n1435), .Z(n4195) );
  XOR U4426 ( .A(n4198), .B(n3979), .Z(out[217]) );
  XOR U4427 ( .A(n4199), .B(n1682), .Z(n3979) );
  NOR U4428 ( .A(n3978), .B(n1482), .Z(n4198) );
  XNOR U4429 ( .A(n4200), .B(n3981), .Z(out[216]) );
  XNOR U4430 ( .A(n4201), .B(n1686), .Z(n3981) );
  IV U4431 ( .A(n4202), .Z(n1516) );
  XNOR U4432 ( .A(n4203), .B(n3987), .Z(out[215]) );
  IV U4433 ( .A(n4122), .Z(n3987) );
  XOR U4434 ( .A(n4204), .B(n1690), .Z(n4122) );
  ANDN U4435 ( .B(n1542), .A(n3986), .Z(n4203) );
  IV U4436 ( .A(n4205), .Z(n1542) );
  XNOR U4437 ( .A(n4206), .B(n3990), .Z(out[214]) );
  IV U4438 ( .A(n4158), .Z(n3990) );
  XOR U4439 ( .A(n4207), .B(n1694), .Z(n4158) );
  ANDN U4440 ( .B(n1565), .A(n3989), .Z(n4206) );
  IV U4441 ( .A(n4208), .Z(n1565) );
  XOR U4442 ( .A(n4209), .B(n3993), .Z(out[213]) );
  XOR U4443 ( .A(n4210), .B(n1698), .Z(n3993) );
  NOR U4444 ( .A(n3992), .B(n1589), .Z(n4209) );
  XNOR U4445 ( .A(n4211), .B(n3995), .Z(out[212]) );
  AND U4446 ( .A(n3996), .B(n4212), .Z(n4211) );
  XOR U4447 ( .A(n4213), .B(n3999), .Z(out[211]) );
  ANDN U4448 ( .B(n1638), .A(n3998), .Z(n4213) );
  XOR U4449 ( .A(n4214), .B(n4002), .Z(out[210]) );
  NOR U4450 ( .A(n4001), .B(n1667), .Z(n4214) );
  XOR U4451 ( .A(n4215), .B(n1615), .Z(out[20]) );
  ANDN U4452 ( .B(n1616), .A(n3995), .Z(n4215) );
  XOR U4453 ( .A(n4216), .B(n1703), .Z(n3995) );
  XNOR U4454 ( .A(n2461), .B(n4217), .Z(n1616) );
  XOR U4455 ( .A(n4218), .B(n4005), .Z(out[209]) );
  NOR U4456 ( .A(n4004), .B(n1715), .Z(n4218) );
  XNOR U4457 ( .A(n4219), .B(n4007), .Z(out[208]) );
  ANDN U4458 ( .B(n4220), .A(n1765), .Z(n4219) );
  XNOR U4459 ( .A(n4221), .B(n4010), .Z(out[207]) );
  AND U4460 ( .A(n1816), .B(n4222), .Z(n4221) );
  XNOR U4461 ( .A(n4223), .B(n4014), .Z(out[206]) );
  NOR U4462 ( .A(n1862), .B(n4013), .Z(n4223) );
  XOR U4463 ( .A(n4224), .B(n4020), .Z(out[205]) );
  XNOR U4464 ( .A(n4225), .B(n4022), .Z(out[204]) );
  AND U4465 ( .A(n4023), .B(n4226), .Z(n4225) );
  XNOR U4466 ( .A(n4227), .B(n4026), .Z(out[203]) );
  NOR U4467 ( .A(n1992), .B(n4025), .Z(n4227) );
  XNOR U4468 ( .A(n4228), .B(n4028), .Z(out[202]) );
  ANDN U4469 ( .B(n4029), .A(n2026), .Z(n4228) );
  XOR U4470 ( .A(n4229), .B(n1035), .Z(out[201]) );
  XNOR U4471 ( .A(n1756), .B(n4230), .Z(n1035) );
  ANDN U4472 ( .B(n4231), .A(n4033), .Z(n4229) );
  XOR U4473 ( .A(n4232), .B(n1479), .Z(out[200]) );
  XOR U4474 ( .A(n4233), .B(n1762), .Z(n1479) );
  NOR U4475 ( .A(n4037), .B(n2101), .Z(n4232) );
  XNOR U4476 ( .A(n4234), .B(n2524), .Z(out[1]) );
  ANDN U4477 ( .B(n4235), .A(n2523), .Z(n4234) );
  XOR U4478 ( .A(n4236), .B(n2605), .Z(n2523) );
  XOR U4479 ( .A(n4237), .B(n1639), .Z(out[19]) );
  AND U4480 ( .A(n3999), .B(n1640), .Z(n4237) );
  XOR U4481 ( .A(n2468), .B(n4238), .Z(n1640) );
  XNOR U4482 ( .A(n4239), .B(n1707), .Z(n3999) );
  XNOR U4483 ( .A(n4240), .B(n1813), .Z(out[199]) );
  XNOR U4484 ( .A(n4241), .B(n1770), .Z(n1813) );
  ANDN U4485 ( .B(n4242), .A(n2138), .Z(n4240) );
  XOR U4486 ( .A(n4243), .B(n2224), .Z(out[198]) );
  XOR U4487 ( .A(n4244), .B(n1775), .Z(n2224) );
  XOR U4488 ( .A(n4245), .B(n2846), .Z(out[197]) );
  XOR U4489 ( .A(n4246), .B(n1780), .Z(n2846) );
  NOR U4490 ( .A(n4046), .B(n2226), .Z(n4245) );
  XOR U4491 ( .A(n4247), .B(n3167), .Z(out[196]) );
  IV U4492 ( .A(n4050), .Z(n3167) );
  XOR U4493 ( .A(n4248), .B(n1784), .Z(n4050) );
  IV U4494 ( .A(n4249), .Z(n1784) );
  IV U4495 ( .A(n4250), .Z(n2300) );
  XNOR U4496 ( .A(n4251), .B(n3508), .Z(out[195]) );
  XOR U4497 ( .A(n4252), .B(n1788), .Z(n3508) );
  NOR U4498 ( .A(n2374), .B(n4056), .Z(n4251) );
  XOR U4499 ( .A(n4253), .B(n3923), .Z(out[194]) );
  XNOR U4500 ( .A(n3860), .B(n4254), .Z(n3923) );
  NOR U4501 ( .A(n4059), .B(n2448), .Z(n4253) );
  XNOR U4502 ( .A(n4255), .B(n4062), .Z(out[193]) );
  IV U4503 ( .A(n4235), .Z(n4062) );
  XOR U4504 ( .A(n4256), .B(n1797), .Z(n4235) );
  NOR U4505 ( .A(n4061), .B(n2522), .Z(n4255) );
  XOR U4506 ( .A(n4257), .B(n4065), .Z(out[192]) );
  NOR U4507 ( .A(n4064), .B(n2596), .Z(n4257) );
  XOR U4508 ( .A(n4258), .B(n3880), .Z(out[191]) );
  XOR U4509 ( .A(n4259), .B(n2079), .Z(n3880) );
  XOR U4510 ( .A(n4260), .B(n3882), .Z(out[190]) );
  XNOR U4511 ( .A(n4261), .B(n2082), .Z(n3882) );
  NOR U4512 ( .A(n4071), .B(n2714), .Z(n4260) );
  XOR U4513 ( .A(n4262), .B(n1669), .Z(out[18]) );
  AND U4514 ( .A(n1668), .B(n4002), .Z(n4262) );
  XNOR U4515 ( .A(n4263), .B(n1711), .Z(n4002) );
  XOR U4516 ( .A(n4265), .B(n3884), .Z(out[189]) );
  XOR U4517 ( .A(n4266), .B(n2085), .Z(n3884) );
  XOR U4518 ( .A(n4267), .B(n3886), .Z(out[188]) );
  IV U4519 ( .A(n4078), .Z(n3886) );
  XNOR U4520 ( .A(n4268), .B(n2088), .Z(n4078) );
  ANDN U4521 ( .B(n2802), .A(n4077), .Z(n4267) );
  IV U4522 ( .A(n4269), .Z(n2802) );
  XNOR U4523 ( .A(n4270), .B(n3888), .Z(out[187]) );
  XOR U4524 ( .A(n4271), .B(n2092), .Z(n3888) );
  NOR U4525 ( .A(n2848), .B(n4081), .Z(n4270) );
  XOR U4526 ( .A(n4272), .B(n3890), .Z(out[186]) );
  XOR U4527 ( .A(n2094), .B(n4273), .Z(n3890) );
  ANDN U4528 ( .B(n2892), .A(n4084), .Z(n4272) );
  XOR U4529 ( .A(n4274), .B(n3892), .Z(out[185]) );
  XOR U4530 ( .A(n3646), .B(n4275), .Z(n3892) );
  ANDN U4531 ( .B(n2936), .A(n4090), .Z(n4274) );
  IV U4532 ( .A(n4276), .Z(n2936) );
  XNOR U4533 ( .A(n4277), .B(n3894), .Z(out[184]) );
  XNOR U4534 ( .A(n4278), .B(n2105), .Z(n3894) );
  NOR U4535 ( .A(n2968), .B(n4093), .Z(n4277) );
  XNOR U4536 ( .A(n4279), .B(n3896), .Z(out[183]) );
  XNOR U4537 ( .A(n2107), .B(n4280), .Z(n3896) );
  ANDN U4538 ( .B(n4096), .A(n2995), .Z(n4279) );
  XOR U4539 ( .A(n4281), .B(n3898), .Z(out[182]) );
  XOR U4540 ( .A(n3664), .B(n4282), .Z(n3898) );
  XOR U4541 ( .A(n4283), .B(n3902), .Z(out[181]) );
  XNOR U4542 ( .A(n4284), .B(n4285), .Z(n3902) );
  NOR U4543 ( .A(n3048), .B(n4104), .Z(n4283) );
  XOR U4544 ( .A(n4286), .B(n3904), .Z(out[180]) );
  XNOR U4545 ( .A(n3672), .B(n4287), .Z(n3904) );
  ANDN U4546 ( .B(n4107), .A(n3074), .Z(n4286) );
  XNOR U4547 ( .A(n4288), .B(n1716), .Z(out[17]) );
  AND U4548 ( .A(n4005), .B(n1717), .Z(n4288) );
  XOR U4549 ( .A(n4289), .B(n4290), .Z(n1717) );
  XOR U4550 ( .A(n4291), .B(n1720), .Z(n4005) );
  XOR U4551 ( .A(n4292), .B(n3906), .Z(out[179]) );
  XNOR U4552 ( .A(n3679), .B(n4293), .Z(n3906) );
  NOR U4553 ( .A(n4110), .B(n3099), .Z(n4292) );
  XOR U4554 ( .A(n4294), .B(n3909), .Z(out[178]) );
  XOR U4555 ( .A(n2126), .B(n4295), .Z(n3909) );
  NOR U4556 ( .A(n3127), .B(n4113), .Z(n4294) );
  XNOR U4557 ( .A(n4296), .B(n3911), .Z(out[177]) );
  XNOR U4558 ( .A(n4297), .B(n2130), .Z(n3911) );
  XOR U4559 ( .A(n4298), .B(n3913), .Z(out[176]) );
  XOR U4560 ( .A(n4299), .B(n2133), .Z(n3913) );
  NOR U4561 ( .A(n3203), .B(n4120), .Z(n4298) );
  XOR U4562 ( .A(n4300), .B(n3915), .Z(out[175]) );
  XOR U4563 ( .A(n4301), .B(n2136), .Z(n3915) );
  ANDN U4564 ( .B(n4302), .A(n3240), .Z(n4300) );
  XNOR U4565 ( .A(n4303), .B(n3917), .Z(out[174]) );
  XNOR U4566 ( .A(n4304), .B(n2142), .Z(n3917) );
  NOR U4567 ( .A(n4129), .B(n3278), .Z(n4303) );
  XNOR U4568 ( .A(n4305), .B(n3919), .Z(out[173]) );
  XNOR U4569 ( .A(n4306), .B(n2146), .Z(n3919) );
  ANDN U4570 ( .B(n4307), .A(n3316), .Z(n4305) );
  XOR U4571 ( .A(n4308), .B(n3921), .Z(out[172]) );
  XOR U4572 ( .A(n4309), .B(n2149), .Z(n3921) );
  NOR U4573 ( .A(n3358), .B(n4135), .Z(n4308) );
  XOR U4574 ( .A(n4310), .B(n3927), .Z(out[171]) );
  IV U4575 ( .A(n4139), .Z(n3927) );
  XOR U4576 ( .A(n4311), .B(n2152), .Z(n4139) );
  ANDN U4577 ( .B(n3388), .A(n4138), .Z(n4310) );
  IV U4578 ( .A(n4312), .Z(n3388) );
  XNOR U4579 ( .A(n4313), .B(n4143), .Z(out[170]) );
  XOR U4580 ( .A(n4314), .B(n2155), .Z(n4143) );
  AND U4581 ( .A(n4142), .B(n3419), .Z(n4313) );
  XNOR U4582 ( .A(n4315), .B(n1766), .Z(out[16]) );
  ANDN U4583 ( .B(n1767), .A(n4007), .Z(n4315) );
  XOR U4584 ( .A(n4316), .B(n1725), .Z(n4007) );
  XNOR U4585 ( .A(n4317), .B(n2492), .Z(n1767) );
  XOR U4586 ( .A(n4318), .B(n3931), .Z(out[169]) );
  XOR U4587 ( .A(n4319), .B(n2159), .Z(n3931) );
  ANDN U4588 ( .B(n4320), .A(n3448), .Z(n4318) );
  XNOR U4589 ( .A(n4321), .B(n3934), .Z(out[168]) );
  XOR U4590 ( .A(n4322), .B(n2163), .Z(n3934) );
  NOR U4591 ( .A(n3477), .B(n4149), .Z(n4321) );
  XNOR U4592 ( .A(n4323), .B(n3936), .Z(out[167]) );
  XNOR U4593 ( .A(n4324), .B(n2166), .Z(n3936) );
  AND U4594 ( .A(n4152), .B(n3510), .Z(n4323) );
  XNOR U4595 ( .A(n4325), .B(n3938), .Z(out[166]) );
  XNOR U4596 ( .A(n4326), .B(n2169), .Z(n3938) );
  ANDN U4597 ( .B(n3537), .A(n4156), .Z(n4325) );
  IV U4598 ( .A(n4327), .Z(n3537) );
  XOR U4599 ( .A(n4328), .B(n3940), .Z(out[165]) );
  XNOR U4600 ( .A(n4329), .B(n2172), .Z(n3940) );
  ANDN U4601 ( .B(n3572), .A(n4162), .Z(n4328) );
  XNOR U4602 ( .A(n4330), .B(n3942), .Z(out[164]) );
  XNOR U4603 ( .A(n4331), .B(n2179), .Z(n3942) );
  AND U4604 ( .A(n4165), .B(n3620), .Z(n4330) );
  XOR U4605 ( .A(n4332), .B(n3945), .Z(out[163]) );
  XNOR U4606 ( .A(n4333), .B(n2182), .Z(n3945) );
  AND U4607 ( .A(n1040), .B(n1038), .Z(n4332) );
  XNOR U4608 ( .A(n2575), .B(n4334), .Z(n1038) );
  XNOR U4609 ( .A(n2415), .B(n4335), .Z(n1040) );
  IV U4610 ( .A(n4336), .Z(n2415) );
  XOR U4611 ( .A(n4337), .B(n3949), .Z(out[162]) );
  IV U4612 ( .A(n4170), .Z(n3949) );
  XOR U4613 ( .A(n4338), .B(n2185), .Z(n4170) );
  ANDN U4614 ( .B(n1082), .A(n1083), .Z(n4337) );
  XNOR U4615 ( .A(n2424), .B(n4339), .Z(n1083) );
  XNOR U4616 ( .A(n2582), .B(n4340), .Z(n1082) );
  XOR U4617 ( .A(n4341), .B(n3954), .Z(out[161]) );
  XOR U4618 ( .A(n4342), .B(n2188), .Z(n3954) );
  ANDN U4619 ( .B(n1128), .A(n1126), .Z(n4341) );
  XNOR U4620 ( .A(n4343), .B(n4344), .Z(n1126) );
  XOR U4621 ( .A(n4345), .B(n4346), .Z(n1128) );
  XOR U4622 ( .A(n4347), .B(n3957), .Z(out[160]) );
  XOR U4623 ( .A(n4348), .B(n2191), .Z(n3957) );
  ANDN U4624 ( .B(n1170), .A(n1171), .Z(n4347) );
  XNOR U4625 ( .A(n4349), .B(n3211), .Z(n1171) );
  XNOR U4626 ( .A(n4350), .B(n2601), .Z(n1170) );
  XOR U4627 ( .A(n4351), .B(n1817), .Z(out[15]) );
  ANDN U4628 ( .B(n1818), .A(n4010), .Z(n4351) );
  XNOR U4629 ( .A(n4352), .B(n1729), .Z(n4010) );
  XNOR U4630 ( .A(n2496), .B(n4353), .Z(n1818) );
  IV U4631 ( .A(n4354), .Z(n2496) );
  XOR U4632 ( .A(n4355), .B(n3960), .Z(out[159]) );
  XNOR U4633 ( .A(n4356), .B(n4357), .Z(n3960) );
  AND U4634 ( .A(n1216), .B(n1214), .Z(n4355) );
  IV U4635 ( .A(n4178), .Z(n1214) );
  XOR U4636 ( .A(n4358), .B(n2608), .Z(n4178) );
  XNOR U4637 ( .A(n4359), .B(n2446), .Z(n1216) );
  XOR U4638 ( .A(n4360), .B(n4361), .Z(out[1599]) );
  XOR U4639 ( .A(n4362), .B(n4363), .Z(n4361) );
  AND U4640 ( .A(n4364), .B(n4365), .Z(n4363) );
  XNOR U4641 ( .A(n4368), .B(n4369), .Z(out[1598]) );
  XNOR U4642 ( .A(n4372), .B(n4373), .Z(out[1597]) );
  ANDN U4643 ( .B(n4374), .A(n4375), .Z(n4372) );
  XOR U4644 ( .A(n4376), .B(n4377), .Z(out[1596]) );
  AND U4645 ( .A(n4378), .B(n4379), .Z(n4376) );
  XNOR U4646 ( .A(n4380), .B(n4381), .Z(out[1595]) );
  AND U4647 ( .A(n4382), .B(n4383), .Z(n4380) );
  XOR U4648 ( .A(n4384), .B(n4385), .Z(out[1594]) );
  ANDN U4649 ( .B(n4386), .A(n4387), .Z(n4384) );
  XOR U4650 ( .A(n4388), .B(n4389), .Z(out[1593]) );
  XNOR U4651 ( .A(n4392), .B(n4393), .Z(out[1592]) );
  AND U4652 ( .A(n4394), .B(n4395), .Z(n4392) );
  XNOR U4653 ( .A(n4396), .B(n4397), .Z(out[1591]) );
  AND U4654 ( .A(n4398), .B(n4399), .Z(n4396) );
  XNOR U4655 ( .A(n4400), .B(n4401), .Z(out[1590]) );
  AND U4656 ( .A(n4402), .B(n4403), .Z(n4400) );
  XNOR U4657 ( .A(n4404), .B(n3963), .Z(out[158]) );
  XNOR U4658 ( .A(n4405), .B(n3783), .Z(n3963) );
  ANDN U4659 ( .B(n4182), .A(n1260), .Z(n4404) );
  XOR U4660 ( .A(n4406), .B(n2455), .Z(n1260) );
  XNOR U4661 ( .A(n4407), .B(n2615), .Z(n4182) );
  XNOR U4662 ( .A(n4408), .B(n4409), .Z(out[1589]) );
  ANDN U4663 ( .B(n4410), .A(n4411), .Z(n4408) );
  XOR U4664 ( .A(n4412), .B(n4413), .Z(out[1588]) );
  ANDN U4665 ( .B(n4414), .A(n4415), .Z(n4412) );
  XOR U4666 ( .A(n4416), .B(n4417), .Z(out[1587]) );
  AND U4667 ( .A(n4418), .B(n4419), .Z(n4416) );
  XNOR U4668 ( .A(n4420), .B(n4421), .Z(out[1586]) );
  AND U4669 ( .A(n4422), .B(n4423), .Z(n4420) );
  XOR U4670 ( .A(n4424), .B(n4425), .Z(out[1585]) );
  ANDN U4671 ( .B(n4426), .A(n4427), .Z(n4424) );
  XOR U4672 ( .A(n4428), .B(n4429), .Z(out[1584]) );
  ANDN U4673 ( .B(n4430), .A(n4431), .Z(n4428) );
  XOR U4674 ( .A(n4432), .B(n4433), .Z(out[1583]) );
  AND U4675 ( .A(n4434), .B(n4435), .Z(n4432) );
  XOR U4676 ( .A(n4436), .B(n4437), .Z(out[1582]) );
  AND U4677 ( .A(n4438), .B(n4439), .Z(n4436) );
  XOR U4678 ( .A(n4440), .B(n4441), .Z(out[1581]) );
  AND U4679 ( .A(n4442), .B(n4443), .Z(n4440) );
  XOR U4680 ( .A(n4444), .B(n4445), .Z(out[1580]) );
  AND U4681 ( .A(n4446), .B(n4447), .Z(n4444) );
  XNOR U4682 ( .A(n4448), .B(n3966), .Z(out[157]) );
  XOR U4683 ( .A(n4449), .B(n3788), .Z(n3966) );
  AND U4684 ( .A(n1305), .B(n1303), .Z(n4448) );
  IV U4685 ( .A(n4186), .Z(n1303) );
  XOR U4686 ( .A(n4450), .B(n2622), .Z(n4186) );
  XOR U4687 ( .A(n4451), .B(n2464), .Z(n1305) );
  XNOR U4688 ( .A(n4452), .B(n4453), .Z(out[1579]) );
  AND U4689 ( .A(n4454), .B(n4455), .Z(n4452) );
  XNOR U4690 ( .A(n4456), .B(n4457), .Z(out[1578]) );
  AND U4691 ( .A(n4458), .B(n4459), .Z(n4456) );
  XOR U4692 ( .A(n4460), .B(n4461), .Z(out[1577]) );
  XNOR U4693 ( .A(n4464), .B(n4465), .Z(out[1576]) );
  AND U4694 ( .A(n4466), .B(n4467), .Z(n4464) );
  XOR U4695 ( .A(n4468), .B(n4469), .Z(out[1575]) );
  XOR U4696 ( .A(n4472), .B(n4473), .Z(out[1574]) );
  XOR U4697 ( .A(n4476), .B(n4477), .Z(out[1573]) );
  NOR U4698 ( .A(n4478), .B(n4479), .Z(n4476) );
  XNOR U4699 ( .A(n4480), .B(n4481), .Z(out[1572]) );
  AND U4700 ( .A(n4482), .B(n4483), .Z(n4480) );
  XOR U4701 ( .A(n4484), .B(n4485), .Z(out[1571]) );
  AND U4702 ( .A(n4486), .B(n4487), .Z(n4484) );
  XOR U4703 ( .A(n4488), .B(n4489), .Z(out[1570]) );
  AND U4704 ( .A(n4490), .B(n4491), .Z(n4488) );
  XOR U4705 ( .A(n4492), .B(n3969), .Z(out[156]) );
  XNOR U4706 ( .A(n4493), .B(n4494), .Z(n3969) );
  ANDN U4707 ( .B(n1347), .A(n1349), .Z(n4492) );
  XNOR U4708 ( .A(n4495), .B(n2471), .Z(n1349) );
  XNOR U4709 ( .A(n4496), .B(n3758), .Z(n1347) );
  XNOR U4710 ( .A(n4497), .B(n4498), .Z(out[1569]) );
  ANDN U4711 ( .B(n4499), .A(n4500), .Z(n4497) );
  XNOR U4712 ( .A(n4501), .B(n4502), .Z(out[1568]) );
  AND U4713 ( .A(n4503), .B(n4504), .Z(n4501) );
  XNOR U4714 ( .A(n4505), .B(n4506), .Z(out[1567]) );
  XOR U4715 ( .A(n4507), .B(n4508), .Z(n4506) );
  AND U4716 ( .A(n4509), .B(n4510), .Z(n4508) );
  XNOR U4717 ( .A(n4513), .B(n4514), .Z(out[1566]) );
  AND U4718 ( .A(n4515), .B(n4516), .Z(n4513) );
  XNOR U4719 ( .A(n4517), .B(n4518), .Z(out[1565]) );
  AND U4720 ( .A(n4519), .B(n4520), .Z(n4517) );
  XNOR U4721 ( .A(n4521), .B(n4522), .Z(out[1564]) );
  ANDN U4722 ( .B(n4523), .A(n4524), .Z(n4521) );
  XOR U4723 ( .A(n4525), .B(n4526), .Z(out[1563]) );
  AND U4724 ( .A(n4527), .B(n4528), .Z(n4525) );
  XOR U4725 ( .A(n4529), .B(n4530), .Z(out[1562]) );
  ANDN U4726 ( .B(n4531), .A(n4532), .Z(n4529) );
  XOR U4727 ( .A(n4533), .B(n4534), .Z(out[1561]) );
  AND U4728 ( .A(n4535), .B(n4536), .Z(n4533) );
  XOR U4729 ( .A(n4537), .B(n4538), .Z(out[1560]) );
  AND U4730 ( .A(n4539), .B(n4540), .Z(n4537) );
  XOR U4731 ( .A(n4541), .B(n3973), .Z(out[155]) );
  XOR U4732 ( .A(n4542), .B(n1978), .Z(n3973) );
  ANDN U4733 ( .B(n1391), .A(n1393), .Z(n4541) );
  XOR U4734 ( .A(n4543), .B(n2476), .Z(n1393) );
  XOR U4735 ( .A(n4544), .B(n3763), .Z(n1391) );
  IV U4736 ( .A(n2636), .Z(n3763) );
  XOR U4737 ( .A(n4545), .B(n4546), .Z(out[1559]) );
  XOR U4738 ( .A(n4549), .B(n4550), .Z(out[1558]) );
  XNOR U4739 ( .A(n4553), .B(n4554), .Z(out[1557]) );
  XNOR U4740 ( .A(n4557), .B(n4558), .Z(out[1556]) );
  AND U4741 ( .A(n4559), .B(n4560), .Z(n4557) );
  XNOR U4742 ( .A(n4561), .B(n4562), .Z(out[1555]) );
  AND U4743 ( .A(n4563), .B(n4564), .Z(n4561) );
  XNOR U4744 ( .A(n4565), .B(n4566), .Z(out[1554]) );
  XNOR U4745 ( .A(n4569), .B(n4570), .Z(out[1553]) );
  AND U4746 ( .A(n4571), .B(n4572), .Z(n4569) );
  XNOR U4747 ( .A(n4573), .B(n4574), .Z(out[1552]) );
  AND U4748 ( .A(n4575), .B(n4576), .Z(n4573) );
  XOR U4749 ( .A(n4578), .B(n4579), .Z(n4577) );
  XNOR U4750 ( .A(n4583), .B(n4584), .Z(out[1550]) );
  XOR U4751 ( .A(n4587), .B(n3976), .Z(out[154]) );
  IV U4752 ( .A(n4197), .Z(n3976) );
  XNOR U4753 ( .A(n4588), .B(n1981), .Z(n4197) );
  ANDN U4754 ( .B(n1435), .A(n1436), .Z(n4587) );
  XNOR U4755 ( .A(n4589), .B(n2483), .Z(n1436) );
  XNOR U4756 ( .A(n4590), .B(n4591), .Z(n1435) );
  XNOR U4757 ( .A(n4592), .B(n4593), .Z(out[1549]) );
  ANDN U4758 ( .B(n4594), .A(n4595), .Z(n4592) );
  XOR U4759 ( .A(n4596), .B(n4597), .Z(out[1548]) );
  XNOR U4760 ( .A(n4600), .B(n4601), .Z(out[1547]) );
  XOR U4761 ( .A(n4604), .B(n4605), .Z(out[1546]) );
  ANDN U4762 ( .B(n4606), .A(n4607), .Z(n4604) );
  XOR U4763 ( .A(n4608), .B(n4609), .Z(out[1545]) );
  AND U4764 ( .A(n4610), .B(n4611), .Z(n4608) );
  XNOR U4765 ( .A(n4612), .B(n4613), .Z(out[1544]) );
  AND U4766 ( .A(n4614), .B(n4615), .Z(n4612) );
  XOR U4767 ( .A(n4616), .B(n4617), .Z(out[1543]) );
  AND U4768 ( .A(n4618), .B(n4619), .Z(n4616) );
  XOR U4769 ( .A(n4620), .B(n4621), .Z(out[1542]) );
  XNOR U4770 ( .A(n4624), .B(n4625), .Z(out[1541]) );
  ANDN U4771 ( .B(n4626), .A(n4627), .Z(n4624) );
  XOR U4772 ( .A(n4628), .B(n4629), .Z(out[1540]) );
  XOR U4773 ( .A(n4632), .B(n3978), .Z(out[153]) );
  XOR U4774 ( .A(n4633), .B(n1984), .Z(n3978) );
  ANDN U4775 ( .B(n1482), .A(n1484), .Z(n4632) );
  XNOR U4776 ( .A(n4634), .B(n2490), .Z(n1484) );
  XOR U4777 ( .A(n4635), .B(n3773), .Z(n1482) );
  XOR U4778 ( .A(n4636), .B(n4637), .Z(out[1539]) );
  XOR U4779 ( .A(n4638), .B(n4639), .Z(n4637) );
  NAND U4780 ( .A(n4640), .B(n4510), .Z(n4639) );
  AND U4781 ( .A(n4641), .B(n4642), .Z(n4638) );
  XOR U4782 ( .A(n4643), .B(n4644), .Z(out[1538]) );
  AND U4783 ( .A(n4645), .B(n4646), .Z(n4643) );
  XOR U4784 ( .A(n4647), .B(n4648), .Z(out[1537]) );
  XOR U4785 ( .A(n4649), .B(n4650), .Z(n4648) );
  ANDN U4786 ( .B(n4651), .A(n4652), .Z(n4649) );
  XOR U4787 ( .A(n4653), .B(n4654), .Z(out[1536]) );
  XOR U4788 ( .A(n4655), .B(n4656), .Z(n4654) );
  AND U4789 ( .A(n4657), .B(n4658), .Z(n4655) );
  XOR U4790 ( .A(n4659), .B(n4367), .Z(out[1535]) );
  ANDN U4791 ( .B(n4660), .A(n4366), .Z(n4659) );
  XOR U4792 ( .A(n4661), .B(n4371), .Z(out[1534]) );
  ANDN U4793 ( .B(n4662), .A(n4370), .Z(n4661) );
  XOR U4794 ( .A(n4663), .B(n4375), .Z(out[1533]) );
  ANDN U4795 ( .B(n4664), .A(n4374), .Z(n4663) );
  XNOR U4796 ( .A(n4665), .B(n4379), .Z(out[1532]) );
  ANDN U4797 ( .B(n4666), .A(n4378), .Z(n4665) );
  XNOR U4798 ( .A(n4667), .B(n4382), .Z(out[1531]) );
  AND U4799 ( .A(n4668), .B(n4669), .Z(n4667) );
  XNOR U4800 ( .A(n4670), .B(n4386), .Z(out[1530]) );
  AND U4801 ( .A(n4387), .B(n4671), .Z(n4670) );
  XOR U4802 ( .A(n4672), .B(n3982), .Z(out[152]) );
  XOR U4803 ( .A(n4673), .B(n1987), .Z(n3982) );
  AND U4804 ( .A(n1517), .B(n4202), .Z(n4672) );
  XOR U4805 ( .A(n4674), .B(n2657), .Z(n4202) );
  XNOR U4806 ( .A(n4675), .B(n4676), .Z(n1517) );
  XNOR U4807 ( .A(n4677), .B(n4390), .Z(out[1529]) );
  AND U4808 ( .A(n4678), .B(n4391), .Z(n4677) );
  XNOR U4809 ( .A(n4679), .B(n4395), .Z(out[1528]) );
  NOR U4810 ( .A(n4680), .B(n4394), .Z(n4679) );
  XNOR U4811 ( .A(n4681), .B(n4398), .Z(out[1527]) );
  XNOR U4812 ( .A(n4683), .B(n4403), .Z(out[1526]) );
  ANDN U4813 ( .B(n4684), .A(n4402), .Z(n4683) );
  XOR U4814 ( .A(n4685), .B(n4411), .Z(out[1525]) );
  XOR U4815 ( .A(n4687), .B(n4415), .Z(out[1524]) );
  XNOR U4816 ( .A(n4689), .B(n4418), .Z(out[1523]) );
  XNOR U4817 ( .A(n4691), .B(n4423), .Z(out[1522]) );
  ANDN U4818 ( .B(n4692), .A(n4422), .Z(n4691) );
  XOR U4819 ( .A(n4693), .B(n4427), .Z(out[1521]) );
  ANDN U4820 ( .B(n4694), .A(n4426), .Z(n4693) );
  XOR U4821 ( .A(n4695), .B(n4431), .Z(out[1520]) );
  XOR U4822 ( .A(n4697), .B(n3986), .Z(out[151]) );
  XOR U4823 ( .A(n4698), .B(n1990), .Z(n3986) );
  IV U4824 ( .A(n3820), .Z(n1990) );
  AND U4825 ( .A(n1544), .B(n4205), .Z(n4697) );
  XOR U4826 ( .A(n4699), .B(n2664), .Z(n4205) );
  XOR U4827 ( .A(n4700), .B(n4701), .Z(n1544) );
  XNOR U4828 ( .A(n4702), .B(n4435), .Z(out[1519]) );
  ANDN U4829 ( .B(n4703), .A(n4434), .Z(n4702) );
  XNOR U4830 ( .A(n4704), .B(n4439), .Z(out[1518]) );
  ANDN U4831 ( .B(n4705), .A(n4438), .Z(n4704) );
  XNOR U4832 ( .A(n4706), .B(n4443), .Z(out[1517]) );
  XNOR U4833 ( .A(n4708), .B(n4446), .Z(out[1516]) );
  AND U4834 ( .A(n4709), .B(n4710), .Z(n4708) );
  XNOR U4835 ( .A(n4711), .B(n4455), .Z(out[1515]) );
  ANDN U4836 ( .B(n4712), .A(n4454), .Z(n4711) );
  XNOR U4837 ( .A(n4713), .B(n4458), .Z(out[1514]) );
  NOR U4838 ( .A(n4459), .B(n4714), .Z(n4713) );
  IV U4839 ( .A(n4715), .Z(n4459) );
  XNOR U4840 ( .A(n4716), .B(n4462), .Z(out[1513]) );
  AND U4841 ( .A(n4717), .B(n4463), .Z(n4716) );
  XNOR U4842 ( .A(n4718), .B(n4467), .Z(out[1512]) );
  ANDN U4843 ( .B(n4719), .A(n4466), .Z(n4718) );
  XNOR U4844 ( .A(n4720), .B(n4470), .Z(out[1511]) );
  XOR U4845 ( .A(n4722), .B(n4475), .Z(out[1510]) );
  ANDN U4846 ( .B(n4723), .A(n4474), .Z(n4722) );
  XOR U4847 ( .A(n4724), .B(n3989), .Z(out[150]) );
  XOR U4848 ( .A(n4725), .B(n1997), .Z(n3989) );
  AND U4849 ( .A(n1566), .B(n4208), .Z(n4724) );
  XNOR U4850 ( .A(n4726), .B(n2197), .Z(n4208) );
  XOR U4851 ( .A(n4727), .B(n4728), .Z(n1566) );
  XOR U4852 ( .A(n4729), .B(n4479), .Z(out[1509]) );
  AND U4853 ( .A(n4478), .B(n4730), .Z(n4729) );
  XNOR U4854 ( .A(n4731), .B(n4483), .Z(out[1508]) );
  ANDN U4855 ( .B(n4732), .A(n4482), .Z(n4731) );
  XNOR U4856 ( .A(n4733), .B(n4487), .Z(out[1507]) );
  ANDN U4857 ( .B(n4734), .A(n4486), .Z(n4733) );
  XNOR U4858 ( .A(n4735), .B(n4491), .Z(out[1506]) );
  ANDN U4859 ( .B(n4736), .A(n4490), .Z(n4735) );
  XNOR U4860 ( .A(n4737), .B(n4499), .Z(out[1505]) );
  AND U4861 ( .A(n4500), .B(n4738), .Z(n4737) );
  XNOR U4862 ( .A(n4739), .B(n4504), .Z(out[1504]) );
  ANDN U4863 ( .B(n4740), .A(n4503), .Z(n4739) );
  XOR U4864 ( .A(n4741), .B(n4511), .Z(out[1503]) );
  AND U4865 ( .A(n4742), .B(n4512), .Z(n4741) );
  XNOR U4866 ( .A(n4743), .B(n4515), .Z(out[1502]) );
  AND U4867 ( .A(n4744), .B(n4745), .Z(n4743) );
  XNOR U4868 ( .A(n4746), .B(n4519), .Z(out[1501]) );
  AND U4869 ( .A(n4747), .B(n4748), .Z(n4746) );
  XOR U4870 ( .A(n4749), .B(n4524), .Z(out[1500]) );
  ANDN U4871 ( .B(n4750), .A(n4523), .Z(n4749) );
  XNOR U4872 ( .A(n4751), .B(n1864), .Z(out[14]) );
  NOR U4873 ( .A(n4014), .B(n1863), .Z(n4751) );
  XNOR U4874 ( .A(n2503), .B(n4752), .Z(n1863) );
  XOR U4875 ( .A(n4753), .B(n1733), .Z(n4014) );
  XOR U4876 ( .A(n4754), .B(n3992), .Z(out[149]) );
  XOR U4877 ( .A(n4755), .B(n2000), .Z(n3992) );
  ANDN U4878 ( .B(n1589), .A(n1591), .Z(n4754) );
  XNOR U4879 ( .A(n4756), .B(n2518), .Z(n1591) );
  XNOR U4880 ( .A(n4757), .B(n3793), .Z(n1589) );
  XNOR U4881 ( .A(n4758), .B(n4527), .Z(out[1499]) );
  AND U4882 ( .A(n4759), .B(n4760), .Z(n4758) );
  XOR U4883 ( .A(n4761), .B(n4532), .Z(out[1498]) );
  ANDN U4884 ( .B(n4762), .A(n4531), .Z(n4761) );
  XNOR U4885 ( .A(n4763), .B(n4535), .Z(out[1497]) );
  AND U4886 ( .A(n4764), .B(n4765), .Z(n4763) );
  XNOR U4887 ( .A(n4766), .B(n4539), .Z(out[1496]) );
  AND U4888 ( .A(n4767), .B(n4768), .Z(n4766) );
  XNOR U4889 ( .A(n4769), .B(n4547), .Z(out[1495]) );
  AND U4890 ( .A(n4770), .B(n4548), .Z(n4769) );
  XOR U4891 ( .A(n4771), .B(n4552), .Z(out[1494]) );
  ANDN U4892 ( .B(n4772), .A(n4551), .Z(n4771) );
  XOR U4893 ( .A(n4773), .B(n4556), .Z(out[1493]) );
  NOR U4894 ( .A(n4774), .B(n4555), .Z(n4773) );
  XNOR U4895 ( .A(n4775), .B(n4559), .Z(out[1492]) );
  ANDN U4896 ( .B(n4776), .A(n4560), .Z(n4775) );
  XNOR U4897 ( .A(n4777), .B(n4563), .Z(out[1491]) );
  NOR U4898 ( .A(n4778), .B(n4564), .Z(n4777) );
  XOR U4899 ( .A(n4779), .B(n4568), .Z(out[1490]) );
  ANDN U4900 ( .B(n4780), .A(n4567), .Z(n4779) );
  XNOR U4901 ( .A(n4781), .B(n3996), .Z(out[148]) );
  XNOR U4902 ( .A(n4782), .B(n2003), .Z(n3996) );
  AND U4903 ( .A(n1615), .B(n1614), .Z(n4781) );
  IV U4904 ( .A(n4212), .Z(n1614) );
  XOR U4905 ( .A(n4783), .B(n2211), .Z(n4212) );
  XOR U4906 ( .A(n4784), .B(n2531), .Z(n1615) );
  XNOR U4907 ( .A(n4785), .B(n4571), .Z(out[1489]) );
  NOR U4908 ( .A(n4786), .B(n4572), .Z(n4785) );
  XNOR U4909 ( .A(n4787), .B(n4576), .Z(out[1488]) );
  ANDN U4910 ( .B(n4788), .A(n4575), .Z(n4787) );
  XOR U4911 ( .A(n4789), .B(n4581), .Z(out[1487]) );
  NOR U4912 ( .A(n4790), .B(n4580), .Z(n4789) );
  XOR U4913 ( .A(n4791), .B(n4586), .Z(out[1486]) );
  NOR U4914 ( .A(n4792), .B(n4585), .Z(n4791) );
  XOR U4915 ( .A(n4793), .B(n4595), .Z(out[1485]) );
  ANDN U4916 ( .B(n4794), .A(n4594), .Z(n4793) );
  XOR U4917 ( .A(n4795), .B(n4599), .Z(out[1484]) );
  NOR U4918 ( .A(n4796), .B(n4598), .Z(n4795) );
  XOR U4919 ( .A(n4797), .B(n4603), .Z(out[1483]) );
  NOR U4920 ( .A(n4798), .B(n4602), .Z(n4797) );
  XOR U4921 ( .A(n4799), .B(n4607), .Z(out[1482]) );
  NOR U4922 ( .A(n4606), .B(n4800), .Z(n4799) );
  XNOR U4923 ( .A(n4801), .B(n4610), .Z(out[1481]) );
  ANDN U4924 ( .B(n4802), .A(n4611), .Z(n4801) );
  XNOR U4925 ( .A(n4803), .B(n4614), .Z(out[1480]) );
  ANDN U4926 ( .B(n4804), .A(n4615), .Z(n4803) );
  XOR U4927 ( .A(n4805), .B(n3998), .Z(out[147]) );
  XOR U4928 ( .A(n4806), .B(n2006), .Z(n3998) );
  ANDN U4929 ( .B(n1639), .A(n1638), .Z(n4805) );
  XNOR U4930 ( .A(n4807), .B(n3803), .Z(n1638) );
  XNOR U4931 ( .A(n4808), .B(n2538), .Z(n1639) );
  XNOR U4932 ( .A(n4809), .B(n4618), .Z(out[1479]) );
  NOR U4933 ( .A(n4810), .B(n4619), .Z(n4809) );
  XOR U4934 ( .A(n4811), .B(n4623), .Z(out[1478]) );
  ANDN U4935 ( .B(n4812), .A(n4622), .Z(n4811) );
  XNOR U4936 ( .A(n4813), .B(n4626), .Z(out[1477]) );
  AND U4937 ( .A(n4627), .B(n4814), .Z(n4813) );
  XOR U4938 ( .A(n4815), .B(n4631), .Z(out[1476]) );
  NOR U4939 ( .A(n4816), .B(n4630), .Z(n4815) );
  XNOR U4940 ( .A(n4817), .B(n4641), .Z(out[1475]) );
  NOR U4941 ( .A(n4818), .B(n4642), .Z(n4817) );
  XNOR U4942 ( .A(n4819), .B(n4645), .Z(out[1474]) );
  NOR U4943 ( .A(n4820), .B(n4646), .Z(n4819) );
  XOR U4944 ( .A(n4821), .B(n4652), .Z(out[1473]) );
  ANDN U4945 ( .B(n4822), .A(n4651), .Z(n4821) );
  XNOR U4946 ( .A(n4823), .B(n4657), .Z(out[1472]) );
  ANDN U4947 ( .B(n4824), .A(n4658), .Z(n4823) );
  XOR U4948 ( .A(n4825), .B(n4366), .Z(out[1471]) );
  XNOR U4949 ( .A(n2477), .B(n4826), .Z(n4366) );
  AND U4950 ( .A(n4827), .B(n4828), .Z(n4825) );
  XOR U4951 ( .A(n4829), .B(n4370), .Z(out[1470]) );
  XNOR U4952 ( .A(n4289), .B(n4830), .Z(n4370) );
  IV U4953 ( .A(n2484), .Z(n4289) );
  ANDN U4954 ( .B(n4831), .A(n4662), .Z(n4829) );
  XOR U4955 ( .A(n4832), .B(n4001), .Z(out[146]) );
  XNOR U4956 ( .A(n4833), .B(n4834), .Z(n4001) );
  AND U4957 ( .A(n1667), .B(n1669), .Z(n4832) );
  XNOR U4958 ( .A(n4835), .B(n2543), .Z(n1669) );
  XNOR U4959 ( .A(n4836), .B(n3809), .Z(n1667) );
  XOR U4960 ( .A(n4837), .B(n4374), .Z(out[1469]) );
  XOR U4961 ( .A(n4838), .B(n2492), .Z(n4374) );
  AND U4962 ( .A(n4839), .B(n4840), .Z(n4837) );
  XOR U4963 ( .A(n4841), .B(n4378), .Z(out[1468]) );
  XOR U4964 ( .A(n4354), .B(n4842), .Z(n4378) );
  ANDN U4965 ( .B(n4843), .A(n4666), .Z(n4841) );
  XOR U4966 ( .A(n4844), .B(n4383), .Z(out[1467]) );
  IV U4967 ( .A(n4669), .Z(n4383) );
  XOR U4968 ( .A(n2503), .B(n4845), .Z(n4669) );
  NOR U4969 ( .A(n4846), .B(n4668), .Z(n4844) );
  XNOR U4970 ( .A(n4847), .B(n4387), .Z(out[1466]) );
  XNOR U4971 ( .A(n3465), .B(n4848), .Z(n4387) );
  ANDN U4972 ( .B(n4849), .A(n4671), .Z(n4847) );
  XNOR U4973 ( .A(n4850), .B(n4391), .Z(out[1465]) );
  XOR U4974 ( .A(n3468), .B(n4851), .Z(n4391) );
  ANDN U4975 ( .B(n4852), .A(n4678), .Z(n4850) );
  XOR U4976 ( .A(n4853), .B(n4394), .Z(out[1464]) );
  XNOR U4977 ( .A(n4854), .B(n4855), .Z(n4394) );
  AND U4978 ( .A(n4680), .B(n4856), .Z(n4853) );
  XOR U4979 ( .A(n4857), .B(n4399), .Z(out[1463]) );
  XOR U4980 ( .A(n4858), .B(n4859), .Z(n4399) );
  XOR U4981 ( .A(n4861), .B(n4402), .Z(out[1462]) );
  XNOR U4982 ( .A(n2544), .B(n4862), .Z(n4402) );
  ANDN U4983 ( .B(n4863), .A(n4684), .Z(n4861) );
  XOR U4984 ( .A(n4864), .B(n4410), .Z(out[1461]) );
  XNOR U4985 ( .A(n4865), .B(n2552), .Z(n4410) );
  AND U4986 ( .A(n4866), .B(n4686), .Z(n4864) );
  XOR U4987 ( .A(n4867), .B(n4414), .Z(out[1460]) );
  XNOR U4988 ( .A(n4868), .B(n2559), .Z(n4414) );
  AND U4989 ( .A(n4869), .B(n4688), .Z(n4867) );
  XOR U4990 ( .A(n4870), .B(n4004), .Z(out[145]) );
  XNOR U4991 ( .A(n4871), .B(n2012), .Z(n4004) );
  ANDN U4992 ( .B(n1715), .A(n1716), .Z(n4870) );
  XOR U4993 ( .A(n4872), .B(n3265), .Z(n1716) );
  XNOR U4994 ( .A(n4873), .B(n3815), .Z(n1715) );
  XOR U4995 ( .A(n4874), .B(n4419), .Z(out[1459]) );
  XOR U4996 ( .A(n4875), .B(n3487), .Z(n4419) );
  ANDN U4997 ( .B(n4876), .A(n4690), .Z(n4874) );
  XOR U4998 ( .A(n4877), .B(n4422), .Z(out[1458]) );
  XOR U4999 ( .A(n4878), .B(n2573), .Z(n4422) );
  ANDN U5000 ( .B(n4879), .A(n4692), .Z(n4877) );
  XOR U5001 ( .A(n4880), .B(n4426), .Z(out[1457]) );
  XNOR U5002 ( .A(n4881), .B(n2578), .Z(n4426) );
  ANDN U5003 ( .B(n4882), .A(n4694), .Z(n4880) );
  XOR U5004 ( .A(n4883), .B(n4430), .Z(out[1456]) );
  XNOR U5005 ( .A(n4884), .B(n2587), .Z(n4430) );
  AND U5006 ( .A(n4885), .B(n4696), .Z(n4883) );
  XOR U5007 ( .A(n4886), .B(n4434), .Z(out[1455]) );
  XOR U5008 ( .A(n4887), .B(n2592), .Z(n4434) );
  ANDN U5009 ( .B(n4888), .A(n4703), .Z(n4886) );
  XOR U5010 ( .A(n4889), .B(n4438), .Z(out[1454]) );
  XNOR U5011 ( .A(n4890), .B(n3501), .Z(n4438) );
  ANDN U5012 ( .B(n4891), .A(n4705), .Z(n4889) );
  XOR U5013 ( .A(n4892), .B(n4442), .Z(out[1453]) );
  XOR U5014 ( .A(n4893), .B(n2610), .Z(n4442) );
  AND U5015 ( .A(n4894), .B(n4707), .Z(n4892) );
  XOR U5016 ( .A(n4895), .B(n4447), .Z(out[1452]) );
  IV U5017 ( .A(n4710), .Z(n4447) );
  XOR U5018 ( .A(n4896), .B(n2617), .Z(n4710) );
  ANDN U5019 ( .B(n4897), .A(n4709), .Z(n4895) );
  XOR U5020 ( .A(n4898), .B(n4454), .Z(out[1451]) );
  XNOR U5021 ( .A(n4899), .B(n2624), .Z(n4454) );
  ANDN U5022 ( .B(n4900), .A(n4712), .Z(n4898) );
  XNOR U5023 ( .A(n4901), .B(n4715), .Z(out[1450]) );
  XOR U5024 ( .A(n4902), .B(n2631), .Z(n4715) );
  AND U5025 ( .A(n4714), .B(n4903), .Z(n4901) );
  XOR U5026 ( .A(n4904), .B(n4008), .Z(out[144]) );
  IV U5027 ( .A(n4220), .Z(n4008) );
  XNOR U5028 ( .A(n4905), .B(n2015), .Z(n4220) );
  ANDN U5029 ( .B(n1765), .A(n1766), .Z(n4904) );
  XNOR U5030 ( .A(n4906), .B(n2557), .Z(n1766) );
  XNOR U5031 ( .A(n4907), .B(n2245), .Z(n1765) );
  IV U5032 ( .A(n3822), .Z(n2245) );
  XNOR U5033 ( .A(n4908), .B(n4463), .Z(out[1449]) );
  XOR U5034 ( .A(n4909), .B(n2638), .Z(n4463) );
  ANDN U5035 ( .B(n4910), .A(n4717), .Z(n4908) );
  XOR U5036 ( .A(n4911), .B(n4466), .Z(out[1448]) );
  XOR U5037 ( .A(n4912), .B(n2645), .Z(n4466) );
  ANDN U5038 ( .B(n4913), .A(n4719), .Z(n4911) );
  XNOR U5039 ( .A(n4914), .B(n4471), .Z(out[1447]) );
  XOR U5040 ( .A(n4915), .B(n2652), .Z(n4471) );
  AND U5041 ( .A(n4916), .B(n4721), .Z(n4914) );
  XOR U5042 ( .A(n4917), .B(n4474), .Z(out[1446]) );
  XNOR U5043 ( .A(n4918), .B(n2659), .Z(n4474) );
  XNOR U5044 ( .A(n4920), .B(n4478), .Z(out[1445]) );
  XOR U5045 ( .A(n4921), .B(n2666), .Z(n4478) );
  XOR U5046 ( .A(n4923), .B(n4482), .Z(out[1444]) );
  XOR U5047 ( .A(n4924), .B(n4925), .Z(n4482) );
  XOR U5048 ( .A(n4927), .B(n4486), .Z(out[1443]) );
  XNOR U5049 ( .A(n4928), .B(n4929), .Z(n4486) );
  XOR U5050 ( .A(n4931), .B(n4490), .Z(out[1442]) );
  XOR U5051 ( .A(n4932), .B(n2213), .Z(n4490) );
  ANDN U5052 ( .B(n4933), .A(n4736), .Z(n4931) );
  XNOR U5053 ( .A(n4934), .B(n4500), .Z(out[1441]) );
  XNOR U5054 ( .A(n4935), .B(n2220), .Z(n4500) );
  AND U5055 ( .A(n4936), .B(n4937), .Z(n4934) );
  XOR U5056 ( .A(n4938), .B(n4503), .Z(out[1440]) );
  XNOR U5057 ( .A(n4939), .B(n2235), .Z(n4503) );
  NOR U5058 ( .A(n4940), .B(n4740), .Z(n4938) );
  XOR U5059 ( .A(n4941), .B(n4011), .Z(out[143]) );
  IV U5060 ( .A(n4222), .Z(n4011) );
  XOR U5061 ( .A(n4942), .B(n2018), .Z(n4222) );
  ANDN U5062 ( .B(n1817), .A(n1816), .Z(n4941) );
  XNOR U5063 ( .A(n4943), .B(n2252), .Z(n1816) );
  XOR U5064 ( .A(n4944), .B(n2566), .Z(n1817) );
  XNOR U5065 ( .A(n4945), .B(n4512), .Z(out[1439]) );
  XOR U5066 ( .A(n4946), .B(n2240), .Z(n4512) );
  ANDN U5067 ( .B(n4947), .A(n4742), .Z(n4945) );
  XOR U5068 ( .A(n4948), .B(n4516), .Z(out[1438]) );
  IV U5069 ( .A(n4745), .Z(n4516) );
  XOR U5070 ( .A(n4949), .B(n2247), .Z(n4745) );
  ANDN U5071 ( .B(n4950), .A(n4744), .Z(n4948) );
  XOR U5072 ( .A(n4951), .B(n4520), .Z(out[1437]) );
  IV U5073 ( .A(n4748), .Z(n4520) );
  XOR U5074 ( .A(n4952), .B(n2254), .Z(n4748) );
  XOR U5075 ( .A(n4954), .B(n4523), .Z(out[1436]) );
  XNOR U5076 ( .A(n4955), .B(n2263), .Z(n4523) );
  XOR U5077 ( .A(n4957), .B(n4528), .Z(out[1435]) );
  IV U5078 ( .A(n4760), .Z(n4528) );
  XNOR U5079 ( .A(n4958), .B(n2270), .Z(n4760) );
  NOR U5080 ( .A(n4959), .B(n4759), .Z(n4957) );
  XOR U5081 ( .A(n4960), .B(n4531), .Z(out[1434]) );
  XOR U5082 ( .A(n4961), .B(n2275), .Z(n4531) );
  ANDN U5083 ( .B(n4962), .A(n4762), .Z(n4960) );
  XOR U5084 ( .A(n4963), .B(n4536), .Z(out[1433]) );
  IV U5085 ( .A(n4765), .Z(n4536) );
  XOR U5086 ( .A(n4964), .B(n2282), .Z(n4765) );
  ANDN U5087 ( .B(n4965), .A(n4764), .Z(n4963) );
  XOR U5088 ( .A(n4966), .B(n4540), .Z(out[1432]) );
  IV U5089 ( .A(n4768), .Z(n4540) );
  XOR U5090 ( .A(n4967), .B(n2289), .Z(n4768) );
  ANDN U5091 ( .B(n4968), .A(n4767), .Z(n4966) );
  XNOR U5092 ( .A(n4969), .B(n4548), .Z(out[1431]) );
  XOR U5093 ( .A(n4970), .B(n2296), .Z(n4548) );
  ANDN U5094 ( .B(n4971), .A(n4770), .Z(n4969) );
  XOR U5095 ( .A(n4972), .B(n4551), .Z(out[1430]) );
  XNOR U5096 ( .A(n4973), .B(n2307), .Z(n4551) );
  ANDN U5097 ( .B(n4974), .A(n4772), .Z(n4972) );
  XOR U5098 ( .A(n4975), .B(n4013), .Z(out[142]) );
  XNOR U5099 ( .A(n4976), .B(n2021), .Z(n4013) );
  ANDN U5100 ( .B(n1862), .A(n1864), .Z(n4975) );
  XOR U5101 ( .A(n4977), .B(n2571), .Z(n1864) );
  XNOR U5102 ( .A(n4978), .B(n2259), .Z(n1862) );
  XOR U5103 ( .A(n4979), .B(n4555), .Z(out[1429]) );
  XNOR U5104 ( .A(n3382), .B(n4980), .Z(n4555) );
  ANDN U5105 ( .B(n4774), .A(n4981), .Z(n4979) );
  XOR U5106 ( .A(n4982), .B(n4560), .Z(out[1428]) );
  XNOR U5107 ( .A(n4983), .B(n4984), .Z(n4560) );
  AND U5108 ( .A(n4985), .B(n4986), .Z(n4982) );
  XOR U5109 ( .A(n4987), .B(n4564), .Z(out[1427]) );
  XOR U5110 ( .A(n3392), .B(n4988), .Z(n4564) );
  IV U5111 ( .A(n2329), .Z(n3392) );
  AND U5112 ( .A(n4778), .B(n4989), .Z(n4987) );
  XOR U5113 ( .A(n4990), .B(n4567), .Z(out[1426]) );
  XNOR U5114 ( .A(n3395), .B(n4991), .Z(n4567) );
  ANDN U5115 ( .B(n4992), .A(n4780), .Z(n4990) );
  XOR U5116 ( .A(n4993), .B(n4572), .Z(out[1425]) );
  XOR U5117 ( .A(n2341), .B(n4994), .Z(n4572) );
  AND U5118 ( .A(n4786), .B(n4995), .Z(n4993) );
  XOR U5119 ( .A(n4996), .B(n4575), .Z(out[1424]) );
  XOR U5120 ( .A(n2350), .B(n4997), .Z(n4575) );
  ANDN U5121 ( .B(n4998), .A(n4788), .Z(n4996) );
  XOR U5122 ( .A(n4999), .B(n4580), .Z(out[1423]) );
  XNOR U5123 ( .A(n2357), .B(n5000), .Z(n4580) );
  AND U5124 ( .A(n5001), .B(n4790), .Z(n4999) );
  IV U5125 ( .A(n5002), .Z(n4790) );
  XOR U5126 ( .A(n5003), .B(n4585), .Z(out[1422]) );
  XNOR U5127 ( .A(n2364), .B(n5004), .Z(n4585) );
  AND U5128 ( .A(n4792), .B(n5005), .Z(n5003) );
  XOR U5129 ( .A(n5006), .B(n4594), .Z(out[1421]) );
  XNOR U5130 ( .A(n5007), .B(n5008), .Z(n4594) );
  XOR U5131 ( .A(n5010), .B(n4598), .Z(out[1420]) );
  XNOR U5132 ( .A(n2382), .B(n5011), .Z(n4598) );
  AND U5133 ( .A(n4796), .B(n5012), .Z(n5010) );
  XOR U5134 ( .A(n5013), .B(n4019), .Z(out[141]) );
  XNOR U5135 ( .A(n5014), .B(n2024), .Z(n4019) );
  AND U5136 ( .A(n1910), .B(n1908), .Z(n5013) );
  XOR U5137 ( .A(n5015), .B(n2266), .Z(n1908) );
  IV U5138 ( .A(n3839), .Z(n2266) );
  XOR U5139 ( .A(n5016), .B(n4602), .Z(out[1419]) );
  XOR U5140 ( .A(n5017), .B(n2388), .Z(n4602) );
  AND U5141 ( .A(n4798), .B(n5018), .Z(n5016) );
  XOR U5142 ( .A(n5019), .B(n4606), .Z(out[1418]) );
  XNOR U5143 ( .A(n5020), .B(n2395), .Z(n4606) );
  AND U5144 ( .A(n4800), .B(n5021), .Z(n5019) );
  XOR U5145 ( .A(n5022), .B(n4611), .Z(out[1417]) );
  XNOR U5146 ( .A(n2403), .B(n5023), .Z(n4611) );
  AND U5147 ( .A(n5024), .B(n5025), .Z(n5022) );
  XOR U5148 ( .A(n5026), .B(n4615), .Z(out[1416]) );
  XOR U5149 ( .A(n2408), .B(n5027), .Z(n4615) );
  XOR U5150 ( .A(n5029), .B(n4619), .Z(out[1415]) );
  XOR U5151 ( .A(n4016), .B(n5030), .Z(n4619) );
  AND U5152 ( .A(n4810), .B(n5031), .Z(n5029) );
  XOR U5153 ( .A(n5032), .B(n4622), .Z(out[1414]) );
  XNOR U5154 ( .A(n4053), .B(n5033), .Z(n4622) );
  ANDN U5155 ( .B(n5034), .A(n4812), .Z(n5032) );
  XNOR U5156 ( .A(n5035), .B(n4627), .Z(out[1413]) );
  XNOR U5157 ( .A(n4087), .B(n5036), .Z(n4627) );
  AND U5158 ( .A(n5037), .B(n5038), .Z(n5035) );
  XOR U5159 ( .A(n5039), .B(n4630), .Z(out[1412]) );
  XNOR U5160 ( .A(n5040), .B(n5041), .Z(n4630) );
  AND U5161 ( .A(n4816), .B(n5042), .Z(n5039) );
  XOR U5162 ( .A(n5043), .B(n4642), .Z(out[1411]) );
  XNOR U5163 ( .A(n2443), .B(n5044), .Z(n4642) );
  AND U5164 ( .A(n4818), .B(n5045), .Z(n5043) );
  XOR U5165 ( .A(n5046), .B(n4646), .Z(out[1410]) );
  XNOR U5166 ( .A(n4191), .B(n5047), .Z(n4646) );
  AND U5167 ( .A(n4820), .B(n5048), .Z(n5046) );
  XNOR U5168 ( .A(n5049), .B(n4023), .Z(out[140]) );
  XOR U5169 ( .A(n5050), .B(n2031), .Z(n4023) );
  AND U5170 ( .A(n1957), .B(n1956), .Z(n5049) );
  IV U5171 ( .A(n4226), .Z(n1956) );
  XOR U5172 ( .A(n5051), .B(n2273), .Z(n4226) );
  IV U5173 ( .A(n3845), .Z(n2273) );
  XOR U5174 ( .A(n5052), .B(n4651), .Z(out[1409]) );
  XNOR U5175 ( .A(n5053), .B(n5054), .Z(n4651) );
  AND U5176 ( .A(n5055), .B(n5056), .Z(n5052) );
  XOR U5177 ( .A(n5057), .B(n4658), .Z(out[1408]) );
  XNOR U5178 ( .A(n2468), .B(n5058), .Z(n4658) );
  AND U5179 ( .A(n5059), .B(n5060), .Z(n5057) );
  XOR U5180 ( .A(n5061), .B(n4660), .Z(out[1407]) );
  IV U5181 ( .A(n4828), .Z(n4660) );
  XOR U5182 ( .A(n1947), .B(n5062), .Z(n4828) );
  XOR U5183 ( .A(n5063), .B(n4662), .Z(out[1406]) );
  XNOR U5184 ( .A(n5064), .B(n1953), .Z(n4662) );
  NOR U5185 ( .A(n4831), .B(n4369), .Z(n5063) );
  XOR U5186 ( .A(n5065), .B(n4664), .Z(out[1405]) );
  IV U5187 ( .A(n4840), .Z(n4664) );
  XNOR U5188 ( .A(n5066), .B(n1961), .Z(n4840) );
  NOR U5189 ( .A(n4839), .B(n4373), .Z(n5065) );
  XOR U5190 ( .A(n5067), .B(n4666), .Z(out[1404]) );
  XOR U5191 ( .A(n5068), .B(n1965), .Z(n4666) );
  ANDN U5192 ( .B(n4377), .A(n4843), .Z(n5067) );
  XOR U5193 ( .A(n5069), .B(n4668), .Z(out[1403]) );
  XNOR U5194 ( .A(n5070), .B(n1660), .Z(n4668) );
  ANDN U5195 ( .B(n4846), .A(n4381), .Z(n5069) );
  XOR U5196 ( .A(n5071), .B(n4671), .Z(out[1402]) );
  XOR U5197 ( .A(n5072), .B(n1664), .Z(n4671) );
  ANDN U5198 ( .B(n4385), .A(n4849), .Z(n5071) );
  XOR U5199 ( .A(n5073), .B(n4678), .Z(out[1401]) );
  XOR U5200 ( .A(n5074), .B(n1672), .Z(n4678) );
  AND U5201 ( .A(n4389), .B(n5075), .Z(n5073) );
  XNOR U5202 ( .A(n5076), .B(n4680), .Z(out[1400]) );
  XNOR U5203 ( .A(n5077), .B(n3735), .Z(n4680) );
  NOR U5204 ( .A(n4856), .B(n4393), .Z(n5076) );
  XOR U5205 ( .A(n5078), .B(n1910), .Z(out[13]) );
  XNOR U5206 ( .A(n5079), .B(n2580), .Z(n1910) );
  AND U5207 ( .A(n1909), .B(n4020), .Z(n5078) );
  XNOR U5208 ( .A(n5080), .B(n1738), .Z(n4020) );
  XNOR U5209 ( .A(n2510), .B(n5081), .Z(n1909) );
  XOR U5210 ( .A(n5082), .B(n4025), .Z(out[139]) );
  XNOR U5211 ( .A(n5083), .B(n2034), .Z(n4025) );
  AND U5212 ( .A(n1994), .B(n1992), .Z(n5082) );
  XOR U5213 ( .A(n5084), .B(n2280), .Z(n1992) );
  IV U5214 ( .A(n3849), .Z(n2280) );
  XOR U5215 ( .A(n5085), .B(n4682), .Z(out[1399]) );
  XOR U5216 ( .A(n5086), .B(n1682), .Z(n4682) );
  ANDN U5217 ( .B(n4860), .A(n4397), .Z(n5085) );
  XOR U5218 ( .A(n5087), .B(n4684), .Z(out[1398]) );
  XOR U5219 ( .A(n5088), .B(n1686), .Z(n4684) );
  NOR U5220 ( .A(n4863), .B(n4401), .Z(n5087) );
  XNOR U5221 ( .A(n5089), .B(n4686), .Z(out[1397]) );
  XNOR U5222 ( .A(n5090), .B(n1690), .Z(n4686) );
  XNOR U5223 ( .A(n5091), .B(n4688), .Z(out[1396]) );
  XNOR U5224 ( .A(n5092), .B(n1694), .Z(n4688) );
  ANDN U5225 ( .B(n4413), .A(n4869), .Z(n5091) );
  XOR U5226 ( .A(n5093), .B(n4690), .Z(out[1395]) );
  XOR U5227 ( .A(n5094), .B(n1698), .Z(n4690) );
  AND U5228 ( .A(n4417), .B(n5095), .Z(n5093) );
  XOR U5229 ( .A(n5096), .B(n4692), .Z(out[1394]) );
  XOR U5230 ( .A(n5097), .B(n1703), .Z(n4692) );
  NOR U5231 ( .A(n4879), .B(n4421), .Z(n5096) );
  XOR U5232 ( .A(n5098), .B(n4694), .Z(out[1393]) );
  XOR U5233 ( .A(n5099), .B(n1707), .Z(n4694) );
  AND U5234 ( .A(n4425), .B(n5100), .Z(n5098) );
  XNOR U5235 ( .A(n5101), .B(n4696), .Z(out[1392]) );
  XNOR U5236 ( .A(n5102), .B(n1711), .Z(n4696) );
  ANDN U5237 ( .B(n4429), .A(n4885), .Z(n5101) );
  XOR U5238 ( .A(n5103), .B(n4703), .Z(out[1391]) );
  XNOR U5239 ( .A(n5104), .B(n1720), .Z(n4703) );
  AND U5240 ( .A(n4433), .B(n5105), .Z(n5103) );
  XOR U5241 ( .A(n5106), .B(n4705), .Z(out[1390]) );
  XNOR U5242 ( .A(n5107), .B(n1725), .Z(n4705) );
  ANDN U5243 ( .B(n4437), .A(n4891), .Z(n5106) );
  XNOR U5244 ( .A(n5108), .B(n4029), .Z(out[138]) );
  XNOR U5245 ( .A(n5109), .B(n2037), .Z(n4029) );
  AND U5246 ( .A(n2026), .B(n2028), .Z(n5108) );
  XNOR U5247 ( .A(n5110), .B(n2287), .Z(n2026) );
  XNOR U5248 ( .A(n5111), .B(n4707), .Z(out[1389]) );
  XNOR U5249 ( .A(n5112), .B(n1729), .Z(n4707) );
  ANDN U5250 ( .B(n4441), .A(n4894), .Z(n5111) );
  XOR U5251 ( .A(n5113), .B(n4709), .Z(out[1388]) );
  XNOR U5252 ( .A(n5114), .B(n1733), .Z(n4709) );
  AND U5253 ( .A(n4445), .B(n5115), .Z(n5113) );
  XOR U5254 ( .A(n5116), .B(n4712), .Z(out[1387]) );
  XNOR U5255 ( .A(n5117), .B(n1738), .Z(n4712) );
  NOR U5256 ( .A(n4900), .B(n4453), .Z(n5116) );
  XNOR U5257 ( .A(n5118), .B(n4714), .Z(out[1386]) );
  XNOR U5258 ( .A(n5119), .B(n3806), .Z(n4714) );
  NOR U5259 ( .A(n4903), .B(n4457), .Z(n5118) );
  XOR U5260 ( .A(n5120), .B(n4717), .Z(out[1385]) );
  XNOR U5261 ( .A(n5121), .B(n1747), .Z(n4717) );
  ANDN U5262 ( .B(n4461), .A(n4910), .Z(n5120) );
  XOR U5263 ( .A(n5122), .B(n4719), .Z(out[1384]) );
  XNOR U5264 ( .A(n5123), .B(n3818), .Z(n4719) );
  NOR U5265 ( .A(n4913), .B(n4465), .Z(n5122) );
  XNOR U5266 ( .A(n5124), .B(n4721), .Z(out[1383]) );
  XOR U5267 ( .A(n1756), .B(n5125), .Z(n4721) );
  ANDN U5268 ( .B(n4469), .A(n4916), .Z(n5124) );
  XOR U5269 ( .A(n5126), .B(n4723), .Z(out[1382]) );
  XOR U5270 ( .A(n5127), .B(n1762), .Z(n4723) );
  IV U5271 ( .A(n5128), .Z(n1762) );
  ANDN U5272 ( .B(n4473), .A(n4919), .Z(n5126) );
  XOR U5273 ( .A(n5129), .B(n4730), .Z(out[1381]) );
  XOR U5274 ( .A(n5130), .B(n1770), .Z(n4730) );
  IV U5275 ( .A(n5131), .Z(n1770) );
  ANDN U5276 ( .B(n4477), .A(n4922), .Z(n5129) );
  XOR U5277 ( .A(n5132), .B(n4732), .Z(out[1380]) );
  XOR U5278 ( .A(n5133), .B(n1775), .Z(n4732) );
  IV U5279 ( .A(n3842), .Z(n1775) );
  NOR U5280 ( .A(n4926), .B(n4481), .Z(n5132) );
  XOR U5281 ( .A(n5134), .B(n4033), .Z(out[137]) );
  XNOR U5282 ( .A(n5135), .B(n5136), .Z(n4033) );
  AND U5283 ( .A(n1034), .B(n2066), .Z(n5134) );
  IV U5284 ( .A(n4231), .Z(n2066) );
  XOR U5285 ( .A(n5137), .B(n5138), .Z(n4231) );
  XNOR U5286 ( .A(n5139), .B(n2611), .Z(n1034) );
  XOR U5287 ( .A(n5140), .B(n4734), .Z(out[1379]) );
  XOR U5288 ( .A(n5141), .B(n1780), .Z(n4734) );
  IV U5289 ( .A(n5142), .Z(n1780) );
  ANDN U5290 ( .B(n4485), .A(n4930), .Z(n5140) );
  XOR U5291 ( .A(n5143), .B(n4736), .Z(out[1378]) );
  XOR U5292 ( .A(n5144), .B(n4249), .Z(n4736) );
  AND U5293 ( .A(n4489), .B(n5145), .Z(n5143) );
  XOR U5294 ( .A(n5146), .B(n4738), .Z(out[1377]) );
  IV U5295 ( .A(n4937), .Z(n4738) );
  XOR U5296 ( .A(n5147), .B(n1788), .Z(n4937) );
  IV U5297 ( .A(n5148), .Z(n1788) );
  XOR U5298 ( .A(n5149), .B(n4740), .Z(out[1376]) );
  XOR U5299 ( .A(n1792), .B(n5150), .Z(n4740) );
  ANDN U5300 ( .B(n4940), .A(n4502), .Z(n5149) );
  XOR U5301 ( .A(n5151), .B(n4742), .Z(out[1375]) );
  XNOR U5302 ( .A(n5152), .B(n1797), .Z(n4742) );
  ANDN U5303 ( .B(n4505), .A(n4947), .Z(n5151) );
  XOR U5304 ( .A(n5153), .B(n4744), .Z(out[1374]) );
  XNOR U5305 ( .A(n1800), .B(n5154), .Z(n4744) );
  XOR U5306 ( .A(n5155), .B(n4747), .Z(out[1373]) );
  XNOR U5307 ( .A(n1804), .B(n5156), .Z(n4747) );
  ANDN U5308 ( .B(n4953), .A(n4518), .Z(n5155) );
  XOR U5309 ( .A(n5157), .B(n4750), .Z(out[1372]) );
  XOR U5310 ( .A(n5158), .B(n5159), .Z(n4750) );
  NOR U5311 ( .A(n4522), .B(n4956), .Z(n5157) );
  XOR U5312 ( .A(n5160), .B(n4759), .Z(out[1371]) );
  XNOR U5313 ( .A(n5161), .B(n5162), .Z(n4759) );
  AND U5314 ( .A(n4959), .B(n4526), .Z(n5160) );
  IV U5315 ( .A(n5163), .Z(n4526) );
  XOR U5316 ( .A(n5164), .B(n4762), .Z(out[1370]) );
  XNOR U5317 ( .A(n3561), .B(n5165), .Z(n4762) );
  XOR U5318 ( .A(n5166), .B(n4037), .Z(out[136]) );
  XNOR U5319 ( .A(n5167), .B(n2046), .Z(n4037) );
  AND U5320 ( .A(n2101), .B(n1478), .Z(n5166) );
  IV U5321 ( .A(n2102), .Z(n1478) );
  XOR U5322 ( .A(n5168), .B(n3298), .Z(n2102) );
  XNOR U5323 ( .A(n5169), .B(n5170), .Z(n2101) );
  XOR U5324 ( .A(n5171), .B(n4764), .Z(out[1369]) );
  XOR U5325 ( .A(n1828), .B(n5172), .Z(n4764) );
  ANDN U5326 ( .B(n4534), .A(n4965), .Z(n5171) );
  XOR U5327 ( .A(n5173), .B(n4767), .Z(out[1368]) );
  XOR U5328 ( .A(n1832), .B(n5174), .Z(n4767) );
  ANDN U5329 ( .B(n4538), .A(n4968), .Z(n5173) );
  XOR U5330 ( .A(n5175), .B(n4770), .Z(out[1367]) );
  XOR U5331 ( .A(n1837), .B(n5176), .Z(n4770) );
  ANDN U5332 ( .B(n4546), .A(n4971), .Z(n5175) );
  XOR U5333 ( .A(n5177), .B(n4772), .Z(out[1366]) );
  XNOR U5334 ( .A(n3585), .B(n5178), .Z(n4772) );
  AND U5335 ( .A(n4550), .B(n5179), .Z(n5177) );
  XNOR U5336 ( .A(n5180), .B(n4774), .Z(out[1365]) );
  XNOR U5337 ( .A(n1845), .B(n5181), .Z(n4774) );
  ANDN U5338 ( .B(n4981), .A(n4554), .Z(n5180) );
  XOR U5339 ( .A(n5182), .B(n4776), .Z(out[1364]) );
  IV U5340 ( .A(n4986), .Z(n4776) );
  XOR U5341 ( .A(n4098), .B(n5183), .Z(n4986) );
  NOR U5342 ( .A(n4558), .B(n4985), .Z(n5182) );
  XNOR U5343 ( .A(n5184), .B(n4778), .Z(out[1363]) );
  XNOR U5344 ( .A(n4102), .B(n5185), .Z(n4778) );
  NOR U5345 ( .A(n4562), .B(n4989), .Z(n5184) );
  XOR U5346 ( .A(n5186), .B(n4780), .Z(out[1362]) );
  XNOR U5347 ( .A(n5187), .B(n5188), .Z(n4780) );
  NOR U5348 ( .A(n4566), .B(n4992), .Z(n5186) );
  XNOR U5349 ( .A(n5189), .B(n4786), .Z(out[1361]) );
  XNOR U5350 ( .A(n5190), .B(n5191), .Z(n4786) );
  NOR U5351 ( .A(n4995), .B(n4570), .Z(n5189) );
  XOR U5352 ( .A(n5192), .B(n4788), .Z(out[1360]) );
  XNOR U5353 ( .A(n5193), .B(n5194), .Z(n4788) );
  NOR U5354 ( .A(n4574), .B(n4998), .Z(n5192) );
  XOR U5355 ( .A(n5195), .B(n4040), .Z(out[135]) );
  IV U5356 ( .A(n4242), .Z(n4040) );
  XNOR U5357 ( .A(n5196), .B(n2049), .Z(n4242) );
  AND U5358 ( .A(n2138), .B(n1812), .Z(n5195) );
  IV U5359 ( .A(n2139), .Z(n1812) );
  XOR U5360 ( .A(n5197), .B(n3302), .Z(n2139) );
  IV U5361 ( .A(n2626), .Z(n3302) );
  XOR U5362 ( .A(n5198), .B(n2312), .Z(n2138) );
  XOR U5363 ( .A(n5199), .B(n5002), .Z(out[1359]) );
  XOR U5364 ( .A(n4115), .B(n5200), .Z(n5002) );
  NOR U5365 ( .A(n4582), .B(n5001), .Z(n5199) );
  XNOR U5366 ( .A(n5201), .B(n4792), .Z(out[1358]) );
  XOR U5367 ( .A(n5202), .B(n5203), .Z(n4792) );
  XOR U5368 ( .A(n5204), .B(n4794), .Z(out[1357]) );
  XOR U5369 ( .A(n1883), .B(n5205), .Z(n4794) );
  NOR U5370 ( .A(n4593), .B(n5009), .Z(n5204) );
  XNOR U5371 ( .A(n5206), .B(n4796), .Z(out[1356]) );
  XOR U5372 ( .A(n1888), .B(n5207), .Z(n4796) );
  AND U5373 ( .A(n4597), .B(n5208), .Z(n5206) );
  XNOR U5374 ( .A(n5209), .B(n4798), .Z(out[1355]) );
  XNOR U5375 ( .A(n3639), .B(n5210), .Z(n4798) );
  NOR U5376 ( .A(n4601), .B(n5018), .Z(n5209) );
  XNOR U5377 ( .A(n5211), .B(n4800), .Z(out[1354]) );
  XNOR U5378 ( .A(n5212), .B(n5213), .Z(n4800) );
  ANDN U5379 ( .B(n4605), .A(n5021), .Z(n5211) );
  XOR U5380 ( .A(n5214), .B(n4802), .Z(out[1353]) );
  IV U5381 ( .A(n5025), .Z(n4802) );
  XOR U5382 ( .A(n5215), .B(n5216), .Z(n5025) );
  ANDN U5383 ( .B(n4609), .A(n5024), .Z(n5214) );
  XOR U5384 ( .A(n5217), .B(n4804), .Z(out[1352]) );
  XOR U5385 ( .A(n3656), .B(n5218), .Z(n4804) );
  NOR U5386 ( .A(n5028), .B(n4613), .Z(n5217) );
  XNOR U5387 ( .A(n5219), .B(n4810), .Z(out[1351]) );
  XNOR U5388 ( .A(n5220), .B(n5221), .Z(n4810) );
  XOR U5389 ( .A(n5222), .B(n4812), .Z(out[1350]) );
  XNOR U5390 ( .A(n5223), .B(n5224), .Z(n4812) );
  ANDN U5391 ( .B(n4621), .A(n5034), .Z(n5222) );
  XOR U5392 ( .A(n5225), .B(n4043), .Z(out[134]) );
  XOR U5393 ( .A(n5226), .B(n2052), .Z(n4043) );
  AND U5394 ( .A(n2174), .B(n2176), .Z(n5225) );
  XOR U5395 ( .A(n5227), .B(n3306), .Z(n2176) );
  IV U5396 ( .A(n2633), .Z(n3306) );
  XOR U5397 ( .A(n5228), .B(n5229), .Z(n2174) );
  XOR U5398 ( .A(n5230), .B(n4814), .Z(out[1349]) );
  IV U5399 ( .A(n5038), .Z(n4814) );
  XOR U5400 ( .A(n5231), .B(n5232), .Z(n5038) );
  XNOR U5401 ( .A(n5233), .B(n4816), .Z(out[1348]) );
  XNOR U5402 ( .A(n1926), .B(n5234), .Z(n4816) );
  XNOR U5403 ( .A(n5235), .B(n4818), .Z(out[1347]) );
  XNOR U5404 ( .A(n5236), .B(n5237), .Z(n4818) );
  ANDN U5405 ( .B(n4636), .A(n5045), .Z(n5235) );
  XNOR U5406 ( .A(n5238), .B(n4820), .Z(out[1346]) );
  XNOR U5407 ( .A(n3689), .B(n5239), .Z(n4820) );
  ANDN U5408 ( .B(n4644), .A(n5048), .Z(n5238) );
  XOR U5409 ( .A(n5240), .B(n4822), .Z(out[1345]) );
  IV U5410 ( .A(n5056), .Z(n4822) );
  XNOR U5411 ( .A(n1939), .B(n5241), .Z(n5056) );
  NOR U5412 ( .A(n4647), .B(n5055), .Z(n5240) );
  XOR U5413 ( .A(n5242), .B(n4824), .Z(out[1344]) );
  IV U5414 ( .A(n5060), .Z(n4824) );
  XOR U5415 ( .A(n1943), .B(n5243), .Z(n5060) );
  NOR U5416 ( .A(n5059), .B(n4653), .Z(n5242) );
  XOR U5417 ( .A(n5244), .B(n4827), .Z(out[1343]) );
  XOR U5418 ( .A(n5245), .B(n1987), .Z(n4827) );
  IV U5419 ( .A(n3813), .Z(n1987) );
  AND U5420 ( .A(n4360), .B(n4367), .Z(n5244) );
  XOR U5421 ( .A(n5246), .B(n2518), .Z(n4367) );
  XNOR U5422 ( .A(n5247), .B(n2541), .Z(n4360) );
  XOR U5423 ( .A(n5248), .B(n4831), .Z(out[1342]) );
  XNOR U5424 ( .A(n5249), .B(n3820), .Z(n4831) );
  AND U5425 ( .A(n4369), .B(n4371), .Z(n5248) );
  XNOR U5426 ( .A(n5250), .B(n2531), .Z(n4371) );
  XOR U5427 ( .A(n5251), .B(n2548), .Z(n4369) );
  XOR U5428 ( .A(n5252), .B(n4839), .Z(out[1341]) );
  XNOR U5429 ( .A(n5253), .B(n1997), .Z(n4839) );
  AND U5430 ( .A(n4375), .B(n4373), .Z(n5252) );
  XOR U5431 ( .A(n5254), .B(n2555), .Z(n4373) );
  XNOR U5432 ( .A(n5255), .B(n3258), .Z(n4375) );
  IV U5433 ( .A(n2538), .Z(n3258) );
  XOR U5434 ( .A(n5256), .B(n4843), .Z(out[1340]) );
  XOR U5435 ( .A(n5257), .B(n2000), .Z(n4843) );
  NOR U5436 ( .A(n4379), .B(n4377), .Z(n5256) );
  XNOR U5437 ( .A(n5258), .B(n2562), .Z(n4377) );
  XOR U5438 ( .A(n5259), .B(n2543), .Z(n4379) );
  XOR U5439 ( .A(n5260), .B(n4046), .Z(out[133]) );
  XNOR U5440 ( .A(n5261), .B(n2056), .Z(n4046) );
  AND U5441 ( .A(n2226), .B(n2228), .Z(n5260) );
  XOR U5442 ( .A(n5262), .B(n2640), .Z(n2228) );
  XNOR U5443 ( .A(n5263), .B(n5264), .Z(n2226) );
  XNOR U5444 ( .A(n5265), .B(n4846), .Z(out[1339]) );
  XNOR U5445 ( .A(n5266), .B(n2003), .Z(n4846) );
  IV U5446 ( .A(n3837), .Z(n2003) );
  ANDN U5447 ( .B(n4381), .A(n4382), .Z(n5265) );
  XOR U5448 ( .A(n5267), .B(n3265), .Z(n4382) );
  IV U5449 ( .A(n2550), .Z(n3265) );
  XOR U5450 ( .A(n5268), .B(n2569), .Z(n4381) );
  XOR U5451 ( .A(n5269), .B(n4849), .Z(out[1338]) );
  XOR U5452 ( .A(n5270), .B(n2006), .Z(n4849) );
  NOR U5453 ( .A(n4386), .B(n4385), .Z(n5269) );
  XOR U5454 ( .A(n2575), .B(n5271), .Z(n4385) );
  IV U5455 ( .A(n5272), .Z(n2575) );
  XNOR U5456 ( .A(n5273), .B(n2557), .Z(n4386) );
  XOR U5457 ( .A(n5274), .B(n4852), .Z(out[1337]) );
  IV U5458 ( .A(n5075), .Z(n4852) );
  XOR U5459 ( .A(n5275), .B(n2009), .Z(n5075) );
  IV U5460 ( .A(n4834), .Z(n2009) );
  NOR U5461 ( .A(n4390), .B(n4389), .Z(n5274) );
  XOR U5462 ( .A(n2582), .B(n5276), .Z(n4389) );
  IV U5463 ( .A(n5277), .Z(n2582) );
  XOR U5464 ( .A(n5278), .B(n2566), .Z(n4390) );
  XOR U5465 ( .A(n5279), .B(n4856), .Z(out[1336]) );
  XOR U5466 ( .A(n5280), .B(n5281), .Z(n4856) );
  ANDN U5467 ( .B(n4393), .A(n4395), .Z(n5279) );
  XNOR U5468 ( .A(n5282), .B(n2571), .Z(n4395) );
  IV U5469 ( .A(n5283), .Z(n2571) );
  XNOR U5470 ( .A(n2589), .B(n5284), .Z(n4393) );
  IV U5471 ( .A(n4343), .Z(n2589) );
  XNOR U5472 ( .A(n5285), .B(n4860), .Z(out[1335]) );
  XOR U5473 ( .A(n5286), .B(n2015), .Z(n4860) );
  ANDN U5474 ( .B(n4397), .A(n4398), .Z(n5285) );
  XNOR U5475 ( .A(n5287), .B(n2580), .Z(n4398) );
  XOR U5476 ( .A(n5288), .B(n2601), .Z(n4397) );
  XOR U5477 ( .A(n5289), .B(n4863), .Z(out[1334]) );
  XOR U5478 ( .A(n5290), .B(n2018), .Z(n4863) );
  ANDN U5479 ( .B(n4401), .A(n4403), .Z(n5289) );
  XNOR U5480 ( .A(n5291), .B(n2585), .Z(n4403) );
  IV U5481 ( .A(n5292), .Z(n2585) );
  XOR U5482 ( .A(n5293), .B(n2608), .Z(n4401) );
  XOR U5483 ( .A(n5294), .B(n4866), .Z(out[1333]) );
  XNOR U5484 ( .A(n5295), .B(n2021), .Z(n4866) );
  AND U5485 ( .A(n4411), .B(n4409), .Z(n5294) );
  XOR U5486 ( .A(n5296), .B(n2615), .Z(n4409) );
  XNOR U5487 ( .A(n5297), .B(n5298), .Z(n4411) );
  XOR U5488 ( .A(n5299), .B(n4869), .Z(out[1332]) );
  XOR U5489 ( .A(n5300), .B(n2024), .Z(n4869) );
  ANDN U5490 ( .B(n4415), .A(n4413), .Z(n5299) );
  XOR U5491 ( .A(n5301), .B(n2622), .Z(n4413) );
  XNOR U5492 ( .A(n5302), .B(n5303), .Z(n4415) );
  XOR U5493 ( .A(n5304), .B(n4876), .Z(out[1331]) );
  IV U5494 ( .A(n5095), .Z(n4876) );
  XOR U5495 ( .A(n5305), .B(n2031), .Z(n5095) );
  NOR U5496 ( .A(n4418), .B(n4417), .Z(n5304) );
  XNOR U5497 ( .A(n5306), .B(n3758), .Z(n4417) );
  XOR U5498 ( .A(n2611), .B(n5307), .Z(n4418) );
  IV U5499 ( .A(n5308), .Z(n2611) );
  XOR U5500 ( .A(n5309), .B(n4879), .Z(out[1330]) );
  XOR U5501 ( .A(n5310), .B(n2034), .Z(n4879) );
  ANDN U5502 ( .B(n4421), .A(n4423), .Z(n5309) );
  XNOR U5503 ( .A(n5311), .B(n3298), .Z(n4423) );
  IV U5504 ( .A(n2619), .Z(n3298) );
  XOR U5505 ( .A(n5312), .B(n2636), .Z(n4421) );
  XOR U5506 ( .A(n5313), .B(n4049), .Z(out[132]) );
  XOR U5507 ( .A(n5314), .B(n2059), .Z(n4049) );
  ANDN U5508 ( .B(n4250), .A(n2302), .Z(n5313) );
  XNOR U5509 ( .A(n5315), .B(n2647), .Z(n2302) );
  XOR U5510 ( .A(n5316), .B(n2333), .Z(n4250) );
  XOR U5511 ( .A(n5317), .B(n4882), .Z(out[1329]) );
  IV U5512 ( .A(n5100), .Z(n4882) );
  XOR U5513 ( .A(n5318), .B(n2037), .Z(n5100) );
  ANDN U5514 ( .B(n4427), .A(n4425), .Z(n5317) );
  XOR U5515 ( .A(n5319), .B(n4591), .Z(n4425) );
  IV U5516 ( .A(n2643), .Z(n4591) );
  XNOR U5517 ( .A(n5320), .B(n2626), .Z(n4427) );
  XOR U5518 ( .A(n5321), .B(n4885), .Z(out[1328]) );
  XOR U5519 ( .A(n5322), .B(n5136), .Z(n4885) );
  ANDN U5520 ( .B(n4431), .A(n4429), .Z(n5321) );
  XOR U5521 ( .A(n5323), .B(n3773), .Z(n4429) );
  XNOR U5522 ( .A(n5324), .B(n2633), .Z(n4431) );
  XOR U5523 ( .A(n5325), .B(n4888), .Z(out[1327]) );
  IV U5524 ( .A(n5105), .Z(n4888) );
  XOR U5525 ( .A(n5326), .B(n2046), .Z(n5105) );
  NOR U5526 ( .A(n4435), .B(n4433), .Z(n5325) );
  XNOR U5527 ( .A(n5327), .B(n2657), .Z(n4433) );
  XNOR U5528 ( .A(n5328), .B(n2640), .Z(n4435) );
  IV U5529 ( .A(n5329), .Z(n2640) );
  XOR U5530 ( .A(n5330), .B(n4891), .Z(out[1326]) );
  XNOR U5531 ( .A(n5331), .B(n2049), .Z(n4891) );
  NOR U5532 ( .A(n4439), .B(n4437), .Z(n5330) );
  XOR U5533 ( .A(n5332), .B(n2664), .Z(n4437) );
  XOR U5534 ( .A(n5333), .B(n2647), .Z(n4439) );
  IV U5535 ( .A(n5334), .Z(n2647) );
  XOR U5536 ( .A(n5335), .B(n4894), .Z(out[1325]) );
  XOR U5537 ( .A(n5336), .B(n2052), .Z(n4894) );
  IV U5538 ( .A(n5337), .Z(n2052) );
  NOR U5539 ( .A(n4443), .B(n4441), .Z(n5335) );
  XNOR U5540 ( .A(n5338), .B(n2197), .Z(n4441) );
  XOR U5541 ( .A(n5339), .B(n2654), .Z(n4443) );
  XOR U5542 ( .A(n5340), .B(n4897), .Z(out[1324]) );
  IV U5543 ( .A(n5115), .Z(n4897) );
  XNOR U5544 ( .A(n5341), .B(n2056), .Z(n5115) );
  NOR U5545 ( .A(n4446), .B(n4445), .Z(n5340) );
  XNOR U5546 ( .A(n5342), .B(n2204), .Z(n4445) );
  XOR U5547 ( .A(n5343), .B(n3324), .Z(n4446) );
  XOR U5548 ( .A(n5344), .B(n4900), .Z(out[1323]) );
  XNOR U5549 ( .A(n5345), .B(n2059), .Z(n4900) );
  IV U5550 ( .A(n5346), .Z(n2059) );
  ANDN U5551 ( .B(n4453), .A(n4455), .Z(n5344) );
  XNOR U5552 ( .A(n5347), .B(n2668), .Z(n4455) );
  XOR U5553 ( .A(n5348), .B(n2211), .Z(n4453) );
  IV U5554 ( .A(n5349), .Z(n2211) );
  XOR U5555 ( .A(n5350), .B(n4903), .Z(out[1322]) );
  XOR U5556 ( .A(n5351), .B(n2062), .Z(n4903) );
  ANDN U5557 ( .B(n4457), .A(n4458), .Z(n5350) );
  XNOR U5558 ( .A(n2200), .B(n5352), .Z(n4458) );
  XOR U5559 ( .A(n5353), .B(n2218), .Z(n4457) );
  IV U5560 ( .A(n3803), .Z(n2218) );
  XOR U5561 ( .A(n5354), .B(n4910), .Z(out[1321]) );
  XNOR U5562 ( .A(n5355), .B(n2069), .Z(n4910) );
  NOR U5563 ( .A(n4462), .B(n4461), .Z(n5354) );
  XNOR U5564 ( .A(n5356), .B(n3809), .Z(n4461) );
  XOR U5565 ( .A(n2207), .B(n5357), .Z(n4462) );
  XOR U5566 ( .A(n5358), .B(n4913), .Z(out[1320]) );
  XOR U5567 ( .A(n5359), .B(n2072), .Z(n4913) );
  ANDN U5568 ( .B(n4465), .A(n4467), .Z(n5358) );
  XOR U5569 ( .A(n2214), .B(n5360), .Z(n4467) );
  XOR U5570 ( .A(n5361), .B(n2238), .Z(n4465) );
  XOR U5571 ( .A(n5362), .B(n4056), .Z(out[131]) );
  XNOR U5572 ( .A(n5363), .B(n2062), .Z(n4056) );
  AND U5573 ( .A(n2374), .B(n2376), .Z(n5362) );
  XOR U5574 ( .A(n5364), .B(n2654), .Z(n2376) );
  IV U5575 ( .A(n5365), .Z(n2654) );
  XNOR U5576 ( .A(n5366), .B(n2340), .Z(n2374) );
  IV U5577 ( .A(n5367), .Z(n2340) );
  XOR U5578 ( .A(n5368), .B(n4916), .Z(out[1319]) );
  XNOR U5579 ( .A(n5369), .B(n2076), .Z(n4916) );
  NOR U5580 ( .A(n4470), .B(n4469), .Z(n5368) );
  XNOR U5581 ( .A(n5370), .B(n3822), .Z(n4469) );
  XNOR U5582 ( .A(n3343), .B(n5371), .Z(n4470) );
  XOR U5583 ( .A(n5372), .B(n4919), .Z(out[1318]) );
  XNOR U5584 ( .A(n5373), .B(n2079), .Z(n4919) );
  ANDN U5585 ( .B(n4475), .A(n4473), .Z(n5372) );
  XNOR U5586 ( .A(n5374), .B(n2252), .Z(n4473) );
  XOR U5587 ( .A(n2232), .B(n5375), .Z(n4475) );
  XOR U5588 ( .A(n5376), .B(n4922), .Z(out[1317]) );
  XOR U5589 ( .A(n5377), .B(n2082), .Z(n4922) );
  ANDN U5590 ( .B(n4479), .A(n4477), .Z(n5376) );
  XNOR U5591 ( .A(n5378), .B(n5379), .Z(n4477) );
  XNOR U5592 ( .A(n5380), .B(n5381), .Z(n4479) );
  XOR U5593 ( .A(n5382), .B(n4926), .Z(out[1316]) );
  XNOR U5594 ( .A(n5383), .B(n2085), .Z(n4926) );
  ANDN U5595 ( .B(n4481), .A(n4483), .Z(n5382) );
  XNOR U5596 ( .A(n5384), .B(n2249), .Z(n4483) );
  XNOR U5597 ( .A(n5385), .B(n3839), .Z(n4481) );
  XOR U5598 ( .A(n5386), .B(n4930), .Z(out[1315]) );
  XOR U5599 ( .A(n5387), .B(n2088), .Z(n4930) );
  NOR U5600 ( .A(n4487), .B(n4485), .Z(n5386) );
  XOR U5601 ( .A(n5388), .B(n3845), .Z(n4485) );
  XNOR U5602 ( .A(n5389), .B(n3363), .Z(n4487) );
  XOR U5603 ( .A(n5390), .B(n4933), .Z(out[1314]) );
  IV U5604 ( .A(n5145), .Z(n4933) );
  XNOR U5605 ( .A(n5391), .B(n2092), .Z(n5145) );
  NOR U5606 ( .A(n4491), .B(n4489), .Z(n5390) );
  XNOR U5607 ( .A(n5392), .B(n3849), .Z(n4489) );
  XNOR U5608 ( .A(n5393), .B(n2261), .Z(n4491) );
  XOR U5609 ( .A(n5394), .B(n4936), .Z(out[1313]) );
  XOR U5610 ( .A(n5395), .B(n5396), .Z(n4936) );
  ANDN U5611 ( .B(n4498), .A(n4499), .Z(n5394) );
  XOR U5612 ( .A(n5397), .B(n2268), .Z(n4499) );
  IV U5613 ( .A(n5398), .Z(n2268) );
  XOR U5614 ( .A(n5399), .B(n5400), .Z(n4498) );
  XNOR U5615 ( .A(n5401), .B(n4940), .Z(out[1312]) );
  XNOR U5616 ( .A(n3646), .B(n5402), .Z(n4940) );
  ANDN U5617 ( .B(n4502), .A(n4504), .Z(n5401) );
  XOR U5618 ( .A(n5403), .B(n2277), .Z(n4504) );
  XNOR U5619 ( .A(n5404), .B(n5138), .Z(n4502) );
  IV U5620 ( .A(n2294), .Z(n5138) );
  XOR U5621 ( .A(n5405), .B(n4947), .Z(out[1311]) );
  XOR U5622 ( .A(n5406), .B(n2105), .Z(n4947) );
  ANDN U5623 ( .B(n4511), .A(n4505), .Z(n5405) );
  XNOR U5624 ( .A(n5407), .B(n2305), .Z(n4505) );
  XOR U5625 ( .A(n5408), .B(n2284), .Z(n4511) );
  XOR U5626 ( .A(n5409), .B(n4950), .Z(out[1310]) );
  XOR U5627 ( .A(n2107), .B(n5410), .Z(n4950) );
  ANDN U5628 ( .B(n4514), .A(n4515), .Z(n5409) );
  XOR U5629 ( .A(n5412), .B(n2312), .Z(n4514) );
  IV U5630 ( .A(n5413), .Z(n2312) );
  XOR U5631 ( .A(n5414), .B(n4059), .Z(out[130]) );
  XOR U5632 ( .A(n5415), .B(n2069), .Z(n4059) );
  AND U5633 ( .A(n2448), .B(n2450), .Z(n5414) );
  XOR U5634 ( .A(n5416), .B(n3324), .Z(n2450) );
  IV U5635 ( .A(n2661), .Z(n3324) );
  XNOR U5636 ( .A(n5417), .B(n3565), .Z(n2448) );
  XNOR U5637 ( .A(n5418), .B(n4953), .Z(out[1309]) );
  XOR U5638 ( .A(n3664), .B(n5419), .Z(n4953) );
  ANDN U5639 ( .B(n4518), .A(n4519), .Z(n5418) );
  XOR U5640 ( .A(n5420), .B(n3140), .Z(n4519) );
  IV U5641 ( .A(n2298), .Z(n3140) );
  XOR U5642 ( .A(n5421), .B(n5229), .Z(n4518) );
  XOR U5643 ( .A(n5422), .B(n4956), .Z(out[1308]) );
  XNOR U5644 ( .A(n4284), .B(n5423), .Z(n4956) );
  AND U5645 ( .A(n4522), .B(n4524), .Z(n5422) );
  XNOR U5646 ( .A(n5424), .B(n2309), .Z(n4524) );
  XNOR U5647 ( .A(n5425), .B(n2326), .Z(n4522) );
  XNOR U5648 ( .A(n5426), .B(n4959), .Z(out[1307]) );
  XNOR U5649 ( .A(n2118), .B(n5427), .Z(n4959) );
  IV U5650 ( .A(n3672), .Z(n2118) );
  ANDN U5651 ( .B(n5163), .A(n4527), .Z(n5426) );
  XNOR U5652 ( .A(n5428), .B(n2316), .Z(n4527) );
  XOR U5653 ( .A(n5429), .B(n2333), .Z(n5163) );
  XOR U5654 ( .A(n5430), .B(n4962), .Z(out[1306]) );
  XOR U5655 ( .A(n2122), .B(n5431), .Z(n4962) );
  IV U5656 ( .A(n3679), .Z(n2122) );
  ANDN U5657 ( .B(n4532), .A(n4530), .Z(n5430) );
  XNOR U5658 ( .A(n5432), .B(n5367), .Z(n4530) );
  XNOR U5659 ( .A(n5433), .B(n5434), .Z(n4532) );
  XOR U5660 ( .A(n5435), .B(n4965), .Z(out[1305]) );
  XOR U5661 ( .A(n2126), .B(n5436), .Z(n4965) );
  NOR U5662 ( .A(n4535), .B(n4534), .Z(n5435) );
  XOR U5663 ( .A(n5437), .B(n3565), .Z(n4534) );
  XOR U5664 ( .A(n5438), .B(n2328), .Z(n4535) );
  XOR U5665 ( .A(n5439), .B(n4968), .Z(out[1304]) );
  XOR U5666 ( .A(n5440), .B(n2130), .Z(n4968) );
  NOR U5667 ( .A(n4539), .B(n4538), .Z(n5439) );
  XNOR U5668 ( .A(n5441), .B(n5442), .Z(n4538) );
  XOR U5669 ( .A(n5443), .B(n2335), .Z(n4539) );
  XOR U5670 ( .A(n5444), .B(n4971), .Z(out[1303]) );
  XOR U5671 ( .A(n5445), .B(n2133), .Z(n4971) );
  NOR U5672 ( .A(n4547), .B(n4546), .Z(n5444) );
  XNOR U5673 ( .A(n5446), .B(n3579), .Z(n4546) );
  XNOR U5674 ( .A(n5447), .B(n2344), .Z(n4547) );
  XOR U5675 ( .A(n5448), .B(n4974), .Z(out[1302]) );
  IV U5676 ( .A(n5179), .Z(n4974) );
  XNOR U5677 ( .A(n5449), .B(n2136), .Z(n5179) );
  ANDN U5678 ( .B(n4552), .A(n4550), .Z(n5448) );
  XNOR U5679 ( .A(n5450), .B(n5451), .Z(n4550) );
  XOR U5680 ( .A(n5452), .B(n2349), .Z(n4552) );
  XNOR U5681 ( .A(n5453), .B(n4981), .Z(out[1301]) );
  XNOR U5682 ( .A(n5454), .B(n2142), .Z(n4981) );
  AND U5683 ( .A(n4554), .B(n4556), .Z(n5453) );
  XOR U5684 ( .A(n5455), .B(n2356), .Z(n4556) );
  XOR U5685 ( .A(n5456), .B(n3588), .Z(n4554) );
  XOR U5686 ( .A(n5457), .B(n4985), .Z(out[1300]) );
  XOR U5687 ( .A(n5458), .B(n2146), .Z(n4985) );
  ANDN U5688 ( .B(n4558), .A(n4559), .Z(n5457) );
  XOR U5689 ( .A(n5459), .B(n2363), .Z(n4559) );
  XNOR U5690 ( .A(n5460), .B(n2386), .Z(n4558) );
  XOR U5691 ( .A(n5461), .B(n1957), .Z(out[12]) );
  XNOR U5692 ( .A(n5462), .B(n5292), .Z(n1957) );
  ANDN U5693 ( .B(n1958), .A(n4022), .Z(n5461) );
  XOR U5694 ( .A(n5463), .B(n1742), .Z(n4022) );
  XNOR U5695 ( .A(n2519), .B(n5464), .Z(n1958) );
  IV U5696 ( .A(n3468), .Z(n2519) );
  XOR U5697 ( .A(n5465), .B(n4061), .Z(out[129]) );
  XNOR U5698 ( .A(n5466), .B(n2072), .Z(n4061) );
  ANDN U5699 ( .B(n2522), .A(n2524), .Z(n5465) );
  XNOR U5700 ( .A(n5467), .B(n2668), .Z(n2524) );
  IV U5701 ( .A(n5468), .Z(n2668) );
  XNOR U5702 ( .A(n5469), .B(n2354), .Z(n2522) );
  IV U5703 ( .A(n5442), .Z(n2354) );
  XOR U5704 ( .A(n5470), .B(n4989), .Z(out[1299]) );
  XOR U5705 ( .A(n5471), .B(n2149), .Z(n4989) );
  ANDN U5706 ( .B(n4562), .A(n4563), .Z(n5470) );
  XOR U5707 ( .A(n5472), .B(n2372), .Z(n4563) );
  XNOR U5708 ( .A(n5473), .B(n2393), .Z(n4562) );
  XOR U5709 ( .A(n5474), .B(n4992), .Z(out[1298]) );
  XNOR U5710 ( .A(n5475), .B(n2152), .Z(n4992) );
  AND U5711 ( .A(n4566), .B(n4568), .Z(n5474) );
  XOR U5712 ( .A(n5476), .B(n2381), .Z(n4568) );
  XOR U5713 ( .A(n5477), .B(n2400), .Z(n4566) );
  XOR U5714 ( .A(n5478), .B(n4995), .Z(out[1297]) );
  XNOR U5715 ( .A(n5479), .B(n2155), .Z(n4995) );
  ANDN U5716 ( .B(n4570), .A(n4571), .Z(n5478) );
  XNOR U5717 ( .A(n5480), .B(n2390), .Z(n4571) );
  XOR U5718 ( .A(n5481), .B(n2407), .Z(n4570) );
  XOR U5719 ( .A(n5482), .B(n4998), .Z(out[1296]) );
  XOR U5720 ( .A(n5483), .B(n2159), .Z(n4998) );
  IV U5721 ( .A(n3728), .Z(n2159) );
  ANDN U5722 ( .B(n4574), .A(n4576), .Z(n5482) );
  XOR U5723 ( .A(n5484), .B(n2397), .Z(n4576) );
  XOR U5724 ( .A(n5485), .B(n2414), .Z(n4574) );
  XOR U5725 ( .A(n5486), .B(n5001), .Z(out[1295]) );
  XNOR U5726 ( .A(n5487), .B(n2163), .Z(n5001) );
  AND U5727 ( .A(n4581), .B(n4582), .Z(n5486) );
  XNOR U5728 ( .A(n5488), .B(n2421), .Z(n4582) );
  XOR U5729 ( .A(n5489), .B(n2402), .Z(n4581) );
  XOR U5730 ( .A(n5490), .B(n5005), .Z(out[1294]) );
  XOR U5731 ( .A(n5491), .B(n2166), .Z(n5005) );
  IV U5732 ( .A(n3737), .Z(n2166) );
  AND U5733 ( .A(n4584), .B(n4586), .Z(n5490) );
  XOR U5734 ( .A(n5492), .B(n2411), .Z(n4586) );
  XOR U5735 ( .A(n5493), .B(n2428), .Z(n4584) );
  XOR U5736 ( .A(n5494), .B(n5009), .Z(out[1293]) );
  XNOR U5737 ( .A(n5495), .B(n2169), .Z(n5009) );
  IV U5738 ( .A(n3743), .Z(n2169) );
  AND U5739 ( .A(n4593), .B(n4595), .Z(n5494) );
  XOR U5740 ( .A(n4336), .B(n5496), .Z(n4595) );
  XNOR U5741 ( .A(n5497), .B(n2435), .Z(n4593) );
  XOR U5742 ( .A(n5498), .B(n5012), .Z(out[1292]) );
  IV U5743 ( .A(n5208), .Z(n5012) );
  XOR U5744 ( .A(n5499), .B(n2172), .Z(n5208) );
  ANDN U5745 ( .B(n4599), .A(n4597), .Z(n5498) );
  XOR U5746 ( .A(n5500), .B(n3632), .Z(n4597) );
  XOR U5747 ( .A(n2424), .B(n5501), .Z(n4599) );
  XOR U5748 ( .A(n5502), .B(n5018), .Z(out[1291]) );
  XOR U5749 ( .A(n5503), .B(n2179), .Z(n5018) );
  IV U5750 ( .A(n3751), .Z(n2179) );
  AND U5751 ( .A(n4601), .B(n4603), .Z(n5502) );
  XOR U5752 ( .A(n5504), .B(n4346), .Z(n4603) );
  XNOR U5753 ( .A(n5505), .B(n2453), .Z(n4601) );
  XOR U5754 ( .A(n5506), .B(n5021), .Z(out[1290]) );
  XNOR U5755 ( .A(n5507), .B(n2182), .Z(n5021) );
  IV U5756 ( .A(n3756), .Z(n2182) );
  ANDN U5757 ( .B(n4607), .A(n4605), .Z(n5506) );
  XOR U5758 ( .A(n5508), .B(n2460), .Z(n4605) );
  XNOR U5759 ( .A(n5509), .B(n2439), .Z(n4607) );
  IV U5760 ( .A(n3211), .Z(n2439) );
  XOR U5761 ( .A(n5510), .B(n4064), .Z(out[128]) );
  XNOR U5762 ( .A(n5511), .B(n2076), .Z(n4064) );
  AND U5763 ( .A(n2598), .B(n2596), .Z(n5510) );
  XNOR U5764 ( .A(n5512), .B(n3579), .Z(n2596) );
  XOR U5765 ( .A(n5513), .B(n5024), .Z(out[1289]) );
  XNOR U5766 ( .A(n5514), .B(n2185), .Z(n5024) );
  NOR U5767 ( .A(n4610), .B(n4609), .Z(n5513) );
  XOR U5768 ( .A(n5515), .B(n3649), .Z(n4609) );
  IV U5769 ( .A(n2467), .Z(n3649) );
  XNOR U5770 ( .A(n5516), .B(n2446), .Z(n4610) );
  IV U5771 ( .A(n3215), .Z(n2446) );
  XOR U5772 ( .A(n5517), .B(n5028), .Z(out[1288]) );
  XOR U5773 ( .A(n5518), .B(n2188), .Z(n5028) );
  ANDN U5774 ( .B(n4613), .A(n4614), .Z(n5517) );
  XOR U5775 ( .A(n5519), .B(n2455), .Z(n4614) );
  XNOR U5776 ( .A(n5520), .B(n3654), .Z(n4613) );
  XOR U5777 ( .A(n5521), .B(n5031), .Z(out[1287]) );
  XOR U5778 ( .A(n5522), .B(n2191), .Z(n5031) );
  IV U5779 ( .A(n3771), .Z(n2191) );
  NOR U5780 ( .A(n4618), .B(n4617), .Z(n5521) );
  XOR U5781 ( .A(n5523), .B(n2481), .Z(n4617) );
  XNOR U5782 ( .A(n5524), .B(n2464), .Z(n4618) );
  IV U5783 ( .A(n3222), .Z(n2464) );
  XOR U5784 ( .A(n5525), .B(n5034), .Z(out[1286]) );
  XNOR U5785 ( .A(n5526), .B(n4357), .Z(n5034) );
  ANDN U5786 ( .B(n4623), .A(n4621), .Z(n5525) );
  XOR U5787 ( .A(n5527), .B(n2488), .Z(n4621) );
  XOR U5788 ( .A(n5528), .B(n2471), .Z(n4623) );
  XOR U5789 ( .A(n5529), .B(n5037), .Z(out[1285]) );
  XOR U5790 ( .A(n5530), .B(n1969), .Z(n5037) );
  ANDN U5791 ( .B(n4625), .A(n4626), .Z(n5529) );
  XOR U5792 ( .A(n5531), .B(n2476), .Z(n4626) );
  XOR U5793 ( .A(n5532), .B(n2495), .Z(n4625) );
  XOR U5794 ( .A(n5533), .B(n5042), .Z(out[1284]) );
  XOR U5795 ( .A(n5534), .B(n1972), .Z(n5042) );
  ANDN U5796 ( .B(n4631), .A(n4629), .Z(n5533) );
  XNOR U5797 ( .A(n5535), .B(n2502), .Z(n4629) );
  XOR U5798 ( .A(n5536), .B(n2483), .Z(n4631) );
  XOR U5799 ( .A(n5537), .B(n5045), .Z(out[1283]) );
  XNOR U5800 ( .A(n5538), .B(n4494), .Z(n5045) );
  NOR U5801 ( .A(n4641), .B(n4636), .Z(n5537) );
  XNOR U5802 ( .A(n5539), .B(n3682), .Z(n4636) );
  IV U5803 ( .A(n2509), .Z(n3682) );
  XOR U5804 ( .A(n5540), .B(n2490), .Z(n4641) );
  XOR U5805 ( .A(n5541), .B(n5048), .Z(out[1282]) );
  XOR U5806 ( .A(n5542), .B(n1978), .Z(n5048) );
  NOR U5807 ( .A(n4645), .B(n4644), .Z(n5541) );
  XOR U5808 ( .A(n5543), .B(n3687), .Z(n4644) );
  XNOR U5809 ( .A(n5544), .B(n4676), .Z(n4645) );
  XOR U5810 ( .A(n5545), .B(n5055), .Z(out[1281]) );
  XOR U5811 ( .A(n5546), .B(n1981), .Z(n5055) );
  AND U5812 ( .A(n4652), .B(n4647), .Z(n5545) );
  XOR U5813 ( .A(n5547), .B(n2527), .Z(n4647) );
  XNOR U5814 ( .A(n5548), .B(n4701), .Z(n4652) );
  XOR U5815 ( .A(n5549), .B(n5059), .Z(out[1280]) );
  XNOR U5816 ( .A(n5550), .B(n1984), .Z(n5059) );
  ANDN U5817 ( .B(n4653), .A(n4657), .Z(n5549) );
  XNOR U5818 ( .A(n5551), .B(n4728), .Z(n4657) );
  XOR U5819 ( .A(n5552), .B(n2534), .Z(n4653) );
  XOR U5820 ( .A(n5553), .B(n4068), .Z(out[127]) );
  XOR U5821 ( .A(n5554), .B(n2368), .Z(n4068) );
  IV U5822 ( .A(n5451), .Z(n2368) );
  NOR U5823 ( .A(n2672), .B(n2670), .Z(n5553) );
  XOR U5824 ( .A(n5555), .B(n5556), .Z(n2670) );
  XOR U5825 ( .A(n5557), .B(n2617), .Z(n2672) );
  XOR U5826 ( .A(n5558), .B(n5559), .Z(out[1279]) );
  XOR U5827 ( .A(n5562), .B(n5563), .Z(out[1278]) );
  ANDN U5828 ( .B(n5564), .A(n5565), .Z(n5562) );
  XOR U5829 ( .A(n5566), .B(n5567), .Z(out[1277]) );
  XOR U5830 ( .A(n5570), .B(n5571), .Z(out[1276]) );
  AND U5831 ( .A(n5572), .B(n5573), .Z(n5570) );
  XOR U5832 ( .A(n5574), .B(n5575), .Z(out[1275]) );
  AND U5833 ( .A(n5576), .B(n5577), .Z(n5574) );
  XOR U5834 ( .A(n5578), .B(n5579), .Z(out[1274]) );
  AND U5835 ( .A(n5580), .B(n5581), .Z(n5578) );
  XOR U5836 ( .A(n5582), .B(n5583), .Z(out[1273]) );
  ANDN U5837 ( .B(n5584), .A(n5585), .Z(n5582) );
  XOR U5838 ( .A(n5586), .B(n5587), .Z(out[1272]) );
  ANDN U5839 ( .B(n5588), .A(n5589), .Z(n5586) );
  XOR U5840 ( .A(n5590), .B(n5591), .Z(out[1271]) );
  ANDN U5841 ( .B(n5592), .A(n5593), .Z(n5590) );
  XOR U5842 ( .A(n5594), .B(n5595), .Z(out[1270]) );
  ANDN U5843 ( .B(n5596), .A(n5597), .Z(n5594) );
  XOR U5844 ( .A(n5598), .B(n4071), .Z(out[126]) );
  XNOR U5845 ( .A(n5599), .B(n3588), .Z(n4071) );
  ANDN U5846 ( .B(n2714), .A(n2716), .Z(n5598) );
  XOR U5847 ( .A(n5600), .B(n2624), .Z(n2716) );
  XNOR U5848 ( .A(n2214), .B(n5601), .Z(n2714) );
  IV U5849 ( .A(n3339), .Z(n2214) );
  XOR U5850 ( .A(n5602), .B(n5603), .Z(out[1269]) );
  ANDN U5851 ( .B(n5604), .A(n5605), .Z(n5602) );
  XOR U5852 ( .A(n5606), .B(n5607), .Z(out[1268]) );
  ANDN U5853 ( .B(n5608), .A(n5609), .Z(n5606) );
  XNOR U5854 ( .A(n5610), .B(n5611), .Z(out[1267]) );
  ANDN U5855 ( .B(n5612), .A(n5613), .Z(n5610) );
  XOR U5856 ( .A(n5614), .B(n5615), .Z(out[1266]) );
  ANDN U5857 ( .B(n5616), .A(n5617), .Z(n5614) );
  XNOR U5858 ( .A(n5618), .B(n5619), .Z(out[1265]) );
  XOR U5859 ( .A(n5622), .B(n5623), .Z(out[1264]) );
  ANDN U5860 ( .B(n5624), .A(n5625), .Z(n5622) );
  XOR U5861 ( .A(n5626), .B(n5627), .Z(out[1263]) );
  AND U5862 ( .A(n5628), .B(n5629), .Z(n5626) );
  XNOR U5863 ( .A(n5630), .B(n5631), .Z(out[1262]) );
  AND U5864 ( .A(n5632), .B(n5633), .Z(n5630) );
  XOR U5865 ( .A(n5634), .B(n5635), .Z(out[1261]) );
  ANDN U5866 ( .B(n5636), .A(n5637), .Z(n5634) );
  XOR U5867 ( .A(n5638), .B(n5639), .Z(out[1260]) );
  ANDN U5868 ( .B(n5640), .A(n5641), .Z(n5638) );
  XOR U5869 ( .A(n5642), .B(n4074), .Z(out[125]) );
  XOR U5870 ( .A(n5643), .B(n2386), .Z(n4074) );
  IV U5871 ( .A(n5644), .Z(n2386) );
  NOR U5872 ( .A(n2760), .B(n2758), .Z(n5642) );
  XOR U5873 ( .A(n3343), .B(n5645), .Z(n2758) );
  IV U5874 ( .A(n2221), .Z(n3343) );
  XOR U5875 ( .A(n5646), .B(n2631), .Z(n2760) );
  XOR U5876 ( .A(n5647), .B(n5648), .Z(out[1259]) );
  ANDN U5877 ( .B(n5649), .A(n5650), .Z(n5647) );
  XOR U5878 ( .A(n5651), .B(n5652), .Z(out[1258]) );
  XNOR U5879 ( .A(n5655), .B(n5656), .Z(out[1257]) );
  XOR U5880 ( .A(n5659), .B(n5660), .Z(out[1256]) );
  ANDN U5881 ( .B(n5661), .A(n5662), .Z(n5659) );
  XNOR U5882 ( .A(n5663), .B(n1044), .Z(out[1255]) );
  ANDN U5883 ( .B(n5664), .A(n1043), .Z(n5663) );
  XOR U5884 ( .A(n5665), .B(n1048), .Z(out[1254]) );
  XOR U5885 ( .A(n5667), .B(n1052), .Z(out[1253]) );
  ANDN U5886 ( .B(n5668), .A(n1051), .Z(n5667) );
  XNOR U5887 ( .A(n5669), .B(n1055), .Z(out[1252]) );
  AND U5888 ( .A(n5670), .B(n1056), .Z(n5669) );
  XOR U5889 ( .A(n5671), .B(n1060), .Z(out[1251]) );
  ANDN U5890 ( .B(n5672), .A(n1059), .Z(n5671) );
  XNOR U5891 ( .A(n5673), .B(n1064), .Z(out[1250]) );
  ANDN U5892 ( .B(n5674), .A(n1063), .Z(n5673) );
  XOR U5893 ( .A(n5675), .B(n4077), .Z(out[124]) );
  XNOR U5894 ( .A(n5676), .B(n3598), .Z(n4077) );
  AND U5895 ( .A(n2804), .B(n4269), .Z(n5675) );
  XOR U5896 ( .A(n5677), .B(n5678), .Z(n4269) );
  XNOR U5897 ( .A(n5679), .B(n2638), .Z(n2804) );
  XNOR U5898 ( .A(n5680), .B(n1068), .Z(out[1249]) );
  ANDN U5899 ( .B(n5681), .A(n1067), .Z(n5680) );
  XOR U5900 ( .A(n5682), .B(n1072), .Z(out[1248]) );
  ANDN U5901 ( .B(n5683), .A(n1071), .Z(n5682) );
  XNOR U5902 ( .A(n5684), .B(n1076), .Z(out[1247]) );
  ANDN U5903 ( .B(n5685), .A(n1075), .Z(n5684) );
  XNOR U5904 ( .A(n5686), .B(n1080), .Z(out[1246]) );
  ANDN U5905 ( .B(n5687), .A(n1079), .Z(n5686) );
  XOR U5906 ( .A(n5688), .B(n1088), .Z(out[1245]) );
  ANDN U5907 ( .B(n5689), .A(n1087), .Z(n5688) );
  XOR U5908 ( .A(n5690), .B(n1092), .Z(out[1244]) );
  ANDN U5909 ( .B(n5691), .A(n1091), .Z(n5690) );
  XNOR U5910 ( .A(n5692), .B(n1096), .Z(out[1243]) );
  ANDN U5911 ( .B(n5693), .A(n1095), .Z(n5692) );
  XOR U5912 ( .A(n5694), .B(n1099), .Z(out[1242]) );
  AND U5913 ( .A(n1100), .B(n5695), .Z(n5694) );
  XOR U5914 ( .A(n5696), .B(n1104), .Z(out[1241]) );
  ANDN U5915 ( .B(n5697), .A(n1103), .Z(n5696) );
  XNOR U5916 ( .A(n5698), .B(n1107), .Z(out[1240]) );
  AND U5917 ( .A(n5699), .B(n5700), .Z(n5698) );
  XOR U5918 ( .A(n5701), .B(n4081), .Z(out[123]) );
  XNOR U5919 ( .A(n5702), .B(n2400), .Z(n4081) );
  ANDN U5920 ( .B(n2848), .A(n2849), .Z(n5701) );
  XNOR U5921 ( .A(n5703), .B(n2645), .Z(n2849) );
  XOR U5922 ( .A(n5704), .B(n5381), .Z(n2848) );
  IV U5923 ( .A(n2242), .Z(n5381) );
  XNOR U5924 ( .A(n5705), .B(n1112), .Z(out[1239]) );
  ANDN U5925 ( .B(n5706), .A(n1111), .Z(n5705) );
  XOR U5926 ( .A(n5707), .B(n1116), .Z(out[1238]) );
  ANDN U5927 ( .B(n5708), .A(n1115), .Z(n5707) );
  XOR U5928 ( .A(n5709), .B(n1119), .Z(out[1237]) );
  AND U5929 ( .A(n1120), .B(n5710), .Z(n5709) );
  XNOR U5930 ( .A(n5711), .B(n1124), .Z(out[1236]) );
  ANDN U5931 ( .B(n5712), .A(n1123), .Z(n5711) );
  XNOR U5932 ( .A(n5713), .B(n1131), .Z(out[1235]) );
  XOR U5933 ( .A(n5715), .B(n1135), .Z(out[1234]) );
  AND U5934 ( .A(n1136), .B(n5716), .Z(n5715) );
  XOR U5935 ( .A(n5717), .B(n1140), .Z(out[1233]) );
  ANDN U5936 ( .B(n5718), .A(n1139), .Z(n5717) );
  XOR U5937 ( .A(n5719), .B(n1144), .Z(out[1232]) );
  AND U5938 ( .A(n5720), .B(n1143), .Z(n5719) );
  IV U5939 ( .A(n5721), .Z(n1143) );
  XOR U5940 ( .A(n5722), .B(n1147), .Z(out[1231]) );
  AND U5941 ( .A(n1148), .B(n5723), .Z(n5722) );
  XOR U5942 ( .A(n5724), .B(n1151), .Z(out[1230]) );
  AND U5943 ( .A(n1152), .B(n5725), .Z(n5724) );
  XOR U5944 ( .A(n5726), .B(n4084), .Z(out[122]) );
  XNOR U5945 ( .A(n5727), .B(n2407), .Z(n4084) );
  NOR U5946 ( .A(n2894), .B(n2892), .Z(n5726) );
  XNOR U5947 ( .A(n5728), .B(n2249), .Z(n2892) );
  IV U5948 ( .A(n5729), .Z(n2249) );
  XNOR U5949 ( .A(n5730), .B(n2652), .Z(n2894) );
  XNOR U5950 ( .A(n5731), .B(n1156), .Z(out[1229]) );
  ANDN U5951 ( .B(n5732), .A(n1155), .Z(n5731) );
  XNOR U5952 ( .A(n5733), .B(n1160), .Z(out[1228]) );
  ANDN U5953 ( .B(n5734), .A(n1159), .Z(n5733) );
  XNOR U5954 ( .A(n5735), .B(n1164), .Z(out[1227]) );
  ANDN U5955 ( .B(n5736), .A(n1163), .Z(n5735) );
  XNOR U5956 ( .A(n5737), .B(n1168), .Z(out[1226]) );
  ANDN U5957 ( .B(n5738), .A(n1167), .Z(n5737) );
  XOR U5958 ( .A(n5739), .B(n1176), .Z(out[1225]) );
  XNOR U5959 ( .A(n5741), .B(n1179), .Z(out[1224]) );
  AND U5960 ( .A(n1180), .B(n5742), .Z(n5741) );
  XNOR U5961 ( .A(n5743), .B(n1183), .Z(out[1223]) );
  AND U5962 ( .A(n5744), .B(n5745), .Z(n5743) );
  XNOR U5963 ( .A(n5746), .B(n1188), .Z(out[1222]) );
  ANDN U5964 ( .B(n5747), .A(n1187), .Z(n5746) );
  XOR U5965 ( .A(n5748), .B(n1192), .Z(out[1221]) );
  AND U5966 ( .A(n5749), .B(n5750), .Z(n5748) );
  XNOR U5967 ( .A(n5751), .B(n1195), .Z(out[1220]) );
  XOR U5968 ( .A(n5753), .B(n4090), .Z(out[121]) );
  XNOR U5969 ( .A(n5754), .B(n2414), .Z(n4090) );
  AND U5970 ( .A(n2938), .B(n4276), .Z(n5753) );
  XOR U5971 ( .A(n5755), .B(n3363), .Z(n4276) );
  IV U5972 ( .A(n2256), .Z(n3363) );
  XNOR U5973 ( .A(n5756), .B(n2659), .Z(n2938) );
  XOR U5974 ( .A(n5757), .B(n1200), .Z(out[1219]) );
  AND U5975 ( .A(n1199), .B(n5758), .Z(n5757) );
  XOR U5976 ( .A(n5759), .B(n1204), .Z(out[1218]) );
  AND U5977 ( .A(n5760), .B(n5761), .Z(n5759) );
  XOR U5978 ( .A(n5762), .B(n1207), .Z(out[1217]) );
  AND U5979 ( .A(n5763), .B(n1208), .Z(n5762) );
  XNOR U5980 ( .A(n5764), .B(n1212), .Z(out[1216]) );
  ANDN U5981 ( .B(n5765), .A(n1211), .Z(n5764) );
  XOR U5982 ( .A(n5766), .B(n5561), .Z(out[1215]) );
  ANDN U5983 ( .B(n5767), .A(n5560), .Z(n5766) );
  XOR U5984 ( .A(n5768), .B(n5565), .Z(out[1214]) );
  ANDN U5985 ( .B(n5769), .A(n5564), .Z(n5768) );
  XOR U5986 ( .A(n5770), .B(n5569), .Z(out[1213]) );
  ANDN U5987 ( .B(n5771), .A(n5568), .Z(n5770) );
  XNOR U5988 ( .A(n5772), .B(n5573), .Z(out[1212]) );
  ANDN U5989 ( .B(n5773), .A(n5572), .Z(n5772) );
  XNOR U5990 ( .A(n5774), .B(n5577), .Z(out[1211]) );
  ANDN U5991 ( .B(n5775), .A(n5576), .Z(n5774) );
  XNOR U5992 ( .A(n5776), .B(n5581), .Z(out[1210]) );
  ANDN U5993 ( .B(n5777), .A(n5580), .Z(n5776) );
  XOR U5994 ( .A(n5778), .B(n4093), .Z(out[120]) );
  XOR U5995 ( .A(n5779), .B(n2421), .Z(n4093) );
  AND U5996 ( .A(n2968), .B(n2970), .Z(n5778) );
  XNOR U5997 ( .A(n5780), .B(n2666), .Z(n2970) );
  XNOR U5998 ( .A(n5781), .B(n2261), .Z(n2968) );
  IV U5999 ( .A(n3367), .Z(n2261) );
  XOR U6000 ( .A(n5782), .B(n5585), .Z(out[1209]) );
  ANDN U6001 ( .B(n5783), .A(n5584), .Z(n5782) );
  XOR U6002 ( .A(n5784), .B(n5589), .Z(out[1208]) );
  NOR U6003 ( .A(n5785), .B(n5588), .Z(n5784) );
  XOR U6004 ( .A(n5786), .B(n5593), .Z(out[1207]) );
  ANDN U6005 ( .B(n5787), .A(n5592), .Z(n5786) );
  XOR U6006 ( .A(n5788), .B(n5597), .Z(out[1206]) );
  ANDN U6007 ( .B(n5789), .A(n5596), .Z(n5788) );
  XOR U6008 ( .A(n5790), .B(n5605), .Z(out[1205]) );
  ANDN U6009 ( .B(n5791), .A(n5604), .Z(n5790) );
  XOR U6010 ( .A(n5792), .B(n5609), .Z(out[1204]) );
  ANDN U6011 ( .B(n5793), .A(n5608), .Z(n5792) );
  XOR U6012 ( .A(n5794), .B(n5613), .Z(out[1203]) );
  ANDN U6013 ( .B(n5795), .A(n5612), .Z(n5794) );
  XOR U6014 ( .A(n5796), .B(n5617), .Z(out[1202]) );
  AND U6015 ( .A(n5797), .B(n5798), .Z(n5796) );
  XOR U6016 ( .A(n5799), .B(n5621), .Z(out[1201]) );
  ANDN U6017 ( .B(n5800), .A(n5620), .Z(n5799) );
  XOR U6018 ( .A(n5801), .B(n5625), .Z(out[1200]) );
  ANDN U6019 ( .B(n5802), .A(n5624), .Z(n5801) );
  XOR U6020 ( .A(n5803), .B(n1994), .Z(out[11]) );
  XNOR U6021 ( .A(n5804), .B(n2594), .Z(n1994) );
  IV U6022 ( .A(n5298), .Z(n2594) );
  ANDN U6023 ( .B(n1993), .A(n4026), .Z(n5803) );
  XOR U6024 ( .A(n5805), .B(n1747), .Z(n4026) );
  XNOR U6025 ( .A(n2528), .B(n5806), .Z(n1993) );
  IV U6026 ( .A(n4854), .Z(n2528) );
  XNOR U6027 ( .A(n5807), .B(n4096), .Z(out[119]) );
  XOR U6028 ( .A(n5808), .B(n2428), .Z(n4096) );
  ANDN U6029 ( .B(n2995), .A(n2997), .Z(n5807) );
  XOR U6030 ( .A(n5809), .B(n2199), .Z(n2997) );
  IV U6031 ( .A(n4925), .Z(n2199) );
  XNOR U6032 ( .A(n5810), .B(n5398), .Z(n2995) );
  XNOR U6033 ( .A(n5811), .B(n5628), .Z(out[1199]) );
  AND U6034 ( .A(n5812), .B(n5813), .Z(n5811) );
  XNOR U6035 ( .A(n5814), .B(n5632), .Z(out[1198]) );
  AND U6036 ( .A(n5815), .B(n5816), .Z(n5814) );
  XOR U6037 ( .A(n5817), .B(n5637), .Z(out[1197]) );
  ANDN U6038 ( .B(n5818), .A(n5636), .Z(n5817) );
  XOR U6039 ( .A(n5819), .B(n5641), .Z(out[1196]) );
  ANDN U6040 ( .B(n5820), .A(n5640), .Z(n5819) );
  XNOR U6041 ( .A(n5821), .B(n5649), .Z(out[1195]) );
  XOR U6042 ( .A(n5823), .B(n5654), .Z(out[1194]) );
  NOR U6043 ( .A(n5824), .B(n5653), .Z(n5823) );
  XOR U6044 ( .A(n5825), .B(n5658), .Z(out[1193]) );
  ANDN U6045 ( .B(n5826), .A(n5657), .Z(n5825) );
  XNOR U6046 ( .A(n5827), .B(n5661), .Z(out[1192]) );
  AND U6047 ( .A(n5662), .B(n5828), .Z(n5827) );
  XOR U6048 ( .A(n5829), .B(n1043), .Z(out[1191]) );
  XNOR U6049 ( .A(n2094), .B(n5830), .Z(n1043) );
  IV U6050 ( .A(n5395), .Z(n2094) );
  XOR U6051 ( .A(n5831), .B(n5832), .Z(n5395) );
  ANDN U6052 ( .B(n5833), .A(n5664), .Z(n5829) );
  XOR U6053 ( .A(n5834), .B(n1047), .Z(out[1190]) );
  XOR U6054 ( .A(n3646), .B(n5835), .Z(n1047) );
  IV U6055 ( .A(n2097), .Z(n3646) );
  XOR U6056 ( .A(n5836), .B(n5837), .Z(n2097) );
  ANDN U6057 ( .B(n5838), .A(n5666), .Z(n5834) );
  XOR U6058 ( .A(n5839), .B(n4100), .Z(out[118]) );
  XOR U6059 ( .A(n5840), .B(n2435), .Z(n4100) );
  IV U6060 ( .A(n5841), .Z(n2435) );
  AND U6061 ( .A(n3022), .B(n3024), .Z(n5839) );
  XOR U6062 ( .A(n5842), .B(n2206), .Z(n3024) );
  IV U6063 ( .A(n4929), .Z(n2206) );
  XNOR U6064 ( .A(n5843), .B(n2277), .Z(n3022) );
  XOR U6065 ( .A(n5844), .B(n1051), .Z(out[1189]) );
  XOR U6066 ( .A(n5845), .B(n2105), .Z(n1051) );
  XOR U6067 ( .A(n5846), .B(n5847), .Z(n2105) );
  ANDN U6068 ( .B(n5848), .A(n5668), .Z(n5844) );
  XNOR U6069 ( .A(n5849), .B(n1056), .Z(out[1188]) );
  XOR U6070 ( .A(n5851), .B(n5852), .Z(n2107) );
  ANDN U6071 ( .B(n5853), .A(n5670), .Z(n5849) );
  XOR U6072 ( .A(n5854), .B(n1059), .Z(out[1187]) );
  XNOR U6073 ( .A(n2111), .B(n5855), .Z(n1059) );
  IV U6074 ( .A(n3664), .Z(n2111) );
  XOR U6075 ( .A(n5856), .B(n5857), .Z(n3664) );
  NOR U6076 ( .A(n5858), .B(n5672), .Z(n5854) );
  XOR U6077 ( .A(n5859), .B(n1063), .Z(out[1186]) );
  XNOR U6078 ( .A(n2114), .B(n5860), .Z(n1063) );
  IV U6079 ( .A(n4284), .Z(n2114) );
  XOR U6080 ( .A(n5861), .B(n5862), .Z(n4284) );
  XOR U6081 ( .A(n5864), .B(n1067), .Z(out[1185]) );
  XNOR U6082 ( .A(n3672), .B(n5865), .Z(n1067) );
  XOR U6083 ( .A(n5866), .B(n5867), .Z(n3672) );
  NOR U6084 ( .A(n5868), .B(n5681), .Z(n5864) );
  XOR U6085 ( .A(n5869), .B(n1071), .Z(out[1184]) );
  XNOR U6086 ( .A(n3679), .B(n5870), .Z(n1071) );
  XOR U6087 ( .A(n5871), .B(n5872), .Z(n3679) );
  ANDN U6088 ( .B(n5873), .A(n5683), .Z(n5869) );
  XOR U6089 ( .A(n5874), .B(n1075), .Z(out[1183]) );
  XNOR U6090 ( .A(n2126), .B(n5875), .Z(n1075) );
  XOR U6091 ( .A(n5876), .B(n5877), .Z(n2126) );
  ANDN U6092 ( .B(n5878), .A(n5685), .Z(n5874) );
  XOR U6093 ( .A(n5879), .B(n1079), .Z(out[1182]) );
  XOR U6094 ( .A(n5880), .B(n2130), .Z(n1079) );
  XNOR U6095 ( .A(n5881), .B(n5882), .Z(n2130) );
  ANDN U6096 ( .B(n5883), .A(n5687), .Z(n5879) );
  XOR U6097 ( .A(n5884), .B(n1087), .Z(out[1181]) );
  XOR U6098 ( .A(n5885), .B(n2133), .Z(n1087) );
  XNOR U6099 ( .A(n5886), .B(n5887), .Z(n2133) );
  ANDN U6100 ( .B(n5888), .A(n5689), .Z(n5884) );
  XOR U6101 ( .A(n5889), .B(n1091), .Z(out[1180]) );
  XOR U6102 ( .A(n5890), .B(n2136), .Z(n1091) );
  XNOR U6103 ( .A(n5891), .B(n5892), .Z(n2136) );
  ANDN U6104 ( .B(n5893), .A(n5691), .Z(n5889) );
  XOR U6105 ( .A(n5894), .B(n4104), .Z(out[117]) );
  XNOR U6106 ( .A(n5895), .B(n2442), .Z(n4104) );
  AND U6107 ( .A(n3048), .B(n3050), .Z(n5894) );
  XOR U6108 ( .A(n5896), .B(n2213), .Z(n3050) );
  IV U6109 ( .A(n5897), .Z(n2213) );
  XNOR U6110 ( .A(n5898), .B(n3132), .Z(n3048) );
  IV U6111 ( .A(n2284), .Z(n3132) );
  XOR U6112 ( .A(n5899), .B(n1095), .Z(out[1179]) );
  XOR U6113 ( .A(n5900), .B(n2142), .Z(n1095) );
  XNOR U6114 ( .A(n5901), .B(n5902), .Z(n2142) );
  ANDN U6115 ( .B(n5903), .A(n5693), .Z(n5899) );
  XNOR U6116 ( .A(n5904), .B(n1100), .Z(out[1178]) );
  XNOR U6117 ( .A(n5905), .B(n2146), .Z(n1100) );
  XNOR U6118 ( .A(n5906), .B(n5907), .Z(n2146) );
  ANDN U6119 ( .B(n5908), .A(n5695), .Z(n5904) );
  XOR U6120 ( .A(n5909), .B(n1103), .Z(out[1177]) );
  XOR U6121 ( .A(n5910), .B(n2149), .Z(n1103) );
  XNOR U6122 ( .A(n5911), .B(n5912), .Z(n2149) );
  NOR U6123 ( .A(n5913), .B(n5697), .Z(n5909) );
  XOR U6124 ( .A(n5914), .B(n1108), .Z(out[1176]) );
  IV U6125 ( .A(n5700), .Z(n1108) );
  XOR U6126 ( .A(n5915), .B(n2152), .Z(n5700) );
  XNOR U6127 ( .A(n5916), .B(n5917), .Z(n2152) );
  ANDN U6128 ( .B(n5918), .A(n5699), .Z(n5914) );
  XOR U6129 ( .A(n5919), .B(n1111), .Z(out[1175]) );
  XNOR U6130 ( .A(n5920), .B(n2155), .Z(n1111) );
  XNOR U6131 ( .A(n5921), .B(n5922), .Z(n2155) );
  ANDN U6132 ( .B(n5923), .A(n5706), .Z(n5919) );
  XOR U6133 ( .A(n5924), .B(n1115), .Z(out[1174]) );
  XNOR U6134 ( .A(n5925), .B(n3728), .Z(n1115) );
  XNOR U6135 ( .A(n5926), .B(n5927), .Z(n3728) );
  ANDN U6136 ( .B(n5928), .A(n5708), .Z(n5924) );
  XNOR U6137 ( .A(n5929), .B(n1120), .Z(out[1173]) );
  XOR U6138 ( .A(n5930), .B(n2163), .Z(n1120) );
  XNOR U6139 ( .A(n5931), .B(n5932), .Z(n2163) );
  ANDN U6140 ( .B(n5933), .A(n5710), .Z(n5929) );
  XOR U6141 ( .A(n5934), .B(n1123), .Z(out[1172]) );
  XNOR U6142 ( .A(n5935), .B(n3737), .Z(n1123) );
  XNOR U6143 ( .A(n5936), .B(n5937), .Z(n3737) );
  ANDN U6144 ( .B(n5938), .A(n5712), .Z(n5934) );
  XOR U6145 ( .A(n5939), .B(n1132), .Z(out[1171]) );
  XOR U6146 ( .A(n5940), .B(n3743), .Z(n1132) );
  ANDN U6147 ( .B(n5943), .A(n5714), .Z(n5939) );
  XNOR U6148 ( .A(n5944), .B(n1136), .Z(out[1170]) );
  XOR U6149 ( .A(n5945), .B(n2172), .Z(n1136) );
  XNOR U6150 ( .A(n5946), .B(n5947), .Z(n2172) );
  ANDN U6151 ( .B(n5948), .A(n5716), .Z(n5944) );
  XNOR U6152 ( .A(n5949), .B(n4107), .Z(out[116]) );
  XNOR U6153 ( .A(n5950), .B(n2453), .Z(n4107) );
  ANDN U6154 ( .B(n3074), .A(n3075), .Z(n5949) );
  XNOR U6155 ( .A(n5951), .B(n2220), .Z(n3075) );
  IV U6156 ( .A(n5952), .Z(n2220) );
  XNOR U6157 ( .A(n5953), .B(n2291), .Z(n3074) );
  XOR U6158 ( .A(n5954), .B(n1139), .Z(out[1169]) );
  XNOR U6159 ( .A(n5955), .B(n3751), .Z(n1139) );
  XNOR U6160 ( .A(n5956), .B(n5957), .Z(n3751) );
  ANDN U6161 ( .B(n5958), .A(n5718), .Z(n5954) );
  XOR U6162 ( .A(n5959), .B(n5721), .Z(out[1168]) );
  XOR U6163 ( .A(n5960), .B(n3756), .Z(n5721) );
  XNOR U6164 ( .A(n5961), .B(n5962), .Z(n3756) );
  NOR U6165 ( .A(n5720), .B(n5963), .Z(n5959) );
  XNOR U6166 ( .A(n5964), .B(n1148), .Z(out[1167]) );
  XOR U6167 ( .A(n5965), .B(n2185), .Z(n1148) );
  XNOR U6168 ( .A(n5966), .B(n5967), .Z(n2185) );
  ANDN U6169 ( .B(n5968), .A(n5723), .Z(n5964) );
  XNOR U6170 ( .A(n5969), .B(n1152), .Z(out[1166]) );
  XOR U6171 ( .A(n5970), .B(n2188), .Z(n1152) );
  XNOR U6172 ( .A(n5971), .B(n5972), .Z(n2188) );
  NOR U6173 ( .A(n5973), .B(n5725), .Z(n5969) );
  XOR U6174 ( .A(n5974), .B(n1155), .Z(out[1165]) );
  XNOR U6175 ( .A(n5975), .B(n3771), .Z(n1155) );
  XNOR U6176 ( .A(n5976), .B(n5977), .Z(n3771) );
  ANDN U6177 ( .B(n5978), .A(n5732), .Z(n5974) );
  XOR U6178 ( .A(n5979), .B(n1159), .Z(out[1164]) );
  XOR U6179 ( .A(n5980), .B(n2194), .Z(n1159) );
  IV U6180 ( .A(n4357), .Z(n2194) );
  ANDN U6181 ( .B(n5983), .A(n5734), .Z(n5979) );
  XOR U6182 ( .A(n5984), .B(n1163), .Z(out[1163]) );
  XNOR U6183 ( .A(n5985), .B(n3783), .Z(n1163) );
  IV U6184 ( .A(n1969), .Z(n3783) );
  ANDN U6185 ( .B(n5988), .A(n5736), .Z(n5984) );
  XOR U6186 ( .A(n5989), .B(n1167), .Z(out[1162]) );
  XNOR U6187 ( .A(n5990), .B(n3788), .Z(n1167) );
  IV U6188 ( .A(n1972), .Z(n3788) );
  ANDN U6189 ( .B(n5993), .A(n5738), .Z(n5989) );
  XOR U6190 ( .A(n5994), .B(n1175), .Z(out[1161]) );
  XOR U6191 ( .A(n5995), .B(n1975), .Z(n1175) );
  IV U6192 ( .A(n4494), .Z(n1975) );
  ANDN U6193 ( .B(n5998), .A(n5740), .Z(n5994) );
  XNOR U6194 ( .A(n5999), .B(n1180), .Z(out[1160]) );
  XOR U6195 ( .A(n6000), .B(n1978), .Z(n1180) );
  XNOR U6196 ( .A(n6001), .B(n6002), .Z(n1978) );
  ANDN U6197 ( .B(n6003), .A(n5742), .Z(n5999) );
  XOR U6198 ( .A(n6004), .B(n4110), .Z(out[115]) );
  XNOR U6199 ( .A(n6005), .B(n2460), .Z(n4110) );
  ANDN U6200 ( .B(n3099), .A(n3100), .Z(n6004) );
  XNOR U6201 ( .A(n6006), .B(n2235), .Z(n3100) );
  IV U6202 ( .A(n6007), .Z(n2235) );
  XNOR U6203 ( .A(n6008), .B(n2298), .Z(n3099) );
  XOR U6204 ( .A(n6009), .B(n1184), .Z(out[1159]) );
  IV U6205 ( .A(n5745), .Z(n1184) );
  XNOR U6206 ( .A(n6010), .B(n1981), .Z(n5745) );
  XNOR U6207 ( .A(n6011), .B(n6012), .Z(n1981) );
  ANDN U6208 ( .B(n6013), .A(n5744), .Z(n6009) );
  XOR U6209 ( .A(n6014), .B(n1187), .Z(out[1158]) );
  XOR U6210 ( .A(n6015), .B(n1984), .Z(n1187) );
  XNOR U6211 ( .A(n6016), .B(n6017), .Z(n1984) );
  XOR U6212 ( .A(n6019), .B(n1191), .Z(out[1157]) );
  IV U6213 ( .A(n5750), .Z(n1191) );
  XOR U6214 ( .A(n6020), .B(n3813), .Z(n5750) );
  XNOR U6215 ( .A(n6021), .B(n6022), .Z(n3813) );
  ANDN U6216 ( .B(n6023), .A(n5749), .Z(n6019) );
  XOR U6217 ( .A(n6024), .B(n1196), .Z(out[1156]) );
  XOR U6218 ( .A(n6025), .B(n3820), .Z(n1196) );
  XNOR U6219 ( .A(n6026), .B(n6027), .Z(n3820) );
  ANDN U6220 ( .B(n6028), .A(n5752), .Z(n6024) );
  XNOR U6221 ( .A(n6029), .B(n1199), .Z(out[1155]) );
  XOR U6222 ( .A(n6030), .B(n1997), .Z(n1199) );
  XNOR U6223 ( .A(n6031), .B(n6032), .Z(n1997) );
  AND U6224 ( .A(n6033), .B(n6034), .Z(n6029) );
  XOR U6225 ( .A(n6035), .B(n1203), .Z(out[1154]) );
  IV U6226 ( .A(n5761), .Z(n1203) );
  XNOR U6227 ( .A(n6036), .B(n2000), .Z(n5761) );
  XOR U6228 ( .A(n6037), .B(n6038), .Z(n2000) );
  NOR U6229 ( .A(n6039), .B(n5760), .Z(n6035) );
  XNOR U6230 ( .A(n6040), .B(n1208), .Z(out[1153]) );
  XOR U6231 ( .A(n6041), .B(n3837), .Z(n1208) );
  XNOR U6232 ( .A(n6042), .B(n6043), .Z(n3837) );
  NOR U6233 ( .A(n6044), .B(n5763), .Z(n6040) );
  XOR U6234 ( .A(n6045), .B(n1211), .Z(out[1152]) );
  XOR U6235 ( .A(n6046), .B(n2006), .Z(n1211) );
  XNOR U6236 ( .A(n6047), .B(n6048), .Z(n2006) );
  NOR U6237 ( .A(n6049), .B(n5765), .Z(n6045) );
  XOR U6238 ( .A(n6050), .B(n5560), .Z(out[1151]) );
  XNOR U6239 ( .A(n6051), .B(n2562), .Z(n5560) );
  ANDN U6240 ( .B(n6052), .A(n5767), .Z(n6050) );
  XOR U6241 ( .A(n6053), .B(n5564), .Z(out[1150]) );
  XOR U6242 ( .A(n6054), .B(n2569), .Z(n5564) );
  ANDN U6243 ( .B(n6055), .A(n5769), .Z(n6053) );
  XOR U6244 ( .A(n6056), .B(n4113), .Z(out[114]) );
  XOR U6245 ( .A(n6057), .B(n2467), .Z(n4113) );
  ANDN U6246 ( .B(n3127), .A(n3128), .Z(n6056) );
  XNOR U6247 ( .A(n6058), .B(n2240), .Z(n3128) );
  XNOR U6248 ( .A(n6059), .B(n3144), .Z(n3127) );
  IV U6249 ( .A(n2309), .Z(n3144) );
  XOR U6250 ( .A(n6060), .B(n5568), .Z(out[1149]) );
  XNOR U6251 ( .A(n5272), .B(n6061), .Z(n5568) );
  XOR U6252 ( .A(n6062), .B(n6063), .Z(n5272) );
  ANDN U6253 ( .B(n6064), .A(n5771), .Z(n6060) );
  XOR U6254 ( .A(n6065), .B(n5572), .Z(out[1148]) );
  XNOR U6255 ( .A(n5277), .B(n6066), .Z(n5572) );
  XOR U6256 ( .A(n6067), .B(n6068), .Z(n5277) );
  ANDN U6257 ( .B(n6069), .A(n5773), .Z(n6065) );
  XOR U6258 ( .A(n6070), .B(n5576), .Z(out[1147]) );
  XOR U6259 ( .A(n4343), .B(n6071), .Z(n5576) );
  XOR U6260 ( .A(n6072), .B(n6073), .Z(n4343) );
  XOR U6261 ( .A(n6075), .B(n5580), .Z(out[1146]) );
  XOR U6262 ( .A(n6076), .B(n2601), .Z(n5580) );
  XOR U6263 ( .A(n6077), .B(n6078), .Z(n2601) );
  ANDN U6264 ( .B(n6079), .A(n5777), .Z(n6075) );
  XOR U6265 ( .A(n6080), .B(n5584), .Z(out[1145]) );
  XOR U6266 ( .A(n6081), .B(n2608), .Z(n5584) );
  XNOR U6267 ( .A(n6082), .B(n6083), .Z(n2608) );
  ANDN U6268 ( .B(n6084), .A(n5783), .Z(n6080) );
  XOR U6269 ( .A(n6085), .B(n5588), .Z(out[1144]) );
  XOR U6270 ( .A(n6086), .B(n2615), .Z(n5588) );
  XOR U6271 ( .A(n6087), .B(n6088), .Z(n2615) );
  AND U6272 ( .A(n5785), .B(n6089), .Z(n6085) );
  XOR U6273 ( .A(n6090), .B(n5592), .Z(out[1143]) );
  XOR U6274 ( .A(n6091), .B(n2622), .Z(n5592) );
  XNOR U6275 ( .A(n6092), .B(n6093), .Z(n2622) );
  ANDN U6276 ( .B(n6094), .A(n5787), .Z(n6090) );
  XOR U6277 ( .A(n6095), .B(n5596), .Z(out[1142]) );
  XOR U6278 ( .A(n6096), .B(n3758), .Z(n5596) );
  IV U6279 ( .A(n2629), .Z(n3758) );
  XNOR U6280 ( .A(n6097), .B(n6098), .Z(n2629) );
  ANDN U6281 ( .B(n6099), .A(n5789), .Z(n6095) );
  XOR U6282 ( .A(n6100), .B(n5604), .Z(out[1141]) );
  XOR U6283 ( .A(n6101), .B(n2636), .Z(n5604) );
  XNOR U6284 ( .A(n6102), .B(n6103), .Z(n2636) );
  ANDN U6285 ( .B(n6104), .A(n5791), .Z(n6100) );
  XOR U6286 ( .A(n6105), .B(n5608), .Z(out[1140]) );
  XNOR U6287 ( .A(n6106), .B(n2643), .Z(n5608) );
  XNOR U6288 ( .A(n6107), .B(n6108), .Z(n2643) );
  XOR U6289 ( .A(n6110), .B(n4117), .Z(out[113]) );
  XOR U6290 ( .A(n6111), .B(n3654), .Z(n4117) );
  AND U6291 ( .A(n3169), .B(n3171), .Z(n6110) );
  XNOR U6292 ( .A(n6112), .B(n2247), .Z(n3171) );
  XNOR U6293 ( .A(n6113), .B(n2316), .Z(n3169) );
  IV U6294 ( .A(n6114), .Z(n2316) );
  XOR U6295 ( .A(n6115), .B(n5612), .Z(out[1139]) );
  XNOR U6296 ( .A(n6116), .B(n3773), .Z(n5612) );
  IV U6297 ( .A(n2650), .Z(n3773) );
  XNOR U6298 ( .A(n6117), .B(n6118), .Z(n2650) );
  ANDN U6299 ( .B(n6119), .A(n5795), .Z(n6115) );
  XOR U6300 ( .A(n6120), .B(n5616), .Z(out[1138]) );
  IV U6301 ( .A(n5798), .Z(n5616) );
  XOR U6302 ( .A(n6121), .B(n2657), .Z(n5798) );
  XNOR U6303 ( .A(n6122), .B(n6123), .Z(n2657) );
  ANDN U6304 ( .B(n6124), .A(n5797), .Z(n6120) );
  XOR U6305 ( .A(n6125), .B(n5620), .Z(out[1137]) );
  XNOR U6306 ( .A(n6126), .B(n2664), .Z(n5620) );
  XNOR U6307 ( .A(n6127), .B(n6128), .Z(n2664) );
  ANDN U6308 ( .B(n6129), .A(n5800), .Z(n6125) );
  XOR U6309 ( .A(n6130), .B(n5624), .Z(out[1136]) );
  XOR U6310 ( .A(n6131), .B(n2197), .Z(n5624) );
  XNOR U6311 ( .A(n6132), .B(n6133), .Z(n2197) );
  ANDN U6312 ( .B(n6134), .A(n5802), .Z(n6130) );
  XOR U6313 ( .A(n6135), .B(n5629), .Z(out[1135]) );
  IV U6314 ( .A(n5813), .Z(n5629) );
  XOR U6315 ( .A(n6136), .B(n2204), .Z(n5813) );
  IV U6316 ( .A(n3793), .Z(n2204) );
  XNOR U6317 ( .A(n6137), .B(n6138), .Z(n3793) );
  ANDN U6318 ( .B(n6139), .A(n5812), .Z(n6135) );
  XOR U6319 ( .A(n6140), .B(n5633), .Z(out[1134]) );
  IV U6320 ( .A(n5816), .Z(n5633) );
  XOR U6321 ( .A(n6141), .B(n5349), .Z(n5816) );
  XOR U6322 ( .A(n6142), .B(n6143), .Z(n5349) );
  ANDN U6323 ( .B(n6144), .A(n5815), .Z(n6140) );
  XOR U6324 ( .A(n6145), .B(n5636), .Z(out[1133]) );
  XNOR U6325 ( .A(n6146), .B(n3803), .Z(n5636) );
  XOR U6326 ( .A(n6147), .B(n6148), .Z(n3803) );
  ANDN U6327 ( .B(n6149), .A(n5818), .Z(n6145) );
  XOR U6328 ( .A(n6150), .B(n5640), .Z(out[1132]) );
  XOR U6329 ( .A(n6151), .B(n2231), .Z(n5640) );
  IV U6330 ( .A(n3809), .Z(n2231) );
  XOR U6331 ( .A(n6152), .B(n6153), .Z(n3809) );
  ANDN U6332 ( .B(n6154), .A(n5820), .Z(n6150) );
  XNOR U6333 ( .A(n6155), .B(n5650), .Z(out[1131]) );
  XNOR U6334 ( .A(n6156), .B(n2238), .Z(n5650) );
  IV U6335 ( .A(n3815), .Z(n2238) );
  XOR U6336 ( .A(n6157), .B(n6158), .Z(n3815) );
  AND U6337 ( .A(n5822), .B(n6159), .Z(n6155) );
  XOR U6338 ( .A(n6160), .B(n5653), .Z(out[1130]) );
  XNOR U6339 ( .A(n6161), .B(n3822), .Z(n5653) );
  XOR U6340 ( .A(n6162), .B(n6163), .Z(n3822) );
  AND U6341 ( .A(n5824), .B(n6164), .Z(n6160) );
  XOR U6342 ( .A(n6165), .B(n4120), .Z(out[112]) );
  XOR U6343 ( .A(n6166), .B(n2481), .Z(n4120) );
  ANDN U6344 ( .B(n3203), .A(n3205), .Z(n6165) );
  XNOR U6345 ( .A(n6167), .B(n2254), .Z(n3205) );
  XOR U6346 ( .A(n6168), .B(n2323), .Z(n3203) );
  IV U6347 ( .A(n5434), .Z(n2323) );
  XOR U6348 ( .A(n6169), .B(n5657), .Z(out[1129]) );
  XNOR U6349 ( .A(n6170), .B(n2252), .Z(n5657) );
  XOR U6350 ( .A(n6171), .B(n6172), .Z(n2252) );
  XNOR U6351 ( .A(n6174), .B(n5662), .Z(out[1128]) );
  XNOR U6352 ( .A(n6175), .B(n2259), .Z(n5662) );
  IV U6353 ( .A(n5379), .Z(n2259) );
  XOR U6354 ( .A(n6176), .B(n6177), .Z(n5379) );
  XOR U6355 ( .A(n6179), .B(n5664), .Z(out[1127]) );
  XNOR U6356 ( .A(n6180), .B(n3839), .Z(n5664) );
  XOR U6357 ( .A(n6181), .B(n6182), .Z(n3839) );
  XOR U6358 ( .A(n6183), .B(n5666), .Z(out[1126]) );
  XNOR U6359 ( .A(n6184), .B(n3845), .Z(n5666) );
  XOR U6360 ( .A(n6185), .B(n6186), .Z(n3845) );
  NOR U6361 ( .A(n1046), .B(n5838), .Z(n6183) );
  XOR U6362 ( .A(n6187), .B(n5668), .Z(out[1125]) );
  XNOR U6363 ( .A(n6188), .B(n3849), .Z(n5668) );
  XOR U6364 ( .A(n6189), .B(n6190), .Z(n3849) );
  XOR U6365 ( .A(n6191), .B(n5670), .Z(out[1124]) );
  XOR U6366 ( .A(n6192), .B(n2287), .Z(n5670) );
  IV U6367 ( .A(n5400), .Z(n2287) );
  XOR U6368 ( .A(n6193), .B(n6194), .Z(n5400) );
  NOR U6369 ( .A(n1054), .B(n5853), .Z(n6191) );
  XOR U6370 ( .A(n6195), .B(n5672), .Z(out[1123]) );
  XNOR U6371 ( .A(n6196), .B(n2294), .Z(n5672) );
  XOR U6372 ( .A(n6197), .B(n6198), .Z(n2294) );
  ANDN U6373 ( .B(n5858), .A(n1058), .Z(n6195) );
  XOR U6374 ( .A(n6199), .B(n5674), .Z(out[1122]) );
  XNOR U6375 ( .A(n6200), .B(n2305), .Z(n5674) );
  IV U6376 ( .A(n5170), .Z(n2305) );
  XOR U6377 ( .A(n6201), .B(n6202), .Z(n5170) );
  ANDN U6378 ( .B(n5863), .A(n1062), .Z(n6199) );
  XOR U6379 ( .A(n6203), .B(n5681), .Z(out[1121]) );
  XOR U6380 ( .A(n6204), .B(n5413), .Z(n5681) );
  XOR U6381 ( .A(n6205), .B(n6206), .Z(n5413) );
  ANDN U6382 ( .B(n5868), .A(n1066), .Z(n6203) );
  XOR U6383 ( .A(n6207), .B(n5683), .Z(out[1120]) );
  XOR U6384 ( .A(n6208), .B(n2319), .Z(n5683) );
  IV U6385 ( .A(n5229), .Z(n2319) );
  XOR U6386 ( .A(n6209), .B(n6210), .Z(n5229) );
  ANDN U6387 ( .B(n1070), .A(n5873), .Z(n6207) );
  XOR U6388 ( .A(n6211), .B(n4126), .Z(out[111]) );
  IV U6389 ( .A(n4302), .Z(n4126) );
  XOR U6390 ( .A(n6212), .B(n3663), .Z(n4302) );
  ANDN U6391 ( .B(n3240), .A(n3241), .Z(n6211) );
  XOR U6392 ( .A(n6213), .B(n2263), .Z(n3241) );
  XNOR U6393 ( .A(n6214), .B(n2328), .Z(n3240) );
  XOR U6394 ( .A(n6215), .B(n5685), .Z(out[1119]) );
  XNOR U6395 ( .A(n6216), .B(n2326), .Z(n5685) );
  IV U6396 ( .A(n5264), .Z(n2326) );
  XOR U6397 ( .A(n6217), .B(n6218), .Z(n5264) );
  NOR U6398 ( .A(n1074), .B(n5878), .Z(n6215) );
  XOR U6399 ( .A(n6219), .B(n5687), .Z(out[1118]) );
  XNOR U6400 ( .A(n6220), .B(n2333), .Z(n5687) );
  XNOR U6401 ( .A(n6221), .B(n6222), .Z(n2333) );
  XOR U6402 ( .A(n6223), .B(n5689), .Z(out[1117]) );
  XNOR U6403 ( .A(n6224), .B(n5367), .Z(n5689) );
  XOR U6404 ( .A(n6225), .B(n6226), .Z(n5367) );
  ANDN U6405 ( .B(n6227), .A(n1086), .Z(n6223) );
  XOR U6406 ( .A(n6228), .B(n5691), .Z(out[1116]) );
  XNOR U6407 ( .A(n6229), .B(n2347), .Z(n5691) );
  IV U6408 ( .A(n3565), .Z(n2347) );
  XOR U6409 ( .A(n6230), .B(n6231), .Z(n3565) );
  NOR U6410 ( .A(n1090), .B(n5893), .Z(n6228) );
  XOR U6411 ( .A(n6232), .B(n5693), .Z(out[1115]) );
  XNOR U6412 ( .A(n6233), .B(n5442), .Z(n5693) );
  XOR U6413 ( .A(n6234), .B(n6235), .Z(n5442) );
  XOR U6414 ( .A(n6236), .B(n5695), .Z(out[1114]) );
  XNOR U6415 ( .A(n6237), .B(n2361), .Z(n5695) );
  IV U6416 ( .A(n3579), .Z(n2361) );
  XOR U6417 ( .A(n6238), .B(n6239), .Z(n3579) );
  NOR U6418 ( .A(n1098), .B(n5908), .Z(n6236) );
  XOR U6419 ( .A(n6240), .B(n5697), .Z(out[1113]) );
  XNOR U6420 ( .A(n6241), .B(n5451), .Z(n5697) );
  XOR U6421 ( .A(n6242), .B(n6243), .Z(n5451) );
  ANDN U6422 ( .B(n5913), .A(n1102), .Z(n6240) );
  XOR U6423 ( .A(n6244), .B(n5699), .Z(out[1112]) );
  XNOR U6424 ( .A(n6245), .B(n3588), .Z(n5699) );
  XOR U6425 ( .A(n6246), .B(n6247), .Z(n3588) );
  XOR U6426 ( .A(n6248), .B(n5706), .Z(out[1111]) );
  XNOR U6427 ( .A(n6249), .B(n5644), .Z(n5706) );
  XOR U6428 ( .A(n6250), .B(n6251), .Z(n5644) );
  NOR U6429 ( .A(n5923), .B(n1110), .Z(n6248) );
  XOR U6430 ( .A(n6252), .B(n5708), .Z(out[1110]) );
  XOR U6431 ( .A(n6253), .B(n2393), .Z(n5708) );
  IV U6432 ( .A(n3598), .Z(n2393) );
  XOR U6433 ( .A(n6254), .B(n6255), .Z(n3598) );
  ANDN U6434 ( .B(n6256), .A(n1114), .Z(n6252) );
  XOR U6435 ( .A(n6257), .B(n4129), .Z(out[110]) );
  XNOR U6436 ( .A(n6258), .B(n2495), .Z(n4129) );
  ANDN U6437 ( .B(n3278), .A(n3279), .Z(n6257) );
  XNOR U6438 ( .A(n6259), .B(n2270), .Z(n3279) );
  XOR U6439 ( .A(n6260), .B(n2335), .Z(n3278) );
  XOR U6440 ( .A(n6261), .B(n5710), .Z(out[1109]) );
  XNOR U6441 ( .A(n6262), .B(n2400), .Z(n5710) );
  XNOR U6442 ( .A(n6263), .B(n6264), .Z(n2400) );
  NOR U6443 ( .A(n5933), .B(n1118), .Z(n6261) );
  XOR U6444 ( .A(n6265), .B(n5712), .Z(out[1108]) );
  XNOR U6445 ( .A(n6266), .B(n2407), .Z(n5712) );
  XNOR U6446 ( .A(n6267), .B(n6268), .Z(n2407) );
  ANDN U6447 ( .B(n6269), .A(n1122), .Z(n6265) );
  XOR U6448 ( .A(n6270), .B(n5714), .Z(out[1107]) );
  XNOR U6449 ( .A(n6271), .B(n2414), .Z(n5714) );
  XNOR U6450 ( .A(n6272), .B(n6273), .Z(n2414) );
  ANDN U6451 ( .B(n6274), .A(n1130), .Z(n6270) );
  XOR U6452 ( .A(n6275), .B(n5716), .Z(out[1106]) );
  XOR U6453 ( .A(n6276), .B(n2421), .Z(n5716) );
  XNOR U6454 ( .A(n6277), .B(n6278), .Z(n2421) );
  ANDN U6455 ( .B(n6279), .A(n1134), .Z(n6275) );
  XOR U6456 ( .A(n6280), .B(n5718), .Z(out[1105]) );
  XNOR U6457 ( .A(n6281), .B(n2428), .Z(n5718) );
  XNOR U6458 ( .A(n6282), .B(n6283), .Z(n2428) );
  NOR U6459 ( .A(n5958), .B(n1138), .Z(n6280) );
  XOR U6460 ( .A(n6284), .B(n5720), .Z(out[1104]) );
  XNOR U6461 ( .A(n6285), .B(n5841), .Z(n5720) );
  XOR U6462 ( .A(n6286), .B(n6287), .Z(n5841) );
  ANDN U6463 ( .B(n5963), .A(n1142), .Z(n6284) );
  XOR U6464 ( .A(n6288), .B(n5723), .Z(out[1103]) );
  XNOR U6465 ( .A(n6289), .B(n2442), .Z(n5723) );
  IV U6466 ( .A(n3632), .Z(n2442) );
  XOR U6467 ( .A(n6290), .B(n6291), .Z(n3632) );
  NOR U6468 ( .A(n1146), .B(n5968), .Z(n6288) );
  XOR U6469 ( .A(n6292), .B(n5725), .Z(out[1102]) );
  XOR U6470 ( .A(n6293), .B(n2453), .Z(n5725) );
  XNOR U6471 ( .A(n6294), .B(n6295), .Z(n2453) );
  ANDN U6472 ( .B(n5973), .A(n1150), .Z(n6292) );
  XOR U6473 ( .A(n6296), .B(n5732), .Z(out[1101]) );
  XNOR U6474 ( .A(n6297), .B(n2460), .Z(n5732) );
  IV U6475 ( .A(n3642), .Z(n2460) );
  XNOR U6476 ( .A(n6298), .B(n6299), .Z(n3642) );
  NOR U6477 ( .A(n1154), .B(n5978), .Z(n6296) );
  XOR U6478 ( .A(n6300), .B(n5734), .Z(out[1100]) );
  XOR U6479 ( .A(n6301), .B(n2467), .Z(n5734) );
  XNOR U6480 ( .A(n6302), .B(n6303), .Z(n2467) );
  NOR U6481 ( .A(n1158), .B(n5983), .Z(n6300) );
  XOR U6482 ( .A(n6304), .B(n2028), .Z(out[10]) );
  XOR U6483 ( .A(n6305), .B(n2603), .Z(n2028) );
  IV U6484 ( .A(n5303), .Z(n2603) );
  NOR U6485 ( .A(n4028), .B(n2027), .Z(n6304) );
  XNOR U6486 ( .A(n2535), .B(n6306), .Z(n2027) );
  XNOR U6487 ( .A(n6307), .B(n1752), .Z(n4028) );
  XOR U6488 ( .A(n6308), .B(n4132), .Z(out[109]) );
  IV U6489 ( .A(n4307), .Z(n4132) );
  XOR U6490 ( .A(n6309), .B(n6310), .Z(n4307) );
  ANDN U6491 ( .B(n3316), .A(n3318), .Z(n6308) );
  XNOR U6492 ( .A(n6311), .B(n2275), .Z(n3318) );
  XNOR U6493 ( .A(n6312), .B(n3161), .Z(n3316) );
  XOR U6494 ( .A(n6313), .B(n5736), .Z(out[1099]) );
  XOR U6495 ( .A(n6314), .B(n3654), .Z(n5736) );
  XNOR U6496 ( .A(n6315), .B(n6316), .Z(n3654) );
  NOR U6497 ( .A(n5988), .B(n1162), .Z(n6313) );
  XOR U6498 ( .A(n6317), .B(n5738), .Z(out[1098]) );
  XOR U6499 ( .A(n6318), .B(n2481), .Z(n5738) );
  XNOR U6500 ( .A(n6319), .B(n6320), .Z(n2481) );
  NOR U6501 ( .A(n5993), .B(n1166), .Z(n6317) );
  XOR U6502 ( .A(n6321), .B(n5740), .Z(out[1097]) );
  XOR U6503 ( .A(n6322), .B(n2488), .Z(n5740) );
  IV U6504 ( .A(n3663), .Z(n2488) );
  XNOR U6505 ( .A(n6323), .B(n6324), .Z(n3663) );
  NOR U6506 ( .A(n1174), .B(n5998), .Z(n6321) );
  XOR U6507 ( .A(n6325), .B(n5742), .Z(out[1096]) );
  XNOR U6508 ( .A(n6326), .B(n2495), .Z(n5742) );
  XNOR U6509 ( .A(n6327), .B(n6328), .Z(n2495) );
  NOR U6510 ( .A(n6003), .B(n1178), .Z(n6325) );
  XOR U6511 ( .A(n6329), .B(n5744), .Z(out[1095]) );
  XOR U6512 ( .A(n6330), .B(n2502), .Z(n5744) );
  IV U6513 ( .A(n6310), .Z(n2502) );
  XNOR U6514 ( .A(n6331), .B(n6332), .Z(n6310) );
  NOR U6515 ( .A(n6013), .B(n1182), .Z(n6329) );
  XOR U6516 ( .A(n6333), .B(n5747), .Z(out[1094]) );
  XNOR U6517 ( .A(n6334), .B(n2509), .Z(n5747) );
  ANDN U6518 ( .B(n6018), .A(n1186), .Z(n6333) );
  XOR U6519 ( .A(n6335), .B(n5749), .Z(out[1093]) );
  XNOR U6520 ( .A(n6336), .B(n3687), .Z(n5749) );
  IV U6521 ( .A(n2516), .Z(n3687) );
  ANDN U6522 ( .B(n1190), .A(n6023), .Z(n6335) );
  XOR U6523 ( .A(n6337), .B(n5752), .Z(out[1092]) );
  XNOR U6524 ( .A(n6338), .B(n3693), .Z(n5752) );
  IV U6525 ( .A(n2527), .Z(n3693) );
  NOR U6526 ( .A(n1194), .B(n6028), .Z(n6337) );
  XOR U6527 ( .A(n6339), .B(n5758), .Z(out[1091]) );
  IV U6528 ( .A(n6034), .Z(n5758) );
  XOR U6529 ( .A(n6340), .B(n2534), .Z(n6034) );
  ANDN U6530 ( .B(n6341), .A(n6033), .Z(n6339) );
  XOR U6531 ( .A(n6342), .B(n5760), .Z(out[1090]) );
  XNOR U6532 ( .A(n6343), .B(n2541), .Z(n5760) );
  AND U6533 ( .A(n1202), .B(n6039), .Z(n6342) );
  IV U6534 ( .A(n6344), .Z(n6039) );
  XOR U6535 ( .A(n6345), .B(n4135), .Z(out[108]) );
  XNOR U6536 ( .A(n6346), .B(n2509), .Z(n4135) );
  XNOR U6537 ( .A(n6347), .B(n6348), .Z(n2509) );
  ANDN U6538 ( .B(n3358), .A(n3359), .Z(n6345) );
  XOR U6539 ( .A(n6349), .B(n2282), .Z(n3359) );
  XNOR U6540 ( .A(n6350), .B(n2349), .Z(n3358) );
  XOR U6541 ( .A(n6351), .B(n5763), .Z(out[1089]) );
  XOR U6542 ( .A(n6352), .B(n2548), .Z(n5763) );
  AND U6543 ( .A(n6044), .B(n6353), .Z(n6351) );
  XOR U6544 ( .A(n6354), .B(n5765), .Z(out[1088]) );
  XOR U6545 ( .A(n6355), .B(n2555), .Z(n5765) );
  ANDN U6546 ( .B(n6049), .A(n1210), .Z(n6354) );
  XOR U6547 ( .A(n6356), .B(n5767), .Z(out[1087]) );
  XOR U6548 ( .A(n6357), .B(n2531), .Z(n5767) );
  XNOR U6549 ( .A(n5831), .B(n6358), .Z(n2531) );
  XOR U6550 ( .A(n6359), .B(n6360), .Z(n5831) );
  XNOR U6551 ( .A(n6262), .B(n2399), .Z(n6360) );
  XOR U6552 ( .A(n6361), .B(n6362), .Z(n2399) );
  ANDN U6553 ( .B(n6363), .A(n6364), .Z(n6361) );
  XOR U6554 ( .A(n6365), .B(n6366), .Z(n6262) );
  NOR U6555 ( .A(n6367), .B(n6368), .Z(n6365) );
  XOR U6556 ( .A(n3601), .B(n6369), .Z(n6359) );
  XNOR U6557 ( .A(n5702), .B(n5477), .Z(n6369) );
  XNOR U6558 ( .A(n6370), .B(n6371), .Z(n5477) );
  ANDN U6559 ( .B(n6372), .A(n6373), .Z(n6370) );
  XNOR U6560 ( .A(n6374), .B(n6375), .Z(n5702) );
  ANDN U6561 ( .B(n6376), .A(n6377), .Z(n6374) );
  XNOR U6562 ( .A(n6378), .B(n6379), .Z(n3601) );
  ANDN U6563 ( .B(n6380), .A(n6381), .Z(n6378) );
  ANDN U6564 ( .B(n5559), .A(n6052), .Z(n6356) );
  XOR U6565 ( .A(n6382), .B(n5769), .Z(out[1086]) );
  XOR U6566 ( .A(n6383), .B(n2538), .Z(n5769) );
  XOR U6567 ( .A(n5836), .B(n6384), .Z(n2538) );
  XOR U6568 ( .A(n6385), .B(n6386), .Z(n5836) );
  XOR U6569 ( .A(n6266), .B(n2406), .Z(n6386) );
  XNOR U6570 ( .A(n6387), .B(n6388), .Z(n2406) );
  XOR U6571 ( .A(n6391), .B(n6392), .Z(n6266) );
  XNOR U6572 ( .A(n3605), .B(n6395), .Z(n6385) );
  XNOR U6573 ( .A(n5727), .B(n5481), .Z(n6395) );
  XOR U6574 ( .A(n6396), .B(n6397), .Z(n5481) );
  ANDN U6575 ( .B(n6398), .A(n6399), .Z(n6396) );
  XOR U6576 ( .A(n6400), .B(n6401), .Z(n5727) );
  ANDN U6577 ( .B(n6402), .A(n6403), .Z(n6400) );
  XOR U6578 ( .A(n6404), .B(n6405), .Z(n3605) );
  AND U6579 ( .A(n6406), .B(n6407), .Z(n6404) );
  AND U6580 ( .A(n5563), .B(n6408), .Z(n6382) );
  XOR U6581 ( .A(n6409), .B(n5771), .Z(out[1085]) );
  XNOR U6582 ( .A(n6410), .B(n2543), .Z(n5771) );
  XNOR U6583 ( .A(n5846), .B(n6411), .Z(n2543) );
  XOR U6584 ( .A(n6412), .B(n6413), .Z(n5846) );
  XNOR U6585 ( .A(n6271), .B(n2413), .Z(n6413) );
  XOR U6586 ( .A(n6414), .B(n6415), .Z(n2413) );
  NOR U6587 ( .A(n6416), .B(n6417), .Z(n6414) );
  XOR U6588 ( .A(n6418), .B(n6419), .Z(n6271) );
  AND U6589 ( .A(n6420), .B(n6421), .Z(n6418) );
  XOR U6590 ( .A(n3609), .B(n6422), .Z(n6412) );
  XNOR U6591 ( .A(n5754), .B(n5485), .Z(n6422) );
  XNOR U6592 ( .A(n6423), .B(n6424), .Z(n5485) );
  ANDN U6593 ( .B(n6425), .A(n6426), .Z(n6423) );
  XOR U6594 ( .A(n6427), .B(n6428), .Z(n5754) );
  NOR U6595 ( .A(n6429), .B(n6430), .Z(n6427) );
  XOR U6596 ( .A(n6431), .B(n6432), .Z(n3609) );
  ANDN U6597 ( .B(n6433), .A(n6434), .Z(n6431) );
  AND U6598 ( .A(n5567), .B(n6435), .Z(n6409) );
  XOR U6599 ( .A(n6436), .B(n5773), .Z(out[1084]) );
  XOR U6600 ( .A(n6437), .B(n2550), .Z(n5773) );
  XOR U6601 ( .A(n5851), .B(n6438), .Z(n2550) );
  XOR U6602 ( .A(n6439), .B(n6440), .Z(n5851) );
  XOR U6603 ( .A(n6276), .B(n2420), .Z(n6440) );
  XOR U6604 ( .A(n6441), .B(n6442), .Z(n2420) );
  ANDN U6605 ( .B(n6443), .A(n6444), .Z(n6441) );
  XNOR U6606 ( .A(n6445), .B(n6446), .Z(n6276) );
  XOR U6607 ( .A(n3613), .B(n6449), .Z(n6439) );
  XNOR U6608 ( .A(n5779), .B(n5488), .Z(n6449) );
  XOR U6609 ( .A(n6450), .B(n6451), .Z(n5488) );
  XOR U6610 ( .A(n6452), .B(n6453), .Z(n6451) );
  NAND U6611 ( .A(n4364), .B(n4650), .Z(n6453) );
  AND U6612 ( .A(n6454), .B(n6455), .Z(n4650) );
  NOR U6613 ( .A(n6456), .B(n6457), .Z(n6452) );
  XNOR U6614 ( .A(n6458), .B(n6459), .Z(n5779) );
  XNOR U6615 ( .A(n6462), .B(n6463), .Z(n3613) );
  ANDN U6616 ( .B(n6464), .A(n6465), .Z(n6462) );
  ANDN U6617 ( .B(n5571), .A(n6069), .Z(n6436) );
  XOR U6618 ( .A(n6466), .B(n5775), .Z(out[1083]) );
  XOR U6619 ( .A(n6467), .B(n2557), .Z(n5775) );
  XNOR U6620 ( .A(n5856), .B(n6468), .Z(n2557) );
  XOR U6621 ( .A(n6469), .B(n6470), .Z(n5856) );
  XNOR U6622 ( .A(n6281), .B(n2427), .Z(n6470) );
  XOR U6623 ( .A(n6471), .B(n6472), .Z(n2427) );
  NOR U6624 ( .A(n6473), .B(n6474), .Z(n6471) );
  XNOR U6625 ( .A(n6475), .B(n6476), .Z(n6281) );
  NOR U6626 ( .A(n6477), .B(n6478), .Z(n6475) );
  XOR U6627 ( .A(n3618), .B(n6479), .Z(n6469) );
  XNOR U6628 ( .A(n5808), .B(n5493), .Z(n6479) );
  XNOR U6629 ( .A(n6480), .B(n6481), .Z(n5493) );
  AND U6630 ( .A(n6482), .B(n6483), .Z(n6480) );
  XOR U6631 ( .A(n6484), .B(n6485), .Z(n5808) );
  AND U6632 ( .A(n6486), .B(n6487), .Z(n6484) );
  XNOR U6633 ( .A(n6488), .B(n6489), .Z(n3618) );
  NOR U6634 ( .A(n6490), .B(n6491), .Z(n6488) );
  AND U6635 ( .A(n5575), .B(n6074), .Z(n6466) );
  XOR U6636 ( .A(n6492), .B(n5777), .Z(out[1082]) );
  XOR U6637 ( .A(n6493), .B(n2566), .Z(n5777) );
  XNOR U6638 ( .A(n5861), .B(n6494), .Z(n2566) );
  XOR U6639 ( .A(n6495), .B(n6496), .Z(n5861) );
  XOR U6640 ( .A(n6285), .B(n2434), .Z(n6496) );
  XOR U6641 ( .A(n6497), .B(n6498), .Z(n2434) );
  ANDN U6642 ( .B(n6499), .A(n6500), .Z(n6497) );
  XNOR U6643 ( .A(n6501), .B(n6502), .Z(n6285) );
  AND U6644 ( .A(n6503), .B(n6504), .Z(n6501) );
  XOR U6645 ( .A(n3625), .B(n6505), .Z(n6495) );
  XOR U6646 ( .A(n5840), .B(n5497), .Z(n6505) );
  XNOR U6647 ( .A(n6506), .B(n6507), .Z(n5497) );
  ANDN U6648 ( .B(n6508), .A(n6509), .Z(n6506) );
  XOR U6649 ( .A(n6510), .B(n6511), .Z(n5840) );
  ANDN U6650 ( .B(n6512), .A(n6513), .Z(n6510) );
  XOR U6651 ( .A(n6514), .B(n6515), .Z(n3625) );
  ANDN U6652 ( .B(n6516), .A(n6517), .Z(n6514) );
  ANDN U6653 ( .B(n5579), .A(n6079), .Z(n6492) );
  XOR U6654 ( .A(n6518), .B(n5783), .Z(out[1081]) );
  XOR U6655 ( .A(n6519), .B(n5283), .Z(n5783) );
  XOR U6656 ( .A(n6520), .B(n5867), .Z(n5283) );
  XNOR U6657 ( .A(n6521), .B(n6522), .Z(n5867) );
  XOR U6658 ( .A(n5500), .B(n3631), .Z(n6522) );
  XOR U6659 ( .A(n6523), .B(n6524), .Z(n3631) );
  AND U6660 ( .A(n6525), .B(n6526), .Z(n6523) );
  XNOR U6661 ( .A(n6527), .B(n6528), .Z(n5500) );
  AND U6662 ( .A(n6529), .B(n6530), .Z(n6527) );
  XOR U6663 ( .A(n6289), .B(n6531), .Z(n6521) );
  XOR U6664 ( .A(n2441), .B(n5895), .Z(n6531) );
  XNOR U6665 ( .A(n6532), .B(n6533), .Z(n5895) );
  NOR U6666 ( .A(n6534), .B(n6535), .Z(n6532) );
  XOR U6667 ( .A(n6536), .B(n6537), .Z(n2441) );
  XNOR U6668 ( .A(n6540), .B(n6541), .Z(n6289) );
  ANDN U6669 ( .B(n6542), .A(n6543), .Z(n6540) );
  AND U6670 ( .A(n5583), .B(n6544), .Z(n6518) );
  XNOR U6671 ( .A(n6545), .B(n5785), .Z(out[1080]) );
  XNOR U6672 ( .A(n6546), .B(n2580), .Z(n5785) );
  XNOR U6673 ( .A(n6547), .B(n5872), .Z(n2580) );
  XNOR U6674 ( .A(n6548), .B(n6549), .Z(n5872) );
  XNOR U6675 ( .A(n5505), .B(n3636), .Z(n6549) );
  XOR U6676 ( .A(n6550), .B(n6551), .Z(n3636) );
  NOR U6677 ( .A(n6552), .B(n6553), .Z(n6550) );
  XOR U6678 ( .A(n6554), .B(n6555), .Z(n5505) );
  NOR U6679 ( .A(n6556), .B(n6557), .Z(n6554) );
  XNOR U6680 ( .A(n6293), .B(n6558), .Z(n6548) );
  XNOR U6681 ( .A(n2452), .B(n5950), .Z(n6558) );
  XNOR U6682 ( .A(n6559), .B(n6560), .Z(n5950) );
  XNOR U6683 ( .A(n6563), .B(n6564), .Z(n2452) );
  AND U6684 ( .A(n6565), .B(n6566), .Z(n6563) );
  XNOR U6685 ( .A(n6567), .B(n6568), .Z(n6293) );
  AND U6686 ( .A(n6569), .B(n6570), .Z(n6567) );
  AND U6687 ( .A(n5587), .B(n6571), .Z(n6545) );
  XOR U6688 ( .A(n6572), .B(n4138), .Z(out[107]) );
  XOR U6689 ( .A(n6573), .B(n2516), .Z(n4138) );
  XNOR U6690 ( .A(n6574), .B(n6575), .Z(n2516) );
  AND U6691 ( .A(n3390), .B(n4312), .Z(n6572) );
  XNOR U6692 ( .A(n6576), .B(n2356), .Z(n4312) );
  XNOR U6693 ( .A(n6577), .B(n2289), .Z(n3390) );
  XOR U6694 ( .A(n6578), .B(n5787), .Z(out[1079]) );
  XNOR U6695 ( .A(n6579), .B(n5292), .Z(n5787) );
  XOR U6696 ( .A(n6580), .B(n5877), .Z(n5292) );
  XNOR U6697 ( .A(n6581), .B(n6582), .Z(n5877) );
  XNOR U6698 ( .A(n5508), .B(n3641), .Z(n6582) );
  XOR U6699 ( .A(n6583), .B(n6584), .Z(n3641) );
  AND U6700 ( .A(n6585), .B(n6586), .Z(n6583) );
  XNOR U6701 ( .A(n6587), .B(n6588), .Z(n5508) );
  AND U6702 ( .A(n6589), .B(n6590), .Z(n6587) );
  XOR U6703 ( .A(n6297), .B(n6591), .Z(n6581) );
  XOR U6704 ( .A(n2459), .B(n6005), .Z(n6591) );
  XOR U6705 ( .A(n6592), .B(n6593), .Z(n6005) );
  XNOR U6706 ( .A(n6596), .B(n6597), .Z(n2459) );
  ANDN U6707 ( .B(n6598), .A(n6599), .Z(n6596) );
  XNOR U6708 ( .A(n6600), .B(n6601), .Z(n6297) );
  AND U6709 ( .A(n5591), .B(n6604), .Z(n6578) );
  IV U6710 ( .A(n6605), .Z(n5591) );
  XOR U6711 ( .A(n6606), .B(n5789), .Z(out[1078]) );
  XNOR U6712 ( .A(n6607), .B(n5298), .Z(n5789) );
  XOR U6713 ( .A(n6608), .B(n5882), .Z(n5298) );
  XNOR U6714 ( .A(n6609), .B(n6610), .Z(n5882) );
  XNOR U6715 ( .A(n5515), .B(n3648), .Z(n6610) );
  XOR U6716 ( .A(n6611), .B(n6612), .Z(n3648) );
  AND U6717 ( .A(n6613), .B(n6614), .Z(n6611) );
  XNOR U6718 ( .A(n6615), .B(n6616), .Z(n5515) );
  AND U6719 ( .A(n6617), .B(n6618), .Z(n6615) );
  XNOR U6720 ( .A(n6301), .B(n6619), .Z(n6609) );
  XOR U6721 ( .A(n2466), .B(n6057), .Z(n6619) );
  XNOR U6722 ( .A(n6620), .B(n6621), .Z(n6057) );
  ANDN U6723 ( .B(n6622), .A(n6623), .Z(n6620) );
  XOR U6724 ( .A(n6624), .B(n6625), .Z(n2466) );
  AND U6725 ( .A(n6626), .B(n6627), .Z(n6624) );
  XNOR U6726 ( .A(n6628), .B(n6629), .Z(n6301) );
  NOR U6727 ( .A(n6630), .B(n6631), .Z(n6628) );
  ANDN U6728 ( .B(n5595), .A(n6099), .Z(n6606) );
  IV U6729 ( .A(n6632), .Z(n5595) );
  XOR U6730 ( .A(n6633), .B(n5791), .Z(out[1077]) );
  XOR U6731 ( .A(n6634), .B(n5303), .Z(n5791) );
  XOR U6732 ( .A(n6635), .B(n5887), .Z(n5303) );
  XNOR U6733 ( .A(n6636), .B(n6637), .Z(n5887) );
  XNOR U6734 ( .A(n5520), .B(n3653), .Z(n6637) );
  XOR U6735 ( .A(n6638), .B(n6639), .Z(n3653) );
  ANDN U6736 ( .B(n6640), .A(n6641), .Z(n6638) );
  XNOR U6737 ( .A(n6642), .B(n6643), .Z(n5520) );
  NOR U6738 ( .A(n6644), .B(n6645), .Z(n6642) );
  XNOR U6739 ( .A(n6314), .B(n6646), .Z(n6636) );
  XOR U6740 ( .A(n2473), .B(n6111), .Z(n6646) );
  XNOR U6741 ( .A(n6647), .B(n6648), .Z(n6111) );
  ANDN U6742 ( .B(n6649), .A(n6650), .Z(n6647) );
  XNOR U6743 ( .A(n6651), .B(n6652), .Z(n2473) );
  XNOR U6744 ( .A(n6655), .B(n6656), .Z(n6314) );
  AND U6745 ( .A(n6657), .B(n6658), .Z(n6655) );
  ANDN U6746 ( .B(n5603), .A(n6104), .Z(n6633) );
  IV U6747 ( .A(n6659), .Z(n5603) );
  XOR U6748 ( .A(n6660), .B(n5793), .Z(out[1076]) );
  XOR U6749 ( .A(n5308), .B(n6661), .Z(n5793) );
  XOR U6750 ( .A(n5891), .B(n6662), .Z(n5308) );
  XOR U6751 ( .A(n6663), .B(n6664), .Z(n5891) );
  XOR U6752 ( .A(n6318), .B(n2480), .Z(n6664) );
  XNOR U6753 ( .A(n6665), .B(n6666), .Z(n2480) );
  ANDN U6754 ( .B(n6667), .A(n6668), .Z(n6665) );
  XNOR U6755 ( .A(n6669), .B(n6670), .Z(n6318) );
  NOR U6756 ( .A(n6671), .B(n6672), .Z(n6669) );
  XOR U6757 ( .A(n3658), .B(n6673), .Z(n6663) );
  XNOR U6758 ( .A(n6166), .B(n5523), .Z(n6673) );
  XOR U6759 ( .A(n6674), .B(n6675), .Z(n5523) );
  XOR U6760 ( .A(n6676), .B(n6677), .Z(n6675) );
  NOR U6761 ( .A(n6678), .B(n6679), .Z(n6676) );
  XNOR U6762 ( .A(n6680), .B(n6681), .Z(n6166) );
  ANDN U6763 ( .B(n6682), .A(n6683), .Z(n6680) );
  XOR U6764 ( .A(n6684), .B(n6685), .Z(n3658) );
  ANDN U6765 ( .B(n5607), .A(n6109), .Z(n6660) );
  XOR U6766 ( .A(n6688), .B(n5795), .Z(out[1075]) );
  XOR U6767 ( .A(n6689), .B(n2619), .Z(n5795) );
  XOR U6768 ( .A(n6690), .B(n5902), .Z(n2619) );
  XNOR U6769 ( .A(n6691), .B(n6692), .Z(n5902) );
  XNOR U6770 ( .A(n5527), .B(n3662), .Z(n6692) );
  XNOR U6771 ( .A(n6693), .B(n6694), .Z(n3662) );
  ANDN U6772 ( .B(n6695), .A(n6696), .Z(n6693) );
  XNOR U6773 ( .A(n6697), .B(n6698), .Z(n5527) );
  ANDN U6774 ( .B(n6699), .A(n6700), .Z(n6697) );
  XNOR U6775 ( .A(n6322), .B(n6701), .Z(n6691) );
  XOR U6776 ( .A(n2487), .B(n6212), .Z(n6701) );
  XNOR U6777 ( .A(n6702), .B(n6703), .Z(n6212) );
  NOR U6778 ( .A(n6704), .B(n6705), .Z(n6702) );
  XOR U6779 ( .A(n6706), .B(n6707), .Z(n2487) );
  ANDN U6780 ( .B(n6708), .A(n6709), .Z(n6706) );
  XNOR U6781 ( .A(n6710), .B(n6711), .Z(n6322) );
  ANDN U6782 ( .B(n6712), .A(n6713), .Z(n6710) );
  NOR U6783 ( .A(n6119), .B(n5611), .Z(n6688) );
  XOR U6784 ( .A(n6714), .B(n5797), .Z(out[1074]) );
  XNOR U6785 ( .A(n6715), .B(n2626), .Z(n5797) );
  XOR U6786 ( .A(n6716), .B(n5907), .Z(n2626) );
  XNOR U6787 ( .A(n6717), .B(n6718), .Z(n5907) );
  XOR U6788 ( .A(n5532), .B(n3668), .Z(n6718) );
  XOR U6789 ( .A(n6719), .B(n6720), .Z(n3668) );
  AND U6790 ( .A(n6721), .B(n6722), .Z(n6719) );
  XNOR U6791 ( .A(n6723), .B(n6724), .Z(n5532) );
  AND U6792 ( .A(n6725), .B(n6726), .Z(n6723) );
  XOR U6793 ( .A(n6326), .B(n6727), .Z(n6717) );
  XOR U6794 ( .A(n2494), .B(n6258), .Z(n6727) );
  XOR U6795 ( .A(n6728), .B(n6729), .Z(n6258) );
  NOR U6796 ( .A(n6730), .B(n6731), .Z(n6728) );
  XNOR U6797 ( .A(n6732), .B(n6733), .Z(n2494) );
  XNOR U6798 ( .A(n6736), .B(n6737), .Z(n6326) );
  ANDN U6799 ( .B(n6738), .A(n6739), .Z(n6736) );
  XOR U6800 ( .A(n6740), .B(n5800), .Z(out[1073]) );
  XNOR U6801 ( .A(n6741), .B(n2633), .Z(n5800) );
  XOR U6802 ( .A(n6742), .B(n5912), .Z(n2633) );
  XNOR U6803 ( .A(n6743), .B(n6744), .Z(n5912) );
  XNOR U6804 ( .A(n5535), .B(n3674), .Z(n6744) );
  XOR U6805 ( .A(n6745), .B(n6746), .Z(n3674) );
  AND U6806 ( .A(n6747), .B(n6748), .Z(n6745) );
  XNOR U6807 ( .A(n6749), .B(n6750), .Z(n5535) );
  NOR U6808 ( .A(n6751), .B(n6752), .Z(n6749) );
  XNOR U6809 ( .A(n6330), .B(n6753), .Z(n6743) );
  XOR U6810 ( .A(n2501), .B(n6309), .Z(n6753) );
  XNOR U6811 ( .A(n6754), .B(n6755), .Z(n6309) );
  AND U6812 ( .A(n6756), .B(n6757), .Z(n6754) );
  XOR U6813 ( .A(n6758), .B(n6759), .Z(n2501) );
  ANDN U6814 ( .B(n6760), .A(n6761), .Z(n6758) );
  XNOR U6815 ( .A(n6762), .B(n6763), .Z(n6330) );
  ANDN U6816 ( .B(n6764), .A(n6765), .Z(n6762) );
  ANDN U6817 ( .B(n6766), .A(n5619), .Z(n6740) );
  XOR U6818 ( .A(n6767), .B(n5802), .Z(out[1072]) );
  XNOR U6819 ( .A(n6768), .B(n5329), .Z(n5802) );
  XOR U6820 ( .A(n6769), .B(n5917), .Z(n5329) );
  XNOR U6821 ( .A(n6770), .B(n6771), .Z(n5917) );
  XOR U6822 ( .A(n5539), .B(n3681), .Z(n6771) );
  XOR U6823 ( .A(n6772), .B(n6773), .Z(n3681) );
  ANDN U6824 ( .B(n6774), .A(n6775), .Z(n6772) );
  XNOR U6825 ( .A(n6776), .B(n6777), .Z(n5539) );
  XOR U6826 ( .A(n6778), .B(n6779), .Z(n6777) );
  NAND U6827 ( .A(n4509), .B(n6454), .Z(n6779) );
  XOR U6828 ( .A(n6334), .B(n6782), .Z(n6770) );
  XNOR U6829 ( .A(n2508), .B(n6346), .Z(n6782) );
  XNOR U6830 ( .A(n6783), .B(n6784), .Z(n6346) );
  AND U6831 ( .A(n6785), .B(n6786), .Z(n6783) );
  XOR U6832 ( .A(n6787), .B(n6788), .Z(n2508) );
  ANDN U6833 ( .B(n6789), .A(n6790), .Z(n6787) );
  XNOR U6834 ( .A(n6791), .B(n6792), .Z(n6334) );
  AND U6835 ( .A(n6793), .B(n6794), .Z(n6791) );
  AND U6836 ( .A(n5623), .B(n6795), .Z(n6767) );
  XOR U6837 ( .A(n6796), .B(n5812), .Z(out[1071]) );
  XNOR U6838 ( .A(n6797), .B(n5334), .Z(n5812) );
  XOR U6839 ( .A(n6798), .B(n5922), .Z(n5334) );
  XNOR U6840 ( .A(n6799), .B(n6800), .Z(n5922) );
  XNOR U6841 ( .A(n5543), .B(n3686), .Z(n6800) );
  XOR U6842 ( .A(n6801), .B(n6802), .Z(n3686) );
  AND U6843 ( .A(n6803), .B(n6804), .Z(n6801) );
  XNOR U6844 ( .A(n6805), .B(n6806), .Z(n5543) );
  ANDN U6845 ( .B(n6807), .A(n6808), .Z(n6805) );
  XOR U6846 ( .A(n6336), .B(n6809), .Z(n6799) );
  XOR U6847 ( .A(n2515), .B(n6573), .Z(n6809) );
  XOR U6848 ( .A(n6810), .B(n6811), .Z(n6573) );
  XOR U6849 ( .A(n6814), .B(n6815), .Z(n2515) );
  ANDN U6850 ( .B(n6816), .A(n6817), .Z(n6814) );
  XNOR U6851 ( .A(n6818), .B(n6819), .Z(n6336) );
  NOR U6852 ( .A(n6820), .B(n6821), .Z(n6818) );
  ANDN U6853 ( .B(n5627), .A(n6139), .Z(n6796) );
  XOR U6854 ( .A(n6822), .B(n5815), .Z(out[1070]) );
  XOR U6855 ( .A(n6823), .B(n5365), .Z(n5815) );
  XOR U6856 ( .A(n6824), .B(n5927), .Z(n5365) );
  XNOR U6857 ( .A(n6825), .B(n6826), .Z(n5927) );
  XOR U6858 ( .A(n5547), .B(n3692), .Z(n6826) );
  XOR U6859 ( .A(n6827), .B(n6828), .Z(n3692) );
  XNOR U6860 ( .A(n6831), .B(n6832), .Z(n5547) );
  XOR U6861 ( .A(n6833), .B(n6834), .Z(n6832) );
  NAND U6862 ( .A(n6835), .B(n6836), .Z(n6834) );
  ANDN U6863 ( .B(n6837), .A(n6838), .Z(n6833) );
  XOR U6864 ( .A(n6338), .B(n6839), .Z(n6825) );
  XOR U6865 ( .A(n2526), .B(n6840), .Z(n6839) );
  XOR U6866 ( .A(n6841), .B(n6842), .Z(n2526) );
  ANDN U6867 ( .B(n6843), .A(n6844), .Z(n6841) );
  XOR U6868 ( .A(n6845), .B(n6846), .Z(n6338) );
  AND U6869 ( .A(n6847), .B(n6848), .Z(n6845) );
  NOR U6870 ( .A(n6144), .B(n5631), .Z(n6822) );
  XNOR U6871 ( .A(n6849), .B(n4142), .Z(out[106]) );
  XNOR U6872 ( .A(n6840), .B(n2527), .Z(n4142) );
  XNOR U6873 ( .A(n6850), .B(n6851), .Z(n2527) );
  XNOR U6874 ( .A(n6852), .B(n6853), .Z(n6840) );
  AND U6875 ( .A(n6854), .B(n6855), .Z(n6852) );
  NOR U6876 ( .A(n3420), .B(n3419), .Z(n6849) );
  XNOR U6877 ( .A(n6856), .B(n2363), .Z(n3419) );
  XNOR U6878 ( .A(n6857), .B(n2296), .Z(n3420) );
  XOR U6879 ( .A(n6858), .B(n5818), .Z(out[1069]) );
  XNOR U6880 ( .A(n6859), .B(n2661), .Z(n5818) );
  XOR U6881 ( .A(n6860), .B(n5932), .Z(n2661) );
  XNOR U6882 ( .A(n6861), .B(n6862), .Z(n5932) );
  XOR U6883 ( .A(n5552), .B(n3696), .Z(n6862) );
  XOR U6884 ( .A(n6863), .B(n6864), .Z(n3696) );
  AND U6885 ( .A(n6865), .B(n6866), .Z(n6863) );
  XNOR U6886 ( .A(n6867), .B(n6868), .Z(n5552) );
  XOR U6887 ( .A(n6869), .B(n6870), .Z(n6868) );
  ANDN U6888 ( .B(n6871), .A(n6872), .Z(n6869) );
  XNOR U6889 ( .A(n6340), .B(n6873), .Z(n6861) );
  XOR U6890 ( .A(n2533), .B(n6874), .Z(n6873) );
  XOR U6891 ( .A(n6875), .B(n6876), .Z(n2533) );
  AND U6892 ( .A(n6877), .B(n6878), .Z(n6875) );
  XNOR U6893 ( .A(n6879), .B(n6880), .Z(n6340) );
  ANDN U6894 ( .B(n6881), .A(n6882), .Z(n6879) );
  ANDN U6895 ( .B(n5635), .A(n6149), .Z(n6858) );
  XOR U6896 ( .A(n6883), .B(n5820), .Z(out[1068]) );
  XNOR U6897 ( .A(n6884), .B(n5468), .Z(n5820) );
  XOR U6898 ( .A(n6885), .B(n5937), .Z(n5468) );
  XNOR U6899 ( .A(n6886), .B(n6887), .Z(n5937) );
  XNOR U6900 ( .A(n5247), .B(n3700), .Z(n6887) );
  XOR U6901 ( .A(n6888), .B(n6889), .Z(n3700) );
  XNOR U6902 ( .A(n6892), .B(n6893), .Z(n5247) );
  XOR U6903 ( .A(n6894), .B(n6677), .Z(n6893) );
  NAND U6904 ( .A(n6835), .B(n4656), .Z(n6677) );
  XNOR U6905 ( .A(n6343), .B(n6897), .Z(n6886) );
  XNOR U6906 ( .A(n2540), .B(n6898), .Z(n6897) );
  XOR U6907 ( .A(n6899), .B(n6900), .Z(n2540) );
  XNOR U6908 ( .A(n6903), .B(n6904), .Z(n6343) );
  ANDN U6909 ( .B(n6905), .A(n6906), .Z(n6903) );
  AND U6910 ( .A(n5639), .B(n6907), .Z(n6883) );
  XNOR U6911 ( .A(n6908), .B(n5822), .Z(out[1067]) );
  XOR U6912 ( .A(n3331), .B(n6909), .Z(n5822) );
  IV U6913 ( .A(n2200), .Z(n3331) );
  AND U6914 ( .A(n5648), .B(n6910), .Z(n6908) );
  XNOR U6915 ( .A(n6911), .B(n5824), .Z(out[1066]) );
  XNOR U6916 ( .A(n2207), .B(n6912), .Z(n5824) );
  IV U6917 ( .A(n5555), .Z(n2207) );
  XOR U6918 ( .A(n6913), .B(n5947), .Z(n5555) );
  XNOR U6919 ( .A(n6914), .B(n6915), .Z(n5947) );
  XOR U6920 ( .A(n5254), .B(n3709), .Z(n6915) );
  XOR U6921 ( .A(n6916), .B(n6917), .Z(n3709) );
  AND U6922 ( .A(n6918), .B(n6919), .Z(n6916) );
  XNOR U6923 ( .A(n6920), .B(n6921), .Z(n5254) );
  ANDN U6924 ( .B(n6922), .A(n6923), .Z(n6920) );
  XNOR U6925 ( .A(n6355), .B(n6924), .Z(n6914) );
  XOR U6926 ( .A(n2554), .B(n6925), .Z(n6924) );
  XOR U6927 ( .A(n6926), .B(n6927), .Z(n2554) );
  AND U6928 ( .A(n6928), .B(n6929), .Z(n6926) );
  XOR U6929 ( .A(n6930), .B(n6931), .Z(n6355) );
  AND U6930 ( .A(n6932), .B(n6933), .Z(n6930) );
  AND U6931 ( .A(n5652), .B(n6934), .Z(n6911) );
  XOR U6932 ( .A(n6935), .B(n5826), .Z(out[1065]) );
  XNOR U6933 ( .A(n3339), .B(n6936), .Z(n5826) );
  XNOR U6934 ( .A(n6937), .B(n5957), .Z(n3339) );
  XNOR U6935 ( .A(n6938), .B(n6939), .Z(n5957) );
  XOR U6936 ( .A(n5258), .B(n3713), .Z(n6939) );
  XOR U6937 ( .A(n6940), .B(n6941), .Z(n3713) );
  ANDN U6938 ( .B(n6942), .A(n6943), .Z(n6940) );
  XNOR U6939 ( .A(n6944), .B(n6945), .Z(n5258) );
  AND U6940 ( .A(n6946), .B(n6947), .Z(n6944) );
  XNOR U6941 ( .A(n6051), .B(n6948), .Z(n6938) );
  XNOR U6942 ( .A(n2561), .B(n6949), .Z(n6948) );
  XNOR U6943 ( .A(n6950), .B(n6951), .Z(n2561) );
  AND U6944 ( .A(n6952), .B(n6953), .Z(n6950) );
  XNOR U6945 ( .A(n6954), .B(n6955), .Z(n6051) );
  NOR U6946 ( .A(n6956), .B(n6957), .Z(n6954) );
  ANDN U6947 ( .B(n6173), .A(n5656), .Z(n6935) );
  XOR U6948 ( .A(n6958), .B(n5828), .Z(out[1064]) );
  XOR U6949 ( .A(n2221), .B(n6959), .Z(n5828) );
  XNOR U6950 ( .A(n6960), .B(n5962), .Z(n2221) );
  XNOR U6951 ( .A(n6961), .B(n6962), .Z(n5962) );
  XNOR U6952 ( .A(n5268), .B(n3716), .Z(n6962) );
  XNOR U6953 ( .A(n6963), .B(n6964), .Z(n3716) );
  AND U6954 ( .A(n6965), .B(n6966), .Z(n6963) );
  XNOR U6955 ( .A(n6967), .B(n6968), .Z(n5268) );
  AND U6956 ( .A(n6969), .B(n6970), .Z(n6967) );
  XNOR U6957 ( .A(n6054), .B(n6971), .Z(n6961) );
  XNOR U6958 ( .A(n2568), .B(n6972), .Z(n6971) );
  XNOR U6959 ( .A(n6973), .B(n6974), .Z(n2568) );
  AND U6960 ( .A(n6975), .B(n6976), .Z(n6973) );
  XOR U6961 ( .A(n6977), .B(n6978), .Z(n6054) );
  ANDN U6962 ( .B(n6979), .A(n6980), .Z(n6977) );
  ANDN U6963 ( .B(n5660), .A(n6178), .Z(n6958) );
  XOR U6964 ( .A(n6981), .B(n5833), .Z(out[1063]) );
  XOR U6965 ( .A(n2232), .B(n6982), .Z(n5833) );
  IV U6966 ( .A(n5677), .Z(n2232) );
  XOR U6967 ( .A(n6983), .B(n5967), .Z(n5677) );
  XNOR U6968 ( .A(n6984), .B(n6985), .Z(n5967) );
  XNOR U6969 ( .A(n5271), .B(n3720), .Z(n6985) );
  XNOR U6970 ( .A(n6986), .B(n6987), .Z(n3720) );
  AND U6971 ( .A(n6988), .B(n6989), .Z(n6986) );
  XOR U6972 ( .A(n6990), .B(n6991), .Z(n5271) );
  ANDN U6973 ( .B(n6992), .A(n6993), .Z(n6990) );
  XNOR U6974 ( .A(n6061), .B(n6994), .Z(n6984) );
  XOR U6975 ( .A(n4334), .B(n2576), .Z(n6994) );
  XOR U6976 ( .A(n6995), .B(n6996), .Z(n2576) );
  XOR U6977 ( .A(n6999), .B(n7000), .Z(n4334) );
  ANDN U6978 ( .B(n7001), .A(n7002), .Z(n6999) );
  XOR U6979 ( .A(n7003), .B(n7004), .Z(n6061) );
  ANDN U6980 ( .B(n7005), .A(n7006), .Z(n7003) );
  ANDN U6981 ( .B(n1042), .A(n1044), .Z(n6981) );
  XNOR U6982 ( .A(n3860), .B(n7007), .Z(n1044) );
  IV U6983 ( .A(n1792), .Z(n3860) );
  XOR U6984 ( .A(n6520), .B(n6298), .Z(n1792) );
  XOR U6985 ( .A(n7008), .B(n7009), .Z(n6298) );
  XNOR U6986 ( .A(n5880), .B(n2129), .Z(n7009) );
  XOR U6987 ( .A(n7010), .B(n7011), .Z(n2129) );
  XOR U6988 ( .A(n7012), .B(n7013), .Z(n5880) );
  ANDN U6989 ( .B(n6584), .A(n6585), .Z(n7012) );
  XNOR U6990 ( .A(n5440), .B(n7014), .Z(n7008) );
  XOR U6991 ( .A(n4297), .B(n3691), .Z(n7014) );
  XOR U6992 ( .A(n7015), .B(n7016), .Z(n3691) );
  ANDN U6993 ( .B(n7017), .A(n6588), .Z(n7015) );
  XOR U6994 ( .A(n7018), .B(n7019), .Z(n4297) );
  AND U6995 ( .A(n6601), .B(n6603), .Z(n7018) );
  XOR U6996 ( .A(n7020), .B(n7021), .Z(n5440) );
  AND U6997 ( .A(n6599), .B(n6597), .Z(n7020) );
  XOR U6998 ( .A(n7022), .B(n7023), .Z(n6520) );
  XOR U6999 ( .A(n3475), .B(n4862), .Z(n7023) );
  XNOR U7000 ( .A(n7024), .B(n6569), .Z(n4862) );
  ANDN U7001 ( .B(n7025), .A(n7026), .Z(n7024) );
  XOR U7002 ( .A(n7027), .B(n6561), .Z(n3475) );
  AND U7003 ( .A(n7028), .B(n7029), .Z(n7027) );
  XOR U7004 ( .A(n7030), .B(n7031), .Z(n7022) );
  XNOR U7005 ( .A(n4032), .B(n2545), .Z(n7031) );
  XOR U7006 ( .A(n7032), .B(n6552), .Z(n2545) );
  XOR U7007 ( .A(n7035), .B(n6556), .Z(n4032) );
  XOR U7008 ( .A(n3382), .B(n7038), .Z(n1042) );
  XOR U7009 ( .A(n7039), .B(n5838), .Z(out[1062]) );
  XNOR U7010 ( .A(n7040), .B(n2242), .Z(n5838) );
  XOR U7011 ( .A(n7041), .B(n5972), .Z(n2242) );
  XNOR U7012 ( .A(n7042), .B(n7043), .Z(n5972) );
  XNOR U7013 ( .A(n5276), .B(n3726), .Z(n7043) );
  XOR U7014 ( .A(n7044), .B(n7045), .Z(n3726) );
  ANDN U7015 ( .B(n7046), .A(n7047), .Z(n7044) );
  XOR U7016 ( .A(n7048), .B(n7049), .Z(n5276) );
  AND U7017 ( .A(n7050), .B(n7051), .Z(n7048) );
  XOR U7018 ( .A(n6066), .B(n7052), .Z(n7042) );
  XNOR U7019 ( .A(n4340), .B(n2583), .Z(n7052) );
  XOR U7020 ( .A(n7053), .B(n7054), .Z(n2583) );
  AND U7021 ( .A(n7055), .B(n7056), .Z(n7053) );
  XOR U7022 ( .A(n7057), .B(n7058), .Z(n4340) );
  AND U7023 ( .A(n7059), .B(n7060), .Z(n7057) );
  XOR U7024 ( .A(n7061), .B(n7062), .Z(n6066) );
  ANDN U7025 ( .B(n7063), .A(n7064), .Z(n7061) );
  AND U7026 ( .A(n1046), .B(n1048), .Z(n7039) );
  XOR U7027 ( .A(n7065), .B(n1797), .Z(n1048) );
  XOR U7028 ( .A(n6547), .B(n6302), .Z(n1797) );
  XOR U7029 ( .A(n7066), .B(n7067), .Z(n6302) );
  XNOR U7030 ( .A(n5445), .B(n4299), .Z(n7067) );
  XOR U7031 ( .A(n7068), .B(n7069), .Z(n4299) );
  ANDN U7032 ( .B(n6631), .A(n6629), .Z(n7068) );
  XNOR U7033 ( .A(n7070), .B(n7071), .Z(n5445) );
  ANDN U7034 ( .B(n6625), .A(n6626), .Z(n7070) );
  XOR U7035 ( .A(n3697), .B(n7072), .Z(n7066) );
  XOR U7036 ( .A(n5885), .B(n2132), .Z(n7072) );
  XNOR U7037 ( .A(n7073), .B(n7074), .Z(n2132) );
  ANDN U7038 ( .B(n6623), .A(n6621), .Z(n7073) );
  XNOR U7039 ( .A(n7075), .B(n7076), .Z(n5885) );
  ANDN U7040 ( .B(n6612), .A(n6613), .Z(n7075) );
  XNOR U7041 ( .A(n7077), .B(n7078), .Z(n3697) );
  ANDN U7042 ( .B(n6616), .A(n6617), .Z(n7077) );
  XOR U7043 ( .A(n7079), .B(n7080), .Z(n6547) );
  XNOR U7044 ( .A(n4865), .B(n4035), .Z(n7080) );
  XOR U7045 ( .A(n7081), .B(n6589), .Z(n4035) );
  IV U7046 ( .A(n7082), .Z(n6589) );
  NOR U7047 ( .A(n7016), .B(n7083), .Z(n7081) );
  XNOR U7048 ( .A(n7084), .B(n6602), .Z(n4865) );
  NOR U7049 ( .A(n7085), .B(n7019), .Z(n7084) );
  XOR U7050 ( .A(n2551), .B(n7086), .Z(n7079) );
  XNOR U7051 ( .A(n3481), .B(n7087), .Z(n7086) );
  XNOR U7052 ( .A(n7088), .B(n6594), .Z(n3481) );
  ANDN U7053 ( .B(n7011), .A(n7089), .Z(n7088) );
  XOR U7054 ( .A(n7090), .B(n6586), .Z(n2551) );
  IV U7055 ( .A(n7091), .Z(n6586) );
  ANDN U7056 ( .B(n7092), .A(n7013), .Z(n7090) );
  XNOR U7057 ( .A(n4983), .B(n7093), .Z(n1046) );
  IV U7058 ( .A(n2320), .Z(n4983) );
  XOR U7059 ( .A(n7094), .B(n5848), .Z(out[1061]) );
  XOR U7060 ( .A(n7095), .B(n5729), .Z(n5848) );
  XOR U7061 ( .A(n7096), .B(n5977), .Z(n5729) );
  XNOR U7062 ( .A(n7097), .B(n7098), .Z(n5977) );
  XOR U7063 ( .A(n5284), .B(n3732), .Z(n7098) );
  XOR U7064 ( .A(n7099), .B(n7100), .Z(n3732) );
  AND U7065 ( .A(n7101), .B(n7102), .Z(n7099) );
  XNOR U7066 ( .A(n7103), .B(n7104), .Z(n5284) );
  AND U7067 ( .A(n7105), .B(n7106), .Z(n7103) );
  XNOR U7068 ( .A(n6071), .B(n7107), .Z(n7097) );
  XOR U7069 ( .A(n4344), .B(n2590), .Z(n7107) );
  XNOR U7070 ( .A(n7108), .B(n7109), .Z(n2590) );
  AND U7071 ( .A(n7110), .B(n7111), .Z(n7108) );
  XOR U7072 ( .A(n7112), .B(n7113), .Z(n4344) );
  ANDN U7073 ( .B(n7114), .A(n7115), .Z(n7112) );
  XOR U7074 ( .A(n7116), .B(n7117), .Z(n6071) );
  AND U7075 ( .A(n7118), .B(n7119), .Z(n7116) );
  AND U7076 ( .A(n1052), .B(n1050), .Z(n7094) );
  XNOR U7077 ( .A(n2329), .B(n7120), .Z(n1050) );
  XNOR U7078 ( .A(n1800), .B(n7121), .Z(n1052) );
  XOR U7079 ( .A(n7122), .B(n5853), .Z(out[1060]) );
  XNOR U7080 ( .A(n7123), .B(n2256), .Z(n5853) );
  XOR U7081 ( .A(n7124), .B(n5981), .Z(n2256) );
  XNOR U7082 ( .A(n7125), .B(n7126), .Z(n5981) );
  XOR U7083 ( .A(n5288), .B(n3738), .Z(n7126) );
  XOR U7084 ( .A(n7127), .B(n7128), .Z(n3738) );
  AND U7085 ( .A(n7129), .B(n7130), .Z(n7127) );
  XNOR U7086 ( .A(n7131), .B(n7132), .Z(n5288) );
  AND U7087 ( .A(n7133), .B(n7134), .Z(n7131) );
  XNOR U7088 ( .A(n6076), .B(n7135), .Z(n7125) );
  XNOR U7089 ( .A(n2600), .B(n4350), .Z(n7135) );
  XNOR U7090 ( .A(n7136), .B(n7137), .Z(n4350) );
  AND U7091 ( .A(n7138), .B(n7139), .Z(n7136) );
  XNOR U7092 ( .A(n7140), .B(n7141), .Z(n2600) );
  ANDN U7093 ( .B(n7142), .A(n7143), .Z(n7140) );
  XOR U7094 ( .A(n7144), .B(n7145), .Z(n6076) );
  ANDN U7095 ( .B(n7146), .A(n7147), .Z(n7144) );
  ANDN U7096 ( .B(n1054), .A(n1055), .Z(n7122) );
  XOR U7097 ( .A(n1804), .B(n7148), .Z(n1055) );
  XNOR U7098 ( .A(n6608), .B(n6319), .Z(n1804) );
  XOR U7099 ( .A(n7149), .B(n7150), .Z(n6319) );
  XNOR U7100 ( .A(n5900), .B(n4304), .Z(n7150) );
  XNOR U7101 ( .A(n7151), .B(n7152), .Z(n4304) );
  AND U7102 ( .A(n6671), .B(n7153), .Z(n7151) );
  XNOR U7103 ( .A(n7154), .B(n7155), .Z(n5900) );
  AND U7104 ( .A(n6685), .B(n6687), .Z(n7154) );
  XOR U7105 ( .A(n3705), .B(n7156), .Z(n7149) );
  XNOR U7106 ( .A(n5454), .B(n2141), .Z(n7156) );
  XNOR U7107 ( .A(n7157), .B(n7158), .Z(n2141) );
  XOR U7108 ( .A(n7159), .B(n7160), .Z(n5454) );
  NOR U7109 ( .A(n6667), .B(n6666), .Z(n7159) );
  XNOR U7110 ( .A(n7161), .B(n7162), .Z(n3705) );
  AND U7111 ( .A(n6674), .B(n6679), .Z(n7161) );
  XOR U7112 ( .A(n7163), .B(n7164), .Z(n6608) );
  XNOR U7113 ( .A(n4875), .B(n4042), .Z(n7164) );
  XNOR U7114 ( .A(n7165), .B(n6645), .Z(n4042) );
  ANDN U7115 ( .B(n7166), .A(n7167), .Z(n7165) );
  XOR U7116 ( .A(n7168), .B(n6658), .Z(n4875) );
  IV U7117 ( .A(n7169), .Z(n6658) );
  NOR U7118 ( .A(n7170), .B(n7171), .Z(n7168) );
  XNOR U7119 ( .A(n2563), .B(n7172), .Z(n7163) );
  XNOR U7120 ( .A(n3486), .B(n7173), .Z(n7172) );
  XNOR U7121 ( .A(n7174), .B(n6650), .Z(n3486) );
  ANDN U7122 ( .B(n7175), .A(n7176), .Z(n7174) );
  XNOR U7123 ( .A(n7177), .B(n7178), .Z(n2563) );
  ANDN U7124 ( .B(n7179), .A(n7180), .Z(n7177) );
  XNOR U7125 ( .A(n2336), .B(n7181), .Z(n1054) );
  XOR U7126 ( .A(n7182), .B(n4146), .Z(out[105]) );
  IV U7127 ( .A(n4320), .Z(n4146) );
  XOR U7128 ( .A(n6874), .B(n2534), .Z(n4320) );
  XNOR U7129 ( .A(n7183), .B(n7184), .Z(n2534) );
  XNOR U7130 ( .A(n7185), .B(n7186), .Z(n6874) );
  AND U7131 ( .A(n7187), .B(n7188), .Z(n7185) );
  ANDN U7132 ( .B(n3448), .A(n3449), .Z(n7182) );
  XNOR U7133 ( .A(n7189), .B(n2307), .Z(n3449) );
  XOR U7134 ( .A(n7190), .B(n2372), .Z(n3448) );
  XNOR U7135 ( .A(n7191), .B(n5858), .Z(out[1059]) );
  XNOR U7136 ( .A(n7192), .B(n3367), .Z(n5858) );
  XOR U7137 ( .A(n7193), .B(n5986), .Z(n3367) );
  XNOR U7138 ( .A(n7194), .B(n7195), .Z(n5986) );
  XOR U7139 ( .A(n5293), .B(n3741), .Z(n7195) );
  XOR U7140 ( .A(n7196), .B(n7197), .Z(n3741) );
  XNOR U7141 ( .A(n7200), .B(n7201), .Z(n5293) );
  AND U7142 ( .A(n7202), .B(n7203), .Z(n7200) );
  XNOR U7143 ( .A(n6081), .B(n7204), .Z(n7194) );
  XOR U7144 ( .A(n2607), .B(n4358), .Z(n7204) );
  XNOR U7145 ( .A(n7205), .B(n7206), .Z(n4358) );
  NOR U7146 ( .A(n7207), .B(n7208), .Z(n7205) );
  XNOR U7147 ( .A(n7209), .B(n7210), .Z(n2607) );
  NOR U7148 ( .A(n7211), .B(n7212), .Z(n7209) );
  XNOR U7149 ( .A(n7213), .B(n7214), .Z(n6081) );
  AND U7150 ( .A(n1060), .B(n1058), .Z(n7191) );
  XNOR U7151 ( .A(n2341), .B(n7217), .Z(n1058) );
  IV U7152 ( .A(n3398), .Z(n2341) );
  XNOR U7153 ( .A(n1808), .B(n7218), .Z(n1060) );
  IV U7154 ( .A(n5158), .Z(n1808) );
  XOR U7155 ( .A(n6635), .B(n6323), .Z(n5158) );
  XOR U7156 ( .A(n7219), .B(n7220), .Z(n6323) );
  XNOR U7157 ( .A(n5905), .B(n4306), .Z(n7220) );
  XOR U7158 ( .A(n7221), .B(n7222), .Z(n4306) );
  NOR U7159 ( .A(n6711), .B(n6712), .Z(n7221) );
  XOR U7160 ( .A(n7223), .B(n7224), .Z(n5905) );
  ANDN U7161 ( .B(n7225), .A(n6694), .Z(n7223) );
  XOR U7162 ( .A(n3708), .B(n7226), .Z(n7219) );
  XNOR U7163 ( .A(n5458), .B(n2145), .Z(n7226) );
  XNOR U7164 ( .A(n7227), .B(n7228), .Z(n2145) );
  XNOR U7165 ( .A(n7229), .B(n7230), .Z(n5458) );
  AND U7166 ( .A(n6707), .B(n6709), .Z(n7229) );
  XNOR U7167 ( .A(n7231), .B(n7232), .Z(n3708) );
  ANDN U7168 ( .B(n6700), .A(n6698), .Z(n7231) );
  XOR U7169 ( .A(n7233), .B(n7234), .Z(n6635) );
  XOR U7170 ( .A(n4878), .B(n4045), .Z(n7234) );
  XOR U7171 ( .A(n7235), .B(n7236), .Z(n4045) );
  NOR U7172 ( .A(n7162), .B(n7237), .Z(n7235) );
  XNOR U7173 ( .A(n7238), .B(n6672), .Z(n4878) );
  ANDN U7174 ( .B(n7239), .A(n7152), .Z(n7238) );
  XNOR U7175 ( .A(n2572), .B(n7240), .Z(n7233) );
  XOR U7176 ( .A(n3490), .B(n7241), .Z(n7240) );
  XNOR U7177 ( .A(n7242), .B(n6683), .Z(n3490) );
  NOR U7178 ( .A(n7243), .B(n7158), .Z(n7242) );
  XNOR U7179 ( .A(n7244), .B(n6686), .Z(n2572) );
  XNOR U7180 ( .A(n7246), .B(n5863), .Z(out[1058]) );
  XOR U7181 ( .A(n7247), .B(n5398), .Z(n5863) );
  XOR U7182 ( .A(n7248), .B(n5991), .Z(n5398) );
  XNOR U7183 ( .A(n7249), .B(n7250), .Z(n5991) );
  XNOR U7184 ( .A(n5296), .B(n3747), .Z(n7250) );
  XOR U7185 ( .A(n7251), .B(n7252), .Z(n3747) );
  XNOR U7186 ( .A(n7255), .B(n7256), .Z(n5296) );
  XNOR U7187 ( .A(n6086), .B(n7259), .Z(n7249) );
  XOR U7188 ( .A(n2614), .B(n4407), .Z(n7259) );
  XNOR U7189 ( .A(n7260), .B(n7261), .Z(n4407) );
  NOR U7190 ( .A(n7262), .B(n7263), .Z(n7260) );
  XNOR U7191 ( .A(n7264), .B(n7265), .Z(n2614) );
  AND U7192 ( .A(n7266), .B(n7267), .Z(n7264) );
  XNOR U7193 ( .A(n7268), .B(n7269), .Z(n6086) );
  ANDN U7194 ( .B(n7270), .A(n7271), .Z(n7268) );
  ANDN U7195 ( .B(n1062), .A(n1064), .Z(n7246) );
  XNOR U7196 ( .A(n1820), .B(n7272), .Z(n1064) );
  IV U7197 ( .A(n5161), .Z(n1820) );
  XOR U7198 ( .A(n6662), .B(n6327), .Z(n5161) );
  XOR U7199 ( .A(n7273), .B(n7274), .Z(n6327) );
  XNOR U7200 ( .A(n5910), .B(n5471), .Z(n7274) );
  XOR U7201 ( .A(n7275), .B(n7276), .Z(n5471) );
  NOR U7202 ( .A(n6734), .B(n6733), .Z(n7275) );
  IV U7203 ( .A(n7277), .Z(n6734) );
  XNOR U7204 ( .A(n7278), .B(n7279), .Z(n5910) );
  ANDN U7205 ( .B(n6720), .A(n6721), .Z(n7278) );
  XOR U7206 ( .A(n3712), .B(n7280), .Z(n7273) );
  XNOR U7207 ( .A(n4309), .B(n2148), .Z(n7280) );
  XNOR U7208 ( .A(n7281), .B(n7282), .Z(n2148) );
  AND U7209 ( .A(n6729), .B(n6730), .Z(n7281) );
  XOR U7210 ( .A(n7283), .B(n7284), .Z(n4309) );
  NOR U7211 ( .A(n6737), .B(n6738), .Z(n7283) );
  XOR U7212 ( .A(n7285), .B(n7286), .Z(n3712) );
  NOR U7213 ( .A(n6725), .B(n6724), .Z(n7285) );
  XOR U7214 ( .A(n7287), .B(n7288), .Z(n6662) );
  XNOR U7215 ( .A(n4881), .B(n4048), .Z(n7288) );
  XOR U7216 ( .A(n7289), .B(n6699), .Z(n4048) );
  IV U7217 ( .A(n7290), .Z(n6699) );
  NOR U7218 ( .A(n7291), .B(n7232), .Z(n7289) );
  XNOR U7219 ( .A(n7292), .B(n6713), .Z(n4881) );
  ANDN U7220 ( .B(n7222), .A(n7293), .Z(n7292) );
  XOR U7221 ( .A(n2577), .B(n7294), .Z(n7287) );
  XOR U7222 ( .A(n3493), .B(n7295), .Z(n7294) );
  XNOR U7223 ( .A(n7296), .B(n6705), .Z(n3493) );
  ANDN U7224 ( .B(n7297), .A(n7228), .Z(n7296) );
  XOR U7225 ( .A(n7298), .B(n6696), .Z(n2577) );
  AND U7226 ( .A(n7224), .B(n7299), .Z(n7298) );
  XNOR U7227 ( .A(n2350), .B(n7300), .Z(n1062) );
  XOR U7228 ( .A(n6171), .B(n7301), .Z(n2350) );
  XOR U7229 ( .A(n7302), .B(n7303), .Z(n6171) );
  XOR U7230 ( .A(n3185), .B(n7304), .Z(n7303) );
  XOR U7231 ( .A(n7305), .B(n7306), .Z(n3185) );
  ANDN U7232 ( .B(n7307), .A(n7308), .Z(n7305) );
  XNOR U7233 ( .A(n5480), .B(n7309), .Z(n7302) );
  XOR U7234 ( .A(n7310), .B(n2389), .Z(n7309) );
  XNOR U7235 ( .A(n7311), .B(n7312), .Z(n2389) );
  AND U7236 ( .A(n7313), .B(n7314), .Z(n7311) );
  XNOR U7237 ( .A(n7315), .B(n7316), .Z(n5480) );
  AND U7238 ( .A(n7317), .B(n7318), .Z(n7315) );
  XNOR U7239 ( .A(n7319), .B(n5868), .Z(out[1057]) );
  XNOR U7240 ( .A(n7320), .B(n2277), .Z(n5868) );
  XNOR U7241 ( .A(n7321), .B(n5996), .Z(n2277) );
  XNOR U7242 ( .A(n7322), .B(n7323), .Z(n5996) );
  XOR U7243 ( .A(n5301), .B(n3752), .Z(n7323) );
  XOR U7244 ( .A(n7324), .B(n7325), .Z(n3752) );
  AND U7245 ( .A(n7326), .B(n7327), .Z(n7324) );
  XNOR U7246 ( .A(n7328), .B(n7329), .Z(n5301) );
  XOR U7247 ( .A(n6091), .B(n7332), .Z(n7322) );
  XOR U7248 ( .A(n2621), .B(n4450), .Z(n7332) );
  XOR U7249 ( .A(n7333), .B(n7334), .Z(n4450) );
  NOR U7250 ( .A(n7335), .B(n7336), .Z(n7333) );
  XNOR U7251 ( .A(n7337), .B(n7338), .Z(n2621) );
  ANDN U7252 ( .B(n7339), .A(n7340), .Z(n7337) );
  XNOR U7253 ( .A(n7341), .B(n7342), .Z(n6091) );
  AND U7254 ( .A(n7343), .B(n7344), .Z(n7341) );
  ANDN U7255 ( .B(n1066), .A(n1068), .Z(n7319) );
  XNOR U7256 ( .A(n1824), .B(n7345), .Z(n1068) );
  IV U7257 ( .A(n3561), .Z(n1824) );
  XOR U7258 ( .A(n6690), .B(n6331), .Z(n3561) );
  XOR U7259 ( .A(n7346), .B(n7347), .Z(n6331) );
  XNOR U7260 ( .A(n5915), .B(n5475), .Z(n7347) );
  XNOR U7261 ( .A(n7348), .B(n7349), .Z(n5475) );
  XNOR U7262 ( .A(n7350), .B(n7351), .Z(n5915) );
  AND U7263 ( .A(n6746), .B(n7352), .Z(n7350) );
  IV U7264 ( .A(n7353), .Z(n6746) );
  XOR U7265 ( .A(n3717), .B(n7354), .Z(n7346) );
  XOR U7266 ( .A(n4311), .B(n2151), .Z(n7354) );
  XNOR U7267 ( .A(n7355), .B(n7356), .Z(n2151) );
  NOR U7268 ( .A(n6755), .B(n6756), .Z(n7355) );
  XOR U7269 ( .A(n7357), .B(n7358), .Z(n4311) );
  ANDN U7270 ( .B(n7359), .A(n6763), .Z(n7357) );
  XNOR U7271 ( .A(n7360), .B(n7361), .Z(n3717) );
  AND U7272 ( .A(n6751), .B(n6750), .Z(n7360) );
  XOR U7273 ( .A(n7362), .B(n7363), .Z(n6690) );
  XNOR U7274 ( .A(n4884), .B(n4055), .Z(n7363) );
  XOR U7275 ( .A(n7364), .B(n6726), .Z(n4055) );
  IV U7276 ( .A(n7365), .Z(n6726) );
  ANDN U7277 ( .B(n7286), .A(n7366), .Z(n7364) );
  XNOR U7278 ( .A(n7367), .B(n6739), .Z(n4884) );
  ANDN U7279 ( .B(n7284), .A(n7368), .Z(n7367) );
  IV U7280 ( .A(n7369), .Z(n7284) );
  XOR U7281 ( .A(n2586), .B(n7370), .Z(n7362) );
  XOR U7282 ( .A(n3495), .B(n7371), .Z(n7370) );
  XNOR U7283 ( .A(n7372), .B(n6731), .Z(n3495) );
  ANDN U7284 ( .B(n7373), .A(n7282), .Z(n7372) );
  XOR U7285 ( .A(n7374), .B(n6722), .Z(n2586) );
  IV U7286 ( .A(n7375), .Z(n6722) );
  NOR U7287 ( .A(n7279), .B(n7376), .Z(n7374) );
  XNOR U7288 ( .A(n3947), .B(n7377), .Z(n1066) );
  IV U7289 ( .A(n2357), .Z(n3947) );
  XOR U7290 ( .A(n6176), .B(n7378), .Z(n2357) );
  XOR U7291 ( .A(n7379), .B(n7380), .Z(n6176) );
  XNOR U7292 ( .A(n3188), .B(n7381), .Z(n7380) );
  XOR U7293 ( .A(n7382), .B(n7383), .Z(n3188) );
  NOR U7294 ( .A(n7384), .B(n7385), .Z(n7382) );
  XNOR U7295 ( .A(n5484), .B(n7386), .Z(n7379) );
  XOR U7296 ( .A(n7387), .B(n2396), .Z(n7386) );
  XOR U7297 ( .A(n7388), .B(n7389), .Z(n2396) );
  ANDN U7298 ( .B(n7390), .A(n7391), .Z(n7388) );
  XNOR U7299 ( .A(n7392), .B(n7393), .Z(n5484) );
  ANDN U7300 ( .B(n7394), .A(n7395), .Z(n7392) );
  XOR U7301 ( .A(n7396), .B(n5873), .Z(out[1056]) );
  XNOR U7302 ( .A(n7397), .B(n2284), .Z(n5873) );
  XOR U7303 ( .A(n7398), .B(n6002), .Z(n2284) );
  XNOR U7304 ( .A(n7399), .B(n7400), .Z(n6002) );
  XOR U7305 ( .A(n5306), .B(n3757), .Z(n7400) );
  XOR U7306 ( .A(n7401), .B(n7402), .Z(n3757) );
  XNOR U7307 ( .A(n7405), .B(n7406), .Z(n5306) );
  NOR U7308 ( .A(n7407), .B(n7408), .Z(n7405) );
  XNOR U7309 ( .A(n6096), .B(n7409), .Z(n7399) );
  XOR U7310 ( .A(n2628), .B(n4496), .Z(n7409) );
  XOR U7311 ( .A(n7410), .B(n7411), .Z(n4496) );
  XOR U7312 ( .A(n7414), .B(n7415), .Z(n2628) );
  ANDN U7313 ( .B(n7416), .A(n7417), .Z(n7414) );
  XNOR U7314 ( .A(n7418), .B(n7419), .Z(n6096) );
  AND U7315 ( .A(n7420), .B(n7421), .Z(n7418) );
  ANDN U7316 ( .B(n1072), .A(n1070), .Z(n7396) );
  XOR U7317 ( .A(n7422), .B(n3407), .Z(n1070) );
  IV U7318 ( .A(n2364), .Z(n3407) );
  XOR U7319 ( .A(n7423), .B(n7424), .Z(n6181) );
  XOR U7320 ( .A(n3191), .B(n7425), .Z(n7424) );
  XNOR U7321 ( .A(n7426), .B(n7427), .Z(n3191) );
  ANDN U7322 ( .B(n7428), .A(n7429), .Z(n7426) );
  XOR U7323 ( .A(n5489), .B(n7430), .Z(n7423) );
  XOR U7324 ( .A(n7431), .B(n2401), .Z(n7430) );
  XNOR U7325 ( .A(n7432), .B(n7433), .Z(n2401) );
  ANDN U7326 ( .B(n7434), .A(n7435), .Z(n7432) );
  XNOR U7327 ( .A(n7436), .B(n7437), .Z(n5489) );
  ANDN U7328 ( .B(n7438), .A(n7439), .Z(n7436) );
  XNOR U7329 ( .A(n3567), .B(n7441), .Z(n1072) );
  IV U7330 ( .A(n1828), .Z(n3567) );
  XOR U7331 ( .A(n6716), .B(n6347), .Z(n1828) );
  XOR U7332 ( .A(n7442), .B(n7443), .Z(n6347) );
  XOR U7333 ( .A(n5920), .B(n5479), .Z(n7443) );
  XNOR U7334 ( .A(n7444), .B(n7445), .Z(n5479) );
  XOR U7335 ( .A(n7446), .B(n7447), .Z(n5920) );
  ANDN U7336 ( .B(n7448), .A(n6773), .Z(n7446) );
  XOR U7337 ( .A(n3721), .B(n7449), .Z(n7442) );
  XNOR U7338 ( .A(n4314), .B(n2154), .Z(n7449) );
  XNOR U7339 ( .A(n7450), .B(n7451), .Z(n2154) );
  NOR U7340 ( .A(n6786), .B(n6784), .Z(n7450) );
  XOR U7341 ( .A(n7452), .B(n7453), .Z(n4314) );
  NOR U7342 ( .A(n6792), .B(n6793), .Z(n7452) );
  XOR U7343 ( .A(n7454), .B(n7455), .Z(n3721) );
  AND U7344 ( .A(n6776), .B(n6781), .Z(n7454) );
  XOR U7345 ( .A(n7456), .B(n7457), .Z(n6716) );
  XNOR U7346 ( .A(n4887), .B(n4058), .Z(n7457) );
  XNOR U7347 ( .A(n7458), .B(n6752), .Z(n4058) );
  ANDN U7348 ( .B(n7459), .A(n7361), .Z(n7458) );
  XNOR U7349 ( .A(n7460), .B(n6765), .Z(n4887) );
  AND U7350 ( .A(n7461), .B(n7358), .Z(n7460) );
  IV U7351 ( .A(n7462), .Z(n7358) );
  XOR U7352 ( .A(n2591), .B(n7463), .Z(n7456) );
  XNOR U7353 ( .A(n3498), .B(n7464), .Z(n7463) );
  XOR U7354 ( .A(n7465), .B(n6757), .Z(n3498) );
  IV U7355 ( .A(n7466), .Z(n6757) );
  NOR U7356 ( .A(n7356), .B(n7467), .Z(n7465) );
  XOR U7357 ( .A(n7468), .B(n6747), .Z(n2591) );
  XOR U7358 ( .A(n7470), .B(n5878), .Z(out[1055]) );
  XNOR U7359 ( .A(n7471), .B(n2291), .Z(n5878) );
  XOR U7360 ( .A(n7472), .B(n6012), .Z(n2291) );
  XNOR U7361 ( .A(n7473), .B(n7474), .Z(n6012) );
  XOR U7362 ( .A(n5312), .B(n3762), .Z(n7474) );
  XOR U7363 ( .A(n7475), .B(n7476), .Z(n3762) );
  XNOR U7364 ( .A(n7479), .B(n7480), .Z(n5312) );
  NOR U7365 ( .A(n7481), .B(n7482), .Z(n7479) );
  XNOR U7366 ( .A(n6101), .B(n7483), .Z(n7473) );
  XNOR U7367 ( .A(n2635), .B(n4544), .Z(n7483) );
  XOR U7368 ( .A(n7484), .B(n7485), .Z(n4544) );
  NOR U7369 ( .A(n7486), .B(n7487), .Z(n7484) );
  XNOR U7370 ( .A(n7488), .B(n7489), .Z(n2635) );
  ANDN U7371 ( .B(n7490), .A(n7491), .Z(n7488) );
  XOR U7372 ( .A(n7492), .B(n7493), .Z(n6101) );
  ANDN U7373 ( .B(n7494), .A(n7495), .Z(n7492) );
  ANDN U7374 ( .B(n1074), .A(n1076), .Z(n7470) );
  XNOR U7375 ( .A(n1832), .B(n7496), .Z(n1076) );
  XNOR U7376 ( .A(n6742), .B(n6574), .Z(n1832) );
  XOR U7377 ( .A(n7497), .B(n7498), .Z(n6574) );
  XNOR U7378 ( .A(n5925), .B(n2158), .Z(n7498) );
  XOR U7379 ( .A(n7499), .B(n7500), .Z(n2158) );
  AND U7380 ( .A(n6811), .B(n6812), .Z(n7499) );
  XOR U7381 ( .A(n7501), .B(n7502), .Z(n5925) );
  AND U7382 ( .A(n6802), .B(n7503), .Z(n7501) );
  XNOR U7383 ( .A(n3727), .B(n7504), .Z(n7497) );
  XOR U7384 ( .A(n4319), .B(n5483), .Z(n7504) );
  XNOR U7385 ( .A(n7505), .B(n7506), .Z(n5483) );
  AND U7386 ( .A(n6815), .B(n6817), .Z(n7505) );
  XNOR U7387 ( .A(n7507), .B(n7508), .Z(n4319) );
  ANDN U7388 ( .B(n6821), .A(n6819), .Z(n7507) );
  XNOR U7389 ( .A(n7509), .B(n7510), .Z(n3727) );
  AND U7390 ( .A(n6808), .B(n6806), .Z(n7509) );
  IV U7391 ( .A(n7511), .Z(n6806) );
  XOR U7392 ( .A(n7512), .B(n7513), .Z(n6742) );
  XOR U7393 ( .A(n4890), .B(n4236), .Z(n7513) );
  XNOR U7394 ( .A(n7514), .B(n6780), .Z(n4236) );
  AND U7395 ( .A(n7515), .B(n7455), .Z(n7514) );
  IV U7396 ( .A(n7516), .Z(n7455) );
  XOR U7397 ( .A(n7517), .B(n6794), .Z(n4890) );
  AND U7398 ( .A(n7518), .B(n7453), .Z(n7517) );
  IV U7399 ( .A(n7519), .Z(n7453) );
  XOR U7400 ( .A(n2604), .B(n7520), .Z(n7512) );
  XOR U7401 ( .A(n3500), .B(n7521), .Z(n7520) );
  XOR U7402 ( .A(n7522), .B(n6785), .Z(n3500) );
  ANDN U7403 ( .B(n7523), .A(n7524), .Z(n7522) );
  XOR U7404 ( .A(n7525), .B(n6775), .Z(n2604) );
  IV U7405 ( .A(n7527), .Z(n7447) );
  XNOR U7406 ( .A(n2369), .B(n7528), .Z(n1074) );
  IV U7407 ( .A(n5007), .Z(n2369) );
  XOR U7408 ( .A(n6185), .B(n7529), .Z(n5007) );
  XOR U7409 ( .A(n7530), .B(n7531), .Z(n6185) );
  XNOR U7410 ( .A(n3194), .B(n7532), .Z(n7531) );
  XOR U7411 ( .A(n7533), .B(n7534), .Z(n3194) );
  AND U7412 ( .A(n7535), .B(n7536), .Z(n7533) );
  XOR U7413 ( .A(n5492), .B(n7537), .Z(n7530) );
  XOR U7414 ( .A(n7538), .B(n2410), .Z(n7537) );
  XNOR U7415 ( .A(n7539), .B(n7540), .Z(n2410) );
  ANDN U7416 ( .B(n7541), .A(n7542), .Z(n7539) );
  XNOR U7417 ( .A(n7543), .B(n7544), .Z(n5492) );
  AND U7418 ( .A(n7545), .B(n7546), .Z(n7543) );
  XOR U7419 ( .A(n7547), .B(n5883), .Z(out[1054]) );
  XOR U7420 ( .A(n7548), .B(n2298), .Z(n5883) );
  XOR U7421 ( .A(n7549), .B(n6017), .Z(n2298) );
  XNOR U7422 ( .A(n7550), .B(n7551), .Z(n6017) );
  XNOR U7423 ( .A(n5319), .B(n3766), .Z(n7551) );
  XOR U7424 ( .A(n7552), .B(n7553), .Z(n3766) );
  ANDN U7425 ( .B(n7554), .A(n7555), .Z(n7552) );
  XNOR U7426 ( .A(n7556), .B(n7557), .Z(n5319) );
  NOR U7427 ( .A(n7558), .B(n7559), .Z(n7556) );
  XOR U7428 ( .A(n6106), .B(n7560), .Z(n7550) );
  XOR U7429 ( .A(n2642), .B(n4590), .Z(n7560) );
  XOR U7430 ( .A(n7561), .B(n7562), .Z(n4590) );
  ANDN U7431 ( .B(n7563), .A(n7564), .Z(n7561) );
  XNOR U7432 ( .A(n7565), .B(n7566), .Z(n2642) );
  AND U7433 ( .A(n7567), .B(n7568), .Z(n7565) );
  XNOR U7434 ( .A(n7569), .B(n7570), .Z(n6106) );
  NOR U7435 ( .A(n7571), .B(n7572), .Z(n7569) );
  ANDN U7436 ( .B(n1078), .A(n1080), .Z(n7547) );
  XNOR U7437 ( .A(n1837), .B(n7573), .Z(n1080) );
  XNOR U7438 ( .A(n6769), .B(n6850), .Z(n1837) );
  XOR U7439 ( .A(n7574), .B(n7575), .Z(n6850) );
  XOR U7440 ( .A(n5930), .B(n2162), .Z(n7575) );
  XNOR U7441 ( .A(n7576), .B(n7577), .Z(n2162) );
  NOR U7442 ( .A(n6853), .B(n6854), .Z(n7576) );
  XNOR U7443 ( .A(n7578), .B(n7579), .Z(n5930) );
  AND U7444 ( .A(n6828), .B(n6830), .Z(n7578) );
  XOR U7445 ( .A(n3731), .B(n7580), .Z(n7574) );
  XOR U7446 ( .A(n4322), .B(n5487), .Z(n7580) );
  XOR U7447 ( .A(n7581), .B(n7582), .Z(n5487) );
  AND U7448 ( .A(n6844), .B(n6842), .Z(n7581) );
  XOR U7449 ( .A(n7583), .B(n7584), .Z(n4322) );
  XOR U7450 ( .A(n7585), .B(n7586), .Z(n3731) );
  XOR U7451 ( .A(n7587), .B(n7588), .Z(n6769) );
  XNOR U7452 ( .A(n4893), .B(n7589), .Z(n7588) );
  XNOR U7453 ( .A(n7590), .B(n6820), .Z(n4893) );
  ANDN U7454 ( .B(n7591), .A(n7592), .Z(n7590) );
  XOR U7455 ( .A(n2609), .B(n7593), .Z(n7587) );
  XNOR U7456 ( .A(n3503), .B(n7594), .Z(n7593) );
  XNOR U7457 ( .A(n7595), .B(n6813), .Z(n3503) );
  ANDN U7458 ( .B(n7500), .A(n7596), .Z(n7595) );
  IV U7459 ( .A(n7597), .Z(n7500) );
  XOR U7460 ( .A(n7598), .B(n6803), .Z(n2609) );
  AND U7461 ( .A(n7599), .B(n7502), .Z(n7598) );
  IV U7462 ( .A(n7600), .Z(n7502) );
  XNOR U7463 ( .A(n3412), .B(n7601), .Z(n1078) );
  IV U7464 ( .A(n2382), .Z(n3412) );
  XOR U7465 ( .A(n6189), .B(n7602), .Z(n2382) );
  XOR U7466 ( .A(n7603), .B(n7604), .Z(n6189) );
  XNOR U7467 ( .A(n7605), .B(n3197), .Z(n7604) );
  XOR U7468 ( .A(n7606), .B(n7607), .Z(n3197) );
  AND U7469 ( .A(n7608), .B(n7609), .Z(n7606) );
  XNOR U7470 ( .A(n2416), .B(n7610), .Z(n7603) );
  XOR U7471 ( .A(n4335), .B(n5496), .Z(n7610) );
  XNOR U7472 ( .A(n7611), .B(n7612), .Z(n5496) );
  NOR U7473 ( .A(n7613), .B(n7614), .Z(n7611) );
  XNOR U7474 ( .A(n7615), .B(n7616), .Z(n4335) );
  ANDN U7475 ( .B(n7617), .A(n7618), .Z(n7615) );
  XNOR U7476 ( .A(n7619), .B(n7620), .Z(n2416) );
  ANDN U7477 ( .B(n7621), .A(n7622), .Z(n7619) );
  XOR U7478 ( .A(n7623), .B(n5888), .Z(out[1053]) );
  IV U7479 ( .A(n6227), .Z(n5888) );
  XOR U7480 ( .A(n7624), .B(n2309), .Z(n6227) );
  XOR U7481 ( .A(n7625), .B(n6022), .Z(n2309) );
  XNOR U7482 ( .A(n7626), .B(n7627), .Z(n6022) );
  XNOR U7483 ( .A(n5323), .B(n3772), .Z(n7627) );
  XOR U7484 ( .A(n7628), .B(n7629), .Z(n3772) );
  NOR U7485 ( .A(n7630), .B(n7631), .Z(n7628) );
  XNOR U7486 ( .A(n7632), .B(n7633), .Z(n5323) );
  AND U7487 ( .A(n7634), .B(n7635), .Z(n7632) );
  XOR U7488 ( .A(n6116), .B(n7636), .Z(n7626) );
  XOR U7489 ( .A(n2649), .B(n4635), .Z(n7636) );
  XNOR U7490 ( .A(n7637), .B(n7638), .Z(n4635) );
  AND U7491 ( .A(n7639), .B(n7640), .Z(n7637) );
  XNOR U7492 ( .A(n7641), .B(n7642), .Z(n2649) );
  AND U7493 ( .A(n7643), .B(n7644), .Z(n7641) );
  XNOR U7494 ( .A(n7645), .B(n7646), .Z(n6116) );
  AND U7495 ( .A(n1088), .B(n1086), .Z(n7623) );
  XNOR U7496 ( .A(n7649), .B(n2388), .Z(n1086) );
  XOR U7497 ( .A(n6193), .B(n7650), .Z(n2388) );
  XOR U7498 ( .A(n7651), .B(n7652), .Z(n6193) );
  XOR U7499 ( .A(n7653), .B(n3200), .Z(n7652) );
  XOR U7500 ( .A(n7654), .B(n7655), .Z(n3200) );
  AND U7501 ( .A(n7656), .B(n7657), .Z(n7654) );
  XOR U7502 ( .A(n2425), .B(n7658), .Z(n7651) );
  XOR U7503 ( .A(n4339), .B(n5501), .Z(n7658) );
  XNOR U7504 ( .A(n7659), .B(n7660), .Z(n5501) );
  ANDN U7505 ( .B(n7661), .A(n7662), .Z(n7659) );
  XNOR U7506 ( .A(n7663), .B(n7664), .Z(n4339) );
  ANDN U7507 ( .B(n7665), .A(n7666), .Z(n7663) );
  XNOR U7508 ( .A(n7667), .B(n7668), .Z(n2425) );
  AND U7509 ( .A(n7669), .B(n7670), .Z(n7667) );
  XNOR U7510 ( .A(n3585), .B(n7671), .Z(n1088) );
  IV U7511 ( .A(n1841), .Z(n3585) );
  XOR U7512 ( .A(n6798), .B(n7183), .Z(n1841) );
  XOR U7513 ( .A(n7672), .B(n7673), .Z(n7183) );
  XNOR U7514 ( .A(n5935), .B(n2165), .Z(n7673) );
  XOR U7515 ( .A(n7674), .B(n7675), .Z(n2165) );
  NOR U7516 ( .A(n7186), .B(n7187), .Z(n7674) );
  XOR U7517 ( .A(n7676), .B(n7677), .Z(n5935) );
  ANDN U7518 ( .B(n6864), .A(n6866), .Z(n7676) );
  XOR U7519 ( .A(n5491), .B(n7678), .Z(n7672) );
  XOR U7520 ( .A(n4324), .B(n3736), .Z(n7678) );
  XOR U7521 ( .A(n7679), .B(n7680), .Z(n3736) );
  ANDN U7522 ( .B(n6872), .A(n6867), .Z(n7679) );
  XOR U7523 ( .A(n7681), .B(n7682), .Z(n4324) );
  NOR U7524 ( .A(n6881), .B(n6880), .Z(n7681) );
  IV U7525 ( .A(n7683), .Z(n6881) );
  XNOR U7526 ( .A(n7684), .B(n7685), .Z(n5491) );
  XOR U7527 ( .A(n7686), .B(n7687), .Z(n6798) );
  XOR U7528 ( .A(n4896), .B(n5557), .Z(n7687) );
  XNOR U7529 ( .A(n7688), .B(n6838), .Z(n5557) );
  AND U7530 ( .A(n7586), .B(n7689), .Z(n7688) );
  XOR U7531 ( .A(n7690), .B(n6847), .Z(n4896) );
  AND U7532 ( .A(n7691), .B(n7584), .Z(n7690) );
  IV U7533 ( .A(n7692), .Z(n7584) );
  XOR U7534 ( .A(n2616), .B(n7693), .Z(n7686) );
  XOR U7535 ( .A(n3506), .B(n7694), .Z(n7693) );
  XOR U7536 ( .A(n7695), .B(n6855), .Z(n3506) );
  IV U7537 ( .A(n7696), .Z(n6855) );
  ANDN U7538 ( .B(n7697), .A(n7577), .Z(n7695) );
  XOR U7539 ( .A(n7698), .B(n6829), .Z(n2616) );
  ANDN U7540 ( .B(n7699), .A(n7579), .Z(n7698) );
  XOR U7541 ( .A(n7700), .B(n5893), .Z(out[1052]) );
  XNOR U7542 ( .A(n7701), .B(n6114), .Z(n5893) );
  XOR U7543 ( .A(n7702), .B(n6027), .Z(n6114) );
  XNOR U7544 ( .A(n7703), .B(n7704), .Z(n6027) );
  XOR U7545 ( .A(n5327), .B(n3778), .Z(n7704) );
  XOR U7546 ( .A(n7705), .B(n7706), .Z(n3778) );
  XNOR U7547 ( .A(n7709), .B(n7710), .Z(n5327) );
  ANDN U7548 ( .B(n7711), .A(n7712), .Z(n7709) );
  XNOR U7549 ( .A(n6121), .B(n7713), .Z(n7703) );
  XNOR U7550 ( .A(n2656), .B(n4674), .Z(n7713) );
  XOR U7551 ( .A(n7714), .B(n7715), .Z(n4674) );
  XOR U7552 ( .A(n7718), .B(n7719), .Z(n2656) );
  XOR U7553 ( .A(n7722), .B(n7723), .Z(n6121) );
  ANDN U7554 ( .B(n7724), .A(n7725), .Z(n7722) );
  AND U7555 ( .A(n1092), .B(n1090), .Z(n7700) );
  XNOR U7556 ( .A(n7726), .B(n2395), .Z(n1090) );
  XOR U7557 ( .A(n6197), .B(n7727), .Z(n2395) );
  XOR U7558 ( .A(n7728), .B(n7729), .Z(n6197) );
  XNOR U7559 ( .A(n3207), .B(n4345), .Z(n7729) );
  XNOR U7560 ( .A(n7730), .B(n7731), .Z(n4345) );
  NOR U7561 ( .A(n7732), .B(n7733), .Z(n7730) );
  XNOR U7562 ( .A(n7734), .B(n7735), .Z(n3207) );
  NOR U7563 ( .A(n7736), .B(n7737), .Z(n7734) );
  XNOR U7564 ( .A(n5504), .B(n7738), .Z(n7728) );
  XOR U7565 ( .A(n7739), .B(n2429), .Z(n7738) );
  XOR U7566 ( .A(n7740), .B(n7741), .Z(n2429) );
  ANDN U7567 ( .B(n7742), .A(n7743), .Z(n7740) );
  XNOR U7568 ( .A(n7744), .B(n7745), .Z(n5504) );
  ANDN U7569 ( .B(n7746), .A(n7747), .Z(n7744) );
  XNOR U7570 ( .A(n1845), .B(n7748), .Z(n1092) );
  XNOR U7571 ( .A(n6824), .B(n7749), .Z(n1845) );
  XOR U7572 ( .A(n7750), .B(n7751), .Z(n6824) );
  XNOR U7573 ( .A(n4899), .B(n5600), .Z(n7751) );
  XOR U7574 ( .A(n7752), .B(n6871), .Z(n5600) );
  ANDN U7575 ( .B(n7680), .A(n7753), .Z(n7752) );
  IV U7576 ( .A(n7754), .Z(n7680) );
  XNOR U7577 ( .A(n7755), .B(n6882), .Z(n4899) );
  IV U7578 ( .A(n7757), .Z(n7682) );
  XOR U7579 ( .A(n2623), .B(n7758), .Z(n7750) );
  XOR U7580 ( .A(n3514), .B(n7759), .Z(n7758) );
  XOR U7581 ( .A(n7760), .B(n7188), .Z(n3514) );
  IV U7582 ( .A(n7761), .Z(n7188) );
  ANDN U7583 ( .B(n7675), .A(n7762), .Z(n7760) );
  IV U7584 ( .A(n7763), .Z(n7675) );
  XOR U7585 ( .A(n7764), .B(n6865), .Z(n2623) );
  ANDN U7586 ( .B(n7677), .A(n7765), .Z(n7764) );
  IV U7587 ( .A(n7766), .Z(n7677) );
  XOR U7588 ( .A(n7767), .B(n5903), .Z(out[1051]) );
  XOR U7589 ( .A(n7768), .B(n5434), .Z(n5903) );
  XOR U7590 ( .A(n7769), .B(n6032), .Z(n5434) );
  XNOR U7591 ( .A(n7770), .B(n7771), .Z(n6032) );
  XNOR U7592 ( .A(n5332), .B(n3784), .Z(n7771) );
  XOR U7593 ( .A(n7772), .B(n7773), .Z(n3784) );
  AND U7594 ( .A(n7774), .B(n7775), .Z(n7772) );
  XOR U7595 ( .A(n7776), .B(n7777), .Z(n5332) );
  ANDN U7596 ( .B(n7778), .A(n7779), .Z(n7776) );
  XOR U7597 ( .A(n6126), .B(n7780), .Z(n7770) );
  XOR U7598 ( .A(n2663), .B(n4699), .Z(n7780) );
  XNOR U7599 ( .A(n7781), .B(n7782), .Z(n4699) );
  XOR U7600 ( .A(n7785), .B(n7786), .Z(n2663) );
  AND U7601 ( .A(n7787), .B(n7788), .Z(n7785) );
  XNOR U7602 ( .A(n7789), .B(n7790), .Z(n6126) );
  ANDN U7603 ( .B(n7791), .A(n7792), .Z(n7789) );
  ANDN U7604 ( .B(n1094), .A(n1096), .Z(n7767) );
  XNOR U7605 ( .A(n1850), .B(n7793), .Z(n1096) );
  IV U7606 ( .A(n4098), .Z(n1850) );
  XOR U7607 ( .A(n6860), .B(n7794), .Z(n4098) );
  XOR U7608 ( .A(n7795), .B(n7796), .Z(n6860) );
  XOR U7609 ( .A(n4902), .B(n7797), .Z(n7796) );
  XNOR U7610 ( .A(n7798), .B(n6906), .Z(n4902) );
  NOR U7611 ( .A(n7799), .B(n7800), .Z(n7798) );
  XNOR U7612 ( .A(n2630), .B(n7801), .Z(n7795) );
  XNOR U7613 ( .A(n3516), .B(n5646), .Z(n7801) );
  XNOR U7614 ( .A(n7802), .B(n6895), .Z(n5646) );
  AND U7615 ( .A(n7803), .B(n7804), .Z(n7802) );
  XOR U7616 ( .A(n7805), .B(n7806), .Z(n3516) );
  ANDN U7617 ( .B(n7807), .A(n7808), .Z(n7805) );
  XNOR U7618 ( .A(n7809), .B(n6891), .Z(n2630) );
  ANDN U7619 ( .B(n7810), .A(n7811), .Z(n7809) );
  XOR U7620 ( .A(n2403), .B(n7812), .Z(n1094) );
  XNOR U7621 ( .A(n6201), .B(n7813), .Z(n2403) );
  XOR U7622 ( .A(n7814), .B(n7815), .Z(n6201) );
  XNOR U7623 ( .A(n3210), .B(n4349), .Z(n7815) );
  XOR U7624 ( .A(n7816), .B(n7817), .Z(n4349) );
  ANDN U7625 ( .B(n7818), .A(n7819), .Z(n7816) );
  XOR U7626 ( .A(n7820), .B(n7821), .Z(n3210) );
  NOR U7627 ( .A(n7822), .B(n7823), .Z(n7820) );
  XOR U7628 ( .A(n5509), .B(n7824), .Z(n7814) );
  XNOR U7629 ( .A(n7825), .B(n2438), .Z(n7824) );
  XOR U7630 ( .A(n7826), .B(n7827), .Z(n2438) );
  XOR U7631 ( .A(n7830), .B(n7831), .Z(n5509) );
  ANDN U7632 ( .B(n7832), .A(n7833), .Z(n7830) );
  XOR U7633 ( .A(n7834), .B(n5908), .Z(out[1050]) );
  XOR U7634 ( .A(n7835), .B(n2328), .Z(n5908) );
  XNOR U7635 ( .A(n7836), .B(n6038), .Z(n2328) );
  XNOR U7636 ( .A(n7837), .B(n7838), .Z(n6038) );
  XNOR U7637 ( .A(n5338), .B(n3789), .Z(n7838) );
  XNOR U7638 ( .A(n7839), .B(n7840), .Z(n3789) );
  AND U7639 ( .A(n7841), .B(n7842), .Z(n7839) );
  XNOR U7640 ( .A(n7843), .B(n7844), .Z(n5338) );
  AND U7641 ( .A(n7845), .B(n7846), .Z(n7843) );
  XNOR U7642 ( .A(n6131), .B(n7847), .Z(n7837) );
  XNOR U7643 ( .A(n2196), .B(n4726), .Z(n7847) );
  XNOR U7644 ( .A(n7848), .B(n7849), .Z(n4726) );
  ANDN U7645 ( .B(n7850), .A(n7851), .Z(n7848) );
  XOR U7646 ( .A(n7852), .B(n7853), .Z(n2196) );
  AND U7647 ( .A(n7854), .B(n7855), .Z(n7852) );
  XNOR U7648 ( .A(n7856), .B(n7857), .Z(n6131) );
  AND U7649 ( .A(n1099), .B(n1098), .Z(n7834) );
  XNOR U7650 ( .A(n2408), .B(n7860), .Z(n1098) );
  XNOR U7651 ( .A(n6205), .B(n7861), .Z(n2408) );
  XOR U7652 ( .A(n7862), .B(n7863), .Z(n6205) );
  XOR U7653 ( .A(n3214), .B(n4359), .Z(n7863) );
  XNOR U7654 ( .A(n7864), .B(n7865), .Z(n4359) );
  ANDN U7655 ( .B(n7866), .A(n7867), .Z(n7864) );
  XOR U7656 ( .A(n7868), .B(n7869), .Z(n3214) );
  XOR U7657 ( .A(n5516), .B(n7872), .Z(n7862) );
  XNOR U7658 ( .A(n7873), .B(n2445), .Z(n7872) );
  AND U7659 ( .A(n7876), .B(n7877), .Z(n7874) );
  XOR U7660 ( .A(n7878), .B(n7879), .Z(n5516) );
  ANDN U7661 ( .B(n7880), .A(n7881), .Z(n7878) );
  XNOR U7662 ( .A(n1854), .B(n7882), .Z(n1099) );
  IV U7663 ( .A(n4102), .Z(n1854) );
  XOR U7664 ( .A(n6885), .B(n7883), .Z(n4102) );
  XOR U7665 ( .A(n7884), .B(n7885), .Z(n6885) );
  XNOR U7666 ( .A(n4909), .B(n7886), .Z(n7885) );
  XNOR U7667 ( .A(n7887), .B(n7888), .Z(n4909) );
  NOR U7668 ( .A(n7889), .B(n7890), .Z(n7887) );
  XOR U7669 ( .A(n2637), .B(n7891), .Z(n7884) );
  XOR U7670 ( .A(n3519), .B(n5679), .Z(n7891) );
  XOR U7671 ( .A(n7892), .B(n7893), .Z(n5679) );
  NOR U7672 ( .A(n7894), .B(n7895), .Z(n7892) );
  XNOR U7673 ( .A(n7896), .B(n7897), .Z(n3519) );
  NOR U7674 ( .A(n7898), .B(n7899), .Z(n7896) );
  XOR U7675 ( .A(n7900), .B(n7901), .Z(n2637) );
  ANDN U7676 ( .B(n7902), .A(n7903), .Z(n7900) );
  XOR U7677 ( .A(n7904), .B(n4149), .Z(out[104]) );
  XNOR U7678 ( .A(n6898), .B(n2541), .Z(n4149) );
  XNOR U7679 ( .A(n7749), .B(n7905), .Z(n2541) );
  XOR U7680 ( .A(n7906), .B(n7907), .Z(n7749) );
  XNOR U7681 ( .A(n4326), .B(n2168), .Z(n7907) );
  XOR U7682 ( .A(n7908), .B(n7909), .Z(n2168) );
  NOR U7683 ( .A(n7910), .B(n7911), .Z(n7908) );
  XOR U7684 ( .A(n7912), .B(n7800), .Z(n4326) );
  NOR U7685 ( .A(n6904), .B(n6905), .Z(n7912) );
  XOR U7686 ( .A(n5940), .B(n7913), .Z(n7906) );
  XOR U7687 ( .A(n5495), .B(n3742), .Z(n7913) );
  XOR U7688 ( .A(n7914), .B(n7803), .Z(n3742) );
  AND U7689 ( .A(n6892), .B(n6896), .Z(n7914) );
  XNOR U7690 ( .A(n7915), .B(n7916), .Z(n5495) );
  AND U7691 ( .A(n6900), .B(n6902), .Z(n7915) );
  XOR U7692 ( .A(n7917), .B(n7810), .Z(n5940) );
  ANDN U7693 ( .B(n6889), .A(n6890), .Z(n7917) );
  XNOR U7694 ( .A(n7918), .B(n7911), .Z(n6898) );
  AND U7695 ( .A(n7910), .B(n7806), .Z(n7918) );
  IV U7696 ( .A(n7919), .Z(n7806) );
  AND U7697 ( .A(n3477), .B(n3479), .Z(n7904) );
  XOR U7698 ( .A(n2313), .B(n7920), .Z(n3479) );
  IV U7699 ( .A(n3382), .Z(n2313) );
  XOR U7700 ( .A(n6142), .B(n7921), .Z(n3382) );
  XOR U7701 ( .A(n7922), .B(n7923), .Z(n6142) );
  XOR U7702 ( .A(n3164), .B(n6350), .Z(n7923) );
  XNOR U7703 ( .A(n7924), .B(n7925), .Z(n6350) );
  AND U7704 ( .A(n7926), .B(n7927), .Z(n7924) );
  XNOR U7705 ( .A(n7928), .B(n7929), .Z(n3164) );
  ANDN U7706 ( .B(n7930), .A(n7931), .Z(n7928) );
  XOR U7707 ( .A(n5452), .B(n7932), .Z(n7922) );
  XOR U7708 ( .A(n7933), .B(n2348), .Z(n7932) );
  XNOR U7709 ( .A(n7934), .B(n7935), .Z(n2348) );
  ANDN U7710 ( .B(n7936), .A(n7937), .Z(n7934) );
  XOR U7711 ( .A(n7938), .B(n7939), .Z(n5452) );
  NOR U7712 ( .A(n7940), .B(n7941), .Z(n7938) );
  XNOR U7713 ( .A(n7942), .B(n2381), .Z(n3477) );
  XNOR U7714 ( .A(n7943), .B(n5913), .Z(out[1049]) );
  XOR U7715 ( .A(n7944), .B(n2335), .Z(n5913) );
  XNOR U7716 ( .A(n7945), .B(n6043), .Z(n2335) );
  XNOR U7717 ( .A(n7946), .B(n7947), .Z(n6043) );
  XNOR U7718 ( .A(n5342), .B(n3792), .Z(n7947) );
  XOR U7719 ( .A(n7948), .B(n7949), .Z(n3792) );
  NOR U7720 ( .A(n7950), .B(n7951), .Z(n7948) );
  XNOR U7721 ( .A(n7952), .B(n7953), .Z(n5342) );
  AND U7722 ( .A(n7954), .B(n7955), .Z(n7952) );
  XNOR U7723 ( .A(n6136), .B(n7956), .Z(n7946) );
  XOR U7724 ( .A(n2203), .B(n4757), .Z(n7956) );
  XNOR U7725 ( .A(n7957), .B(n7958), .Z(n4757) );
  XNOR U7726 ( .A(n7961), .B(n7962), .Z(n2203) );
  XNOR U7727 ( .A(n7965), .B(n7966), .Z(n6136) );
  ANDN U7728 ( .B(n7967), .A(n7968), .Z(n7965) );
  AND U7729 ( .A(n1104), .B(n1102), .Z(n7943) );
  XNOR U7730 ( .A(n4016), .B(n7969), .Z(n1102) );
  IV U7731 ( .A(n2417), .Z(n4016) );
  XOR U7732 ( .A(n6209), .B(n7970), .Z(n2417) );
  XOR U7733 ( .A(n7971), .B(n7972), .Z(n6209) );
  XOR U7734 ( .A(n3218), .B(n4406), .Z(n7972) );
  XNOR U7735 ( .A(n7973), .B(n7974), .Z(n4406) );
  NOR U7736 ( .A(n7975), .B(n7976), .Z(n7973) );
  XNOR U7737 ( .A(n7977), .B(n7978), .Z(n3218) );
  NOR U7738 ( .A(n7979), .B(n7980), .Z(n7977) );
  XNOR U7739 ( .A(n5519), .B(n7981), .Z(n7971) );
  XNOR U7740 ( .A(n7982), .B(n2454), .Z(n7981) );
  XNOR U7741 ( .A(n7983), .B(n7984), .Z(n2454) );
  ANDN U7742 ( .B(n7985), .A(n7986), .Z(n7983) );
  XOR U7743 ( .A(n7987), .B(n7988), .Z(n5519) );
  NOR U7744 ( .A(n7989), .B(n7990), .Z(n7987) );
  XNOR U7745 ( .A(n1858), .B(n7991), .Z(n1104) );
  IV U7746 ( .A(n5187), .Z(n1858) );
  XOR U7747 ( .A(n7992), .B(n7993), .Z(n5187) );
  XOR U7748 ( .A(n7994), .B(n5918), .Z(out[1048]) );
  XOR U7749 ( .A(n7995), .B(n2344), .Z(n5918) );
  IV U7750 ( .A(n3161), .Z(n2344) );
  XNOR U7751 ( .A(n7996), .B(n6048), .Z(n3161) );
  XNOR U7752 ( .A(n7997), .B(n7998), .Z(n6048) );
  XOR U7753 ( .A(n5348), .B(n3797), .Z(n7998) );
  XOR U7754 ( .A(n7999), .B(n8000), .Z(n3797) );
  XNOR U7755 ( .A(n8003), .B(n8004), .Z(n5348) );
  NOR U7756 ( .A(n8005), .B(n8006), .Z(n8003) );
  XNOR U7757 ( .A(n6141), .B(n8007), .Z(n7997) );
  XOR U7758 ( .A(n2210), .B(n4783), .Z(n8007) );
  XNOR U7759 ( .A(n8008), .B(n8009), .Z(n4783) );
  AND U7760 ( .A(n8010), .B(n8011), .Z(n8008) );
  XNOR U7761 ( .A(n8012), .B(n8013), .Z(n2210) );
  ANDN U7762 ( .B(n8014), .A(n8015), .Z(n8012) );
  XNOR U7763 ( .A(n8016), .B(n8017), .Z(n6141) );
  NOR U7764 ( .A(n8018), .B(n8019), .Z(n8016) );
  ANDN U7765 ( .B(n1106), .A(n1107), .Z(n7994) );
  XNOR U7766 ( .A(n1866), .B(n8020), .Z(n1107) );
  IV U7767 ( .A(n5190), .Z(n1866) );
  XOR U7768 ( .A(n6913), .B(n8021), .Z(n5190) );
  XOR U7769 ( .A(n8022), .B(n8023), .Z(n6913) );
  XNOR U7770 ( .A(n4915), .B(n8024), .Z(n8023) );
  XNOR U7771 ( .A(n8025), .B(n6957), .Z(n4915) );
  XOR U7772 ( .A(n2651), .B(n8028), .Z(n8022) );
  XOR U7773 ( .A(n3524), .B(n5730), .Z(n8028) );
  XOR U7774 ( .A(n8029), .B(n8030), .Z(n5730) );
  XNOR U7775 ( .A(n8033), .B(n8034), .Z(n3524) );
  ANDN U7776 ( .B(n8035), .A(n8036), .Z(n8033) );
  XOR U7777 ( .A(n8037), .B(n6942), .Z(n2651) );
  XNOR U7778 ( .A(n4053), .B(n8040), .Z(n1106) );
  XOR U7779 ( .A(n6217), .B(n8041), .Z(n4053) );
  XOR U7780 ( .A(n8042), .B(n8043), .Z(n6217) );
  XOR U7781 ( .A(n3221), .B(n4451), .Z(n8043) );
  XOR U7782 ( .A(n8044), .B(n8045), .Z(n4451) );
  ANDN U7783 ( .B(n8046), .A(n8047), .Z(n8044) );
  XNOR U7784 ( .A(n8048), .B(n8049), .Z(n3221) );
  NOR U7785 ( .A(n8050), .B(n8051), .Z(n8048) );
  XOR U7786 ( .A(n5524), .B(n8052), .Z(n8042) );
  XOR U7787 ( .A(n8053), .B(n2463), .Z(n8052) );
  XOR U7788 ( .A(n8054), .B(n8055), .Z(n2463) );
  NOR U7789 ( .A(n8056), .B(n8057), .Z(n8054) );
  XOR U7790 ( .A(n8058), .B(n8059), .Z(n5524) );
  ANDN U7791 ( .B(n8060), .A(n8061), .Z(n8058) );
  XOR U7792 ( .A(n8062), .B(n5923), .Z(out[1047]) );
  XOR U7793 ( .A(n7933), .B(n2349), .Z(n5923) );
  XNOR U7794 ( .A(n8063), .B(n8064), .Z(n2349) );
  XOR U7795 ( .A(n8065), .B(n8066), .Z(n7933) );
  NOR U7796 ( .A(n8067), .B(n8068), .Z(n8065) );
  ANDN U7797 ( .B(n1110), .A(n1112), .Z(n8062) );
  XNOR U7798 ( .A(n1870), .B(n8069), .Z(n1112) );
  IV U7799 ( .A(n5193), .Z(n1870) );
  XOR U7800 ( .A(n6063), .B(n6937), .Z(n5193) );
  XOR U7801 ( .A(n8070), .B(n8071), .Z(n6937) );
  XOR U7802 ( .A(n4918), .B(n8072), .Z(n8071) );
  XNOR U7803 ( .A(n8073), .B(n6980), .Z(n4918) );
  AND U7804 ( .A(n8074), .B(n8075), .Z(n8073) );
  XOR U7805 ( .A(n2658), .B(n8076), .Z(n8070) );
  XOR U7806 ( .A(n3526), .B(n5756), .Z(n8076) );
  XOR U7807 ( .A(n8077), .B(n6969), .Z(n5756) );
  NOR U7808 ( .A(n8078), .B(n8079), .Z(n8077) );
  XOR U7809 ( .A(n8080), .B(n8081), .Z(n3526) );
  NOR U7810 ( .A(n8082), .B(n8083), .Z(n8080) );
  XOR U7811 ( .A(n8084), .B(n6965), .Z(n2658) );
  AND U7812 ( .A(n8085), .B(n8086), .Z(n8084) );
  XOR U7813 ( .A(n8087), .B(n8088), .Z(n6063) );
  XOR U7814 ( .A(n4342), .B(n2187), .Z(n8088) );
  XNOR U7815 ( .A(n8089), .B(n8090), .Z(n2187) );
  ANDN U7816 ( .B(n7000), .A(n7001), .Z(n8089) );
  XNOR U7817 ( .A(n8091), .B(n8092), .Z(n4342) );
  AND U7818 ( .A(n7004), .B(n7006), .Z(n8091) );
  XOR U7819 ( .A(n5970), .B(n8093), .Z(n8087) );
  XNOR U7820 ( .A(n5518), .B(n3767), .Z(n8093) );
  XNOR U7821 ( .A(n8094), .B(n8095), .Z(n3767) );
  AND U7822 ( .A(n6993), .B(n6991), .Z(n8094) );
  XNOR U7823 ( .A(n8096), .B(n8097), .Z(n5518) );
  AND U7824 ( .A(n6996), .B(n6998), .Z(n8096) );
  XOR U7825 ( .A(n8098), .B(n8099), .Z(n5970) );
  NOR U7826 ( .A(n6989), .B(n6987), .Z(n8098) );
  IV U7827 ( .A(n8100), .Z(n6989) );
  XNOR U7828 ( .A(n4087), .B(n8101), .Z(n1110) );
  XOR U7829 ( .A(n6221), .B(n8102), .Z(n4087) );
  XOR U7830 ( .A(n8103), .B(n8104), .Z(n6221) );
  XNOR U7831 ( .A(n3225), .B(n4495), .Z(n8104) );
  XOR U7832 ( .A(n8105), .B(n8106), .Z(n4495) );
  AND U7833 ( .A(n8107), .B(n8108), .Z(n8105) );
  XOR U7834 ( .A(n8109), .B(n8110), .Z(n3225) );
  ANDN U7835 ( .B(n8111), .A(n8112), .Z(n8109) );
  XOR U7836 ( .A(n5528), .B(n8113), .Z(n8103) );
  XOR U7837 ( .A(n8114), .B(n2470), .Z(n8113) );
  XNOR U7838 ( .A(n8115), .B(n8116), .Z(n2470) );
  AND U7839 ( .A(n8117), .B(n8118), .Z(n8115) );
  XOR U7840 ( .A(n8119), .B(n8120), .Z(n5528) );
  ANDN U7841 ( .B(n8121), .A(n8122), .Z(n8119) );
  XOR U7842 ( .A(n8123), .B(n5928), .Z(out[1046]) );
  IV U7843 ( .A(n6256), .Z(n5928) );
  XOR U7844 ( .A(n8124), .B(n2356), .Z(n6256) );
  XNOR U7845 ( .A(n8125), .B(n8126), .Z(n2356) );
  AND U7846 ( .A(n1116), .B(n1114), .Z(n8123) );
  XNOR U7847 ( .A(n2436), .B(n8127), .Z(n1114) );
  IV U7848 ( .A(n5040), .Z(n2436) );
  XOR U7849 ( .A(n6225), .B(n8128), .Z(n5040) );
  XOR U7850 ( .A(n8129), .B(n8130), .Z(n6225) );
  XOR U7851 ( .A(n3228), .B(n4543), .Z(n8130) );
  XNOR U7852 ( .A(n8131), .B(n8132), .Z(n4543) );
  ANDN U7853 ( .B(n8133), .A(n8134), .Z(n8131) );
  XNOR U7854 ( .A(n8135), .B(n8136), .Z(n3228) );
  AND U7855 ( .A(n8137), .B(n8138), .Z(n8135) );
  XNOR U7856 ( .A(n5531), .B(n8139), .Z(n8129) );
  XNOR U7857 ( .A(n8140), .B(n2475), .Z(n8139) );
  XOR U7858 ( .A(n8141), .B(n8142), .Z(n2475) );
  NOR U7859 ( .A(n8143), .B(n8144), .Z(n8141) );
  XNOR U7860 ( .A(n8145), .B(n8146), .Z(n5531) );
  NOR U7861 ( .A(n8147), .B(n8148), .Z(n8145) );
  XNOR U7862 ( .A(n1874), .B(n8149), .Z(n1116) );
  IV U7863 ( .A(n4115), .Z(n1874) );
  XOR U7864 ( .A(n6068), .B(n6960), .Z(n4115) );
  XOR U7865 ( .A(n8150), .B(n8151), .Z(n6960) );
  XNOR U7866 ( .A(n4921), .B(n8152), .Z(n8151) );
  XOR U7867 ( .A(n8153), .B(n7005), .Z(n4921) );
  IV U7868 ( .A(n8154), .Z(n7005) );
  NOR U7869 ( .A(n8155), .B(n8092), .Z(n8153) );
  XOR U7870 ( .A(n2665), .B(n8156), .Z(n8150) );
  XNOR U7871 ( .A(n3528), .B(n5780), .Z(n8156) );
  XOR U7872 ( .A(n8157), .B(n6992), .Z(n5780) );
  NOR U7873 ( .A(n8158), .B(n8095), .Z(n8157) );
  XNOR U7874 ( .A(n8159), .B(n7002), .Z(n3528) );
  ANDN U7875 ( .B(n8160), .A(n8090), .Z(n8159) );
  XOR U7876 ( .A(n8161), .B(n6988), .Z(n2665) );
  XOR U7877 ( .A(n8163), .B(n8164), .Z(n6068) );
  XNOR U7878 ( .A(n4348), .B(n2190), .Z(n8164) );
  XOR U7879 ( .A(n8165), .B(n8166), .Z(n2190) );
  ANDN U7880 ( .B(n7058), .A(n7059), .Z(n8165) );
  XNOR U7881 ( .A(n8167), .B(n8168), .Z(n4348) );
  ANDN U7882 ( .B(n7062), .A(n7063), .Z(n8167) );
  IV U7883 ( .A(n8169), .Z(n7062) );
  XOR U7884 ( .A(n5975), .B(n8170), .Z(n8163) );
  XOR U7885 ( .A(n5522), .B(n3770), .Z(n8170) );
  XNOR U7886 ( .A(n8171), .B(n8172), .Z(n3770) );
  ANDN U7887 ( .B(n7049), .A(n7050), .Z(n8171) );
  XOR U7888 ( .A(n8173), .B(n8174), .Z(n5522) );
  ANDN U7889 ( .B(n7054), .A(n7055), .Z(n8173) );
  XOR U7890 ( .A(n8175), .B(n8176), .Z(n5975) );
  ANDN U7891 ( .B(n7045), .A(n7046), .Z(n8175) );
  XOR U7892 ( .A(n8177), .B(n5933), .Z(out[1045]) );
  XNOR U7893 ( .A(n8178), .B(n2363), .Z(n5933) );
  XNOR U7894 ( .A(n8179), .B(n8180), .Z(n2363) );
  AND U7895 ( .A(n1119), .B(n1118), .Z(n8177) );
  XOR U7896 ( .A(n2443), .B(n8181), .Z(n1118) );
  XNOR U7897 ( .A(n6230), .B(n8182), .Z(n2443) );
  XOR U7898 ( .A(n8183), .B(n8184), .Z(n6230) );
  XNOR U7899 ( .A(n3231), .B(n4589), .Z(n8184) );
  XOR U7900 ( .A(n8185), .B(n8186), .Z(n4589) );
  NOR U7901 ( .A(n8187), .B(n8188), .Z(n8185) );
  XNOR U7902 ( .A(n8189), .B(n8190), .Z(n3231) );
  ANDN U7903 ( .B(n8191), .A(n8192), .Z(n8189) );
  XOR U7904 ( .A(n5536), .B(n8193), .Z(n8183) );
  XNOR U7905 ( .A(n8194), .B(n2482), .Z(n8193) );
  XOR U7906 ( .A(n8195), .B(n8196), .Z(n2482) );
  XOR U7907 ( .A(n8199), .B(n8200), .Z(n5536) );
  NOR U7908 ( .A(n8201), .B(n8202), .Z(n8199) );
  XNOR U7909 ( .A(n1878), .B(n8203), .Z(n1119) );
  IV U7910 ( .A(n5202), .Z(n1878) );
  XOR U7911 ( .A(n6983), .B(n6072), .Z(n5202) );
  XOR U7912 ( .A(n8204), .B(n8205), .Z(n6072) );
  XNOR U7913 ( .A(n4356), .B(n2193), .Z(n8205) );
  XOR U7914 ( .A(n8206), .B(n8207), .Z(n2193) );
  NOR U7915 ( .A(n7114), .B(n7113), .Z(n8206) );
  XOR U7916 ( .A(n8208), .B(n8209), .Z(n4356) );
  ANDN U7917 ( .B(n7117), .A(n7119), .Z(n8208) );
  XNOR U7918 ( .A(n5980), .B(n8210), .Z(n8204) );
  XOR U7919 ( .A(n5526), .B(n3779), .Z(n8210) );
  XOR U7920 ( .A(n8211), .B(n8212), .Z(n3779) );
  ANDN U7921 ( .B(n7104), .A(n7106), .Z(n8211) );
  XOR U7922 ( .A(n8213), .B(n8214), .Z(n5526) );
  XNOR U7923 ( .A(n8216), .B(n8217), .Z(n5980) );
  ANDN U7924 ( .B(n7100), .A(n7101), .Z(n8216) );
  XOR U7925 ( .A(n8218), .B(n8219), .Z(n6983) );
  XNOR U7926 ( .A(n4924), .B(n8220), .Z(n8219) );
  XOR U7927 ( .A(n8221), .B(n7064), .Z(n4924) );
  ANDN U7928 ( .B(n8222), .A(n8168), .Z(n8221) );
  XNOR U7929 ( .A(n2198), .B(n8223), .Z(n8218) );
  XOR U7930 ( .A(n3530), .B(n5809), .Z(n8223) );
  XNOR U7931 ( .A(n8224), .B(n7051), .Z(n5809) );
  ANDN U7932 ( .B(n8225), .A(n8172), .Z(n8224) );
  XNOR U7933 ( .A(n8226), .B(n7060), .Z(n3530) );
  AND U7934 ( .A(n8227), .B(n8166), .Z(n8226) );
  IV U7935 ( .A(n8228), .Z(n8166) );
  XOR U7936 ( .A(n8229), .B(n7047), .Z(n2198) );
  XOR U7937 ( .A(n8231), .B(n5938), .Z(out[1044]) );
  IV U7938 ( .A(n6269), .Z(n5938) );
  XOR U7939 ( .A(n8232), .B(n2372), .Z(n6269) );
  XNOR U7940 ( .A(n8233), .B(n8234), .Z(n2372) );
  ANDN U7941 ( .B(n1122), .A(n1124), .Z(n8231) );
  XNOR U7942 ( .A(n3628), .B(n8235), .Z(n1124) );
  IV U7943 ( .A(n1883), .Z(n3628) );
  XOR U7944 ( .A(n7041), .B(n6077), .Z(n1883) );
  XOR U7945 ( .A(n8236), .B(n8237), .Z(n6077) );
  XNOR U7946 ( .A(n4405), .B(n1968), .Z(n8237) );
  XNOR U7947 ( .A(n8238), .B(n8239), .Z(n1968) );
  ANDN U7948 ( .B(n8240), .A(n7137), .Z(n8238) );
  XOR U7949 ( .A(n8241), .B(n8242), .Z(n4405) );
  AND U7950 ( .A(n7147), .B(n7145), .Z(n8241) );
  XOR U7951 ( .A(n5985), .B(n8243), .Z(n8236) );
  XOR U7952 ( .A(n5530), .B(n3782), .Z(n8243) );
  XOR U7953 ( .A(n8244), .B(n8245), .Z(n3782) );
  ANDN U7954 ( .B(n7132), .A(n7133), .Z(n8244) );
  XOR U7955 ( .A(n8246), .B(n8247), .Z(n5530) );
  NOR U7956 ( .A(n7141), .B(n7142), .Z(n8246) );
  XNOR U7957 ( .A(n8248), .B(n8249), .Z(n5985) );
  AND U7958 ( .A(n7128), .B(n8250), .Z(n8248) );
  XOR U7959 ( .A(n8251), .B(n8252), .Z(n7041) );
  XNOR U7960 ( .A(n4928), .B(n8253), .Z(n8252) );
  XNOR U7961 ( .A(n8254), .B(n7118), .Z(n4928) );
  ANDN U7962 ( .B(n8209), .A(n8255), .Z(n8254) );
  XOR U7963 ( .A(n2205), .B(n8256), .Z(n8251) );
  XOR U7964 ( .A(n3532), .B(n5842), .Z(n8256) );
  XNOR U7965 ( .A(n8257), .B(n7105), .Z(n5842) );
  AND U7966 ( .A(n8212), .B(n8258), .Z(n8257) );
  XOR U7967 ( .A(n8259), .B(n7115), .Z(n3532) );
  AND U7968 ( .A(n8260), .B(n8207), .Z(n8259) );
  IV U7969 ( .A(n8261), .Z(n8207) );
  XOR U7970 ( .A(n8262), .B(n8263), .Z(n2205) );
  ANDN U7971 ( .B(n8264), .A(n8217), .Z(n8262) );
  XNOR U7972 ( .A(n4191), .B(n8265), .Z(n1122) );
  IV U7973 ( .A(n2456), .Z(n4191) );
  XOR U7974 ( .A(n6234), .B(n8266), .Z(n2456) );
  XOR U7975 ( .A(n8267), .B(n8268), .Z(n6234) );
  XNOR U7976 ( .A(n3234), .B(n4634), .Z(n8268) );
  XOR U7977 ( .A(n8269), .B(n8270), .Z(n4634) );
  NOR U7978 ( .A(n8271), .B(n8272), .Z(n8269) );
  XOR U7979 ( .A(n8273), .B(n8274), .Z(n3234) );
  ANDN U7980 ( .B(n8275), .A(n8276), .Z(n8273) );
  XOR U7981 ( .A(n5540), .B(n8277), .Z(n8267) );
  XOR U7982 ( .A(n8278), .B(n2489), .Z(n8277) );
  XOR U7983 ( .A(n8279), .B(n8280), .Z(n2489) );
  ANDN U7984 ( .B(n8281), .A(n8282), .Z(n8279) );
  XOR U7985 ( .A(n8283), .B(n8284), .Z(n5540) );
  ANDN U7986 ( .B(n8285), .A(n8286), .Z(n8283) );
  XOR U7987 ( .A(n8287), .B(n5943), .Z(out[1043]) );
  IV U7988 ( .A(n6274), .Z(n5943) );
  XOR U7989 ( .A(n8288), .B(n2381), .Z(n6274) );
  XNOR U7990 ( .A(n8289), .B(n8290), .Z(n2381) );
  ANDN U7991 ( .B(n1130), .A(n1131), .Z(n8287) );
  XNOR U7992 ( .A(n3634), .B(n8291), .Z(n1131) );
  IV U7993 ( .A(n1888), .Z(n3634) );
  XOR U7994 ( .A(n7096), .B(n6082), .Z(n1888) );
  XOR U7995 ( .A(n8292), .B(n8293), .Z(n6082) );
  XNOR U7996 ( .A(n4449), .B(n1971), .Z(n8293) );
  XOR U7997 ( .A(n8294), .B(n8295), .Z(n1971) );
  XNOR U7998 ( .A(n8296), .B(n8297), .Z(n4449) );
  XOR U7999 ( .A(n5990), .B(n8298), .Z(n8292) );
  XNOR U8000 ( .A(n5534), .B(n3787), .Z(n8298) );
  XNOR U8001 ( .A(n8299), .B(n8300), .Z(n3787) );
  ANDN U8002 ( .B(n7201), .A(n7202), .Z(n8299) );
  XNOR U8003 ( .A(n8301), .B(n8302), .Z(n5534) );
  ANDN U8004 ( .B(n7212), .A(n7210), .Z(n8301) );
  XOR U8005 ( .A(n8303), .B(n8304), .Z(n5990) );
  AND U8006 ( .A(n7197), .B(n7199), .Z(n8303) );
  XOR U8007 ( .A(n8305), .B(n8306), .Z(n7096) );
  XOR U8008 ( .A(n4932), .B(n8307), .Z(n8306) );
  XNOR U8009 ( .A(n8308), .B(n7146), .Z(n4932) );
  ANDN U8010 ( .B(n8309), .A(n8242), .Z(n8308) );
  XOR U8011 ( .A(n2212), .B(n8310), .Z(n8305) );
  XOR U8012 ( .A(n3535), .B(n5896), .Z(n8310) );
  XNOR U8013 ( .A(n8311), .B(n7134), .Z(n5896) );
  ANDN U8014 ( .B(n8245), .A(n8312), .Z(n8311) );
  XNOR U8015 ( .A(n8313), .B(n7138), .Z(n3535) );
  ANDN U8016 ( .B(n8314), .A(n8239), .Z(n8313) );
  XNOR U8017 ( .A(n8315), .B(n7129), .Z(n2212) );
  NOR U8018 ( .A(n8249), .B(n8316), .Z(n8315) );
  XNOR U8019 ( .A(n2461), .B(n8317), .Z(n1130) );
  IV U8020 ( .A(n5053), .Z(n2461) );
  XOR U8021 ( .A(n6238), .B(n8318), .Z(n5053) );
  XOR U8022 ( .A(n8319), .B(n8320), .Z(n6238) );
  XOR U8023 ( .A(n3237), .B(n4675), .Z(n8320) );
  XNOR U8024 ( .A(n8321), .B(n8322), .Z(n4675) );
  ANDN U8025 ( .B(n8323), .A(n8324), .Z(n8321) );
  XOR U8026 ( .A(n8325), .B(n8326), .Z(n3237) );
  ANDN U8027 ( .B(n8327), .A(n8328), .Z(n8325) );
  XOR U8028 ( .A(n5544), .B(n8329), .Z(n8319) );
  XOR U8029 ( .A(n8330), .B(n2498), .Z(n8329) );
  XNOR U8030 ( .A(n8331), .B(n8332), .Z(n2498) );
  AND U8031 ( .A(n8333), .B(n8334), .Z(n8331) );
  XOR U8032 ( .A(n8335), .B(n8336), .Z(n5544) );
  XOR U8033 ( .A(n8339), .B(n5948), .Z(out[1042]) );
  IV U8034 ( .A(n6279), .Z(n5948) );
  XOR U8035 ( .A(n7310), .B(n2390), .Z(n6279) );
  XOR U8036 ( .A(n8340), .B(n8341), .Z(n7310) );
  NOR U8037 ( .A(n8342), .B(n8343), .Z(n8340) );
  AND U8038 ( .A(n1135), .B(n1134), .Z(n8339) );
  XNOR U8039 ( .A(n2468), .B(n8344), .Z(n1134) );
  XNOR U8040 ( .A(n6242), .B(n8345), .Z(n2468) );
  XOR U8041 ( .A(n8346), .B(n8347), .Z(n6242) );
  XNOR U8042 ( .A(n3244), .B(n4700), .Z(n8347) );
  XOR U8043 ( .A(n8348), .B(n8349), .Z(n4700) );
  NOR U8044 ( .A(n8350), .B(n8351), .Z(n8348) );
  XOR U8045 ( .A(n8352), .B(n8353), .Z(n3244) );
  ANDN U8046 ( .B(n8354), .A(n8355), .Z(n8352) );
  XOR U8047 ( .A(n5548), .B(n8356), .Z(n8346) );
  XNOR U8048 ( .A(n8357), .B(n2505), .Z(n8356) );
  XNOR U8049 ( .A(n8358), .B(n8359), .Z(n2505) );
  ANDN U8050 ( .B(n8360), .A(n8361), .Z(n8358) );
  XOR U8051 ( .A(n8362), .B(n8363), .Z(n5548) );
  NOR U8052 ( .A(n8364), .B(n8365), .Z(n8362) );
  XNOR U8053 ( .A(n1892), .B(n8366), .Z(n1135) );
  IV U8054 ( .A(n3639), .Z(n1892) );
  XOR U8055 ( .A(n7124), .B(n6087), .Z(n3639) );
  XOR U8056 ( .A(n8367), .B(n8368), .Z(n6087) );
  XOR U8057 ( .A(n4493), .B(n1974), .Z(n8368) );
  XOR U8058 ( .A(n8369), .B(n8370), .Z(n1974) );
  XNOR U8059 ( .A(n8371), .B(n8372), .Z(n4493) );
  NOR U8060 ( .A(n7270), .B(n7269), .Z(n8371) );
  XOR U8061 ( .A(n5995), .B(n8373), .Z(n8367) );
  XOR U8062 ( .A(n5538), .B(n3794), .Z(n8373) );
  XOR U8063 ( .A(n8374), .B(n8375), .Z(n3794) );
  AND U8064 ( .A(n7256), .B(n7258), .Z(n8374) );
  XOR U8065 ( .A(n8376), .B(n8377), .Z(n5538) );
  NOR U8066 ( .A(n7267), .B(n7265), .Z(n8376) );
  XOR U8067 ( .A(n8378), .B(n8379), .Z(n5995) );
  ANDN U8068 ( .B(n7254), .A(n7252), .Z(n8378) );
  XOR U8069 ( .A(n8380), .B(n8381), .Z(n7124) );
  XNOR U8070 ( .A(n4935), .B(n8382), .Z(n8381) );
  XOR U8071 ( .A(n8383), .B(n7215), .Z(n4935) );
  IV U8072 ( .A(n8384), .Z(n7215) );
  ANDN U8073 ( .B(n8385), .A(n8297), .Z(n8383) );
  XOR U8074 ( .A(n2219), .B(n8386), .Z(n8380) );
  XNOR U8075 ( .A(n3541), .B(n5951), .Z(n8386) );
  XOR U8076 ( .A(n8387), .B(n7203), .Z(n5951) );
  IV U8077 ( .A(n8388), .Z(n7203) );
  NOR U8078 ( .A(n8389), .B(n8300), .Z(n8387) );
  XNOR U8079 ( .A(n8390), .B(n7208), .Z(n3541) );
  AND U8080 ( .A(n8391), .B(n8295), .Z(n8390) );
  XOR U8081 ( .A(n8392), .B(n7198), .Z(n2219) );
  ANDN U8082 ( .B(n8304), .A(n8393), .Z(n8392) );
  XOR U8083 ( .A(n8394), .B(n5958), .Z(out[1041]) );
  XNOR U8084 ( .A(n7387), .B(n2397), .Z(n5958) );
  XOR U8085 ( .A(n8395), .B(n8396), .Z(n7387) );
  NOR U8086 ( .A(n8397), .B(n8398), .Z(n8395) );
  AND U8087 ( .A(n1140), .B(n1138), .Z(n8394) );
  XNOR U8088 ( .A(n2477), .B(n8399), .Z(n1138) );
  XOR U8089 ( .A(n5832), .B(n6246), .Z(n2477) );
  XOR U8090 ( .A(n8400), .B(n8401), .Z(n6246) );
  XNOR U8091 ( .A(n3248), .B(n4727), .Z(n8401) );
  XOR U8092 ( .A(n8402), .B(n8403), .Z(n4727) );
  ANDN U8093 ( .B(n8404), .A(n8405), .Z(n8402) );
  XOR U8094 ( .A(n8406), .B(n8407), .Z(n3248) );
  ANDN U8095 ( .B(n8408), .A(n8409), .Z(n8406) );
  XOR U8096 ( .A(n5551), .B(n8410), .Z(n8400) );
  XOR U8097 ( .A(n8411), .B(n2512), .Z(n8410) );
  XNOR U8098 ( .A(n8412), .B(n8413), .Z(n2512) );
  ANDN U8099 ( .B(n8414), .A(n8415), .Z(n8412) );
  XOR U8100 ( .A(n8416), .B(n8417), .Z(n5551) );
  ANDN U8101 ( .B(n8418), .A(n8419), .Z(n8416) );
  XOR U8102 ( .A(n8420), .B(n8421), .Z(n5832) );
  XNOR U8103 ( .A(n3817), .B(n5123), .Z(n8421) );
  XNOR U8104 ( .A(n8422), .B(n8423), .Z(n5123) );
  NOR U8105 ( .A(n8424), .B(n8425), .Z(n8422) );
  XOR U8106 ( .A(n8426), .B(n8427), .Z(n3817) );
  AND U8107 ( .A(n8428), .B(n8429), .Z(n8426) );
  XOR U8108 ( .A(n6307), .B(n8430), .Z(n8420) );
  XOR U8109 ( .A(n1751), .B(n8431), .Z(n8430) );
  XOR U8110 ( .A(n8432), .B(n8433), .Z(n1751) );
  XNOR U8111 ( .A(n8436), .B(n8437), .Z(n6307) );
  ANDN U8112 ( .B(n8438), .A(n8439), .Z(n8436) );
  XNOR U8113 ( .A(n1896), .B(n8440), .Z(n1140) );
  IV U8114 ( .A(n5212), .Z(n1896) );
  XOR U8115 ( .A(n7193), .B(n6092), .Z(n5212) );
  XOR U8116 ( .A(n8441), .B(n8442), .Z(n6092) );
  XNOR U8117 ( .A(n4542), .B(n1977), .Z(n8442) );
  XNOR U8118 ( .A(n8443), .B(n8444), .Z(n1977) );
  AND U8119 ( .A(n7334), .B(n7335), .Z(n8443) );
  IV U8120 ( .A(n8445), .Z(n7335) );
  XOR U8121 ( .A(n8446), .B(n8447), .Z(n4542) );
  XOR U8122 ( .A(n6000), .B(n8448), .Z(n8441) );
  XOR U8123 ( .A(n5542), .B(n3798), .Z(n8448) );
  XOR U8124 ( .A(n8449), .B(n8450), .Z(n3798) );
  NOR U8125 ( .A(n7330), .B(n7329), .Z(n8449) );
  XNOR U8126 ( .A(n8451), .B(n8452), .Z(n5542) );
  NOR U8127 ( .A(n7338), .B(n7339), .Z(n8451) );
  XOR U8128 ( .A(n8453), .B(n8454), .Z(n6000) );
  ANDN U8129 ( .B(n7325), .A(n7327), .Z(n8453) );
  XOR U8130 ( .A(n8455), .B(n8456), .Z(n7193) );
  XNOR U8131 ( .A(n4939), .B(n8457), .Z(n8456) );
  XNOR U8132 ( .A(n8458), .B(n7271), .Z(n4939) );
  ANDN U8133 ( .B(n8459), .A(n8372), .Z(n8458) );
  XOR U8134 ( .A(n2234), .B(n8460), .Z(n8455) );
  XNOR U8135 ( .A(n3543), .B(n6006), .Z(n8460) );
  XOR U8136 ( .A(n8461), .B(n7257), .Z(n6006) );
  AND U8137 ( .A(n8375), .B(n8462), .Z(n8461) );
  XNOR U8138 ( .A(n8463), .B(n7263), .Z(n3543) );
  ANDN U8139 ( .B(n8464), .A(n8370), .Z(n8463) );
  XOR U8140 ( .A(n8465), .B(n7253), .Z(n2234) );
  ANDN U8141 ( .B(n8379), .A(n8466), .Z(n8465) );
  XNOR U8142 ( .A(n8467), .B(n5963), .Z(out[1040]) );
  XNOR U8143 ( .A(n7431), .B(n2402), .Z(n5963) );
  XOR U8144 ( .A(n8468), .B(n8469), .Z(n7431) );
  ANDN U8145 ( .B(n8470), .A(n8471), .Z(n8468) );
  AND U8146 ( .A(n1144), .B(n1142), .Z(n8467) );
  XNOR U8147 ( .A(n2484), .B(n8472), .Z(n1142) );
  XOR U8148 ( .A(n5837), .B(n6250), .Z(n2484) );
  XOR U8149 ( .A(n8473), .B(n8474), .Z(n6250) );
  XNOR U8150 ( .A(n3251), .B(n4756), .Z(n8474) );
  XOR U8151 ( .A(n8475), .B(n8476), .Z(n4756) );
  AND U8152 ( .A(n8477), .B(n8427), .Z(n8475) );
  IV U8153 ( .A(n8478), .Z(n8427) );
  XOR U8154 ( .A(n8479), .B(n8480), .Z(n3251) );
  AND U8155 ( .A(n8481), .B(n8433), .Z(n8479) );
  IV U8156 ( .A(n8482), .Z(n8433) );
  XOR U8157 ( .A(n5246), .B(n8483), .Z(n8473) );
  XOR U8158 ( .A(n8484), .B(n2517), .Z(n8483) );
  XOR U8159 ( .A(n8485), .B(n8486), .Z(n2517) );
  NOR U8160 ( .A(n8487), .B(n8488), .Z(n8485) );
  XNOR U8161 ( .A(n8489), .B(n8490), .Z(n5246) );
  ANDN U8162 ( .B(n8491), .A(n8437), .Z(n8489) );
  XOR U8163 ( .A(n8492), .B(n8493), .Z(n5837) );
  XNOR U8164 ( .A(n3825), .B(n5125), .Z(n8493) );
  XNOR U8165 ( .A(n8494), .B(n8495), .Z(n5125) );
  ANDN U8166 ( .B(n8496), .A(n6375), .Z(n8494) );
  XOR U8167 ( .A(n8497), .B(n8498), .Z(n3825) );
  ANDN U8168 ( .B(n8499), .A(n6362), .Z(n8497) );
  XNOR U8169 ( .A(n8500), .B(n8501), .Z(n8492) );
  XNOR U8170 ( .A(n4230), .B(n1757), .Z(n8501) );
  XNOR U8171 ( .A(n8502), .B(n8503), .Z(n1757) );
  AND U8172 ( .A(n8504), .B(n6366), .Z(n8502) );
  IV U8173 ( .A(n8505), .Z(n6366) );
  XOR U8174 ( .A(n8506), .B(n8507), .Z(n4230) );
  ANDN U8175 ( .B(n8508), .A(n6379), .Z(n8506) );
  XNOR U8176 ( .A(n1900), .B(n8509), .Z(n1144) );
  IV U8177 ( .A(n5215), .Z(n1900) );
  XOR U8178 ( .A(n7248), .B(n6097), .Z(n5215) );
  XOR U8179 ( .A(n8510), .B(n8511), .Z(n6097) );
  XOR U8180 ( .A(n4588), .B(n1980), .Z(n8511) );
  XOR U8181 ( .A(n8512), .B(n8513), .Z(n1980) );
  AND U8182 ( .A(n7411), .B(n7412), .Z(n8512) );
  XNOR U8183 ( .A(n8514), .B(n8515), .Z(n4588) );
  NOR U8184 ( .A(n7421), .B(n7419), .Z(n8514) );
  IV U8185 ( .A(n8516), .Z(n7421) );
  XOR U8186 ( .A(n6010), .B(n8517), .Z(n8510) );
  XOR U8187 ( .A(n5546), .B(n3801), .Z(n8517) );
  XNOR U8188 ( .A(n8518), .B(n8519), .Z(n3801) );
  AND U8189 ( .A(n7408), .B(n7406), .Z(n8518) );
  AND U8190 ( .A(n7415), .B(n7417), .Z(n8520) );
  XOR U8191 ( .A(n8522), .B(n8523), .Z(n6010) );
  ANDN U8192 ( .B(n7404), .A(n7402), .Z(n8522) );
  XOR U8193 ( .A(n8524), .B(n8525), .Z(n7248) );
  XOR U8194 ( .A(n4946), .B(n8526), .Z(n8525) );
  XOR U8195 ( .A(n8527), .B(n7343), .Z(n4946) );
  AND U8196 ( .A(n8528), .B(n8447), .Z(n8527) );
  IV U8197 ( .A(n8529), .Z(n8447) );
  XOR U8198 ( .A(n2239), .B(n8530), .Z(n8524) );
  XOR U8199 ( .A(n3545), .B(n6058), .Z(n8530) );
  XOR U8200 ( .A(n8531), .B(n7331), .Z(n6058) );
  AND U8201 ( .A(n8532), .B(n8450), .Z(n8531) );
  IV U8202 ( .A(n8533), .Z(n8450) );
  XNOR U8203 ( .A(n8534), .B(n7336), .Z(n3545) );
  ANDN U8204 ( .B(n8535), .A(n8444), .Z(n8534) );
  XOR U8205 ( .A(n8536), .B(n7326), .Z(n2239) );
  NOR U8206 ( .A(n8537), .B(n8454), .Z(n8536) );
  XNOR U8207 ( .A(n8538), .B(n4152), .Z(out[103]) );
  XNOR U8208 ( .A(n8539), .B(n2548), .Z(n4152) );
  XNOR U8209 ( .A(n7794), .B(n8540), .Z(n2548) );
  XOR U8210 ( .A(n8541), .B(n8542), .Z(n7794) );
  XNOR U8211 ( .A(n4329), .B(n2171), .Z(n8542) );
  XNOR U8212 ( .A(n8543), .B(n7899), .Z(n2171) );
  ANDN U8213 ( .B(n8544), .A(n8545), .Z(n8543) );
  XNOR U8214 ( .A(n8546), .B(n7890), .Z(n4329) );
  ANDN U8215 ( .B(n8547), .A(n8548), .Z(n8546) );
  XOR U8216 ( .A(n5945), .B(n8549), .Z(n8541) );
  XNOR U8217 ( .A(n5499), .B(n3746), .Z(n8549) );
  XNOR U8218 ( .A(n8550), .B(n7895), .Z(n3746) );
  ANDN U8219 ( .B(n8551), .A(n8552), .Z(n8550) );
  XOR U8220 ( .A(n8553), .B(n8554), .Z(n5499) );
  AND U8221 ( .A(n8555), .B(n8556), .Z(n8553) );
  XOR U8222 ( .A(n8557), .B(n7902), .Z(n5945) );
  ANDN U8223 ( .B(n8558), .A(n8559), .Z(n8557) );
  ANDN U8224 ( .B(n3512), .A(n3510), .Z(n8538) );
  XOR U8225 ( .A(n7304), .B(n2390), .Z(n3510) );
  XNOR U8226 ( .A(n8560), .B(n8561), .Z(n2390) );
  XNOR U8227 ( .A(n8562), .B(n8563), .Z(n7304) );
  AND U8228 ( .A(n8564), .B(n8565), .Z(n8562) );
  XOR U8229 ( .A(n2320), .B(n8566), .Z(n3512) );
  XOR U8230 ( .A(n6147), .B(n8567), .Z(n2320) );
  XOR U8231 ( .A(n8568), .B(n8569), .Z(n6147) );
  XNOR U8232 ( .A(n3173), .B(n6576), .Z(n8569) );
  XOR U8233 ( .A(n8570), .B(n8571), .Z(n6576) );
  ANDN U8234 ( .B(n8572), .A(n8573), .Z(n8570) );
  XNOR U8235 ( .A(n8574), .B(n8575), .Z(n3173) );
  NOR U8236 ( .A(n8576), .B(n8577), .Z(n8574) );
  XOR U8237 ( .A(n5455), .B(n8578), .Z(n8568) );
  XOR U8238 ( .A(n8124), .B(n2355), .Z(n8578) );
  XOR U8239 ( .A(n8579), .B(n8580), .Z(n2355) );
  ANDN U8240 ( .B(n8581), .A(n8582), .Z(n8579) );
  XOR U8241 ( .A(n8583), .B(n8584), .Z(n8124) );
  NOR U8242 ( .A(n8585), .B(n8586), .Z(n8583) );
  XOR U8243 ( .A(n8587), .B(n8588), .Z(n5455) );
  AND U8244 ( .A(n8589), .B(n8590), .Z(n8587) );
  XOR U8245 ( .A(n8591), .B(n5968), .Z(out[1039]) );
  XOR U8246 ( .A(n7538), .B(n2411), .Z(n5968) );
  XNOR U8247 ( .A(n8592), .B(n8593), .Z(n7538) );
  AND U8248 ( .A(n8594), .B(n8595), .Z(n8592) );
  AND U8249 ( .A(n1147), .B(n1146), .Z(n8591) );
  XNOR U8250 ( .A(n8596), .B(n2492), .Z(n1146) );
  XOR U8251 ( .A(n5847), .B(n6254), .Z(n2492) );
  XOR U8252 ( .A(n8597), .B(n8598), .Z(n6254) );
  XNOR U8253 ( .A(n3254), .B(n4784), .Z(n8598) );
  XOR U8254 ( .A(n8599), .B(n6363), .Z(n4784) );
  ANDN U8255 ( .B(n6364), .A(n8498), .Z(n8599) );
  XNOR U8256 ( .A(n8600), .B(n6368), .Z(n3254) );
  AND U8257 ( .A(n6367), .B(n8503), .Z(n8600) );
  XOR U8258 ( .A(n5250), .B(n8601), .Z(n8597) );
  XOR U8259 ( .A(n6357), .B(n2530), .Z(n8601) );
  XOR U8260 ( .A(n8602), .B(n6372), .Z(n2530) );
  AND U8261 ( .A(n8603), .B(n6373), .Z(n8602) );
  XOR U8262 ( .A(n8604), .B(n6376), .Z(n6357) );
  AND U8263 ( .A(n6377), .B(n8495), .Z(n8604) );
  XNOR U8264 ( .A(n8605), .B(n6380), .Z(n5250) );
  ANDN U8265 ( .B(n6381), .A(n8507), .Z(n8605) );
  XOR U8266 ( .A(n8606), .B(n8607), .Z(n5847) );
  XNOR U8267 ( .A(n3831), .B(n5127), .Z(n8607) );
  XOR U8268 ( .A(n8608), .B(n8609), .Z(n5127) );
  ANDN U8269 ( .B(n8610), .A(n6401), .Z(n8608) );
  XNOR U8270 ( .A(n8611), .B(n8612), .Z(n3831) );
  AND U8271 ( .A(n6388), .B(n8613), .Z(n8611) );
  XOR U8272 ( .A(n4233), .B(n8614), .Z(n8606) );
  XOR U8273 ( .A(n1761), .B(n8615), .Z(n8614) );
  XNOR U8274 ( .A(n8616), .B(n8617), .Z(n1761) );
  XOR U8275 ( .A(n8619), .B(n8620), .Z(n4233) );
  ANDN U8276 ( .B(n8621), .A(n6405), .Z(n8619) );
  XNOR U8277 ( .A(n1904), .B(n8622), .Z(n1147) );
  IV U8278 ( .A(n3656), .Z(n1904) );
  XOR U8279 ( .A(n7321), .B(n6102), .Z(n3656) );
  XOR U8280 ( .A(n8623), .B(n8624), .Z(n6102) );
  XNOR U8281 ( .A(n4633), .B(n1983), .Z(n8624) );
  XOR U8282 ( .A(n8625), .B(n8626), .Z(n1983) );
  AND U8283 ( .A(n7485), .B(n7486), .Z(n8625) );
  XNOR U8284 ( .A(n8627), .B(n8628), .Z(n4633) );
  XNOR U8285 ( .A(n6015), .B(n8629), .Z(n8623) );
  XOR U8286 ( .A(n5550), .B(n3807), .Z(n8629) );
  XOR U8287 ( .A(n8630), .B(n8631), .Z(n3807) );
  AND U8288 ( .A(n7482), .B(n7480), .Z(n8630) );
  XOR U8289 ( .A(n8632), .B(n8633), .Z(n5550) );
  NOR U8290 ( .A(n7489), .B(n7490), .Z(n8632) );
  XNOR U8291 ( .A(n8634), .B(n8635), .Z(n6015) );
  AND U8292 ( .A(n7476), .B(n7478), .Z(n8634) );
  XOR U8293 ( .A(n8636), .B(n8637), .Z(n7321) );
  XNOR U8294 ( .A(n4949), .B(n8638), .Z(n8637) );
  XOR U8295 ( .A(n8639), .B(n7420), .Z(n4949) );
  NOR U8296 ( .A(n8640), .B(n8515), .Z(n8639) );
  XNOR U8297 ( .A(n2246), .B(n8641), .Z(n8636) );
  XNOR U8298 ( .A(n3547), .B(n6112), .Z(n8641) );
  XNOR U8299 ( .A(n8642), .B(n7407), .Z(n6112) );
  ANDN U8300 ( .B(n8643), .A(n8519), .Z(n8642) );
  XNOR U8301 ( .A(n8644), .B(n7413), .Z(n3547) );
  ANDN U8302 ( .B(n8513), .A(n8645), .Z(n8644) );
  XNOR U8303 ( .A(n8646), .B(n7403), .Z(n2246) );
  XNOR U8304 ( .A(n8648), .B(n5973), .Z(out[1038]) );
  XNOR U8305 ( .A(n4336), .B(n7605), .Z(n5973) );
  XOR U8306 ( .A(n8649), .B(n8650), .Z(n7605) );
  ANDN U8307 ( .B(n8651), .A(n8652), .Z(n8649) );
  XOR U8308 ( .A(n8653), .B(n8654), .Z(n4336) );
  AND U8309 ( .A(n1151), .B(n1150), .Z(n8648) );
  XNOR U8310 ( .A(n4354), .B(n8655), .Z(n1150) );
  XOR U8311 ( .A(n5852), .B(n6263), .Z(n4354) );
  XOR U8312 ( .A(n8656), .B(n8657), .Z(n6263) );
  XOR U8313 ( .A(n3257), .B(n4808), .Z(n8657) );
  XOR U8314 ( .A(n8658), .B(n6389), .Z(n4808) );
  ANDN U8315 ( .B(n6390), .A(n8612), .Z(n8658) );
  XNOR U8316 ( .A(n8659), .B(n6393), .Z(n3257) );
  ANDN U8317 ( .B(n6394), .A(n8617), .Z(n8659) );
  XOR U8318 ( .A(n5255), .B(n8660), .Z(n8656) );
  XNOR U8319 ( .A(n6383), .B(n2537), .Z(n8660) );
  XNOR U8320 ( .A(n8661), .B(n6398), .Z(n2537) );
  AND U8321 ( .A(n6399), .B(n8662), .Z(n8661) );
  XNOR U8322 ( .A(n8663), .B(n6402), .Z(n6383) );
  AND U8323 ( .A(n6403), .B(n8609), .Z(n8663) );
  IV U8324 ( .A(n8664), .Z(n8609) );
  XNOR U8325 ( .A(n8665), .B(n6407), .Z(n5255) );
  ANDN U8326 ( .B(n8620), .A(n6406), .Z(n8665) );
  IV U8327 ( .A(n8666), .Z(n8620) );
  XOR U8328 ( .A(n8667), .B(n8668), .Z(n5852) );
  XNOR U8329 ( .A(n3835), .B(n5130), .Z(n8668) );
  XNOR U8330 ( .A(n8669), .B(n8670), .Z(n5130) );
  ANDN U8331 ( .B(n6428), .A(n8671), .Z(n8669) );
  IV U8332 ( .A(n8672), .Z(n6428) );
  XOR U8333 ( .A(n8673), .B(n8674), .Z(n3835) );
  ANDN U8334 ( .B(n6415), .A(n8675), .Z(n8673) );
  IV U8335 ( .A(n8676), .Z(n6415) );
  XNOR U8336 ( .A(n4241), .B(n8677), .Z(n8667) );
  XNOR U8337 ( .A(n1769), .B(n8678), .Z(n8677) );
  XNOR U8338 ( .A(n8679), .B(n8680), .Z(n1769) );
  AND U8339 ( .A(n8681), .B(n6419), .Z(n8679) );
  XNOR U8340 ( .A(n8682), .B(n8683), .Z(n4241) );
  AND U8341 ( .A(n8684), .B(n6432), .Z(n8682) );
  IV U8342 ( .A(n8685), .Z(n6432) );
  XNOR U8343 ( .A(n1912), .B(n8686), .Z(n1151) );
  IV U8344 ( .A(n5220), .Z(n1912) );
  XOR U8345 ( .A(n7398), .B(n6107), .Z(n5220) );
  XOR U8346 ( .A(n8687), .B(n8688), .Z(n6107) );
  XNOR U8347 ( .A(n4673), .B(n1986), .Z(n8688) );
  XOR U8348 ( .A(n8689), .B(n8690), .Z(n1986) );
  ANDN U8349 ( .B(n7562), .A(n7563), .Z(n8689) );
  XOR U8350 ( .A(n8691), .B(n8692), .Z(n4673) );
  ANDN U8351 ( .B(n7571), .A(n7570), .Z(n8691) );
  XNOR U8352 ( .A(n6020), .B(n8693), .Z(n8687) );
  XOR U8353 ( .A(n5245), .B(n3812), .Z(n8693) );
  XNOR U8354 ( .A(n8694), .B(n8695), .Z(n3812) );
  XOR U8355 ( .A(n8696), .B(n8697), .Z(n5245) );
  NOR U8356 ( .A(n7567), .B(n7566), .Z(n8696) );
  XNOR U8357 ( .A(n8698), .B(n8699), .Z(n6020) );
  NOR U8358 ( .A(n8700), .B(n7554), .Z(n8698) );
  XOR U8359 ( .A(n8701), .B(n8702), .Z(n7398) );
  XOR U8360 ( .A(n4952), .B(n8703), .Z(n8702) );
  XOR U8361 ( .A(n8704), .B(n7495), .Z(n4952) );
  ANDN U8362 ( .B(n8705), .A(n8628), .Z(n8704) );
  XOR U8363 ( .A(n2253), .B(n8706), .Z(n8701) );
  XOR U8364 ( .A(n3549), .B(n6167), .Z(n8706) );
  XNOR U8365 ( .A(n8707), .B(n7481), .Z(n6167) );
  ANDN U8366 ( .B(n8708), .A(n8631), .Z(n8707) );
  XOR U8367 ( .A(n8709), .B(n7487), .Z(n3549) );
  AND U8368 ( .A(n8710), .B(n8626), .Z(n8709) );
  XOR U8369 ( .A(n8711), .B(n7477), .Z(n2253) );
  XOR U8370 ( .A(n8713), .B(n5978), .Z(out[1037]) );
  XOR U8371 ( .A(n2424), .B(n7653), .Z(n5978) );
  XNOR U8372 ( .A(n8714), .B(n8715), .Z(n7653) );
  NOR U8373 ( .A(n8716), .B(n8717), .Z(n8714) );
  XOR U8374 ( .A(n8718), .B(n8719), .Z(n2424) );
  ANDN U8375 ( .B(n1154), .A(n1156), .Z(n8713) );
  XNOR U8376 ( .A(n1917), .B(n8720), .Z(n1156) );
  IV U8377 ( .A(n5223), .Z(n1917) );
  XOR U8378 ( .A(n7472), .B(n6117), .Z(n5223) );
  XOR U8379 ( .A(n8721), .B(n8722), .Z(n6117) );
  XOR U8380 ( .A(n4698), .B(n1989), .Z(n8722) );
  XOR U8381 ( .A(n8723), .B(n8724), .Z(n1989) );
  XNOR U8382 ( .A(n8725), .B(n8726), .Z(n4698) );
  NOR U8383 ( .A(n7647), .B(n7646), .Z(n8725) );
  XOR U8384 ( .A(n6025), .B(n8727), .Z(n8721) );
  XOR U8385 ( .A(n5249), .B(n3819), .Z(n8727) );
  XOR U8386 ( .A(n8728), .B(n8729), .Z(n3819) );
  XOR U8387 ( .A(n8730), .B(n8731), .Z(n5249) );
  NOR U8388 ( .A(n7642), .B(n7644), .Z(n8730) );
  XOR U8389 ( .A(n8732), .B(n8733), .Z(n6025) );
  AND U8390 ( .A(n7630), .B(n7629), .Z(n8732) );
  IV U8391 ( .A(n8734), .Z(n7629) );
  XOR U8392 ( .A(n8735), .B(n8736), .Z(n7472) );
  XOR U8393 ( .A(n4955), .B(n8737), .Z(n8736) );
  XNOR U8394 ( .A(n8738), .B(n7572), .Z(n4955) );
  AND U8395 ( .A(n8692), .B(n8739), .Z(n8738) );
  XOR U8396 ( .A(n2262), .B(n8740), .Z(n8735) );
  XOR U8397 ( .A(n3551), .B(n6213), .Z(n8740) );
  XNOR U8398 ( .A(n8741), .B(n7558), .Z(n6213) );
  NOR U8399 ( .A(n8742), .B(n8695), .Z(n8741) );
  XNOR U8400 ( .A(n8743), .B(n7564), .Z(n3551) );
  AND U8401 ( .A(n8690), .B(n8744), .Z(n8743) );
  XNOR U8402 ( .A(n8745), .B(n7555), .Z(n2262) );
  NOR U8403 ( .A(n8746), .B(n8699), .Z(n8745) );
  XNOR U8404 ( .A(n2503), .B(n8747), .Z(n1154) );
  XOR U8405 ( .A(n5857), .B(n6268), .Z(n2503) );
  XNOR U8406 ( .A(n8748), .B(n8749), .Z(n6268) );
  XOR U8407 ( .A(n2542), .B(n5259), .Z(n8749) );
  XNOR U8408 ( .A(n8750), .B(n6434), .Z(n5259) );
  NOR U8409 ( .A(n6433), .B(n8683), .Z(n8750) );
  XOR U8410 ( .A(n8751), .B(n6425), .Z(n2542) );
  IV U8411 ( .A(n8752), .Z(n6425) );
  AND U8412 ( .A(n6426), .B(n8753), .Z(n8751) );
  XOR U8413 ( .A(n3261), .B(n8754), .Z(n8748) );
  XOR U8414 ( .A(n4835), .B(n6410), .Z(n8754) );
  XNOR U8415 ( .A(n8755), .B(n6429), .Z(n6410) );
  ANDN U8416 ( .B(n6430), .A(n8670), .Z(n8755) );
  XNOR U8417 ( .A(n8756), .B(n6416), .Z(n4835) );
  AND U8418 ( .A(n8674), .B(n6417), .Z(n8756) );
  XOR U8419 ( .A(n8757), .B(n6420), .Z(n3261) );
  ANDN U8420 ( .B(n8758), .A(n8680), .Z(n8757) );
  XOR U8421 ( .A(n8759), .B(n8760), .Z(n5857) );
  XNOR U8422 ( .A(n3841), .B(n5133), .Z(n8760) );
  XOR U8423 ( .A(n8761), .B(n8762), .Z(n5133) );
  NOR U8424 ( .A(n8763), .B(n6459), .Z(n8761) );
  XNOR U8425 ( .A(n8764), .B(n8765), .Z(n3841) );
  ANDN U8426 ( .B(n8766), .A(n6442), .Z(n8764) );
  XOR U8427 ( .A(n4244), .B(n8767), .Z(n8759) );
  XOR U8428 ( .A(n1774), .B(n8768), .Z(n8767) );
  XOR U8429 ( .A(n8769), .B(n8770), .Z(n1774) );
  ANDN U8430 ( .B(n8771), .A(n8772), .Z(n8769) );
  XNOR U8431 ( .A(n8773), .B(n8774), .Z(n4244) );
  ANDN U8432 ( .B(n8775), .A(n6463), .Z(n8773) );
  XOR U8433 ( .A(n8776), .B(n5983), .Z(out[1036]) );
  XNOR U8434 ( .A(n7739), .B(n4346), .Z(n5983) );
  IV U8435 ( .A(n2430), .Z(n4346) );
  XNOR U8436 ( .A(n8777), .B(n8778), .Z(n2430) );
  XOR U8437 ( .A(n8779), .B(n8780), .Z(n7739) );
  NOR U8438 ( .A(n8781), .B(n8782), .Z(n8779) );
  ANDN U8439 ( .B(n1158), .A(n1160), .Z(n8776) );
  XNOR U8440 ( .A(n1921), .B(n8783), .Z(n1160) );
  IV U8441 ( .A(n5231), .Z(n1921) );
  XOR U8442 ( .A(n7549), .B(n6122), .Z(n5231) );
  XOR U8443 ( .A(n8784), .B(n8785), .Z(n6122) );
  XOR U8444 ( .A(n4725), .B(n1996), .Z(n8785) );
  XNOR U8445 ( .A(n8786), .B(n8787), .Z(n1996) );
  AND U8446 ( .A(n7715), .B(n7717), .Z(n8786) );
  XOR U8447 ( .A(n8788), .B(n8789), .Z(n4725) );
  ANDN U8448 ( .B(n7723), .A(n7724), .Z(n8788) );
  XOR U8449 ( .A(n6030), .B(n8790), .Z(n8784) );
  XOR U8450 ( .A(n5253), .B(n3827), .Z(n8790) );
  XOR U8451 ( .A(n8791), .B(n8792), .Z(n3827) );
  XOR U8452 ( .A(n8793), .B(n8794), .Z(n5253) );
  AND U8453 ( .A(n7719), .B(n7721), .Z(n8793) );
  XOR U8454 ( .A(n8795), .B(n8796), .Z(n6030) );
  ANDN U8455 ( .B(n7706), .A(n7707), .Z(n8795) );
  XOR U8456 ( .A(n8797), .B(n8798), .Z(n7549) );
  XOR U8457 ( .A(n4958), .B(n8799), .Z(n8798) );
  XNOR U8458 ( .A(n8800), .B(n7648), .Z(n4958) );
  ANDN U8459 ( .B(n8801), .A(n8802), .Z(n8800) );
  XOR U8460 ( .A(n2269), .B(n8803), .Z(n8797) );
  XOR U8461 ( .A(n3370), .B(n6259), .Z(n8803) );
  XOR U8462 ( .A(n8804), .B(n7635), .Z(n6259) );
  IV U8463 ( .A(n8805), .Z(n7635) );
  ANDN U8464 ( .B(n8729), .A(n8806), .Z(n8804) );
  XOR U8465 ( .A(n8807), .B(n7639), .Z(n3370) );
  AND U8466 ( .A(n8724), .B(n8808), .Z(n8807) );
  XOR U8467 ( .A(n8809), .B(n7631), .Z(n2269) );
  ANDN U8468 ( .B(n8810), .A(n8733), .Z(n8809) );
  XNOR U8469 ( .A(n2510), .B(n8811), .Z(n1158) );
  IV U8470 ( .A(n3465), .Z(n2510) );
  XOR U8471 ( .A(n5862), .B(n6272), .Z(n3465) );
  XOR U8472 ( .A(n8812), .B(n8813), .Z(n6272) );
  XOR U8473 ( .A(n3264), .B(n4872), .Z(n8813) );
  XOR U8474 ( .A(n8814), .B(n6443), .Z(n4872) );
  ANDN U8475 ( .B(n6444), .A(n8765), .Z(n8814) );
  XNOR U8476 ( .A(n8815), .B(n6447), .Z(n3264) );
  AND U8477 ( .A(n8770), .B(n6448), .Z(n8815) );
  IV U8478 ( .A(n8816), .Z(n8770) );
  XNOR U8479 ( .A(n5267), .B(n8817), .Z(n8812) );
  XNOR U8480 ( .A(n6437), .B(n2549), .Z(n8817) );
  XNOR U8481 ( .A(n8818), .B(n6456), .Z(n2549) );
  AND U8482 ( .A(n6457), .B(n8819), .Z(n8818) );
  XOR U8483 ( .A(n8820), .B(n6460), .Z(n6437) );
  AND U8484 ( .A(n8762), .B(n6461), .Z(n8820) );
  IV U8485 ( .A(n8821), .Z(n8762) );
  XNOR U8486 ( .A(n8822), .B(n6465), .Z(n5267) );
  NOR U8487 ( .A(n8774), .B(n6464), .Z(n8822) );
  XOR U8488 ( .A(n8823), .B(n8824), .Z(n5862) );
  XOR U8489 ( .A(n3847), .B(n5141), .Z(n8824) );
  XOR U8490 ( .A(n8825), .B(n8826), .Z(n5141) );
  AND U8491 ( .A(n8827), .B(n6485), .Z(n8825) );
  XNOR U8492 ( .A(n8828), .B(n8829), .Z(n3847) );
  ANDN U8493 ( .B(n6472), .A(n8830), .Z(n8828) );
  IV U8494 ( .A(n8831), .Z(n6472) );
  XOR U8495 ( .A(n4246), .B(n8832), .Z(n8823) );
  XOR U8496 ( .A(n1779), .B(n8833), .Z(n8832) );
  XOR U8497 ( .A(n8834), .B(n8835), .Z(n1779) );
  NOR U8498 ( .A(n6476), .B(n8836), .Z(n8834) );
  XOR U8499 ( .A(n8837), .B(n8838), .Z(n4246) );
  NOR U8500 ( .A(n6489), .B(n8839), .Z(n8837) );
  XOR U8501 ( .A(n8840), .B(n5988), .Z(out[1035]) );
  XOR U8502 ( .A(n7825), .B(n3211), .Z(n5988) );
  XNOR U8503 ( .A(n8843), .B(n8844), .Z(n7825) );
  AND U8504 ( .A(n8845), .B(n8846), .Z(n8843) );
  ANDN U8505 ( .B(n1162), .A(n1164), .Z(n8840) );
  XNOR U8506 ( .A(n1926), .B(n8847), .Z(n1164) );
  IV U8507 ( .A(n4154), .Z(n1926) );
  XOR U8508 ( .A(n7625), .B(n6127), .Z(n4154) );
  XOR U8509 ( .A(n8848), .B(n8849), .Z(n6127) );
  XNOR U8510 ( .A(n4755), .B(n1999), .Z(n8849) );
  XOR U8511 ( .A(n8850), .B(n8851), .Z(n1999) );
  ANDN U8512 ( .B(n7784), .A(n7782), .Z(n8850) );
  XOR U8513 ( .A(n8852), .B(n8853), .Z(n4755) );
  NOR U8514 ( .A(n7790), .B(n7791), .Z(n8852) );
  XNOR U8515 ( .A(n6036), .B(n8854), .Z(n8848) );
  XNOR U8516 ( .A(n5257), .B(n3833), .Z(n8854) );
  XNOR U8517 ( .A(n8855), .B(n8856), .Z(n3833) );
  ANDN U8518 ( .B(n7779), .A(n7777), .Z(n8855) );
  XNOR U8519 ( .A(n8857), .B(n8858), .Z(n5257) );
  ANDN U8520 ( .B(n7786), .A(n7787), .Z(n8857) );
  XNOR U8521 ( .A(n8859), .B(n8860), .Z(n6036) );
  ANDN U8522 ( .B(n7773), .A(n7775), .Z(n8859) );
  XOR U8523 ( .A(n8861), .B(n8862), .Z(n7625) );
  XOR U8524 ( .A(n4961), .B(n8863), .Z(n8862) );
  XNOR U8525 ( .A(n8864), .B(n7725), .Z(n4961) );
  NOR U8526 ( .A(n8865), .B(n8789), .Z(n8864) );
  XNOR U8527 ( .A(n2274), .B(n8866), .Z(n8861) );
  XOR U8528 ( .A(n3372), .B(n6311), .Z(n8866) );
  XOR U8529 ( .A(n8867), .B(n7711), .Z(n6311) );
  IV U8530 ( .A(n8868), .Z(n7711) );
  ANDN U8531 ( .B(n8792), .A(n8869), .Z(n8867) );
  XOR U8532 ( .A(n8870), .B(n7716), .Z(n3372) );
  NOR U8533 ( .A(n8871), .B(n8787), .Z(n8870) );
  XNOR U8534 ( .A(n8872), .B(n7708), .Z(n2274) );
  AND U8535 ( .A(n8796), .B(n8873), .Z(n8872) );
  XOR U8536 ( .A(n3468), .B(n8874), .Z(n1162) );
  XOR U8537 ( .A(n5866), .B(n6277), .Z(n3468) );
  XOR U8538 ( .A(n8875), .B(n8876), .Z(n6277) );
  XOR U8539 ( .A(n3269), .B(n4906), .Z(n8876) );
  XNOR U8540 ( .A(n8877), .B(n6473), .Z(n4906) );
  AND U8541 ( .A(n6474), .B(n8878), .Z(n8877) );
  XNOR U8542 ( .A(n8879), .B(n6477), .Z(n3269) );
  AND U8543 ( .A(n8835), .B(n6478), .Z(n8879) );
  XNOR U8544 ( .A(n5273), .B(n8880), .Z(n8875) );
  XOR U8545 ( .A(n6467), .B(n2556), .Z(n8880) );
  XOR U8546 ( .A(n8881), .B(n6482), .Z(n2556) );
  XOR U8547 ( .A(n8883), .B(n6486), .Z(n6467) );
  ANDN U8548 ( .B(n8826), .A(n6487), .Z(n8883) );
  XNOR U8549 ( .A(n8884), .B(n6490), .Z(n5273) );
  AND U8550 ( .A(n6491), .B(n8838), .Z(n8884) );
  IV U8551 ( .A(n8885), .Z(n8838) );
  XOR U8552 ( .A(n8886), .B(n8887), .Z(n5866) );
  XNOR U8553 ( .A(n3852), .B(n5144), .Z(n8887) );
  XOR U8554 ( .A(n8888), .B(n8889), .Z(n5144) );
  ANDN U8555 ( .B(n6511), .A(n8890), .Z(n8888) );
  IV U8556 ( .A(n8891), .Z(n6511) );
  XOR U8557 ( .A(n8892), .B(n8893), .Z(n3852) );
  ANDN U8558 ( .B(n6498), .A(n8894), .Z(n8892) );
  IV U8559 ( .A(n8895), .Z(n6498) );
  XNOR U8560 ( .A(n4248), .B(n8896), .Z(n8886) );
  XOR U8561 ( .A(n1783), .B(n8897), .Z(n8896) );
  XOR U8562 ( .A(n8898), .B(n8899), .Z(n1783) );
  ANDN U8563 ( .B(n8900), .A(n6502), .Z(n8898) );
  XNOR U8564 ( .A(n8901), .B(n8902), .Z(n4248) );
  AND U8565 ( .A(n8903), .B(n6515), .Z(n8901) );
  XOR U8566 ( .A(n8904), .B(n5993), .Z(out[1034]) );
  XOR U8567 ( .A(n7873), .B(n3215), .Z(n5993) );
  XNOR U8568 ( .A(n8905), .B(n8906), .Z(n3215) );
  XNOR U8569 ( .A(n8907), .B(n8908), .Z(n7873) );
  AND U8570 ( .A(n8909), .B(n8910), .Z(n8907) );
  ANDN U8571 ( .B(n1166), .A(n1168), .Z(n8904) );
  XNOR U8572 ( .A(n1930), .B(n8911), .Z(n1168) );
  IV U8573 ( .A(n5236), .Z(n1930) );
  XOR U8574 ( .A(n7702), .B(n6132), .Z(n5236) );
  XOR U8575 ( .A(n8912), .B(n8913), .Z(n6132) );
  XNOR U8576 ( .A(n4782), .B(n2002), .Z(n8913) );
  XOR U8577 ( .A(n8914), .B(n8915), .Z(n2002) );
  XOR U8578 ( .A(n8916), .B(n8917), .Z(n4782) );
  XOR U8579 ( .A(n6041), .B(n8918), .Z(n8912) );
  XNOR U8580 ( .A(n5266), .B(n3836), .Z(n8918) );
  XOR U8581 ( .A(n8919), .B(n8920), .Z(n3836) );
  XNOR U8582 ( .A(n8921), .B(n8922), .Z(n5266) );
  ANDN U8583 ( .B(n7853), .A(n7855), .Z(n8921) );
  XOR U8584 ( .A(n8923), .B(n8924), .Z(n6041) );
  NOR U8585 ( .A(n7842), .B(n7840), .Z(n8923) );
  XOR U8586 ( .A(n8925), .B(n8926), .Z(n7702) );
  XNOR U8587 ( .A(n4964), .B(n8927), .Z(n8926) );
  XNOR U8588 ( .A(n8928), .B(n7792), .Z(n4964) );
  ANDN U8589 ( .B(n8853), .A(n8929), .Z(n8928) );
  XOR U8590 ( .A(n2281), .B(n8930), .Z(n8925) );
  XOR U8591 ( .A(n3374), .B(n6349), .Z(n8930) );
  XOR U8592 ( .A(n8931), .B(n7778), .Z(n6349) );
  ANDN U8593 ( .B(n8932), .A(n8856), .Z(n8931) );
  XNOR U8594 ( .A(n8933), .B(n7783), .Z(n3374) );
  XOR U8595 ( .A(n8935), .B(n7774), .Z(n2281) );
  XNOR U8596 ( .A(n4854), .B(n8937), .Z(n1166) );
  XOR U8597 ( .A(n5871), .B(n6282), .Z(n4854) );
  XOR U8598 ( .A(n8938), .B(n8939), .Z(n6282) );
  XNOR U8599 ( .A(n3272), .B(n4944), .Z(n8939) );
  XOR U8600 ( .A(n8940), .B(n6499), .Z(n4944) );
  AND U8601 ( .A(n8893), .B(n6500), .Z(n8940) );
  XOR U8602 ( .A(n8941), .B(n6503), .Z(n3272) );
  ANDN U8603 ( .B(n8942), .A(n8899), .Z(n8941) );
  XOR U8604 ( .A(n5278), .B(n8943), .Z(n8938) );
  XOR U8605 ( .A(n6493), .B(n2565), .Z(n8943) );
  XOR U8606 ( .A(n8944), .B(n6508), .Z(n2565) );
  AND U8607 ( .A(n6509), .B(n8945), .Z(n8944) );
  XOR U8608 ( .A(n8946), .B(n6512), .Z(n6493) );
  AND U8609 ( .A(n6513), .B(n8889), .Z(n8946) );
  IV U8610 ( .A(n8947), .Z(n8889) );
  XNOR U8611 ( .A(n8948), .B(n6516), .Z(n5278) );
  ANDN U8612 ( .B(n6517), .A(n8902), .Z(n8948) );
  XOR U8613 ( .A(n8949), .B(n8950), .Z(n5871) );
  XOR U8614 ( .A(n3856), .B(n5147), .Z(n8950) );
  XNOR U8615 ( .A(n8951), .B(n8952), .Z(n5147) );
  ANDN U8616 ( .B(n8953), .A(n6533), .Z(n8951) );
  XOR U8617 ( .A(n8954), .B(n8955), .Z(n3856) );
  ANDN U8618 ( .B(n6537), .A(n8956), .Z(n8954) );
  IV U8619 ( .A(n8957), .Z(n6537) );
  XOR U8620 ( .A(n4252), .B(n8958), .Z(n8949) );
  XNOR U8621 ( .A(n1787), .B(n8959), .Z(n8958) );
  XOR U8622 ( .A(n8960), .B(n8961), .Z(n1787) );
  NOR U8623 ( .A(n6541), .B(n8962), .Z(n8960) );
  XOR U8624 ( .A(n8963), .B(n8964), .Z(n4252) );
  AND U8625 ( .A(n8965), .B(n6524), .Z(n8963) );
  IV U8626 ( .A(n8966), .Z(n6524) );
  XOR U8627 ( .A(n8967), .B(n5998), .Z(out[1033]) );
  XNOR U8628 ( .A(n7982), .B(n2455), .Z(n5998) );
  XOR U8629 ( .A(n8970), .B(n8971), .Z(n7982) );
  NOR U8630 ( .A(n8972), .B(n8973), .Z(n8970) );
  AND U8631 ( .A(n1174), .B(n1176), .Z(n8967) );
  XNOR U8632 ( .A(n1934), .B(n8974), .Z(n1176) );
  IV U8633 ( .A(n3689), .Z(n1934) );
  XOR U8634 ( .A(n7769), .B(n6137), .Z(n3689) );
  XOR U8635 ( .A(n8975), .B(n8976), .Z(n6137) );
  XNOR U8636 ( .A(n4806), .B(n2005), .Z(n8976) );
  XOR U8637 ( .A(n8977), .B(n8978), .Z(n2005) );
  ANDN U8638 ( .B(n7960), .A(n7958), .Z(n8977) );
  XNOR U8639 ( .A(n8979), .B(n8980), .Z(n4806) );
  ANDN U8640 ( .B(n7968), .A(n7966), .Z(n8979) );
  XNOR U8641 ( .A(n6046), .B(n8981), .Z(n8975) );
  XOR U8642 ( .A(n5270), .B(n3843), .Z(n8981) );
  XNOR U8643 ( .A(n8982), .B(n8983), .Z(n3843) );
  NOR U8644 ( .A(n7954), .B(n7953), .Z(n8982) );
  XOR U8645 ( .A(n8984), .B(n8985), .Z(n5270) );
  ANDN U8646 ( .B(n7964), .A(n7962), .Z(n8984) );
  XNOR U8647 ( .A(n8986), .B(n8987), .Z(n6046) );
  AND U8648 ( .A(n7951), .B(n7949), .Z(n8986) );
  IV U8649 ( .A(n8988), .Z(n7949) );
  XOR U8650 ( .A(n8989), .B(n8990), .Z(n7769) );
  XNOR U8651 ( .A(n4967), .B(n8991), .Z(n8990) );
  XNOR U8652 ( .A(n8992), .B(n7858), .Z(n4967) );
  AND U8653 ( .A(n8993), .B(n8917), .Z(n8992) );
  XOR U8654 ( .A(n2288), .B(n8994), .Z(n8989) );
  XOR U8655 ( .A(n3376), .B(n6577), .Z(n8994) );
  XOR U8656 ( .A(n8995), .B(n7846), .Z(n6577) );
  IV U8657 ( .A(n8996), .Z(n7846) );
  ANDN U8658 ( .B(n8920), .A(n8997), .Z(n8995) );
  IV U8659 ( .A(n8998), .Z(n8920) );
  XOR U8660 ( .A(n8999), .B(n7851), .Z(n3376) );
  AND U8661 ( .A(n8915), .B(n9000), .Z(n8999) );
  XOR U8662 ( .A(n9001), .B(n7841), .Z(n2288) );
  AND U8663 ( .A(n8924), .B(n9002), .Z(n9001) );
  XNOR U8664 ( .A(n2535), .B(n9003), .Z(n1174) );
  IV U8665 ( .A(n4858), .Z(n2535) );
  XOR U8666 ( .A(n5876), .B(n6286), .Z(n4858) );
  XOR U8667 ( .A(n9004), .B(n9005), .Z(n6286) );
  XNOR U8668 ( .A(n3275), .B(n4977), .Z(n9005) );
  XOR U8669 ( .A(n9006), .B(n6538), .Z(n4977) );
  AND U8670 ( .A(n6539), .B(n9007), .Z(n9006) );
  XNOR U8671 ( .A(n9008), .B(n6543), .Z(n3275) );
  AND U8672 ( .A(n8961), .B(n9009), .Z(n9008) );
  IV U8673 ( .A(n9010), .Z(n8961) );
  XOR U8674 ( .A(n5282), .B(n9011), .Z(n9004) );
  XNOR U8675 ( .A(n6519), .B(n2570), .Z(n9011) );
  XOR U8676 ( .A(n9012), .B(n6529), .Z(n2570) );
  ANDN U8677 ( .B(n9013), .A(n9014), .Z(n9012) );
  XNOR U8678 ( .A(n9015), .B(n6535), .Z(n6519) );
  ANDN U8679 ( .B(n6534), .A(n8952), .Z(n9015) );
  IV U8680 ( .A(n9016), .Z(n6534) );
  XNOR U8681 ( .A(n9017), .B(n6526), .Z(n5282) );
  ANDN U8682 ( .B(n8964), .A(n6525), .Z(n9017) );
  XOR U8683 ( .A(n9018), .B(n9019), .Z(n5876) );
  XNOR U8684 ( .A(n3861), .B(n5150), .Z(n9019) );
  XNOR U8685 ( .A(n9020), .B(n7029), .Z(n5150) );
  NOR U8686 ( .A(n7028), .B(n6560), .Z(n9020) );
  XOR U8687 ( .A(n9021), .B(n9022), .Z(n3861) );
  ANDN U8688 ( .B(n9023), .A(n6564), .Z(n9021) );
  XOR U8689 ( .A(n4254), .B(n9024), .Z(n9018) );
  XNOR U8690 ( .A(n7007), .B(n1793), .Z(n9024) );
  XNOR U8691 ( .A(n9025), .B(n7026), .Z(n1793) );
  XOR U8692 ( .A(n9026), .B(n7036), .Z(n7007) );
  AND U8693 ( .A(n6555), .B(n7037), .Z(n9026) );
  XNOR U8694 ( .A(n9027), .B(n7033), .Z(n4254) );
  AND U8695 ( .A(n6551), .B(n7034), .Z(n9027) );
  XOR U8696 ( .A(n9028), .B(n6003), .Z(out[1032]) );
  XNOR U8697 ( .A(n8053), .B(n3222), .Z(n6003) );
  XNOR U8698 ( .A(n9029), .B(n9030), .Z(n3222) );
  XNOR U8699 ( .A(n9031), .B(n9032), .Z(n8053) );
  ANDN U8700 ( .B(n1178), .A(n1179), .Z(n9028) );
  XOR U8701 ( .A(n9035), .B(n1939), .Z(n1179) );
  XOR U8702 ( .A(n9036), .B(n9037), .Z(n7836) );
  XOR U8703 ( .A(n4970), .B(n9038), .Z(n9037) );
  XNOR U8704 ( .A(n9039), .B(n7967), .Z(n4970) );
  NOR U8705 ( .A(n8980), .B(n9040), .Z(n9039) );
  XOR U8706 ( .A(n2295), .B(n9041), .Z(n9036) );
  XOR U8707 ( .A(n3378), .B(n6857), .Z(n9041) );
  XOR U8708 ( .A(n9042), .B(n7955), .Z(n6857) );
  IV U8709 ( .A(n9043), .Z(n7955) );
  AND U8710 ( .A(n9044), .B(n8983), .Z(n9042) );
  XNOR U8711 ( .A(n9045), .B(n7959), .Z(n3378) );
  ANDN U8712 ( .B(n8978), .A(n9046), .Z(n9045) );
  XNOR U8713 ( .A(n9047), .B(n7950), .Z(n2295) );
  XNOR U8714 ( .A(n9049), .B(n9050), .Z(n6143) );
  XOR U8715 ( .A(n9051), .B(n3850), .Z(n9050) );
  XOR U8716 ( .A(n9052), .B(n9053), .Z(n3850) );
  AND U8717 ( .A(n8006), .B(n8004), .Z(n9052) );
  XOR U8718 ( .A(n4833), .B(n9054), .Z(n9049) );
  XNOR U8719 ( .A(n2008), .B(n5275), .Z(n9054) );
  XNOR U8720 ( .A(n9055), .B(n9056), .Z(n5275) );
  XNOR U8721 ( .A(n9057), .B(n9058), .Z(n2008) );
  XOR U8722 ( .A(n9059), .B(n9060), .Z(n4833) );
  XNOR U8723 ( .A(n4031), .B(n7030), .Z(n1178) );
  XNOR U8724 ( .A(n9061), .B(n6565), .Z(n7030) );
  ANDN U8725 ( .B(n9062), .A(n9022), .Z(n9061) );
  IV U8726 ( .A(n2544), .Z(n4031) );
  XOR U8727 ( .A(n6290), .B(n5881), .Z(n2544) );
  XOR U8728 ( .A(n9063), .B(n9064), .Z(n5881) );
  XOR U8729 ( .A(n3865), .B(n5152), .Z(n9064) );
  XOR U8730 ( .A(n9065), .B(n7089), .Z(n5152) );
  ANDN U8731 ( .B(n6593), .A(n7011), .Z(n9065) );
  XNOR U8732 ( .A(n9066), .B(n9067), .Z(n7011) );
  XOR U8733 ( .A(n9068), .B(n9069), .Z(n6593) );
  XOR U8734 ( .A(n9070), .B(n9071), .Z(n3865) );
  ANDN U8735 ( .B(n7021), .A(n6597), .Z(n9070) );
  XNOR U8736 ( .A(n9072), .B(n9073), .Z(n6597) );
  XOR U8737 ( .A(n4256), .B(n9074), .Z(n9063) );
  XNOR U8738 ( .A(n1796), .B(n7065), .Z(n9074) );
  XNOR U8739 ( .A(n9075), .B(n7083), .Z(n7065) );
  AND U8740 ( .A(n6588), .B(n7016), .Z(n9075) );
  XOR U8741 ( .A(n9076), .B(n9077), .Z(n7016) );
  XOR U8742 ( .A(n9078), .B(n9079), .Z(n6588) );
  XNOR U8743 ( .A(n9080), .B(n7085), .Z(n1796) );
  ANDN U8744 ( .B(n7019), .A(n6601), .Z(n9080) );
  XOR U8745 ( .A(n9081), .B(n9082), .Z(n6601) );
  XNOR U8746 ( .A(n9083), .B(n9084), .Z(n7019) );
  XOR U8747 ( .A(n9085), .B(n7092), .Z(n4256) );
  ANDN U8748 ( .B(n7013), .A(n6584), .Z(n9085) );
  XNOR U8749 ( .A(n9086), .B(n9087), .Z(n6584) );
  XNOR U8750 ( .A(n9088), .B(n9089), .Z(n7013) );
  XOR U8751 ( .A(n9090), .B(n9091), .Z(n6290) );
  XNOR U8752 ( .A(n3282), .B(n5079), .Z(n9091) );
  XOR U8753 ( .A(n9092), .B(n9093), .Z(n5079) );
  ANDN U8754 ( .B(n9022), .A(n6565), .Z(n9092) );
  XNOR U8755 ( .A(n9094), .B(n9095), .Z(n6565) );
  XOR U8756 ( .A(n9096), .B(n9097), .Z(n9022) );
  XOR U8757 ( .A(n9098), .B(n9099), .Z(n3282) );
  ANDN U8758 ( .B(n7026), .A(n6569), .Z(n9098) );
  XOR U8759 ( .A(n9100), .B(n9101), .Z(n6569) );
  XNOR U8760 ( .A(n9102), .B(n9103), .Z(n7026) );
  XNOR U8761 ( .A(n5287), .B(n9104), .Z(n9090) );
  XOR U8762 ( .A(n6546), .B(n2579), .Z(n9104) );
  XNOR U8763 ( .A(n9105), .B(n6557), .Z(n2579) );
  ANDN U8764 ( .B(n6556), .A(n7036), .Z(n9105) );
  XNOR U8765 ( .A(n9106), .B(n9107), .Z(n7036) );
  XNOR U8766 ( .A(n9108), .B(n9109), .Z(n6556) );
  XNOR U8767 ( .A(n9110), .B(n6562), .Z(n6546) );
  ANDN U8768 ( .B(n6561), .A(n7029), .Z(n9110) );
  XNOR U8769 ( .A(n9111), .B(n9112), .Z(n7029) );
  XNOR U8770 ( .A(n9113), .B(n9114), .Z(n6561) );
  XNOR U8771 ( .A(n9115), .B(n6553), .Z(n5287) );
  ANDN U8772 ( .B(n6552), .A(n7033), .Z(n9115) );
  XNOR U8773 ( .A(n9116), .B(n9117), .Z(n7033) );
  XOR U8774 ( .A(n9118), .B(n9119), .Z(n6552) );
  XOR U8775 ( .A(n9120), .B(n6013), .Z(out[1031]) );
  XOR U8776 ( .A(n8114), .B(n2471), .Z(n6013) );
  XNOR U8777 ( .A(n9121), .B(n9122), .Z(n2471) );
  XNOR U8778 ( .A(n9123), .B(n9124), .Z(n8114) );
  AND U8779 ( .A(n9125), .B(n9126), .Z(n9123) );
  ANDN U8780 ( .B(n1182), .A(n1183), .Z(n9120) );
  XOR U8781 ( .A(n9127), .B(n1943), .Z(n1183) );
  XOR U8782 ( .A(n9128), .B(n9129), .Z(n7945) );
  XNOR U8783 ( .A(n4973), .B(n9130), .Z(n9129) );
  XOR U8784 ( .A(n9131), .B(n8019), .Z(n4973) );
  NOR U8785 ( .A(n9132), .B(n9060), .Z(n9131) );
  XOR U8786 ( .A(n2306), .B(n9133), .Z(n9128) );
  XOR U8787 ( .A(n3380), .B(n7189), .Z(n9133) );
  XNOR U8788 ( .A(n9134), .B(n8005), .Z(n7189) );
  XOR U8789 ( .A(n9136), .B(n8010), .Z(n3380) );
  NOR U8790 ( .A(n9058), .B(n9137), .Z(n9136) );
  XOR U8791 ( .A(n9138), .B(n8001), .Z(n2306) );
  IV U8792 ( .A(n9139), .Z(n8001) );
  ANDN U8793 ( .B(n9140), .A(n9141), .Z(n9138) );
  XNOR U8794 ( .A(n9142), .B(n9143), .Z(n6148) );
  XNOR U8795 ( .A(n9144), .B(n3854), .Z(n9143) );
  XNOR U8796 ( .A(n9145), .B(n9146), .Z(n3854) );
  ANDN U8797 ( .B(n9147), .A(n7935), .Z(n9145) );
  XOR U8798 ( .A(n4871), .B(n9148), .Z(n9142) );
  XNOR U8799 ( .A(n2011), .B(n5280), .Z(n9148) );
  XOR U8800 ( .A(n9149), .B(n9150), .Z(n5280) );
  NOR U8801 ( .A(n7925), .B(n9151), .Z(n9149) );
  XNOR U8802 ( .A(n9152), .B(n9153), .Z(n2011) );
  AND U8803 ( .A(n8066), .B(n9154), .Z(n9152) );
  IV U8804 ( .A(n9155), .Z(n8066) );
  XOR U8805 ( .A(n9156), .B(n9157), .Z(n4871) );
  NOR U8806 ( .A(n9158), .B(n7929), .Z(n9156) );
  XNOR U8807 ( .A(n7087), .B(n4036), .Z(n1182) );
  IV U8808 ( .A(n2552), .Z(n4036) );
  XOR U8809 ( .A(n5886), .B(n6294), .Z(n2552) );
  XOR U8810 ( .A(n9159), .B(n9160), .Z(n6294) );
  XNOR U8811 ( .A(n3285), .B(n5462), .Z(n9160) );
  XOR U8812 ( .A(n9161), .B(n6599), .Z(n5462) );
  XNOR U8813 ( .A(n9162), .B(n9163), .Z(n6599) );
  ANDN U8814 ( .B(n9164), .A(n9071), .Z(n9161) );
  XNOR U8815 ( .A(n9165), .B(n6603), .Z(n3285) );
  XOR U8816 ( .A(n9166), .B(n9167), .Z(n6603) );
  AND U8817 ( .A(n7085), .B(n6602), .Z(n9165) );
  XOR U8818 ( .A(n9168), .B(n9169), .Z(n6602) );
  XNOR U8819 ( .A(n9170), .B(n9171), .Z(n7085) );
  XOR U8820 ( .A(n5291), .B(n9172), .Z(n9159) );
  XNOR U8821 ( .A(n6579), .B(n2584), .Z(n9172) );
  XNOR U8822 ( .A(n9173), .B(n7017), .Z(n2584) );
  IV U8823 ( .A(n6590), .Z(n7017) );
  XNOR U8824 ( .A(n9116), .B(n9174), .Z(n6590) );
  AND U8825 ( .A(n7083), .B(n7082), .Z(n9173) );
  XOR U8826 ( .A(n9175), .B(n9176), .Z(n7082) );
  XNOR U8827 ( .A(n9177), .B(n9178), .Z(n7083) );
  XOR U8828 ( .A(n9179), .B(n6595), .Z(n6579) );
  XOR U8829 ( .A(n9180), .B(n9181), .Z(n6595) );
  AND U8830 ( .A(n7089), .B(n6594), .Z(n9179) );
  XOR U8831 ( .A(n9182), .B(n9183), .Z(n6594) );
  XOR U8832 ( .A(n9184), .B(n9185), .Z(n7089) );
  XNOR U8833 ( .A(n9186), .B(n6585), .Z(n5291) );
  XNOR U8834 ( .A(n9187), .B(n9188), .Z(n6585) );
  ANDN U8835 ( .B(n7091), .A(n7092), .Z(n9186) );
  XNOR U8836 ( .A(n9189), .B(n9190), .Z(n7092) );
  XNOR U8837 ( .A(n9191), .B(n9192), .Z(n7091) );
  XOR U8838 ( .A(n9193), .B(n9194), .Z(n5886) );
  XNOR U8839 ( .A(n3870), .B(n5154), .Z(n9194) );
  XNOR U8840 ( .A(n9195), .B(n9196), .Z(n5154) );
  AND U8841 ( .A(n7074), .B(n6621), .Z(n9195) );
  XNOR U8842 ( .A(n9197), .B(n9198), .Z(n6621) );
  XOR U8843 ( .A(n9199), .B(n9200), .Z(n3870) );
  ANDN U8844 ( .B(n7071), .A(n6625), .Z(n9199) );
  XNOR U8845 ( .A(n9201), .B(n9202), .Z(n6625) );
  XOR U8846 ( .A(n9203), .B(n9204), .Z(n9193) );
  XNOR U8847 ( .A(n7121), .B(n1801), .Z(n9204) );
  XNOR U8848 ( .A(n9205), .B(n9206), .Z(n1801) );
  AND U8849 ( .A(n6629), .B(n9207), .Z(n9205) );
  XNOR U8850 ( .A(n9208), .B(n9209), .Z(n6629) );
  XOR U8851 ( .A(n9210), .B(n9211), .Z(n7121) );
  ANDN U8852 ( .B(n7078), .A(n6616), .Z(n9210) );
  XNOR U8853 ( .A(n9212), .B(n9213), .Z(n6616) );
  XOR U8854 ( .A(n9214), .B(n6598), .Z(n7087) );
  IV U8855 ( .A(n9164), .Z(n6598) );
  XOR U8856 ( .A(n9215), .B(n9216), .Z(n9164) );
  ANDN U8857 ( .B(n9071), .A(n7021), .Z(n9214) );
  XNOR U8858 ( .A(n9208), .B(n9217), .Z(n7021) );
  XOR U8859 ( .A(n9218), .B(n9219), .Z(n9071) );
  XNOR U8860 ( .A(n9220), .B(n6018), .Z(out[1030]) );
  XOR U8861 ( .A(n8140), .B(n2476), .Z(n6018) );
  XNOR U8862 ( .A(n9221), .B(n9222), .Z(n2476) );
  XNOR U8863 ( .A(n9223), .B(n9224), .Z(n8140) );
  ANDN U8864 ( .B(n1186), .A(n1188), .Z(n9220) );
  XNOR U8865 ( .A(n9227), .B(n1947), .Z(n1188) );
  XOR U8866 ( .A(n9228), .B(n9229), .Z(n7996) );
  XOR U8867 ( .A(n3383), .B(n4980), .Z(n9229) );
  XOR U8868 ( .A(n9230), .B(n7930), .Z(n4980) );
  AND U8869 ( .A(n9157), .B(n7931), .Z(n9230) );
  XNOR U8870 ( .A(n9231), .B(n8068), .Z(n3383) );
  ANDN U8871 ( .B(n8067), .A(n9153), .Z(n9231) );
  XNOR U8872 ( .A(n7920), .B(n9232), .Z(n9228) );
  XNOR U8873 ( .A(n7038), .B(n2314), .Z(n9232) );
  XNOR U8874 ( .A(n9233), .B(n7940), .Z(n2314) );
  AND U8875 ( .A(n9234), .B(n7941), .Z(n9233) );
  XOR U8876 ( .A(n9235), .B(n7926), .Z(n7038) );
  IV U8877 ( .A(n9236), .Z(n7926) );
  XOR U8878 ( .A(n9237), .B(n7936), .Z(n7920) );
  AND U8879 ( .A(n9146), .B(n7937), .Z(n9237) );
  XNOR U8880 ( .A(n9238), .B(n9239), .Z(n6153) );
  XOR U8881 ( .A(n9240), .B(n3857), .Z(n9239) );
  XOR U8882 ( .A(n9241), .B(n9242), .Z(n3857) );
  AND U8883 ( .A(n9243), .B(n8580), .Z(n9241) );
  IV U8884 ( .A(n9244), .Z(n8580) );
  XOR U8885 ( .A(n4905), .B(n9245), .Z(n9238) );
  XNOR U8886 ( .A(n2014), .B(n5286), .Z(n9245) );
  XNOR U8887 ( .A(n9246), .B(n9247), .Z(n5286) );
  AND U8888 ( .A(n9248), .B(n8571), .Z(n9246) );
  XNOR U8889 ( .A(n9249), .B(n9250), .Z(n2014) );
  ANDN U8890 ( .B(n9251), .A(n9252), .Z(n9249) );
  ANDN U8891 ( .B(n9255), .A(n8575), .Z(n9253) );
  XNOR U8892 ( .A(n9256), .B(n3484), .Z(n1186) );
  IV U8893 ( .A(n2559), .Z(n3484) );
  XNOR U8894 ( .A(n5892), .B(n6299), .Z(n2559) );
  XNOR U8895 ( .A(n9257), .B(n9258), .Z(n6299) );
  XNOR U8896 ( .A(n2593), .B(n5297), .Z(n9258) );
  XOR U8897 ( .A(n9259), .B(n6613), .Z(n5297) );
  XNOR U8898 ( .A(n9260), .B(n9261), .Z(n6613) );
  AND U8899 ( .A(n9262), .B(n9263), .Z(n9259) );
  XNOR U8900 ( .A(n9264), .B(n6617), .Z(n2593) );
  XNOR U8901 ( .A(n9265), .B(n9190), .Z(n6617) );
  ANDN U8902 ( .B(n9266), .A(n9211), .Z(n9264) );
  XNOR U8903 ( .A(n3288), .B(n9267), .Z(n9257) );
  XNOR U8904 ( .A(n5804), .B(n6607), .Z(n9267) );
  XNOR U8905 ( .A(n9268), .B(n6623), .Z(n6607) );
  XOR U8906 ( .A(n9269), .B(n9270), .Z(n6623) );
  AND U8907 ( .A(n9196), .B(n9271), .Z(n9268) );
  XNOR U8908 ( .A(n9272), .B(n6626), .Z(n5804) );
  XNOR U8909 ( .A(n9273), .B(n9274), .Z(n6626) );
  ANDN U8910 ( .B(n9275), .A(n9200), .Z(n9272) );
  XNOR U8911 ( .A(n9276), .B(n6631), .Z(n3288) );
  XNOR U8912 ( .A(n9277), .B(n9278), .Z(n6631) );
  AND U8913 ( .A(n6630), .B(n9206), .Z(n9276) );
  XOR U8914 ( .A(n9279), .B(n9280), .Z(n5892) );
  XOR U8915 ( .A(n3874), .B(n5156), .Z(n9280) );
  XNOR U8916 ( .A(n9281), .B(n7176), .Z(n5156) );
  AND U8917 ( .A(n6648), .B(n9282), .Z(n9281) );
  XNOR U8918 ( .A(n9283), .B(n9284), .Z(n3874) );
  AND U8919 ( .A(n6652), .B(n9285), .Z(n9283) );
  XOR U8920 ( .A(n4067), .B(n9286), .Z(n9279) );
  XOR U8921 ( .A(n7148), .B(n1805), .Z(n9286) );
  XNOR U8922 ( .A(n9287), .B(n7171), .Z(n1805) );
  AND U8923 ( .A(n7170), .B(n6656), .Z(n9287) );
  XNOR U8924 ( .A(n9288), .B(n7167), .Z(n7148) );
  AND U8925 ( .A(n6643), .B(n9289), .Z(n9288) );
  XNOR U8926 ( .A(n9290), .B(n7180), .Z(n4067) );
  NOR U8927 ( .A(n6639), .B(n7179), .Z(n9290) );
  XOR U8928 ( .A(n9291), .B(n4156), .Z(out[102]) );
  XOR U8929 ( .A(n6925), .B(n2555), .Z(n4156) );
  XNOR U8930 ( .A(n7883), .B(n9292), .Z(n2555) );
  XOR U8931 ( .A(n9293), .B(n9294), .Z(n7883) );
  XOR U8932 ( .A(n4331), .B(n2178), .Z(n9294) );
  XOR U8933 ( .A(n9295), .B(n9296), .Z(n2178) );
  AND U8934 ( .A(n9297), .B(n9298), .Z(n9295) );
  XNOR U8935 ( .A(n9299), .B(n9300), .Z(n4331) );
  ANDN U8936 ( .B(n6931), .A(n6932), .Z(n9299) );
  XOR U8937 ( .A(n5955), .B(n9301), .Z(n9293) );
  XNOR U8938 ( .A(n5503), .B(n3750), .Z(n9301) );
  XNOR U8939 ( .A(n9302), .B(n9303), .Z(n3750) );
  AND U8940 ( .A(n6923), .B(n6921), .Z(n9302) );
  XNOR U8941 ( .A(n9304), .B(n9305), .Z(n5503) );
  AND U8942 ( .A(n6927), .B(n9306), .Z(n9304) );
  XOR U8943 ( .A(n9307), .B(n9308), .Z(n5955) );
  ANDN U8944 ( .B(n6917), .A(n6919), .Z(n9307) );
  XOR U8945 ( .A(n9309), .B(n9297), .Z(n6925) );
  ANDN U8946 ( .B(n9310), .A(n9298), .Z(n9309) );
  AND U8947 ( .A(n3539), .B(n4327), .Z(n9291) );
  XNOR U8948 ( .A(n7381), .B(n2397), .Z(n4327) );
  XNOR U8949 ( .A(n9311), .B(n9312), .Z(n2397) );
  XOR U8950 ( .A(n9313), .B(n9314), .Z(n7381) );
  ANDN U8951 ( .B(n9315), .A(n9316), .Z(n9313) );
  XNOR U8952 ( .A(n2329), .B(n9317), .Z(n3539) );
  XOR U8953 ( .A(n6152), .B(n9318), .Z(n2329) );
  XOR U8954 ( .A(n9319), .B(n9320), .Z(n6152) );
  XNOR U8955 ( .A(n3176), .B(n6856), .Z(n9320) );
  XOR U8956 ( .A(n9321), .B(n9322), .Z(n6856) );
  NOR U8957 ( .A(n9323), .B(n9324), .Z(n9321) );
  XOR U8958 ( .A(n9325), .B(n9326), .Z(n3176) );
  NOR U8959 ( .A(n9327), .B(n9328), .Z(n9325) );
  XOR U8960 ( .A(n5459), .B(n9329), .Z(n9319) );
  XOR U8961 ( .A(n8178), .B(n2362), .Z(n9329) );
  XOR U8962 ( .A(n9330), .B(n9331), .Z(n2362) );
  AND U8963 ( .A(n9332), .B(n9333), .Z(n9330) );
  XOR U8964 ( .A(n9334), .B(n9335), .Z(n8178) );
  ANDN U8965 ( .B(n9336), .A(n9337), .Z(n9334) );
  XOR U8966 ( .A(n9338), .B(n9339), .Z(n5459) );
  NOR U8967 ( .A(n9340), .B(n9341), .Z(n9338) );
  XOR U8968 ( .A(n9342), .B(n6023), .Z(out[1029]) );
  XOR U8969 ( .A(n8194), .B(n2483), .Z(n6023) );
  XNOR U8970 ( .A(n9343), .B(n9344), .Z(n2483) );
  XNOR U8971 ( .A(n9345), .B(n9346), .Z(n8194) );
  NOR U8972 ( .A(n9347), .B(n9348), .Z(n9345) );
  ANDN U8973 ( .B(n1192), .A(n1190), .Z(n9342) );
  XOR U8974 ( .A(n7173), .B(n3487), .Z(n1190) );
  IV U8975 ( .A(n2564), .Z(n3487) );
  XNOR U8976 ( .A(n5901), .B(n6303), .Z(n2564) );
  XNOR U8977 ( .A(n9349), .B(n9350), .Z(n6303) );
  XNOR U8978 ( .A(n2602), .B(n5302), .Z(n9350) );
  XOR U8979 ( .A(n9351), .B(n6641), .Z(n5302) );
  AND U8980 ( .A(n7180), .B(n7178), .Z(n9351) );
  IV U8981 ( .A(n6640), .Z(n7178) );
  XNOR U8982 ( .A(n9352), .B(n9353), .Z(n6640) );
  XOR U8983 ( .A(n9354), .B(n9355), .Z(n7180) );
  XNOR U8984 ( .A(n9356), .B(n6644), .Z(n2602) );
  AND U8985 ( .A(n6645), .B(n7167), .Z(n9356) );
  XNOR U8986 ( .A(n9357), .B(n9358), .Z(n7167) );
  XNOR U8987 ( .A(n9359), .B(n9360), .Z(n6645) );
  XOR U8988 ( .A(n3291), .B(n9361), .Z(n9349) );
  XNOR U8989 ( .A(n6305), .B(n6634), .Z(n9361) );
  XOR U8990 ( .A(n9362), .B(n6649), .Z(n6634) );
  AND U8991 ( .A(n6650), .B(n7176), .Z(n9362) );
  XNOR U8992 ( .A(n9363), .B(n9364), .Z(n7176) );
  XNOR U8993 ( .A(n9365), .B(n9366), .Z(n6650) );
  XNOR U8994 ( .A(n9367), .B(n6653), .Z(n6305) );
  AND U8995 ( .A(n9284), .B(n6654), .Z(n9367) );
  XNOR U8996 ( .A(n9368), .B(n6657), .Z(n3291) );
  AND U8997 ( .A(n7171), .B(n7169), .Z(n9368) );
  XNOR U8998 ( .A(n9369), .B(n9370), .Z(n7169) );
  XNOR U8999 ( .A(n9371), .B(n9372), .Z(n7171) );
  XOR U9000 ( .A(n9373), .B(n9374), .Z(n5901) );
  XOR U9001 ( .A(n3553), .B(n5159), .Z(n9374) );
  XNOR U9002 ( .A(n9375), .B(n7243), .Z(n5159) );
  AND U9003 ( .A(n7158), .B(n6681), .Z(n9375) );
  XOR U9004 ( .A(n9376), .B(n9377), .Z(n6681) );
  XNOR U9005 ( .A(n9378), .B(n9379), .Z(n7158) );
  XNOR U9006 ( .A(n9380), .B(n9381), .Z(n3553) );
  AND U9007 ( .A(n6666), .B(n9382), .Z(n9380) );
  XNOR U9008 ( .A(n9383), .B(n9384), .Z(n6666) );
  XOR U9009 ( .A(n4070), .B(n9385), .Z(n9373) );
  XOR U9010 ( .A(n7218), .B(n1809), .Z(n9385) );
  XOR U9011 ( .A(n9386), .B(n7239), .Z(n1809) );
  AND U9012 ( .A(n7152), .B(n6670), .Z(n9386) );
  IV U9013 ( .A(n7153), .Z(n6670) );
  XNOR U9014 ( .A(n9387), .B(n9388), .Z(n7153) );
  XOR U9015 ( .A(n9389), .B(n9390), .Z(n7152) );
  XNOR U9016 ( .A(n9391), .B(n7237), .Z(n7218) );
  ANDN U9017 ( .B(n7162), .A(n6674), .Z(n9391) );
  XNOR U9018 ( .A(n9392), .B(n9191), .Z(n6674) );
  XNOR U9019 ( .A(n9393), .B(n9394), .Z(n7162) );
  XOR U9020 ( .A(n9395), .B(n7245), .Z(n4070) );
  IV U9021 ( .A(n9396), .Z(n7245) );
  ANDN U9022 ( .B(n7155), .A(n6685), .Z(n9395) );
  XNOR U9023 ( .A(n9397), .B(n9398), .Z(n6685) );
  XOR U9024 ( .A(n9399), .B(n9400), .Z(n7155) );
  XNOR U9025 ( .A(n9401), .B(n6654), .Z(n7173) );
  XOR U9026 ( .A(n9402), .B(n9403), .Z(n6654) );
  ANDN U9027 ( .B(n9404), .A(n9284), .Z(n9401) );
  XOR U9028 ( .A(n9405), .B(n9406), .Z(n9284) );
  XOR U9029 ( .A(n9407), .B(n4175), .Z(n1192) );
  IV U9030 ( .A(n1953), .Z(n4175) );
  XOR U9031 ( .A(n9408), .B(n9409), .Z(n8063) );
  XNOR U9032 ( .A(n3386), .B(n4984), .Z(n9409) );
  XNOR U9033 ( .A(n9410), .B(n8576), .Z(n4984) );
  AND U9034 ( .A(n8577), .B(n9254), .Z(n9410) );
  XNOR U9035 ( .A(n9411), .B(n8586), .Z(n3386) );
  AND U9036 ( .A(n8585), .B(n9250), .Z(n9411) );
  XNOR U9037 ( .A(n8566), .B(n9412), .Z(n9408) );
  XOR U9038 ( .A(n7093), .B(n2321), .Z(n9412) );
  XOR U9039 ( .A(n9413), .B(n8589), .Z(n2321) );
  ANDN U9040 ( .B(n9414), .A(n8590), .Z(n9413) );
  XOR U9041 ( .A(n9415), .B(n8573), .Z(n7093) );
  ANDN U9042 ( .B(n9416), .A(n9247), .Z(n9415) );
  XNOR U9043 ( .A(n9417), .B(n8582), .Z(n8566) );
  ANDN U9044 ( .B(n9418), .A(n9242), .Z(n9417) );
  XNOR U9045 ( .A(n9419), .B(n9420), .Z(n6158) );
  XNOR U9046 ( .A(n9421), .B(n3863), .Z(n9420) );
  XOR U9047 ( .A(n9422), .B(n9423), .Z(n3863) );
  AND U9048 ( .A(n9424), .B(n9331), .Z(n9422) );
  IV U9049 ( .A(n9425), .Z(n9331) );
  XNOR U9050 ( .A(n4942), .B(n9426), .Z(n9419) );
  XNOR U9051 ( .A(n2017), .B(n5290), .Z(n9426) );
  XNOR U9052 ( .A(n9427), .B(n9428), .Z(n5290) );
  AND U9053 ( .A(n9322), .B(n9429), .Z(n9427) );
  XNOR U9054 ( .A(n9430), .B(n9431), .Z(n2017) );
  AND U9055 ( .A(n9432), .B(n9335), .Z(n9430) );
  IV U9056 ( .A(n9433), .Z(n9335) );
  XNOR U9057 ( .A(n9434), .B(n9435), .Z(n4942) );
  AND U9058 ( .A(n9326), .B(n9436), .Z(n9434) );
  IV U9059 ( .A(n9437), .Z(n9326) );
  XOR U9060 ( .A(n9438), .B(n6028), .Z(out[1028]) );
  XOR U9061 ( .A(n8278), .B(n2490), .Z(n6028) );
  XNOR U9062 ( .A(n9439), .B(n9440), .Z(n2490) );
  XNOR U9063 ( .A(n9441), .B(n9442), .Z(n8278) );
  ANDN U9064 ( .B(n9443), .A(n9444), .Z(n9441) );
  ANDN U9065 ( .B(n1194), .A(n1195), .Z(n9438) );
  XOR U9066 ( .A(n9445), .B(n1961), .Z(n1195) );
  XOR U9067 ( .A(n9446), .B(n9447), .Z(n8125) );
  XOR U9068 ( .A(n3393), .B(n4988), .Z(n9447) );
  XNOR U9069 ( .A(n9448), .B(n9328), .Z(n4988) );
  AND U9070 ( .A(n9327), .B(n9435), .Z(n9448) );
  XNOR U9071 ( .A(n9449), .B(n9337), .Z(n3393) );
  AND U9072 ( .A(n9431), .B(n9450), .Z(n9449) );
  XOR U9073 ( .A(n9317), .B(n9451), .Z(n9446) );
  XNOR U9074 ( .A(n7120), .B(n2330), .Z(n9451) );
  XNOR U9075 ( .A(n9452), .B(n9340), .Z(n2330) );
  ANDN U9076 ( .B(n9341), .A(n9453), .Z(n9452) );
  XOR U9077 ( .A(n9454), .B(n9324), .Z(n7120) );
  ANDN U9078 ( .B(n9323), .A(n9428), .Z(n9454) );
  XOR U9079 ( .A(n9455), .B(n9332), .Z(n9317) );
  ANDN U9080 ( .B(n9456), .A(n9423), .Z(n9455) );
  XNOR U9081 ( .A(n9457), .B(n9458), .Z(n6163) );
  XNOR U9082 ( .A(n2020), .B(n3867), .Z(n9458) );
  XOR U9083 ( .A(n9459), .B(n9460), .Z(n3867) );
  AND U9084 ( .A(n9461), .B(n9462), .Z(n9459) );
  XOR U9085 ( .A(n9463), .B(n9464), .Z(n2020) );
  ANDN U9086 ( .B(n9465), .A(n9466), .Z(n9463) );
  XNOR U9087 ( .A(n9467), .B(n9468), .Z(n9457) );
  XNOR U9088 ( .A(n5295), .B(n4976), .Z(n9468) );
  XNOR U9089 ( .A(n9469), .B(n9470), .Z(n4976) );
  XNOR U9090 ( .A(n9473), .B(n9474), .Z(n5295) );
  NOR U9091 ( .A(n9475), .B(n9476), .Z(n9473) );
  XNOR U9092 ( .A(n7241), .B(n2573), .Z(n1194) );
  XNOR U9093 ( .A(n5906), .B(n6316), .Z(n2573) );
  XNOR U9094 ( .A(n9477), .B(n9478), .Z(n6316) );
  XOR U9095 ( .A(n2612), .B(n5307), .Z(n9478) );
  XOR U9096 ( .A(n9479), .B(n6687), .Z(n5307) );
  XOR U9097 ( .A(n9480), .B(n9481), .Z(n6687) );
  AND U9098 ( .A(n6686), .B(n9396), .Z(n9479) );
  XNOR U9099 ( .A(n9482), .B(n9483), .Z(n9396) );
  XNOR U9100 ( .A(n9484), .B(n9485), .Z(n6686) );
  XOR U9101 ( .A(n9486), .B(n6679), .Z(n2612) );
  XOR U9102 ( .A(n9354), .B(n9487), .Z(n6679) );
  AND U9103 ( .A(n7237), .B(n6678), .Z(n9486) );
  IV U9104 ( .A(n7236), .Z(n6678) );
  XOR U9105 ( .A(n9488), .B(n9489), .Z(n7236) );
  XOR U9106 ( .A(n9101), .B(n9490), .Z(n7237) );
  XOR U9107 ( .A(n6661), .B(n9491), .Z(n9477) );
  XOR U9108 ( .A(n5139), .B(n3294), .Z(n9491) );
  XNOR U9109 ( .A(n9492), .B(n6671), .Z(n3294) );
  XNOR U9110 ( .A(n9493), .B(n9494), .Z(n6671) );
  ANDN U9111 ( .B(n6672), .A(n7239), .Z(n9492) );
  XNOR U9112 ( .A(n9495), .B(n9496), .Z(n7239) );
  XNOR U9113 ( .A(n9497), .B(n9086), .Z(n6672) );
  XOR U9114 ( .A(n9499), .B(n9500), .Z(n6667) );
  AND U9115 ( .A(n6668), .B(n9381), .Z(n9498) );
  XNOR U9116 ( .A(n9501), .B(n6682), .Z(n6661) );
  XOR U9117 ( .A(n9502), .B(n9503), .Z(n6682) );
  AND U9118 ( .A(n6683), .B(n7243), .Z(n9501) );
  XOR U9119 ( .A(n9504), .B(n9505), .Z(n7243) );
  XNOR U9120 ( .A(n9506), .B(n9507), .Z(n6683) );
  XOR U9121 ( .A(n9508), .B(n9509), .Z(n5906) );
  XNOR U9122 ( .A(n1821), .B(n5162), .Z(n9509) );
  XOR U9123 ( .A(n9510), .B(n7297), .Z(n5162) );
  AND U9124 ( .A(n7228), .B(n6703), .Z(n9510) );
  XOR U9125 ( .A(n9511), .B(n9512), .Z(n6703) );
  XNOR U9126 ( .A(n9513), .B(n9514), .Z(n7228) );
  XNOR U9127 ( .A(n9515), .B(n7293), .Z(n1821) );
  ANDN U9128 ( .B(n6711), .A(n7222), .Z(n9515) );
  XNOR U9129 ( .A(n9516), .B(n9517), .Z(n7222) );
  XNOR U9130 ( .A(n9518), .B(n9519), .Z(n6711) );
  XNOR U9131 ( .A(n4073), .B(n9520), .Z(n9508) );
  XOR U9132 ( .A(n7272), .B(n3557), .Z(n9520) );
  XNOR U9133 ( .A(n9521), .B(n9522), .Z(n3557) );
  ANDN U9134 ( .B(n7230), .A(n6707), .Z(n9521) );
  XNOR U9135 ( .A(n9523), .B(n9524), .Z(n6707) );
  XNOR U9136 ( .A(n9525), .B(n7291), .Z(n7272) );
  AND U9137 ( .A(n6698), .B(n7232), .Z(n9525) );
  XNOR U9138 ( .A(n9526), .B(n9527), .Z(n7232) );
  XOR U9139 ( .A(n9528), .B(n9529), .Z(n6698) );
  XOR U9140 ( .A(n9530), .B(n7299), .Z(n4073) );
  ANDN U9141 ( .B(n6694), .A(n7224), .Z(n9530) );
  XNOR U9142 ( .A(n9383), .B(n9531), .Z(n7224) );
  XOR U9143 ( .A(n9532), .B(n9533), .Z(n6694) );
  XNOR U9144 ( .A(n9534), .B(n6668), .Z(n7241) );
  XNOR U9145 ( .A(n9535), .B(n9536), .Z(n6668) );
  ANDN U9146 ( .B(n7160), .A(n9381), .Z(n9534) );
  XNOR U9147 ( .A(n9537), .B(n9538), .Z(n9381) );
  IV U9148 ( .A(n9382), .Z(n7160) );
  XOR U9149 ( .A(n9539), .B(n9519), .Z(n9382) );
  XOR U9150 ( .A(n9540), .B(n6033), .Z(out[1027]) );
  XNOR U9151 ( .A(n8330), .B(n4676), .Z(n6033) );
  IV U9152 ( .A(n2499), .Z(n4676) );
  XNOR U9153 ( .A(n9541), .B(n9542), .Z(n2499) );
  XOR U9154 ( .A(n9543), .B(n9544), .Z(n8330) );
  ANDN U9155 ( .B(n9545), .A(n9546), .Z(n9543) );
  AND U9156 ( .A(n1200), .B(n1198), .Z(n9540) );
  IV U9157 ( .A(n6341), .Z(n1198) );
  XNOR U9158 ( .A(n7295), .B(n2578), .Z(n6341) );
  XNOR U9159 ( .A(n5911), .B(n6320), .Z(n2578) );
  XNOR U9160 ( .A(n9547), .B(n9548), .Z(n6320) );
  XNOR U9161 ( .A(n2618), .B(n5311), .Z(n9548) );
  XOR U9162 ( .A(n9549), .B(n7225), .Z(n5311) );
  IV U9163 ( .A(n6695), .Z(n7225) );
  XNOR U9164 ( .A(n9550), .B(n9551), .Z(n6695) );
  ANDN U9165 ( .B(n6696), .A(n7299), .Z(n9549) );
  XNOR U9166 ( .A(n9552), .B(n9553), .Z(n7299) );
  XNOR U9167 ( .A(n9554), .B(n9555), .Z(n6696) );
  XNOR U9168 ( .A(n9556), .B(n6700), .Z(n2618) );
  XNOR U9169 ( .A(n9557), .B(n9483), .Z(n6700) );
  AND U9170 ( .A(n7291), .B(n7290), .Z(n9556) );
  XNOR U9171 ( .A(n9558), .B(n9559), .Z(n7290) );
  XNOR U9172 ( .A(n9168), .B(n9560), .Z(n7291) );
  XOR U9173 ( .A(n3297), .B(n9561), .Z(n9547) );
  XNOR U9174 ( .A(n5168), .B(n6689), .Z(n9561) );
  XNOR U9175 ( .A(n9562), .B(n6704), .Z(n6689) );
  XOR U9176 ( .A(n9097), .B(n9563), .Z(n6704) );
  ANDN U9177 ( .B(n6705), .A(n7297), .Z(n9562) );
  XNOR U9178 ( .A(n9564), .B(n9565), .Z(n7297) );
  XOR U9179 ( .A(n9566), .B(n9567), .Z(n6705) );
  XNOR U9180 ( .A(n9568), .B(n6709), .Z(n5168) );
  XNOR U9181 ( .A(n9378), .B(n9569), .Z(n6709) );
  AND U9182 ( .A(n9522), .B(n9570), .Z(n9568) );
  XNOR U9183 ( .A(n9571), .B(n6712), .Z(n3297) );
  XNOR U9184 ( .A(n9572), .B(n9573), .Z(n6712) );
  AND U9185 ( .A(n6713), .B(n7293), .Z(n9571) );
  XNOR U9186 ( .A(n9574), .B(n9575), .Z(n7293) );
  XNOR U9187 ( .A(n9576), .B(n9577), .Z(n6713) );
  XOR U9188 ( .A(n9578), .B(n9579), .Z(n5911) );
  XNOR U9189 ( .A(n1825), .B(n5165), .Z(n9579) );
  XOR U9190 ( .A(n9580), .B(n7373), .Z(n5165) );
  ANDN U9191 ( .B(n7282), .A(n6729), .Z(n9580) );
  XNOR U9192 ( .A(n9581), .B(n9582), .Z(n6729) );
  XOR U9193 ( .A(n9583), .B(n9584), .Z(n7282) );
  XNOR U9194 ( .A(n9585), .B(n7368), .Z(n1825) );
  AND U9195 ( .A(n6737), .B(n7369), .Z(n9585) );
  XNOR U9196 ( .A(n9586), .B(n9587), .Z(n7369) );
  XNOR U9197 ( .A(n9588), .B(n9589), .Z(n6737) );
  XNOR U9198 ( .A(n4076), .B(n9590), .Z(n9578) );
  XNOR U9199 ( .A(n7345), .B(n3562), .Z(n9590) );
  XNOR U9200 ( .A(n9591), .B(n9592), .Z(n3562) );
  AND U9201 ( .A(n6733), .B(n9593), .Z(n9591) );
  XNOR U9202 ( .A(n9594), .B(n9595), .Z(n6733) );
  XNOR U9203 ( .A(n9596), .B(n7366), .Z(n7345) );
  ANDN U9204 ( .B(n6724), .A(n7286), .Z(n9596) );
  XNOR U9205 ( .A(n9597), .B(n9598), .Z(n7286) );
  XNOR U9206 ( .A(n9599), .B(n9353), .Z(n6724) );
  XNOR U9207 ( .A(n9600), .B(n7376), .Z(n4076) );
  ANDN U9208 ( .B(n7279), .A(n6720), .Z(n9600) );
  XNOR U9209 ( .A(n9601), .B(n9602), .Z(n6720) );
  XNOR U9210 ( .A(n9603), .B(n9524), .Z(n7279) );
  XOR U9211 ( .A(n9604), .B(n6708), .Z(n7295) );
  IV U9212 ( .A(n9570), .Z(n6708) );
  XNOR U9213 ( .A(n9605), .B(n9606), .Z(n9570) );
  NOR U9214 ( .A(n7230), .B(n9522), .Z(n9604) );
  XNOR U9215 ( .A(n9607), .B(n9608), .Z(n9522) );
  XOR U9216 ( .A(n9609), .B(n9588), .Z(n7230) );
  XOR U9217 ( .A(n9610), .B(n4181), .Z(n1200) );
  IV U9218 ( .A(n1965), .Z(n4181) );
  XOR U9219 ( .A(n9611), .B(n9612), .Z(n8179) );
  XOR U9220 ( .A(n3396), .B(n4991), .Z(n9612) );
  XNOR U9221 ( .A(n9613), .B(n9614), .Z(n4991) );
  ANDN U9222 ( .B(n9470), .A(n9615), .Z(n9613) );
  XOR U9223 ( .A(n9616), .B(n9617), .Z(n3396) );
  ANDN U9224 ( .B(n9618), .A(n9464), .Z(n9616) );
  XNOR U9225 ( .A(n9619), .B(n9620), .Z(n9611) );
  XOR U9226 ( .A(n7181), .B(n2337), .Z(n9620) );
  XOR U9227 ( .A(n9621), .B(n9622), .Z(n2337) );
  ANDN U9228 ( .B(n9623), .A(n9624), .Z(n9621) );
  XOR U9229 ( .A(n9625), .B(n9626), .Z(n7181) );
  AND U9230 ( .A(n9474), .B(n9627), .Z(n9625) );
  XNOR U9231 ( .A(n9628), .B(n9629), .Z(n6172) );
  XNOR U9232 ( .A(n2023), .B(n3871), .Z(n9629) );
  XOR U9233 ( .A(n9630), .B(n9631), .Z(n3871) );
  AND U9234 ( .A(n9632), .B(n9633), .Z(n9630) );
  XNOR U9235 ( .A(n9634), .B(n9635), .Z(n2023) );
  AND U9236 ( .A(n9636), .B(n9637), .Z(n9634) );
  XNOR U9237 ( .A(n9638), .B(n9639), .Z(n9628) );
  XNOR U9238 ( .A(n5300), .B(n5014), .Z(n9639) );
  XOR U9239 ( .A(n9640), .B(n9641), .Z(n5014) );
  ANDN U9240 ( .B(n9642), .A(n9643), .Z(n9640) );
  XNOR U9241 ( .A(n9644), .B(n9645), .Z(n5300) );
  AND U9242 ( .A(n9646), .B(n9647), .Z(n9644) );
  XOR U9243 ( .A(n9648), .B(n6344), .Z(out[1026]) );
  XOR U9244 ( .A(n8357), .B(n4701), .Z(n6344) );
  IV U9245 ( .A(n2506), .Z(n4701) );
  XNOR U9246 ( .A(n9649), .B(n9650), .Z(n2506) );
  XOR U9247 ( .A(n9651), .B(n9652), .Z(n8357) );
  ANDN U9248 ( .B(n9653), .A(n9654), .Z(n9651) );
  ANDN U9249 ( .B(n1204), .A(n1202), .Z(n9648) );
  XOR U9250 ( .A(n7371), .B(n3496), .Z(n1202) );
  IV U9251 ( .A(n2587), .Z(n3496) );
  XNOR U9252 ( .A(n5916), .B(n6324), .Z(n2587) );
  XNOR U9253 ( .A(n9655), .B(n9656), .Z(n6324) );
  XOR U9254 ( .A(n2625), .B(n5320), .Z(n9656) );
  XOR U9255 ( .A(n9657), .B(n6721), .Z(n5320) );
  XNOR U9256 ( .A(n9658), .B(n9659), .Z(n6721) );
  AND U9257 ( .A(n7376), .B(n7375), .Z(n9657) );
  XOR U9258 ( .A(n9660), .B(n9661), .Z(n7375) );
  XNOR U9259 ( .A(n9662), .B(n9663), .Z(n7376) );
  XNOR U9260 ( .A(n9664), .B(n6725), .Z(n2625) );
  XNOR U9261 ( .A(n9665), .B(n9666), .Z(n6725) );
  AND U9262 ( .A(n7366), .B(n7365), .Z(n9664) );
  XOR U9263 ( .A(n9667), .B(n9668), .Z(n7365) );
  XNOR U9264 ( .A(n9669), .B(n9670), .Z(n7366) );
  XOR U9265 ( .A(n3301), .B(n9671), .Z(n9655) );
  XOR U9266 ( .A(n5197), .B(n6715), .Z(n9671) );
  XNOR U9267 ( .A(n9672), .B(n6730), .Z(n6715) );
  XOR U9268 ( .A(n9673), .B(n9674), .Z(n6730) );
  ANDN U9269 ( .B(n6731), .A(n7373), .Z(n9672) );
  XNOR U9270 ( .A(n9675), .B(n9676), .Z(n7373) );
  XOR U9271 ( .A(n9677), .B(n9678), .Z(n6731) );
  XOR U9272 ( .A(n9679), .B(n7277), .Z(n5197) );
  XNOR U9273 ( .A(n9513), .B(n9680), .Z(n7277) );
  AND U9274 ( .A(n9592), .B(n6735), .Z(n9679) );
  XNOR U9275 ( .A(n9681), .B(n6738), .Z(n3301) );
  XNOR U9276 ( .A(n9682), .B(n9683), .Z(n6738) );
  AND U9277 ( .A(n6739), .B(n7368), .Z(n9681) );
  XNOR U9278 ( .A(n9684), .B(n9685), .Z(n7368) );
  XOR U9279 ( .A(n9686), .B(n9687), .Z(n6739) );
  XOR U9280 ( .A(n9688), .B(n9689), .Z(n5916) );
  XOR U9281 ( .A(n1829), .B(n5172), .Z(n9689) );
  XNOR U9282 ( .A(n9690), .B(n7467), .Z(n5172) );
  AND U9283 ( .A(n7356), .B(n6755), .Z(n9690) );
  XOR U9284 ( .A(n9691), .B(n9692), .Z(n6755) );
  XOR U9285 ( .A(n9693), .B(n9694), .Z(n7356) );
  XOR U9286 ( .A(n9695), .B(n7461), .Z(n1829) );
  AND U9287 ( .A(n6763), .B(n7462), .Z(n9695) );
  XNOR U9288 ( .A(n9696), .B(n9697), .Z(n7462) );
  XOR U9289 ( .A(n9698), .B(n9699), .Z(n6763) );
  XNOR U9290 ( .A(n4080), .B(n9700), .Z(n9688) );
  XNOR U9291 ( .A(n7441), .B(n3568), .Z(n9700) );
  XOR U9292 ( .A(n9701), .B(n9702), .Z(n3568) );
  ANDN U9293 ( .B(n7349), .A(n6759), .Z(n9701) );
  XOR U9294 ( .A(n9703), .B(n9704), .Z(n6759) );
  XOR U9295 ( .A(n9705), .B(n7459), .Z(n7441) );
  IV U9296 ( .A(n9706), .Z(n7459) );
  ANDN U9297 ( .B(n7361), .A(n6750), .Z(n9705) );
  XNOR U9298 ( .A(n9485), .B(n9707), .Z(n6750) );
  XNOR U9299 ( .A(n9187), .B(n9708), .Z(n7361) );
  XNOR U9300 ( .A(n9709), .B(n7469), .Z(n4080) );
  AND U9301 ( .A(n7351), .B(n7353), .Z(n9709) );
  XOR U9302 ( .A(n9710), .B(n9711), .Z(n7353) );
  XNOR U9303 ( .A(n9712), .B(n9713), .Z(n7351) );
  XNOR U9304 ( .A(n9714), .B(n6735), .Z(n7371) );
  XOR U9305 ( .A(n9715), .B(n9716), .Z(n6735) );
  ANDN U9306 ( .B(n7276), .A(n9592), .Z(n9714) );
  XOR U9307 ( .A(n9717), .B(n9718), .Z(n9592) );
  IV U9308 ( .A(n9593), .Z(n7276) );
  XOR U9309 ( .A(n9719), .B(n9720), .Z(n9593) );
  XOR U9310 ( .A(n9721), .B(n4185), .Z(n1204) );
  IV U9311 ( .A(n1660), .Z(n4185) );
  XOR U9312 ( .A(n9722), .B(n9723), .Z(n8233) );
  XNOR U9313 ( .A(n3399), .B(n4994), .Z(n9723) );
  XNOR U9314 ( .A(n9724), .B(n9725), .Z(n4994) );
  ANDN U9315 ( .B(n9726), .A(n9641), .Z(n9724) );
  XNOR U9316 ( .A(n9727), .B(n9728), .Z(n3399) );
  AND U9317 ( .A(n9635), .B(n9729), .Z(n9727) );
  XOR U9318 ( .A(n9730), .B(n9731), .Z(n9722) );
  XOR U9319 ( .A(n7217), .B(n2342), .Z(n9731) );
  XNOR U9320 ( .A(n9732), .B(n9733), .Z(n2342) );
  AND U9321 ( .A(n9734), .B(n9735), .Z(n9732) );
  XNOR U9322 ( .A(n9736), .B(n9737), .Z(n7217) );
  ANDN U9323 ( .B(n9738), .A(n9645), .Z(n9736) );
  XNOR U9324 ( .A(n9739), .B(n9740), .Z(n6177) );
  XNOR U9325 ( .A(n2030), .B(n3876), .Z(n9740) );
  XOR U9326 ( .A(n9741), .B(n9742), .Z(n3876) );
  NOR U9327 ( .A(n7312), .B(n9743), .Z(n9741) );
  XNOR U9328 ( .A(n9744), .B(n9745), .Z(n2030) );
  XOR U9329 ( .A(n9747), .B(n9748), .Z(n9739) );
  XNOR U9330 ( .A(n5305), .B(n5050), .Z(n9748) );
  XNOR U9331 ( .A(n9749), .B(n9750), .Z(n5050) );
  ANDN U9332 ( .B(n7306), .A(n9751), .Z(n9749) );
  XOR U9333 ( .A(n9752), .B(n9753), .Z(n5305) );
  NOR U9334 ( .A(n9754), .B(n8563), .Z(n9752) );
  XNOR U9335 ( .A(n9755), .B(n6044), .Z(out[1025]) );
  XNOR U9336 ( .A(n8411), .B(n4728), .Z(n6044) );
  IV U9337 ( .A(n2513), .Z(n4728) );
  XNOR U9338 ( .A(n9756), .B(n9757), .Z(n2513) );
  XNOR U9339 ( .A(n9758), .B(n9759), .Z(n8411) );
  ANDN U9340 ( .B(n9760), .A(n9761), .Z(n9758) );
  AND U9341 ( .A(n1207), .B(n1206), .Z(n9755) );
  IV U9342 ( .A(n6353), .Z(n1206) );
  XOR U9343 ( .A(n7464), .B(n2592), .Z(n6353) );
  XNOR U9344 ( .A(n5921), .B(n6328), .Z(n2592) );
  XNOR U9345 ( .A(n9762), .B(n9763), .Z(n6328) );
  XOR U9346 ( .A(n2632), .B(n5324), .Z(n9763) );
  XOR U9347 ( .A(n9764), .B(n7352), .Z(n5324) );
  IV U9348 ( .A(n6748), .Z(n7352) );
  XOR U9349 ( .A(n9765), .B(n9766), .Z(n6748) );
  ANDN U9350 ( .B(n7469), .A(n6747), .Z(n9764) );
  XNOR U9351 ( .A(n9767), .B(n9768), .Z(n6747) );
  XOR U9352 ( .A(n9769), .B(n9770), .Z(n7469) );
  XNOR U9353 ( .A(n9771), .B(n6751), .Z(n2632) );
  XOR U9354 ( .A(n9772), .B(n9773), .Z(n6751) );
  AND U9355 ( .A(n6752), .B(n9706), .Z(n9771) );
  XOR U9356 ( .A(n9774), .B(n9370), .Z(n9706) );
  XNOR U9357 ( .A(n9775), .B(n9776), .Z(n6752) );
  XOR U9358 ( .A(n3305), .B(n9777), .Z(n9762) );
  XNOR U9359 ( .A(n5227), .B(n6741), .Z(n9777) );
  XNOR U9360 ( .A(n9778), .B(n6756), .Z(n6741) );
  XNOR U9361 ( .A(n9779), .B(n9780), .Z(n6756) );
  AND U9362 ( .A(n7467), .B(n7466), .Z(n9778) );
  XNOR U9363 ( .A(n9781), .B(n9782), .Z(n7466) );
  XNOR U9364 ( .A(n9783), .B(n9784), .Z(n7467) );
  XNOR U9365 ( .A(n9785), .B(n6760), .Z(n5227) );
  XOR U9366 ( .A(n9786), .B(n9584), .Z(n6760) );
  AND U9367 ( .A(n6761), .B(n9787), .Z(n9785) );
  XOR U9368 ( .A(n9788), .B(n7359), .Z(n3305) );
  IV U9369 ( .A(n6764), .Z(n7359) );
  XOR U9370 ( .A(n9789), .B(n9790), .Z(n6764) );
  ANDN U9371 ( .B(n6765), .A(n7461), .Z(n9788) );
  XOR U9372 ( .A(n9791), .B(n9077), .Z(n7461) );
  XOR U9373 ( .A(n9792), .B(n9793), .Z(n6765) );
  XOR U9374 ( .A(n9794), .B(n9795), .Z(n5921) );
  XOR U9375 ( .A(n1833), .B(n5174), .Z(n9795) );
  XNOR U9376 ( .A(n9796), .B(n7524), .Z(n5174) );
  AND U9377 ( .A(n6784), .B(n7451), .Z(n9796) );
  IV U9378 ( .A(n7523), .Z(n7451) );
  XOR U9379 ( .A(n9797), .B(n9798), .Z(n7523) );
  XNOR U9380 ( .A(n9799), .B(n9800), .Z(n6784) );
  XOR U9381 ( .A(n9801), .B(n7518), .Z(n1833) );
  AND U9382 ( .A(n6792), .B(n7519), .Z(n9801) );
  XNOR U9383 ( .A(n9802), .B(n9803), .Z(n7519) );
  XOR U9384 ( .A(n9804), .B(n9805), .Z(n6792) );
  XNOR U9385 ( .A(n4083), .B(n9806), .Z(n9794) );
  XOR U9386 ( .A(n7496), .B(n3576), .Z(n9806) );
  XOR U9387 ( .A(n9807), .B(n9808), .Z(n3576) );
  ANDN U9388 ( .B(n7445), .A(n6788), .Z(n9807) );
  XOR U9389 ( .A(n9809), .B(n9810), .Z(n6788) );
  XOR U9390 ( .A(n9811), .B(n7515), .Z(n7496) );
  ANDN U9391 ( .B(n7516), .A(n6776), .Z(n9811) );
  XNOR U9392 ( .A(n9555), .B(n9812), .Z(n6776) );
  XNOR U9393 ( .A(n9813), .B(n9261), .Z(n7516) );
  XNOR U9394 ( .A(n9814), .B(n7526), .Z(n4083) );
  AND U9395 ( .A(n6773), .B(n7527), .Z(n9814) );
  XNOR U9396 ( .A(n9815), .B(n9704), .Z(n7527) );
  XNOR U9397 ( .A(n9816), .B(n9817), .Z(n6773) );
  XNOR U9398 ( .A(n9818), .B(n6761), .Z(n7464) );
  XNOR U9399 ( .A(n9819), .B(n9820), .Z(n6761) );
  ANDN U9400 ( .B(n9702), .A(n7349), .Z(n9818) );
  XOR U9401 ( .A(n9821), .B(n9822), .Z(n7349) );
  IV U9402 ( .A(n9787), .Z(n9702) );
  XOR U9403 ( .A(n9823), .B(n9824), .Z(n9787) );
  XNOR U9404 ( .A(n9825), .B(n4189), .Z(n1207) );
  IV U9405 ( .A(n1664), .Z(n4189) );
  XOR U9406 ( .A(n9826), .B(n9827), .Z(n8289) );
  XNOR U9407 ( .A(n3402), .B(n4997), .Z(n9827) );
  XNOR U9408 ( .A(n9828), .B(n7308), .Z(n4997) );
  ANDN U9409 ( .B(n9750), .A(n7307), .Z(n9828) );
  XNOR U9410 ( .A(n9829), .B(n8342), .Z(n3402) );
  AND U9411 ( .A(n8343), .B(n9745), .Z(n9829) );
  XNOR U9412 ( .A(n2351), .B(n9830), .Z(n9826) );
  XOR U9413 ( .A(n3944), .B(n7300), .Z(n9830) );
  XOR U9414 ( .A(n9831), .B(n8564), .Z(n7300) );
  XOR U9415 ( .A(n9832), .B(n7313), .Z(n3944) );
  NOR U9416 ( .A(n7314), .B(n9742), .Z(n9832) );
  XOR U9417 ( .A(n9833), .B(n7317), .Z(n2351) );
  ANDN U9418 ( .B(n9834), .A(n7318), .Z(n9833) );
  XNOR U9419 ( .A(n9835), .B(n9836), .Z(n6182) );
  XNOR U9420 ( .A(n2033), .B(n3555), .Z(n9836) );
  XOR U9421 ( .A(n9837), .B(n9838), .Z(n3555) );
  XOR U9422 ( .A(n9840), .B(n9841), .Z(n2033) );
  AND U9423 ( .A(n9842), .B(n8396), .Z(n9840) );
  IV U9424 ( .A(n9843), .Z(n8396) );
  XOR U9425 ( .A(n9844), .B(n9845), .Z(n9835) );
  XOR U9426 ( .A(n5310), .B(n5083), .Z(n9845) );
  XNOR U9427 ( .A(n9846), .B(n9847), .Z(n5083) );
  ANDN U9428 ( .B(n7383), .A(n9848), .Z(n9846) );
  IV U9429 ( .A(n9849), .Z(n7383) );
  XNOR U9430 ( .A(n9850), .B(n9851), .Z(n5310) );
  XNOR U9431 ( .A(n9853), .B(n6049), .Z(out[1024]) );
  XNOR U9432 ( .A(n8484), .B(n2518), .Z(n6049) );
  XNOR U9433 ( .A(n9854), .B(n9855), .Z(n2518) );
  XOR U9434 ( .A(n9856), .B(n9857), .Z(n8484) );
  NOR U9435 ( .A(n8423), .B(n9858), .Z(n9856) );
  ANDN U9436 ( .B(n1210), .A(n1212), .Z(n9853) );
  XNOR U9437 ( .A(n9859), .B(n1672), .Z(n1212) );
  XOR U9438 ( .A(n9860), .B(n9861), .Z(n8560) );
  XNOR U9439 ( .A(n3405), .B(n5000), .Z(n9861) );
  XNOR U9440 ( .A(n9862), .B(n7384), .Z(n5000) );
  AND U9441 ( .A(n9847), .B(n7385), .Z(n9862) );
  XNOR U9442 ( .A(n9863), .B(n8397), .Z(n3405) );
  ANDN U9443 ( .B(n8398), .A(n9841), .Z(n9863) );
  XOR U9444 ( .A(n2358), .B(n9864), .Z(n9860) );
  XOR U9445 ( .A(n7377), .B(n3948), .Z(n9864) );
  XOR U9446 ( .A(n9865), .B(n7390), .Z(n3948) );
  ANDN U9447 ( .B(n7391), .A(n9838), .Z(n9865) );
  XOR U9448 ( .A(n9866), .B(n9315), .Z(n7377) );
  ANDN U9449 ( .B(n9316), .A(n9851), .Z(n9866) );
  XNOR U9450 ( .A(n9867), .B(n7395), .Z(n2358) );
  AND U9451 ( .A(n9868), .B(n9869), .Z(n9867) );
  XNOR U9452 ( .A(n9870), .B(n9871), .Z(n6186) );
  XOR U9453 ( .A(n2036), .B(n3558), .Z(n9871) );
  XOR U9454 ( .A(n9872), .B(n9873), .Z(n3558) );
  NOR U9455 ( .A(n7433), .B(n9874), .Z(n9872) );
  XNOR U9456 ( .A(n9875), .B(n9876), .Z(n2036) );
  AND U9457 ( .A(n9877), .B(n8469), .Z(n9875) );
  IV U9458 ( .A(n9878), .Z(n8469) );
  XNOR U9459 ( .A(n9879), .B(n9880), .Z(n9870) );
  XOR U9460 ( .A(n5318), .B(n5109), .Z(n9880) );
  XNOR U9461 ( .A(n9881), .B(n9882), .Z(n5109) );
  ANDN U9462 ( .B(n9883), .A(n7427), .Z(n9881) );
  XNOR U9463 ( .A(n9884), .B(n9885), .Z(n5318) );
  ANDN U9464 ( .B(n9886), .A(n9887), .Z(n9884) );
  XNOR U9465 ( .A(n7521), .B(n3501), .Z(n1210) );
  IV U9466 ( .A(n2605), .Z(n3501) );
  XNOR U9467 ( .A(n5926), .B(n6332), .Z(n2605) );
  XNOR U9468 ( .A(n9888), .B(n9889), .Z(n6332) );
  XNOR U9469 ( .A(n2639), .B(n5328), .Z(n9889) );
  XOR U9470 ( .A(n9890), .B(n7448), .Z(n5328) );
  IV U9471 ( .A(n6774), .Z(n7448) );
  XOR U9472 ( .A(n9069), .B(n9891), .Z(n6774) );
  AND U9473 ( .A(n6775), .B(n7526), .Z(n9890) );
  XNOR U9474 ( .A(n9892), .B(n9893), .Z(n7526) );
  XNOR U9475 ( .A(n9894), .B(n9895), .Z(n6775) );
  XOR U9476 ( .A(n9896), .B(n6781), .Z(n2639) );
  XNOR U9477 ( .A(n9769), .B(n9897), .Z(n6781) );
  ANDN U9478 ( .B(n6780), .A(n7515), .Z(n9896) );
  XNOR U9479 ( .A(n9086), .B(n9898), .Z(n7515) );
  XNOR U9480 ( .A(n9899), .B(n9900), .Z(n6780) );
  XNOR U9481 ( .A(n3309), .B(n9901), .Z(n9888) );
  XNOR U9482 ( .A(n5262), .B(n6768), .Z(n9901) );
  XNOR U9483 ( .A(n9902), .B(n6786), .Z(n6768) );
  XOR U9484 ( .A(n9903), .B(n9904), .Z(n6786) );
  ANDN U9485 ( .B(n7524), .A(n6785), .Z(n9902) );
  XNOR U9486 ( .A(n9905), .B(n9906), .Z(n6785) );
  XNOR U9487 ( .A(n9907), .B(n9908), .Z(n7524) );
  XNOR U9488 ( .A(n9909), .B(n6789), .Z(n5262) );
  XNOR U9489 ( .A(n9910), .B(n9694), .Z(n6789) );
  ANDN U9490 ( .B(n6790), .A(n9808), .Z(n9909) );
  XNOR U9491 ( .A(n9911), .B(n6793), .Z(n3309) );
  XNOR U9492 ( .A(n9912), .B(n9913), .Z(n6793) );
  NOR U9493 ( .A(n7518), .B(n6794), .Z(n9911) );
  XNOR U9494 ( .A(n9914), .B(n9915), .Z(n6794) );
  XOR U9495 ( .A(n9916), .B(n9917), .Z(n7518) );
  XOR U9496 ( .A(n9918), .B(n9919), .Z(n5926) );
  XOR U9497 ( .A(n1838), .B(n5176), .Z(n9919) );
  XNOR U9498 ( .A(n9920), .B(n7596), .Z(n5176) );
  ANDN U9499 ( .B(n7597), .A(n6811), .Z(n9920) );
  XNOR U9500 ( .A(n9921), .B(n9922), .Z(n6811) );
  XNOR U9501 ( .A(n9923), .B(n9924), .Z(n7597) );
  XNOR U9502 ( .A(n9925), .B(n7592), .Z(n1838) );
  AND U9503 ( .A(n6819), .B(n7508), .Z(n9925) );
  IV U9504 ( .A(n7591), .Z(n7508) );
  XOR U9505 ( .A(n9926), .B(n9927), .Z(n7591) );
  XOR U9506 ( .A(n9928), .B(n9114), .Z(n6819) );
  XNOR U9507 ( .A(n4089), .B(n9929), .Z(n9918) );
  XNOR U9508 ( .A(n7573), .B(n3581), .Z(n9929) );
  XOR U9509 ( .A(n9930), .B(n9931), .Z(n3581) );
  ANDN U9510 ( .B(n7506), .A(n6815), .Z(n9930) );
  XOR U9511 ( .A(n9166), .B(n9932), .Z(n6815) );
  AND U9512 ( .A(n7510), .B(n7511), .Z(n9933) );
  XNOR U9513 ( .A(n9935), .B(n9661), .Z(n7511) );
  XOR U9514 ( .A(n9936), .B(n7599), .Z(n4089) );
  ANDN U9515 ( .B(n7600), .A(n6802), .Z(n9936) );
  XOR U9516 ( .A(n9937), .B(n9938), .Z(n6802) );
  XOR U9517 ( .A(n9939), .B(n9810), .Z(n7600) );
  XOR U9518 ( .A(n9940), .B(n6790), .Z(n7521) );
  XOR U9519 ( .A(n9941), .B(n9942), .Z(n6790) );
  ANDN U9520 ( .B(n9808), .A(n7445), .Z(n9940) );
  XOR U9521 ( .A(n9943), .B(n9944), .Z(n7445) );
  XNOR U9522 ( .A(n9945), .B(n9946), .Z(n9808) );
  XOR U9523 ( .A(n9947), .B(n6052), .Z(out[1023]) );
  XOR U9524 ( .A(n7594), .B(n2610), .Z(n6052) );
  XOR U9525 ( .A(n9948), .B(n6816), .Z(n7594) );
  ANDN U9526 ( .B(n9931), .A(n7506), .Z(n9948) );
  XOR U9527 ( .A(n9949), .B(n9950), .Z(n7506) );
  IV U9528 ( .A(n9951), .Z(n9931) );
  ANDN U9529 ( .B(n5561), .A(n5559), .Z(n9947) );
  XNOR U9530 ( .A(n9952), .B(n3735), .Z(n5559) );
  IV U9531 ( .A(n1677), .Z(n3735) );
  XOR U9532 ( .A(n9953), .B(n9954), .Z(n9311) );
  XOR U9533 ( .A(n3408), .B(n5004), .Z(n9954) );
  XNOR U9534 ( .A(n9955), .B(n7429), .Z(n5004) );
  AND U9535 ( .A(n9882), .B(n9956), .Z(n9955) );
  XNOR U9536 ( .A(n9957), .B(n8471), .Z(n3408) );
  ANDN U9537 ( .B(n9876), .A(n8470), .Z(n9957) );
  XOR U9538 ( .A(n2365), .B(n9958), .Z(n9953) );
  XOR U9539 ( .A(n7422), .B(n3953), .Z(n9958) );
  XNOR U9540 ( .A(n9959), .B(n7435), .Z(n3953) );
  XNOR U9541 ( .A(n9960), .B(n9961), .Z(n7422) );
  NOR U9542 ( .A(n9962), .B(n9885), .Z(n9960) );
  XNOR U9543 ( .A(n9963), .B(n7439), .Z(n2365) );
  AND U9544 ( .A(n9964), .B(n9965), .Z(n9963) );
  XNOR U9545 ( .A(n9966), .B(n9967), .Z(n6190) );
  XNOR U9546 ( .A(n5322), .B(n3563), .Z(n9967) );
  XOR U9547 ( .A(n9968), .B(n9969), .Z(n3563) );
  ANDN U9548 ( .B(n9970), .A(n7540), .Z(n9968) );
  XNOR U9549 ( .A(n9971), .B(n9972), .Z(n5322) );
  ANDN U9550 ( .B(n9973), .A(n9974), .Z(n9971) );
  XNOR U9551 ( .A(n9975), .B(n9976), .Z(n9966) );
  XNOR U9552 ( .A(n2040), .B(n5135), .Z(n9976) );
  XNOR U9553 ( .A(n9977), .B(n9978), .Z(n5135) );
  XNOR U9554 ( .A(n9980), .B(n9981), .Z(n2040) );
  NOR U9555 ( .A(n9982), .B(n8593), .Z(n9980) );
  XOR U9556 ( .A(n9051), .B(n4834), .Z(n5561) );
  XOR U9557 ( .A(n9983), .B(n8064), .Z(n4834) );
  XNOR U9558 ( .A(n9984), .B(n9985), .Z(n8064) );
  XOR U9559 ( .A(n5353), .B(n3802), .Z(n9985) );
  XOR U9560 ( .A(n9986), .B(n9987), .Z(n3802) );
  AND U9561 ( .A(n7940), .B(n9988), .Z(n9986) );
  XNOR U9562 ( .A(n9989), .B(n9990), .Z(n7940) );
  XNOR U9563 ( .A(n9991), .B(n9147), .Z(n5353) );
  ANDN U9564 ( .B(n7935), .A(n7936), .Z(n9991) );
  XNOR U9565 ( .A(n9682), .B(n9992), .Z(n7936) );
  XNOR U9566 ( .A(n9993), .B(n9994), .Z(n7935) );
  XOR U9567 ( .A(n6146), .B(n9995), .Z(n9984) );
  XOR U9568 ( .A(n2217), .B(n4807), .Z(n9995) );
  XOR U9569 ( .A(n9996), .B(n9154), .Z(n4807) );
  IV U9570 ( .A(n9997), .Z(n9154) );
  AND U9571 ( .A(n8068), .B(n9155), .Z(n9996) );
  XOR U9572 ( .A(n9998), .B(n9529), .Z(n9155) );
  XNOR U9573 ( .A(n9999), .B(n10000), .Z(n8068) );
  XNOR U9574 ( .A(n10001), .B(n9151), .Z(n2217) );
  AND U9575 ( .A(n7925), .B(n9236), .Z(n10001) );
  XOR U9576 ( .A(n10002), .B(n10003), .Z(n9236) );
  XNOR U9577 ( .A(n10004), .B(n10005), .Z(n7925) );
  XNOR U9578 ( .A(n10006), .B(n9158), .Z(n6146) );
  ANDN U9579 ( .B(n7929), .A(n7930), .Z(n10006) );
  XNOR U9580 ( .A(n10007), .B(n10008), .Z(n7930) );
  XNOR U9581 ( .A(n10009), .B(n10010), .Z(n7929) );
  XOR U9582 ( .A(n10011), .B(n9140), .Z(n9051) );
  ANDN U9583 ( .B(n8002), .A(n8000), .Z(n10011) );
  XOR U9584 ( .A(n10012), .B(n6055), .Z(out[1022]) );
  IV U9585 ( .A(n6408), .Z(n6055) );
  XOR U9586 ( .A(n7694), .B(n2617), .Z(n6408) );
  XNOR U9587 ( .A(n5936), .B(n6575), .Z(n2617) );
  XNOR U9588 ( .A(n10013), .B(n10014), .Z(n6575) );
  XNOR U9589 ( .A(n2653), .B(n5339), .Z(n10014) );
  XOR U9590 ( .A(n10015), .B(n6830), .Z(n5339) );
  XNOR U9591 ( .A(n10016), .B(n10017), .Z(n6830) );
  NOR U9592 ( .A(n7699), .B(n6829), .Z(n10015) );
  XNOR U9593 ( .A(n10018), .B(n10019), .Z(n6829) );
  XNOR U9594 ( .A(n10020), .B(n6837), .Z(n2653) );
  XOR U9595 ( .A(n10021), .B(n10022), .Z(n6837) );
  AND U9596 ( .A(n6838), .B(n10023), .Z(n10020) );
  XNOR U9597 ( .A(n10024), .B(n10025), .Z(n6838) );
  XNOR U9598 ( .A(n3320), .B(n10026), .Z(n10013) );
  XOR U9599 ( .A(n5364), .B(n6823), .Z(n10026) );
  XNOR U9600 ( .A(n10027), .B(n6854), .Z(n6823) );
  XNOR U9601 ( .A(n9608), .B(n10028), .Z(n6854) );
  ANDN U9602 ( .B(n7696), .A(n7697), .Z(n10027) );
  XOR U9603 ( .A(n10029), .B(n10030), .Z(n7696) );
  XNOR U9604 ( .A(n10031), .B(n6844), .Z(n5364) );
  XOR U9605 ( .A(n10032), .B(n9924), .Z(n6844) );
  AND U9606 ( .A(n10033), .B(n10034), .Z(n10031) );
  XNOR U9607 ( .A(n10035), .B(n6848), .Z(n3320) );
  XOR U9608 ( .A(n10036), .B(n10037), .Z(n6848) );
  NOR U9609 ( .A(n7691), .B(n6847), .Z(n10035) );
  XNOR U9610 ( .A(n9710), .B(n10038), .Z(n6847) );
  XOR U9611 ( .A(n10039), .B(n10040), .Z(n5936) );
  XOR U9612 ( .A(n1846), .B(n5181), .Z(n10040) );
  XNOR U9613 ( .A(n10041), .B(n7762), .Z(n5181) );
  AND U9614 ( .A(n7186), .B(n7763), .Z(n10041) );
  XNOR U9615 ( .A(n10042), .B(n10043), .Z(n7763) );
  XOR U9616 ( .A(n10044), .B(n10045), .Z(n7186) );
  XNOR U9617 ( .A(n10046), .B(n7756), .Z(n1846) );
  AND U9618 ( .A(n6880), .B(n7757), .Z(n10046) );
  XOR U9619 ( .A(n10047), .B(n10048), .Z(n7757) );
  XNOR U9620 ( .A(n10049), .B(n10050), .Z(n6880) );
  XNOR U9621 ( .A(n4095), .B(n10051), .Z(n10039) );
  XNOR U9622 ( .A(n7748), .B(n3591), .Z(n10051) );
  XNOR U9623 ( .A(n10052), .B(n10053), .Z(n3591) );
  ANDN U9624 ( .B(n7685), .A(n6876), .Z(n10052) );
  XOR U9625 ( .A(n10054), .B(n10055), .Z(n6876) );
  XOR U9626 ( .A(n10056), .B(n7753), .Z(n7748) );
  AND U9627 ( .A(n6867), .B(n7754), .Z(n10056) );
  XNOR U9628 ( .A(n10057), .B(n9551), .Z(n7754) );
  XNOR U9629 ( .A(n9894), .B(n10058), .Z(n6867) );
  XNOR U9630 ( .A(n10059), .B(n7765), .Z(n4095) );
  ANDN U9631 ( .B(n7766), .A(n6864), .Z(n10059) );
  XOR U9632 ( .A(n10060), .B(n10061), .Z(n6864) );
  XOR U9633 ( .A(n10062), .B(n9278), .Z(n7766) );
  XOR U9634 ( .A(n10063), .B(n6843), .Z(n7694) );
  IV U9635 ( .A(n10034), .Z(n6843) );
  XOR U9636 ( .A(n10064), .B(n10065), .Z(n10034) );
  ANDN U9637 ( .B(n7582), .A(n10033), .Z(n10063) );
  IV U9638 ( .A(n10066), .Z(n7582) );
  ANDN U9639 ( .B(n5565), .A(n5563), .Z(n10012) );
  XOR U9640 ( .A(n10067), .B(n1682), .Z(n5563) );
  XNOR U9641 ( .A(n10068), .B(n6194), .Z(n1682) );
  XNOR U9642 ( .A(n10069), .B(n10070), .Z(n6194) );
  XNOR U9643 ( .A(n5326), .B(n3570), .Z(n10070) );
  XOR U9644 ( .A(n10071), .B(n10072), .Z(n3570) );
  AND U9645 ( .A(n10073), .B(n7620), .Z(n10071) );
  XNOR U9646 ( .A(n10074), .B(n10075), .Z(n5326) );
  AND U9647 ( .A(n10076), .B(n7616), .Z(n10074) );
  XOR U9648 ( .A(n10077), .B(n10078), .Z(n10069) );
  XNOR U9649 ( .A(n2045), .B(n5167), .Z(n10078) );
  XNOR U9650 ( .A(n10079), .B(n10080), .Z(n5167) );
  ANDN U9651 ( .B(n10081), .A(n7607), .Z(n10079) );
  XNOR U9652 ( .A(n10082), .B(n10083), .Z(n2045) );
  NOR U9653 ( .A(n8650), .B(n10084), .Z(n10082) );
  XNOR U9654 ( .A(n9144), .B(n2012), .Z(n5565) );
  IV U9655 ( .A(n5281), .Z(n2012) );
  XOR U9656 ( .A(n10085), .B(n8126), .Z(n5281) );
  XNOR U9657 ( .A(n10086), .B(n10087), .Z(n8126) );
  XOR U9658 ( .A(n5356), .B(n3808), .Z(n10087) );
  XNOR U9659 ( .A(n10088), .B(n10089), .Z(n3808) );
  ANDN U9660 ( .B(n10090), .A(n8589), .Z(n10088) );
  XNOR U9661 ( .A(n10091), .B(n9181), .Z(n8589) );
  XNOR U9662 ( .A(n10092), .B(n9243), .Z(n5356) );
  AND U9663 ( .A(n8582), .B(n9244), .Z(n10092) );
  XOR U9664 ( .A(n9506), .B(n10093), .Z(n9244) );
  IV U9665 ( .A(n10094), .Z(n9506) );
  XOR U9666 ( .A(n10095), .B(n10096), .Z(n8582) );
  XNOR U9667 ( .A(n6151), .B(n10097), .Z(n10086) );
  XNOR U9668 ( .A(n2230), .B(n4836), .Z(n10097) );
  XNOR U9669 ( .A(n10098), .B(n9252), .Z(n4836) );
  AND U9670 ( .A(n8586), .B(n8584), .Z(n10098) );
  IV U9671 ( .A(n9251), .Z(n8584) );
  XNOR U9672 ( .A(n10099), .B(n9353), .Z(n9251) );
  XNOR U9673 ( .A(n10100), .B(n10101), .Z(n8586) );
  XNOR U9674 ( .A(n10102), .B(n9248), .Z(n2230) );
  ANDN U9675 ( .B(n8573), .A(n8571), .Z(n10102) );
  XOR U9676 ( .A(n9101), .B(n10103), .Z(n8571) );
  XNOR U9677 ( .A(n10104), .B(n10105), .Z(n8573) );
  XNOR U9678 ( .A(n10106), .B(n9255), .Z(n6151) );
  AND U9679 ( .A(n8576), .B(n8575), .Z(n10106) );
  XNOR U9680 ( .A(n10107), .B(n10108), .Z(n8575) );
  XNOR U9681 ( .A(n9499), .B(n10109), .Z(n8576) );
  IV U9682 ( .A(n10110), .Z(n9499) );
  XOR U9683 ( .A(n10111), .B(n9234), .Z(n9144) );
  AND U9684 ( .A(n9987), .B(n7939), .Z(n10111) );
  IV U9685 ( .A(n9988), .Z(n7939) );
  XOR U9686 ( .A(n10112), .B(n10113), .Z(n9988) );
  XOR U9687 ( .A(n10114), .B(n6064), .Z(out[1021]) );
  IV U9688 ( .A(n6435), .Z(n6064) );
  XOR U9689 ( .A(n7759), .B(n2624), .Z(n6435) );
  XNOR U9690 ( .A(n5941), .B(n6851), .Z(n2624) );
  XNOR U9691 ( .A(n10115), .B(n10116), .Z(n6851) );
  XOR U9692 ( .A(n2660), .B(n5343), .Z(n10116) );
  XOR U9693 ( .A(n10117), .B(n6866), .Z(n5343) );
  XOR U9694 ( .A(n10118), .B(n10119), .Z(n6866) );
  ANDN U9695 ( .B(n7765), .A(n6865), .Z(n10117) );
  XOR U9696 ( .A(n10120), .B(n10121), .Z(n6865) );
  XNOR U9697 ( .A(n10122), .B(n10123), .Z(n7765) );
  XNOR U9698 ( .A(n10124), .B(n6872), .Z(n2660) );
  XNOR U9699 ( .A(n10125), .B(n10126), .Z(n6872) );
  ANDN U9700 ( .B(n7753), .A(n6871), .Z(n10124) );
  XOR U9701 ( .A(n10127), .B(n10128), .Z(n6871) );
  XOR U9702 ( .A(n9398), .B(n10129), .Z(n7753) );
  XOR U9703 ( .A(n3323), .B(n10130), .Z(n10115) );
  XNOR U9704 ( .A(n5416), .B(n6859), .Z(n10130) );
  XNOR U9705 ( .A(n10131), .B(n7187), .Z(n6859) );
  XOR U9706 ( .A(n10132), .B(n9718), .Z(n7187) );
  AND U9707 ( .A(n7762), .B(n7761), .Z(n10131) );
  XOR U9708 ( .A(n10133), .B(n10134), .Z(n7761) );
  XNOR U9709 ( .A(n10135), .B(n10136), .Z(n7762) );
  XNOR U9710 ( .A(n10137), .B(n6877), .Z(n5416) );
  XOR U9711 ( .A(n10138), .B(n10139), .Z(n6877) );
  AND U9712 ( .A(n10053), .B(n10140), .Z(n10137) );
  XOR U9713 ( .A(n10141), .B(n7683), .Z(n3323) );
  XOR U9714 ( .A(n10142), .B(n10143), .Z(n7683) );
  AND U9715 ( .A(n6882), .B(n7756), .Z(n10141) );
  XOR U9716 ( .A(n9526), .B(n10144), .Z(n7756) );
  XNOR U9717 ( .A(n10145), .B(n9817), .Z(n6882) );
  XOR U9718 ( .A(n10146), .B(n10147), .Z(n5941) );
  XNOR U9719 ( .A(n5183), .B(n1851), .Z(n10147) );
  XNOR U9720 ( .A(n10148), .B(n7799), .Z(n1851) );
  AND U9721 ( .A(n6904), .B(n7800), .Z(n10148) );
  XOR U9722 ( .A(n10149), .B(n10150), .Z(n7800) );
  XNOR U9723 ( .A(n10151), .B(n9994), .Z(n6904) );
  XNOR U9724 ( .A(n10152), .B(n7808), .Z(n5183) );
  AND U9725 ( .A(n7911), .B(n7909), .Z(n10152) );
  IV U9726 ( .A(n7807), .Z(n7909) );
  XOR U9727 ( .A(n9094), .B(n10155), .Z(n7911) );
  XNOR U9728 ( .A(n3595), .B(n10156), .Z(n10146) );
  XNOR U9729 ( .A(n7793), .B(n4099), .Z(n10156) );
  XNOR U9730 ( .A(n10157), .B(n7811), .Z(n4099) );
  NOR U9731 ( .A(n6889), .B(n7810), .Z(n10157) );
  XOR U9732 ( .A(n10158), .B(n10055), .Z(n7810) );
  XNOR U9733 ( .A(n10159), .B(n10160), .Z(n6889) );
  XOR U9734 ( .A(n10161), .B(n7804), .Z(n7793) );
  NOR U9735 ( .A(n7803), .B(n6892), .Z(n10161) );
  XOR U9736 ( .A(n10162), .B(n10163), .Z(n6892) );
  XNOR U9737 ( .A(n10164), .B(n10165), .Z(n7803) );
  XNOR U9738 ( .A(n10166), .B(n10167), .Z(n3595) );
  ANDN U9739 ( .B(n7916), .A(n6900), .Z(n10166) );
  XOR U9740 ( .A(n10168), .B(n10169), .Z(n6900) );
  XOR U9741 ( .A(n10170), .B(n6878), .Z(n7759) );
  IV U9742 ( .A(n10140), .Z(n6878) );
  XNOR U9743 ( .A(n10171), .B(n10172), .Z(n10140) );
  NOR U9744 ( .A(n7685), .B(n10053), .Z(n10170) );
  XNOR U9745 ( .A(n10173), .B(n10174), .Z(n10053) );
  XNOR U9746 ( .A(n10175), .B(n9366), .Z(n7685) );
  IV U9747 ( .A(n9994), .Z(n9366) );
  ANDN U9748 ( .B(n5569), .A(n5567), .Z(n10114) );
  XOR U9749 ( .A(n10176), .B(n1686), .Z(n5567) );
  XNOR U9750 ( .A(n10177), .B(n6198), .Z(n1686) );
  XNOR U9751 ( .A(n10178), .B(n10179), .Z(n6198) );
  XOR U9752 ( .A(n5331), .B(n3577), .Z(n10179) );
  XOR U9753 ( .A(n10180), .B(n10181), .Z(n3577) );
  ANDN U9754 ( .B(n7668), .A(n10182), .Z(n10180) );
  XNOR U9755 ( .A(n10183), .B(n10184), .Z(n5331) );
  AND U9756 ( .A(n7664), .B(n10185), .Z(n10183) );
  XOR U9757 ( .A(n10186), .B(n10187), .Z(n10178) );
  XNOR U9758 ( .A(n2048), .B(n5196), .Z(n10187) );
  XNOR U9759 ( .A(n10188), .B(n10189), .Z(n5196) );
  ANDN U9760 ( .B(n10190), .A(n7655), .Z(n10188) );
  XNOR U9761 ( .A(n10191), .B(n10192), .Z(n2048) );
  AND U9762 ( .A(n10193), .B(n8715), .Z(n10191) );
  XOR U9763 ( .A(n9240), .B(n2015), .Z(n5569) );
  XNOR U9764 ( .A(n7921), .B(n8180), .Z(n2015) );
  XNOR U9765 ( .A(n10194), .B(n10195), .Z(n8180) );
  XOR U9766 ( .A(n5361), .B(n3814), .Z(n10195) );
  XOR U9767 ( .A(n10196), .B(n10197), .Z(n3814) );
  AND U9768 ( .A(n9340), .B(n10198), .Z(n10196) );
  XNOR U9769 ( .A(n10199), .B(n10200), .Z(n9340) );
  XNOR U9770 ( .A(n10201), .B(n9424), .Z(n5361) );
  ANDN U9771 ( .B(n9425), .A(n9332), .Z(n10201) );
  XOR U9772 ( .A(n10202), .B(n10203), .Z(n9332) );
  XOR U9773 ( .A(n10204), .B(n10205), .Z(n9425) );
  XNOR U9774 ( .A(n6156), .B(n10206), .Z(n10194) );
  XOR U9775 ( .A(n2237), .B(n4873), .Z(n10206) );
  XNOR U9776 ( .A(n10207), .B(n9432), .Z(n4873) );
  AND U9777 ( .A(n9337), .B(n9433), .Z(n10207) );
  XOR U9778 ( .A(n10208), .B(n10209), .Z(n9433) );
  XNOR U9779 ( .A(n9116), .B(n10210), .Z(n9337) );
  XNOR U9780 ( .A(n10211), .B(n9429), .Z(n2237) );
  ANDN U9781 ( .B(n9324), .A(n9322), .Z(n10211) );
  XOR U9782 ( .A(n10212), .B(n10213), .Z(n9322) );
  XNOR U9783 ( .A(n10214), .B(n10215), .Z(n9324) );
  XNOR U9784 ( .A(n10216), .B(n10217), .Z(n6156) );
  AND U9785 ( .A(n9328), .B(n9437), .Z(n10216) );
  XNOR U9786 ( .A(n10218), .B(n10219), .Z(n9437) );
  XNOR U9787 ( .A(n10220), .B(n10221), .Z(n9328) );
  XOR U9788 ( .A(n10222), .B(n10223), .Z(n7921) );
  XOR U9789 ( .A(n1952), .B(n9407), .Z(n10223) );
  XOR U9790 ( .A(n10224), .B(n8581), .Z(n9407) );
  IV U9791 ( .A(n9418), .Z(n8581) );
  XOR U9792 ( .A(n10225), .B(n10226), .Z(n9418) );
  ANDN U9793 ( .B(n9242), .A(n9243), .Z(n10224) );
  XNOR U9794 ( .A(n10227), .B(n10228), .Z(n9243) );
  XNOR U9795 ( .A(n10229), .B(n10230), .Z(n9242) );
  XNOR U9796 ( .A(n10231), .B(n8577), .Z(n1952) );
  XNOR U9797 ( .A(n10232), .B(n10233), .Z(n8577) );
  NOR U9798 ( .A(n9254), .B(n9255), .Z(n10231) );
  XOR U9799 ( .A(n10234), .B(n10235), .Z(n9255) );
  XNOR U9800 ( .A(n10236), .B(n10174), .Z(n9254) );
  XOR U9801 ( .A(n3707), .B(n10237), .Z(n10222) );
  XOR U9802 ( .A(n5064), .B(n4174), .Z(n10237) );
  XOR U9803 ( .A(n10238), .B(n8590), .Z(n4174) );
  XNOR U9804 ( .A(n10204), .B(n10239), .Z(n8590) );
  NOR U9805 ( .A(n10089), .B(n9414), .Z(n10238) );
  XNOR U9806 ( .A(n10241), .B(n9668), .Z(n8585) );
  AND U9807 ( .A(n9252), .B(n10242), .Z(n10240) );
  IV U9808 ( .A(n9250), .Z(n10242) );
  XOR U9809 ( .A(n10212), .B(n10243), .Z(n9250) );
  IV U9810 ( .A(n9168), .Z(n10212) );
  XNOR U9811 ( .A(n10244), .B(n10245), .Z(n9252) );
  XOR U9812 ( .A(n10246), .B(n8572), .Z(n3707) );
  IV U9813 ( .A(n9416), .Z(n8572) );
  XNOR U9814 ( .A(n9894), .B(n10247), .Z(n9416) );
  ANDN U9815 ( .B(n9247), .A(n9248), .Z(n10246) );
  XOR U9816 ( .A(n10248), .B(n10249), .Z(n9248) );
  XNOR U9817 ( .A(n10250), .B(n10251), .Z(n9247) );
  XNOR U9818 ( .A(n10252), .B(n9414), .Z(n9240) );
  XNOR U9819 ( .A(n10253), .B(n10254), .Z(n9414) );
  AND U9820 ( .A(n10089), .B(n8588), .Z(n10252) );
  IV U9821 ( .A(n10090), .Z(n8588) );
  XNOR U9822 ( .A(n10255), .B(n10256), .Z(n10090) );
  XOR U9823 ( .A(n10257), .B(n9584), .Z(n10089) );
  XOR U9824 ( .A(n10258), .B(n6069), .Z(out[1020]) );
  XNOR U9825 ( .A(n7797), .B(n2631), .Z(n6069) );
  XNOR U9826 ( .A(n5946), .B(n7184), .Z(n2631) );
  XNOR U9827 ( .A(n10259), .B(n10260), .Z(n7184) );
  XNOR U9828 ( .A(n2667), .B(n5347), .Z(n10260) );
  XNOR U9829 ( .A(n10261), .B(n6890), .Z(n5347) );
  XNOR U9830 ( .A(n10262), .B(n10263), .Z(n6890) );
  AND U9831 ( .A(n7811), .B(n6891), .Z(n10261) );
  XOR U9832 ( .A(n10264), .B(n10265), .Z(n6891) );
  XNOR U9833 ( .A(n10266), .B(n10267), .Z(n7811) );
  XOR U9834 ( .A(n10268), .B(n6896), .Z(n2667) );
  XOR U9835 ( .A(n10269), .B(n10270), .Z(n6896) );
  ANDN U9836 ( .B(n6895), .A(n7804), .Z(n10268) );
  XNOR U9837 ( .A(n9532), .B(n10271), .Z(n7804) );
  XOR U9838 ( .A(n10272), .B(n10273), .Z(n6895) );
  XOR U9839 ( .A(n3327), .B(n10274), .Z(n10259) );
  XOR U9840 ( .A(n5467), .B(n6884), .Z(n10274) );
  XNOR U9841 ( .A(n10275), .B(n7910), .Z(n6884) );
  XNOR U9842 ( .A(n10276), .B(n10277), .Z(n7910) );
  AND U9843 ( .A(n7808), .B(n7919), .Z(n10275) );
  XNOR U9844 ( .A(n10278), .B(n10279), .Z(n7919) );
  XNOR U9845 ( .A(n10280), .B(n10281), .Z(n7808) );
  XOR U9846 ( .A(n10282), .B(n6902), .Z(n5467) );
  XNOR U9847 ( .A(n10283), .B(n10043), .Z(n6902) );
  AND U9848 ( .A(n10167), .B(n6901), .Z(n10282) );
  XNOR U9849 ( .A(n10284), .B(n6905), .Z(n3327) );
  XOR U9850 ( .A(n10285), .B(n10286), .Z(n6905) );
  AND U9851 ( .A(n6906), .B(n7799), .Z(n10284) );
  XNOR U9852 ( .A(n9597), .B(n10287), .Z(n7799) );
  XNOR U9853 ( .A(n10288), .B(n9938), .Z(n6906) );
  XOR U9854 ( .A(n10289), .B(n10290), .Z(n5946) );
  XNOR U9855 ( .A(n5185), .B(n1855), .Z(n10290) );
  XNOR U9856 ( .A(n10291), .B(n7889), .Z(n1855) );
  ANDN U9857 ( .B(n7890), .A(n8547), .Z(n10291) );
  XOR U9858 ( .A(n10292), .B(n10293), .Z(n7890) );
  XNOR U9859 ( .A(n10294), .B(n7898), .Z(n5185) );
  ANDN U9860 ( .B(n7899), .A(n8544), .Z(n10294) );
  XOR U9861 ( .A(n10295), .B(n10296), .Z(n7899) );
  XOR U9862 ( .A(n3600), .B(n10297), .Z(n10289) );
  XOR U9863 ( .A(n7882), .B(n4103), .Z(n10297) );
  XNOR U9864 ( .A(n10298), .B(n7903), .Z(n4103) );
  ANDN U9865 ( .B(n10299), .A(n7902), .Z(n10298) );
  XNOR U9866 ( .A(n10168), .B(n10300), .Z(n7902) );
  XNOR U9867 ( .A(n10301), .B(n7894), .Z(n7882) );
  ANDN U9868 ( .B(n7895), .A(n8551), .Z(n10301) );
  XOR U9869 ( .A(n10302), .B(n9766), .Z(n7895) );
  XNOR U9870 ( .A(n10303), .B(n10304), .Z(n3600) );
  NOR U9871 ( .A(n8555), .B(n8554), .Z(n10303) );
  XNOR U9872 ( .A(n10305), .B(n6901), .Z(n7797) );
  XOR U9873 ( .A(n10306), .B(n10307), .Z(n6901) );
  NOR U9874 ( .A(n10167), .B(n7916), .Z(n10305) );
  XNOR U9875 ( .A(n10094), .B(n10308), .Z(n7916) );
  XNOR U9876 ( .A(n10309), .B(n10310), .Z(n10167) );
  NOR U9877 ( .A(n5573), .B(n5571), .Z(n10258) );
  XOR U9878 ( .A(n10311), .B(n1690), .Z(n5571) );
  XNOR U9879 ( .A(n8654), .B(n6202), .Z(n1690) );
  XNOR U9880 ( .A(n10312), .B(n10313), .Z(n6202) );
  XOR U9881 ( .A(n5336), .B(n3583), .Z(n10313) );
  XNOR U9882 ( .A(n10314), .B(n10315), .Z(n3583) );
  AND U9883 ( .A(n10316), .B(n7741), .Z(n10314) );
  IV U9884 ( .A(n10317), .Z(n7741) );
  XNOR U9885 ( .A(n10318), .B(n10319), .Z(n5336) );
  AND U9886 ( .A(n7731), .B(n10320), .Z(n10318) );
  XOR U9887 ( .A(n10321), .B(n10322), .Z(n10312) );
  XNOR U9888 ( .A(n2051), .B(n5226), .Z(n10322) );
  XNOR U9889 ( .A(n10323), .B(n10324), .Z(n5226) );
  AND U9890 ( .A(n7735), .B(n10325), .Z(n10323) );
  XNOR U9891 ( .A(n10326), .B(n10327), .Z(n2051) );
  AND U9892 ( .A(n10328), .B(n8780), .Z(n10326) );
  XOR U9893 ( .A(n10329), .B(n10330), .Z(n8654) );
  XOR U9894 ( .A(n5017), .B(n7649), .Z(n10330) );
  XNOR U9895 ( .A(n10331), .B(n7665), .Z(n7649) );
  ANDN U9896 ( .B(n7666), .A(n10184), .Z(n10331) );
  XNOR U9897 ( .A(n10332), .B(n7656), .Z(n5017) );
  AND U9898 ( .A(n10189), .B(n10333), .Z(n10332) );
  XOR U9899 ( .A(n2387), .B(n10334), .Z(n10329) );
  XNOR U9900 ( .A(n3415), .B(n3962), .Z(n10334) );
  XNOR U9901 ( .A(n10335), .B(n7670), .Z(n3962) );
  NOR U9902 ( .A(n10181), .B(n7669), .Z(n10335) );
  XOR U9903 ( .A(n10336), .B(n8717), .Z(n3415) );
  AND U9904 ( .A(n8716), .B(n10337), .Z(n10336) );
  XOR U9905 ( .A(n10338), .B(n7661), .Z(n2387) );
  ANDN U9906 ( .B(n7662), .A(n10339), .Z(n10338) );
  XOR U9907 ( .A(n9421), .B(n2018), .Z(n5573) );
  XNOR U9908 ( .A(n8567), .B(n8234), .Z(n2018) );
  XNOR U9909 ( .A(n10340), .B(n10341), .Z(n8234) );
  XOR U9910 ( .A(n5370), .B(n3821), .Z(n10341) );
  XNOR U9911 ( .A(n10342), .B(n10343), .Z(n3821) );
  ANDN U9912 ( .B(n10344), .A(n9622), .Z(n10342) );
  XNOR U9913 ( .A(n10345), .B(n9461), .Z(n5370) );
  ANDN U9914 ( .B(n10346), .A(n10347), .Z(n10345) );
  XOR U9915 ( .A(n6161), .B(n10348), .Z(n10340) );
  XOR U9916 ( .A(n2244), .B(n4907), .Z(n10348) );
  XOR U9917 ( .A(n10349), .B(n10350), .Z(n4907) );
  AND U9918 ( .A(n9466), .B(n10351), .Z(n10349) );
  XNOR U9919 ( .A(n10352), .B(n9475), .Z(n2244) );
  ANDN U9920 ( .B(n9476), .A(n9626), .Z(n10352) );
  XOR U9921 ( .A(n10353), .B(n9472), .Z(n6161) );
  AND U9922 ( .A(n9614), .B(n10354), .Z(n10353) );
  XOR U9923 ( .A(n10355), .B(n10356), .Z(n8567) );
  XNOR U9924 ( .A(n1960), .B(n9445), .Z(n10356) );
  XOR U9925 ( .A(n10357), .B(n9456), .Z(n9445) );
  IV U9926 ( .A(n9333), .Z(n9456) );
  XNOR U9927 ( .A(n10358), .B(n9163), .Z(n9333) );
  ANDN U9928 ( .B(n9423), .A(n9424), .Z(n10357) );
  XOR U9929 ( .A(n10359), .B(n10360), .Z(n9424) );
  XNOR U9930 ( .A(n10361), .B(n10065), .Z(n9423) );
  XNOR U9931 ( .A(n10362), .B(n9327), .Z(n1960) );
  XNOR U9932 ( .A(n9535), .B(n10363), .Z(n9327) );
  ANDN U9933 ( .B(n10217), .A(n9435), .Z(n10362) );
  XNOR U9934 ( .A(n10309), .B(n10364), .Z(n9435) );
  IV U9935 ( .A(n9436), .Z(n10217) );
  XNOR U9936 ( .A(n10365), .B(n10251), .Z(n9436) );
  XOR U9937 ( .A(n3711), .B(n10366), .Z(n10355) );
  XNOR U9938 ( .A(n5066), .B(n4177), .Z(n10366) );
  XNOR U9939 ( .A(n10367), .B(n9341), .Z(n4177) );
  XOR U9940 ( .A(n10368), .B(n9678), .Z(n9341) );
  ANDN U9941 ( .B(n9453), .A(n10197), .Z(n10367) );
  XOR U9942 ( .A(n10369), .B(n9336), .Z(n5066) );
  IV U9943 ( .A(n9450), .Z(n9336) );
  XOR U9944 ( .A(n10370), .B(n10371), .Z(n9450) );
  NOR U9945 ( .A(n9431), .B(n9432), .Z(n10369) );
  XOR U9946 ( .A(n10372), .B(n10373), .Z(n9432) );
  XNOR U9947 ( .A(n10374), .B(n10375), .Z(n9431) );
  XNOR U9948 ( .A(n10376), .B(n9323), .Z(n3711) );
  XNOR U9949 ( .A(n10377), .B(n10378), .Z(n9323) );
  ANDN U9950 ( .B(n9428), .A(n9429), .Z(n10376) );
  XNOR U9951 ( .A(n10379), .B(n10380), .Z(n9429) );
  XOR U9952 ( .A(n10381), .B(n10382), .Z(n9428) );
  XOR U9953 ( .A(n10383), .B(n9453), .Z(n9421) );
  XNOR U9954 ( .A(n10384), .B(n10249), .Z(n9453) );
  AND U9955 ( .A(n10197), .B(n9339), .Z(n10383) );
  IV U9956 ( .A(n10198), .Z(n9339) );
  XNOR U9957 ( .A(n10385), .B(n10386), .Z(n10198) );
  XOR U9958 ( .A(n10387), .B(n9694), .Z(n10197) );
  XOR U9959 ( .A(n10388), .B(n4162), .Z(out[101]) );
  XNOR U9960 ( .A(n6949), .B(n2562), .Z(n4162) );
  XOR U9961 ( .A(n7993), .B(n10389), .Z(n2562) );
  XOR U9962 ( .A(n10390), .B(n10391), .Z(n7993) );
  XOR U9963 ( .A(n4333), .B(n2181), .Z(n10391) );
  XOR U9964 ( .A(n10392), .B(n8035), .Z(n2181) );
  NOR U9965 ( .A(n10393), .B(n10394), .Z(n10392) );
  XOR U9966 ( .A(n10395), .B(n8026), .Z(n4333) );
  IV U9967 ( .A(n10396), .Z(n8026) );
  ANDN U9968 ( .B(n6956), .A(n6955), .Z(n10395) );
  IV U9969 ( .A(n10397), .Z(n6956) );
  XOR U9970 ( .A(n5960), .B(n10398), .Z(n10390) );
  XNOR U9971 ( .A(n5507), .B(n3755), .Z(n10398) );
  XNOR U9972 ( .A(n10399), .B(n8032), .Z(n3755) );
  NOR U9973 ( .A(n6946), .B(n6945), .Z(n10399) );
  XOR U9974 ( .A(n10400), .B(n10401), .Z(n5507) );
  NOR U9975 ( .A(n6951), .B(n6953), .Z(n10400) );
  XNOR U9976 ( .A(n10402), .B(n8038), .Z(n5960) );
  AND U9977 ( .A(n6941), .B(n6943), .Z(n10402) );
  XNOR U9978 ( .A(n10403), .B(n10393), .Z(n6949) );
  ANDN U9979 ( .B(n10394), .A(n8034), .Z(n10403) );
  ANDN U9980 ( .B(n3574), .A(n3572), .Z(n10388) );
  XOR U9981 ( .A(n7425), .B(n2402), .Z(n3572) );
  XNOR U9982 ( .A(n10068), .B(n10404), .Z(n2402) );
  XOR U9983 ( .A(n10405), .B(n10406), .Z(n10068) );
  XNOR U9984 ( .A(n3410), .B(n5008), .Z(n10406) );
  XOR U9985 ( .A(n10407), .B(n7535), .Z(n5008) );
  AND U9986 ( .A(n9978), .B(n10408), .Z(n10407) );
  XOR U9987 ( .A(n10409), .B(n8594), .Z(n3410) );
  ANDN U9988 ( .B(n9981), .A(n8595), .Z(n10409) );
  XNOR U9989 ( .A(n2370), .B(n10410), .Z(n10405) );
  XOR U9990 ( .A(n7528), .B(n3956), .Z(n10410) );
  XOR U9991 ( .A(n10411), .B(n7541), .Z(n3956) );
  IV U9992 ( .A(n10412), .Z(n7541) );
  ANDN U9993 ( .B(n10415), .A(n9972), .Z(n10413) );
  XOR U9994 ( .A(n10416), .B(n7545), .Z(n2370) );
  ANDN U9995 ( .B(n10417), .A(n10418), .Z(n10416) );
  XNOR U9996 ( .A(n10419), .B(n9887), .Z(n7425) );
  XOR U9997 ( .A(n2336), .B(n9619), .Z(n3574) );
  XOR U9998 ( .A(n10420), .B(n10347), .Z(n9619) );
  ANDN U9999 ( .B(n10421), .A(n9460), .Z(n10420) );
  IV U10000 ( .A(n3395), .Z(n2336) );
  XOR U10001 ( .A(n6157), .B(n10422), .Z(n3395) );
  XOR U10002 ( .A(n10423), .B(n10424), .Z(n6157) );
  XOR U10003 ( .A(n3179), .B(n7190), .Z(n10424) );
  XNOR U10004 ( .A(n10425), .B(n9476), .Z(n7190) );
  XNOR U10005 ( .A(n10374), .B(n10426), .Z(n9476) );
  AND U10006 ( .A(n9626), .B(n10427), .Z(n10425) );
  XNOR U10007 ( .A(n10428), .B(n9372), .Z(n9626) );
  XOR U10008 ( .A(n10429), .B(n9471), .Z(n3179) );
  IV U10009 ( .A(n10354), .Z(n9471) );
  XOR U10010 ( .A(n10430), .B(n10431), .Z(n10354) );
  ANDN U10011 ( .B(n9615), .A(n9614), .Z(n10429) );
  XNOR U10012 ( .A(n9513), .B(n10432), .Z(n9614) );
  XOR U10013 ( .A(n5472), .B(n10433), .Z(n10423) );
  XNOR U10014 ( .A(n8232), .B(n2371), .Z(n10433) );
  XOR U10015 ( .A(n10434), .B(n10346), .Z(n2371) );
  IV U10016 ( .A(n9462), .Z(n10346) );
  XOR U10017 ( .A(n10435), .B(n10436), .Z(n9462) );
  AND U10018 ( .A(n10347), .B(n10437), .Z(n10434) );
  XNOR U10019 ( .A(n10438), .B(n10439), .Z(n10347) );
  XNOR U10020 ( .A(n10440), .B(n9466), .Z(n8232) );
  XOR U10021 ( .A(n10441), .B(n10442), .Z(n9466) );
  ANDN U10022 ( .B(n9617), .A(n9618), .Z(n10440) );
  IV U10023 ( .A(n10351), .Z(n9617) );
  XOR U10024 ( .A(n10443), .B(n9190), .Z(n10351) );
  XOR U10025 ( .A(n10444), .B(n10445), .Z(n5472) );
  AND U10026 ( .A(n9622), .B(n10446), .Z(n10444) );
  XNOR U10027 ( .A(n10447), .B(n10448), .Z(n9622) );
  XNOR U10028 ( .A(n10449), .B(n6074), .Z(out[1019]) );
  XOR U10029 ( .A(n7886), .B(n2638), .Z(n6074) );
  XNOR U10030 ( .A(n5956), .B(n7905), .Z(n2638) );
  XNOR U10031 ( .A(n10450), .B(n10451), .Z(n7905) );
  XNOR U10032 ( .A(n10452), .B(n5352), .Z(n10451) );
  XNOR U10033 ( .A(n10453), .B(n8559), .Z(n5352) );
  ANDN U10034 ( .B(n7903), .A(n7901), .Z(n10453) );
  XOR U10035 ( .A(n10454), .B(n10455), .Z(n7903) );
  XOR U10036 ( .A(n6909), .B(n10456), .Z(n10450) );
  XNOR U10037 ( .A(n2201), .B(n3332), .Z(n10456) );
  XNOR U10038 ( .A(n10457), .B(n8548), .Z(n3332) );
  AND U10039 ( .A(n7888), .B(n7889), .Z(n10457) );
  XOR U10040 ( .A(n9187), .B(n10458), .Z(n7889) );
  XNOR U10041 ( .A(n10459), .B(n8552), .Z(n2201) );
  ANDN U10042 ( .B(n7894), .A(n7893), .Z(n10459) );
  XNOR U10043 ( .A(n10460), .B(n10461), .Z(n7894) );
  XNOR U10044 ( .A(n10462), .B(n8545), .Z(n6909) );
  AND U10045 ( .A(n7897), .B(n7898), .Z(n10462) );
  XOR U10046 ( .A(n10463), .B(n10464), .Z(n7898) );
  XOR U10047 ( .A(n10465), .B(n10466), .Z(n5956) );
  XOR U10048 ( .A(n5188), .B(n1859), .Z(n10466) );
  XNOR U10049 ( .A(n10467), .B(n10468), .Z(n1859) );
  ANDN U10050 ( .B(n9300), .A(n6931), .Z(n10467) );
  XNOR U10051 ( .A(n9567), .B(n10469), .Z(n6931) );
  XNOR U10052 ( .A(n10470), .B(n10471), .Z(n5188) );
  ANDN U10053 ( .B(n9296), .A(n9297), .Z(n10470) );
  XOR U10054 ( .A(n10472), .B(n10473), .Z(n9297) );
  XNOR U10055 ( .A(n3604), .B(n10474), .Z(n10465) );
  XNOR U10056 ( .A(n7991), .B(n4106), .Z(n10474) );
  XNOR U10057 ( .A(n10475), .B(n10476), .Z(n4106) );
  NOR U10058 ( .A(n6917), .B(n9308), .Z(n10475) );
  XNOR U10059 ( .A(n10477), .B(n10478), .Z(n6917) );
  XOR U10060 ( .A(n10479), .B(n10480), .Z(n7991) );
  ANDN U10061 ( .B(n9303), .A(n6921), .Z(n10479) );
  XNOR U10062 ( .A(n10481), .B(n10121), .Z(n6921) );
  XOR U10063 ( .A(n10482), .B(n10483), .Z(n3604) );
  ANDN U10064 ( .B(n9305), .A(n6927), .Z(n10482) );
  XNOR U10065 ( .A(n9682), .B(n10484), .Z(n6927) );
  XOR U10066 ( .A(n10485), .B(n10486), .Z(n7886) );
  ANDN U10067 ( .B(n8554), .A(n10304), .Z(n10485) );
  XNOR U10068 ( .A(n10204), .B(n10487), .Z(n8554) );
  IV U10069 ( .A(n9567), .Z(n10204) );
  XOR U10070 ( .A(n10488), .B(n10489), .Z(n9567) );
  NOR U10071 ( .A(n5577), .B(n5575), .Z(n10449) );
  XOR U10072 ( .A(n10490), .B(n1694), .Z(n5575) );
  XNOR U10073 ( .A(n8719), .B(n6206), .Z(n1694) );
  XNOR U10074 ( .A(n10491), .B(n10492), .Z(n6206) );
  XOR U10075 ( .A(n5341), .B(n3589), .Z(n10492) );
  XOR U10076 ( .A(n10493), .B(n10494), .Z(n3589) );
  ANDN U10077 ( .B(n7827), .A(n10495), .Z(n10493) );
  IV U10078 ( .A(n10496), .Z(n7827) );
  XOR U10079 ( .A(n10497), .B(n10498), .Z(n5341) );
  ANDN U10080 ( .B(n10499), .A(n7817), .Z(n10497) );
  XNOR U10081 ( .A(n10500), .B(n10501), .Z(n10491) );
  XOR U10082 ( .A(n2055), .B(n5261), .Z(n10501) );
  XNOR U10083 ( .A(n10502), .B(n10503), .Z(n5261) );
  ANDN U10084 ( .B(n10504), .A(n10505), .Z(n10502) );
  XNOR U10085 ( .A(n10506), .B(n10507), .Z(n2055) );
  ANDN U10086 ( .B(n8844), .A(n10508), .Z(n10506) );
  XOR U10087 ( .A(n10509), .B(n10510), .Z(n8719) );
  XNOR U10088 ( .A(n5020), .B(n7726), .Z(n10510) );
  XOR U10089 ( .A(n10511), .B(n7732), .Z(n7726) );
  XNOR U10090 ( .A(n10512), .B(n7737), .Z(n5020) );
  ANDN U10091 ( .B(n7736), .A(n10324), .Z(n10512) );
  IV U10092 ( .A(n10513), .Z(n7736) );
  XNOR U10093 ( .A(n2394), .B(n10514), .Z(n10509) );
  XNOR U10094 ( .A(n3417), .B(n3965), .Z(n10514) );
  XOR U10095 ( .A(n10515), .B(n7742), .Z(n3965) );
  ANDN U10096 ( .B(n7743), .A(n10315), .Z(n10515) );
  XNOR U10097 ( .A(n10516), .B(n8781), .Z(n3417) );
  XNOR U10098 ( .A(n10517), .B(n10518), .Z(n2394) );
  AND U10099 ( .A(n7747), .B(n10519), .Z(n10517) );
  XOR U10100 ( .A(n9467), .B(n2021), .Z(n5577) );
  XNOR U10101 ( .A(n9318), .B(n8290), .Z(n2021) );
  XNOR U10102 ( .A(n10520), .B(n10521), .Z(n8290) );
  XOR U10103 ( .A(n5374), .B(n3826), .Z(n10521) );
  XOR U10104 ( .A(n10522), .B(n10523), .Z(n3826) );
  AND U10105 ( .A(n10524), .B(n9733), .Z(n10522) );
  XNOR U10106 ( .A(n10525), .B(n9632), .Z(n5374) );
  AND U10107 ( .A(n10526), .B(n10527), .Z(n10525) );
  XOR U10108 ( .A(n6170), .B(n10528), .Z(n10520) );
  XNOR U10109 ( .A(n2251), .B(n4943), .Z(n10528) );
  XNOR U10110 ( .A(n10529), .B(n9636), .Z(n4943) );
  AND U10111 ( .A(n9728), .B(n10530), .Z(n10529) );
  XNOR U10112 ( .A(n10531), .B(n10532), .Z(n2251) );
  AND U10113 ( .A(n9737), .B(n10533), .Z(n10531) );
  XNOR U10114 ( .A(n10534), .B(n9642), .Z(n6170) );
  AND U10115 ( .A(n9643), .B(n9725), .Z(n10534) );
  XOR U10116 ( .A(n10535), .B(n10536), .Z(n9318) );
  XNOR U10117 ( .A(n1964), .B(n9610), .Z(n10536) );
  XOR U10118 ( .A(n10537), .B(n10421), .Z(n9610) );
  IV U10119 ( .A(n10437), .Z(n10421) );
  XOR U10120 ( .A(n10538), .B(n9274), .Z(n10437) );
  ANDN U10121 ( .B(n9460), .A(n9461), .Z(n10537) );
  XNOR U10122 ( .A(n10539), .B(n10540), .Z(n9461) );
  XOR U10123 ( .A(n10541), .B(n10172), .Z(n9460) );
  XOR U10124 ( .A(n10542), .B(n9615), .Z(n1964) );
  XNOR U10125 ( .A(n9605), .B(n10543), .Z(n9615) );
  ANDN U10126 ( .B(n9472), .A(n9470), .Z(n10542) );
  XNOR U10127 ( .A(n10544), .B(n10545), .Z(n9470) );
  XNOR U10128 ( .A(n10546), .B(n10382), .Z(n9472) );
  XOR U10129 ( .A(n3715), .B(n10547), .Z(n10535) );
  XNOR U10130 ( .A(n5068), .B(n4180), .Z(n10547) );
  XOR U10131 ( .A(n10548), .B(n10446), .Z(n4180) );
  IV U10132 ( .A(n9623), .Z(n10446) );
  XNOR U10133 ( .A(n10549), .B(n9782), .Z(n9623) );
  ANDN U10134 ( .B(n9624), .A(n10343), .Z(n10548) );
  XNOR U10135 ( .A(n10550), .B(n9618), .Z(n5068) );
  XNOR U10136 ( .A(n10551), .B(n9900), .Z(n9618) );
  AND U10137 ( .A(n9464), .B(n10350), .Z(n10550) );
  IV U10138 ( .A(n9465), .Z(n10350) );
  XOR U10139 ( .A(n10552), .B(n10553), .Z(n9465) );
  XOR U10140 ( .A(n10554), .B(n9370), .Z(n9464) );
  XOR U10141 ( .A(n10555), .B(n10427), .Z(n3715) );
  IV U10142 ( .A(n9627), .Z(n10427) );
  XNOR U10143 ( .A(n10556), .B(n10019), .Z(n9627) );
  ANDN U10144 ( .B(n9475), .A(n9474), .Z(n10555) );
  XOR U10145 ( .A(n10557), .B(n10558), .Z(n9474) );
  XOR U10146 ( .A(n10559), .B(n10560), .Z(n9475) );
  XOR U10147 ( .A(n10561), .B(n9624), .Z(n9467) );
  XOR U10148 ( .A(n10562), .B(n10563), .Z(n9624) );
  AND U10149 ( .A(n10343), .B(n10445), .Z(n10561) );
  IV U10150 ( .A(n10344), .Z(n10445) );
  XOR U10151 ( .A(n10564), .B(n10565), .Z(n10344) );
  XNOR U10152 ( .A(n10566), .B(n9798), .Z(n10343) );
  XOR U10153 ( .A(n10567), .B(n6079), .Z(out[1018]) );
  XOR U10154 ( .A(n10568), .B(n2645), .Z(n6079) );
  XNOR U10155 ( .A(n5961), .B(n8540), .Z(n2645) );
  XNOR U10156 ( .A(n10569), .B(n10570), .Z(n8540) );
  XOR U10157 ( .A(n5556), .B(n5357), .Z(n10570) );
  XNOR U10158 ( .A(n10571), .B(n6919), .Z(n5357) );
  XOR U10159 ( .A(n10572), .B(n9692), .Z(n6919) );
  ANDN U10160 ( .B(n10476), .A(n6918), .Z(n10571) );
  XOR U10161 ( .A(n10573), .B(n9306), .Z(n5556) );
  IV U10162 ( .A(n6929), .Z(n9306) );
  XOR U10163 ( .A(n10574), .B(n10296), .Z(n6929) );
  NOR U10164 ( .A(n10483), .B(n6928), .Z(n10573) );
  XOR U10165 ( .A(n6912), .B(n10575), .Z(n10569) );
  XNOR U10166 ( .A(n2208), .B(n3336), .Z(n10575) );
  XNOR U10167 ( .A(n10576), .B(n6932), .Z(n3336) );
  XNOR U10168 ( .A(n10577), .B(n10578), .Z(n6932) );
  AND U10169 ( .A(n10468), .B(n10579), .Z(n10576) );
  XNOR U10170 ( .A(n10580), .B(n6923), .Z(n2208) );
  XOR U10171 ( .A(n10581), .B(n10455), .Z(n6923) );
  ANDN U10172 ( .B(n10480), .A(n6922), .Z(n10580) );
  XNOR U10173 ( .A(n10582), .B(n9298), .Z(n6912) );
  XNOR U10174 ( .A(n10583), .B(n10584), .Z(n9298) );
  AND U10175 ( .A(n10471), .B(n10585), .Z(n10582) );
  XOR U10176 ( .A(n10586), .B(n10587), .Z(n5961) );
  XOR U10177 ( .A(n5191), .B(n1867), .Z(n10587) );
  XNOR U10178 ( .A(n10588), .B(n8027), .Z(n1867) );
  AND U10179 ( .A(n6955), .B(n10396), .Z(n10588) );
  XOR U10180 ( .A(n10589), .B(n10590), .Z(n10396) );
  XNOR U10181 ( .A(n10591), .B(n9678), .Z(n6955) );
  IV U10182 ( .A(n10436), .Z(n9678) );
  XNOR U10183 ( .A(n10592), .B(n8036), .Z(n5191) );
  ANDN U10184 ( .B(n10393), .A(n8035), .Z(n10592) );
  XNOR U10185 ( .A(n10593), .B(n10594), .Z(n8035) );
  XOR U10186 ( .A(n10595), .B(n10233), .Z(n10393) );
  XNOR U10187 ( .A(n3608), .B(n10596), .Z(n10586) );
  XOR U10188 ( .A(n8020), .B(n4109), .Z(n10596) );
  XNOR U10189 ( .A(n10597), .B(n8039), .Z(n4109) );
  ANDN U10190 ( .B(n8038), .A(n6941), .Z(n10597) );
  XNOR U10191 ( .A(n10598), .B(n10599), .Z(n6941) );
  XOR U10192 ( .A(n9682), .B(n10600), .Z(n8038) );
  XOR U10193 ( .A(n10601), .B(n8031), .Z(n8020) );
  AND U10194 ( .A(n6945), .B(n8032), .Z(n10601) );
  XOR U10195 ( .A(n10602), .B(n10603), .Z(n8032) );
  XNOR U10196 ( .A(n10604), .B(n10265), .Z(n6945) );
  XNOR U10197 ( .A(n10605), .B(n10606), .Z(n3608) );
  ANDN U10198 ( .B(n6951), .A(n10401), .Z(n10605) );
  XOR U10199 ( .A(n10607), .B(n10096), .Z(n6951) );
  NOR U10200 ( .A(n5581), .B(n5579), .Z(n10567) );
  XOR U10201 ( .A(n10608), .B(n1698), .Z(n5579) );
  XNOR U10202 ( .A(n8778), .B(n6210), .Z(n1698) );
  XNOR U10203 ( .A(n10609), .B(n10610), .Z(n6210) );
  XOR U10204 ( .A(n5345), .B(n3593), .Z(n10610) );
  XOR U10205 ( .A(n10611), .B(n10612), .Z(n3593) );
  NOR U10206 ( .A(n7875), .B(n10613), .Z(n10611) );
  XOR U10207 ( .A(n10614), .B(n10615), .Z(n5345) );
  AND U10208 ( .A(n7865), .B(n10616), .Z(n10614) );
  XNOR U10209 ( .A(n10617), .B(n10618), .Z(n10609) );
  XNOR U10210 ( .A(n2058), .B(n5314), .Z(n10618) );
  XOR U10211 ( .A(n10619), .B(n10620), .Z(n5314) );
  ANDN U10212 ( .B(n7869), .A(n10621), .Z(n10619) );
  XNOR U10213 ( .A(n10622), .B(n10623), .Z(n2058) );
  AND U10214 ( .A(n10624), .B(n8908), .Z(n10622) );
  XOR U10215 ( .A(n10625), .B(n10626), .Z(n8778) );
  XNOR U10216 ( .A(n3423), .B(n5023), .Z(n10626) );
  XNOR U10217 ( .A(n10627), .B(n7823), .Z(n5023) );
  XOR U10218 ( .A(n10628), .B(n8845), .Z(n3423) );
  AND U10219 ( .A(n10507), .B(n10629), .Z(n10628) );
  XOR U10220 ( .A(n3968), .B(n10630), .Z(n10625) );
  XOR U10221 ( .A(n7812), .B(n2404), .Z(n10630) );
  XOR U10222 ( .A(n10631), .B(n7832), .Z(n2404) );
  AND U10223 ( .A(n7833), .B(n10632), .Z(n10631) );
  XOR U10224 ( .A(n10633), .B(n7818), .Z(n7812) );
  AND U10225 ( .A(n7819), .B(n10634), .Z(n10633) );
  XOR U10226 ( .A(n10635), .B(n7828), .Z(n3968) );
  AND U10227 ( .A(n10494), .B(n7829), .Z(n10635) );
  XOR U10228 ( .A(n9638), .B(n2024), .Z(n5581) );
  XNOR U10229 ( .A(n10422), .B(n8561), .Z(n2024) );
  XNOR U10230 ( .A(n10636), .B(n10637), .Z(n8561) );
  XOR U10231 ( .A(n5378), .B(n3832), .Z(n10637) );
  XOR U10232 ( .A(n10638), .B(n10639), .Z(n3832) );
  ANDN U10233 ( .B(n7316), .A(n7317), .Z(n10638) );
  XNOR U10234 ( .A(n9097), .B(n10640), .Z(n7317) );
  XNOR U10235 ( .A(n10641), .B(n9743), .Z(n5378) );
  ANDN U10236 ( .B(n7312), .A(n7313), .Z(n10641) );
  XNOR U10237 ( .A(n10142), .B(n10642), .Z(n7313) );
  XOR U10238 ( .A(n10643), .B(n9906), .Z(n7312) );
  XNOR U10239 ( .A(n6175), .B(n10644), .Z(n10636) );
  XOR U10240 ( .A(n2258), .B(n4978), .Z(n10644) );
  XNOR U10241 ( .A(n10645), .B(n9746), .Z(n4978) );
  AND U10242 ( .A(n8342), .B(n8341), .Z(n10645) );
  XNOR U10243 ( .A(n10646), .B(n9768), .Z(n8341) );
  XOR U10244 ( .A(n9354), .B(n10647), .Z(n8342) );
  XOR U10245 ( .A(n10648), .B(n9754), .Z(n2258) );
  ANDN U10246 ( .B(n8563), .A(n8564), .Z(n10648) );
  XNOR U10247 ( .A(n10649), .B(n10650), .Z(n8564) );
  XNOR U10248 ( .A(n10651), .B(n10652), .Z(n8563) );
  XNOR U10249 ( .A(n10653), .B(n9751), .Z(n6175) );
  ANDN U10250 ( .B(n7308), .A(n7306), .Z(n10653) );
  XOR U10251 ( .A(n10654), .B(n9176), .Z(n7306) );
  XOR U10252 ( .A(n10655), .B(n9694), .Z(n7308) );
  XOR U10253 ( .A(n10656), .B(n10657), .Z(n10422) );
  XOR U10254 ( .A(n1659), .B(n9721), .Z(n10657) );
  XOR U10255 ( .A(n10658), .B(n10659), .Z(n9721) );
  NOR U10256 ( .A(n9632), .B(n9631), .Z(n10658) );
  XNOR U10257 ( .A(n10660), .B(n10661), .Z(n9632) );
  XNOR U10258 ( .A(n10662), .B(n9726), .Z(n1659) );
  ANDN U10259 ( .B(n9641), .A(n9642), .Z(n10662) );
  XNOR U10260 ( .A(n10557), .B(n10663), .Z(n9642) );
  XNOR U10261 ( .A(n10664), .B(n10665), .Z(n9641) );
  XOR U10262 ( .A(n3719), .B(n10666), .Z(n10656) );
  XOR U10263 ( .A(n5070), .B(n4184), .Z(n10666) );
  XOR U10264 ( .A(n10667), .B(n10668), .Z(n4184) );
  NOR U10265 ( .A(n9734), .B(n10523), .Z(n10667) );
  XOR U10266 ( .A(n10669), .B(n10670), .Z(n5070) );
  NOR U10267 ( .A(n9636), .B(n9635), .Z(n10669) );
  XOR U10268 ( .A(n9086), .B(n10671), .Z(n9635) );
  IV U10269 ( .A(n10651), .Z(n9086) );
  XOR U10270 ( .A(n10672), .B(n10673), .Z(n10651) );
  XOR U10271 ( .A(n10674), .B(n10675), .Z(n9636) );
  XOR U10272 ( .A(n10676), .B(n10677), .Z(n3719) );
  AND U10273 ( .A(n9645), .B(n10532), .Z(n10676) );
  IV U10274 ( .A(n9647), .Z(n10532) );
  XOR U10275 ( .A(n10678), .B(n10679), .Z(n9647) );
  XOR U10276 ( .A(n10680), .B(n10681), .Z(n9645) );
  XNOR U10277 ( .A(n10682), .B(n9734), .Z(n9638) );
  XNOR U10278 ( .A(n10559), .B(n10683), .Z(n9734) );
  ANDN U10279 ( .B(n10523), .A(n10524), .Z(n10682) );
  XNOR U10280 ( .A(n10684), .B(n9924), .Z(n10523) );
  XOR U10281 ( .A(n10685), .B(n6084), .Z(out[1017]) );
  IV U10282 ( .A(n6544), .Z(n6084) );
  XOR U10283 ( .A(n8024), .B(n2652), .Z(n6544) );
  XNOR U10284 ( .A(n5966), .B(n9292), .Z(n2652) );
  XNOR U10285 ( .A(n10686), .B(n10687), .Z(n9292) );
  XNOR U10286 ( .A(n5601), .B(n5360), .Z(n10687) );
  XNOR U10287 ( .A(n10688), .B(n6943), .Z(n5360) );
  XNOR U10288 ( .A(n10689), .B(n9800), .Z(n6943) );
  ANDN U10289 ( .B(n8039), .A(n6942), .Z(n10688) );
  XNOR U10290 ( .A(n10690), .B(n10691), .Z(n6942) );
  XNOR U10291 ( .A(n10692), .B(n10693), .Z(n8039) );
  XNOR U10292 ( .A(n10694), .B(n6953), .Z(n5601) );
  XNOR U10293 ( .A(n10695), .B(n10696), .Z(n6953) );
  ANDN U10294 ( .B(n10606), .A(n6952), .Z(n10694) );
  XOR U10295 ( .A(n6936), .B(n10697), .Z(n10686) );
  XOR U10296 ( .A(n2215), .B(n3340), .Z(n10697) );
  XOR U10297 ( .A(n10698), .B(n10397), .Z(n3340) );
  XNOR U10298 ( .A(n10699), .B(n9676), .Z(n10397) );
  AND U10299 ( .A(n6957), .B(n8027), .Z(n10698) );
  XOR U10300 ( .A(n10700), .B(n10701), .Z(n8027) );
  XNOR U10301 ( .A(n10702), .B(n10160), .Z(n6957) );
  XNOR U10302 ( .A(n10703), .B(n6946), .Z(n2215) );
  XNOR U10303 ( .A(n10704), .B(n10705), .Z(n6946) );
  AND U10304 ( .A(n8031), .B(n8030), .Z(n10703) );
  IV U10305 ( .A(n6947), .Z(n8030) );
  XOR U10306 ( .A(n10706), .B(n10707), .Z(n6947) );
  XOR U10307 ( .A(n10708), .B(n10709), .Z(n8031) );
  XNOR U10308 ( .A(n10710), .B(n10394), .Z(n6936) );
  XNOR U10309 ( .A(n10711), .B(n10712), .Z(n10394) );
  AND U10310 ( .A(n8034), .B(n8036), .Z(n10710) );
  XNOR U10311 ( .A(n10713), .B(n10714), .Z(n8036) );
  XNOR U10312 ( .A(n10715), .B(n10716), .Z(n8034) );
  XOR U10313 ( .A(n10717), .B(n10718), .Z(n5966) );
  XOR U10314 ( .A(n5194), .B(n1871), .Z(n10718) );
  XOR U10315 ( .A(n10719), .B(n8074), .Z(n1871) );
  NOR U10316 ( .A(n6978), .B(n8075), .Z(n10719) );
  XNOR U10317 ( .A(n10720), .B(n8082), .Z(n5194) );
  ANDN U10318 ( .B(n8083), .A(n10721), .Z(n10720) );
  XOR U10319 ( .A(n3612), .B(n10722), .Z(n10717) );
  XNOR U10320 ( .A(n8069), .B(n4112), .Z(n10722) );
  XOR U10321 ( .A(n10723), .B(n8086), .Z(n4112) );
  ANDN U10322 ( .B(n6964), .A(n8085), .Z(n10723) );
  XNOR U10323 ( .A(n10724), .B(n8078), .Z(n8069) );
  ANDN U10324 ( .B(n8079), .A(n6968), .Z(n10724) );
  XNOR U10325 ( .A(n10725), .B(n10726), .Z(n3612) );
  ANDN U10326 ( .B(n6974), .A(n10727), .Z(n10725) );
  XOR U10327 ( .A(n10728), .B(n6952), .Z(n8024) );
  XOR U10328 ( .A(n10729), .B(n10256), .Z(n6952) );
  ANDN U10329 ( .B(n10401), .A(n10606), .Z(n10728) );
  XNOR U10330 ( .A(n10730), .B(n10731), .Z(n10606) );
  XOR U10331 ( .A(n10732), .B(n9782), .Z(n10401) );
  ANDN U10332 ( .B(n5585), .A(n5583), .Z(n10685) );
  XOR U10333 ( .A(n10733), .B(n1703), .Z(n5583) );
  XNOR U10334 ( .A(n8841), .B(n6218), .Z(n1703) );
  XNOR U10335 ( .A(n10734), .B(n10735), .Z(n6218) );
  XOR U10336 ( .A(n5351), .B(n3596), .Z(n10735) );
  XOR U10337 ( .A(n10736), .B(n10737), .Z(n3596) );
  XOR U10338 ( .A(n10739), .B(n10740), .Z(n5351) );
  NOR U10339 ( .A(n7974), .B(n10741), .Z(n10739) );
  XNOR U10340 ( .A(n10742), .B(n10743), .Z(n10734) );
  XNOR U10341 ( .A(n2061), .B(n5363), .Z(n10743) );
  XOR U10342 ( .A(n10744), .B(n10745), .Z(n5363) );
  XNOR U10343 ( .A(n10747), .B(n10748), .Z(n2061) );
  ANDN U10344 ( .B(n8971), .A(n10749), .Z(n10747) );
  IV U10345 ( .A(n10750), .Z(n8971) );
  XOR U10346 ( .A(n10751), .B(n10752), .Z(n8841) );
  XOR U10347 ( .A(n3426), .B(n5027), .Z(n10752) );
  XNOR U10348 ( .A(n10753), .B(n7871), .Z(n5027) );
  AND U10349 ( .A(n10620), .B(n10754), .Z(n10753) );
  XOR U10350 ( .A(n10755), .B(n8909), .Z(n3426) );
  AND U10351 ( .A(n10623), .B(n10756), .Z(n10755) );
  XNOR U10352 ( .A(n3984), .B(n10757), .Z(n10751) );
  XOR U10353 ( .A(n7860), .B(n2409), .Z(n10757) );
  XOR U10354 ( .A(n10758), .B(n7880), .Z(n2409) );
  AND U10355 ( .A(n10759), .B(n7881), .Z(n10758) );
  XOR U10356 ( .A(n10760), .B(n7866), .Z(n7860) );
  XOR U10357 ( .A(n10761), .B(n7876), .Z(n3984) );
  ANDN U10358 ( .B(n10762), .A(n7877), .Z(n10761) );
  XNOR U10359 ( .A(n9747), .B(n2031), .Z(n5585) );
  XNOR U10360 ( .A(n10763), .B(n9312), .Z(n2031) );
  XNOR U10361 ( .A(n10764), .B(n10765), .Z(n9312) );
  XNOR U10362 ( .A(n5385), .B(n3838), .Z(n10765) );
  XNOR U10363 ( .A(n10766), .B(n10767), .Z(n3838) );
  AND U10364 ( .A(n7395), .B(n7393), .Z(n10766) );
  IV U10365 ( .A(n10768), .Z(n7393) );
  XOR U10366 ( .A(n9673), .B(n10769), .Z(n7395) );
  XOR U10367 ( .A(n10770), .B(n9839), .Z(n5385) );
  ANDN U10368 ( .B(n7389), .A(n7390), .Z(n10770) );
  XNOR U10369 ( .A(n10771), .B(n10286), .Z(n7390) );
  XNOR U10370 ( .A(n10772), .B(n10773), .Z(n7389) );
  XOR U10371 ( .A(n6180), .B(n10774), .Z(n10764) );
  XOR U10372 ( .A(n2265), .B(n5015), .Z(n10774) );
  XNOR U10373 ( .A(n10775), .B(n9842), .Z(n5015) );
  AND U10374 ( .A(n8397), .B(n9843), .Z(n10775) );
  XOR U10375 ( .A(n9894), .B(n10776), .Z(n9843) );
  XNOR U10376 ( .A(n10777), .B(n9483), .Z(n8397) );
  XOR U10377 ( .A(n10778), .B(n9852), .Z(n2265) );
  ANDN U10378 ( .B(n9314), .A(n9315), .Z(n10778) );
  XOR U10379 ( .A(n9684), .B(n10779), .Z(n9315) );
  XNOR U10380 ( .A(n9576), .B(n10780), .Z(n9314) );
  XNOR U10381 ( .A(n10781), .B(n9848), .Z(n6180) );
  AND U10382 ( .A(n7384), .B(n9849), .Z(n10781) );
  XNOR U10383 ( .A(n10782), .B(n10783), .Z(n9849) );
  XNOR U10384 ( .A(n10784), .B(n10785), .Z(n7384) );
  XNOR U10385 ( .A(n10786), .B(n9834), .Z(n9747) );
  XNOR U10386 ( .A(n10787), .B(n10788), .Z(n7316) );
  XOR U10387 ( .A(n10789), .B(n6089), .Z(out[1016]) );
  IV U10388 ( .A(n6571), .Z(n6089) );
  XOR U10389 ( .A(n8072), .B(n2659), .Z(n6571) );
  XNOR U10390 ( .A(n5971), .B(n10389), .Z(n2659) );
  XNOR U10391 ( .A(n10790), .B(n10791), .Z(n10389) );
  XOR U10392 ( .A(n5645), .B(n5371), .Z(n10791) );
  XNOR U10393 ( .A(n10792), .B(n6966), .Z(n5371) );
  NOR U10394 ( .A(n6965), .B(n8086), .Z(n10792) );
  XOR U10395 ( .A(n10793), .B(n10794), .Z(n8086) );
  XOR U10396 ( .A(n9083), .B(n10795), .Z(n6965) );
  XOR U10397 ( .A(n10796), .B(n10797), .Z(n5645) );
  ANDN U10398 ( .B(n10726), .A(n6975), .Z(n10796) );
  XOR U10399 ( .A(n6959), .B(n10798), .Z(n10790) );
  XOR U10400 ( .A(n2222), .B(n3344), .Z(n10798) );
  XOR U10401 ( .A(n10799), .B(n10800), .Z(n3344) );
  ANDN U10402 ( .B(n6980), .A(n8074), .Z(n10799) );
  XOR U10403 ( .A(n9480), .B(n10801), .Z(n8074) );
  XNOR U10404 ( .A(n10802), .B(n10803), .Z(n6980) );
  XOR U10405 ( .A(n10804), .B(n6970), .Z(n2222) );
  ANDN U10406 ( .B(n8078), .A(n6969), .Z(n10804) );
  XNOR U10407 ( .A(n10805), .B(n10806), .Z(n6969) );
  XNOR U10408 ( .A(n10807), .B(n10808), .Z(n8078) );
  XNOR U10409 ( .A(n10809), .B(n10810), .Z(n6959) );
  AND U10410 ( .A(n8082), .B(n10811), .Z(n10809) );
  XNOR U10411 ( .A(n10812), .B(n10254), .Z(n8082) );
  XOR U10412 ( .A(n10813), .B(n10814), .Z(n5971) );
  XOR U10413 ( .A(n5200), .B(n1875), .Z(n10814) );
  XNOR U10414 ( .A(n10815), .B(n8155), .Z(n1875) );
  ANDN U10415 ( .B(n8092), .A(n7004), .Z(n10815) );
  XOR U10416 ( .A(n10816), .B(n10817), .Z(n7004) );
  XOR U10417 ( .A(n10819), .B(n8160), .Z(n5200) );
  IV U10418 ( .A(n10820), .Z(n8160) );
  ANDN U10419 ( .B(n8090), .A(n7000), .Z(n10819) );
  XOR U10420 ( .A(n9605), .B(n10821), .Z(n7000) );
  XNOR U10421 ( .A(n10822), .B(n10823), .Z(n8090) );
  XOR U10422 ( .A(n3616), .B(n10824), .Z(n10813) );
  XOR U10423 ( .A(n8149), .B(n4116), .Z(n10824) );
  XNOR U10424 ( .A(n10825), .B(n8162), .Z(n4116) );
  AND U10425 ( .A(n6987), .B(n8099), .Z(n10825) );
  XOR U10426 ( .A(n10826), .B(n10203), .Z(n8099) );
  XNOR U10427 ( .A(n10827), .B(n10828), .Z(n6987) );
  XNOR U10428 ( .A(n10829), .B(n8158), .Z(n8149) );
  XNOR U10429 ( .A(n10830), .B(n10831), .Z(n6991) );
  XOR U10430 ( .A(n10118), .B(n10832), .Z(n8095) );
  XNOR U10431 ( .A(n10833), .B(n10834), .Z(n3616) );
  ANDN U10432 ( .B(n8097), .A(n6996), .Z(n10833) );
  XNOR U10433 ( .A(n10835), .B(n10439), .Z(n6996) );
  XOR U10434 ( .A(n10836), .B(n6975), .Z(n8072) );
  XOR U10435 ( .A(n10837), .B(n10386), .Z(n6975) );
  ANDN U10436 ( .B(n10727), .A(n10726), .Z(n10836) );
  XOR U10437 ( .A(n10838), .B(n10839), .Z(n10726) );
  ANDN U10438 ( .B(n5589), .A(n5587), .Z(n10789) );
  XOR U10439 ( .A(n10840), .B(n1707), .Z(n5587) );
  XNOR U10440 ( .A(n8906), .B(n6222), .Z(n1707) );
  XNOR U10441 ( .A(n10841), .B(n10842), .Z(n6222) );
  XNOR U10442 ( .A(n5355), .B(n3602), .Z(n10842) );
  XOR U10443 ( .A(n10843), .B(n10844), .Z(n3602) );
  ANDN U10444 ( .B(n8055), .A(n10845), .Z(n10843) );
  IV U10445 ( .A(n10846), .Z(n8055) );
  XNOR U10446 ( .A(n10847), .B(n10848), .Z(n5355) );
  AND U10447 ( .A(n8045), .B(n10849), .Z(n10847) );
  XNOR U10448 ( .A(n10850), .B(n10851), .Z(n10841) );
  XOR U10449 ( .A(n2068), .B(n5415), .Z(n10851) );
  XNOR U10450 ( .A(n10852), .B(n10853), .Z(n5415) );
  ANDN U10451 ( .B(n10854), .A(n10855), .Z(n10852) );
  XNOR U10452 ( .A(n10856), .B(n10857), .Z(n2068) );
  XOR U10453 ( .A(n10859), .B(n10860), .Z(n8906) );
  XNOR U10454 ( .A(n3429), .B(n5030), .Z(n10860) );
  XNOR U10455 ( .A(n10861), .B(n7980), .Z(n5030) );
  AND U10456 ( .A(n7979), .B(n10745), .Z(n10861) );
  XNOR U10457 ( .A(n10862), .B(n8972), .Z(n3429) );
  AND U10458 ( .A(n8973), .B(n10748), .Z(n10862) );
  XOR U10459 ( .A(n4017), .B(n10863), .Z(n10859) );
  XNOR U10460 ( .A(n7969), .B(n2418), .Z(n10863) );
  XNOR U10461 ( .A(n10864), .B(n7990), .Z(n2418) );
  AND U10462 ( .A(n7989), .B(n10865), .Z(n10864) );
  XNOR U10463 ( .A(n10866), .B(n7976), .Z(n7969) );
  XOR U10464 ( .A(n10867), .B(n7985), .Z(n4017) );
  IV U10465 ( .A(n10868), .Z(n7985) );
  AND U10466 ( .A(n7986), .B(n10869), .Z(n10867) );
  XNOR U10467 ( .A(n9844), .B(n2034), .Z(n5589) );
  XNOR U10468 ( .A(n7301), .B(n10404), .Z(n2034) );
  XNOR U10469 ( .A(n10870), .B(n10871), .Z(n10404) );
  XNOR U10470 ( .A(n5388), .B(n3844), .Z(n10871) );
  XOR U10471 ( .A(n10872), .B(n10873), .Z(n3844) );
  AND U10472 ( .A(n7437), .B(n7439), .Z(n10872) );
  XNOR U10473 ( .A(n10874), .B(n10875), .Z(n7439) );
  XNOR U10474 ( .A(n10876), .B(n9874), .Z(n5388) );
  AND U10475 ( .A(n7433), .B(n7435), .Z(n10876) );
  XNOR U10476 ( .A(n10877), .B(n9505), .Z(n7435) );
  XNOR U10477 ( .A(n10878), .B(n10030), .Z(n7433) );
  XOR U10478 ( .A(n6184), .B(n10879), .Z(n10870) );
  XNOR U10479 ( .A(n2272), .B(n5051), .Z(n10879) );
  XNOR U10480 ( .A(n10880), .B(n9877), .Z(n5051) );
  AND U10481 ( .A(n8471), .B(n9878), .Z(n10880) );
  XOR U10482 ( .A(n10377), .B(n10881), .Z(n9878) );
  XNOR U10483 ( .A(n9552), .B(n10882), .Z(n8471) );
  XOR U10484 ( .A(n10883), .B(n10884), .Z(n2272) );
  AND U10485 ( .A(n9887), .B(n9961), .Z(n10883) );
  XNOR U10486 ( .A(n10885), .B(n9077), .Z(n9961) );
  XOR U10487 ( .A(n10886), .B(n9687), .Z(n9887) );
  XNOR U10488 ( .A(n10887), .B(n9883), .Z(n6184) );
  AND U10489 ( .A(n7427), .B(n7429), .Z(n10887) );
  XOR U10490 ( .A(n10888), .B(n9924), .Z(n7429) );
  XNOR U10491 ( .A(n10889), .B(n9360), .Z(n7427) );
  XOR U10492 ( .A(n10890), .B(n10891), .Z(n7301) );
  XNOR U10493 ( .A(n1671), .B(n9859), .Z(n10891) );
  XNOR U10494 ( .A(n10892), .B(n7391), .Z(n9859) );
  XNOR U10495 ( .A(n9378), .B(n10893), .Z(n7391) );
  IV U10496 ( .A(n10220), .Z(n9378) );
  AND U10497 ( .A(n9838), .B(n9839), .Z(n10892) );
  XNOR U10498 ( .A(n10894), .B(n10448), .Z(n9839) );
  XOR U10499 ( .A(n10895), .B(n10896), .Z(n9838) );
  XNOR U10500 ( .A(n10897), .B(n7385), .Z(n1671) );
  XOR U10501 ( .A(n10898), .B(n10899), .Z(n7385) );
  ANDN U10502 ( .B(n9848), .A(n9847), .Z(n10897) );
  XNOR U10503 ( .A(n10900), .B(n10901), .Z(n9847) );
  XNOR U10504 ( .A(n10902), .B(n10903), .Z(n9848) );
  XNOR U10505 ( .A(n3730), .B(n10904), .Z(n10890) );
  XNOR U10506 ( .A(n5074), .B(n4194), .Z(n10904) );
  XOR U10507 ( .A(n10905), .B(n7394), .Z(n4194) );
  IV U10508 ( .A(n9869), .Z(n7394) );
  XOR U10509 ( .A(n10906), .B(n10030), .Z(n9869) );
  NOR U10510 ( .A(n9868), .B(n10767), .Z(n10905) );
  IV U10511 ( .A(n10907), .Z(n9868) );
  XNOR U10512 ( .A(n10908), .B(n8398), .Z(n5074) );
  XNOR U10513 ( .A(n10909), .B(n10910), .Z(n8398) );
  ANDN U10514 ( .B(n9841), .A(n9842), .Z(n10908) );
  XNOR U10515 ( .A(n10911), .B(n10912), .Z(n9842) );
  XOR U10516 ( .A(n10913), .B(n9687), .Z(n9841) );
  XNOR U10517 ( .A(n10914), .B(n9316), .Z(n3730) );
  XOR U10518 ( .A(n10915), .B(n10916), .Z(n9316) );
  AND U10519 ( .A(n9851), .B(n9852), .Z(n10914) );
  XNOR U10520 ( .A(n10917), .B(n10918), .Z(n9852) );
  XOR U10521 ( .A(n10921), .B(n10907), .Z(n9844) );
  XOR U10522 ( .A(n10922), .B(n10923), .Z(n10907) );
  AND U10523 ( .A(n10767), .B(n10768), .Z(n10921) );
  XNOR U10524 ( .A(n10924), .B(n10925), .Z(n10768) );
  XOR U10525 ( .A(n10926), .B(n10043), .Z(n10767) );
  XOR U10526 ( .A(n10927), .B(n6094), .Z(out[1015]) );
  IV U10527 ( .A(n6604), .Z(n6094) );
  XOR U10528 ( .A(n8152), .B(n2666), .Z(n6604) );
  XNOR U10529 ( .A(n5976), .B(n10928), .Z(n2666) );
  XOR U10530 ( .A(n10929), .B(n10930), .Z(n5976) );
  XNOR U10531 ( .A(n5203), .B(n1879), .Z(n10930) );
  XNOR U10532 ( .A(n10931), .B(n8222), .Z(n1879) );
  AND U10533 ( .A(n8168), .B(n8169), .Z(n10931) );
  XOR U10534 ( .A(n10932), .B(n10933), .Z(n8169) );
  XNOR U10535 ( .A(n10539), .B(n10934), .Z(n8168) );
  XNOR U10536 ( .A(n10935), .B(n8227), .Z(n5203) );
  ANDN U10537 ( .B(n8228), .A(n7058), .Z(n10935) );
  XOR U10538 ( .A(n10936), .B(n9716), .Z(n7058) );
  XNOR U10539 ( .A(n10937), .B(n10938), .Z(n8228) );
  XOR U10540 ( .A(n3624), .B(n10939), .Z(n10929) );
  XOR U10541 ( .A(n8203), .B(n4119), .Z(n10939) );
  XOR U10542 ( .A(n10940), .B(n8230), .Z(n4119) );
  NOR U10543 ( .A(n7045), .B(n8176), .Z(n10940) );
  XOR U10544 ( .A(n10941), .B(n9112), .Z(n8176) );
  XNOR U10545 ( .A(n10942), .B(n10943), .Z(n7045) );
  XOR U10546 ( .A(n10944), .B(n8225), .Z(n8203) );
  ANDN U10547 ( .B(n8172), .A(n7049), .Z(n10944) );
  XOR U10548 ( .A(n10945), .B(n10691), .Z(n7049) );
  XOR U10549 ( .A(n10262), .B(n10946), .Z(n8172) );
  XNOR U10550 ( .A(n10947), .B(n10948), .Z(n3624) );
  ANDN U10551 ( .B(n10949), .A(n7054), .Z(n10947) );
  XNOR U10552 ( .A(n10950), .B(n9185), .Z(n7054) );
  IV U10553 ( .A(n10037), .Z(n9185) );
  XOR U10554 ( .A(n10951), .B(n6997), .Z(n8152) );
  NOR U10555 ( .A(n10834), .B(n8097), .Z(n10951) );
  XNOR U10556 ( .A(n10932), .B(n10952), .Z(n8097) );
  AND U10557 ( .A(n5593), .B(n6605), .Z(n10927) );
  XOR U10558 ( .A(n10953), .B(n1711), .Z(n6605) );
  XNOR U10559 ( .A(n8968), .B(n6226), .Z(n1711) );
  XNOR U10560 ( .A(n10954), .B(n10955), .Z(n6226) );
  XOR U10561 ( .A(n5359), .B(n3606), .Z(n10955) );
  XOR U10562 ( .A(n10956), .B(n10957), .Z(n3606) );
  XOR U10563 ( .A(n10959), .B(n10960), .Z(n5359) );
  ANDN U10564 ( .B(n8106), .A(n10961), .Z(n10959) );
  XNOR U10565 ( .A(n10962), .B(n10963), .Z(n10954) );
  XNOR U10566 ( .A(n2071), .B(n5466), .Z(n10963) );
  XOR U10567 ( .A(n10964), .B(n10965), .Z(n5466) );
  AND U10568 ( .A(n10966), .B(n10967), .Z(n10964) );
  XNOR U10569 ( .A(n10968), .B(n10969), .Z(n2071) );
  ANDN U10570 ( .B(n10970), .A(n9124), .Z(n10968) );
  XOR U10571 ( .A(n10971), .B(n10972), .Z(n8968) );
  XOR U10572 ( .A(n3431), .B(n5033), .Z(n10972) );
  XNOR U10573 ( .A(n10973), .B(n8051), .Z(n5033) );
  AND U10574 ( .A(n8050), .B(n10974), .Z(n10973) );
  XNOR U10575 ( .A(n10975), .B(n9034), .Z(n3431) );
  AND U10576 ( .A(n9033), .B(n10857), .Z(n10975) );
  XNOR U10577 ( .A(n4052), .B(n10976), .Z(n10971) );
  XOR U10578 ( .A(n8040), .B(n2423), .Z(n10976) );
  XNOR U10579 ( .A(n10977), .B(n8061), .Z(n2423) );
  AND U10580 ( .A(n10978), .B(n10979), .Z(n10977) );
  XOR U10581 ( .A(n10980), .B(n8047), .Z(n8040) );
  AND U10582 ( .A(n10848), .B(n10981), .Z(n10980) );
  XNOR U10583 ( .A(n10982), .B(n8056), .Z(n4052) );
  XOR U10584 ( .A(n9879), .B(n2037), .Z(n5593) );
  XNOR U10585 ( .A(n7378), .B(n10983), .Z(n2037) );
  XOR U10586 ( .A(n10984), .B(n10985), .Z(n7378) );
  XNOR U10587 ( .A(n3734), .B(n5077), .Z(n10985) );
  XNOR U10588 ( .A(n10986), .B(n8470), .Z(n5077) );
  XNOR U10589 ( .A(n10987), .B(n10988), .Z(n8470) );
  NOR U10590 ( .A(n9877), .B(n9876), .Z(n10986) );
  XNOR U10591 ( .A(n9792), .B(n10989), .Z(n9876) );
  XOR U10592 ( .A(n10990), .B(n10991), .Z(n9877) );
  XOR U10593 ( .A(n10992), .B(n9962), .Z(n3734) );
  XNOR U10594 ( .A(n10830), .B(n10993), .Z(n9962) );
  AND U10595 ( .A(n9885), .B(n10884), .Z(n10992) );
  IV U10596 ( .A(n9886), .Z(n10884) );
  XNOR U10597 ( .A(n10994), .B(n10995), .Z(n9886) );
  XNOR U10598 ( .A(n10996), .B(n10997), .Z(n9885) );
  XOR U10599 ( .A(n4196), .B(n10998), .Z(n10984) );
  XOR U10600 ( .A(n1676), .B(n9952), .Z(n10998) );
  XOR U10601 ( .A(n10999), .B(n7434), .Z(n9952) );
  XNOR U10602 ( .A(n9513), .B(n11000), .Z(n7434) );
  AND U10603 ( .A(n9874), .B(n9873), .Z(n10999) );
  XOR U10604 ( .A(n11001), .B(n10256), .Z(n9873) );
  XNOR U10605 ( .A(n11002), .B(n11003), .Z(n9874) );
  XOR U10606 ( .A(n11004), .B(n7428), .Z(n1676) );
  IV U10607 ( .A(n9956), .Z(n7428) );
  XNOR U10608 ( .A(n10229), .B(n11005), .Z(n9956) );
  NOR U10609 ( .A(n9882), .B(n9883), .Z(n11004) );
  XNOR U10610 ( .A(n11006), .B(n10920), .Z(n9883) );
  XOR U10611 ( .A(n11007), .B(n11008), .Z(n9882) );
  XOR U10612 ( .A(n11009), .B(n7438), .Z(n4196) );
  IV U10613 ( .A(n9965), .Z(n7438) );
  XOR U10614 ( .A(n11010), .B(n10134), .Z(n9965) );
  ANDN U10615 ( .B(n10873), .A(n9964), .Z(n11009) );
  XNOR U10616 ( .A(n11011), .B(n9964), .Z(n9879) );
  XOR U10617 ( .A(n10917), .B(n11012), .Z(n9964) );
  NOR U10618 ( .A(n7437), .B(n10873), .Z(n11011) );
  XNOR U10619 ( .A(n10154), .B(n11013), .Z(n10873) );
  XNOR U10620 ( .A(n11014), .B(n11015), .Z(n7437) );
  XOR U10621 ( .A(n11016), .B(n6099), .Z(out[1014]) );
  XOR U10622 ( .A(n8220), .B(n4925), .Z(n6099) );
  XOR U10623 ( .A(n6062), .B(n5982), .Z(n4925) );
  XNOR U10624 ( .A(n11017), .B(n11018), .Z(n5982) );
  XNOR U10625 ( .A(n3629), .B(n4125), .Z(n11018) );
  XOR U10626 ( .A(n11019), .B(n8264), .Z(n4125) );
  ANDN U10627 ( .B(n8217), .A(n7100), .Z(n11019) );
  XOR U10628 ( .A(n11020), .B(n11021), .Z(n7100) );
  XNOR U10629 ( .A(n11022), .B(n10037), .Z(n8217) );
  XNOR U10630 ( .A(n11023), .B(n11024), .Z(n3629) );
  ANDN U10631 ( .B(n7109), .A(n8214), .Z(n11023) );
  XNOR U10632 ( .A(n10142), .B(n11025), .Z(n7109) );
  XOR U10633 ( .A(n5205), .B(n11026), .Z(n11017) );
  XNOR U10634 ( .A(n8235), .B(n1884), .Z(n11026) );
  XNOR U10635 ( .A(n11027), .B(n8255), .Z(n1884) );
  NOR U10636 ( .A(n7117), .B(n8209), .Z(n11027) );
  XOR U10637 ( .A(n11028), .B(n10661), .Z(n8209) );
  XNOR U10638 ( .A(n11029), .B(n11030), .Z(n7117) );
  XOR U10639 ( .A(n11031), .B(n8258), .Z(n8235) );
  NOR U10640 ( .A(n8212), .B(n7104), .Z(n11031) );
  XNOR U10641 ( .A(n11032), .B(n11033), .Z(n7104) );
  XOR U10642 ( .A(n11034), .B(n9582), .Z(n8212) );
  XNOR U10643 ( .A(n11035), .B(n8260), .Z(n5205) );
  AND U10644 ( .A(n7113), .B(n8261), .Z(n11035) );
  XOR U10645 ( .A(n11036), .B(n11037), .Z(n8261) );
  XNOR U10646 ( .A(n11038), .B(n9820), .Z(n7113) );
  XOR U10647 ( .A(n11039), .B(n11040), .Z(n6062) );
  XNOR U10648 ( .A(n3351), .B(n5704), .Z(n11040) );
  XNOR U10649 ( .A(n11041), .B(n7055), .Z(n5704) );
  XNOR U10650 ( .A(n11042), .B(n10823), .Z(n7055) );
  AND U10651 ( .A(n10948), .B(n11043), .Z(n11041) );
  XNOR U10652 ( .A(n11044), .B(n7063), .Z(n3351) );
  XOR U10653 ( .A(n11045), .B(n11046), .Z(n7063) );
  ANDN U10654 ( .B(n7064), .A(n8222), .Z(n11044) );
  XOR U10655 ( .A(n11047), .B(n10165), .Z(n8222) );
  XNOR U10656 ( .A(n11048), .B(n10599), .Z(n7064) );
  XOR U10657 ( .A(n5380), .B(n11049), .Z(n11039) );
  XOR U10658 ( .A(n7040), .B(n2241), .Z(n11049) );
  XNOR U10659 ( .A(n11050), .B(n7050), .Z(n2241) );
  XNOR U10660 ( .A(n11051), .B(n11052), .Z(n7050) );
  NOR U10661 ( .A(n7051), .B(n8225), .Z(n11050) );
  XNOR U10662 ( .A(n11053), .B(n10061), .Z(n8225) );
  XOR U10663 ( .A(n11054), .B(n11055), .Z(n7051) );
  XOR U10664 ( .A(n11056), .B(n7059), .Z(n7040) );
  XNOR U10665 ( .A(n10379), .B(n11058), .Z(n8227) );
  XOR U10666 ( .A(n11059), .B(n11060), .Z(n7060) );
  XNOR U10667 ( .A(n11061), .B(n7046), .Z(n5380) );
  XNOR U10668 ( .A(n11062), .B(n11063), .Z(n7046) );
  AND U10669 ( .A(n7047), .B(n8230), .Z(n11061) );
  XOR U10670 ( .A(n11064), .B(n11065), .Z(n8230) );
  XNOR U10671 ( .A(n11066), .B(n11067), .Z(n7047) );
  XOR U10672 ( .A(n11068), .B(n11043), .Z(n8220) );
  IV U10673 ( .A(n7056), .Z(n11043) );
  XOR U10674 ( .A(n11069), .B(n11070), .Z(n7056) );
  ANDN U10675 ( .B(n8174), .A(n10948), .Z(n11068) );
  XOR U10676 ( .A(n11071), .B(n11072), .Z(n10948) );
  IV U10677 ( .A(n10949), .Z(n8174) );
  XOR U10678 ( .A(n11073), .B(n10030), .Z(n10949) );
  IV U10679 ( .A(n11030), .Z(n10030) );
  XOR U10680 ( .A(n11074), .B(n11075), .Z(n11030) );
  AND U10681 ( .A(n5597), .B(n6632), .Z(n11016) );
  XNOR U10682 ( .A(n11076), .B(n1720), .Z(n6632) );
  XOR U10683 ( .A(n11077), .B(n11078), .Z(n9029) );
  XOR U10684 ( .A(n3433), .B(n5036), .Z(n11078) );
  XNOR U10685 ( .A(n11079), .B(n8112), .Z(n5036) );
  ANDN U10686 ( .B(n11080), .A(n10965), .Z(n11079) );
  XOR U10687 ( .A(n11081), .B(n9125), .Z(n3433) );
  IV U10688 ( .A(n11082), .Z(n9125) );
  AND U10689 ( .A(n10969), .B(n11083), .Z(n11081) );
  XNOR U10690 ( .A(n4086), .B(n11084), .Z(n11077) );
  XNOR U10691 ( .A(n8101), .B(n2432), .Z(n11084) );
  XOR U10692 ( .A(n11085), .B(n8121), .Z(n2432) );
  AND U10693 ( .A(n8122), .B(n11086), .Z(n11085) );
  XOR U10694 ( .A(n11087), .B(n8107), .Z(n8101) );
  AND U10695 ( .A(n10960), .B(n11088), .Z(n11087) );
  XOR U10696 ( .A(n11089), .B(n8117), .Z(n4086) );
  ANDN U10697 ( .B(n11090), .A(n10957), .Z(n11089) );
  XNOR U10698 ( .A(n11091), .B(n11092), .Z(n6231) );
  XNOR U10699 ( .A(n5369), .B(n3610), .Z(n11092) );
  XOR U10700 ( .A(n11093), .B(n11094), .Z(n3610) );
  AND U10701 ( .A(n11095), .B(n8142), .Z(n11093) );
  IV U10702 ( .A(n11096), .Z(n8142) );
  XNOR U10703 ( .A(n11097), .B(n11098), .Z(n5369) );
  NOR U10704 ( .A(n11099), .B(n8132), .Z(n11097) );
  XOR U10705 ( .A(n11100), .B(n11101), .Z(n11091) );
  XOR U10706 ( .A(n2075), .B(n5511), .Z(n11101) );
  XOR U10707 ( .A(n11102), .B(n11103), .Z(n5511) );
  ANDN U10708 ( .B(n11104), .A(n8136), .Z(n11102) );
  XOR U10709 ( .A(n11105), .B(n11106), .Z(n2075) );
  ANDN U10710 ( .B(n11107), .A(n9224), .Z(n11105) );
  XOR U10711 ( .A(n9975), .B(n2041), .Z(n5597) );
  IV U10712 ( .A(n5136), .Z(n2041) );
  XOR U10713 ( .A(n8653), .B(n7440), .Z(n5136) );
  XNOR U10714 ( .A(n11108), .B(n11109), .Z(n7440) );
  XOR U10715 ( .A(n10067), .B(n4199), .Z(n11109) );
  XOR U10716 ( .A(n11110), .B(n7546), .Z(n4199) );
  IV U10717 ( .A(n10417), .Z(n7546) );
  XOR U10718 ( .A(n11111), .B(n10279), .Z(n10417) );
  AND U10719 ( .A(n11112), .B(n10418), .Z(n11110) );
  XNOR U10720 ( .A(n11113), .B(n7542), .Z(n10067) );
  XNOR U10721 ( .A(n11114), .B(n9584), .Z(n7542) );
  ANDN U10722 ( .B(n9969), .A(n9970), .Z(n11113) );
  XNOR U10723 ( .A(n11115), .B(n10386), .Z(n9969) );
  XOR U10724 ( .A(n3740), .B(n11116), .Z(n11108) );
  XOR U10725 ( .A(n5086), .B(n1681), .Z(n11116) );
  XOR U10726 ( .A(n11117), .B(n7536), .Z(n1681) );
  IV U10727 ( .A(n10408), .Z(n7536) );
  XOR U10728 ( .A(n11118), .B(n10065), .Z(n10408) );
  ANDN U10729 ( .B(n9979), .A(n9978), .Z(n11117) );
  XNOR U10730 ( .A(n11119), .B(n11072), .Z(n9978) );
  XOR U10731 ( .A(n11120), .B(n8595), .Z(n5086) );
  XOR U10732 ( .A(n11121), .B(n11122), .Z(n8595) );
  ANDN U10733 ( .B(n9982), .A(n9981), .Z(n11120) );
  XNOR U10734 ( .A(n9914), .B(n11123), .Z(n9981) );
  XNOR U10735 ( .A(n11124), .B(n10415), .Z(n3740) );
  XOR U10736 ( .A(n11125), .B(n11126), .Z(n9972) );
  XOR U10737 ( .A(n11127), .B(n11128), .Z(n8653) );
  XOR U10738 ( .A(n6192), .B(n2286), .Z(n11128) );
  XNOR U10739 ( .A(n11129), .B(n10076), .Z(n2286) );
  NOR U10740 ( .A(n7616), .B(n7617), .Z(n11129) );
  XOR U10741 ( .A(n11130), .B(n9532), .Z(n7616) );
  IV U10742 ( .A(n9914), .Z(n9532) );
  XOR U10743 ( .A(n11131), .B(n11132), .Z(n9914) );
  XNOR U10744 ( .A(n11133), .B(n10081), .Z(n6192) );
  ANDN U10745 ( .B(n7607), .A(n7608), .Z(n11133) );
  XNOR U10746 ( .A(n9558), .B(n11134), .Z(n7607) );
  XOR U10747 ( .A(n3853), .B(n11135), .Z(n11127) );
  XNOR U10748 ( .A(n5110), .B(n5399), .Z(n11135) );
  XNOR U10749 ( .A(n11136), .B(n10073), .Z(n5399) );
  XNOR U10750 ( .A(n11137), .B(n10279), .Z(n7620) );
  XOR U10751 ( .A(n11138), .B(n10084), .Z(n5110) );
  AND U10752 ( .A(n8652), .B(n8650), .Z(n11138) );
  XOR U10753 ( .A(n11139), .B(n10121), .Z(n8650) );
  XOR U10754 ( .A(n11140), .B(n11141), .Z(n3853) );
  ANDN U10755 ( .B(n7614), .A(n7612), .Z(n11140) );
  XOR U10756 ( .A(n11142), .B(n10418), .Z(n9975) );
  XOR U10757 ( .A(n11143), .B(n10995), .Z(n10418) );
  NOR U10758 ( .A(n7544), .B(n11112), .Z(n11142) );
  XOR U10759 ( .A(n11144), .B(n6104), .Z(out[1013]) );
  XNOR U10760 ( .A(n8253), .B(n4929), .Z(n6104) );
  XOR U10761 ( .A(n6067), .B(n5987), .Z(n4929) );
  XNOR U10762 ( .A(n11145), .B(n11146), .Z(n5987) );
  XNOR U10763 ( .A(n3635), .B(n4128), .Z(n11146) );
  XNOR U10764 ( .A(n11147), .B(n8316), .Z(n4128) );
  ANDN U10765 ( .B(n8249), .A(n7128), .Z(n11147) );
  XNOR U10766 ( .A(n11148), .B(n11149), .Z(n7128) );
  XOR U10767 ( .A(n10142), .B(n11150), .Z(n8249) );
  XNOR U10768 ( .A(n11151), .B(n11152), .Z(n3635) );
  ANDN U10769 ( .B(n7141), .A(n8247), .Z(n11151) );
  XOR U10770 ( .A(n11153), .B(n10286), .Z(n7141) );
  IV U10771 ( .A(n9364), .Z(n10286) );
  XOR U10772 ( .A(n5207), .B(n11154), .Z(n11145) );
  XNOR U10773 ( .A(n8291), .B(n1889), .Z(n11154) );
  XOR U10774 ( .A(n11155), .B(n11156), .Z(n1889) );
  ANDN U10775 ( .B(n8242), .A(n7145), .Z(n11155) );
  XOR U10776 ( .A(n11157), .B(n10134), .Z(n7145) );
  XNOR U10777 ( .A(n11158), .B(n9270), .Z(n8242) );
  XOR U10778 ( .A(n11159), .B(n8312), .Z(n8291) );
  NOR U10779 ( .A(n7132), .B(n8245), .Z(n11159) );
  XNOR U10780 ( .A(n11160), .B(n9692), .Z(n8245) );
  XNOR U10781 ( .A(n11161), .B(n11162), .Z(n7132) );
  XNOR U10782 ( .A(n11163), .B(n8314), .Z(n5207) );
  AND U10783 ( .A(n8239), .B(n7137), .Z(n11163) );
  XOR U10784 ( .A(n9941), .B(n11164), .Z(n7137) );
  IV U10785 ( .A(n10898), .Z(n9941) );
  XNOR U10786 ( .A(n11165), .B(n11166), .Z(n8239) );
  XOR U10787 ( .A(n11167), .B(n11168), .Z(n6067) );
  XNOR U10788 ( .A(n3354), .B(n5728), .Z(n11168) );
  XOR U10789 ( .A(n11169), .B(n8215), .Z(n5728) );
  IV U10790 ( .A(n7111), .Z(n8215) );
  XNOR U10791 ( .A(n11170), .B(n10938), .Z(n7111) );
  ANDN U10792 ( .B(n11024), .A(n7110), .Z(n11169) );
  XNOR U10793 ( .A(n11171), .B(n7119), .Z(n3354) );
  XNOR U10794 ( .A(n11172), .B(n11173), .Z(n7119) );
  ANDN U10795 ( .B(n8255), .A(n7118), .Z(n11171) );
  XNOR U10796 ( .A(n11174), .B(n11175), .Z(n7118) );
  XOR U10797 ( .A(n11176), .B(n11177), .Z(n8255) );
  XOR U10798 ( .A(n5384), .B(n11178), .Z(n11167) );
  XNOR U10799 ( .A(n7095), .B(n2248), .Z(n11178) );
  XNOR U10800 ( .A(n11179), .B(n7106), .Z(n2248) );
  XOR U10801 ( .A(n11180), .B(n11065), .Z(n7106) );
  NOR U10802 ( .A(n7105), .B(n8258), .Z(n11179) );
  XOR U10803 ( .A(n11181), .B(n11182), .Z(n8258) );
  XNOR U10804 ( .A(n9088), .B(n11183), .Z(n7105) );
  XNOR U10805 ( .A(n11184), .B(n7114), .Z(n7095) );
  XNOR U10806 ( .A(n11185), .B(n10665), .Z(n7114) );
  ANDN U10807 ( .B(n7115), .A(n8260), .Z(n11184) );
  XNOR U10808 ( .A(n10559), .B(n11186), .Z(n8260) );
  XNOR U10809 ( .A(n11187), .B(n11188), .Z(n7115) );
  XOR U10810 ( .A(n11189), .B(n7101), .Z(n5384) );
  XNOR U10811 ( .A(n9094), .B(n11190), .Z(n7101) );
  XOR U10812 ( .A(n11191), .B(n11192), .Z(n8264) );
  IV U10813 ( .A(n7102), .Z(n8263) );
  XOR U10814 ( .A(n11193), .B(n11194), .Z(n7102) );
  XNOR U10815 ( .A(n11195), .B(n7110), .Z(n8253) );
  XNOR U10816 ( .A(n11196), .B(n10788), .Z(n7110) );
  IV U10817 ( .A(n11197), .Z(n10788) );
  ANDN U10818 ( .B(n8214), .A(n11024), .Z(n11195) );
  XOR U10819 ( .A(n11198), .B(n11199), .Z(n11024) );
  XNOR U10820 ( .A(n11200), .B(n10134), .Z(n8214) );
  AND U10821 ( .A(n5605), .B(n6659), .Z(n11144) );
  XOR U10822 ( .A(n11201), .B(n1725), .Z(n6659) );
  XOR U10823 ( .A(n11202), .B(n11203), .Z(n9121) );
  XNOR U10824 ( .A(n3435), .B(n5041), .Z(n11203) );
  XOR U10825 ( .A(n11204), .B(n8137), .Z(n5041) );
  ANDN U10826 ( .B(n11205), .A(n11103), .Z(n11204) );
  XNOR U10827 ( .A(n11206), .B(n9226), .Z(n3435) );
  NOR U10828 ( .A(n11106), .B(n9225), .Z(n11206) );
  XOR U10829 ( .A(n4123), .B(n11207), .Z(n11202) );
  XOR U10830 ( .A(n8127), .B(n2437), .Z(n11207) );
  XNOR U10831 ( .A(n11208), .B(n8147), .Z(n2437) );
  AND U10832 ( .A(n8148), .B(n11209), .Z(n11208) );
  XOR U10833 ( .A(n11210), .B(n8133), .Z(n8127) );
  AND U10834 ( .A(n11098), .B(n8134), .Z(n11210) );
  XNOR U10835 ( .A(n11211), .B(n8143), .Z(n4123) );
  AND U10836 ( .A(n8144), .B(n11212), .Z(n11211) );
  XNOR U10837 ( .A(n11213), .B(n11214), .Z(n6235) );
  XOR U10838 ( .A(n5373), .B(n3614), .Z(n11214) );
  XOR U10839 ( .A(n11215), .B(n11216), .Z(n3614) );
  AND U10840 ( .A(n11217), .B(n11218), .Z(n11215) );
  XOR U10841 ( .A(n11219), .B(n11220), .Z(n5373) );
  ANDN U10842 ( .B(n8186), .A(n11221), .Z(n11219) );
  XNOR U10843 ( .A(n11222), .B(n11223), .Z(n11213) );
  XOR U10844 ( .A(n2078), .B(n4259), .Z(n11223) );
  XNOR U10845 ( .A(n11224), .B(n11225), .Z(n4259) );
  ANDN U10846 ( .B(n11226), .A(n8190), .Z(n11224) );
  XOR U10847 ( .A(n11227), .B(n11228), .Z(n2078) );
  AND U10848 ( .A(n11229), .B(n11230), .Z(n11227) );
  XNOR U10849 ( .A(n10077), .B(n2046), .Z(n5605) );
  XNOR U10850 ( .A(n7529), .B(n8718), .Z(n2046) );
  XNOR U10851 ( .A(n11231), .B(n11232), .Z(n8718) );
  XOR U10852 ( .A(n5404), .B(n3858), .Z(n11232) );
  XOR U10853 ( .A(n11233), .B(n11234), .Z(n3858) );
  NOR U10854 ( .A(n7660), .B(n7661), .Z(n11233) );
  XNOR U10855 ( .A(n9608), .B(n11235), .Z(n7661) );
  XOR U10856 ( .A(n11236), .B(n10182), .Z(n5404) );
  XNOR U10857 ( .A(n11237), .B(n11238), .Z(n7668) );
  XOR U10858 ( .A(n11239), .B(n9784), .Z(n7670) );
  XOR U10859 ( .A(n6196), .B(n11240), .Z(n11231) );
  XNOR U10860 ( .A(n2293), .B(n5137), .Z(n11240) );
  XNOR U10861 ( .A(n11241), .B(n10193), .Z(n5137) );
  ANDN U10862 ( .B(n8717), .A(n8715), .Z(n11241) );
  XOR U10863 ( .A(n11242), .B(n10265), .Z(n8715) );
  XNOR U10864 ( .A(n9892), .B(n11243), .Z(n8717) );
  XOR U10865 ( .A(n11244), .B(n11245), .Z(n2293) );
  NOR U10866 ( .A(n7665), .B(n7664), .Z(n11244) );
  XOR U10867 ( .A(n11246), .B(n9602), .Z(n7664) );
  XNOR U10868 ( .A(n11247), .B(n11248), .Z(n7665) );
  XNOR U10869 ( .A(n11249), .B(n10190), .Z(n6196) );
  ANDN U10870 ( .B(n7655), .A(n7656), .Z(n11249) );
  XNOR U10871 ( .A(n10154), .B(n11250), .Z(n7656) );
  XOR U10872 ( .A(n11251), .B(n9668), .Z(n7655) );
  XOR U10873 ( .A(n11252), .B(n11253), .Z(n7529) );
  XNOR U10874 ( .A(n3745), .B(n5088), .Z(n11253) );
  XOR U10875 ( .A(n11254), .B(n8651), .Z(n5088) );
  IV U10876 ( .A(n11255), .Z(n8651) );
  ANDN U10877 ( .B(n10084), .A(n10083), .Z(n11254) );
  XOR U10878 ( .A(n11256), .B(n11257), .Z(n10084) );
  XNOR U10879 ( .A(n11258), .B(n7618), .Z(n3745) );
  NOR U10880 ( .A(n10076), .B(n10075), .Z(n11258) );
  XNOR U10881 ( .A(n10107), .B(n11259), .Z(n10076) );
  XOR U10882 ( .A(n4201), .B(n11260), .Z(n11252) );
  XOR U10883 ( .A(n1685), .B(n10176), .Z(n11260) );
  XOR U10884 ( .A(n11261), .B(n7621), .Z(n10176) );
  ANDN U10885 ( .B(n10072), .A(n10073), .Z(n11261) );
  XNOR U10886 ( .A(n9673), .B(n11262), .Z(n10073) );
  XOR U10887 ( .A(n11263), .B(n7609), .Z(n1685) );
  IV U10888 ( .A(n11264), .Z(n7609) );
  NOR U10889 ( .A(n10080), .B(n10081), .Z(n11263) );
  XNOR U10890 ( .A(n11265), .B(n11126), .Z(n10081) );
  XNOR U10891 ( .A(n11266), .B(n7613), .Z(n4201) );
  AND U10892 ( .A(n11267), .B(n11141), .Z(n11266) );
  IV U10893 ( .A(n11268), .Z(n11141) );
  XOR U10894 ( .A(n11269), .B(n11267), .Z(n10077) );
  AND U10895 ( .A(n7612), .B(n11268), .Z(n11269) );
  XNOR U10896 ( .A(n10695), .B(n11270), .Z(n11268) );
  XNOR U10897 ( .A(n11271), .B(n10373), .Z(n7612) );
  XOR U10898 ( .A(n11272), .B(n6109), .Z(out[1012]) );
  XNOR U10899 ( .A(n8307), .B(n5897), .Z(n6109) );
  XOR U10900 ( .A(n6073), .B(n5992), .Z(n5897) );
  XNOR U10901 ( .A(n11273), .B(n11274), .Z(n5992) );
  XNOR U10902 ( .A(n3640), .B(n4131), .Z(n11274) );
  XNOR U10903 ( .A(n11275), .B(n8393), .Z(n4131) );
  NOR U10904 ( .A(n7197), .B(n8304), .Z(n11275) );
  XNOR U10905 ( .A(n11276), .B(n9364), .Z(n8304) );
  XOR U10906 ( .A(n11277), .B(n11278), .Z(n9364) );
  XOR U10907 ( .A(n11279), .B(n11280), .Z(n7197) );
  XNOR U10908 ( .A(n11281), .B(n11282), .Z(n3640) );
  AND U10909 ( .A(n7210), .B(n8302), .Z(n11281) );
  XNOR U10910 ( .A(n11283), .B(n9505), .Z(n7210) );
  XNOR U10911 ( .A(n5210), .B(n11284), .Z(n11273) );
  XNOR U10912 ( .A(n8366), .B(n1893), .Z(n11284) );
  XOR U10913 ( .A(n11285), .B(n8385), .Z(n1893) );
  AND U10914 ( .A(n8297), .B(n7214), .Z(n11285) );
  XOR U10915 ( .A(n11286), .B(n10279), .Z(n7214) );
  XOR U10916 ( .A(n11287), .B(n10448), .Z(n8297) );
  XNOR U10917 ( .A(n11288), .B(n8389), .Z(n8366) );
  ANDN U10918 ( .B(n8300), .A(n7201), .Z(n11288) );
  XOR U10919 ( .A(n11289), .B(n11067), .Z(n7201) );
  XNOR U10920 ( .A(n11290), .B(n9800), .Z(n8300) );
  XOR U10921 ( .A(n11291), .B(n8391), .Z(n5210) );
  ANDN U10922 ( .B(n7206), .A(n8295), .Z(n11291) );
  XNOR U10923 ( .A(n11292), .B(n11293), .Z(n8295) );
  XNOR U10924 ( .A(n10229), .B(n11294), .Z(n7206) );
  XOR U10925 ( .A(n11295), .B(n11296), .Z(n6073) );
  XNOR U10926 ( .A(n3362), .B(n5755), .Z(n11296) );
  XOR U10927 ( .A(n11297), .B(n7142), .Z(n5755) );
  XOR U10928 ( .A(n11298), .B(n11037), .Z(n7142) );
  AND U10929 ( .A(n7143), .B(n11152), .Z(n11297) );
  XOR U10930 ( .A(n11299), .B(n7147), .Z(n3362) );
  XNOR U10931 ( .A(n11300), .B(n10136), .Z(n7147) );
  ANDN U10932 ( .B(n11156), .A(n7146), .Z(n11299) );
  XOR U10933 ( .A(n11301), .B(n11302), .Z(n7146) );
  IV U10934 ( .A(n8309), .Z(n11156) );
  XOR U10935 ( .A(n9069), .B(n11303), .Z(n8309) );
  XOR U10936 ( .A(n5389), .B(n11304), .Z(n11295) );
  XNOR U10937 ( .A(n7123), .B(n2255), .Z(n11304) );
  XNOR U10938 ( .A(n11305), .B(n7133), .Z(n2255) );
  XNOR U10939 ( .A(n11306), .B(n11307), .Z(n7133) );
  ANDN U10940 ( .B(n8312), .A(n7134), .Z(n11305) );
  XOR U10941 ( .A(n9072), .B(n11308), .Z(n7134) );
  IV U10942 ( .A(n11309), .Z(n9072) );
  XOR U10943 ( .A(n11310), .B(n10803), .Z(n8312) );
  XOR U10944 ( .A(n11311), .B(n8240), .Z(n7123) );
  IV U10945 ( .A(n7139), .Z(n8240) );
  XOR U10946 ( .A(n10730), .B(n11312), .Z(n7139) );
  NOR U10947 ( .A(n7138), .B(n8314), .Z(n11311) );
  XOR U10948 ( .A(n11313), .B(n10679), .Z(n8314) );
  XOR U10949 ( .A(n11314), .B(n11315), .Z(n7138) );
  XOR U10950 ( .A(n11316), .B(n8250), .Z(n5389) );
  IV U10951 ( .A(n7130), .Z(n8250) );
  XOR U10952 ( .A(n11317), .B(n9216), .Z(n7130) );
  ANDN U10953 ( .B(n8316), .A(n7129), .Z(n11316) );
  XNOR U10954 ( .A(n9516), .B(n11318), .Z(n7129) );
  XNOR U10955 ( .A(n11319), .B(n11320), .Z(n8316) );
  XOR U10956 ( .A(n11321), .B(n7143), .Z(n8307) );
  XOR U10957 ( .A(n11322), .B(n10925), .Z(n7143) );
  ANDN U10958 ( .B(n8247), .A(n11152), .Z(n11321) );
  XOR U10959 ( .A(n11323), .B(n11324), .Z(n11152) );
  XOR U10960 ( .A(n11325), .B(n10279), .Z(n8247) );
  XOR U10961 ( .A(n11326), .B(n11327), .Z(n10279) );
  ANDN U10962 ( .B(n5609), .A(n5607), .Z(n11272) );
  XOR U10963 ( .A(n11328), .B(n1729), .Z(n5607) );
  XOR U10964 ( .A(n11329), .B(n11330), .Z(n9221) );
  XOR U10965 ( .A(n3437), .B(n5044), .Z(n11330) );
  XOR U10966 ( .A(n11331), .B(n8191), .Z(n5044) );
  AND U10967 ( .A(n8192), .B(n11225), .Z(n11331) );
  XNOR U10968 ( .A(n11332), .B(n9348), .Z(n3437) );
  ANDN U10969 ( .B(n9347), .A(n11228), .Z(n11332) );
  XNOR U10970 ( .A(n4159), .B(n11333), .Z(n11329) );
  XNOR U10971 ( .A(n8181), .B(n2444), .Z(n11333) );
  XNOR U10972 ( .A(n11334), .B(n8201), .Z(n2444) );
  ANDN U10973 ( .B(n8202), .A(n11335), .Z(n11334) );
  XNOR U10974 ( .A(n11336), .B(n8188), .Z(n8181) );
  AND U10975 ( .A(n8187), .B(n11220), .Z(n11336) );
  XOR U10976 ( .A(n11337), .B(n8197), .Z(n4159) );
  AND U10977 ( .A(n11216), .B(n8198), .Z(n11337) );
  XNOR U10978 ( .A(n11338), .B(n11339), .Z(n6239) );
  XOR U10979 ( .A(n5377), .B(n3617), .Z(n11339) );
  XOR U10980 ( .A(n11340), .B(n11341), .Z(n3617) );
  ANDN U10981 ( .B(n11342), .A(n11343), .Z(n11340) );
  XNOR U10982 ( .A(n11344), .B(n11345), .Z(n5377) );
  AND U10983 ( .A(n11346), .B(n8270), .Z(n11344) );
  XNOR U10984 ( .A(n11347), .B(n11348), .Z(n11338) );
  XOR U10985 ( .A(n2081), .B(n4261), .Z(n11348) );
  XOR U10986 ( .A(n11349), .B(n11350), .Z(n4261) );
  XNOR U10987 ( .A(n11352), .B(n11353), .Z(n2081) );
  ANDN U10988 ( .B(n11354), .A(n9442), .Z(n11352) );
  XNOR U10989 ( .A(n10186), .B(n2049), .Z(n5609) );
  XNOR U10990 ( .A(n7602), .B(n8777), .Z(n2049) );
  XNOR U10991 ( .A(n11355), .B(n11356), .Z(n8777) );
  XOR U10992 ( .A(n5407), .B(n3862), .Z(n11356) );
  XOR U10993 ( .A(n11357), .B(n11358), .Z(n3862) );
  ANDN U10994 ( .B(n10518), .A(n7745), .Z(n11357) );
  IV U10995 ( .A(n7746), .Z(n10518) );
  XNOR U10996 ( .A(n11359), .B(n9718), .Z(n7746) );
  XNOR U10997 ( .A(n10316), .B(n11360), .Z(n5407) );
  XOR U10998 ( .A(n11361), .B(n11362), .Z(n11360) );
  NAND U10999 ( .A(n11363), .B(n11364), .Z(n11362) );
  AND U11000 ( .A(n6455), .B(n11365), .Z(n11364) );
  ANDN U11001 ( .B(n10317), .A(n7742), .Z(n11361) );
  XOR U11002 ( .A(n11366), .B(n11367), .Z(n7742) );
  XNOR U11003 ( .A(n11368), .B(n11369), .Z(n10317) );
  XOR U11004 ( .A(n6200), .B(n11370), .Z(n11355) );
  XOR U11005 ( .A(n2304), .B(n5169), .Z(n11370) );
  XNOR U11006 ( .A(n11371), .B(n10328), .Z(n5169) );
  XOR U11007 ( .A(n11372), .B(n11373), .Z(n8780) );
  XOR U11008 ( .A(n11374), .B(n10022), .Z(n8781) );
  XNOR U11009 ( .A(n11375), .B(n10320), .Z(n2304) );
  ANDN U11010 ( .B(n7732), .A(n7731), .Z(n11375) );
  XNOR U11011 ( .A(n11376), .B(n11377), .Z(n7731) );
  XNOR U11012 ( .A(n11379), .B(n10325), .Z(n6200) );
  ANDN U11013 ( .B(n7737), .A(n7735), .Z(n11379) );
  XNOR U11014 ( .A(n11380), .B(n10371), .Z(n7735) );
  XNOR U11015 ( .A(n11381), .B(n10296), .Z(n7737) );
  XOR U11016 ( .A(n11382), .B(n11383), .Z(n7602) );
  XNOR U11017 ( .A(n3749), .B(n5090), .Z(n11383) );
  XOR U11018 ( .A(n11384), .B(n8716), .Z(n5090) );
  XNOR U11019 ( .A(n10706), .B(n11385), .Z(n8716) );
  NOR U11020 ( .A(n10337), .B(n10193), .Z(n11384) );
  XNOR U11021 ( .A(n11386), .B(n11387), .Z(n10193) );
  IV U11022 ( .A(n10192), .Z(n10337) );
  XOR U11023 ( .A(n9710), .B(n11388), .Z(n10192) );
  IV U11024 ( .A(n11376), .Z(n9710) );
  XOR U11025 ( .A(n11389), .B(n7666), .Z(n3749) );
  XNOR U11026 ( .A(n11390), .B(n11162), .Z(n7666) );
  AND U11027 ( .A(n10184), .B(n11245), .Z(n11389) );
  IV U11028 ( .A(n10185), .Z(n11245) );
  XNOR U11029 ( .A(n11391), .B(n10219), .Z(n10185) );
  XNOR U11030 ( .A(n9116), .B(n11392), .Z(n10184) );
  XNOR U11031 ( .A(n4204), .B(n11393), .Z(n11382) );
  XOR U11032 ( .A(n1689), .B(n10311), .Z(n11393) );
  XNOR U11033 ( .A(n11394), .B(n7669), .Z(n10311) );
  XOR U11034 ( .A(n11395), .B(n9798), .Z(n7669) );
  IV U11035 ( .A(n10785), .Z(n9798) );
  AND U11036 ( .A(n10182), .B(n10181), .Z(n11394) );
  XOR U11037 ( .A(n11396), .B(n11397), .Z(n10181) );
  XNOR U11038 ( .A(n11398), .B(n9780), .Z(n10182) );
  IV U11039 ( .A(n10875), .Z(n9780) );
  XOR U11040 ( .A(n11399), .B(n10333), .Z(n1689) );
  IV U11041 ( .A(n7657), .Z(n10333) );
  XNOR U11042 ( .A(n11400), .B(n10307), .Z(n7657) );
  NOR U11043 ( .A(n10189), .B(n10190), .Z(n11399) );
  XOR U11044 ( .A(n11401), .B(n11402), .Z(n10190) );
  XNOR U11045 ( .A(n11403), .B(n11404), .Z(n10189) );
  XOR U11046 ( .A(n11405), .B(n7662), .Z(n4204) );
  XNOR U11047 ( .A(n11406), .B(n11369), .Z(n7662) );
  AND U11048 ( .A(n11234), .B(n10339), .Z(n11405) );
  XNOR U11049 ( .A(n11407), .B(n10339), .Z(n10186) );
  XNOR U11050 ( .A(n10107), .B(n11408), .Z(n10339) );
  IV U11051 ( .A(n11409), .Z(n10107) );
  ANDN U11052 ( .B(n7660), .A(n11234), .Z(n11407) );
  XNOR U11053 ( .A(n11410), .B(n10594), .Z(n11234) );
  XOR U11054 ( .A(n11411), .B(n11412), .Z(n7660) );
  XOR U11055 ( .A(n11413), .B(n6119), .Z(out[1011]) );
  XNOR U11056 ( .A(n8382), .B(n5952), .Z(n6119) );
  XOR U11057 ( .A(n6078), .B(n5997), .Z(n5952) );
  XNOR U11058 ( .A(n11414), .B(n11415), .Z(n5997) );
  XOR U11059 ( .A(n3645), .B(n4134), .Z(n11415) );
  XNOR U11060 ( .A(n11416), .B(n8466), .Z(n4134) );
  ANDN U11061 ( .B(n7252), .A(n8379), .Z(n11416) );
  XOR U11062 ( .A(n11417), .B(n9505), .Z(n8379) );
  XOR U11063 ( .A(n11418), .B(n11419), .Z(n7252) );
  XOR U11064 ( .A(n11420), .B(n11421), .Z(n3645) );
  ANDN U11065 ( .B(n7265), .A(n8377), .Z(n11420) );
  XOR U11066 ( .A(n9564), .B(n11422), .Z(n7265) );
  XNOR U11067 ( .A(n5213), .B(n11423), .Z(n11414) );
  XNOR U11068 ( .A(n8440), .B(n1897), .Z(n11423) );
  XOR U11069 ( .A(n11424), .B(n8459), .Z(n1897) );
  AND U11070 ( .A(n8372), .B(n7269), .Z(n11424) );
  XNOR U11071 ( .A(n11425), .B(n11238), .Z(n7269) );
  XNOR U11072 ( .A(n9502), .B(n11426), .Z(n8372) );
  XOR U11073 ( .A(n11427), .B(n8462), .Z(n8440) );
  IV U11074 ( .A(n11428), .Z(n8462) );
  NOR U11075 ( .A(n8375), .B(n7256), .Z(n11427) );
  XOR U11076 ( .A(n11429), .B(n9390), .Z(n7256) );
  IV U11077 ( .A(n11194), .Z(n9390) );
  XOR U11078 ( .A(n11430), .B(n9922), .Z(n8375) );
  XOR U11079 ( .A(n11431), .B(n8464), .Z(n5213) );
  AND U11080 ( .A(n8370), .B(n7261), .Z(n11431) );
  XOR U11081 ( .A(n11432), .B(n10065), .Z(n7261) );
  XNOR U11082 ( .A(n11433), .B(n11434), .Z(n8370) );
  XOR U11083 ( .A(n11435), .B(n11436), .Z(n6078) );
  XOR U11084 ( .A(n3366), .B(n5781), .Z(n11436) );
  XOR U11085 ( .A(n11437), .B(n7212), .Z(n5781) );
  XNOR U11086 ( .A(n11438), .B(n11439), .Z(n7212) );
  AND U11087 ( .A(n7211), .B(n11282), .Z(n11437) );
  XNOR U11088 ( .A(n11440), .B(n7216), .Z(n3366) );
  XOR U11089 ( .A(n11441), .B(n11442), .Z(n7216) );
  ANDN U11090 ( .B(n8384), .A(n8385), .Z(n11440) );
  XNOR U11091 ( .A(n11443), .B(n9198), .Z(n8385) );
  IV U11092 ( .A(n10603), .Z(n9198) );
  XOR U11093 ( .A(n11444), .B(n10943), .Z(n8384) );
  XOR U11094 ( .A(n5393), .B(n11445), .Z(n11435) );
  XOR U11095 ( .A(n7192), .B(n2260), .Z(n11445) );
  XOR U11096 ( .A(n11446), .B(n7202), .Z(n2260) );
  XNOR U11097 ( .A(n11447), .B(n11448), .Z(n7202) );
  AND U11098 ( .A(n8389), .B(n8388), .Z(n11446) );
  XOR U11099 ( .A(n11449), .B(n11450), .Z(n8388) );
  XNOR U11100 ( .A(n11451), .B(n10478), .Z(n8389) );
  XNOR U11101 ( .A(n11452), .B(n7207), .Z(n7192) );
  XNOR U11102 ( .A(n10838), .B(n11453), .Z(n7207) );
  ANDN U11103 ( .B(n7208), .A(n8391), .Z(n11452) );
  XOR U11104 ( .A(n10922), .B(n11454), .Z(n8391) );
  XNOR U11105 ( .A(n11455), .B(n11456), .Z(n7208) );
  XOR U11106 ( .A(n11457), .B(n7199), .Z(n5393) );
  XOR U11107 ( .A(n11458), .B(n10473), .Z(n7199) );
  ANDN U11108 ( .B(n8393), .A(n7198), .Z(n11457) );
  XOR U11109 ( .A(n11459), .B(n9587), .Z(n7198) );
  XOR U11110 ( .A(n11460), .B(n9082), .Z(n8393) );
  XNOR U11111 ( .A(n11461), .B(n7211), .Z(n8382) );
  XNOR U11112 ( .A(n11462), .B(n11015), .Z(n7211) );
  NOR U11113 ( .A(n8302), .B(n11282), .Z(n11461) );
  XOR U11114 ( .A(n11463), .B(n11464), .Z(n11282) );
  XNOR U11115 ( .A(n11465), .B(n11466), .Z(n8302) );
  AND U11116 ( .A(n5613), .B(n5611), .Z(n11413) );
  XOR U11117 ( .A(n11467), .B(n1733), .Z(n5611) );
  XOR U11118 ( .A(n11468), .B(n11469), .Z(n9343) );
  XNOR U11119 ( .A(n3439), .B(n5047), .Z(n11469) );
  XOR U11120 ( .A(n11470), .B(n8275), .Z(n5047) );
  ANDN U11121 ( .B(n8276), .A(n11350), .Z(n11470) );
  XNOR U11122 ( .A(n11471), .B(n9444), .Z(n3439) );
  ANDN U11123 ( .B(n11353), .A(n9443), .Z(n11471) );
  XOR U11124 ( .A(n4192), .B(n11472), .Z(n11468) );
  XOR U11125 ( .A(n8265), .B(n2457), .Z(n11472) );
  XOR U11126 ( .A(n11473), .B(n8285), .Z(n2457) );
  ANDN U11127 ( .B(n8286), .A(n11474), .Z(n11473) );
  XOR U11128 ( .A(n11475), .B(n8272), .Z(n8265) );
  ANDN U11129 ( .B(n8271), .A(n11345), .Z(n11475) );
  XNOR U11130 ( .A(n11476), .B(n8282), .Z(n4192) );
  AND U11131 ( .A(n11341), .B(n11477), .Z(n11476) );
  XNOR U11132 ( .A(n11478), .B(n11479), .Z(n6243) );
  XNOR U11133 ( .A(n5383), .B(n3626), .Z(n11479) );
  ANDN U11134 ( .B(n11482), .A(n8332), .Z(n11480) );
  XNOR U11135 ( .A(n11483), .B(n11484), .Z(n5383) );
  ANDN U11136 ( .B(n11485), .A(n8322), .Z(n11483) );
  XOR U11137 ( .A(n11486), .B(n11487), .Z(n11478) );
  XOR U11138 ( .A(n2084), .B(n4266), .Z(n11487) );
  XNOR U11139 ( .A(n11488), .B(n11489), .Z(n4266) );
  AND U11140 ( .A(n8326), .B(n11490), .Z(n11488) );
  XNOR U11141 ( .A(n11491), .B(n11492), .Z(n2084) );
  AND U11142 ( .A(n11493), .B(n9544), .Z(n11491) );
  IV U11143 ( .A(n11494), .Z(n9544) );
  XNOR U11144 ( .A(n10321), .B(n5337), .Z(n5613) );
  XOR U11145 ( .A(n7650), .B(n8842), .Z(n5337) );
  XNOR U11146 ( .A(n11495), .B(n11496), .Z(n8842) );
  XNOR U11147 ( .A(n5412), .B(n3866), .Z(n11496) );
  XOR U11148 ( .A(n11497), .B(n11498), .Z(n3866) );
  ANDN U11149 ( .B(n7831), .A(n7832), .Z(n11497) );
  XNOR U11150 ( .A(n11499), .B(n9824), .Z(n7832) );
  IV U11151 ( .A(n11500), .Z(n7831) );
  XOR U11152 ( .A(n11501), .B(n10495), .Z(n5412) );
  ANDN U11153 ( .B(n10496), .A(n7828), .Z(n11501) );
  XNOR U11154 ( .A(n11502), .B(n11503), .Z(n7828) );
  XOR U11155 ( .A(n11504), .B(n10716), .Z(n10496) );
  XNOR U11156 ( .A(n6204), .B(n11505), .Z(n11495) );
  XNOR U11157 ( .A(n2311), .B(n5198), .Z(n11505) );
  XOR U11158 ( .A(n11506), .B(n10508), .Z(n5198) );
  NOR U11159 ( .A(n8845), .B(n8844), .Z(n11506) );
  XNOR U11160 ( .A(n10830), .B(n11507), .Z(n8844) );
  XNOR U11161 ( .A(n11508), .B(n10126), .Z(n8845) );
  XNOR U11162 ( .A(n11509), .B(n10499), .Z(n2311) );
  ANDN U11163 ( .B(n7817), .A(n7818), .Z(n11509) );
  XNOR U11164 ( .A(n11510), .B(n11511), .Z(n7818) );
  XOR U11165 ( .A(n11512), .B(n9817), .Z(n7817) );
  XOR U11166 ( .A(n11513), .B(n10505), .Z(n6204) );
  AND U11167 ( .A(n7823), .B(n7821), .Z(n11513) );
  IV U11168 ( .A(n10504), .Z(n7821) );
  XOR U11169 ( .A(n11514), .B(n11515), .Z(n10504) );
  XNOR U11170 ( .A(n10695), .B(n11516), .Z(n7823) );
  XOR U11171 ( .A(n11517), .B(n11518), .Z(n7650) );
  XNOR U11172 ( .A(n3754), .B(n5092), .Z(n11518) );
  XOR U11173 ( .A(n11519), .B(n8782), .Z(n5092) );
  XNOR U11174 ( .A(n11520), .B(n10806), .Z(n8782) );
  ANDN U11175 ( .B(n10327), .A(n10328), .Z(n11519) );
  XOR U11176 ( .A(n11521), .B(n11522), .Z(n10328) );
  XOR U11177 ( .A(n11523), .B(n10709), .Z(n10327) );
  IV U11178 ( .A(n9817), .Z(n10709) );
  XOR U11179 ( .A(n11524), .B(n11525), .Z(n9817) );
  XOR U11180 ( .A(n11526), .B(n7733), .Z(n3754) );
  XNOR U11181 ( .A(n11527), .B(n11067), .Z(n7733) );
  ANDN U11182 ( .B(n10319), .A(n10320), .Z(n11526) );
  XOR U11183 ( .A(n11528), .B(n10431), .Z(n10320) );
  XNOR U11184 ( .A(n11529), .B(n9190), .Z(n10319) );
  XNOR U11185 ( .A(n4207), .B(n11530), .Z(n11517) );
  XOR U11186 ( .A(n1693), .B(n10490), .Z(n11530) );
  XOR U11187 ( .A(n11531), .B(n7743), .Z(n10490) );
  XNOR U11188 ( .A(n11532), .B(n9924), .Z(n7743) );
  XNOR U11189 ( .A(n11533), .B(n11534), .Z(n9924) );
  ANDN U11190 ( .B(n10315), .A(n10316), .Z(n11531) );
  XNOR U11191 ( .A(n11535), .B(n9904), .Z(n10316) );
  XNOR U11192 ( .A(n11536), .B(n11197), .Z(n10315) );
  XNOR U11193 ( .A(n11537), .B(n10513), .Z(n1693) );
  XOR U11194 ( .A(n11538), .B(n11539), .Z(n10513) );
  ANDN U11195 ( .B(n10324), .A(n10325), .Z(n11537) );
  XOR U11196 ( .A(n9116), .B(n11540), .Z(n10325) );
  XNOR U11197 ( .A(n11541), .B(n11542), .Z(n9116) );
  XNOR U11198 ( .A(n11543), .B(n11544), .Z(n10324) );
  XOR U11199 ( .A(n11545), .B(n7747), .Z(n4207) );
  XOR U11200 ( .A(n11546), .B(n10716), .Z(n7747) );
  XOR U11201 ( .A(n11547), .B(n10519), .Z(n10321) );
  XNOR U11202 ( .A(n11548), .B(n10219), .Z(n10519) );
  ANDN U11203 ( .B(n7745), .A(n11358), .Z(n11547) );
  XNOR U11204 ( .A(n11549), .B(n11550), .Z(n11358) );
  XOR U11205 ( .A(n11551), .B(n10675), .Z(n7745) );
  XOR U11206 ( .A(n11552), .B(n6124), .Z(out[1010]) );
  XOR U11207 ( .A(n8457), .B(n6007), .Z(n6124) );
  XOR U11208 ( .A(n6001), .B(n6083), .Z(n6007) );
  XNOR U11209 ( .A(n11553), .B(n11554), .Z(n6083) );
  XOR U11210 ( .A(n2267), .B(n5397), .Z(n11554) );
  XOR U11211 ( .A(n11555), .B(n7254), .Z(n5397) );
  XOR U11212 ( .A(n11556), .B(n10233), .Z(n7254) );
  ANDN U11213 ( .B(n8466), .A(n7253), .Z(n11555) );
  XOR U11214 ( .A(n11557), .B(n9697), .Z(n7253) );
  XNOR U11215 ( .A(n9208), .B(n11558), .Z(n8466) );
  XOR U11216 ( .A(n11559), .B(n7258), .Z(n2267) );
  XOR U11217 ( .A(n11560), .B(n9082), .Z(n7258) );
  AND U11218 ( .A(n7257), .B(n11428), .Z(n11559) );
  XNOR U11219 ( .A(n11561), .B(n10599), .Z(n11428) );
  XOR U11220 ( .A(n11562), .B(n11563), .Z(n7257) );
  XNOR U11221 ( .A(n3119), .B(n11564), .Z(n11553) );
  XOR U11222 ( .A(n5810), .B(n7247), .Z(n11564) );
  XNOR U11223 ( .A(n11565), .B(n7262), .Z(n7247) );
  XOR U11224 ( .A(n11566), .B(n11567), .Z(n7262) );
  ANDN U11225 ( .B(n7263), .A(n8464), .Z(n11565) );
  XOR U11226 ( .A(n10917), .B(n11568), .Z(n8464) );
  XNOR U11227 ( .A(n11569), .B(n11570), .Z(n7263) );
  XNOR U11228 ( .A(n11571), .B(n7267), .Z(n5810) );
  XNOR U11229 ( .A(n11572), .B(n11573), .Z(n7267) );
  NOR U11230 ( .A(n7266), .B(n11421), .Z(n11571) );
  XOR U11231 ( .A(n11574), .B(n7270), .Z(n3119) );
  XNOR U11232 ( .A(n11575), .B(n10464), .Z(n7270) );
  ANDN U11233 ( .B(n7271), .A(n8459), .Z(n11574) );
  XNOR U11234 ( .A(n11576), .B(n10017), .Z(n8459) );
  XNOR U11235 ( .A(n11577), .B(n11021), .Z(n7271) );
  XOR U11236 ( .A(n11578), .B(n11579), .Z(n6001) );
  XNOR U11237 ( .A(n5216), .B(n1901), .Z(n11579) );
  XOR U11238 ( .A(n11580), .B(n8528), .Z(n1901) );
  AND U11239 ( .A(n7342), .B(n8529), .Z(n11580) );
  XNOR U11240 ( .A(n9097), .B(n11581), .Z(n8529) );
  XNOR U11241 ( .A(n11582), .B(n11369), .Z(n7342) );
  XOR U11242 ( .A(n11583), .B(n8535), .Z(n5216) );
  ANDN U11243 ( .B(n8444), .A(n7334), .Z(n11583) );
  XNOR U11244 ( .A(n11584), .B(n10172), .Z(n7334) );
  XNOR U11245 ( .A(n11585), .B(n11586), .Z(n8444) );
  XNOR U11246 ( .A(n3651), .B(n11587), .Z(n11578) );
  XOR U11247 ( .A(n8509), .B(n4137), .Z(n11587) );
  XNOR U11248 ( .A(n11588), .B(n8537), .Z(n4137) );
  ANDN U11249 ( .B(n8454), .A(n7325), .Z(n11588) );
  XOR U11250 ( .A(n11589), .B(n11590), .Z(n7325) );
  XOR U11251 ( .A(n10577), .B(n11591), .Z(n8454) );
  IV U11252 ( .A(n9564), .Z(n10577) );
  XNOR U11253 ( .A(n11592), .B(n8532), .Z(n8509) );
  AND U11254 ( .A(n7329), .B(n8533), .Z(n11592) );
  XOR U11255 ( .A(n11593), .B(n11594), .Z(n8533) );
  XOR U11256 ( .A(n9516), .B(n11595), .Z(n7329) );
  XNOR U11257 ( .A(n11596), .B(n11597), .Z(n3651) );
  AND U11258 ( .A(n8452), .B(n7338), .Z(n11596) );
  XOR U11259 ( .A(n11598), .B(n9676), .Z(n7338) );
  XOR U11260 ( .A(n11599), .B(n7266), .Z(n8457) );
  XNOR U11261 ( .A(n11600), .B(n10245), .Z(n7266) );
  AND U11262 ( .A(n8377), .B(n11421), .Z(n11599) );
  XNOR U11263 ( .A(n11601), .B(n11602), .Z(n11421) );
  XNOR U11264 ( .A(n11603), .B(n11369), .Z(n8377) );
  ANDN U11265 ( .B(n5617), .A(n5615), .Z(n11552) );
  XNOR U11266 ( .A(n11604), .B(n1738), .Z(n5615) );
  XOR U11267 ( .A(n11605), .B(n11606), .Z(n9439) );
  XOR U11268 ( .A(n3442), .B(n5054), .Z(n11606) );
  XNOR U11269 ( .A(n11607), .B(n8328), .Z(n5054) );
  ANDN U11270 ( .B(n11489), .A(n8327), .Z(n11607) );
  XNOR U11271 ( .A(n11608), .B(n9546), .Z(n3442) );
  ANDN U11272 ( .B(n11492), .A(n9545), .Z(n11608) );
  XOR U11273 ( .A(n4217), .B(n11609), .Z(n11605) );
  XOR U11274 ( .A(n8317), .B(n2462), .Z(n11609) );
  XOR U11275 ( .A(n11610), .B(n8337), .Z(n2462) );
  ANDN U11276 ( .B(n8338), .A(n11611), .Z(n11610) );
  XOR U11277 ( .A(n11612), .B(n8323), .Z(n8317) );
  ANDN U11278 ( .B(n8324), .A(n11484), .Z(n11612) );
  XOR U11279 ( .A(n11613), .B(n8334), .Z(n4217) );
  ANDN U11280 ( .B(n11481), .A(n8333), .Z(n11613) );
  XNOR U11281 ( .A(n11614), .B(n11615), .Z(n6247) );
  XNOR U11282 ( .A(n5387), .B(n3630), .Z(n11615) );
  XNOR U11283 ( .A(n11616), .B(n11617), .Z(n3630) );
  ANDN U11284 ( .B(n11618), .A(n8359), .Z(n11616) );
  XNOR U11285 ( .A(n11619), .B(n11620), .Z(n5387) );
  AND U11286 ( .A(n8349), .B(n11621), .Z(n11619) );
  XOR U11287 ( .A(n11622), .B(n11623), .Z(n11614) );
  XNOR U11288 ( .A(n2087), .B(n4268), .Z(n11623) );
  XNOR U11289 ( .A(n11624), .B(n11625), .Z(n4268) );
  AND U11290 ( .A(n8353), .B(n11626), .Z(n11624) );
  XOR U11291 ( .A(n11627), .B(n11628), .Z(n2087) );
  AND U11292 ( .A(n11629), .B(n9652), .Z(n11627) );
  IV U11293 ( .A(n11630), .Z(n9652) );
  XOR U11294 ( .A(n10500), .B(n2056), .Z(n5617) );
  XNOR U11295 ( .A(n7727), .B(n8905), .Z(n2056) );
  XNOR U11296 ( .A(n11631), .B(n11632), .Z(n8905) );
  XOR U11297 ( .A(n5421), .B(n3872), .Z(n11632) );
  NOR U11298 ( .A(n7880), .B(n7879), .Z(n11633) );
  XNOR U11299 ( .A(n11635), .B(n9946), .Z(n7880) );
  XOR U11300 ( .A(n11636), .B(n10613), .Z(n5421) );
  ANDN U11301 ( .B(n7875), .A(n7876), .Z(n11636) );
  XNOR U11302 ( .A(n11637), .B(n11173), .Z(n7876) );
  XOR U11303 ( .A(n11638), .B(n11639), .Z(n7875) );
  XNOR U11304 ( .A(n6208), .B(n11640), .Z(n11631) );
  XNOR U11305 ( .A(n2318), .B(n5228), .Z(n11640) );
  XNOR U11306 ( .A(n11641), .B(n10624), .Z(n5228) );
  NOR U11307 ( .A(n8909), .B(n8908), .Z(n11641) );
  XOR U11308 ( .A(n11642), .B(n10691), .Z(n8908) );
  XNOR U11309 ( .A(n11643), .B(n10270), .Z(n8909) );
  XOR U11310 ( .A(n11644), .B(n11645), .Z(n2318) );
  NOR U11311 ( .A(n7866), .B(n7865), .Z(n11644) );
  XNOR U11312 ( .A(n11646), .B(n10808), .Z(n7865) );
  XNOR U11313 ( .A(n9187), .B(n11647), .Z(n7866) );
  XOR U11314 ( .A(n11648), .B(n10621), .Z(n6208) );
  ANDN U11315 ( .B(n7871), .A(n7869), .Z(n11648) );
  XNOR U11316 ( .A(n11649), .B(n11650), .Z(n7869) );
  XNOR U11317 ( .A(n11651), .B(n10594), .Z(n7871) );
  XOR U11318 ( .A(n11652), .B(n11653), .Z(n7727) );
  XOR U11319 ( .A(n3760), .B(n5094), .Z(n11653) );
  XOR U11320 ( .A(n11654), .B(n8846), .Z(n5094) );
  IV U11321 ( .A(n10629), .Z(n8846) );
  XNOR U11322 ( .A(n11655), .B(n11656), .Z(n10629) );
  XOR U11323 ( .A(n11657), .B(n9938), .Z(n10507) );
  IV U11324 ( .A(n10808), .Z(n9938) );
  XOR U11325 ( .A(n11658), .B(n11659), .Z(n10808) );
  XNOR U11326 ( .A(n11660), .B(n9103), .Z(n10508) );
  XNOR U11327 ( .A(n11661), .B(n7819), .Z(n3760) );
  XOR U11328 ( .A(n11662), .B(n11194), .Z(n7819) );
  ANDN U11329 ( .B(n10498), .A(n10499), .Z(n11661) );
  XOR U11330 ( .A(n11663), .B(n11664), .Z(n10499) );
  IV U11331 ( .A(n10634), .Z(n10498) );
  XOR U11332 ( .A(n11665), .B(n11666), .Z(n10634) );
  XOR U11333 ( .A(n4210), .B(n11667), .Z(n11652) );
  XNOR U11334 ( .A(n1697), .B(n10608), .Z(n11667) );
  XNOR U11335 ( .A(n11668), .B(n7829), .Z(n10608) );
  XNOR U11336 ( .A(n11669), .B(n10139), .Z(n7829) );
  ANDN U11337 ( .B(n10495), .A(n10494), .Z(n11668) );
  XOR U11338 ( .A(n11670), .B(n10925), .Z(n10494) );
  XOR U11339 ( .A(n11673), .B(n10113), .Z(n7822) );
  AND U11340 ( .A(n10505), .B(n10503), .Z(n11672) );
  XOR U11341 ( .A(n11674), .B(n11675), .Z(n10503) );
  XOR U11342 ( .A(n11676), .B(n9190), .Z(n10505) );
  XOR U11343 ( .A(n11677), .B(n11678), .Z(n9190) );
  XNOR U11344 ( .A(n11679), .B(n7833), .Z(n4210) );
  XNOR U11345 ( .A(n11680), .B(n11639), .Z(n7833) );
  XNOR U11346 ( .A(n11681), .B(n10632), .Z(n10500) );
  XNOR U11347 ( .A(n11682), .B(n10431), .Z(n10632) );
  ANDN U11348 ( .B(n11500), .A(n11498), .Z(n11681) );
  XNOR U11349 ( .A(n11683), .B(n11684), .Z(n11498) );
  XNOR U11350 ( .A(n11687), .B(n4165), .Z(out[100]) );
  XNOR U11351 ( .A(n6972), .B(n2569), .Z(n4165) );
  XNOR U11352 ( .A(n8021), .B(n10928), .Z(n2569) );
  XNOR U11353 ( .A(n11688), .B(n11689), .Z(n10928) );
  XOR U11354 ( .A(n5678), .B(n5375), .Z(n11689) );
  XOR U11355 ( .A(n11690), .B(n8100), .Z(n5375) );
  XOR U11356 ( .A(n11691), .B(n11692), .Z(n8100) );
  ANDN U11357 ( .B(n8162), .A(n6988), .Z(n11690) );
  XOR U11358 ( .A(n11693), .B(n11162), .Z(n6988) );
  XNOR U11359 ( .A(n11694), .B(n11695), .Z(n8162) );
  XOR U11360 ( .A(n11696), .B(n6998), .Z(n5678) );
  XNOR U11361 ( .A(n11697), .B(n11550), .Z(n6998) );
  ANDN U11362 ( .B(n10834), .A(n6997), .Z(n11696) );
  XNOR U11363 ( .A(n11698), .B(n10565), .Z(n6997) );
  XOR U11364 ( .A(n11566), .B(n11699), .Z(n10834) );
  XOR U11365 ( .A(n6982), .B(n11700), .Z(n11688) );
  XNOR U11366 ( .A(n2233), .B(n3347), .Z(n11700) );
  XNOR U11367 ( .A(n11701), .B(n7006), .Z(n3347) );
  XNOR U11368 ( .A(n11702), .B(n9907), .Z(n7006) );
  AND U11369 ( .A(n8155), .B(n8154), .Z(n11701) );
  XNOR U11370 ( .A(n11703), .B(n10478), .Z(n8154) );
  XNOR U11371 ( .A(n11704), .B(n9551), .Z(n8155) );
  XOR U11372 ( .A(n11705), .B(n6993), .Z(n2233) );
  XNOR U11373 ( .A(n11706), .B(n10794), .Z(n6993) );
  ANDN U11374 ( .B(n8158), .A(n6992), .Z(n11705) );
  XOR U11375 ( .A(n11707), .B(n11656), .Z(n6992) );
  XNOR U11376 ( .A(n11708), .B(n11709), .Z(n8158) );
  XNOR U11377 ( .A(n11710), .B(n7001), .Z(n6982) );
  XNOR U11378 ( .A(n11711), .B(n11712), .Z(n7001) );
  AND U11379 ( .A(n7002), .B(n10820), .Z(n11710) );
  XNOR U11380 ( .A(n11713), .B(n10249), .Z(n10820) );
  XOR U11381 ( .A(n11714), .B(n11715), .Z(n7002) );
  XOR U11382 ( .A(n11716), .B(n11717), .Z(n8021) );
  XOR U11383 ( .A(n4338), .B(n2184), .Z(n11717) );
  XNOR U11384 ( .A(n11718), .B(n8083), .Z(n2184) );
  XOR U11385 ( .A(n11719), .B(n11550), .Z(n8083) );
  AND U11386 ( .A(n10721), .B(n10810), .Z(n11718) );
  XOR U11387 ( .A(n11720), .B(n8075), .Z(n4338) );
  XOR U11388 ( .A(n10227), .B(n11721), .Z(n8075) );
  AND U11389 ( .A(n6978), .B(n10800), .Z(n11720) );
  IV U11390 ( .A(n6979), .Z(n10800) );
  XOR U11391 ( .A(n11722), .B(n9784), .Z(n6979) );
  XNOR U11392 ( .A(n11723), .B(n9782), .Z(n6978) );
  XOR U11393 ( .A(n5965), .B(n11724), .Z(n11716) );
  XNOR U11394 ( .A(n5514), .B(n3761), .Z(n11724) );
  XNOR U11395 ( .A(n11725), .B(n8079), .Z(n3761) );
  XOR U11396 ( .A(n11726), .B(n10017), .Z(n8079) );
  ANDN U11397 ( .B(n6968), .A(n6970), .Z(n11725) );
  XOR U11398 ( .A(n10692), .B(n11727), .Z(n6970) );
  XNOR U11399 ( .A(n11728), .B(n11373), .Z(n6968) );
  XOR U11400 ( .A(n11729), .B(n10727), .Z(n5514) );
  XOR U11401 ( .A(n11730), .B(n9906), .Z(n10727) );
  ANDN U11402 ( .B(n10797), .A(n6974), .Z(n11729) );
  XNOR U11403 ( .A(n11731), .B(n10203), .Z(n6974) );
  IV U11404 ( .A(n6976), .Z(n10797) );
  XOR U11405 ( .A(n11732), .B(n10594), .Z(n6976) );
  XOR U11406 ( .A(n11733), .B(n8085), .Z(n5965) );
  XOR U11407 ( .A(n11734), .B(n10096), .Z(n8085) );
  NOR U11408 ( .A(n6964), .B(n6966), .Z(n11733) );
  XNOR U11409 ( .A(n11735), .B(n9922), .Z(n6966) );
  XNOR U11410 ( .A(n11736), .B(n11175), .Z(n6964) );
  XOR U11411 ( .A(n11737), .B(n10721), .Z(n6972) );
  XOR U11412 ( .A(n9535), .B(n11738), .Z(n10721) );
  ANDN U11413 ( .B(n8081), .A(n10810), .Z(n11737) );
  XNOR U11414 ( .A(n11739), .B(n10174), .Z(n10810) );
  IV U11415 ( .A(n10811), .Z(n8081) );
  XOR U11416 ( .A(n11740), .B(n11639), .Z(n10811) );
  ANDN U11417 ( .B(n3622), .A(n3620), .Z(n11687) );
  XNOR U11418 ( .A(n7532), .B(n2411), .Z(n3620) );
  XNOR U11419 ( .A(n10177), .B(n10983), .Z(n2411) );
  XNOR U11420 ( .A(n11741), .B(n11742), .Z(n10983) );
  XOR U11421 ( .A(n5392), .B(n3848), .Z(n11742) );
  XOR U11422 ( .A(n11743), .B(n11112), .Z(n3848) );
  XNOR U11423 ( .A(n11744), .B(n10296), .Z(n11112) );
  ANDN U11424 ( .B(n7544), .A(n7545), .Z(n11743) );
  XNOR U11425 ( .A(n11745), .B(n9406), .Z(n7545) );
  XNOR U11426 ( .A(n11746), .B(n11747), .Z(n7544) );
  XNOR U11427 ( .A(n11748), .B(n9970), .Z(n5392) );
  XNOR U11428 ( .A(n9097), .B(n11749), .Z(n9970) );
  XOR U11429 ( .A(n11750), .B(n11751), .Z(n9097) );
  AND U11430 ( .A(n7540), .B(n10412), .Z(n11748) );
  XOR U11431 ( .A(n9564), .B(n11752), .Z(n10412) );
  XOR U11432 ( .A(n11753), .B(n11754), .Z(n9564) );
  XOR U11433 ( .A(n11755), .B(n10134), .Z(n7540) );
  XNOR U11434 ( .A(n11756), .B(n11757), .Z(n10134) );
  XOR U11435 ( .A(n6188), .B(n11758), .Z(n11741) );
  XOR U11436 ( .A(n2279), .B(n5084), .Z(n11758) );
  XNOR U11437 ( .A(n11759), .B(n9982), .Z(n5084) );
  XOR U11438 ( .A(n11760), .B(n11761), .Z(n9982) );
  ANDN U11439 ( .B(n8593), .A(n8594), .Z(n11759) );
  XNOR U11440 ( .A(n11762), .B(n9773), .Z(n8594) );
  XOR U11441 ( .A(n11763), .B(n10019), .Z(n8593) );
  XNOR U11442 ( .A(n11764), .B(n9973), .Z(n2279) );
  XOR U11443 ( .A(n11765), .B(n11766), .Z(n9973) );
  AND U11444 ( .A(n9974), .B(n10414), .Z(n11764) );
  XOR U11445 ( .A(n11767), .B(n9979), .Z(n6188) );
  XOR U11446 ( .A(n11768), .B(n11769), .Z(n9979) );
  ANDN U11447 ( .B(n7534), .A(n7535), .Z(n11767) );
  XOR U11448 ( .A(n11770), .B(n10139), .Z(n7535) );
  XNOR U11449 ( .A(n9488), .B(n11771), .Z(n7534) );
  XOR U11450 ( .A(n11772), .B(n11773), .Z(n10177) );
  XNOR U11451 ( .A(n3413), .B(n5011), .Z(n11773) );
  XOR U11452 ( .A(n11774), .B(n7608), .Z(n5011) );
  XOR U11453 ( .A(n11775), .B(n10043), .Z(n7608) );
  AND U11454 ( .A(n10080), .B(n11264), .Z(n11774) );
  XNOR U11455 ( .A(n11776), .B(n10172), .Z(n11264) );
  XNOR U11456 ( .A(n11777), .B(n11778), .Z(n10080) );
  XOR U11457 ( .A(n11779), .B(n8652), .Z(n3413) );
  XOR U11458 ( .A(n11780), .B(n9769), .Z(n8652) );
  AND U11459 ( .A(n10083), .B(n11255), .Z(n11779) );
  XNOR U11460 ( .A(n11781), .B(n11782), .Z(n11255) );
  XNOR U11461 ( .A(n11783), .B(n10461), .Z(n10083) );
  IV U11462 ( .A(n9602), .Z(n10461) );
  XOR U11463 ( .A(n2383), .B(n11784), .Z(n11772) );
  XOR U11464 ( .A(n7601), .B(n3959), .Z(n11784) );
  XNOR U11465 ( .A(n11785), .B(n7622), .Z(n3959) );
  XOR U11466 ( .A(n11786), .B(n9676), .Z(n7622) );
  NOR U11467 ( .A(n7621), .B(n10072), .Z(n11785) );
  XNOR U11468 ( .A(n11787), .B(n10565), .Z(n10072) );
  XNOR U11469 ( .A(n11788), .B(n9694), .Z(n7621) );
  XOR U11470 ( .A(n11791), .B(n7617), .Z(n7601) );
  XOR U11471 ( .A(n11792), .B(n11793), .Z(n7617) );
  AND U11472 ( .A(n10075), .B(n7618), .Z(n11791) );
  XNOR U11473 ( .A(n11032), .B(n11794), .Z(n7618) );
  IV U11474 ( .A(n9083), .Z(n11032) );
  XNOR U11475 ( .A(n11401), .B(n11795), .Z(n10075) );
  XNOR U11476 ( .A(n11796), .B(n7614), .Z(n2383) );
  XNOR U11477 ( .A(n9537), .B(n11797), .Z(n7614) );
  ANDN U11478 ( .B(n7613), .A(n11267), .Z(n11796) );
  XNOR U11479 ( .A(n11798), .B(n10010), .Z(n11267) );
  XNOR U11480 ( .A(n11799), .B(n11466), .Z(n7613) );
  XOR U11481 ( .A(n11800), .B(n9974), .Z(n7532) );
  XNOR U11482 ( .A(n9398), .B(n11801), .Z(n9974) );
  IV U11483 ( .A(n9792), .Z(n9398) );
  XOR U11484 ( .A(n11802), .B(n11803), .Z(n9792) );
  NOR U11485 ( .A(n10414), .B(n10415), .Z(n11800) );
  XOR U11486 ( .A(n11804), .B(n10691), .Z(n10415) );
  XOR U11487 ( .A(n11805), .B(n9917), .Z(n10414) );
  XNOR U11488 ( .A(n3398), .B(n9730), .Z(n3622) );
  XNOR U11489 ( .A(n11806), .B(n10526), .Z(n9730) );
  ANDN U11490 ( .B(n9631), .A(n10659), .Z(n11806) );
  XNOR U11491 ( .A(n11807), .B(n10307), .Z(n9631) );
  XOR U11492 ( .A(n6162), .B(n10763), .Z(n3398) );
  XOR U11493 ( .A(n11808), .B(n11809), .Z(n10763) );
  XNOR U11494 ( .A(n1663), .B(n9825), .Z(n11809) );
  XOR U11495 ( .A(n11810), .B(n7314), .Z(n9825) );
  XNOR U11496 ( .A(n10110), .B(n11811), .Z(n7314) );
  AND U11497 ( .A(n9743), .B(n9742), .Z(n11810) );
  XNOR U11498 ( .A(n11538), .B(n11812), .Z(n9742) );
  XNOR U11499 ( .A(n11813), .B(n10200), .Z(n9743) );
  XOR U11500 ( .A(n11814), .B(n7307), .Z(n1663) );
  XOR U11501 ( .A(n11815), .B(n9820), .Z(n7307) );
  ANDN U11502 ( .B(n9751), .A(n9750), .Z(n11814) );
  XNOR U11503 ( .A(n10730), .B(n11816), .Z(n9750) );
  XOR U11504 ( .A(n11817), .B(n10681), .Z(n9751) );
  XNOR U11505 ( .A(n3725), .B(n11818), .Z(n11808) );
  XOR U11506 ( .A(n5072), .B(n4188), .Z(n11818) );
  XOR U11507 ( .A(n11819), .B(n7318), .Z(n4188) );
  XNOR U11508 ( .A(n10772), .B(n11820), .Z(n7318) );
  ANDN U11509 ( .B(n10639), .A(n9834), .Z(n11819) );
  XOR U11510 ( .A(n11822), .B(n10139), .Z(n10639) );
  XNOR U11511 ( .A(n11823), .B(n8343), .Z(n5072) );
  XOR U11512 ( .A(n11824), .B(n11825), .Z(n8343) );
  XOR U11513 ( .A(n9576), .B(n11826), .Z(n9745) );
  XNOR U11514 ( .A(n11686), .B(n11827), .Z(n9746) );
  XOR U11515 ( .A(n11828), .B(n8565), .Z(n3725) );
  XNOR U11516 ( .A(n11829), .B(n10265), .Z(n8565) );
  AND U11517 ( .A(n9754), .B(n9753), .Z(n11828) );
  XOR U11518 ( .A(n11830), .B(n10903), .Z(n9753) );
  XNOR U11519 ( .A(n10922), .B(n11831), .Z(n9754) );
  XOR U11520 ( .A(n11832), .B(n11833), .Z(n6162) );
  XNOR U11521 ( .A(n3182), .B(n7942), .Z(n11833) );
  XOR U11522 ( .A(n11834), .B(n9646), .Z(n7942) );
  IV U11523 ( .A(n10533), .Z(n9646) );
  XOR U11524 ( .A(n11835), .B(n9370), .Z(n10533) );
  ANDN U11525 ( .B(n10677), .A(n9737), .Z(n11834) );
  XOR U11526 ( .A(n11836), .B(n11837), .Z(n9737) );
  IV U11527 ( .A(n9738), .Z(n10677) );
  XNOR U11528 ( .A(n11838), .B(n10121), .Z(n9738) );
  XNOR U11529 ( .A(n11839), .B(n9643), .Z(n3182) );
  XOR U11530 ( .A(n11663), .B(n11840), .Z(n9643) );
  XNOR U11531 ( .A(n11841), .B(n11842), .Z(n9726) );
  XNOR U11532 ( .A(n11843), .B(n9584), .Z(n9725) );
  XNOR U11533 ( .A(n11844), .B(n11845), .Z(n9584) );
  XOR U11534 ( .A(n5476), .B(n11846), .Z(n11832) );
  XOR U11535 ( .A(n8288), .B(n2380), .Z(n11846) );
  XOR U11536 ( .A(n11847), .B(n9633), .Z(n2380) );
  IV U11537 ( .A(n10527), .Z(n9633) );
  XOR U11538 ( .A(n11848), .B(n9782), .Z(n10527) );
  XNOR U11539 ( .A(n11849), .B(n11850), .Z(n9782) );
  ANDN U11540 ( .B(n10659), .A(n10526), .Z(n11847) );
  XNOR U11541 ( .A(n11851), .B(n10037), .Z(n10526) );
  XNOR U11542 ( .A(n11852), .B(n11853), .Z(n10037) );
  XNOR U11543 ( .A(n11854), .B(n11855), .Z(n10659) );
  XOR U11544 ( .A(n11856), .B(n10530), .Z(n8288) );
  IV U11545 ( .A(n9637), .Z(n10530) );
  XNOR U11546 ( .A(n11857), .B(n9661), .Z(n9637) );
  ANDN U11547 ( .B(n10670), .A(n9728), .Z(n11856) );
  XOR U11548 ( .A(n11858), .B(n11859), .Z(n9728) );
  IV U11549 ( .A(n9729), .Z(n10670) );
  XNOR U11550 ( .A(n11649), .B(n11860), .Z(n9729) );
  XNOR U11551 ( .A(n11861), .B(n10524), .Z(n5476) );
  XNOR U11552 ( .A(n11396), .B(n11862), .Z(n10524) );
  XOR U11553 ( .A(n11002), .B(n11863), .Z(n9733) );
  IV U11554 ( .A(n9735), .Z(n10668) );
  XOR U11555 ( .A(n11864), .B(n10817), .Z(n9735) );
  IV U11556 ( .A(n9906), .Z(n10817) );
  XOR U11557 ( .A(n11865), .B(n11866), .Z(n9906) );
  XOR U11558 ( .A(n11867), .B(n6129), .Z(out[1009]) );
  IV U11559 ( .A(n6766), .Z(n6129) );
  XNOR U11560 ( .A(n8526), .B(n2240), .Z(n6766) );
  XNOR U11561 ( .A(n6011), .B(n6088), .Z(n2240) );
  XNOR U11562 ( .A(n11868), .B(n11869), .Z(n6088) );
  XOR U11563 ( .A(n2276), .B(n5403), .Z(n11869) );
  XOR U11564 ( .A(n11870), .B(n7327), .Z(n5403) );
  XNOR U11565 ( .A(n9535), .B(n11871), .Z(n7327) );
  IV U11566 ( .A(n11872), .Z(n9535) );
  ANDN U11567 ( .B(n8537), .A(n7326), .Z(n11870) );
  XOR U11568 ( .A(n11873), .B(n9803), .Z(n7326) );
  XNOR U11569 ( .A(n11874), .B(n11875), .Z(n8537) );
  XNOR U11570 ( .A(n11876), .B(n7330), .Z(n2276) );
  XNOR U11571 ( .A(n11877), .B(n11878), .Z(n7330) );
  ANDN U11572 ( .B(n7331), .A(n8532), .Z(n11876) );
  XNOR U11573 ( .A(n11879), .B(n11880), .Z(n8532) );
  XOR U11574 ( .A(n11881), .B(n11882), .Z(n7331) );
  XNOR U11575 ( .A(n3123), .B(n11883), .Z(n11868) );
  XNOR U11576 ( .A(n5843), .B(n7320), .Z(n11883) );
  XNOR U11577 ( .A(n11884), .B(n8445), .Z(n7320) );
  XNOR U11578 ( .A(n11885), .B(n11072), .Z(n8445) );
  ANDN U11579 ( .B(n7336), .A(n8535), .Z(n11884) );
  XOR U11580 ( .A(n11886), .B(n10995), .Z(n8535) );
  XNOR U11581 ( .A(n11887), .B(n11888), .Z(n7336) );
  XNOR U11582 ( .A(n11889), .B(n7339), .Z(n5843) );
  XOR U11583 ( .A(n11890), .B(n11891), .Z(n7339) );
  AND U11584 ( .A(n11597), .B(n7340), .Z(n11889) );
  XNOR U11585 ( .A(n11892), .B(n7344), .Z(n3123) );
  XOR U11586 ( .A(n11893), .B(n11894), .Z(n7344) );
  NOR U11587 ( .A(n8528), .B(n7343), .Z(n11892) );
  XNOR U11588 ( .A(n11895), .B(n11896), .Z(n7343) );
  XNOR U11589 ( .A(n9377), .B(n11897), .Z(n8528) );
  IV U11590 ( .A(n10118), .Z(n9377) );
  XOR U11591 ( .A(n11898), .B(n11899), .Z(n6011) );
  XOR U11592 ( .A(n5218), .B(n1905), .Z(n11899) );
  XNOR U11593 ( .A(n11900), .B(n8640), .Z(n1905) );
  AND U11594 ( .A(n7419), .B(n8515), .Z(n11900) );
  XOR U11595 ( .A(n9219), .B(n11901), .Z(n8515) );
  IV U11596 ( .A(n9673), .Z(n9219) );
  XOR U11597 ( .A(n11902), .B(n11903), .Z(n9673) );
  XNOR U11598 ( .A(n11904), .B(n11905), .Z(n7419) );
  XNOR U11599 ( .A(n11906), .B(n8645), .Z(n5218) );
  NOR U11600 ( .A(n7411), .B(n8513), .Z(n11906) );
  XOR U11601 ( .A(n11907), .B(n11908), .Z(n8513) );
  XOR U11602 ( .A(n11909), .B(n10307), .Z(n7411) );
  XNOR U11603 ( .A(n3657), .B(n11910), .Z(n11898) );
  XOR U11604 ( .A(n8622), .B(n4141), .Z(n11910) );
  XNOR U11605 ( .A(n11911), .B(n8647), .Z(n4141) );
  ANDN U11606 ( .B(n7402), .A(n8523), .Z(n11911) );
  XOR U11607 ( .A(n11912), .B(n9676), .Z(n8523) );
  XOR U11608 ( .A(n11913), .B(n11914), .Z(n9676) );
  XNOR U11609 ( .A(n11915), .B(n11916), .Z(n7402) );
  XOR U11610 ( .A(n11917), .B(n8643), .Z(n8622) );
  IV U11611 ( .A(n11918), .Z(n8643) );
  ANDN U11612 ( .B(n8519), .A(n7406), .Z(n11917) );
  XNOR U11613 ( .A(n11919), .B(n9587), .Z(n7406) );
  XNOR U11614 ( .A(n10044), .B(n11920), .Z(n8519) );
  XNOR U11615 ( .A(n11921), .B(n11922), .Z(n3657) );
  ANDN U11616 ( .B(n8521), .A(n7415), .Z(n11921) );
  XOR U11617 ( .A(n11924), .B(n7340), .Z(n8526) );
  XNOR U11618 ( .A(n11925), .B(n10373), .Z(n7340) );
  NOR U11619 ( .A(n8452), .B(n11597), .Z(n11924) );
  XNOR U11620 ( .A(n11926), .B(n11927), .Z(n11597) );
  XNOR U11621 ( .A(n11928), .B(n10716), .Z(n8452) );
  IV U11622 ( .A(n11905), .Z(n10716) );
  XOR U11623 ( .A(n11929), .B(n11930), .Z(n11905) );
  AND U11624 ( .A(n5619), .B(n5621), .Z(n11867) );
  XOR U11625 ( .A(n10617), .B(n5346), .Z(n5621) );
  XOR U11626 ( .A(n7813), .B(n8969), .Z(n5346) );
  XNOR U11627 ( .A(n11931), .B(n11932), .Z(n8969) );
  XNOR U11628 ( .A(n5425), .B(n3875), .Z(n11932) );
  XOR U11629 ( .A(n11933), .B(n11934), .Z(n3875) );
  ANDN U11630 ( .B(n7990), .A(n7988), .Z(n11933) );
  XOR U11631 ( .A(n11935), .B(n11936), .Z(n7990) );
  XOR U11632 ( .A(n11937), .B(n10738), .Z(n5425) );
  AND U11633 ( .A(n7984), .B(n10868), .Z(n11937) );
  XNOR U11634 ( .A(n11938), .B(n10136), .Z(n10868) );
  XOR U11635 ( .A(n11715), .B(n11939), .Z(n7984) );
  XOR U11636 ( .A(n6216), .B(n11940), .Z(n11931) );
  XNOR U11637 ( .A(n2325), .B(n5263), .Z(n11940) );
  XNOR U11638 ( .A(n11941), .B(n10749), .Z(n5263) );
  AND U11639 ( .A(n8972), .B(n10750), .Z(n11941) );
  XOR U11640 ( .A(n9083), .B(n11942), .Z(n10750) );
  XNOR U11641 ( .A(n11944), .B(n11945), .Z(n11754) );
  XNOR U11642 ( .A(n10029), .B(n11073), .Z(n11945) );
  XOR U11643 ( .A(n11946), .B(n11947), .Z(n11073) );
  NOR U11644 ( .A(n11948), .B(n11949), .Z(n11946) );
  XNOR U11645 ( .A(n11950), .B(n11951), .Z(n10029) );
  NOR U11646 ( .A(n11952), .B(n11953), .Z(n11950) );
  XOR U11647 ( .A(n10878), .B(n11954), .Z(n11944) );
  XOR U11648 ( .A(n10906), .B(n11029), .Z(n11954) );
  XNOR U11649 ( .A(n11955), .B(n11956), .Z(n11029) );
  NOR U11650 ( .A(n11957), .B(n11958), .Z(n11955) );
  XNOR U11651 ( .A(n11959), .B(n11960), .Z(n10906) );
  AND U11652 ( .A(n11961), .B(n11962), .Z(n11959) );
  XNOR U11653 ( .A(n11963), .B(n11964), .Z(n10878) );
  NOR U11654 ( .A(n11965), .B(n11966), .Z(n11963) );
  XNOR U11655 ( .A(n10266), .B(n11967), .Z(n8972) );
  XNOR U11656 ( .A(n11968), .B(n10741), .Z(n2325) );
  AND U11657 ( .A(n7974), .B(n7976), .Z(n11968) );
  XOR U11658 ( .A(n11969), .B(n9261), .Z(n7976) );
  XNOR U11659 ( .A(n11970), .B(n11971), .Z(n7974) );
  XNOR U11660 ( .A(n11972), .B(n10746), .Z(n6216) );
  AND U11661 ( .A(n7980), .B(n7978), .Z(n11972) );
  XOR U11662 ( .A(n11973), .B(n10025), .Z(n7978) );
  XNOR U11663 ( .A(n11974), .B(n11550), .Z(n7980) );
  XOR U11664 ( .A(n11975), .B(n11976), .Z(n7813) );
  XNOR U11665 ( .A(n3765), .B(n5097), .Z(n11976) );
  XOR U11666 ( .A(n11977), .B(n8910), .Z(n5097) );
  IV U11667 ( .A(n10756), .Z(n8910) );
  XOR U11668 ( .A(n11978), .B(n11979), .Z(n10756) );
  NOR U11669 ( .A(n10623), .B(n10624), .Z(n11977) );
  XNOR U11670 ( .A(n9170), .B(n11980), .Z(n10624) );
  XOR U11671 ( .A(n11981), .B(n11971), .Z(n10623) );
  XOR U11672 ( .A(n11982), .B(n7867), .Z(n3765) );
  XOR U11673 ( .A(n9516), .B(n11983), .Z(n7867) );
  AND U11674 ( .A(n11645), .B(n10615), .Z(n11982) );
  XNOR U11675 ( .A(n9354), .B(n11984), .Z(n10615) );
  IV U11676 ( .A(n10616), .Z(n11645) );
  XNOR U11677 ( .A(n11985), .B(n9176), .Z(n10616) );
  XOR U11678 ( .A(n4216), .B(n11986), .Z(n11975) );
  XOR U11679 ( .A(n1702), .B(n10733), .Z(n11986) );
  XOR U11680 ( .A(n11987), .B(n7877), .Z(n10733) );
  XNOR U11681 ( .A(n11988), .B(n10043), .Z(n7877) );
  XNOR U11682 ( .A(n11989), .B(n11990), .Z(n10043) );
  AND U11683 ( .A(n10613), .B(n10612), .Z(n11987) );
  IV U11684 ( .A(n10762), .Z(n10612) );
  XOR U11685 ( .A(n11991), .B(n11015), .Z(n10762) );
  XNOR U11686 ( .A(n9608), .B(n11992), .Z(n10613) );
  IV U11687 ( .A(n11993), .Z(n9608) );
  XOR U11688 ( .A(n11994), .B(n7870), .Z(n1702) );
  IV U11689 ( .A(n10754), .Z(n7870) );
  XOR U11690 ( .A(n11995), .B(n10256), .Z(n10754) );
  ANDN U11691 ( .B(n10621), .A(n10620), .Z(n11994) );
  XNOR U11692 ( .A(n11926), .B(n11996), .Z(n10620) );
  XNOR U11693 ( .A(n11997), .B(n11666), .Z(n10621) );
  XOR U11694 ( .A(n11998), .B(n7881), .Z(n4216) );
  XNOR U11695 ( .A(n11999), .B(n12000), .Z(n7881) );
  NOR U11696 ( .A(n11634), .B(n10759), .Z(n11998) );
  XNOR U11697 ( .A(n12001), .B(n10759), .Z(n10617) );
  XNOR U11698 ( .A(n9108), .B(n12002), .Z(n10759) );
  AND U11699 ( .A(n7879), .B(n11634), .Z(n12001) );
  XNOR U11700 ( .A(n12003), .B(n10938), .Z(n11634) );
  XOR U11701 ( .A(n10912), .B(n12004), .Z(n7879) );
  IV U11702 ( .A(n12005), .Z(n10912) );
  XNOR U11703 ( .A(n12006), .B(n3806), .Z(n5619) );
  IV U11704 ( .A(n1742), .Z(n3806) );
  XOR U11705 ( .A(n12007), .B(n12008), .Z(n9541) );
  XOR U11706 ( .A(n3445), .B(n5058), .Z(n12008) );
  XNOR U11707 ( .A(n12009), .B(n8355), .Z(n5058) );
  AND U11708 ( .A(n11625), .B(n12010), .Z(n12009) );
  XNOR U11709 ( .A(n12011), .B(n9654), .Z(n3445) );
  ANDN U11710 ( .B(n12012), .A(n11628), .Z(n12011) );
  XNOR U11711 ( .A(n4238), .B(n12013), .Z(n12007) );
  XNOR U11712 ( .A(n8344), .B(n2469), .Z(n12013) );
  XNOR U11713 ( .A(n12014), .B(n8364), .Z(n2469) );
  ANDN U11714 ( .B(n8365), .A(n12015), .Z(n12014) );
  XOR U11715 ( .A(n12016), .B(n8350), .Z(n8344) );
  AND U11716 ( .A(n11620), .B(n8351), .Z(n12016) );
  XNOR U11717 ( .A(n12017), .B(n8361), .Z(n4238) );
  ANDN U11718 ( .B(n11617), .A(n8360), .Z(n12017) );
  XNOR U11719 ( .A(n12018), .B(n12019), .Z(n6251) );
  XNOR U11720 ( .A(n5391), .B(n3637), .Z(n12019) );
  XOR U11721 ( .A(n12020), .B(n12021), .Z(n3637) );
  XNOR U11722 ( .A(n12023), .B(n12024), .Z(n5391) );
  ANDN U11723 ( .B(n8403), .A(n12025), .Z(n12023) );
  XNOR U11724 ( .A(n12026), .B(n12027), .Z(n12018) );
  XNOR U11725 ( .A(n2091), .B(n4271), .Z(n12027) );
  XOR U11726 ( .A(n12028), .B(n12029), .Z(n4271) );
  AND U11727 ( .A(n8407), .B(n12030), .Z(n12028) );
  XOR U11728 ( .A(n12031), .B(n12032), .Z(n2091) );
  AND U11729 ( .A(n12033), .B(n12034), .Z(n12031) );
  XOR U11730 ( .A(n12035), .B(n6134), .Z(out[1008]) );
  IV U11731 ( .A(n6795), .Z(n6134) );
  XOR U11732 ( .A(n8638), .B(n2247), .Z(n6795) );
  XNOR U11733 ( .A(n6016), .B(n6093), .Z(n2247) );
  XNOR U11734 ( .A(n12036), .B(n12037), .Z(n6093) );
  XOR U11735 ( .A(n2283), .B(n5408), .Z(n12037) );
  XOR U11736 ( .A(n12038), .B(n7404), .Z(n5408) );
  XNOR U11737 ( .A(n9605), .B(n12039), .Z(n7404) );
  AND U11738 ( .A(n7403), .B(n8647), .Z(n12038) );
  XNOR U11739 ( .A(n12040), .B(n9388), .Z(n8647) );
  XNOR U11740 ( .A(n12041), .B(n9927), .Z(n7403) );
  XNOR U11741 ( .A(n12042), .B(n7408), .Z(n2283) );
  XNOR U11742 ( .A(n12043), .B(n11875), .Z(n7408) );
  AND U11743 ( .A(n7407), .B(n11918), .Z(n12042) );
  XOR U11744 ( .A(n10827), .B(n12044), .Z(n11918) );
  XNOR U11745 ( .A(n12045), .B(n9524), .Z(n7407) );
  XNOR U11746 ( .A(n3131), .B(n12046), .Z(n12036) );
  XOR U11747 ( .A(n5898), .B(n7397), .Z(n12046) );
  XNOR U11748 ( .A(n12047), .B(n7412), .Z(n7397) );
  XNOR U11749 ( .A(n11777), .B(n12048), .Z(n7412) );
  AND U11750 ( .A(n8645), .B(n7413), .Z(n12047) );
  XOR U11751 ( .A(n12049), .B(n12050), .Z(n7413) );
  XNOR U11752 ( .A(n12051), .B(n11766), .Z(n8645) );
  XNOR U11753 ( .A(n12052), .B(n7417), .Z(n5898) );
  XOR U11754 ( .A(n12053), .B(n11586), .Z(n7417) );
  ANDN U11755 ( .B(n11922), .A(n7416), .Z(n12052) );
  XNOR U11756 ( .A(n12054), .B(n8516), .Z(n3131) );
  XOR U11757 ( .A(n12055), .B(n12056), .Z(n8516) );
  ANDN U11758 ( .B(n8640), .A(n7420), .Z(n12054) );
  XOR U11759 ( .A(n12057), .B(n12058), .Z(n7420) );
  XNOR U11760 ( .A(n9511), .B(n12059), .Z(n8640) );
  XOR U11761 ( .A(n12060), .B(n12061), .Z(n6016) );
  XNOR U11762 ( .A(n5221), .B(n1913), .Z(n12061) );
  XOR U11763 ( .A(n12062), .B(n8705), .Z(n1913) );
  IV U11764 ( .A(n12063), .Z(n8705) );
  ANDN U11765 ( .B(n8628), .A(n7493), .Z(n12062) );
  XNOR U11766 ( .A(n12064), .B(n12065), .Z(n7493) );
  XNOR U11767 ( .A(n12066), .B(n10875), .Z(n8628) );
  XOR U11768 ( .A(n12067), .B(n8710), .Z(n5221) );
  NOR U11769 ( .A(n7485), .B(n8626), .Z(n12067) );
  XOR U11770 ( .A(n12068), .B(n12069), .Z(n8626) );
  XNOR U11771 ( .A(n11538), .B(n12070), .Z(n7485) );
  XOR U11772 ( .A(n3661), .B(n12071), .Z(n12060) );
  XOR U11773 ( .A(n8686), .B(n4145), .Z(n12071) );
  XNOR U11774 ( .A(n12072), .B(n8712), .Z(n4145) );
  ANDN U11775 ( .B(n8635), .A(n7476), .Z(n12072) );
  XNOR U11776 ( .A(n12073), .B(n12074), .Z(n7476) );
  XOR U11777 ( .A(n12075), .B(n9784), .Z(n8635) );
  XOR U11778 ( .A(n12078), .B(n8708), .Z(n8686) );
  IV U11779 ( .A(n12079), .Z(n8708) );
  ANDN U11780 ( .B(n8631), .A(n7480), .Z(n12078) );
  XNOR U11781 ( .A(n12080), .B(n9697), .Z(n7480) );
  XNOR U11782 ( .A(n9094), .B(n12081), .Z(n8631) );
  IV U11783 ( .A(n12082), .Z(n9094) );
  XOR U11784 ( .A(n12083), .B(n12084), .Z(n3661) );
  AND U11785 ( .A(n7489), .B(n8633), .Z(n12083) );
  IV U11786 ( .A(n12085), .Z(n8633) );
  XOR U11787 ( .A(n9907), .B(n12086), .Z(n7489) );
  IV U11788 ( .A(n11366), .Z(n9907) );
  XOR U11789 ( .A(n12087), .B(n7416), .Z(n8638) );
  XOR U11790 ( .A(n12088), .B(n11412), .Z(n7416) );
  NOR U11791 ( .A(n8521), .B(n11922), .Z(n12087) );
  XNOR U11792 ( .A(n9079), .B(n12089), .Z(n11922) );
  XOR U11793 ( .A(n12090), .B(n11639), .Z(n8521) );
  IV U11794 ( .A(n12065), .Z(n11639) );
  XOR U11795 ( .A(n12091), .B(n12092), .Z(n12065) );
  ANDN U11796 ( .B(n5625), .A(n5623), .Z(n12035) );
  XNOR U11797 ( .A(n12093), .B(n1747), .Z(n5623) );
  XOR U11798 ( .A(n12094), .B(n12095), .Z(n9649) );
  XOR U11799 ( .A(n3452), .B(n4826), .Z(n12095) );
  XNOR U11800 ( .A(n12096), .B(n8409), .Z(n4826) );
  NOR U11801 ( .A(n8408), .B(n12029), .Z(n12096) );
  XNOR U11802 ( .A(n12097), .B(n9761), .Z(n3452) );
  NOR U11803 ( .A(n12032), .B(n9760), .Z(n12097) );
  XOR U11804 ( .A(n4264), .B(n12098), .Z(n12094) );
  XNOR U11805 ( .A(n8399), .B(n2478), .Z(n12098) );
  XNOR U11806 ( .A(n12099), .B(n8419), .Z(n2478) );
  ANDN U11807 ( .B(n12100), .A(n12101), .Z(n12099) );
  XOR U11808 ( .A(n12102), .B(n8405), .Z(n8399) );
  ANDN U11809 ( .B(n12103), .A(n12024), .Z(n12102) );
  XOR U11810 ( .A(n12104), .B(n8414), .Z(n4264) );
  AND U11811 ( .A(n8415), .B(n12105), .Z(n12104) );
  XNOR U11812 ( .A(n12106), .B(n12107), .Z(n6255) );
  XOR U11813 ( .A(n5396), .B(n3643), .Z(n12107) );
  XOR U11814 ( .A(n12108), .B(n12109), .Z(n3643) );
  AND U11815 ( .A(n8486), .B(n12110), .Z(n12108) );
  XNOR U11816 ( .A(n12111), .B(n8428), .Z(n5396) );
  ANDN U11817 ( .B(n8476), .A(n8429), .Z(n12111) );
  IV U11818 ( .A(n12112), .Z(n8476) );
  XOR U11819 ( .A(n4273), .B(n12113), .Z(n12106) );
  XOR U11820 ( .A(n5830), .B(n2095), .Z(n12113) );
  XNOR U11821 ( .A(n12114), .B(n8424), .Z(n2095) );
  AND U11822 ( .A(n8425), .B(n9857), .Z(n12114) );
  IV U11823 ( .A(n12115), .Z(n9857) );
  XOR U11824 ( .A(n12116), .B(n8439), .Z(n5830) );
  ANDN U11825 ( .B(n12117), .A(n8490), .Z(n12116) );
  XOR U11826 ( .A(n12118), .B(n8434), .Z(n4273) );
  AND U11827 ( .A(n8480), .B(n8435), .Z(n12118) );
  XOR U11828 ( .A(n10742), .B(n2062), .Z(n5625) );
  XNOR U11829 ( .A(n7861), .B(n9030), .Z(n2062) );
  XNOR U11830 ( .A(n12119), .B(n12120), .Z(n9030) );
  XNOR U11831 ( .A(n5429), .B(n3554), .Z(n12120) );
  XOR U11832 ( .A(n12121), .B(n12122), .Z(n3554) );
  AND U11833 ( .A(n8061), .B(n12123), .Z(n12121) );
  XNOR U11834 ( .A(n12124), .B(n10712), .Z(n8061) );
  XNOR U11835 ( .A(n12125), .B(n10845), .Z(n5429) );
  AND U11836 ( .A(n8056), .B(n10846), .Z(n12125) );
  XOR U11837 ( .A(n11060), .B(n12126), .Z(n10846) );
  XOR U11838 ( .A(n12127), .B(n10281), .Z(n8056) );
  XOR U11839 ( .A(n6220), .B(n12128), .Z(n12119) );
  XOR U11840 ( .A(n2332), .B(n5316), .Z(n12128) );
  XNOR U11841 ( .A(n12129), .B(n10858), .Z(n5316) );
  AND U11842 ( .A(n9032), .B(n9034), .Z(n12129) );
  XOR U11843 ( .A(n12130), .B(n10455), .Z(n9034) );
  XOR U11844 ( .A(n12131), .B(n11162), .Z(n9032) );
  XNOR U11845 ( .A(n12132), .B(n12133), .Z(n2332) );
  ANDN U11846 ( .B(n8047), .A(n8045), .Z(n12132) );
  XOR U11847 ( .A(n12134), .B(n12135), .Z(n8045) );
  XNOR U11848 ( .A(n12136), .B(n12137), .Z(n8047) );
  XNOR U11849 ( .A(n12138), .B(n10855), .Z(n6220) );
  AND U11850 ( .A(n8051), .B(n8049), .Z(n12138) );
  IV U11851 ( .A(n10854), .Z(n8049) );
  XOR U11852 ( .A(n10909), .B(n12139), .Z(n10854) );
  XNOR U11853 ( .A(n12140), .B(n11684), .Z(n8051) );
  XOR U11854 ( .A(n12141), .B(n12142), .Z(n7861) );
  XNOR U11855 ( .A(n3769), .B(n5099), .Z(n12142) );
  XOR U11856 ( .A(n12143), .B(n8973), .Z(n5099) );
  XNOR U11857 ( .A(n9088), .B(n12144), .Z(n8973) );
  IV U11858 ( .A(n12145), .Z(n9088) );
  XOR U11859 ( .A(n12146), .B(n10061), .Z(n10748) );
  XOR U11860 ( .A(n12147), .B(n10215), .Z(n10749) );
  XNOR U11861 ( .A(n12148), .B(n7975), .Z(n3769) );
  XNOR U11862 ( .A(n12149), .B(n9587), .Z(n7975) );
  AND U11863 ( .A(n10741), .B(n10740), .Z(n12148) );
  XOR U11864 ( .A(n12150), .B(n9483), .Z(n10740) );
  XOR U11865 ( .A(n12151), .B(n10783), .Z(n10741) );
  XOR U11866 ( .A(n4239), .B(n12152), .Z(n12141) );
  XOR U11867 ( .A(n1706), .B(n10840), .Z(n12152) );
  XOR U11868 ( .A(n12153), .B(n7986), .Z(n10840) );
  XOR U11869 ( .A(n10154), .B(n12154), .Z(n7986) );
  AND U11870 ( .A(n10738), .B(n10737), .Z(n12153) );
  IV U11871 ( .A(n10869), .Z(n10737) );
  XOR U11872 ( .A(n12155), .B(n11747), .Z(n10869) );
  XOR U11873 ( .A(n12156), .B(n9718), .Z(n10738) );
  XNOR U11874 ( .A(n12157), .B(n7979), .Z(n1706) );
  XNOR U11875 ( .A(n12158), .B(n10386), .Z(n7979) );
  XOR U11876 ( .A(n9079), .B(n12159), .Z(n10745) );
  XOR U11877 ( .A(n9354), .B(n12160), .Z(n10746) );
  XNOR U11878 ( .A(n12161), .B(n12162), .Z(n9354) );
  XNOR U11879 ( .A(n12163), .B(n7989), .Z(n4239) );
  XNOR U11880 ( .A(n12164), .B(n12165), .Z(n7989) );
  XNOR U11881 ( .A(n12166), .B(n10865), .Z(n10742) );
  XNOR U11882 ( .A(n12167), .B(n9176), .Z(n10865) );
  ANDN U11883 ( .B(n7988), .A(n11934), .Z(n12166) );
  XNOR U11884 ( .A(n12168), .B(n11037), .Z(n11934) );
  XNOR U11885 ( .A(n12169), .B(n10991), .Z(n7988) );
  XOR U11886 ( .A(n12170), .B(n6139), .Z(out[1007]) );
  XNOR U11887 ( .A(n8703), .B(n2254), .Z(n6139) );
  XNOR U11888 ( .A(n6021), .B(n6098), .Z(n2254) );
  XNOR U11889 ( .A(n12171), .B(n12172), .Z(n6098) );
  XNOR U11890 ( .A(n2290), .B(n5411), .Z(n12172) );
  XOR U11891 ( .A(n12173), .B(n7478), .Z(n5411) );
  XOR U11892 ( .A(n12174), .B(n11842), .Z(n7478) );
  IV U11893 ( .A(n9716), .Z(n11842) );
  ANDN U11894 ( .B(n8712), .A(n7477), .Z(n12173) );
  XOR U11895 ( .A(n12175), .B(n12176), .Z(n7477) );
  XNOR U11896 ( .A(n12177), .B(n9519), .Z(n8712) );
  XNOR U11897 ( .A(n12178), .B(n7482), .Z(n2290) );
  XOR U11898 ( .A(n12179), .B(n9388), .Z(n7482) );
  AND U11899 ( .A(n7481), .B(n12079), .Z(n12178) );
  XNOR U11900 ( .A(n12180), .B(n10943), .Z(n12079) );
  XOR U11901 ( .A(n12181), .B(n9595), .Z(n7481) );
  XNOR U11902 ( .A(n3135), .B(n12182), .Z(n12171) );
  XOR U11903 ( .A(n5953), .B(n7471), .Z(n12182) );
  XNOR U11904 ( .A(n12183), .B(n7486), .Z(n7471) );
  XOR U11905 ( .A(n12184), .B(n11324), .Z(n7486) );
  ANDN U11906 ( .B(n7487), .A(n8710), .Z(n12183) );
  XOR U11907 ( .A(n11409), .B(n12185), .Z(n8710) );
  XOR U11908 ( .A(n12186), .B(n10235), .Z(n7487) );
  XNOR U11909 ( .A(n12187), .B(n7490), .Z(n5953) );
  XNOR U11910 ( .A(n12188), .B(n11908), .Z(n7490) );
  ANDN U11911 ( .B(n7491), .A(n12084), .Z(n12187) );
  XNOR U11912 ( .A(n12189), .B(n7494), .Z(n3135) );
  XOR U11913 ( .A(n12190), .B(n10254), .Z(n7494) );
  IV U11914 ( .A(n12191), .Z(n10254) );
  AND U11915 ( .A(n7495), .B(n12063), .Z(n12189) );
  XOR U11916 ( .A(n12192), .B(n9582), .Z(n12063) );
  XOR U11917 ( .A(n12193), .B(n12194), .Z(n7495) );
  XOR U11918 ( .A(n12195), .B(n12196), .Z(n6021) );
  XNOR U11919 ( .A(n5224), .B(n1918), .Z(n12196) );
  XOR U11920 ( .A(n12197), .B(n8739), .Z(n1918) );
  IV U11921 ( .A(n12198), .Z(n8739) );
  ANDN U11922 ( .B(n7570), .A(n8692), .Z(n12197) );
  XNOR U11923 ( .A(n12199), .B(n9904), .Z(n8692) );
  IV U11924 ( .A(n9406), .Z(n9904) );
  XNOR U11925 ( .A(n12200), .B(n12201), .Z(n9406) );
  XOR U11926 ( .A(n11999), .B(n12202), .Z(n7570) );
  XOR U11927 ( .A(n12203), .B(n8744), .Z(n5224) );
  NOR U11928 ( .A(n8690), .B(n7562), .Z(n12203) );
  XOR U11929 ( .A(n12204), .B(n10896), .Z(n7562) );
  XOR U11930 ( .A(n12205), .B(n12206), .Z(n8690) );
  XNOR U11931 ( .A(n3667), .B(n12207), .Z(n12195) );
  XNOR U11932 ( .A(n8720), .B(n4148), .Z(n12207) );
  XNOR U11933 ( .A(n12208), .B(n8746), .Z(n4148) );
  AND U11934 ( .A(n8699), .B(n8700), .Z(n12208) );
  IV U11935 ( .A(n7553), .Z(n8700) );
  XOR U11936 ( .A(n12209), .B(n12210), .Z(n7553) );
  XNOR U11937 ( .A(n11366), .B(n12211), .Z(n8699) );
  XOR U11938 ( .A(n12212), .B(n12213), .Z(n11366) );
  AND U11939 ( .A(n8695), .B(n7557), .Z(n12214) );
  XNOR U11940 ( .A(n12215), .B(n9803), .Z(n7557) );
  XNOR U11941 ( .A(n12216), .B(n9216), .Z(n8695) );
  XNOR U11942 ( .A(n12217), .B(n12218), .Z(n3667) );
  ANDN U11943 ( .B(n7566), .A(n8697), .Z(n12217) );
  XNOR U11944 ( .A(n11502), .B(n12219), .Z(n7566) );
  IV U11945 ( .A(n11045), .Z(n11502) );
  XOR U11946 ( .A(n12220), .B(n7491), .Z(n8703) );
  XOR U11947 ( .A(n12221), .B(n10675), .Z(n7491) );
  AND U11948 ( .A(n12084), .B(n12085), .Z(n12220) );
  XOR U11949 ( .A(n11999), .B(n12222), .Z(n12085) );
  IV U11950 ( .A(n11715), .Z(n11999) );
  XOR U11951 ( .A(n12223), .B(n12224), .Z(n11715) );
  XOR U11952 ( .A(n12225), .B(n9213), .Z(n12084) );
  NOR U11953 ( .A(n5628), .B(n5627), .Z(n12170) );
  XNOR U11954 ( .A(n8431), .B(n3818), .Z(n5627) );
  IV U11955 ( .A(n1752), .Z(n3818) );
  XNOR U11956 ( .A(n6264), .B(n9756), .Z(n1752) );
  XOR U11957 ( .A(n12226), .B(n12227), .Z(n9756) );
  XNOR U11958 ( .A(n3454), .B(n4830), .Z(n12227) );
  XOR U11959 ( .A(n12228), .B(n8481), .Z(n4830) );
  ANDN U11960 ( .B(n8482), .A(n8434), .Z(n12228) );
  XNOR U11961 ( .A(n12229), .B(n9768), .Z(n8434) );
  XOR U11962 ( .A(n12230), .B(n10675), .Z(n8482) );
  XNOR U11963 ( .A(n12231), .B(n9858), .Z(n3454) );
  AND U11964 ( .A(n8423), .B(n8424), .Z(n12231) );
  XNOR U11965 ( .A(n12232), .B(n11896), .Z(n8424) );
  XNOR U11966 ( .A(n9166), .B(n12233), .Z(n8423) );
  IV U11967 ( .A(n12234), .Z(n9166) );
  XNOR U11968 ( .A(n4290), .B(n12235), .Z(n12226) );
  XOR U11969 ( .A(n8472), .B(n2485), .Z(n12235) );
  XOR U11970 ( .A(n12236), .B(n8491), .Z(n2485) );
  AND U11971 ( .A(n8437), .B(n8439), .Z(n12236) );
  XOR U11972 ( .A(n12237), .B(n10025), .Z(n8439) );
  IV U11973 ( .A(n11825), .Z(n10025) );
  XOR U11974 ( .A(n12238), .B(n10382), .Z(n8437) );
  XOR U11975 ( .A(n12239), .B(n8477), .Z(n8472) );
  ANDN U11976 ( .B(n8478), .A(n8428), .Z(n12239) );
  XNOR U11977 ( .A(n12240), .B(n10455), .Z(n8428) );
  XOR U11978 ( .A(n12241), .B(n10590), .Z(n8478) );
  XNOR U11979 ( .A(n12242), .B(n8488), .Z(n4290) );
  ANDN U11980 ( .B(n8487), .A(n12109), .Z(n12242) );
  XNOR U11981 ( .A(n12243), .B(n12244), .Z(n6264) );
  XOR U11982 ( .A(n5402), .B(n3647), .Z(n12244) );
  XOR U11983 ( .A(n12245), .B(n12246), .Z(n3647) );
  ANDN U11984 ( .B(n6371), .A(n6372), .Z(n12245) );
  XOR U11985 ( .A(n12247), .B(n10382), .Z(n6372) );
  XOR U11986 ( .A(n12248), .B(n12249), .Z(n5402) );
  ANDN U11987 ( .B(n6362), .A(n6363), .Z(n12248) );
  XNOR U11988 ( .A(n12250), .B(n11149), .Z(n6363) );
  XOR U11989 ( .A(n10987), .B(n12251), .Z(n6362) );
  XOR U11990 ( .A(n4275), .B(n12252), .Z(n12243) );
  XNOR U11991 ( .A(n5835), .B(n2098), .Z(n12252) );
  XNOR U11992 ( .A(n12253), .B(n8496), .Z(n2098) );
  ANDN U11993 ( .B(n6375), .A(n6376), .Z(n12253) );
  XNOR U11994 ( .A(n12254), .B(n10048), .Z(n6376) );
  XOR U11995 ( .A(n11510), .B(n12255), .Z(n6375) );
  XOR U11996 ( .A(n12256), .B(n12257), .Z(n5835) );
  ANDN U11997 ( .B(n6379), .A(n6380), .Z(n12256) );
  XNOR U11998 ( .A(n10649), .B(n12258), .Z(n6380) );
  XOR U11999 ( .A(n12259), .B(n12260), .Z(n6379) );
  XNOR U12000 ( .A(n12261), .B(n8504), .Z(n4275) );
  AND U12001 ( .A(n6368), .B(n8505), .Z(n12261) );
  XNOR U12002 ( .A(n12262), .B(n10455), .Z(n8505) );
  XNOR U12003 ( .A(n12263), .B(n12264), .Z(n10455) );
  XNOR U12004 ( .A(n11309), .B(n12265), .Z(n6368) );
  XNOR U12005 ( .A(n12266), .B(n8487), .Z(n8431) );
  XNOR U12006 ( .A(n12267), .B(n11573), .Z(n8487) );
  ANDN U12007 ( .B(n12109), .A(n12110), .Z(n12266) );
  XNOR U12008 ( .A(n11386), .B(n12268), .Z(n12109) );
  XOR U12009 ( .A(n10850), .B(n2069), .Z(n5628) );
  XNOR U12010 ( .A(n7970), .B(n9122), .Z(n2069) );
  XNOR U12011 ( .A(n12269), .B(n12270), .Z(n9122) );
  XOR U12012 ( .A(n5432), .B(n3559), .Z(n12270) );
  XOR U12013 ( .A(n12271), .B(n12272), .Z(n3559) );
  NOR U12014 ( .A(n8120), .B(n8121), .Z(n12271) );
  XOR U12015 ( .A(n12273), .B(n10174), .Z(n8121) );
  XOR U12016 ( .A(n12274), .B(n10958), .Z(n5432) );
  ANDN U12017 ( .B(n8116), .A(n8117), .Z(n12274) );
  XNOR U12018 ( .A(n12275), .B(n10464), .Z(n8117) );
  XNOR U12019 ( .A(n12276), .B(n12277), .Z(n8116) );
  XOR U12020 ( .A(n6224), .B(n12278), .Z(n12269) );
  XOR U12021 ( .A(n2339), .B(n5366), .Z(n12278) );
  XNOR U12022 ( .A(n12279), .B(n10970), .Z(n5366) );
  AND U12023 ( .A(n9124), .B(n11082), .Z(n12279) );
  XOR U12024 ( .A(n10704), .B(n12280), .Z(n11082) );
  XNOR U12025 ( .A(n12281), .B(n12282), .Z(n9124) );
  XNOR U12026 ( .A(n12283), .B(n10961), .Z(n2339) );
  NOR U12027 ( .A(n8107), .B(n8106), .Z(n12283) );
  XNOR U12028 ( .A(n12284), .B(n11182), .Z(n8106) );
  XNOR U12029 ( .A(n12285), .B(n12286), .Z(n8107) );
  XNOR U12030 ( .A(n12287), .B(n10966), .Z(n6224) );
  AND U12031 ( .A(n8112), .B(n8110), .Z(n12287) );
  IV U12032 ( .A(n10967), .Z(n8110) );
  XOR U12033 ( .A(n10272), .B(n12288), .Z(n10967) );
  XOR U12034 ( .A(n12289), .B(n10938), .Z(n8112) );
  XOR U12035 ( .A(n12290), .B(n12291), .Z(n7970) );
  XOR U12036 ( .A(n3777), .B(n5102), .Z(n12291) );
  XOR U12037 ( .A(n12292), .B(n9033), .Z(n5102) );
  XOR U12038 ( .A(n11309), .B(n12293), .Z(n9033) );
  XOR U12039 ( .A(n12294), .B(n10160), .Z(n10857) );
  IV U12040 ( .A(n11182), .Z(n10160) );
  XOR U12041 ( .A(n11750), .B(n12295), .Z(n11182) );
  XOR U12042 ( .A(n12296), .B(n12297), .Z(n11750) );
  XOR U12043 ( .A(n12298), .B(n10472), .Z(n12297) );
  XOR U12044 ( .A(n12299), .B(n12300), .Z(n10472) );
  XOR U12045 ( .A(n11458), .B(n12303), .Z(n12296) );
  XOR U12046 ( .A(n12304), .B(n12305), .Z(n12303) );
  XOR U12047 ( .A(n12306), .B(n12307), .Z(n11458) );
  ANDN U12048 ( .B(n12308), .A(n12309), .Z(n12306) );
  XOR U12049 ( .A(n12310), .B(n9372), .Z(n10858) );
  XOR U12050 ( .A(n12311), .B(n8046), .Z(n3777) );
  IV U12051 ( .A(n10981), .Z(n8046) );
  XNOR U12052 ( .A(n12312), .B(n9697), .Z(n10981) );
  NOR U12053 ( .A(n10849), .B(n10848), .Z(n12311) );
  XNOR U12054 ( .A(n9552), .B(n12313), .Z(n10848) );
  IV U12055 ( .A(n9665), .Z(n9552) );
  IV U12056 ( .A(n12133), .Z(n10849) );
  XOR U12057 ( .A(n12314), .B(n9360), .Z(n12133) );
  XOR U12058 ( .A(n4263), .B(n12315), .Z(n12290) );
  XNOR U12059 ( .A(n1710), .B(n10953), .Z(n12315) );
  XNOR U12060 ( .A(n12316), .B(n8057), .Z(n10953) );
  XNOR U12061 ( .A(n12317), .B(n10296), .Z(n8057) );
  XNOR U12062 ( .A(n12318), .B(n12319), .Z(n10296) );
  AND U12063 ( .A(n10845), .B(n10844), .Z(n12316) );
  XNOR U12064 ( .A(n12320), .B(n10373), .Z(n10844) );
  XNOR U12065 ( .A(n12321), .B(n10277), .Z(n10845) );
  XNOR U12066 ( .A(n12322), .B(n8050), .Z(n1710) );
  XOR U12067 ( .A(n12323), .B(n10565), .Z(n8050) );
  AND U12068 ( .A(n10855), .B(n10853), .Z(n12322) );
  IV U12069 ( .A(n10974), .Z(n10853) );
  XNOR U12070 ( .A(n12324), .B(n9213), .Z(n10974) );
  XNOR U12071 ( .A(n12325), .B(n9483), .Z(n10855) );
  XNOR U12072 ( .A(n12326), .B(n12327), .Z(n9483) );
  XOR U12073 ( .A(n12328), .B(n8060), .Z(n4263) );
  IV U12074 ( .A(n10979), .Z(n8060) );
  XOR U12075 ( .A(n12329), .B(n11188), .Z(n10979) );
  XNOR U12076 ( .A(n12330), .B(n10978), .Z(n10850) );
  XNOR U12077 ( .A(n12331), .B(n10783), .Z(n10978) );
  AND U12078 ( .A(n12122), .B(n8059), .Z(n12330) );
  IV U12079 ( .A(n12123), .Z(n8059) );
  XNOR U12080 ( .A(n12332), .B(n11761), .Z(n12123) );
  XOR U12081 ( .A(n12333), .B(n11439), .Z(n12122) );
  IV U12082 ( .A(n11166), .Z(n11439) );
  XOR U12083 ( .A(n12334), .B(n6144), .Z(out[1006]) );
  XOR U12084 ( .A(n8737), .B(n2263), .Z(n6144) );
  XNOR U12085 ( .A(n6026), .B(n6103), .Z(n2263) );
  XNOR U12086 ( .A(n12335), .B(n12336), .Z(n6103) );
  XNOR U12087 ( .A(n2297), .B(n5420), .Z(n12336) );
  XNOR U12088 ( .A(n12337), .B(n7554), .Z(n5420) );
  XNOR U12089 ( .A(n12338), .B(n9820), .Z(n7554) );
  AND U12090 ( .A(n7555), .B(n8746), .Z(n12337) );
  XNOR U12091 ( .A(n9588), .B(n12339), .Z(n8746) );
  XNOR U12092 ( .A(n12340), .B(n10048), .Z(n7555) );
  XNOR U12093 ( .A(n12341), .B(n7559), .Z(n2297) );
  XNOR U12094 ( .A(n12342), .B(n9519), .Z(n7559) );
  AND U12095 ( .A(n7558), .B(n8742), .Z(n12341) );
  XOR U12096 ( .A(n12343), .B(n12344), .Z(n8742) );
  XOR U12097 ( .A(n12345), .B(n9704), .Z(n7558) );
  XOR U12098 ( .A(n3139), .B(n12346), .Z(n12335) );
  XOR U12099 ( .A(n6008), .B(n7548), .Z(n12346) );
  XNOR U12100 ( .A(n12347), .B(n7563), .Z(n7548) );
  XNOR U12101 ( .A(n12348), .B(n11464), .Z(n7563) );
  ANDN U12102 ( .B(n7564), .A(n8744), .Z(n12347) );
  XOR U12103 ( .A(n12349), .B(n10219), .Z(n8744) );
  XNOR U12104 ( .A(n12350), .B(n10251), .Z(n7564) );
  XNOR U12105 ( .A(n12351), .B(n7567), .Z(n6008) );
  XNOR U12106 ( .A(n12352), .B(n12069), .Z(n7567) );
  AND U12107 ( .A(n12218), .B(n12353), .Z(n12351) );
  XNOR U12108 ( .A(n12354), .B(n7571), .Z(n3139) );
  XNOR U12109 ( .A(n12355), .B(n10249), .Z(n7571) );
  AND U12110 ( .A(n7572), .B(n12198), .Z(n12354) );
  XOR U12111 ( .A(n12356), .B(n9692), .Z(n12198) );
  XNOR U12112 ( .A(n12357), .B(n12358), .Z(n7572) );
  XOR U12113 ( .A(n12359), .B(n12360), .Z(n6026) );
  XOR U12114 ( .A(n5232), .B(n1922), .Z(n12360) );
  XNOR U12115 ( .A(n12361), .B(n8802), .Z(n1922) );
  AND U12116 ( .A(n7646), .B(n8726), .Z(n12361) );
  IV U12117 ( .A(n8801), .Z(n8726) );
  XOR U12118 ( .A(n9537), .B(n12362), .Z(n8801) );
  XOR U12119 ( .A(n11060), .B(n12363), .Z(n7646) );
  XOR U12120 ( .A(n12364), .B(n8808), .Z(n5232) );
  ANDN U12121 ( .B(n7638), .A(n8724), .Z(n12364) );
  XNOR U12122 ( .A(n12365), .B(n12366), .Z(n8724) );
  XNOR U12123 ( .A(n12367), .B(n10256), .Z(n7638) );
  XNOR U12124 ( .A(n12368), .B(n12369), .Z(n10256) );
  XNOR U12125 ( .A(n3671), .B(n12370), .Z(n12359) );
  XOR U12126 ( .A(n8783), .B(n4151), .Z(n12370) );
  XOR U12127 ( .A(n12371), .B(n8810), .Z(n4151) );
  AND U12128 ( .A(n8733), .B(n8734), .Z(n12371) );
  XNOR U12129 ( .A(n12372), .B(n10226), .Z(n8734) );
  XOR U12130 ( .A(n11045), .B(n12373), .Z(n8733) );
  XNOR U12131 ( .A(n12374), .B(n8806), .Z(n8783) );
  NOR U12132 ( .A(n8729), .B(n7633), .Z(n12374) );
  XOR U12133 ( .A(n12375), .B(n12376), .Z(n7633) );
  XOR U12134 ( .A(n12298), .B(n10473), .Z(n8729) );
  XNOR U12135 ( .A(n12377), .B(n12378), .Z(n12298) );
  NOR U12136 ( .A(n12379), .B(n12380), .Z(n12377) );
  XNOR U12137 ( .A(n12381), .B(n12382), .Z(n3671) );
  AND U12138 ( .A(n7642), .B(n12383), .Z(n12381) );
  XNOR U12139 ( .A(n12384), .B(n12385), .Z(n7642) );
  XOR U12140 ( .A(n12386), .B(n12353), .Z(n8737) );
  IV U12141 ( .A(n7568), .Z(n12353) );
  XOR U12142 ( .A(n11686), .B(n12387), .Z(n7568) );
  XNOR U12143 ( .A(n12388), .B(n9119), .Z(n12218) );
  XOR U12144 ( .A(n11060), .B(n12389), .Z(n8697) );
  IV U12145 ( .A(n12164), .Z(n11060) );
  XOR U12146 ( .A(n10672), .B(n12390), .Z(n12164) );
  XOR U12147 ( .A(n12391), .B(n12392), .Z(n10672) );
  XOR U12148 ( .A(n12393), .B(n12394), .Z(n12392) );
  XOR U12149 ( .A(n11893), .B(n12395), .Z(n12391) );
  XOR U12150 ( .A(n12396), .B(n12397), .Z(n12395) );
  XNOR U12151 ( .A(n12398), .B(n12399), .Z(n11893) );
  NOR U12152 ( .A(n12400), .B(n12401), .Z(n12398) );
  ANDN U12153 ( .B(n5631), .A(n5632), .Z(n12334) );
  XOR U12154 ( .A(n10962), .B(n2072), .Z(n5632) );
  XNOR U12155 ( .A(n8041), .B(n9222), .Z(n2072) );
  XNOR U12156 ( .A(n12402), .B(n12403), .Z(n9222) );
  XOR U12157 ( .A(n5437), .B(n3564), .Z(n12403) );
  XOR U12158 ( .A(n12404), .B(n12405), .Z(n3564) );
  AND U12159 ( .A(n8147), .B(n8146), .Z(n12404) );
  XNOR U12160 ( .A(n10309), .B(n12406), .Z(n8147) );
  IV U12161 ( .A(n11712), .Z(n10309) );
  XNOR U12162 ( .A(n12407), .B(n11095), .Z(n5437) );
  AND U12163 ( .A(n8143), .B(n11096), .Z(n12407) );
  XOR U12164 ( .A(n12408), .B(n11315), .Z(n11096) );
  XNOR U12165 ( .A(n12393), .B(n11894), .Z(n8143) );
  XOR U12166 ( .A(n12409), .B(n12410), .Z(n12393) );
  NOR U12167 ( .A(n12411), .B(n12412), .Z(n12409) );
  XOR U12168 ( .A(n6229), .B(n12413), .Z(n12402) );
  XOR U12169 ( .A(n2346), .B(n5417), .Z(n12413) );
  XOR U12170 ( .A(n12414), .B(n12415), .Z(n5417) );
  AND U12171 ( .A(n9224), .B(n9226), .Z(n12414) );
  XNOR U12172 ( .A(n10692), .B(n12416), .Z(n9226) );
  XNOR U12173 ( .A(n12417), .B(n11194), .Z(n9224) );
  XNOR U12174 ( .A(n12418), .B(n12213), .Z(n11194) );
  XNOR U12175 ( .A(n12419), .B(n12420), .Z(n12213) );
  XOR U12176 ( .A(n11425), .B(n11237), .Z(n12420) );
  XOR U12177 ( .A(n12421), .B(n12422), .Z(n11237) );
  NOR U12178 ( .A(n12423), .B(n12424), .Z(n12421) );
  XNOR U12179 ( .A(n12425), .B(n12426), .Z(n11425) );
  AND U12180 ( .A(n12427), .B(n12428), .Z(n12425) );
  XOR U12181 ( .A(n12429), .B(n12430), .Z(n12419) );
  XOR U12182 ( .A(n11465), .B(n11799), .Z(n12430) );
  XOR U12183 ( .A(n12431), .B(n12432), .Z(n11799) );
  NOR U12184 ( .A(n12433), .B(n12434), .Z(n12431) );
  XNOR U12185 ( .A(n12435), .B(n12436), .Z(n11465) );
  ANDN U12186 ( .B(n12437), .A(n12438), .Z(n12435) );
  XOR U12187 ( .A(n12439), .B(n11099), .Z(n2346) );
  ANDN U12188 ( .B(n8132), .A(n8133), .Z(n12439) );
  XOR U12189 ( .A(n12440), .B(n9551), .Z(n8133) );
  XNOR U12190 ( .A(n12441), .B(n10803), .Z(n8132) );
  XNOR U12191 ( .A(n12442), .B(n11104), .Z(n6229) );
  ANDN U12192 ( .B(n8136), .A(n8137), .Z(n12442) );
  XOR U12193 ( .A(n12443), .B(n11037), .Z(n8137) );
  IV U12194 ( .A(n12444), .Z(n11037) );
  XNOR U12195 ( .A(n11121), .B(n12445), .Z(n8136) );
  XOR U12196 ( .A(n12446), .B(n12447), .Z(n8041) );
  XNOR U12197 ( .A(n3781), .B(n5104), .Z(n12447) );
  XOR U12198 ( .A(n12448), .B(n11083), .Z(n5104) );
  IV U12199 ( .A(n9126), .Z(n11083) );
  XOR U12200 ( .A(n9201), .B(n12449), .Z(n9126) );
  NOR U12201 ( .A(n10970), .B(n10969), .Z(n12448) );
  XNOR U12202 ( .A(n12450), .B(n10803), .Z(n10969) );
  XOR U12203 ( .A(n12451), .B(n9496), .Z(n10970) );
  XOR U12204 ( .A(n12452), .B(n8108), .Z(n3781) );
  IV U12205 ( .A(n11088), .Z(n8108) );
  XNOR U12206 ( .A(n12453), .B(n9803), .Z(n11088) );
  ANDN U12207 ( .B(n10961), .A(n10960), .Z(n12452) );
  XNOR U12208 ( .A(n12454), .B(n9663), .Z(n10960) );
  IV U12209 ( .A(n9773), .Z(n9663) );
  XOR U12210 ( .A(n12455), .B(n12456), .Z(n10961) );
  XOR U12211 ( .A(n4291), .B(n12457), .Z(n12446) );
  XOR U12212 ( .A(n1719), .B(n11076), .Z(n12457) );
  XOR U12213 ( .A(n12458), .B(n8118), .Z(n11076) );
  IV U12214 ( .A(n11090), .Z(n8118) );
  XOR U12215 ( .A(n10695), .B(n12459), .Z(n11090) );
  AND U12216 ( .A(n10957), .B(n10958), .Z(n12458) );
  XOR U12217 ( .A(n12460), .B(n12461), .Z(n10958) );
  XOR U12218 ( .A(n12462), .B(n10553), .Z(n10957) );
  XOR U12219 ( .A(n12463), .B(n8111), .Z(n1719) );
  IV U12220 ( .A(n11080), .Z(n8111) );
  XOR U12221 ( .A(n11396), .B(n12464), .Z(n11080) );
  IV U12222 ( .A(n11069), .Z(n11396) );
  ANDN U12223 ( .B(n10965), .A(n10966), .Z(n12463) );
  XNOR U12224 ( .A(n9665), .B(n12465), .Z(n10966) );
  XOR U12225 ( .A(n12466), .B(n12467), .Z(n9665) );
  XOR U12226 ( .A(n12468), .B(n9119), .Z(n10965) );
  XNOR U12227 ( .A(n12469), .B(n8122), .Z(n4291) );
  XNOR U12228 ( .A(n12470), .B(n11315), .Z(n8122) );
  XNOR U12229 ( .A(n12471), .B(n11086), .Z(n10962) );
  XOR U12230 ( .A(n12472), .B(n9360), .Z(n11086) );
  IV U12231 ( .A(n12473), .Z(n9360) );
  AND U12232 ( .A(n8120), .B(n12272), .Z(n12471) );
  XOR U12233 ( .A(n12474), .B(n11293), .Z(n12272) );
  IV U12234 ( .A(n11573), .Z(n11293) );
  XOR U12235 ( .A(n11257), .B(n12475), .Z(n8120) );
  XOR U12236 ( .A(n1756), .B(n8500), .Z(n5631) );
  XNOR U12237 ( .A(n12476), .B(n8603), .Z(n8500) );
  NOR U12238 ( .A(n12246), .B(n6371), .Z(n12476) );
  XNOR U12239 ( .A(n10838), .B(n12477), .Z(n6371) );
  IV U12240 ( .A(n3824), .Z(n1756) );
  XOR U12241 ( .A(n9854), .B(n6267), .Z(n3824) );
  XOR U12242 ( .A(n12478), .B(n12479), .Z(n6267) );
  XNOR U12243 ( .A(n5845), .B(n2104), .Z(n12479) );
  XOR U12244 ( .A(n12480), .B(n8610), .Z(n2104) );
  XOR U12245 ( .A(n12481), .B(n10149), .Z(n6402) );
  XOR U12246 ( .A(n11753), .B(n11326), .Z(n9187) );
  XOR U12247 ( .A(n12483), .B(n12484), .Z(n11326) );
  XNOR U12248 ( .A(n12417), .B(n11429), .Z(n12484) );
  XOR U12249 ( .A(n12485), .B(n12486), .Z(n11429) );
  ANDN U12250 ( .B(n12487), .A(n12488), .Z(n12485) );
  XNOR U12251 ( .A(n12489), .B(n12490), .Z(n12417) );
  AND U12252 ( .A(n12491), .B(n12492), .Z(n12489) );
  XNOR U12253 ( .A(n11193), .B(n12493), .Z(n12483) );
  XNOR U12254 ( .A(n9389), .B(n11662), .Z(n12493) );
  XNOR U12255 ( .A(n12494), .B(n12495), .Z(n11662) );
  NOR U12256 ( .A(n12496), .B(n12497), .Z(n12494) );
  XNOR U12257 ( .A(n12498), .B(n12499), .Z(n9389) );
  AND U12258 ( .A(n12500), .B(n12501), .Z(n12498) );
  XNOR U12259 ( .A(n12502), .B(n12503), .Z(n11193) );
  AND U12260 ( .A(n12504), .B(n12505), .Z(n12502) );
  XOR U12261 ( .A(n12506), .B(n12507), .Z(n11753) );
  XNOR U12262 ( .A(n12508), .B(n12509), .Z(n12507) );
  XNOR U12263 ( .A(n12510), .B(n12511), .Z(n12506) );
  XOR U12264 ( .A(n12259), .B(n9106), .Z(n12511) );
  XNOR U12265 ( .A(n12512), .B(n12513), .Z(n9106) );
  ANDN U12266 ( .B(n12514), .A(n12515), .Z(n12512) );
  XOR U12267 ( .A(n12516), .B(n12517), .Z(n12259) );
  ANDN U12268 ( .B(n12518), .A(n12519), .Z(n12516) );
  XOR U12269 ( .A(n12520), .B(n8621), .Z(n5845) );
  ANDN U12270 ( .B(n6405), .A(n6407), .Z(n12520) );
  XNOR U12271 ( .A(n9684), .B(n12521), .Z(n6407) );
  XNOR U12272 ( .A(n12522), .B(n12523), .Z(n6405) );
  XOR U12273 ( .A(n3652), .B(n12524), .Z(n12478) );
  XOR U12274 ( .A(n4278), .B(n5406), .Z(n12524) );
  XNOR U12275 ( .A(n12525), .B(n12526), .Z(n5406) );
  NOR U12276 ( .A(n6388), .B(n6389), .Z(n12525) );
  XNOR U12277 ( .A(n12527), .B(n12058), .Z(n6389) );
  XOR U12278 ( .A(n12528), .B(n11121), .Z(n6388) );
  XNOR U12279 ( .A(n12529), .B(n8618), .Z(n4278) );
  ANDN U12280 ( .B(n6392), .A(n6393), .Z(n12529) );
  XNOR U12281 ( .A(n9201), .B(n12530), .Z(n6393) );
  XOR U12282 ( .A(n12531), .B(n12532), .Z(n6392) );
  XOR U12283 ( .A(n12533), .B(n12534), .Z(n3652) );
  ANDN U12284 ( .B(n6397), .A(n6398), .Z(n12533) );
  XNOR U12285 ( .A(n10557), .B(n12535), .Z(n6398) );
  XOR U12286 ( .A(n12536), .B(n12537), .Z(n9854) );
  XNOR U12287 ( .A(n4838), .B(n8596), .Z(n12537) );
  XNOR U12288 ( .A(n12538), .B(n6364), .Z(n8596) );
  XNOR U12289 ( .A(n9511), .B(n12539), .Z(n6364) );
  IV U12290 ( .A(n10262), .Z(n9511) );
  XOR U12291 ( .A(n12540), .B(n12541), .Z(n10262) );
  AND U12292 ( .A(n8498), .B(n12249), .Z(n12538) );
  IV U12293 ( .A(n8499), .Z(n12249) );
  XOR U12294 ( .A(n12531), .B(n12542), .Z(n8499) );
  IV U12295 ( .A(n10704), .Z(n12531) );
  XNOR U12296 ( .A(n12543), .B(n10227), .Z(n8498) );
  XNOR U12297 ( .A(n12544), .B(n6367), .Z(n4838) );
  XNOR U12298 ( .A(n12545), .B(n12205), .Z(n6367) );
  NOR U12299 ( .A(n8503), .B(n8504), .Z(n12544) );
  XNOR U12300 ( .A(n9894), .B(n12546), .Z(n8504) );
  XOR U12301 ( .A(n12549), .B(n11686), .Z(n8503) );
  XNOR U12302 ( .A(n2491), .B(n12550), .Z(n12536) );
  XOR U12303 ( .A(n3457), .B(n4317), .Z(n12550) );
  XNOR U12304 ( .A(n12551), .B(n6373), .Z(n4317) );
  XNOR U12305 ( .A(n10922), .B(n12552), .Z(n6373) );
  IV U12306 ( .A(n12553), .Z(n10922) );
  ANDN U12307 ( .B(n12246), .A(n8603), .Z(n12551) );
  XNOR U12308 ( .A(n12554), .B(n11890), .Z(n8603) );
  XNOR U12309 ( .A(n12555), .B(n11522), .Z(n12246) );
  XNOR U12310 ( .A(n12556), .B(n6377), .Z(n3457) );
  XNOR U12311 ( .A(n9208), .B(n12557), .Z(n6377) );
  IV U12312 ( .A(n11877), .Z(n9208) );
  XOR U12313 ( .A(n12558), .B(n12559), .Z(n11877) );
  NOR U12314 ( .A(n8496), .B(n8495), .Z(n12556) );
  XNOR U12315 ( .A(n12560), .B(n9278), .Z(n8495) );
  XNOR U12316 ( .A(n12561), .B(n12058), .Z(n8496) );
  IV U12317 ( .A(n11280), .Z(n12058) );
  XNOR U12318 ( .A(n12562), .B(n6381), .Z(n2491) );
  XNOR U12319 ( .A(n12563), .B(n11198), .Z(n6381) );
  AND U12320 ( .A(n8507), .B(n12257), .Z(n12562) );
  IV U12321 ( .A(n8508), .Z(n12257) );
  XOR U12322 ( .A(n10127), .B(n12564), .Z(n8508) );
  IV U12323 ( .A(n10909), .Z(n10127) );
  XNOR U12324 ( .A(n10557), .B(n12565), .Z(n8507) );
  XOR U12325 ( .A(n12566), .B(n6149), .Z(out[1005]) );
  XOR U12326 ( .A(n8799), .B(n2270), .Z(n6149) );
  XNOR U12327 ( .A(n6031), .B(n6108), .Z(n2270) );
  XNOR U12328 ( .A(n12567), .B(n12568), .Z(n6108) );
  XNOR U12329 ( .A(n2308), .B(n5424), .Z(n12568) );
  XOR U12330 ( .A(n12569), .B(n7630), .Z(n5424) );
  XNOR U12331 ( .A(n10898), .B(n12570), .Z(n7630) );
  ANDN U12332 ( .B(n7631), .A(n8810), .Z(n12569) );
  XNOR U12333 ( .A(n12571), .B(n9720), .Z(n8810) );
  XOR U12334 ( .A(n10149), .B(n12572), .Z(n7631) );
  XNOR U12335 ( .A(n12573), .B(n7634), .Z(n2308) );
  XOR U12336 ( .A(n9588), .B(n12574), .Z(n7634) );
  AND U12337 ( .A(n8806), .B(n8805), .Z(n12573) );
  XOR U12338 ( .A(n12575), .B(n9810), .Z(n8805) );
  XNOR U12339 ( .A(n12576), .B(n11896), .Z(n8806) );
  IV U12340 ( .A(n11149), .Z(n11896) );
  XOR U12341 ( .A(n3143), .B(n12579), .Z(n12567) );
  XNOR U12342 ( .A(n6059), .B(n7624), .Z(n12579) );
  XNOR U12343 ( .A(n12580), .B(n7640), .Z(n7624) );
  XOR U12344 ( .A(n12581), .B(n11602), .Z(n7640) );
  NOR U12345 ( .A(n8808), .B(n7639), .Z(n12580) );
  XNOR U12346 ( .A(n12582), .B(n10382), .Z(n7639) );
  XOR U12347 ( .A(n12585), .B(n10431), .Z(n8808) );
  XNOR U12348 ( .A(n12586), .B(n7644), .Z(n6059) );
  XNOR U12349 ( .A(n12205), .B(n12587), .Z(n7644) );
  ANDN U12350 ( .B(n12382), .A(n7643), .Z(n12586) );
  XNOR U12351 ( .A(n12588), .B(n7647), .Z(n3143) );
  XNOR U12352 ( .A(n10379), .B(n12589), .Z(n7647) );
  AND U12353 ( .A(n8802), .B(n7648), .Z(n12588) );
  XOR U12354 ( .A(n12590), .B(n11916), .Z(n7648) );
  XNOR U12355 ( .A(n12591), .B(n9800), .Z(n8802) );
  XOR U12356 ( .A(n12592), .B(n12593), .Z(n6031) );
  XNOR U12357 ( .A(n5234), .B(n1927), .Z(n12593) );
  ANDN U12358 ( .B(n8789), .A(n7723), .Z(n12594) );
  XNOR U12359 ( .A(n12595), .B(n12277), .Z(n7723) );
  XOR U12360 ( .A(n11993), .B(n12596), .Z(n8789) );
  XOR U12361 ( .A(n12597), .B(n12598), .Z(n11993) );
  XNOR U12362 ( .A(n12599), .B(n8871), .Z(n5234) );
  ANDN U12363 ( .B(n8787), .A(n7715), .Z(n12599) );
  XOR U12364 ( .A(n12600), .B(n10386), .Z(n7715) );
  XNOR U12365 ( .A(n12601), .B(n12602), .Z(n10386) );
  XNOR U12366 ( .A(n12603), .B(n12604), .Z(n8787) );
  XNOR U12367 ( .A(n3678), .B(n12605), .Z(n12592) );
  XNOR U12368 ( .A(n8847), .B(n4155), .Z(n12605) );
  XOR U12369 ( .A(n12606), .B(n8873), .Z(n4155) );
  NOR U12370 ( .A(n7706), .B(n8796), .Z(n12606) );
  XOR U12371 ( .A(n12607), .B(n12385), .Z(n8796) );
  XNOR U12372 ( .A(n12608), .B(n9163), .Z(n7706) );
  XNOR U12373 ( .A(n12609), .B(n8869), .Z(n8847) );
  ANDN U12374 ( .B(n7710), .A(n8792), .Z(n12609) );
  XOR U12375 ( .A(n12610), .B(n10233), .Z(n8792) );
  IV U12376 ( .A(n9403), .Z(n10233) );
  XNOR U12377 ( .A(n12611), .B(n12612), .Z(n9403) );
  XNOR U12378 ( .A(n12613), .B(n12176), .Z(n7710) );
  XNOR U12379 ( .A(n12614), .B(n12615), .Z(n3678) );
  NOR U12380 ( .A(n8794), .B(n7719), .Z(n12614) );
  XOR U12381 ( .A(n12616), .B(n10136), .Z(n7719) );
  XOR U12382 ( .A(n12617), .B(n7643), .Z(n8799) );
  XNOR U12383 ( .A(n12005), .B(n12618), .Z(n7643) );
  ANDN U12384 ( .B(n8731), .A(n12382), .Z(n12617) );
  XOR U12385 ( .A(n9191), .B(n12619), .Z(n12382) );
  IV U12386 ( .A(n12383), .Z(n8731) );
  XOR U12387 ( .A(n12620), .B(n11188), .Z(n12383) );
  IV U12388 ( .A(n12277), .Z(n11188) );
  XOR U12389 ( .A(n12621), .B(n12622), .Z(n12277) );
  ANDN U12390 ( .B(n5637), .A(n5635), .Z(n12566) );
  XNOR U12391 ( .A(n8615), .B(n5128), .Z(n5635) );
  XNOR U12392 ( .A(n12623), .B(n12624), .Z(n6358) );
  XNOR U12393 ( .A(n4353), .B(n2497), .Z(n12624) );
  XNOR U12394 ( .A(n12625), .B(n6406), .Z(n2497) );
  XOR U12395 ( .A(n12626), .B(n11324), .Z(n6406) );
  IV U12396 ( .A(n11404), .Z(n11324) );
  ANDN U12397 ( .B(n8666), .A(n8621), .Z(n12625) );
  XOR U12398 ( .A(n12627), .B(n10987), .Z(n8621) );
  IV U12399 ( .A(n10272), .Z(n10987) );
  XOR U12400 ( .A(n12628), .B(n12629), .Z(n10272) );
  XOR U12401 ( .A(n12630), .B(n10681), .Z(n8666) );
  XNOR U12402 ( .A(n12631), .B(n6399), .Z(n4353) );
  XNOR U12403 ( .A(n10917), .B(n12632), .Z(n6399) );
  AND U12404 ( .A(n12534), .B(n12633), .Z(n12631) );
  XOR U12405 ( .A(n3460), .B(n12634), .Z(n12623) );
  XOR U12406 ( .A(n8655), .B(n4842), .Z(n12634) );
  XOR U12407 ( .A(n12635), .B(n6394), .Z(n4842) );
  XOR U12408 ( .A(n12636), .B(n12366), .Z(n6394) );
  AND U12409 ( .A(n8617), .B(n8618), .Z(n12635) );
  XOR U12410 ( .A(n10377), .B(n12637), .Z(n8618) );
  XOR U12411 ( .A(n12005), .B(n12638), .Z(n8617) );
  XOR U12412 ( .A(n12639), .B(n6390), .Z(n8655) );
  XNOR U12413 ( .A(n12640), .B(n9582), .Z(n6390) );
  AND U12414 ( .A(n8612), .B(n12526), .Z(n12639) );
  IV U12415 ( .A(n8613), .Z(n12526) );
  XNOR U12416 ( .A(n12641), .B(n10692), .Z(n8613) );
  XOR U12417 ( .A(n10359), .B(n12642), .Z(n8612) );
  XNOR U12418 ( .A(n12643), .B(n6403), .Z(n3460) );
  XNOR U12419 ( .A(n12644), .B(n12645), .Z(n6403) );
  ANDN U12420 ( .B(n8664), .A(n8610), .Z(n12643) );
  XOR U12421 ( .A(n12646), .B(n12193), .Z(n8610) );
  IV U12422 ( .A(n11418), .Z(n12193) );
  XOR U12423 ( .A(n12647), .B(n10055), .Z(n8664) );
  XNOR U12424 ( .A(n12648), .B(n12649), .Z(n6273) );
  XOR U12425 ( .A(n5410), .B(n3659), .Z(n12649) );
  XNOR U12426 ( .A(n12650), .B(n12651), .Z(n3659) );
  AND U12427 ( .A(n6424), .B(n8752), .Z(n12650) );
  XNOR U12428 ( .A(n12652), .B(n10681), .Z(n8752) );
  XNOR U12429 ( .A(n12653), .B(n8675), .Z(n5410) );
  AND U12430 ( .A(n6416), .B(n8676), .Z(n12653) );
  XNOR U12431 ( .A(n12654), .B(n11782), .Z(n8676) );
  XOR U12432 ( .A(n11418), .B(n12655), .Z(n6416) );
  XNOR U12433 ( .A(n4280), .B(n12656), .Z(n12648) );
  XOR U12434 ( .A(n5850), .B(n2108), .Z(n12656) );
  XNOR U12435 ( .A(n12657), .B(n8671), .Z(n2108) );
  AND U12436 ( .A(n6429), .B(n8672), .Z(n12657) );
  XNOR U12437 ( .A(n12658), .B(n9261), .Z(n8672) );
  XOR U12438 ( .A(n12659), .B(n10293), .Z(n6429) );
  XOR U12439 ( .A(n12660), .B(n8684), .Z(n5850) );
  AND U12440 ( .A(n6434), .B(n8685), .Z(n12660) );
  XOR U12441 ( .A(n12661), .B(n12662), .Z(n8685) );
  XNOR U12442 ( .A(n12663), .B(n9077), .Z(n6434) );
  XOR U12443 ( .A(n12664), .B(n8681), .Z(n4280) );
  NOR U12444 ( .A(n6420), .B(n6419), .Z(n12664) );
  XNOR U12445 ( .A(n10692), .B(n12665), .Z(n6419) );
  XOR U12446 ( .A(n9399), .B(n12668), .Z(n6420) );
  XOR U12447 ( .A(n12669), .B(n8662), .Z(n8615) );
  IV U12448 ( .A(n12633), .Z(n8662) );
  XOR U12449 ( .A(n12670), .B(n11586), .Z(n12633) );
  IV U12450 ( .A(n12671), .Z(n11586) );
  NOR U12451 ( .A(n6397), .B(n12534), .Z(n12669) );
  XNOR U12452 ( .A(n12672), .B(n10003), .Z(n12534) );
  XOR U12453 ( .A(n12673), .B(n11007), .Z(n6397) );
  XNOR U12454 ( .A(n11100), .B(n2076), .Z(n5637) );
  XNOR U12455 ( .A(n8102), .B(n9344), .Z(n2076) );
  XNOR U12456 ( .A(n12674), .B(n12675), .Z(n9344) );
  XOR U12457 ( .A(n5441), .B(n3569), .Z(n12675) );
  XOR U12458 ( .A(n12676), .B(n12677), .Z(n3569) );
  AND U12459 ( .A(n8201), .B(n12678), .Z(n12676) );
  XNOR U12460 ( .A(n10544), .B(n12679), .Z(n8201) );
  XNOR U12461 ( .A(n12680), .B(n11217), .Z(n5441) );
  ANDN U12462 ( .B(n8196), .A(n8197), .Z(n12680) );
  XOR U12463 ( .A(n12681), .B(n12056), .Z(n8197) );
  IV U12464 ( .A(n10714), .Z(n12056) );
  IV U12465 ( .A(n11218), .Z(n8196) );
  XOR U12466 ( .A(n6233), .B(n12683), .Z(n12674) );
  XNOR U12467 ( .A(n2353), .B(n5469), .Z(n12683) );
  XNOR U12468 ( .A(n12684), .B(n11229), .Z(n5469) );
  AND U12469 ( .A(n9348), .B(n9346), .Z(n12684) );
  IV U12470 ( .A(n11230), .Z(n9346) );
  XOR U12471 ( .A(n9516), .B(n12685), .Z(n11230) );
  XOR U12472 ( .A(n12686), .B(n12687), .Z(n9516) );
  XNOR U12473 ( .A(n12688), .B(n10794), .Z(n9348) );
  XNOR U12474 ( .A(n12689), .B(n11221), .Z(n2353) );
  ANDN U12475 ( .B(n8188), .A(n8186), .Z(n12689) );
  XOR U12476 ( .A(n12690), .B(n10478), .Z(n8186) );
  XNOR U12477 ( .A(n12691), .B(n10165), .Z(n8188) );
  IV U12478 ( .A(n9659), .Z(n10165) );
  XNOR U12479 ( .A(n12692), .B(n11226), .Z(n6233) );
  ANDN U12480 ( .B(n8190), .A(n8191), .Z(n12692) );
  XNOR U12481 ( .A(n12693), .B(n11166), .Z(n8191) );
  XNOR U12482 ( .A(n12694), .B(n11782), .Z(n8190) );
  XOR U12483 ( .A(n12695), .B(n12696), .Z(n8102) );
  XOR U12484 ( .A(n3786), .B(n5107), .Z(n12696) );
  XOR U12485 ( .A(n12697), .B(n9225), .Z(n5107) );
  XNOR U12486 ( .A(n9399), .B(n12698), .Z(n9225) );
  AND U12487 ( .A(n11106), .B(n12415), .Z(n12697) );
  IV U12488 ( .A(n11107), .Z(n12415) );
  XOR U12489 ( .A(n9574), .B(n12699), .Z(n11107) );
  XNOR U12490 ( .A(n12700), .B(n10478), .Z(n11106) );
  XNOR U12491 ( .A(n12701), .B(n12702), .Z(n10478) );
  XNOR U12492 ( .A(n12703), .B(n8134), .Z(n3786) );
  XOR U12493 ( .A(n12704), .B(n12376), .Z(n8134) );
  IV U12494 ( .A(n9927), .Z(n12376) );
  ANDN U12495 ( .B(n11099), .A(n11098), .Z(n12703) );
  XNOR U12496 ( .A(n9769), .B(n12705), .Z(n11098) );
  XNOR U12497 ( .A(n9558), .B(n12706), .Z(n11099) );
  XNOR U12498 ( .A(n4316), .B(n12707), .Z(n12695) );
  XNOR U12499 ( .A(n1724), .B(n11201), .Z(n12707) );
  XNOR U12500 ( .A(n12708), .B(n8144), .Z(n11201) );
  XOR U12501 ( .A(n12709), .B(n10594), .Z(n8144) );
  XNOR U12502 ( .A(n12710), .B(n12711), .Z(n10594) );
  XOR U12503 ( .A(n12712), .B(n10584), .Z(n11095) );
  IV U12504 ( .A(n11212), .Z(n11094) );
  XNOR U12505 ( .A(n12713), .B(n10675), .Z(n11212) );
  XOR U12506 ( .A(n12714), .B(n12715), .Z(n10675) );
  XOR U12507 ( .A(n12716), .B(n11205), .Z(n1724) );
  IV U12508 ( .A(n8138), .Z(n11205) );
  XOR U12509 ( .A(n12717), .B(n11197), .Z(n8138) );
  ANDN U12510 ( .B(n11103), .A(n11104), .Z(n12716) );
  XNOR U12511 ( .A(n12718), .B(n9773), .Z(n11104) );
  XNOR U12512 ( .A(n12719), .B(n12720), .Z(n9773) );
  XNOR U12513 ( .A(n9191), .B(n12721), .Z(n11103) );
  XNOR U12514 ( .A(n12722), .B(n8148), .Z(n4316) );
  XNOR U12515 ( .A(n12723), .B(n11456), .Z(n8148) );
  AND U12516 ( .A(n12724), .B(n12405), .Z(n12722) );
  IV U12517 ( .A(n12725), .Z(n12405) );
  XOR U12518 ( .A(n12726), .B(n12724), .Z(n11100) );
  IV U12519 ( .A(n11209), .Z(n12724) );
  XOR U12520 ( .A(n9488), .B(n12727), .Z(n11209) );
  IV U12521 ( .A(n12455), .Z(n9488) );
  ANDN U12522 ( .B(n12725), .A(n8146), .Z(n12726) );
  XOR U12523 ( .A(n12728), .B(n12729), .Z(n8146) );
  XOR U12524 ( .A(n11890), .B(n12730), .Z(n12725) );
  XOR U12525 ( .A(n12731), .B(n6154), .Z(out[1004]) );
  IV U12526 ( .A(n6907), .Z(n6154) );
  XNOR U12527 ( .A(n8863), .B(n2275), .Z(n6907) );
  XNOR U12528 ( .A(n6037), .B(n6118), .Z(n2275) );
  XNOR U12529 ( .A(n12732), .B(n12733), .Z(n6118) );
  XOR U12530 ( .A(n2315), .B(n5428), .Z(n12733) );
  XNOR U12531 ( .A(n12734), .B(n7707), .Z(n5428) );
  XOR U12532 ( .A(n10229), .B(n12735), .Z(n7707) );
  ANDN U12533 ( .B(n7708), .A(n8873), .Z(n12734) );
  XNOR U12534 ( .A(n12736), .B(n9822), .Z(n8873) );
  XOR U12535 ( .A(n12737), .B(n10293), .Z(n7708) );
  XNOR U12536 ( .A(n12738), .B(n7712), .Z(n2315) );
  XOR U12537 ( .A(n12739), .B(n9699), .Z(n7712) );
  AND U12538 ( .A(n8869), .B(n8868), .Z(n12738) );
  XOR U12539 ( .A(n12234), .B(n12740), .Z(n8868) );
  XNOR U12540 ( .A(n12741), .B(n11280), .Z(n8869) );
  XNOR U12541 ( .A(n12743), .B(n12744), .Z(n12162) );
  XNOR U12542 ( .A(n9667), .B(n12745), .Z(n12744) );
  XNOR U12543 ( .A(n12746), .B(n12747), .Z(n9667) );
  XNOR U12544 ( .A(n11251), .B(n12750), .Z(n12743) );
  XNOR U12545 ( .A(n10241), .B(n12751), .Z(n12750) );
  XOR U12546 ( .A(n12752), .B(n12753), .Z(n10241) );
  AND U12547 ( .A(n12754), .B(n12755), .Z(n12752) );
  XNOR U12548 ( .A(n12756), .B(n12757), .Z(n11251) );
  NOR U12549 ( .A(n12758), .B(n12759), .Z(n12756) );
  XNOR U12550 ( .A(n3148), .B(n12760), .Z(n12732) );
  XOR U12551 ( .A(n6113), .B(n7701), .Z(n12760) );
  XOR U12552 ( .A(n12761), .B(n7717), .Z(n7701) );
  XOR U12553 ( .A(n12762), .B(n12763), .Z(n7717) );
  ANDN U12554 ( .B(n8871), .A(n7716), .Z(n12761) );
  XOR U12555 ( .A(n10557), .B(n12764), .Z(n7716) );
  XOR U12556 ( .A(n9108), .B(n12767), .Z(n8871) );
  IV U12557 ( .A(n11663), .Z(n9108) );
  XOR U12558 ( .A(n12768), .B(n12769), .Z(n11902) );
  XOR U12559 ( .A(n9999), .B(n11125), .Z(n12769) );
  XNOR U12560 ( .A(n12770), .B(n12771), .Z(n11125) );
  XNOR U12561 ( .A(n12774), .B(n12775), .Z(n9999) );
  ANDN U12562 ( .B(n12776), .A(n12777), .Z(n12774) );
  XOR U12563 ( .A(n11265), .B(n12778), .Z(n12768) );
  XNOR U12564 ( .A(n12779), .B(n12780), .Z(n12778) );
  XOR U12565 ( .A(n12781), .B(n12782), .Z(n11265) );
  ANDN U12566 ( .B(n12783), .A(n12784), .Z(n12781) );
  XOR U12567 ( .A(n12786), .B(n7721), .Z(n6113) );
  XOR U12568 ( .A(n12787), .B(n12366), .Z(n7721) );
  AND U12569 ( .A(n7720), .B(n12615), .Z(n12786) );
  XNOR U12570 ( .A(n12788), .B(n7724), .Z(n3148) );
  XOR U12571 ( .A(n10559), .B(n12789), .Z(n7724) );
  AND U12572 ( .A(n7725), .B(n8865), .Z(n12788) );
  XOR U12573 ( .A(n12790), .B(n9922), .Z(n8865) );
  XNOR U12574 ( .A(n12791), .B(n12074), .Z(n7725) );
  XOR U12575 ( .A(n12792), .B(n12793), .Z(n6037) );
  XNOR U12576 ( .A(n5237), .B(n1931), .Z(n12793) );
  XNOR U12577 ( .A(n12794), .B(n8929), .Z(n1931) );
  ANDN U12578 ( .B(n7790), .A(n8853), .Z(n12794) );
  XOR U12579 ( .A(n12795), .B(n9718), .Z(n8853) );
  XNOR U12580 ( .A(n12796), .B(n12797), .Z(n9718) );
  XOR U12581 ( .A(n12798), .B(n11315), .Z(n7790) );
  XNOR U12582 ( .A(n12799), .B(n8934), .Z(n5237) );
  ANDN U12583 ( .B(n7782), .A(n8851), .Z(n12799) );
  XOR U12584 ( .A(n12509), .B(n9107), .Z(n8851) );
  IV U12585 ( .A(n12260), .Z(n9107) );
  XNOR U12586 ( .A(n12800), .B(n12801), .Z(n12509) );
  ANDN U12587 ( .B(n12802), .A(n12803), .Z(n12800) );
  XNOR U12588 ( .A(n12804), .B(n10565), .Z(n7782) );
  XNOR U12589 ( .A(n12629), .B(n12805), .Z(n10565) );
  XOR U12590 ( .A(n12806), .B(n12807), .Z(n12629) );
  XNOR U12591 ( .A(n12808), .B(n10358), .Z(n12807) );
  NOR U12592 ( .A(n12811), .B(n12812), .Z(n12809) );
  XOR U12593 ( .A(n9162), .B(n12813), .Z(n12806) );
  XNOR U12594 ( .A(n12814), .B(n12608), .Z(n12813) );
  XNOR U12595 ( .A(n12815), .B(n12816), .Z(n12608) );
  ANDN U12596 ( .B(n12817), .A(n12818), .Z(n12815) );
  XNOR U12597 ( .A(n12819), .B(n12820), .Z(n9162) );
  NOR U12598 ( .A(n12821), .B(n12822), .Z(n12819) );
  XOR U12599 ( .A(n3684), .B(n12823), .Z(n12792) );
  XNOR U12600 ( .A(n8911), .B(n4161), .Z(n12823) );
  XOR U12601 ( .A(n12824), .B(n8936), .Z(n4161) );
  IV U12602 ( .A(n12825), .Z(n8936) );
  ANDN U12603 ( .B(n8860), .A(n7773), .Z(n12824) );
  XOR U12604 ( .A(n12826), .B(n9067), .Z(n7773) );
  XNOR U12605 ( .A(n12827), .B(n10136), .Z(n8860) );
  XNOR U12606 ( .A(n12828), .B(n12829), .Z(n10136) );
  XNOR U12607 ( .A(n12830), .B(n8932), .Z(n8911) );
  AND U12608 ( .A(n8856), .B(n7777), .Z(n12830) );
  XNOR U12609 ( .A(n12831), .B(n12832), .Z(n7777) );
  XNOR U12610 ( .A(n11872), .B(n12833), .Z(n8856) );
  XOR U12611 ( .A(n12834), .B(n12835), .Z(n11872) );
  XNOR U12612 ( .A(n12836), .B(n12837), .Z(n3684) );
  ANDN U12613 ( .B(n8858), .A(n7786), .Z(n12836) );
  XNOR U12614 ( .A(n12838), .B(n11442), .Z(n7786) );
  IV U12615 ( .A(n10281), .Z(n11442) );
  XNOR U12616 ( .A(n12839), .B(n7720), .Z(n8863) );
  XOR U12617 ( .A(n12840), .B(n10991), .Z(n7720) );
  XOR U12618 ( .A(n12841), .B(n9529), .Z(n12615) );
  XOR U12619 ( .A(n12842), .B(n11315), .Z(n8794) );
  XNOR U12620 ( .A(n12843), .B(n12844), .Z(n11315) );
  ANDN U12621 ( .B(n5641), .A(n5639), .Z(n12731) );
  XNOR U12622 ( .A(n8678), .B(n5131), .Z(n5639) );
  XNOR U12623 ( .A(n6278), .B(n6384), .Z(n5131) );
  XNOR U12624 ( .A(n12845), .B(n12846), .Z(n6384) );
  XNOR U12625 ( .A(n4752), .B(n2504), .Z(n12846) );
  XOR U12626 ( .A(n12847), .B(n6433), .Z(n2504) );
  XNOR U12627 ( .A(n12848), .B(n11464), .Z(n6433) );
  ANDN U12628 ( .B(n8683), .A(n8684), .Z(n12847) );
  XNOR U12629 ( .A(n11121), .B(n12849), .Z(n8684) );
  XNOR U12630 ( .A(n12850), .B(n10903), .Z(n8683) );
  XNOR U12631 ( .A(n12851), .B(n6426), .Z(n4752) );
  XNOR U12632 ( .A(n12852), .B(n10995), .Z(n6426) );
  AND U12633 ( .A(n12651), .B(n12853), .Z(n12851) );
  XOR U12634 ( .A(n3463), .B(n12854), .Z(n12845) );
  XOR U12635 ( .A(n8747), .B(n4845), .Z(n12854) );
  XOR U12636 ( .A(n12855), .B(n6421), .Z(n4845) );
  IV U12637 ( .A(n8758), .Z(n6421) );
  XOR U12638 ( .A(n12856), .B(n12857), .Z(n8758) );
  ANDN U12639 ( .B(n8680), .A(n8681), .Z(n12855) );
  XNOR U12640 ( .A(n12858), .B(n10019), .Z(n8681) );
  XOR U12641 ( .A(n12859), .B(n10991), .Z(n8680) );
  XOR U12642 ( .A(n12860), .B(n6417), .Z(n8747) );
  XNOR U12643 ( .A(n12861), .B(n9692), .Z(n6417) );
  XOR U12644 ( .A(n12862), .B(n12863), .Z(n9692) );
  ANDN U12645 ( .B(n8675), .A(n8674), .Z(n12860) );
  XOR U12646 ( .A(n10539), .B(n12864), .Z(n8674) );
  XOR U12647 ( .A(n12865), .B(n10794), .Z(n8675) );
  XNOR U12648 ( .A(n12866), .B(n6430), .Z(n3463) );
  XOR U12649 ( .A(n12867), .B(n9388), .Z(n6430) );
  AND U12650 ( .A(n8670), .B(n8671), .Z(n12866) );
  XOR U12651 ( .A(n12868), .B(n12358), .Z(n8671) );
  XNOR U12652 ( .A(n10168), .B(n12869), .Z(n8670) );
  IV U12653 ( .A(n9494), .Z(n10168) );
  XNOR U12654 ( .A(n12870), .B(n12871), .Z(n6278) );
  XOR U12655 ( .A(n5419), .B(n3665), .Z(n12871) );
  XOR U12656 ( .A(n12872), .B(n12873), .Z(n3665) );
  AND U12657 ( .A(n6456), .B(n12874), .Z(n12872) );
  XOR U12658 ( .A(n12875), .B(n12876), .Z(n6456) );
  XNOR U12659 ( .A(n12877), .B(n8766), .Z(n5419) );
  ANDN U12660 ( .B(n6442), .A(n6443), .Z(n12877) );
  XOR U12661 ( .A(n12878), .B(n11590), .Z(n6443) );
  IV U12662 ( .A(n12358), .Z(n11590) );
  XOR U12663 ( .A(n10706), .B(n12879), .Z(n6442) );
  IV U12664 ( .A(n12880), .Z(n10706) );
  XNOR U12665 ( .A(n4282), .B(n12881), .Z(n12870) );
  XNOR U12666 ( .A(n5855), .B(n2112), .Z(n12881) );
  XNOR U12667 ( .A(n12882), .B(n8763), .Z(n2112) );
  ANDN U12668 ( .B(n6459), .A(n6460), .Z(n12882) );
  XOR U12669 ( .A(n12883), .B(n12884), .Z(n6460) );
  XNOR U12670 ( .A(n12885), .B(n10701), .Z(n6459) );
  IV U12671 ( .A(n12137), .Z(n10701) );
  XOR U12672 ( .A(n12886), .B(n8775), .Z(n5855) );
  AND U12673 ( .A(n6465), .B(n6463), .Z(n12886) );
  XOR U12674 ( .A(n12887), .B(n9358), .Z(n6463) );
  XOR U12675 ( .A(n12888), .B(n9917), .Z(n6465) );
  XNOR U12676 ( .A(n12889), .B(n8772), .Z(n4282) );
  AND U12677 ( .A(n6447), .B(n6446), .Z(n12889) );
  IV U12678 ( .A(n8771), .Z(n6446) );
  XNOR U12679 ( .A(n12890), .B(n10794), .Z(n8771) );
  XOR U12680 ( .A(n12891), .B(n11844), .Z(n10794) );
  XOR U12681 ( .A(n12892), .B(n12893), .Z(n11844) );
  XNOR U12682 ( .A(n12894), .B(n12895), .Z(n12893) );
  XOR U12683 ( .A(n12144), .B(n12896), .Z(n12892) );
  XNOR U12684 ( .A(n9089), .B(n11183), .Z(n12896) );
  XNOR U12685 ( .A(n12897), .B(n12898), .Z(n11183) );
  AND U12686 ( .A(n12899), .B(n12900), .Z(n12897) );
  XNOR U12687 ( .A(n12901), .B(n12902), .Z(n9089) );
  XNOR U12688 ( .A(n12905), .B(n12906), .Z(n12144) );
  AND U12689 ( .A(n12907), .B(n12908), .Z(n12905) );
  XNOR U12690 ( .A(n9383), .B(n12909), .Z(n6447) );
  IV U12691 ( .A(n11881), .Z(n9383) );
  XOR U12692 ( .A(n12910), .B(n8753), .Z(n8678) );
  IV U12693 ( .A(n12853), .Z(n8753) );
  XOR U12694 ( .A(n12911), .B(n11908), .Z(n12853) );
  NOR U12695 ( .A(n12651), .B(n6424), .Z(n12910) );
  XNOR U12696 ( .A(n12912), .B(n11072), .Z(n6424) );
  XNOR U12697 ( .A(n9170), .B(n12913), .Z(n12651) );
  IV U12698 ( .A(n10104), .Z(n9170) );
  XOR U12699 ( .A(n11222), .B(n2079), .Z(n5641) );
  XNOR U12700 ( .A(n8128), .B(n9440), .Z(n2079) );
  XNOR U12701 ( .A(n12914), .B(n12915), .Z(n9440) );
  XNOR U12702 ( .A(n5446), .B(n3578), .Z(n12915) );
  XOR U12703 ( .A(n12916), .B(n12917), .Z(n3578) );
  ANDN U12704 ( .B(n8284), .A(n8285), .Z(n12916) );
  XOR U12705 ( .A(n12918), .B(n10665), .Z(n8285) );
  XNOR U12706 ( .A(n12919), .B(n11343), .Z(n5446) );
  AND U12707 ( .A(n8282), .B(n8280), .Z(n12919) );
  IV U12708 ( .A(n11342), .Z(n8280) );
  XOR U12709 ( .A(n12920), .B(n12921), .Z(n11342) );
  XOR U12710 ( .A(n12922), .B(n12191), .Z(n8282) );
  XOR U12711 ( .A(n6237), .B(n12923), .Z(n12914) );
  XNOR U12712 ( .A(n2360), .B(n5512), .Z(n12923) );
  XNOR U12713 ( .A(n12924), .B(n11354), .Z(n5512) );
  AND U12714 ( .A(n9444), .B(n9442), .Z(n12924) );
  XOR U12715 ( .A(n12925), .B(n9587), .Z(n9442) );
  XNOR U12716 ( .A(n12926), .B(n12927), .Z(n9587) );
  XNOR U12717 ( .A(n12928), .B(n11695), .Z(n9444) );
  XNOR U12718 ( .A(n12929), .B(n11346), .Z(n2360) );
  ANDN U12719 ( .B(n8272), .A(n8270), .Z(n12929) );
  XOR U12720 ( .A(n12930), .B(n10599), .Z(n8270) );
  XNOR U12721 ( .A(n12931), .B(n9766), .Z(n8272) );
  XOR U12722 ( .A(n12932), .B(n11351), .Z(n6237) );
  ANDN U12723 ( .B(n8274), .A(n8275), .Z(n12932) );
  XNOR U12724 ( .A(n12933), .B(n11573), .Z(n8275) );
  XOR U12725 ( .A(n12934), .B(n12935), .Z(n11573) );
  XOR U12726 ( .A(n12880), .B(n12936), .Z(n8274) );
  XOR U12727 ( .A(n12937), .B(n12938), .Z(n8128) );
  XNOR U12728 ( .A(n3791), .B(n5112), .Z(n12938) );
  XNOR U12729 ( .A(n12939), .B(n9347), .Z(n5112) );
  XNOR U12730 ( .A(n11881), .B(n12940), .Z(n9347) );
  XOR U12731 ( .A(n12941), .B(n12942), .Z(n11881) );
  ANDN U12732 ( .B(n11228), .A(n11229), .Z(n12939) );
  XOR U12733 ( .A(n9684), .B(n12943), .Z(n11229) );
  XNOR U12734 ( .A(n12944), .B(n10599), .Z(n11228) );
  XOR U12735 ( .A(n12945), .B(n12200), .Z(n10599) );
  XOR U12736 ( .A(n12946), .B(n12947), .Z(n12200) );
  XNOR U12737 ( .A(n12948), .B(n10821), .Z(n12947) );
  XNOR U12738 ( .A(n12949), .B(n12950), .Z(n10821) );
  AND U12739 ( .A(n12951), .B(n12952), .Z(n12949) );
  XOR U12740 ( .A(n12039), .B(n12953), .Z(n12946) );
  XNOR U12741 ( .A(n9606), .B(n10543), .Z(n12953) );
  XNOR U12742 ( .A(n12954), .B(n12955), .Z(n10543) );
  AND U12743 ( .A(n12956), .B(n12957), .Z(n12954) );
  XNOR U12744 ( .A(n12958), .B(n12959), .Z(n9606) );
  ANDN U12745 ( .B(n12960), .A(n12961), .Z(n12958) );
  XNOR U12746 ( .A(n12962), .B(n12963), .Z(n12039) );
  AND U12747 ( .A(n12964), .B(n12965), .Z(n12962) );
  XNOR U12748 ( .A(n12966), .B(n8187), .Z(n3791) );
  XNOR U12749 ( .A(n12967), .B(n12176), .Z(n8187) );
  XNOR U12750 ( .A(n9892), .B(n12968), .Z(n11220) );
  XNOR U12751 ( .A(n12751), .B(n9668), .Z(n11221) );
  XNOR U12752 ( .A(n12969), .B(n12970), .Z(n12751) );
  AND U12753 ( .A(n12971), .B(n12972), .Z(n12969) );
  XNOR U12754 ( .A(n4352), .B(n12973), .Z(n12937) );
  XOR U12755 ( .A(n1728), .B(n11328), .Z(n12973) );
  XNOR U12756 ( .A(n12974), .B(n8198), .Z(n11328) );
  XNOR U12757 ( .A(n12975), .B(n11550), .Z(n8198) );
  XNOR U12758 ( .A(n12976), .B(n12977), .Z(n11550) );
  NOR U12759 ( .A(n11217), .B(n11216), .Z(n12974) );
  XNOR U12760 ( .A(n11686), .B(n12978), .Z(n11216) );
  XOR U12761 ( .A(n12979), .B(n12980), .Z(n11686) );
  XNOR U12762 ( .A(n12981), .B(n10712), .Z(n11217) );
  XNOR U12763 ( .A(n12982), .B(n8192), .Z(n1728) );
  XOR U12764 ( .A(n12983), .B(n10925), .Z(n8192) );
  XNOR U12765 ( .A(n9769), .B(n12984), .Z(n11226) );
  XOR U12766 ( .A(n12987), .B(n9529), .Z(n11225) );
  XNOR U12767 ( .A(n12988), .B(n8202), .Z(n4352) );
  XNOR U12768 ( .A(n12989), .B(n11570), .Z(n8202) );
  ANDN U12769 ( .B(n11335), .A(n12677), .Z(n12988) );
  XOR U12770 ( .A(n12990), .B(n11335), .Z(n11222) );
  XOR U12771 ( .A(n9558), .B(n12991), .Z(n11335) );
  AND U12772 ( .A(n12677), .B(n8200), .Z(n12990) );
  IV U12773 ( .A(n12678), .Z(n8200) );
  XOR U12774 ( .A(n12992), .B(n11522), .Z(n12678) );
  XNOR U12775 ( .A(n12993), .B(n12671), .Z(n12677) );
  XOR U12776 ( .A(n12994), .B(n6159), .Z(out[1003]) );
  IV U12777 ( .A(n6910), .Z(n6159) );
  XOR U12778 ( .A(n8927), .B(n2282), .Z(n6910) );
  XNOR U12779 ( .A(n6042), .B(n6123), .Z(n2282) );
  XNOR U12780 ( .A(n12995), .B(n12996), .Z(n6123) );
  XOR U12781 ( .A(n2322), .B(n5433), .Z(n12996) );
  XOR U12782 ( .A(n12997), .B(n7775), .Z(n5433) );
  XNOR U12783 ( .A(n12998), .B(n10065), .Z(n7775) );
  XNOR U12784 ( .A(n12467), .B(n12999), .Z(n10065) );
  XOR U12785 ( .A(n13000), .B(n13001), .Z(n12467) );
  XNOR U12786 ( .A(n12712), .B(n10583), .Z(n13001) );
  XNOR U12787 ( .A(n13002), .B(n13003), .Z(n10583) );
  ANDN U12788 ( .B(n13004), .A(n13005), .Z(n13002) );
  XOR U12789 ( .A(n13006), .B(n13007), .Z(n12712) );
  ANDN U12790 ( .B(n13008), .A(n13009), .Z(n13006) );
  XNOR U12791 ( .A(n11935), .B(n13010), .Z(n13000) );
  XOR U12792 ( .A(n13011), .B(n13012), .Z(n13010) );
  XNOR U12793 ( .A(n13013), .B(n13014), .Z(n11935) );
  AND U12794 ( .A(n13015), .B(n13016), .Z(n13013) );
  ANDN U12795 ( .B(n12825), .A(n7774), .Z(n12997) );
  XOR U12796 ( .A(n13017), .B(n13018), .Z(n7774) );
  XOR U12797 ( .A(n13019), .B(n9114), .Z(n12825) );
  IV U12798 ( .A(n9944), .Z(n9114) );
  XNOR U12799 ( .A(n13020), .B(n7779), .Z(n2322) );
  XNOR U12800 ( .A(n13021), .B(n9822), .Z(n7779) );
  IV U12801 ( .A(n9805), .Z(n9822) );
  NOR U12802 ( .A(n7778), .B(n8932), .Z(n13020) );
  XOR U12803 ( .A(n11418), .B(n13022), .Z(n8932) );
  XOR U12804 ( .A(n13023), .B(n12326), .Z(n11418) );
  XOR U12805 ( .A(n13024), .B(n13025), .Z(n12326) );
  XNOR U12806 ( .A(n9775), .B(n13026), .Z(n13025) );
  XOR U12807 ( .A(n13027), .B(n13015), .Z(n9775) );
  ANDN U12808 ( .B(n13028), .A(n13029), .Z(n13027) );
  XOR U12809 ( .A(n11380), .B(n13030), .Z(n13024) );
  XNOR U12810 ( .A(n10370), .B(n13031), .Z(n13030) );
  XNOR U12811 ( .A(n13032), .B(n13033), .Z(n10370) );
  XNOR U12812 ( .A(n13036), .B(n13005), .Z(n11380) );
  ANDN U12813 ( .B(n13037), .A(n13038), .Z(n13036) );
  XOR U12814 ( .A(n13039), .B(n13040), .Z(n7778) );
  XOR U12815 ( .A(n3151), .B(n13041), .Z(n12995) );
  XNOR U12816 ( .A(n6168), .B(n7768), .Z(n13041) );
  XOR U12817 ( .A(n13042), .B(n7784), .Z(n7768) );
  XOR U12818 ( .A(n13043), .B(n13044), .Z(n7784) );
  AND U12819 ( .A(n7783), .B(n8934), .Z(n13042) );
  XOR U12820 ( .A(n13045), .B(n9176), .Z(n8934) );
  XNOR U12821 ( .A(n13046), .B(n13047), .Z(n9176) );
  XNOR U12822 ( .A(n13048), .B(n10681), .Z(n7783) );
  XNOR U12823 ( .A(n13049), .B(n12295), .Z(n10681) );
  XNOR U12824 ( .A(n13050), .B(n13051), .Z(n12295) );
  XOR U12825 ( .A(n12185), .B(n13052), .Z(n13051) );
  XOR U12826 ( .A(n13053), .B(n13054), .Z(n12185) );
  ANDN U12827 ( .B(n13055), .A(n13056), .Z(n13053) );
  XNOR U12828 ( .A(n10108), .B(n13057), .Z(n13050) );
  XOR U12829 ( .A(n11259), .B(n11408), .Z(n13057) );
  XNOR U12830 ( .A(n13058), .B(n13059), .Z(n11408) );
  AND U12831 ( .A(n13060), .B(n13061), .Z(n13058) );
  XNOR U12832 ( .A(n13062), .B(n13063), .Z(n11259) );
  ANDN U12833 ( .B(n13064), .A(n13065), .Z(n13062) );
  XOR U12834 ( .A(n13066), .B(n13067), .Z(n10108) );
  AND U12835 ( .A(n13068), .B(n13069), .Z(n13066) );
  XNOR U12836 ( .A(n13070), .B(n7787), .Z(n6168) );
  XNOR U12837 ( .A(n13071), .B(n12604), .Z(n7787) );
  ANDN U12838 ( .B(n12837), .A(n7788), .Z(n13070) );
  XNOR U12839 ( .A(n13072), .B(n7791), .Z(n3151) );
  XOR U12840 ( .A(n13073), .B(n10679), .Z(n7791) );
  AND U12841 ( .A(n8929), .B(n7792), .Z(n13072) );
  XNOR U12842 ( .A(n13074), .B(n13075), .Z(n7792) );
  XNOR U12843 ( .A(n11593), .B(n13076), .Z(n8929) );
  XOR U12844 ( .A(n13077), .B(n13078), .Z(n6042) );
  XNOR U12845 ( .A(n5239), .B(n1935), .Z(n13078) );
  XOR U12846 ( .A(n13079), .B(n8993), .Z(n1935) );
  ANDN U12847 ( .B(n7857), .A(n8917), .Z(n13079) );
  XNOR U12848 ( .A(n13080), .B(n10277), .Z(n8917) );
  IV U12849 ( .A(n9824), .Z(n10277) );
  XNOR U12850 ( .A(n13081), .B(n13082), .Z(n9824) );
  XOR U12851 ( .A(n13083), .B(n11456), .Z(n7857) );
  XOR U12852 ( .A(n13084), .B(n9000), .Z(n5239) );
  ANDN U12853 ( .B(n7849), .A(n8915), .Z(n13084) );
  XOR U12854 ( .A(n12522), .B(n13085), .Z(n8915) );
  IV U12855 ( .A(n9177), .Z(n12522) );
  XOR U12856 ( .A(n11069), .B(n13086), .Z(n7849) );
  XOR U12857 ( .A(n13087), .B(n12264), .Z(n11069) );
  XNOR U12858 ( .A(n13088), .B(n13089), .Z(n12264) );
  XOR U12859 ( .A(n13090), .B(n11008), .Z(n13089) );
  XNOR U12860 ( .A(n13091), .B(n13092), .Z(n11008) );
  ANDN U12861 ( .B(n13093), .A(n13094), .Z(n13091) );
  XNOR U12862 ( .A(n11567), .B(n13095), .Z(n13088) );
  XOR U12863 ( .A(n12673), .B(n11699), .Z(n13095) );
  XNOR U12864 ( .A(n13096), .B(n13097), .Z(n11699) );
  ANDN U12865 ( .B(n13098), .A(n13099), .Z(n13096) );
  XNOR U12866 ( .A(n13100), .B(n13101), .Z(n12673) );
  ANDN U12867 ( .B(n13102), .A(n13103), .Z(n13100) );
  XOR U12868 ( .A(n13104), .B(n13105), .Z(n11567) );
  XNOR U12869 ( .A(n3690), .B(n13108), .Z(n13077) );
  XNOR U12870 ( .A(n8974), .B(n4164), .Z(n13108) );
  XOR U12871 ( .A(n13109), .B(n9002), .Z(n4164) );
  ANDN U12872 ( .B(n7840), .A(n8924), .Z(n13109) );
  XOR U12873 ( .A(n13110), .B(n10281), .Z(n8924) );
  XOR U12874 ( .A(n13111), .B(n13112), .Z(n10281) );
  XNOR U12875 ( .A(n13113), .B(n11855), .Z(n7840) );
  XNOR U12876 ( .A(n13114), .B(n8997), .Z(n8974) );
  ANDN U12877 ( .B(n8998), .A(n7844), .Z(n13114) );
  XOR U12878 ( .A(n13115), .B(n13116), .Z(n7844) );
  XOR U12879 ( .A(n9605), .B(n12948), .Z(n8998) );
  XNOR U12880 ( .A(n13117), .B(n13118), .Z(n12948) );
  AND U12881 ( .A(n13119), .B(n13120), .Z(n13117) );
  XOR U12882 ( .A(n11541), .B(n12785), .Z(n9605) );
  XNOR U12883 ( .A(n13121), .B(n13122), .Z(n12785) );
  XNOR U12884 ( .A(n13123), .B(n11879), .Z(n13122) );
  XNOR U12885 ( .A(n13124), .B(n13125), .Z(n11879) );
  ANDN U12886 ( .B(n12955), .A(n12956), .Z(n13124) );
  XOR U12887 ( .A(n11736), .B(n13126), .Z(n13121) );
  XOR U12888 ( .A(n11174), .B(n13127), .Z(n13126) );
  XOR U12889 ( .A(n13128), .B(n13129), .Z(n11174) );
  NOR U12890 ( .A(n12960), .B(n12959), .Z(n13128) );
  XNOR U12891 ( .A(n13130), .B(n13131), .Z(n11736) );
  ANDN U12892 ( .B(n12950), .A(n12951), .Z(n13130) );
  XOR U12893 ( .A(n13132), .B(n13133), .Z(n11541) );
  XNOR U12894 ( .A(n13134), .B(n11671), .Z(n13133) );
  XOR U12895 ( .A(n13135), .B(n13136), .Z(n11671) );
  ANDN U12896 ( .B(n13137), .A(n13138), .Z(n13135) );
  XOR U12897 ( .A(n11797), .B(n13139), .Z(n13132) );
  XNOR U12898 ( .A(n9538), .B(n12362), .Z(n13139) );
  XOR U12899 ( .A(n13140), .B(n13141), .Z(n12362) );
  ANDN U12900 ( .B(n13142), .A(n13143), .Z(n13140) );
  XOR U12901 ( .A(n13144), .B(n13145), .Z(n9538) );
  NOR U12902 ( .A(n13146), .B(n13147), .Z(n13144) );
  XOR U12903 ( .A(n13148), .B(n13149), .Z(n11797) );
  ANDN U12904 ( .B(n13150), .A(n13151), .Z(n13148) );
  XOR U12905 ( .A(n13152), .B(n13153), .Z(n3690) );
  ANDN U12906 ( .B(n8922), .A(n7853), .Z(n13152) );
  XNOR U12907 ( .A(n13154), .B(n10464), .Z(n7853) );
  XOR U12908 ( .A(n13155), .B(n7788), .Z(n8927) );
  XOR U12909 ( .A(n13156), .B(n11761), .Z(n7788) );
  NOR U12910 ( .A(n12837), .B(n8858), .Z(n13155) );
  XNOR U12911 ( .A(n13157), .B(n11456), .Z(n8858) );
  XOR U12912 ( .A(n11802), .B(n13158), .Z(n11456) );
  XOR U12913 ( .A(n13159), .B(n13160), .Z(n11802) );
  XNOR U12914 ( .A(n13161), .B(n10384), .Z(n13160) );
  XOR U12915 ( .A(n13162), .B(n13163), .Z(n10384) );
  AND U12916 ( .A(n13164), .B(n13165), .Z(n13162) );
  XOR U12917 ( .A(n12355), .B(n13166), .Z(n13159) );
  XOR U12918 ( .A(n11713), .B(n10248), .Z(n13166) );
  XOR U12919 ( .A(n13167), .B(n13168), .Z(n10248) );
  AND U12920 ( .A(n13169), .B(n13170), .Z(n13167) );
  XOR U12921 ( .A(n13171), .B(n13172), .Z(n11713) );
  NOR U12922 ( .A(n13173), .B(n13174), .Z(n13171) );
  XNOR U12923 ( .A(n13175), .B(n13176), .Z(n12355) );
  ANDN U12924 ( .B(n13177), .A(n13178), .Z(n13175) );
  XNOR U12925 ( .A(n13179), .B(n9353), .Z(n12837) );
  NOR U12926 ( .A(n5649), .B(n5648), .Z(n12994) );
  XNOR U12927 ( .A(n8768), .B(n3842), .Z(n5648) );
  XNOR U12928 ( .A(n6283), .B(n6411), .Z(n3842) );
  XNOR U12929 ( .A(n13180), .B(n13181), .Z(n6411) );
  XOR U12930 ( .A(n5081), .B(n2511), .Z(n13181) );
  XNOR U12931 ( .A(n13182), .B(n6464), .Z(n2511) );
  XNOR U12932 ( .A(n13183), .B(n11675), .Z(n6464) );
  ANDN U12933 ( .B(n8774), .A(n8775), .Z(n13182) );
  XNOR U12934 ( .A(n13184), .B(n11782), .Z(n8775) );
  XNOR U12935 ( .A(n13185), .B(n10920), .Z(n8774) );
  XNOR U12936 ( .A(n13186), .B(n6457), .Z(n5081) );
  XNOR U12937 ( .A(n13187), .B(n10010), .Z(n6457) );
  IV U12938 ( .A(n11766), .Z(n10010) );
  XNOR U12939 ( .A(n13188), .B(n13189), .Z(n11766) );
  ANDN U12940 ( .B(n13190), .A(n12873), .Z(n13186) );
  XNOR U12941 ( .A(n3466), .B(n13191), .Z(n13180) );
  XOR U12942 ( .A(n8811), .B(n4848), .Z(n13191) );
  XOR U12943 ( .A(n13192), .B(n6448), .Z(n4848) );
  XOR U12944 ( .A(n12510), .B(n12260), .Z(n6448) );
  XNOR U12945 ( .A(n13193), .B(n13194), .Z(n12510) );
  ANDN U12946 ( .B(n13195), .A(n13196), .Z(n13193) );
  AND U12947 ( .A(n8772), .B(n8816), .Z(n13192) );
  XNOR U12948 ( .A(n13197), .B(n11761), .Z(n8816) );
  XNOR U12949 ( .A(n13198), .B(n10121), .Z(n8772) );
  XOR U12950 ( .A(n13199), .B(n12934), .Z(n10121) );
  XOR U12951 ( .A(n13200), .B(n13201), .Z(n12934) );
  XNOR U12952 ( .A(n10779), .B(n9685), .Z(n13201) );
  XOR U12953 ( .A(n13202), .B(n13203), .Z(n9685) );
  XNOR U12954 ( .A(n13206), .B(n13207), .Z(n10779) );
  AND U12955 ( .A(n13208), .B(n13209), .Z(n13206) );
  XOR U12956 ( .A(n12943), .B(n13210), .Z(n13200) );
  XOR U12957 ( .A(n12521), .B(n13211), .Z(n13210) );
  XOR U12958 ( .A(n13212), .B(n13213), .Z(n12521) );
  ANDN U12959 ( .B(n13214), .A(n13215), .Z(n13212) );
  XNOR U12960 ( .A(n13216), .B(n13217), .Z(n12943) );
  AND U12961 ( .A(n13218), .B(n13219), .Z(n13216) );
  XNOR U12962 ( .A(n13220), .B(n6444), .Z(n8811) );
  XOR U12963 ( .A(n13221), .B(n9800), .Z(n6444) );
  XNOR U12964 ( .A(n13222), .B(n13223), .Z(n9800) );
  ANDN U12965 ( .B(n8765), .A(n8766), .Z(n13220) );
  XNOR U12966 ( .A(n13224), .B(n11052), .Z(n8766) );
  XNOR U12967 ( .A(n13225), .B(n9181), .Z(n8765) );
  IV U12968 ( .A(n10661), .Z(n9181) );
  XNOR U12969 ( .A(n13227), .B(n13228), .Z(n11525) );
  XOR U12970 ( .A(n13229), .B(n13076), .Z(n13228) );
  XOR U12971 ( .A(n13230), .B(n13231), .Z(n13076) );
  ANDN U12972 ( .B(n13232), .A(n13233), .Z(n13230) );
  XNOR U12973 ( .A(n13234), .B(n13235), .Z(n13227) );
  XOR U12974 ( .A(n11692), .B(n11594), .Z(n13235) );
  XOR U12975 ( .A(n13236), .B(n13237), .Z(n11594) );
  AND U12976 ( .A(n13238), .B(n13239), .Z(n13236) );
  XOR U12977 ( .A(n13240), .B(n13241), .Z(n11692) );
  ANDN U12978 ( .B(n13242), .A(n13243), .Z(n13240) );
  XOR U12979 ( .A(n13244), .B(n6461), .Z(n3466) );
  XOR U12980 ( .A(n13245), .B(n9519), .Z(n6461) );
  XNOR U12981 ( .A(n13246), .B(n12711), .Z(n9519) );
  XNOR U12982 ( .A(n13247), .B(n13248), .Z(n12711) );
  XOR U12983 ( .A(n12740), .B(n9932), .Z(n13248) );
  XNOR U12984 ( .A(n13249), .B(n13250), .Z(n9932) );
  ANDN U12985 ( .B(n13251), .A(n13252), .Z(n13249) );
  XOR U12986 ( .A(n13253), .B(n13254), .Z(n12740) );
  ANDN U12987 ( .B(n13255), .A(n13256), .Z(n13253) );
  XOR U12988 ( .A(n13257), .B(n13258), .Z(n13247) );
  XOR U12989 ( .A(n12233), .B(n9167), .Z(n13258) );
  XNOR U12990 ( .A(n13259), .B(n13260), .Z(n9167) );
  AND U12991 ( .A(n13261), .B(n13262), .Z(n13259) );
  XOR U12992 ( .A(n13263), .B(n13264), .Z(n12233) );
  AND U12993 ( .A(n13265), .B(n13266), .Z(n13263) );
  AND U12994 ( .A(n8763), .B(n8821), .Z(n13244) );
  XOR U12995 ( .A(n13267), .B(n9573), .Z(n8821) );
  XNOR U12996 ( .A(n13268), .B(n11916), .Z(n8763) );
  XNOR U12997 ( .A(n13269), .B(n13270), .Z(n6283) );
  XOR U12998 ( .A(n5423), .B(n3669), .Z(n13270) );
  XOR U12999 ( .A(n13271), .B(n13272), .Z(n3669) );
  ANDN U13000 ( .B(n6481), .A(n6482), .Z(n13271) );
  XNOR U13001 ( .A(n13273), .B(n10920), .Z(n6482) );
  XNOR U13002 ( .A(n13274), .B(n8830), .Z(n5423) );
  AND U13003 ( .A(n6473), .B(n8831), .Z(n13274) );
  XNOR U13004 ( .A(n13275), .B(n10806), .Z(n8831) );
  XNOR U13005 ( .A(n13276), .B(n11916), .Z(n6473) );
  XOR U13006 ( .A(n4285), .B(n13277), .Z(n13269) );
  XOR U13007 ( .A(n5860), .B(n2115), .Z(n13277) );
  XOR U13008 ( .A(n13278), .B(n8827), .Z(n2115) );
  NOR U13009 ( .A(n6486), .B(n6485), .Z(n13278) );
  XNOR U13010 ( .A(n9480), .B(n13279), .Z(n6485) );
  XOR U13011 ( .A(n13280), .B(n10590), .Z(n6486) );
  XOR U13012 ( .A(n13281), .B(n8839), .Z(n5860) );
  AND U13013 ( .A(n6490), .B(n6489), .Z(n13281) );
  XNOR U13014 ( .A(n9101), .B(n13282), .Z(n6489) );
  XNOR U13015 ( .A(n13283), .B(n11793), .Z(n6490) );
  XNOR U13016 ( .A(n13284), .B(n8836), .Z(n4285) );
  AND U13017 ( .A(n6476), .B(n6477), .Z(n13284) );
  XNOR U13018 ( .A(n13285), .B(n13286), .Z(n6477) );
  XNOR U13019 ( .A(n13287), .B(n11052), .Z(n6476) );
  IV U13020 ( .A(n11695), .Z(n11052) );
  XOR U13021 ( .A(n13288), .B(n11790), .Z(n11695) );
  XNOR U13022 ( .A(n13289), .B(n13290), .Z(n11790) );
  XNOR U13023 ( .A(n13291), .B(n12265), .Z(n13290) );
  XNOR U13024 ( .A(n13292), .B(n13293), .Z(n12265) );
  AND U13025 ( .A(n13294), .B(n13295), .Z(n13292) );
  XNOR U13026 ( .A(n12293), .B(n13296), .Z(n13289) );
  XOR U13027 ( .A(n9073), .B(n11308), .Z(n13296) );
  XNOR U13028 ( .A(n13297), .B(n13298), .Z(n11308) );
  AND U13029 ( .A(n13299), .B(n13300), .Z(n13297) );
  XNOR U13030 ( .A(n13301), .B(n13302), .Z(n9073) );
  ANDN U13031 ( .B(n13303), .A(n13304), .Z(n13301) );
  XNOR U13032 ( .A(n13305), .B(n13306), .Z(n12293) );
  AND U13033 ( .A(n13307), .B(n13308), .Z(n13305) );
  XOR U13034 ( .A(n13309), .B(n8819), .Z(n8768) );
  IV U13035 ( .A(n13190), .Z(n8819) );
  XNOR U13036 ( .A(n13310), .B(n12069), .Z(n13190) );
  AND U13037 ( .A(n12873), .B(n6450), .Z(n13309) );
  IV U13038 ( .A(n12874), .Z(n6450) );
  XOR U13039 ( .A(n11777), .B(n13311), .Z(n12874) );
  IV U13040 ( .A(n11198), .Z(n11777) );
  XOR U13041 ( .A(n13312), .B(n13313), .Z(n11198) );
  XNOR U13042 ( .A(n13314), .B(n10215), .Z(n12873) );
  IV U13043 ( .A(n13315), .Z(n10215) );
  XOR U13044 ( .A(n11347), .B(n2082), .Z(n5649) );
  XNOR U13045 ( .A(n8182), .B(n9542), .Z(n2082) );
  XNOR U13046 ( .A(n13316), .B(n13317), .Z(n9542) );
  XNOR U13047 ( .A(n5450), .B(n3582), .Z(n13317) );
  XOR U13048 ( .A(n13318), .B(n13319), .Z(n3582) );
  ANDN U13049 ( .B(n8336), .A(n8337), .Z(n13318) );
  XNOR U13050 ( .A(n10730), .B(n13320), .Z(n8337) );
  XNOR U13051 ( .A(n13321), .B(n11482), .Z(n5450) );
  ANDN U13052 ( .B(n8332), .A(n8334), .Z(n13321) );
  XOR U13053 ( .A(n13161), .B(n10249), .Z(n8334) );
  XNOR U13054 ( .A(n13322), .B(n13323), .Z(n10249) );
  XNOR U13055 ( .A(n13324), .B(n13325), .Z(n13161) );
  AND U13056 ( .A(n13326), .B(n13327), .Z(n13324) );
  XNOR U13057 ( .A(n13328), .B(n13329), .Z(n8332) );
  XOR U13058 ( .A(n6241), .B(n13330), .Z(n13316) );
  XNOR U13059 ( .A(n2367), .B(n5554), .Z(n13330) );
  XNOR U13060 ( .A(n13331), .B(n11493), .Z(n5554) );
  AND U13061 ( .A(n9546), .B(n11494), .Z(n13331) );
  XNOR U13062 ( .A(n13332), .B(n9697), .Z(n11494) );
  XOR U13063 ( .A(n13333), .B(n12828), .Z(n9697) );
  XOR U13064 ( .A(n13334), .B(n13335), .Z(n12828) );
  XNOR U13065 ( .A(n12064), .B(n11638), .Z(n13335) );
  XOR U13066 ( .A(n13336), .B(n13337), .Z(n11638) );
  AND U13067 ( .A(n13338), .B(n13339), .Z(n13336) );
  XNOR U13068 ( .A(n13340), .B(n13341), .Z(n12064) );
  AND U13069 ( .A(n13342), .B(n13343), .Z(n13340) );
  XNOR U13070 ( .A(n11740), .B(n13344), .Z(n13334) );
  XNOR U13071 ( .A(n12090), .B(n11680), .Z(n13344) );
  XNOR U13072 ( .A(n13345), .B(n13346), .Z(n11680) );
  ANDN U13073 ( .B(n13347), .A(n13348), .Z(n13345) );
  XNOR U13074 ( .A(n13349), .B(n13350), .Z(n12090) );
  ANDN U13075 ( .B(n13351), .A(n13352), .Z(n13349) );
  XOR U13076 ( .A(n13353), .B(n13354), .Z(n11740) );
  AND U13077 ( .A(n13355), .B(n13356), .Z(n13353) );
  XOR U13078 ( .A(n13357), .B(n11065), .Z(n9546) );
  XNOR U13079 ( .A(n13358), .B(n11485), .Z(n2367) );
  ANDN U13080 ( .B(n8322), .A(n8323), .Z(n13358) );
  XNOR U13081 ( .A(n13359), .B(n13360), .Z(n8323) );
  XNOR U13082 ( .A(n13127), .B(n11880), .Z(n8322) );
  XOR U13083 ( .A(n13361), .B(n13362), .Z(n13127) );
  AND U13084 ( .A(n12963), .B(n13363), .Z(n13361) );
  XNOR U13085 ( .A(n13364), .B(n11490), .Z(n6241) );
  ANDN U13086 ( .B(n8328), .A(n8326), .Z(n13364) );
  XOR U13087 ( .A(n13365), .B(n10806), .Z(n8326) );
  XOR U13088 ( .A(n11890), .B(n13366), .Z(n8328) );
  IV U13089 ( .A(n11433), .Z(n11890) );
  XOR U13090 ( .A(n13367), .B(n13368), .Z(n11433) );
  XOR U13091 ( .A(n13369), .B(n13370), .Z(n8182) );
  XNOR U13092 ( .A(n3796), .B(n5114), .Z(n13370) );
  XOR U13093 ( .A(n13371), .B(n9443), .Z(n5114) );
  XNOR U13094 ( .A(n13372), .B(n13286), .Z(n9443) );
  IV U13095 ( .A(n9524), .Z(n13286) );
  XNOR U13096 ( .A(n13373), .B(n13374), .Z(n9524) );
  NOR U13097 ( .A(n11354), .B(n11353), .Z(n13371) );
  XNOR U13098 ( .A(n13123), .B(n11175), .Z(n11353) );
  IV U13099 ( .A(n11880), .Z(n11175) );
  XOR U13100 ( .A(n13375), .B(n13376), .Z(n11880) );
  XOR U13101 ( .A(n13377), .B(n13378), .Z(n13123) );
  AND U13102 ( .A(n13118), .B(n13379), .Z(n13377) );
  XOR U13103 ( .A(n13380), .B(n9077), .Z(n11354) );
  XOR U13104 ( .A(n13381), .B(n13382), .Z(n9077) );
  XNOR U13105 ( .A(n13383), .B(n8271), .Z(n3796) );
  XNOR U13106 ( .A(n13384), .B(n10048), .Z(n8271) );
  IV U13107 ( .A(n12832), .Z(n10048) );
  ANDN U13108 ( .B(n11345), .A(n11346), .Z(n13383) );
  XNOR U13109 ( .A(n13031), .B(n9776), .Z(n11346) );
  XNOR U13110 ( .A(n13387), .B(n13009), .Z(n13031) );
  AND U13111 ( .A(n13388), .B(n13389), .Z(n13387) );
  XNOR U13112 ( .A(n13390), .B(n13391), .Z(n11345) );
  XOR U13113 ( .A(n4753), .B(n13392), .Z(n13369) );
  XNOR U13114 ( .A(n1732), .B(n11467), .Z(n13392) );
  XNOR U13115 ( .A(n13393), .B(n11477), .Z(n11467) );
  IV U13116 ( .A(n8281), .Z(n11477) );
  XOR U13117 ( .A(n13394), .B(n10823), .Z(n8281) );
  IV U13118 ( .A(n11684), .Z(n10823) );
  ANDN U13119 ( .B(n11343), .A(n11341), .Z(n13393) );
  XNOR U13120 ( .A(n12005), .B(n13397), .Z(n11341) );
  XOR U13121 ( .A(n12559), .B(n13398), .Z(n12005) );
  XOR U13122 ( .A(n13399), .B(n13400), .Z(n12559) );
  XNOR U13123 ( .A(n13401), .B(n13402), .Z(n13400) );
  XNOR U13124 ( .A(n12388), .B(n13403), .Z(n13399) );
  XNOR U13125 ( .A(n12468), .B(n9118), .Z(n13403) );
  XNOR U13126 ( .A(n13404), .B(n13405), .Z(n9118) );
  AND U13127 ( .A(n13406), .B(n13407), .Z(n13404) );
  XNOR U13128 ( .A(n13408), .B(n13409), .Z(n12468) );
  AND U13129 ( .A(n13410), .B(n13411), .Z(n13408) );
  XNOR U13130 ( .A(n13412), .B(n13413), .Z(n12388) );
  ANDN U13131 ( .B(n13414), .A(n13415), .Z(n13412) );
  XNOR U13132 ( .A(n13416), .B(n10174), .Z(n11343) );
  XNOR U13133 ( .A(n13417), .B(n13418), .Z(n10174) );
  XNOR U13134 ( .A(n13419), .B(n8276), .Z(n1732) );
  XNOR U13135 ( .A(n13420), .B(n11015), .Z(n8276) );
  IV U13136 ( .A(n13421), .Z(n11015) );
  AND U13137 ( .A(n11350), .B(n11351), .Z(n13419) );
  XOR U13138 ( .A(n9892), .B(n13422), .Z(n11351) );
  XOR U13139 ( .A(n13423), .B(n9353), .Z(n11350) );
  XOR U13140 ( .A(n13424), .B(n12318), .Z(n9353) );
  XOR U13141 ( .A(n13425), .B(n13426), .Z(n12318) );
  XNOR U13142 ( .A(n13427), .B(n12729), .Z(n13426) );
  XOR U13143 ( .A(n13428), .B(n13429), .Z(n12729) );
  ANDN U13144 ( .B(n13430), .A(n13431), .Z(n13428) );
  XOR U13145 ( .A(n13432), .B(n13433), .Z(n13425) );
  XNOR U13146 ( .A(n12268), .B(n11387), .Z(n13433) );
  XNOR U13147 ( .A(n13434), .B(n13435), .Z(n11387) );
  AND U13148 ( .A(n13436), .B(n13437), .Z(n13434) );
  XNOR U13149 ( .A(n13438), .B(n13439), .Z(n12268) );
  ANDN U13150 ( .B(n13440), .A(n13441), .Z(n13438) );
  XNOR U13151 ( .A(n13442), .B(n8286), .Z(n4753) );
  XNOR U13152 ( .A(n13443), .B(n13329), .Z(n8286) );
  AND U13153 ( .A(n11474), .B(n12917), .Z(n13442) );
  IV U13154 ( .A(n13444), .Z(n12917) );
  XOR U13155 ( .A(n13445), .B(n11474), .Z(n11347) );
  XOR U13156 ( .A(n12745), .B(n9668), .Z(n11474) );
  XOR U13157 ( .A(n13081), .B(n13446), .Z(n9668) );
  XOR U13158 ( .A(n13447), .B(n13448), .Z(n13081) );
  XNOR U13159 ( .A(n10777), .B(n12150), .Z(n13448) );
  XOR U13160 ( .A(n13449), .B(n13450), .Z(n12150) );
  ANDN U13161 ( .B(n13451), .A(n13452), .Z(n13449) );
  XNOR U13162 ( .A(n13453), .B(n13454), .Z(n10777) );
  XOR U13163 ( .A(n9557), .B(n13455), .Z(n13447) );
  XOR U13164 ( .A(n9482), .B(n12325), .Z(n13455) );
  XOR U13165 ( .A(n13456), .B(n13457), .Z(n12325) );
  NOR U13166 ( .A(n12971), .B(n12970), .Z(n13456) );
  XOR U13167 ( .A(n13458), .B(n13459), .Z(n9482) );
  ANDN U13168 ( .B(n13460), .A(n12753), .Z(n13458) );
  XNOR U13169 ( .A(n13461), .B(n13462), .Z(n9557) );
  XNOR U13170 ( .A(n13463), .B(n13452), .Z(n12745) );
  ANDN U13171 ( .B(n13464), .A(n13465), .Z(n13463) );
  ANDN U13172 ( .B(n13444), .A(n8284), .Z(n13445) );
  XOR U13173 ( .A(n13466), .B(n9103), .Z(n8284) );
  IV U13174 ( .A(n10003), .Z(n9103) );
  XOR U13175 ( .A(n13467), .B(n13468), .Z(n10003) );
  XOR U13176 ( .A(n13469), .B(n11908), .Z(n13444) );
  XOR U13177 ( .A(n13470), .B(n6164), .Z(out[1002]) );
  IV U13178 ( .A(n6934), .Z(n6164) );
  XOR U13179 ( .A(n8991), .B(n2289), .Z(n6934) );
  XNOR U13180 ( .A(n6047), .B(n6128), .Z(n2289) );
  XNOR U13181 ( .A(n13471), .B(n13472), .Z(n6128) );
  XNOR U13182 ( .A(n2327), .B(n5438), .Z(n13472) );
  XOR U13183 ( .A(n13473), .B(n7842), .Z(n5438) );
  XNOR U13184 ( .A(n13474), .B(n10172), .Z(n7842) );
  XOR U13185 ( .A(n13446), .B(n12719), .Z(n10172) );
  XOR U13186 ( .A(n13475), .B(n13476), .Z(n12719) );
  XNOR U13187 ( .A(n12981), .B(n10711), .Z(n13476) );
  XOR U13188 ( .A(n13477), .B(n13478), .Z(n10711) );
  AND U13189 ( .A(n13479), .B(n13480), .Z(n13477) );
  XNOR U13190 ( .A(n13481), .B(n13482), .Z(n12981) );
  ANDN U13191 ( .B(n13483), .A(n13484), .Z(n13481) );
  XOR U13192 ( .A(n12124), .B(n13485), .Z(n13475) );
  XOR U13193 ( .A(n13486), .B(n13487), .Z(n13485) );
  XOR U13194 ( .A(n13488), .B(n13489), .Z(n12124) );
  AND U13195 ( .A(n13490), .B(n13491), .Z(n13488) );
  XOR U13196 ( .A(n13492), .B(n13493), .Z(n13446) );
  XOR U13197 ( .A(n12194), .B(n13022), .Z(n13493) );
  XOR U13198 ( .A(n13494), .B(n13035), .Z(n13022) );
  AND U13199 ( .A(n13495), .B(n13496), .Z(n13494) );
  XNOR U13200 ( .A(n13497), .B(n13029), .Z(n12194) );
  AND U13201 ( .A(n13014), .B(n13498), .Z(n13497) );
  XNOR U13202 ( .A(n11419), .B(n13499), .Z(n13492) );
  XOR U13203 ( .A(n12646), .B(n12655), .Z(n13499) );
  XNOR U13204 ( .A(n13500), .B(n13038), .Z(n12655) );
  ANDN U13205 ( .B(n13003), .A(n13037), .Z(n13500) );
  XNOR U13206 ( .A(n13501), .B(n13502), .Z(n12646) );
  XOR U13207 ( .A(n13505), .B(n13388), .Z(n11419) );
  ANDN U13208 ( .B(n13506), .A(n13007), .Z(n13505) );
  NOR U13209 ( .A(n7841), .B(n9002), .Z(n13473) );
  XNOR U13210 ( .A(n13507), .B(n9950), .Z(n9002) );
  XNOR U13211 ( .A(n13508), .B(n10590), .Z(n7841) );
  XNOR U13212 ( .A(n13509), .B(n7845), .Z(n2327) );
  XOR U13213 ( .A(n13510), .B(n9944), .Z(n7845) );
  AND U13214 ( .A(n8997), .B(n8996), .Z(n13509) );
  XOR U13215 ( .A(n13513), .B(n10055), .Z(n8996) );
  XOR U13216 ( .A(n13514), .B(n12358), .Z(n8997) );
  XOR U13217 ( .A(n12466), .B(n13418), .Z(n12358) );
  XNOR U13218 ( .A(n13515), .B(n13516), .Z(n13418) );
  XNOR U13219 ( .A(n11539), .B(n12070), .Z(n13516) );
  XOR U13220 ( .A(n13517), .B(n13518), .Z(n12070) );
  XNOR U13221 ( .A(n13521), .B(n13522), .Z(n11539) );
  AND U13222 ( .A(n13523), .B(n13524), .Z(n13521) );
  XNOR U13223 ( .A(n13525), .B(n13526), .Z(n13515) );
  XOR U13224 ( .A(n11812), .B(n13527), .Z(n13526) );
  XOR U13225 ( .A(n13528), .B(n13529), .Z(n11812) );
  ANDN U13226 ( .B(n13530), .A(n13531), .Z(n13528) );
  XOR U13227 ( .A(n13532), .B(n13533), .Z(n12466) );
  XNOR U13228 ( .A(n9899), .B(n13534), .Z(n13533) );
  XOR U13229 ( .A(n13535), .B(n13491), .Z(n9899) );
  IV U13230 ( .A(n13536), .Z(n13491) );
  AND U13231 ( .A(n13537), .B(n13538), .Z(n13535) );
  XNOR U13232 ( .A(n11514), .B(n13539), .Z(n13532) );
  XOR U13233 ( .A(n10551), .B(n13540), .Z(n13539) );
  XOR U13234 ( .A(n13541), .B(n13542), .Z(n10551) );
  ANDN U13235 ( .B(n13543), .A(n13544), .Z(n13541) );
  XNOR U13236 ( .A(n13545), .B(n13480), .Z(n11514) );
  AND U13237 ( .A(n13546), .B(n13547), .Z(n13545) );
  XNOR U13238 ( .A(n3154), .B(n13548), .Z(n13471) );
  XNOR U13239 ( .A(n6214), .B(n7835), .Z(n13548) );
  XNOR U13240 ( .A(n13549), .B(n7850), .Z(n7835) );
  XOR U13241 ( .A(n13550), .B(n9213), .Z(n7850) );
  ANDN U13242 ( .B(n7851), .A(n9000), .Z(n13549) );
  XOR U13243 ( .A(n13551), .B(n10783), .Z(n9000) );
  XOR U13244 ( .A(n13552), .B(n10903), .Z(n7851) );
  IV U13245 ( .A(n12876), .Z(n10903) );
  XNOR U13246 ( .A(n13553), .B(n13554), .Z(n12876) );
  XNOR U13247 ( .A(n13555), .B(n7855), .Z(n6214) );
  XOR U13248 ( .A(n12508), .B(n12260), .Z(n7855) );
  XOR U13249 ( .A(n13556), .B(n13557), .Z(n12418) );
  XOR U13250 ( .A(n11969), .B(n13558), .Z(n13557) );
  XOR U13251 ( .A(n13559), .B(n13560), .Z(n11969) );
  ANDN U13252 ( .B(n13561), .A(n12505), .Z(n13559) );
  XOR U13253 ( .A(n9260), .B(n13562), .Z(n13556) );
  XOR U13254 ( .A(n9813), .B(n12658), .Z(n13562) );
  XOR U13255 ( .A(n13563), .B(n13564), .Z(n12658) );
  ANDN U13256 ( .B(n12486), .A(n12487), .Z(n13563) );
  XNOR U13257 ( .A(n13565), .B(n13566), .Z(n9813) );
  XNOR U13258 ( .A(n13567), .B(n13568), .Z(n9260) );
  XNOR U13259 ( .A(n13569), .B(n13570), .Z(n11075) );
  XNOR U13260 ( .A(n11786), .B(n11912), .Z(n13570) );
  XOR U13261 ( .A(n13571), .B(n13572), .Z(n11912) );
  NOR U13262 ( .A(n12801), .B(n12802), .Z(n13571) );
  XNOR U13263 ( .A(n13573), .B(n13574), .Z(n11786) );
  XOR U13264 ( .A(n10699), .B(n13575), .Z(n13569) );
  XOR U13265 ( .A(n9675), .B(n11598), .Z(n13575) );
  XNOR U13266 ( .A(n13576), .B(n13577), .Z(n11598) );
  AND U13267 ( .A(n12519), .B(n12517), .Z(n13576) );
  XNOR U13268 ( .A(n13578), .B(n13579), .Z(n9675) );
  XOR U13269 ( .A(n13580), .B(n13581), .Z(n10699) );
  NOR U13270 ( .A(n13582), .B(n13583), .Z(n13580) );
  XNOR U13271 ( .A(n13584), .B(n13583), .Z(n12508) );
  ANDN U13272 ( .B(n13582), .A(n13585), .Z(n13584) );
  NOR U13273 ( .A(n7854), .B(n13153), .Z(n13555) );
  XNOR U13274 ( .A(n13586), .B(n7859), .Z(n3154) );
  XOR U13275 ( .A(n12553), .B(n13587), .Z(n7859) );
  XOR U13276 ( .A(n13588), .B(n13589), .Z(n12553) );
  ANDN U13277 ( .B(n7858), .A(n8993), .Z(n13586) );
  XOR U13278 ( .A(n10044), .B(n13590), .Z(n8993) );
  XOR U13279 ( .A(n13591), .B(n10226), .Z(n7858) );
  XOR U13280 ( .A(n13592), .B(n13593), .Z(n6047) );
  XOR U13281 ( .A(n5241), .B(n1940), .Z(n13593) );
  XNOR U13282 ( .A(n13594), .B(n9040), .Z(n1940) );
  AND U13283 ( .A(n7966), .B(n8980), .Z(n13594) );
  XOR U13284 ( .A(n13595), .B(n9946), .Z(n8980) );
  XNOR U13285 ( .A(n13596), .B(n11570), .Z(n7966) );
  IV U13286 ( .A(n12921), .Z(n11570) );
  XNOR U13287 ( .A(n13597), .B(n9046), .Z(n5241) );
  ANDN U13288 ( .B(n7958), .A(n8978), .Z(n13597) );
  XNOR U13289 ( .A(n13598), .B(n12662), .Z(n8978) );
  XNOR U13290 ( .A(n13599), .B(n11197), .Z(n7958) );
  XOR U13291 ( .A(n13600), .B(n13601), .Z(n11197) );
  XOR U13292 ( .A(n3695), .B(n13602), .Z(n13592) );
  XOR U13293 ( .A(n9035), .B(n4167), .Z(n13602) );
  XNOR U13294 ( .A(n13603), .B(n9048), .Z(n4167) );
  AND U13295 ( .A(n8987), .B(n8988), .Z(n13603) );
  XOR U13296 ( .A(n10110), .B(n13604), .Z(n8988) );
  XNOR U13297 ( .A(n13605), .B(n10464), .Z(n8987) );
  XNOR U13298 ( .A(n13606), .B(n13607), .Z(n10464) );
  XNOR U13299 ( .A(n13608), .B(n9044), .Z(n9035) );
  ANDN U13300 ( .B(n7953), .A(n8983), .Z(n13608) );
  XNOR U13301 ( .A(n13609), .B(n9716), .Z(n8983) );
  XNOR U13302 ( .A(n11678), .B(n13047), .Z(n9716) );
  XNOR U13303 ( .A(n13610), .B(n13611), .Z(n13047) );
  XOR U13304 ( .A(n13612), .B(n12044), .Z(n13611) );
  XNOR U13305 ( .A(n13613), .B(n13614), .Z(n12044) );
  AND U13306 ( .A(n13615), .B(n13145), .Z(n13613) );
  XNOR U13307 ( .A(n13616), .B(n13617), .Z(n13610) );
  XOR U13308 ( .A(n10828), .B(n11302), .Z(n13617) );
  XOR U13309 ( .A(n13618), .B(n13619), .Z(n11302) );
  AND U13310 ( .A(n13149), .B(n13620), .Z(n13618) );
  XOR U13311 ( .A(n13621), .B(n13622), .Z(n10828) );
  AND U13312 ( .A(n13136), .B(n13623), .Z(n13621) );
  XOR U13313 ( .A(n13624), .B(n13625), .Z(n11678) );
  XOR U13314 ( .A(n11992), .B(n10028), .Z(n13625) );
  XOR U13315 ( .A(n13626), .B(n13627), .Z(n10028) );
  NOR U13316 ( .A(n13628), .B(n13629), .Z(n13626) );
  XOR U13317 ( .A(n13630), .B(n13631), .Z(n11992) );
  XOR U13318 ( .A(n11235), .B(n13634), .Z(n13624) );
  XOR U13319 ( .A(n9607), .B(n12596), .Z(n13634) );
  XOR U13320 ( .A(n13635), .B(n13636), .Z(n12596) );
  AND U13321 ( .A(n13637), .B(n13638), .Z(n13635) );
  XOR U13322 ( .A(n13639), .B(n13640), .Z(n9607) );
  AND U13323 ( .A(n13641), .B(n13642), .Z(n13639) );
  XOR U13324 ( .A(n13643), .B(n13644), .Z(n11235) );
  XNOR U13325 ( .A(n13647), .B(n13648), .Z(n7953) );
  XNOR U13326 ( .A(n13649), .B(n13650), .Z(n3695) );
  AND U13327 ( .A(n7962), .B(n13651), .Z(n13649) );
  XNOR U13328 ( .A(n12397), .B(n11894), .Z(n7962) );
  XOR U13329 ( .A(n13652), .B(n13653), .Z(n12397) );
  AND U13330 ( .A(n13654), .B(n13655), .Z(n13652) );
  XOR U13331 ( .A(n13656), .B(n7854), .Z(n8991) );
  XOR U13332 ( .A(n11257), .B(n13657), .Z(n7854) );
  ANDN U13333 ( .B(n13153), .A(n8922), .Z(n13656) );
  XOR U13334 ( .A(n13658), .B(n12921), .Z(n8922) );
  XNOR U13335 ( .A(n13659), .B(n11132), .Z(n12921) );
  XNOR U13336 ( .A(n13660), .B(n13661), .Z(n11132) );
  XNOR U13337 ( .A(n13662), .B(n10563), .Z(n13661) );
  XOR U13338 ( .A(n13663), .B(n13664), .Z(n10563) );
  XOR U13339 ( .A(n10380), .B(n13667), .Z(n13660) );
  XOR U13340 ( .A(n11058), .B(n12589), .Z(n13667) );
  XNOR U13341 ( .A(n13668), .B(n13669), .Z(n12589) );
  AND U13342 ( .A(n13670), .B(n13671), .Z(n13668) );
  XNOR U13343 ( .A(n13672), .B(n13673), .Z(n11058) );
  ANDN U13344 ( .B(n13674), .A(n13675), .Z(n13672) );
  XNOR U13345 ( .A(n13676), .B(n13677), .Z(n10380) );
  XNOR U13346 ( .A(n9485), .B(n13680), .Z(n13153) );
  ANDN U13347 ( .B(n5654), .A(n5652), .Z(n13470) );
  XNOR U13348 ( .A(n8833), .B(n5142), .Z(n5652) );
  XNOR U13349 ( .A(n13681), .B(n13682), .Z(n6438) );
  XNOR U13350 ( .A(n5464), .B(n2520), .Z(n13682) );
  XNOR U13351 ( .A(n13683), .B(n6491), .Z(n2520) );
  XNOR U13352 ( .A(n12762), .B(n13684), .Z(n6491) );
  IV U13353 ( .A(n11926), .Z(n12762) );
  AND U13354 ( .A(n8839), .B(n8885), .Z(n13683) );
  XOR U13355 ( .A(n13685), .B(n11769), .Z(n8885) );
  XNOR U13356 ( .A(n12880), .B(n13686), .Z(n8839) );
  XNOR U13357 ( .A(n13687), .B(n13688), .Z(n12880) );
  XOR U13358 ( .A(n13689), .B(n6483), .Z(n5464) );
  XOR U13359 ( .A(n11409), .B(n13052), .Z(n6483) );
  XOR U13360 ( .A(n13690), .B(n13691), .Z(n13052) );
  AND U13361 ( .A(n13692), .B(n13693), .Z(n13690) );
  XOR U13362 ( .A(n13694), .B(n13695), .Z(n11409) );
  ANDN U13363 ( .B(n8882), .A(n13272), .Z(n13689) );
  XOR U13364 ( .A(n3469), .B(n13696), .Z(n13681) );
  XOR U13365 ( .A(n8874), .B(n4851), .Z(n13696) );
  XNOR U13366 ( .A(n13697), .B(n6478), .Z(n4851) );
  XOR U13367 ( .A(n9177), .B(n13698), .Z(n6478) );
  ANDN U13368 ( .B(n8836), .A(n8835), .Z(n13697) );
  XOR U13369 ( .A(n11257), .B(n13699), .Z(n8835) );
  XOR U13370 ( .A(n13700), .B(n10265), .Z(n8836) );
  XNOR U13371 ( .A(n13368), .B(n11853), .Z(n10265) );
  XNOR U13372 ( .A(n13701), .B(n13702), .Z(n11853) );
  XOR U13373 ( .A(n10591), .B(n10435), .Z(n13702) );
  XNOR U13374 ( .A(n13703), .B(n13704), .Z(n10435) );
  ANDN U13375 ( .B(n13705), .A(n13706), .Z(n13703) );
  XNOR U13376 ( .A(n13707), .B(n13708), .Z(n10591) );
  ANDN U13377 ( .B(n13709), .A(n13710), .Z(n13707) );
  XNOR U13378 ( .A(n9677), .B(n13711), .Z(n13701) );
  XOR U13379 ( .A(n13712), .B(n10368), .Z(n13711) );
  XNOR U13380 ( .A(n13713), .B(n13714), .Z(n10368) );
  AND U13381 ( .A(n13715), .B(n13716), .Z(n13713) );
  XNOR U13382 ( .A(n13717), .B(n13718), .Z(n9677) );
  ANDN U13383 ( .B(n13719), .A(n13720), .Z(n13717) );
  XOR U13384 ( .A(n13721), .B(n13722), .Z(n13368) );
  XNOR U13385 ( .A(n10885), .B(n9791), .Z(n13722) );
  XOR U13386 ( .A(n13723), .B(n13724), .Z(n9791) );
  AND U13387 ( .A(n13725), .B(n13726), .Z(n13723) );
  XNOR U13388 ( .A(n13727), .B(n13728), .Z(n10885) );
  AND U13389 ( .A(n13729), .B(n13730), .Z(n13727) );
  XNOR U13390 ( .A(n13380), .B(n13731), .Z(n13721) );
  XOR U13391 ( .A(n12663), .B(n9076), .Z(n13731) );
  XNOR U13392 ( .A(n13732), .B(n13733), .Z(n9076) );
  ANDN U13393 ( .B(n13734), .A(n13735), .Z(n13732) );
  XNOR U13394 ( .A(n13736), .B(n13737), .Z(n12663) );
  ANDN U13395 ( .B(n13738), .A(n13739), .Z(n13736) );
  XNOR U13396 ( .A(n13740), .B(n13741), .Z(n13380) );
  AND U13397 ( .A(n13742), .B(n13743), .Z(n13740) );
  XNOR U13398 ( .A(n13744), .B(n6474), .Z(n8874) );
  XNOR U13399 ( .A(n13745), .B(n9922), .Z(n6474) );
  XNOR U13400 ( .A(n12583), .B(n13746), .Z(n9922) );
  XOR U13401 ( .A(n13747), .B(n13748), .Z(n12583) );
  XNOR U13402 ( .A(n11028), .B(n10660), .Z(n13748) );
  XOR U13403 ( .A(n13749), .B(n13750), .Z(n10660) );
  ANDN U13404 ( .B(n13751), .A(n13752), .Z(n13749) );
  XNOR U13405 ( .A(n13753), .B(n13754), .Z(n11028) );
  AND U13406 ( .A(n13755), .B(n13756), .Z(n13753) );
  XOR U13407 ( .A(n13225), .B(n13757), .Z(n13747) );
  XOR U13408 ( .A(n10091), .B(n9180), .Z(n13757) );
  XNOR U13409 ( .A(n13758), .B(n13242), .Z(n9180) );
  ANDN U13410 ( .B(n13243), .A(n13759), .Z(n13758) );
  XNOR U13411 ( .A(n13760), .B(n13761), .Z(n10091) );
  XNOR U13412 ( .A(n13764), .B(n13232), .Z(n13225) );
  AND U13413 ( .A(n8830), .B(n8829), .Z(n13744) );
  IV U13414 ( .A(n8878), .Z(n8829) );
  XOR U13415 ( .A(n13766), .B(n9270), .Z(n8878) );
  IV U13416 ( .A(n10200), .Z(n9270) );
  XNOR U13417 ( .A(n13188), .B(n11659), .Z(n10200) );
  XNOR U13418 ( .A(n13767), .B(n13768), .Z(n11659) );
  XOR U13419 ( .A(n13590), .B(n10045), .Z(n13768) );
  XNOR U13420 ( .A(n13769), .B(n13770), .Z(n10045) );
  AND U13421 ( .A(n13771), .B(n13772), .Z(n13769) );
  XOR U13422 ( .A(n13773), .B(n13774), .Z(n13590) );
  ANDN U13423 ( .B(n13775), .A(n13776), .Z(n13773) );
  XOR U13424 ( .A(n13777), .B(n13778), .Z(n13767) );
  XNOR U13425 ( .A(n11063), .B(n11920), .Z(n13778) );
  XNOR U13426 ( .A(n13779), .B(n13780), .Z(n11920) );
  ANDN U13427 ( .B(n13781), .A(n13782), .Z(n13779) );
  XNOR U13428 ( .A(n13783), .B(n13784), .Z(n11063) );
  AND U13429 ( .A(n13785), .B(n13786), .Z(n13783) );
  XOR U13430 ( .A(n13787), .B(n13788), .Z(n13188) );
  XOR U13431 ( .A(n13048), .B(n10680), .Z(n13788) );
  XOR U13432 ( .A(n13789), .B(n13790), .Z(n10680) );
  ANDN U13433 ( .B(n13791), .A(n13792), .Z(n13789) );
  XNOR U13434 ( .A(n13793), .B(n13794), .Z(n13048) );
  ANDN U13435 ( .B(n13795), .A(n13796), .Z(n13793) );
  XOR U13436 ( .A(n12652), .B(n13797), .Z(n13787) );
  XNOR U13437 ( .A(n12630), .B(n11817), .Z(n13797) );
  XNOR U13438 ( .A(n13798), .B(n13799), .Z(n11817) );
  ANDN U13439 ( .B(n13800), .A(n13801), .Z(n13798) );
  XNOR U13440 ( .A(n13802), .B(n13803), .Z(n12630) );
  AND U13441 ( .A(n13804), .B(n13805), .Z(n13802) );
  XNOR U13442 ( .A(n13806), .B(n13807), .Z(n12652) );
  AND U13443 ( .A(n13808), .B(n13809), .Z(n13806) );
  XNOR U13444 ( .A(n13810), .B(n13811), .Z(n8830) );
  XNOR U13445 ( .A(n13812), .B(n6487), .Z(n3469) );
  XNOR U13446 ( .A(n9588), .B(n13813), .Z(n6487) );
  XOR U13447 ( .A(n13814), .B(n12976), .Z(n9588) );
  XOR U13448 ( .A(n13815), .B(n13816), .Z(n12976) );
  XNOR U13449 ( .A(n13039), .B(n13817), .Z(n13816) );
  XNOR U13450 ( .A(n13818), .B(n13819), .Z(n13039) );
  AND U13451 ( .A(n13820), .B(n13821), .Z(n13818) );
  XNOR U13452 ( .A(n9277), .B(n13822), .Z(n13815) );
  XOR U13453 ( .A(n12560), .B(n10062), .Z(n13822) );
  XNOR U13454 ( .A(n13823), .B(n13824), .Z(n10062) );
  ANDN U13455 ( .B(n13825), .A(n13826), .Z(n13823) );
  XNOR U13456 ( .A(n13827), .B(n13828), .Z(n12560) );
  AND U13457 ( .A(n13829), .B(n13830), .Z(n13827) );
  XNOR U13458 ( .A(n13831), .B(n13832), .Z(n9277) );
  AND U13459 ( .A(n13833), .B(n13834), .Z(n13831) );
  NOR U13460 ( .A(n8827), .B(n8826), .Z(n13812) );
  XOR U13461 ( .A(n9682), .B(n13835), .Z(n8826) );
  XOR U13462 ( .A(n13836), .B(n12548), .Z(n9682) );
  XNOR U13463 ( .A(n13837), .B(n13838), .Z(n12548) );
  XOR U13464 ( .A(n13839), .B(n10049), .Z(n13838) );
  XOR U13465 ( .A(n13840), .B(n13841), .Z(n10049) );
  AND U13466 ( .A(n13842), .B(n13843), .Z(n13840) );
  XOR U13467 ( .A(n13844), .B(n13845), .Z(n13837) );
  XOR U13468 ( .A(n13846), .B(n13847), .Z(n13845) );
  XNOR U13469 ( .A(n13848), .B(n12074), .Z(n8827) );
  XNOR U13470 ( .A(n13849), .B(n13850), .Z(n6287) );
  XOR U13471 ( .A(n5427), .B(n3673), .Z(n13850) );
  XNOR U13472 ( .A(n13851), .B(n13852), .Z(n3673) );
  ANDN U13473 ( .B(n6507), .A(n6508), .Z(n13851) );
  XNOR U13474 ( .A(n13853), .B(n11769), .Z(n6508) );
  IV U13475 ( .A(n10997), .Z(n11769) );
  XNOR U13476 ( .A(n13854), .B(n8894), .Z(n5427) );
  ANDN U13477 ( .B(n8895), .A(n6499), .Z(n13854) );
  XNOR U13478 ( .A(n13855), .B(n12074), .Z(n6499) );
  IV U13479 ( .A(n13856), .Z(n12074) );
  XNOR U13480 ( .A(n13857), .B(n11656), .Z(n8895) );
  XNOR U13481 ( .A(n4287), .B(n13858), .Z(n13849) );
  XOR U13482 ( .A(n5865), .B(n2119), .Z(n13858) );
  XNOR U13483 ( .A(n13859), .B(n8890), .Z(n2119) );
  ANDN U13484 ( .B(n8891), .A(n6512), .Z(n13859) );
  XOR U13485 ( .A(n10227), .B(n13860), .Z(n6512) );
  IV U13486 ( .A(n13861), .Z(n10227) );
  XNOR U13487 ( .A(n13862), .B(n9551), .Z(n8891) );
  XNOR U13488 ( .A(n13863), .B(n12092), .Z(n9551) );
  XNOR U13489 ( .A(n13864), .B(n13865), .Z(n12092) );
  XNOR U13490 ( .A(n13866), .B(n12215), .Z(n13865) );
  XOR U13491 ( .A(n13867), .B(n13868), .Z(n12215) );
  NOR U13492 ( .A(n13342), .B(n13341), .Z(n13867) );
  XOR U13493 ( .A(n11873), .B(n13869), .Z(n13864) );
  XOR U13494 ( .A(n9802), .B(n12453), .Z(n13869) );
  XNOR U13495 ( .A(n13870), .B(n13871), .Z(n12453) );
  ANDN U13496 ( .B(n13346), .A(n13347), .Z(n13870) );
  XNOR U13497 ( .A(n13872), .B(n13873), .Z(n9802) );
  XNOR U13498 ( .A(n13874), .B(n13875), .Z(n11873) );
  ANDN U13499 ( .B(n13354), .A(n13355), .Z(n13874) );
  XOR U13500 ( .A(n13876), .B(n8903), .Z(n5865) );
  NOR U13501 ( .A(n6516), .B(n6515), .Z(n13876) );
  XNOR U13502 ( .A(n9168), .B(n13877), .Z(n6515) );
  XNOR U13503 ( .A(n13879), .B(n13880), .Z(n11930) );
  XOR U13504 ( .A(n11938), .B(n12827), .Z(n13880) );
  XOR U13505 ( .A(n13881), .B(n13351), .Z(n12827) );
  XNOR U13506 ( .A(n13882), .B(n13883), .Z(n13351) );
  ANDN U13507 ( .B(n13352), .A(n13884), .Z(n13881) );
  XNOR U13508 ( .A(n13885), .B(n13355), .Z(n11938) );
  XNOR U13509 ( .A(n13886), .B(n13887), .Z(n13355) );
  ANDN U13510 ( .B(n13888), .A(n13356), .Z(n13885) );
  XOR U13511 ( .A(n11300), .B(n13889), .Z(n13879) );
  XOR U13512 ( .A(n10135), .B(n12616), .Z(n13889) );
  XNOR U13513 ( .A(n13890), .B(n13342), .Z(n12616) );
  XNOR U13514 ( .A(n13891), .B(n13892), .Z(n13342) );
  NOR U13515 ( .A(n13343), .B(n13893), .Z(n13890) );
  XNOR U13516 ( .A(n13894), .B(n13347), .Z(n10135) );
  XOR U13517 ( .A(n13895), .B(n13896), .Z(n13347) );
  AND U13518 ( .A(n13348), .B(n13897), .Z(n13894) );
  XNOR U13519 ( .A(n13898), .B(n13338), .Z(n11300) );
  NOR U13520 ( .A(n13899), .B(n13339), .Z(n13898) );
  XNOR U13521 ( .A(n9393), .B(n13900), .Z(n6516) );
  XOR U13522 ( .A(n13901), .B(n8900), .Z(n4287) );
  ANDN U13523 ( .B(n6502), .A(n6503), .Z(n13901) );
  XOR U13524 ( .A(n13902), .B(n9595), .Z(n6503) );
  IV U13525 ( .A(n9713), .Z(n9595) );
  XOR U13526 ( .A(n13903), .B(n13811), .Z(n6502) );
  IV U13527 ( .A(n11065), .Z(n13811) );
  XNOR U13528 ( .A(n13904), .B(n13905), .Z(n11065) );
  XNOR U13529 ( .A(n13906), .B(n8882), .Z(n8833) );
  ANDN U13530 ( .B(n13272), .A(n6481), .Z(n13906) );
  XOR U13531 ( .A(n13908), .B(n11404), .Z(n6481) );
  XOR U13532 ( .A(n13909), .B(n13910), .Z(n11404) );
  XNOR U13533 ( .A(n13911), .B(n9372), .Z(n13272) );
  IV U13534 ( .A(n13912), .Z(n9372) );
  XOR U13535 ( .A(n11486), .B(n2085), .Z(n5654) );
  XNOR U13536 ( .A(n8266), .B(n9650), .Z(n2085) );
  XNOR U13537 ( .A(n13913), .B(n13914), .Z(n9650) );
  XOR U13538 ( .A(n5456), .B(n3587), .Z(n13914) );
  XNOR U13539 ( .A(n13915), .B(n13916), .Z(n3587) );
  AND U13540 ( .A(n8364), .B(n8363), .Z(n13915) );
  IV U13541 ( .A(n13917), .Z(n8363) );
  XOR U13542 ( .A(n10900), .B(n13918), .Z(n8364) );
  IV U13543 ( .A(n10838), .Z(n10900) );
  XOR U13544 ( .A(n13687), .B(n13919), .Z(n10838) );
  XOR U13545 ( .A(n13920), .B(n13921), .Z(n13687) );
  XNOR U13546 ( .A(n12130), .B(n12240), .Z(n13921) );
  XNOR U13547 ( .A(n13922), .B(n13093), .Z(n12240) );
  ANDN U13548 ( .B(n13094), .A(n13923), .Z(n13922) );
  XOR U13549 ( .A(n13924), .B(n13925), .Z(n12130) );
  XOR U13550 ( .A(n10581), .B(n13928), .Z(n13920) );
  XOR U13551 ( .A(n10454), .B(n12262), .Z(n13928) );
  XNOR U13552 ( .A(n13929), .B(n13102), .Z(n12262) );
  ANDN U13553 ( .B(n13103), .A(n13930), .Z(n13929) );
  XNOR U13554 ( .A(n13931), .B(n13098), .Z(n10454) );
  AND U13555 ( .A(n13099), .B(n13932), .Z(n13931) );
  XNOR U13556 ( .A(n13933), .B(n13106), .Z(n10581) );
  ANDN U13557 ( .B(n13107), .A(n13934), .Z(n13933) );
  XNOR U13558 ( .A(n13935), .B(n11618), .Z(n5456) );
  AND U13559 ( .A(n8361), .B(n8359), .Z(n13935) );
  XNOR U13560 ( .A(n10562), .B(n13662), .Z(n8361) );
  XOR U13561 ( .A(n13937), .B(n13938), .Z(n13662) );
  NOR U13562 ( .A(n13939), .B(n13940), .Z(n13937) );
  IV U13563 ( .A(n10379), .Z(n10562) );
  XOR U13564 ( .A(n13941), .B(n12862), .Z(n10379) );
  XOR U13565 ( .A(n13942), .B(n13943), .Z(n12862) );
  XNOR U13566 ( .A(n13944), .B(n9601), .Z(n13943) );
  XOR U13567 ( .A(n13945), .B(n13946), .Z(n9601) );
  ANDN U13568 ( .B(n13947), .A(n13948), .Z(n13945) );
  XOR U13569 ( .A(n11783), .B(n13949), .Z(n13942) );
  XOR U13570 ( .A(n10460), .B(n11246), .Z(n13949) );
  XNOR U13571 ( .A(n13950), .B(n13951), .Z(n11246) );
  XOR U13572 ( .A(n13954), .B(n13955), .Z(n10460) );
  AND U13573 ( .A(n13956), .B(n13957), .Z(n13954) );
  XNOR U13574 ( .A(n13958), .B(n13959), .Z(n11783) );
  AND U13575 ( .A(n13960), .B(n13961), .Z(n13958) );
  XOR U13576 ( .A(n6245), .B(n13962), .Z(n13913) );
  XOR U13577 ( .A(n2378), .B(n5599), .Z(n13962) );
  XNOR U13578 ( .A(n13963), .B(n11629), .Z(n5599) );
  AND U13579 ( .A(n9654), .B(n11630), .Z(n13963) );
  XOR U13580 ( .A(n13866), .B(n9803), .Z(n11630) );
  XNOR U13581 ( .A(n13964), .B(n13112), .Z(n9803) );
  XNOR U13582 ( .A(n13965), .B(n13966), .Z(n13112) );
  XNOR U13583 ( .A(n12202), .B(n11939), .Z(n13966) );
  XNOR U13584 ( .A(n13967), .B(n13968), .Z(n11939) );
  ANDN U13585 ( .B(n13969), .A(n13970), .Z(n13967) );
  XNOR U13586 ( .A(n13971), .B(n13972), .Z(n12202) );
  AND U13587 ( .A(n13973), .B(n13974), .Z(n13971) );
  XOR U13588 ( .A(n12000), .B(n13975), .Z(n13965) );
  XOR U13589 ( .A(n11714), .B(n12222), .Z(n13975) );
  XOR U13590 ( .A(n13976), .B(n13977), .Z(n12222) );
  ANDN U13591 ( .B(n13978), .A(n13979), .Z(n13976) );
  XOR U13592 ( .A(n13980), .B(n13981), .Z(n11714) );
  XNOR U13593 ( .A(n13984), .B(n13985), .Z(n12000) );
  ANDN U13594 ( .B(n13986), .A(n13987), .Z(n13984) );
  XNOR U13595 ( .A(n13988), .B(n13989), .Z(n13866) );
  ANDN U13596 ( .B(n13337), .A(n13338), .Z(n13988) );
  XNOR U13597 ( .A(n13990), .B(n13991), .Z(n13338) );
  XNOR U13598 ( .A(n13992), .B(n11192), .Z(n9654) );
  XNOR U13599 ( .A(n13993), .B(n11621), .Z(n2378) );
  ANDN U13600 ( .B(n8350), .A(n8349), .Z(n13993) );
  XOR U13601 ( .A(n11301), .B(n13616), .Z(n8349) );
  XNOR U13602 ( .A(n13994), .B(n13995), .Z(n13616) );
  AND U13603 ( .A(n13996), .B(n13997), .Z(n13994) );
  XNOR U13604 ( .A(n13998), .B(n10603), .Z(n8350) );
  XNOR U13605 ( .A(n13999), .B(n11626), .Z(n6245) );
  ANDN U13606 ( .B(n8355), .A(n8353), .Z(n13999) );
  XNOR U13607 ( .A(n14000), .B(n11656), .Z(n8353) );
  XNOR U13608 ( .A(n14001), .B(n12671), .Z(n8355) );
  XOR U13609 ( .A(n14002), .B(n14003), .Z(n12671) );
  XOR U13610 ( .A(n14004), .B(n14005), .Z(n8266) );
  XNOR U13611 ( .A(n3800), .B(n5117), .Z(n14005) );
  XOR U13612 ( .A(n14006), .B(n9545), .Z(n5117) );
  XOR U13613 ( .A(n14007), .B(n9713), .Z(n9545) );
  XOR U13614 ( .A(n14008), .B(n14009), .Z(n9713) );
  XOR U13615 ( .A(n14010), .B(n9917), .Z(n11493) );
  XOR U13616 ( .A(n11301), .B(n13612), .Z(n11492) );
  XNOR U13617 ( .A(n14011), .B(n14012), .Z(n13612) );
  ANDN U13618 ( .B(n14013), .A(n13141), .Z(n14011) );
  IV U13619 ( .A(n10827), .Z(n11301) );
  XNOR U13620 ( .A(n12598), .B(n14014), .Z(n10827) );
  XOR U13621 ( .A(n14015), .B(n14016), .Z(n12598) );
  XOR U13622 ( .A(n14017), .B(n11038), .Z(n14016) );
  XOR U13623 ( .A(n14018), .B(n14019), .Z(n11038) );
  AND U13624 ( .A(n13631), .B(n13633), .Z(n14018) );
  XOR U13625 ( .A(n12338), .B(n14020), .Z(n14015) );
  XOR U13626 ( .A(n11815), .B(n9819), .Z(n14020) );
  XNOR U13627 ( .A(n14021), .B(n14022), .Z(n9819) );
  AND U13628 ( .A(n13646), .B(n14023), .Z(n14021) );
  XNOR U13629 ( .A(n14024), .B(n14025), .Z(n11815) );
  AND U13630 ( .A(n13640), .B(n14026), .Z(n14024) );
  XNOR U13631 ( .A(n14027), .B(n14028), .Z(n12338) );
  XOR U13632 ( .A(n14029), .B(n8324), .Z(n3800) );
  XOR U13633 ( .A(n10149), .B(n14030), .Z(n8324) );
  IV U13634 ( .A(n13115), .Z(n10149) );
  XOR U13635 ( .A(n14032), .B(n14033), .Z(n10673) );
  XOR U13636 ( .A(n14034), .B(n11576), .Z(n14033) );
  XOR U13637 ( .A(n14035), .B(n14036), .Z(n11576) );
  XOR U13638 ( .A(n10016), .B(n14039), .Z(n14032) );
  XOR U13639 ( .A(n11726), .B(n14040), .Z(n14039) );
  XNOR U13640 ( .A(n14041), .B(n14042), .Z(n11726) );
  NOR U13641 ( .A(n14043), .B(n14044), .Z(n14041) );
  XOR U13642 ( .A(n14045), .B(n14046), .Z(n10016) );
  NOR U13643 ( .A(n14047), .B(n14048), .Z(n14045) );
  ANDN U13644 ( .B(n11484), .A(n11485), .Z(n14029) );
  XNOR U13645 ( .A(n13540), .B(n9900), .Z(n11485) );
  XOR U13646 ( .A(n14049), .B(n13483), .Z(n13540) );
  ANDN U13647 ( .B(n14050), .A(n14051), .Z(n14049) );
  XNOR U13648 ( .A(n14052), .B(n10126), .Z(n11484) );
  XNOR U13649 ( .A(n5080), .B(n14053), .Z(n14004) );
  XOR U13650 ( .A(n1737), .B(n11604), .Z(n14053) );
  XOR U13651 ( .A(n14054), .B(n8333), .Z(n11604) );
  XOR U13652 ( .A(n14055), .B(n10938), .Z(n8333) );
  XNOR U13653 ( .A(n12547), .B(n14056), .Z(n10938) );
  XOR U13654 ( .A(n14057), .B(n14058), .Z(n12547) );
  XOR U13655 ( .A(n14059), .B(n9371), .Z(n14058) );
  XOR U13656 ( .A(n14060), .B(n14061), .Z(n9371) );
  AND U13657 ( .A(n14062), .B(n14063), .Z(n14060) );
  XOR U13658 ( .A(n13911), .B(n14064), .Z(n14057) );
  XOR U13659 ( .A(n10428), .B(n12310), .Z(n14064) );
  XOR U13660 ( .A(n14065), .B(n14066), .Z(n12310) );
  XOR U13661 ( .A(n14069), .B(n14070), .Z(n10428) );
  NOR U13662 ( .A(n14071), .B(n14072), .Z(n14069) );
  XNOR U13663 ( .A(n14073), .B(n14074), .Z(n13911) );
  AND U13664 ( .A(n14075), .B(n14076), .Z(n14073) );
  NOR U13665 ( .A(n11481), .B(n11482), .Z(n14054) );
  XNOR U13666 ( .A(n11712), .B(n14077), .Z(n11482) );
  XOR U13667 ( .A(n14078), .B(n14079), .Z(n11712) );
  XNOR U13668 ( .A(n14080), .B(n10991), .Z(n11481) );
  XNOR U13669 ( .A(n12942), .B(n14081), .Z(n10991) );
  XOR U13670 ( .A(n14082), .B(n14083), .Z(n12942) );
  XOR U13671 ( .A(n10042), .B(n11988), .Z(n14083) );
  XNOR U13672 ( .A(n14084), .B(n14085), .Z(n11988) );
  AND U13673 ( .A(n13413), .B(n14086), .Z(n14084) );
  IV U13674 ( .A(n14087), .Z(n13413) );
  XOR U13675 ( .A(n14088), .B(n14089), .Z(n10042) );
  AND U13676 ( .A(n13409), .B(n14090), .Z(n14088) );
  XNOR U13677 ( .A(n10283), .B(n14091), .Z(n14082) );
  XNOR U13678 ( .A(n11775), .B(n10926), .Z(n14091) );
  XNOR U13679 ( .A(n14092), .B(n14093), .Z(n10926) );
  AND U13680 ( .A(n14094), .B(n14095), .Z(n14092) );
  XNOR U13681 ( .A(n14096), .B(n14097), .Z(n11775) );
  AND U13682 ( .A(n14098), .B(n13405), .Z(n14096) );
  XNOR U13683 ( .A(n14099), .B(n14100), .Z(n10283) );
  AND U13684 ( .A(n14101), .B(n14102), .Z(n14099) );
  XOR U13685 ( .A(n14103), .B(n8327), .Z(n1737) );
  XNOR U13686 ( .A(n14104), .B(n10245), .Z(n8327) );
  IV U13687 ( .A(n11747), .Z(n10245) );
  XNOR U13688 ( .A(n13288), .B(n14105), .Z(n11747) );
  XOR U13689 ( .A(n14106), .B(n14107), .Z(n13288) );
  XNOR U13690 ( .A(n12848), .B(n11543), .Z(n14107) );
  XOR U13691 ( .A(n14108), .B(n14109), .Z(n11543) );
  AND U13692 ( .A(n12902), .B(n14110), .Z(n14108) );
  XOR U13693 ( .A(n14111), .B(n14112), .Z(n12848) );
  ANDN U13694 ( .B(n14113), .A(n12898), .Z(n14111) );
  XOR U13695 ( .A(n12348), .B(n14114), .Z(n14106) );
  XOR U13696 ( .A(n11463), .B(n14115), .Z(n14114) );
  XNOR U13697 ( .A(n14116), .B(n14117), .Z(n11463) );
  AND U13698 ( .A(n12906), .B(n14118), .Z(n14116) );
  XNOR U13699 ( .A(n14119), .B(n14120), .Z(n12348) );
  ANDN U13700 ( .B(n14121), .A(n14122), .Z(n14119) );
  NOR U13701 ( .A(n11490), .B(n11489), .Z(n14103) );
  XNOR U13702 ( .A(n10208), .B(n14123), .Z(n11489) );
  IV U13703 ( .A(n9485), .Z(n10208) );
  XOR U13704 ( .A(n14124), .B(n14125), .Z(n9485) );
  XOR U13705 ( .A(n14126), .B(n10022), .Z(n11490) );
  XNOR U13706 ( .A(n14127), .B(n8338), .Z(n5080) );
  XOR U13707 ( .A(n14128), .B(n12050), .Z(n8338) );
  AND U13708 ( .A(n11611), .B(n13319), .Z(n14127) );
  IV U13709 ( .A(n14129), .Z(n13319) );
  XOR U13710 ( .A(n14130), .B(n11611), .Z(n11486) );
  XNOR U13711 ( .A(n13026), .B(n9776), .Z(n11611) );
  IV U13712 ( .A(n10371), .Z(n9776) );
  XNOR U13713 ( .A(n14131), .B(n14132), .Z(n10371) );
  XNOR U13714 ( .A(n14133), .B(n14134), .Z(n13026) );
  ANDN U13715 ( .B(n13504), .A(n13502), .Z(n14133) );
  ANDN U13716 ( .B(n14129), .A(n8336), .Z(n14130) );
  XOR U13717 ( .A(n10104), .B(n14135), .Z(n8336) );
  XOR U13718 ( .A(n14136), .B(n13511), .Z(n10104) );
  XNOR U13719 ( .A(n14137), .B(n14138), .Z(n13511) );
  XNOR U13720 ( .A(n14139), .B(n10646), .Z(n14138) );
  XOR U13721 ( .A(n14140), .B(n14141), .Z(n10646) );
  ANDN U13722 ( .B(n14142), .A(n14143), .Z(n14140) );
  XOR U13723 ( .A(n9767), .B(n14144), .Z(n14137) );
  XNOR U13724 ( .A(n12229), .B(n14145), .Z(n14144) );
  XOR U13725 ( .A(n14146), .B(n14147), .Z(n12229) );
  ANDN U13726 ( .B(n14148), .A(n14149), .Z(n14146) );
  XNOR U13727 ( .A(n14150), .B(n14151), .Z(n9767) );
  ANDN U13728 ( .B(n14152), .A(n14153), .Z(n14150) );
  XNOR U13729 ( .A(n14154), .B(n12069), .Z(n14129) );
  XNOR U13730 ( .A(n14155), .B(n6173), .Z(out[1001]) );
  XNOR U13731 ( .A(n9038), .B(n2296), .Z(n6173) );
  XNOR U13732 ( .A(n9983), .B(n6133), .Z(n2296) );
  XNOR U13733 ( .A(n14156), .B(n14157), .Z(n6133) );
  XNOR U13734 ( .A(n2334), .B(n5443), .Z(n14157) );
  XOR U13735 ( .A(n14158), .B(n7951), .Z(n5443) );
  XNOR U13736 ( .A(n14159), .B(n10307), .Z(n7951) );
  XOR U13737 ( .A(n12985), .B(n14131), .Z(n10307) );
  XOR U13738 ( .A(n14160), .B(n14161), .Z(n14131) );
  XNOR U13739 ( .A(n12868), .B(n13514), .Z(n14161) );
  XNOR U13740 ( .A(n14162), .B(n13544), .Z(n13514) );
  ANDN U13741 ( .B(n14163), .A(n13543), .Z(n14162) );
  XNOR U13742 ( .A(n14164), .B(n14165), .Z(n12868) );
  NOR U13743 ( .A(n14166), .B(n14167), .Z(n14164) );
  XNOR U13744 ( .A(n12878), .B(n14168), .Z(n14160) );
  XNOR U13745 ( .A(n12357), .B(n11589), .Z(n14168) );
  XOR U13746 ( .A(n14169), .B(n14050), .Z(n11589) );
  AND U13747 ( .A(n13482), .B(n14051), .Z(n14169) );
  XOR U13748 ( .A(n14170), .B(n13538), .Z(n12357) );
  ANDN U13749 ( .B(n13489), .A(n13537), .Z(n14170) );
  XOR U13750 ( .A(n14171), .B(n13546), .Z(n12878) );
  ANDN U13751 ( .B(n14172), .A(n13478), .Z(n14171) );
  XOR U13752 ( .A(n14173), .B(n14174), .Z(n12985) );
  XNOR U13753 ( .A(n13416), .B(n11739), .Z(n14174) );
  XOR U13754 ( .A(n14175), .B(n14176), .Z(n11739) );
  ANDN U13755 ( .B(n14177), .A(n14178), .Z(n14175) );
  XNOR U13756 ( .A(n14179), .B(n13519), .Z(n13416) );
  ANDN U13757 ( .B(n13520), .A(n14180), .Z(n14179) );
  XOR U13758 ( .A(n12273), .B(n14181), .Z(n14173) );
  XOR U13759 ( .A(n10236), .B(n10173), .Z(n14181) );
  XNOR U13760 ( .A(n14182), .B(n13523), .Z(n10173) );
  AND U13761 ( .A(n14183), .B(n14184), .Z(n14182) );
  XNOR U13762 ( .A(n14185), .B(n13530), .Z(n10236) );
  ANDN U13763 ( .B(n13531), .A(n14186), .Z(n14185) );
  XNOR U13764 ( .A(n14187), .B(n14188), .Z(n12273) );
  AND U13765 ( .A(n7950), .B(n9048), .Z(n14158) );
  XOR U13766 ( .A(n13847), .B(n10050), .Z(n9048) );
  XOR U13767 ( .A(n14191), .B(n14192), .Z(n13847) );
  ANDN U13768 ( .B(n14193), .A(n14194), .Z(n14191) );
  XNOR U13769 ( .A(n13861), .B(n14195), .Z(n7950) );
  XOR U13770 ( .A(n11131), .B(n14196), .Z(n13861) );
  XOR U13771 ( .A(n14197), .B(n14198), .Z(n11131) );
  XOR U13772 ( .A(n9691), .B(n10572), .Z(n14198) );
  XOR U13773 ( .A(n14199), .B(n13953), .Z(n10572) );
  NOR U13774 ( .A(n13952), .B(n14200), .Z(n14199) );
  XNOR U13775 ( .A(n14201), .B(n13948), .Z(n9691) );
  ANDN U13776 ( .B(n14202), .A(n14203), .Z(n14201) );
  XNOR U13777 ( .A(n12861), .B(n14204), .Z(n14197) );
  XNOR U13778 ( .A(n12356), .B(n11160), .Z(n14204) );
  XOR U13779 ( .A(n14205), .B(n14206), .Z(n11160) );
  NOR U13780 ( .A(n14207), .B(n13960), .Z(n14205) );
  XNOR U13781 ( .A(n14208), .B(n14209), .Z(n12356) );
  NOR U13782 ( .A(n13956), .B(n14210), .Z(n14208) );
  XNOR U13783 ( .A(n14211), .B(n14212), .Z(n12861) );
  ANDN U13784 ( .B(n14213), .A(n14214), .Z(n14211) );
  XNOR U13785 ( .A(n14215), .B(n7954), .Z(n2334) );
  XNOR U13786 ( .A(n14216), .B(n9950), .Z(n7954) );
  IV U13787 ( .A(n9183), .Z(n9950) );
  ANDN U13788 ( .B(n9043), .A(n9044), .Z(n14215) );
  XNOR U13789 ( .A(n14217), .B(n11916), .Z(n9044) );
  XNOR U13790 ( .A(n14079), .B(n12720), .Z(n11916) );
  XNOR U13791 ( .A(n14218), .B(n14219), .Z(n12720) );
  XNOR U13792 ( .A(n14220), .B(n14221), .Z(n14219) );
  XOR U13793 ( .A(n14222), .B(n14223), .Z(n14218) );
  XNOR U13794 ( .A(n11860), .B(n11650), .Z(n14223) );
  XNOR U13795 ( .A(n14224), .B(n14178), .Z(n11650) );
  ANDN U13796 ( .B(n14225), .A(n14226), .Z(n14224) );
  XNOR U13797 ( .A(n14227), .B(n14183), .Z(n11860) );
  AND U13798 ( .A(n13522), .B(n14228), .Z(n14227) );
  XOR U13799 ( .A(n14229), .B(n14230), .Z(n14079) );
  XOR U13800 ( .A(n10895), .B(n12204), .Z(n14230) );
  XOR U13801 ( .A(n14231), .B(n14232), .Z(n12204) );
  ANDN U13802 ( .B(n14233), .A(n14234), .Z(n14231) );
  XOR U13803 ( .A(n14235), .B(n14236), .Z(n10895) );
  ANDN U13804 ( .B(n14237), .A(n14238), .Z(n14235) );
  XNOR U13805 ( .A(n10112), .B(n14239), .Z(n14229) );
  XNOR U13806 ( .A(n11673), .B(n14240), .Z(n14239) );
  XNOR U13807 ( .A(n14241), .B(n14242), .Z(n11673) );
  AND U13808 ( .A(n14243), .B(n14244), .Z(n14241) );
  XNOR U13809 ( .A(n14245), .B(n14246), .Z(n10112) );
  NOR U13810 ( .A(n14247), .B(n14248), .Z(n14245) );
  XOR U13811 ( .A(n9494), .B(n14249), .Z(n9043) );
  XOR U13812 ( .A(n14250), .B(n14251), .Z(n9494) );
  XOR U13813 ( .A(n3157), .B(n14252), .Z(n14156) );
  XOR U13814 ( .A(n6260), .B(n7944), .Z(n14252) );
  XOR U13815 ( .A(n14253), .B(n7960), .Z(n7944) );
  XNOR U13816 ( .A(n13402), .B(n9119), .Z(n7960) );
  XNOR U13817 ( .A(n14254), .B(n14101), .Z(n13402) );
  AND U13818 ( .A(n14255), .B(n14256), .Z(n14254) );
  AND U13819 ( .A(n9046), .B(n7959), .Z(n14253) );
  XNOR U13820 ( .A(n14257), .B(n10920), .Z(n7959) );
  XOR U13821 ( .A(n14258), .B(n12701), .Z(n10920) );
  XOR U13822 ( .A(n14259), .B(n14260), .Z(n12701) );
  XNOR U13823 ( .A(n14261), .B(n11682), .Z(n14260) );
  XOR U13824 ( .A(n14262), .B(n14263), .Z(n11682) );
  XNOR U13825 ( .A(n10430), .B(n14266), .Z(n14259) );
  XOR U13826 ( .A(n12585), .B(n11528), .Z(n14266) );
  XNOR U13827 ( .A(n14267), .B(n14268), .Z(n11528) );
  AND U13828 ( .A(n14269), .B(n14270), .Z(n14267) );
  XNOR U13829 ( .A(n14271), .B(n14272), .Z(n12585) );
  ANDN U13830 ( .B(n14273), .A(n14274), .Z(n14271) );
  XOR U13831 ( .A(n14275), .B(n14276), .Z(n10430) );
  ANDN U13832 ( .B(n14277), .A(n14278), .Z(n14275) );
  XNOR U13833 ( .A(n14279), .B(n12473), .Z(n9046) );
  XOR U13834 ( .A(n14280), .B(n14281), .Z(n12473) );
  XOR U13835 ( .A(n14282), .B(n7964), .Z(n6260) );
  XOR U13836 ( .A(n9177), .B(n14283), .Z(n7964) );
  XOR U13837 ( .A(n14284), .B(n14285), .Z(n11756) );
  XNOR U13838 ( .A(n11239), .B(n12075), .Z(n14285) );
  XOR U13839 ( .A(n14286), .B(n12501), .Z(n12075) );
  IV U13840 ( .A(n14287), .Z(n12501) );
  NOR U13841 ( .A(n13566), .B(n14288), .Z(n14286) );
  XOR U13842 ( .A(n14289), .B(n12504), .Z(n11239) );
  ANDN U13843 ( .B(n13560), .A(n14290), .Z(n14289) );
  XOR U13844 ( .A(n11722), .B(n14291), .Z(n14284) );
  XOR U13845 ( .A(n9783), .B(n11923), .Z(n14291) );
  XNOR U13846 ( .A(n14292), .B(n12488), .Z(n11923) );
  AND U13847 ( .A(n14293), .B(n13564), .Z(n14292) );
  XNOR U13848 ( .A(n14294), .B(n12496), .Z(n9783) );
  NOR U13849 ( .A(n14295), .B(n14296), .Z(n14294) );
  XOR U13850 ( .A(n14297), .B(n12492), .Z(n11722) );
  IV U13851 ( .A(n14298), .Z(n12492) );
  ANDN U13852 ( .B(n14299), .A(n13568), .Z(n14297) );
  XNOR U13853 ( .A(n14300), .B(n14301), .Z(n12687) );
  XNOR U13854 ( .A(n12136), .B(n10700), .Z(n14301) );
  XOR U13855 ( .A(n14302), .B(n14303), .Z(n10700) );
  NOR U13856 ( .A(n14304), .B(n14305), .Z(n14302) );
  XNOR U13857 ( .A(n14306), .B(n14307), .Z(n12136) );
  ANDN U13858 ( .B(n14308), .A(n14309), .Z(n14306) );
  XOR U13859 ( .A(n12885), .B(n14310), .Z(n14300) );
  XOR U13860 ( .A(n14311), .B(n14312), .Z(n14310) );
  XNOR U13861 ( .A(n14313), .B(n14314), .Z(n12885) );
  ANDN U13862 ( .B(n14315), .A(n12426), .Z(n14313) );
  ANDN U13863 ( .B(n13650), .A(n7963), .Z(n14282) );
  XOR U13864 ( .A(n14316), .B(n7968), .Z(n3157) );
  XOR U13865 ( .A(n10917), .B(n14317), .Z(n7968) );
  XNOR U13866 ( .A(n14318), .B(n14319), .Z(n10917) );
  ANDN U13867 ( .B(n9040), .A(n7967), .Z(n14316) );
  XNOR U13868 ( .A(n12814), .B(n9163), .Z(n7967) );
  XNOR U13869 ( .A(n14320), .B(n14321), .Z(n12814) );
  XNOR U13870 ( .A(n12082), .B(n14324), .Z(n9040) );
  XOR U13871 ( .A(n13553), .B(n14325), .Z(n12082) );
  XOR U13872 ( .A(n14326), .B(n14327), .Z(n13553) );
  XNOR U13873 ( .A(n11426), .B(n11003), .Z(n14327) );
  XOR U13874 ( .A(n14328), .B(n14329), .Z(n11003) );
  ANDN U13875 ( .B(n13063), .A(n14330), .Z(n14328) );
  XOR U13876 ( .A(n14331), .B(n14332), .Z(n11426) );
  AND U13877 ( .A(n13059), .B(n14333), .Z(n14331) );
  XOR U13878 ( .A(n14334), .B(n14335), .Z(n14326) );
  XOR U13879 ( .A(n9503), .B(n11863), .Z(n14335) );
  XOR U13880 ( .A(n14336), .B(n14337), .Z(n11863) );
  XOR U13881 ( .A(n14339), .B(n14340), .Z(n9503) );
  NOR U13882 ( .A(n14341), .B(n13067), .Z(n14339) );
  XOR U13883 ( .A(n14342), .B(n14343), .Z(n9983) );
  XOR U13884 ( .A(n5243), .B(n1944), .Z(n14343) );
  XNOR U13885 ( .A(n14344), .B(n9132), .Z(n1944) );
  AND U13886 ( .A(n9060), .B(n8017), .Z(n14344) );
  XOR U13887 ( .A(n14345), .B(n11888), .Z(n8017) );
  XOR U13888 ( .A(n13011), .B(n10584), .Z(n9060) );
  IV U13889 ( .A(n11936), .Z(n10584) );
  XNOR U13890 ( .A(n14346), .B(n13503), .Z(n13011) );
  NOR U13891 ( .A(n14134), .B(n14347), .Z(n14346) );
  XNOR U13892 ( .A(n14348), .B(n9137), .Z(n5243) );
  AND U13893 ( .A(n9058), .B(n8009), .Z(n14348) );
  XOR U13894 ( .A(n14349), .B(n10925), .Z(n8009) );
  XNOR U13895 ( .A(n12666), .B(n13688), .Z(n10925) );
  XNOR U13896 ( .A(n14350), .B(n14351), .Z(n13688) );
  XOR U13897 ( .A(n14352), .B(n11811), .Z(n14351) );
  XNOR U13898 ( .A(n14353), .B(n14354), .Z(n11811) );
  ANDN U13899 ( .B(n14355), .A(n14356), .Z(n14353) );
  XNOR U13900 ( .A(n13604), .B(n14357), .Z(n14350) );
  XNOR U13901 ( .A(n9500), .B(n10109), .Z(n14357) );
  XNOR U13902 ( .A(n14358), .B(n14359), .Z(n10109) );
  XOR U13903 ( .A(n14362), .B(n14363), .Z(n9500) );
  ANDN U13904 ( .B(n14364), .A(n14365), .Z(n14362) );
  XOR U13905 ( .A(n14366), .B(n14367), .Z(n13604) );
  AND U13906 ( .A(n14368), .B(n14369), .Z(n14366) );
  XOR U13907 ( .A(n14370), .B(n14371), .Z(n12666) );
  XNOR U13908 ( .A(n11199), .B(n11778), .Z(n14371) );
  XNOR U13909 ( .A(n14372), .B(n14373), .Z(n11778) );
  AND U13910 ( .A(n14374), .B(n14375), .Z(n14372) );
  XOR U13911 ( .A(n14376), .B(n14377), .Z(n11199) );
  ANDN U13912 ( .B(n14378), .A(n14379), .Z(n14376) );
  XNOR U13913 ( .A(n13311), .B(n14380), .Z(n14370) );
  XOR U13914 ( .A(n12563), .B(n12048), .Z(n14380) );
  XNOR U13915 ( .A(n14381), .B(n14382), .Z(n12048) );
  ANDN U13916 ( .B(n14383), .A(n14384), .Z(n14381) );
  XNOR U13917 ( .A(n14385), .B(n14386), .Z(n12563) );
  AND U13918 ( .A(n14387), .B(n14388), .Z(n14385) );
  XOR U13919 ( .A(n14389), .B(n14390), .Z(n13311) );
  XOR U13920 ( .A(n14391), .B(n14392), .Z(n14390) );
  NAND U13921 ( .A(n6835), .B(n11365), .Z(n14392) );
  AND U13922 ( .A(n14393), .B(n14394), .Z(n14391) );
  XNOR U13923 ( .A(n14395), .B(n10005), .Z(n9058) );
  XOR U13924 ( .A(n3699), .B(n14396), .Z(n14342) );
  XOR U13925 ( .A(n9127), .B(n4169), .Z(n14396) );
  XNOR U13926 ( .A(n14397), .B(n9141), .Z(n4169) );
  ANDN U13927 ( .B(n8000), .A(n9140), .Z(n14397) );
  XNOR U13928 ( .A(n12394), .B(n14398), .Z(n9140) );
  XOR U13929 ( .A(n14399), .B(n14400), .Z(n12394) );
  ANDN U13930 ( .B(n14401), .A(n14402), .Z(n14399) );
  XOR U13931 ( .A(n10220), .B(n14403), .Z(n8000) );
  XOR U13932 ( .A(n14404), .B(n13910), .Z(n10220) );
  XNOR U13933 ( .A(n14405), .B(n14406), .Z(n13910) );
  XOR U13934 ( .A(n12155), .B(n10244), .Z(n14406) );
  XNOR U13935 ( .A(n14407), .B(n14408), .Z(n10244) );
  NOR U13936 ( .A(n14409), .B(n14410), .Z(n14407) );
  XNOR U13937 ( .A(n14411), .B(n14412), .Z(n12155) );
  ANDN U13938 ( .B(n14413), .A(n14414), .Z(n14411) );
  XOR U13939 ( .A(n11746), .B(n14415), .Z(n14405) );
  XOR U13940 ( .A(n14104), .B(n11600), .Z(n14415) );
  XOR U13941 ( .A(n14416), .B(n14417), .Z(n11600) );
  ANDN U13942 ( .B(n14418), .A(n14419), .Z(n14416) );
  XOR U13943 ( .A(n14420), .B(n14421), .Z(n14104) );
  NOR U13944 ( .A(n14422), .B(n14423), .Z(n14420) );
  XNOR U13945 ( .A(n14424), .B(n14425), .Z(n11746) );
  XNOR U13946 ( .A(n14428), .B(n9135), .Z(n9127) );
  ANDN U13947 ( .B(n9053), .A(n8004), .Z(n14428) );
  XNOR U13948 ( .A(n14429), .B(n12884), .Z(n8004) );
  XNOR U13949 ( .A(n14017), .B(n9820), .Z(n9053) );
  XNOR U13950 ( .A(n14430), .B(n14431), .Z(n9820) );
  XNOR U13951 ( .A(n14432), .B(n14433), .Z(n14017) );
  XNOR U13952 ( .A(n14434), .B(n14435), .Z(n3699) );
  AND U13953 ( .A(n9056), .B(n8013), .Z(n14434) );
  XOR U13954 ( .A(n14436), .B(n10714), .Z(n8013) );
  XOR U13955 ( .A(n14437), .B(n7963), .Z(n9038) );
  XNOR U13956 ( .A(n12728), .B(n13427), .Z(n7963) );
  XOR U13957 ( .A(n14438), .B(n14439), .Z(n13427) );
  AND U13958 ( .A(n14440), .B(n14441), .Z(n14438) );
  ANDN U13959 ( .B(n8985), .A(n13650), .Z(n14437) );
  XNOR U13960 ( .A(n9555), .B(n14442), .Z(n13650) );
  IV U13961 ( .A(n10441), .Z(n9555) );
  IV U13962 ( .A(n13651), .Z(n8985) );
  XOR U13963 ( .A(n14443), .B(n13329), .Z(n13651) );
  IV U13964 ( .A(n11888), .Z(n13329) );
  XOR U13965 ( .A(n12540), .B(n14444), .Z(n11888) );
  XOR U13966 ( .A(n14445), .B(n14446), .Z(n12540) );
  XNOR U13967 ( .A(n14447), .B(n13280), .Z(n14446) );
  XOR U13968 ( .A(n14448), .B(n14449), .Z(n13280) );
  ANDN U13969 ( .B(n14450), .A(n13669), .Z(n14448) );
  XNOR U13970 ( .A(n13508), .B(n14451), .Z(n14445) );
  XOR U13971 ( .A(n10589), .B(n12241), .Z(n14451) );
  XNOR U13972 ( .A(n14452), .B(n14453), .Z(n12241) );
  ANDN U13973 ( .B(n14454), .A(n13673), .Z(n14452) );
  XNOR U13974 ( .A(n14455), .B(n14456), .Z(n10589) );
  AND U13975 ( .A(n13664), .B(n14457), .Z(n14455) );
  XNOR U13976 ( .A(n14458), .B(n14459), .Z(n13508) );
  ANDN U13977 ( .B(n13938), .A(n14460), .Z(n14458) );
  AND U13978 ( .A(n5656), .B(n5658), .Z(n14155) );
  XOR U13979 ( .A(n11622), .B(n2088), .Z(n5658) );
  XNOR U13980 ( .A(n8318), .B(n9757), .Z(n2088) );
  XNOR U13981 ( .A(n14461), .B(n14462), .Z(n9757) );
  XOR U13982 ( .A(n5460), .B(n3592), .Z(n14462) );
  XOR U13983 ( .A(n14463), .B(n14464), .Z(n3592) );
  ANDN U13984 ( .B(n8419), .A(n8417), .Z(n14463) );
  XNOR U13985 ( .A(n11007), .B(n13090), .Z(n8419) );
  XOR U13986 ( .A(n14465), .B(n14466), .Z(n13090) );
  ANDN U13987 ( .B(n13927), .A(n13925), .Z(n14465) );
  IV U13988 ( .A(n11566), .Z(n11007) );
  XOR U13989 ( .A(n14467), .B(n14468), .Z(n11566) );
  XOR U13990 ( .A(n14469), .B(n12022), .Z(n5460) );
  ANDN U13991 ( .B(n8413), .A(n8414), .Z(n14469) );
  XOR U13992 ( .A(n10559), .B(n14470), .Z(n8414) );
  XNOR U13993 ( .A(n14471), .B(n13223), .Z(n10559) );
  XNOR U13994 ( .A(n14472), .B(n14473), .Z(n13223) );
  XNOR U13995 ( .A(n10038), .B(n9711), .Z(n14473) );
  XOR U13996 ( .A(n14474), .B(n14475), .Z(n9711) );
  ANDN U13997 ( .B(n14476), .A(n14477), .Z(n14474) );
  XOR U13998 ( .A(n14478), .B(n14479), .Z(n10038) );
  AND U13999 ( .A(n14480), .B(n14481), .Z(n14478) );
  XOR U14000 ( .A(n11377), .B(n14482), .Z(n14472) );
  XNOR U14001 ( .A(n11388), .B(n14483), .Z(n14482) );
  XOR U14002 ( .A(n14484), .B(n14485), .Z(n11388) );
  NOR U14003 ( .A(n14486), .B(n14487), .Z(n14484) );
  XNOR U14004 ( .A(n14488), .B(n14489), .Z(n11377) );
  ANDN U14005 ( .B(n14490), .A(n14491), .Z(n14488) );
  XOR U14006 ( .A(n14492), .B(n10235), .Z(n8413) );
  XOR U14007 ( .A(n6249), .B(n14493), .Z(n14461) );
  XOR U14008 ( .A(n2385), .B(n5643), .Z(n14493) );
  XNOR U14009 ( .A(n14494), .B(n12033), .Z(n5643) );
  AND U14010 ( .A(n9761), .B(n9759), .Z(n14494) );
  IV U14011 ( .A(n12034), .Z(n9759) );
  XOR U14012 ( .A(n14495), .B(n9927), .Z(n12034) );
  XNOR U14013 ( .A(n13878), .B(n13607), .Z(n9927) );
  XNOR U14014 ( .A(n14496), .B(n14497), .Z(n13607) );
  XNOR U14015 ( .A(n12363), .B(n12126), .Z(n14497) );
  XNOR U14016 ( .A(n14498), .B(n14499), .Z(n12126) );
  AND U14017 ( .A(n14500), .B(n14501), .Z(n14498) );
  XNOR U14018 ( .A(n14502), .B(n14503), .Z(n12363) );
  AND U14019 ( .A(n14504), .B(n14505), .Z(n14502) );
  XOR U14020 ( .A(n12165), .B(n14506), .Z(n14496) );
  XOR U14021 ( .A(n11059), .B(n12389), .Z(n14506) );
  XOR U14022 ( .A(n14507), .B(n14508), .Z(n12389) );
  ANDN U14023 ( .B(n14509), .A(n14510), .Z(n14507) );
  XNOR U14024 ( .A(n14511), .B(n14512), .Z(n11059) );
  AND U14025 ( .A(n14513), .B(n14514), .Z(n14511) );
  XOR U14026 ( .A(n14515), .B(n14516), .Z(n12165) );
  AND U14027 ( .A(n14517), .B(n14518), .Z(n14515) );
  XOR U14028 ( .A(n14519), .B(n14520), .Z(n13878) );
  XNOR U14029 ( .A(n12931), .B(n11176), .Z(n14520) );
  XOR U14030 ( .A(n14521), .B(n14522), .Z(n11176) );
  NOR U14031 ( .A(n14523), .B(n13985), .Z(n14521) );
  XNOR U14032 ( .A(n14524), .B(n14525), .Z(n12931) );
  NOR U14033 ( .A(n14526), .B(n14527), .Z(n14524) );
  XOR U14034 ( .A(n9765), .B(n14528), .Z(n14519) );
  XOR U14035 ( .A(n10302), .B(n14529), .Z(n14528) );
  XOR U14036 ( .A(n14530), .B(n14531), .Z(n10302) );
  ANDN U14037 ( .B(n13977), .A(n14532), .Z(n14530) );
  XOR U14038 ( .A(n14533), .B(n14534), .Z(n9765) );
  ANDN U14039 ( .B(n14535), .A(n13968), .Z(n14533) );
  XNOR U14040 ( .A(n14536), .B(n11320), .Z(n9761) );
  XNOR U14041 ( .A(n14537), .B(n12025), .Z(n2385) );
  ANDN U14042 ( .B(n8405), .A(n8403), .Z(n14537) );
  XOR U14043 ( .A(n14538), .B(n10943), .Z(n8403) );
  XNOR U14044 ( .A(n14034), .B(n10017), .Z(n8405) );
  XOR U14045 ( .A(n14539), .B(n14540), .Z(n14034) );
  NOR U14046 ( .A(n14541), .B(n14542), .Z(n14539) );
  XNOR U14047 ( .A(n14543), .B(n12030), .Z(n6249) );
  ANDN U14048 ( .B(n8409), .A(n8407), .Z(n14543) );
  XOR U14049 ( .A(n14544), .B(n11055), .Z(n8407) );
  XOR U14050 ( .A(n14545), .B(n11908), .Z(n8409) );
  XNOR U14051 ( .A(n10489), .B(n14546), .Z(n11908) );
  XOR U14052 ( .A(n14547), .B(n14548), .Z(n10489) );
  XOR U14053 ( .A(n11851), .B(n11022), .Z(n14548) );
  XOR U14054 ( .A(n14549), .B(n14550), .Z(n11022) );
  ANDN U14055 ( .B(n14551), .A(n14552), .Z(n14549) );
  XNOR U14056 ( .A(n14553), .B(n13719), .Z(n11851) );
  ANDN U14057 ( .B(n13720), .A(n14554), .Z(n14553) );
  XOR U14058 ( .A(n10036), .B(n14555), .Z(n14547) );
  XOR U14059 ( .A(n9184), .B(n10950), .Z(n14555) );
  XNOR U14060 ( .A(n14556), .B(n13709), .Z(n10950) );
  AND U14061 ( .A(n14557), .B(n13710), .Z(n14556) );
  XNOR U14062 ( .A(n14558), .B(n13715), .Z(n9184) );
  XNOR U14063 ( .A(n14560), .B(n13705), .Z(n10036) );
  ANDN U14064 ( .B(n13706), .A(n14561), .Z(n14560) );
  XOR U14065 ( .A(n14562), .B(n14563), .Z(n8318) );
  XOR U14066 ( .A(n3805), .B(n5119), .Z(n14563) );
  XOR U14067 ( .A(n14564), .B(n9653), .Z(n5119) );
  IV U14068 ( .A(n12012), .Z(n9653) );
  XOR U14069 ( .A(n14565), .B(n9704), .Z(n12012) );
  ANDN U14070 ( .B(n11628), .A(n11629), .Z(n14564) );
  XOR U14071 ( .A(n14566), .B(n11793), .Z(n11629) );
  XOR U14072 ( .A(n14567), .B(n10943), .Z(n11628) );
  XNOR U14073 ( .A(n11542), .B(n12797), .Z(n10943) );
  XNOR U14074 ( .A(n14568), .B(n14569), .Z(n12797) );
  XNOR U14075 ( .A(n14570), .B(n11164), .Z(n14569) );
  XOR U14076 ( .A(n14571), .B(n14572), .Z(n11164) );
  AND U14077 ( .A(n14573), .B(n14574), .Z(n14571) );
  XNOR U14078 ( .A(n9942), .B(n14575), .Z(n14568) );
  XOR U14079 ( .A(n10899), .B(n12570), .Z(n14575) );
  XOR U14080 ( .A(n14576), .B(n14577), .Z(n12570) );
  ANDN U14081 ( .B(n14578), .A(n14579), .Z(n14576) );
  XOR U14082 ( .A(n14580), .B(n14581), .Z(n10899) );
  AND U14083 ( .A(n14582), .B(n14583), .Z(n14580) );
  XOR U14084 ( .A(n14584), .B(n14585), .Z(n9942) );
  AND U14085 ( .A(n14586), .B(n14587), .Z(n14584) );
  XOR U14086 ( .A(n14588), .B(n14589), .Z(n11542) );
  XNOR U14087 ( .A(n9359), .B(n12472), .Z(n14589) );
  XOR U14088 ( .A(n14590), .B(n13638), .Z(n12472) );
  IV U14089 ( .A(n14591), .Z(n13638) );
  NOR U14090 ( .A(n14592), .B(n14433), .Z(n14590) );
  XOR U14091 ( .A(n14593), .B(n13645), .Z(n9359) );
  XOR U14092 ( .A(n10889), .B(n14595), .Z(n14588) );
  XOR U14093 ( .A(n14279), .B(n12314), .Z(n14595) );
  XNOR U14094 ( .A(n14596), .B(n13632), .Z(n12314) );
  ANDN U14095 ( .B(n14597), .A(n14019), .Z(n14596) );
  XOR U14096 ( .A(n14598), .B(n13641), .Z(n14279) );
  NOR U14097 ( .A(n14599), .B(n14025), .Z(n14598) );
  XNOR U14098 ( .A(n14600), .B(n13628), .Z(n10889) );
  ANDN U14099 ( .B(n14601), .A(n14028), .Z(n14600) );
  XNOR U14100 ( .A(n14602), .B(n8351), .Z(n3805) );
  XNOR U14101 ( .A(n14603), .B(n10293), .Z(n8351) );
  IV U14102 ( .A(n13648), .Z(n10293) );
  XNOR U14103 ( .A(n14604), .B(n13323), .Z(n13648) );
  XNOR U14104 ( .A(n14605), .B(n14606), .Z(n13323) );
  XOR U14105 ( .A(n13596), .B(n12920), .Z(n14606) );
  XOR U14106 ( .A(n14607), .B(n14608), .Z(n12920) );
  AND U14107 ( .A(n13176), .B(n13178), .Z(n14607) );
  XNOR U14108 ( .A(n14609), .B(n14610), .Z(n13596) );
  ANDN U14109 ( .B(n14611), .A(n13168), .Z(n14609) );
  XOR U14110 ( .A(n11569), .B(n14612), .Z(n14605) );
  XOR U14111 ( .A(n13658), .B(n12989), .Z(n14612) );
  XNOR U14112 ( .A(n14613), .B(n14614), .Z(n12989) );
  ANDN U14113 ( .B(n13174), .A(n13172), .Z(n14613) );
  XNOR U14114 ( .A(n14615), .B(n14616), .Z(n13658) );
  AND U14115 ( .A(n14617), .B(n13163), .Z(n14615) );
  XNOR U14116 ( .A(n14618), .B(n14619), .Z(n11569) );
  AND U14117 ( .A(n13325), .B(n14620), .Z(n14618) );
  NOR U14118 ( .A(n11620), .B(n11621), .Z(n14602) );
  XOR U14119 ( .A(n11649), .B(n14222), .Z(n11621) );
  XNOR U14120 ( .A(n14621), .B(n14180), .Z(n14222) );
  NOR U14121 ( .A(n14622), .B(n13518), .Z(n14621) );
  XNOR U14122 ( .A(n14623), .B(n10123), .Z(n11620) );
  IV U14123 ( .A(n10270), .Z(n10123) );
  XNOR U14124 ( .A(n5463), .B(n14624), .Z(n14562) );
  XOR U14125 ( .A(n1741), .B(n12006), .Z(n14624) );
  XOR U14126 ( .A(n14625), .B(n8360), .Z(n12006) );
  XOR U14127 ( .A(n14626), .B(n12444), .Z(n8360) );
  XOR U14128 ( .A(n14627), .B(n13512), .Z(n12444) );
  XNOR U14129 ( .A(n14628), .B(n14629), .Z(n13512) );
  XNOR U14130 ( .A(n14630), .B(n14631), .Z(n14629) );
  XOR U14131 ( .A(n9572), .B(n14632), .Z(n14628) );
  XNOR U14132 ( .A(n13267), .B(n14633), .Z(n14632) );
  XNOR U14133 ( .A(n14634), .B(n14635), .Z(n13267) );
  ANDN U14134 ( .B(n14636), .A(n14061), .Z(n14634) );
  XOR U14135 ( .A(n14637), .B(n14638), .Z(n9572) );
  ANDN U14136 ( .B(n14639), .A(n14640), .Z(n14637) );
  XOR U14137 ( .A(n14641), .B(n11761), .Z(n11617) );
  XNOR U14138 ( .A(n14642), .B(n13374), .Z(n11761) );
  XNOR U14139 ( .A(n14643), .B(n14644), .Z(n13374) );
  XNOR U14140 ( .A(n10153), .B(n12154), .Z(n14644) );
  XNOR U14141 ( .A(n14645), .B(n14646), .Z(n12154) );
  AND U14142 ( .A(n14647), .B(n14648), .Z(n14645) );
  XNOR U14143 ( .A(n14649), .B(n14650), .Z(n10153) );
  AND U14144 ( .A(n14651), .B(n14652), .Z(n14649) );
  XNOR U14145 ( .A(n14653), .B(n14654), .Z(n14643) );
  XNOR U14146 ( .A(n11250), .B(n11013), .Z(n14654) );
  XNOR U14147 ( .A(n14655), .B(n14656), .Z(n11013) );
  ANDN U14148 ( .B(n14657), .A(n14658), .Z(n14655) );
  XOR U14149 ( .A(n14659), .B(n14660), .Z(n11250) );
  ANDN U14150 ( .B(n14661), .A(n14662), .Z(n14659) );
  XOR U14151 ( .A(n10544), .B(n14663), .Z(n11618) );
  XOR U14152 ( .A(n14664), .B(n8354), .Z(n1741) );
  IV U14153 ( .A(n12010), .Z(n8354) );
  XOR U14154 ( .A(n14665), .B(n10373), .Z(n12010) );
  XNOR U14155 ( .A(n14666), .B(n14667), .Z(n13905) );
  XOR U14156 ( .A(n14668), .B(n12581), .Z(n14667) );
  XOR U14157 ( .A(n14669), .B(n14670), .Z(n12581) );
  XOR U14158 ( .A(n13183), .B(n14672), .Z(n14666) );
  XOR U14159 ( .A(n11674), .B(n11601), .Z(n14672) );
  XOR U14160 ( .A(n14673), .B(n14674), .Z(n11601) );
  ANDN U14161 ( .B(n13306), .A(n14675), .Z(n14673) );
  XNOR U14162 ( .A(n14676), .B(n14677), .Z(n11674) );
  AND U14163 ( .A(n14678), .B(n14679), .Z(n14676) );
  XOR U14164 ( .A(n14680), .B(n14681), .Z(n13183) );
  ANDN U14165 ( .B(n13298), .A(n14682), .Z(n14680) );
  NOR U14166 ( .A(n11626), .B(n11625), .Z(n14664) );
  XNOR U14167 ( .A(n10441), .B(n14684), .Z(n11625) );
  XOR U14168 ( .A(n14685), .B(n12710), .Z(n10441) );
  XOR U14169 ( .A(n14686), .B(n14687), .Z(n12710) );
  XNOR U14170 ( .A(n13466), .B(n12672), .Z(n14687) );
  XOR U14171 ( .A(n14688), .B(n13825), .Z(n12672) );
  AND U14172 ( .A(n14689), .B(n14690), .Z(n14688) );
  XNOR U14173 ( .A(n14691), .B(n13833), .Z(n13466) );
  ANDN U14174 ( .B(n14692), .A(n14693), .Z(n14691) );
  XNOR U14175 ( .A(n11660), .B(n14694), .Z(n14686) );
  XOR U14176 ( .A(n10002), .B(n9102), .Z(n14694) );
  XNOR U14177 ( .A(n14695), .B(n13829), .Z(n9102) );
  AND U14178 ( .A(n14696), .B(n14697), .Z(n14695) );
  XNOR U14179 ( .A(n14698), .B(n13820), .Z(n10002) );
  AND U14180 ( .A(n14699), .B(n14700), .Z(n14698) );
  XOR U14181 ( .A(n14701), .B(n14702), .Z(n11660) );
  ANDN U14182 ( .B(n14703), .A(n14704), .Z(n14701) );
  XNOR U14183 ( .A(n14705), .B(n10126), .Z(n11626) );
  XNOR U14184 ( .A(n14706), .B(n8365), .Z(n5463) );
  XOR U14185 ( .A(n14707), .B(n10235), .Z(n8365) );
  ANDN U14186 ( .B(n12015), .A(n13916), .Z(n14706) );
  XOR U14187 ( .A(n14708), .B(n12015), .Z(n11622) );
  XNOR U14188 ( .A(n13534), .B(n9900), .Z(n12015) );
  IV U14189 ( .A(n11515), .Z(n9900) );
  XNOR U14190 ( .A(n14709), .B(n14710), .Z(n11515) );
  XOR U14191 ( .A(n14711), .B(n14712), .Z(n13534) );
  ANDN U14192 ( .B(n14167), .A(n14165), .Z(n14711) );
  AND U14193 ( .A(n13916), .B(n13917), .Z(n14708) );
  XOR U14194 ( .A(n14713), .B(n13315), .Z(n13917) );
  XNOR U14195 ( .A(n12205), .B(n14714), .Z(n13916) );
  XOR U14196 ( .A(n14715), .B(n14716), .Z(n11849) );
  XNOR U14197 ( .A(n10771), .B(n11276), .Z(n14716) );
  XOR U14198 ( .A(n14717), .B(n14718), .Z(n11276) );
  AND U14199 ( .A(n14719), .B(n14720), .Z(n14717) );
  NOR U14200 ( .A(n14723), .B(n14724), .Z(n14721) );
  XNOR U14201 ( .A(n10285), .B(n14725), .Z(n14715) );
  XOR U14202 ( .A(n9363), .B(n11153), .Z(n14725) );
  XNOR U14203 ( .A(n14726), .B(n14727), .Z(n11153) );
  ANDN U14204 ( .B(n14728), .A(n14729), .Z(n14726) );
  XNOR U14205 ( .A(n14730), .B(n14731), .Z(n9363) );
  XOR U14206 ( .A(n14734), .B(n14735), .Z(n10285) );
  ANDN U14207 ( .B(n14736), .A(n14737), .Z(n14734) );
  XOR U14208 ( .A(n14738), .B(n14739), .Z(n11943) );
  XOR U14209 ( .A(n11378), .B(n10144), .Z(n14739) );
  XOR U14210 ( .A(n14740), .B(n14741), .Z(n10144) );
  ANDN U14211 ( .B(n14742), .A(n14743), .Z(n14740) );
  XOR U14212 ( .A(n14744), .B(n14745), .Z(n11378) );
  AND U14213 ( .A(n14746), .B(n14747), .Z(n14744) );
  XNOR U14214 ( .A(n14748), .B(n14749), .Z(n14738) );
  XOR U14215 ( .A(n9527), .B(n14750), .Z(n14749) );
  XOR U14216 ( .A(n14751), .B(n14752), .Z(n9527) );
  ANDN U14217 ( .B(n14753), .A(n14754), .Z(n14751) );
  XNOR U14218 ( .A(n8897), .B(n4249), .Z(n5656) );
  XNOR U14219 ( .A(n14755), .B(n14756), .Z(n6468) );
  XNOR U14220 ( .A(n5806), .B(n2529), .Z(n14756) );
  XNOR U14221 ( .A(n14757), .B(n6517), .Z(n2529) );
  XNOR U14222 ( .A(n9079), .B(n14758), .Z(n6517) );
  IV U14223 ( .A(n13043), .Z(n9079) );
  XOR U14224 ( .A(n12941), .B(n14759), .Z(n13043) );
  XOR U14225 ( .A(n14760), .B(n14761), .Z(n12941) );
  XOR U14226 ( .A(n9081), .B(n11560), .Z(n14761) );
  XOR U14227 ( .A(n14762), .B(n14763), .Z(n11560) );
  ANDN U14228 ( .B(n14764), .A(n14765), .Z(n14762) );
  XOR U14229 ( .A(n14766), .B(n14767), .Z(n9081) );
  ANDN U14230 ( .B(n14768), .A(n14769), .Z(n14766) );
  XNOR U14231 ( .A(n14770), .B(n14771), .Z(n14760) );
  XOR U14232 ( .A(n14772), .B(n11460), .Z(n14771) );
  XOR U14233 ( .A(n14773), .B(n14774), .Z(n11460) );
  NOR U14234 ( .A(n14775), .B(n14776), .Z(n14773) );
  ANDN U14235 ( .B(n8902), .A(n8903), .Z(n14757) );
  XNOR U14236 ( .A(n14777), .B(n10806), .Z(n8903) );
  XNOR U14237 ( .A(n14468), .B(n14778), .Z(n10806) );
  XOR U14238 ( .A(n14779), .B(n14780), .Z(n14468) );
  XNOR U14239 ( .A(n14781), .B(n10705), .Z(n14780) );
  XOR U14240 ( .A(n14782), .B(n14783), .Z(n10705) );
  ANDN U14241 ( .B(n14784), .A(n14363), .Z(n14782) );
  XNOR U14242 ( .A(n12280), .B(n14785), .Z(n14779) );
  XOR U14243 ( .A(n12542), .B(n12532), .Z(n14785) );
  XNOR U14244 ( .A(n14786), .B(n14787), .Z(n12532) );
  ANDN U14245 ( .B(n14788), .A(n14367), .Z(n14786) );
  XNOR U14246 ( .A(n14789), .B(n14790), .Z(n12542) );
  XOR U14247 ( .A(n14793), .B(n14794), .Z(n12280) );
  XNOR U14248 ( .A(n12779), .B(n11126), .Z(n8902) );
  XOR U14249 ( .A(n14796), .B(n14797), .Z(n12779) );
  NOR U14250 ( .A(n14798), .B(n14799), .Z(n14796) );
  XNOR U14251 ( .A(n14800), .B(n6509), .Z(n5806) );
  XOR U14252 ( .A(n14801), .B(n10219), .Z(n6509) );
  XNOR U14253 ( .A(n14802), .B(n12612), .Z(n10219) );
  XNOR U14254 ( .A(n14803), .B(n14804), .Z(n12612) );
  XOR U14255 ( .A(n12700), .B(n11451), .Z(n14804) );
  XOR U14256 ( .A(n14805), .B(n14273), .Z(n11451) );
  AND U14257 ( .A(n14274), .B(n14806), .Z(n14805) );
  XOR U14258 ( .A(n14807), .B(n14265), .Z(n12700) );
  AND U14259 ( .A(n14264), .B(n14808), .Z(n14807) );
  XOR U14260 ( .A(n12690), .B(n14809), .Z(n14803) );
  XOR U14261 ( .A(n11703), .B(n10477), .Z(n14809) );
  XNOR U14262 ( .A(n14810), .B(n14269), .Z(n10477) );
  AND U14263 ( .A(n14811), .B(n14812), .Z(n14810) );
  XNOR U14264 ( .A(n14813), .B(n14814), .Z(n11703) );
  AND U14265 ( .A(n14815), .B(n14816), .Z(n14813) );
  XOR U14266 ( .A(n14817), .B(n14818), .Z(n12690) );
  ANDN U14267 ( .B(n14278), .A(n14819), .Z(n14817) );
  AND U14268 ( .A(n13852), .B(n14820), .Z(n14800) );
  XOR U14269 ( .A(n3471), .B(n14821), .Z(n14755) );
  XNOR U14270 ( .A(n8937), .B(n4855), .Z(n14821) );
  XOR U14271 ( .A(n14822), .B(n6504), .Z(n4855) );
  IV U14272 ( .A(n8942), .Z(n6504) );
  XOR U14273 ( .A(n14823), .B(n12662), .Z(n8942) );
  ANDN U14274 ( .B(n8899), .A(n8900), .Z(n14822) );
  XNOR U14275 ( .A(n14824), .B(n11373), .Z(n8900) );
  XNOR U14276 ( .A(n11386), .B(n13432), .Z(n8899) );
  XNOR U14277 ( .A(n14825), .B(n14826), .Z(n13432) );
  AND U14278 ( .A(n14827), .B(n14828), .Z(n14825) );
  IV U14279 ( .A(n12728), .Z(n11386) );
  XNOR U14280 ( .A(n13814), .B(n14829), .Z(n12728) );
  XOR U14281 ( .A(n14830), .B(n14831), .Z(n13814) );
  XNOR U14282 ( .A(n9707), .B(n10209), .Z(n14831) );
  XNOR U14283 ( .A(n14832), .B(n14833), .Z(n10209) );
  AND U14284 ( .A(n13260), .B(n14834), .Z(n14832) );
  XNOR U14285 ( .A(n14835), .B(n14836), .Z(n9707) );
  ANDN U14286 ( .B(n14837), .A(n13250), .Z(n14835) );
  XOR U14287 ( .A(n13680), .B(n14838), .Z(n14830) );
  XNOR U14288 ( .A(n9484), .B(n14123), .Z(n14838) );
  XNOR U14289 ( .A(n14839), .B(n14840), .Z(n14123) );
  AND U14290 ( .A(n14841), .B(n14842), .Z(n14839) );
  XNOR U14291 ( .A(n14843), .B(n14844), .Z(n9484) );
  NOR U14292 ( .A(n13254), .B(n14845), .Z(n14843) );
  XNOR U14293 ( .A(n14846), .B(n14847), .Z(n13680) );
  ANDN U14294 ( .B(n14848), .A(n13264), .Z(n14846) );
  XOR U14295 ( .A(n14849), .B(n6500), .Z(n8937) );
  XOR U14296 ( .A(n11593), .B(n13234), .Z(n6500) );
  XNOR U14297 ( .A(n14850), .B(n14851), .Z(n13234) );
  AND U14298 ( .A(n13761), .B(n13763), .Z(n14850) );
  IV U14299 ( .A(n11691), .Z(n11593) );
  ANDN U14300 ( .B(n8894), .A(n8893), .Z(n14849) );
  XOR U14301 ( .A(n14852), .B(n10448), .Z(n8893) );
  XOR U14302 ( .A(n14853), .B(n11307), .Z(n8894) );
  IV U14303 ( .A(n11192), .Z(n11307) );
  XNOR U14304 ( .A(n14854), .B(n6513), .Z(n3471) );
  XOR U14305 ( .A(n14855), .B(n9720), .Z(n6513) );
  IV U14306 ( .A(n9699), .Z(n9720) );
  XOR U14307 ( .A(n14856), .B(n13396), .Z(n9699) );
  XNOR U14308 ( .A(n14857), .B(n14858), .Z(n13396) );
  XNOR U14309 ( .A(n13513), .B(n10054), .Z(n14858) );
  XOR U14310 ( .A(n14859), .B(n14860), .Z(n10054) );
  AND U14311 ( .A(n14861), .B(n14862), .Z(n14859) );
  XNOR U14312 ( .A(n14863), .B(n14864), .Z(n13513) );
  ANDN U14313 ( .B(n14865), .A(n14866), .Z(n14863) );
  XOR U14314 ( .A(n10158), .B(n14867), .Z(n14857) );
  XNOR U14315 ( .A(n12647), .B(n14868), .Z(n14867) );
  XOR U14316 ( .A(n14869), .B(n14870), .Z(n12647) );
  AND U14317 ( .A(n14871), .B(n14872), .Z(n14869) );
  XNOR U14318 ( .A(n14873), .B(n14874), .Z(n10158) );
  ANDN U14319 ( .B(n14875), .A(n14876), .Z(n14873) );
  AND U14320 ( .A(n8890), .B(n8947), .Z(n14854) );
  XOR U14321 ( .A(n14877), .B(n9790), .Z(n8947) );
  IV U14322 ( .A(n10096), .Z(n9790) );
  XOR U14323 ( .A(n14878), .B(n14879), .Z(n10096) );
  XNOR U14324 ( .A(n14880), .B(n12210), .Z(n8890) );
  XNOR U14325 ( .A(n14881), .B(n14882), .Z(n6291) );
  XOR U14326 ( .A(n5431), .B(n3680), .Z(n14882) );
  XOR U14327 ( .A(n14883), .B(n14884), .Z(n3680) );
  ANDN U14328 ( .B(n6528), .A(n6529), .Z(n14883) );
  XOR U14329 ( .A(n12780), .B(n11126), .Z(n6529) );
  IV U14330 ( .A(n10000), .Z(n11126) );
  XOR U14331 ( .A(n14885), .B(n14886), .Z(n12611) );
  XOR U14332 ( .A(n11398), .B(n9779), .Z(n14886) );
  XOR U14333 ( .A(n14887), .B(n14888), .Z(n9779) );
  AND U14334 ( .A(n14889), .B(n14890), .Z(n14887) );
  XOR U14335 ( .A(n14891), .B(n14892), .Z(n11398) );
  ANDN U14336 ( .B(n14893), .A(n12782), .Z(n14891) );
  XOR U14337 ( .A(n10874), .B(n14894), .Z(n14885) );
  XOR U14338 ( .A(n12066), .B(n14895), .Z(n14894) );
  XOR U14339 ( .A(n14896), .B(n14897), .Z(n12066) );
  ANDN U14340 ( .B(n12773), .A(n12771), .Z(n14896) );
  XNOR U14341 ( .A(n14898), .B(n14899), .Z(n10874) );
  ANDN U14342 ( .B(n12775), .A(n12776), .Z(n14898) );
  XNOR U14343 ( .A(n14900), .B(n14901), .Z(n13376) );
  XNOR U14344 ( .A(n9175), .B(n12167), .Z(n14901) );
  XOR U14345 ( .A(n14902), .B(n14903), .Z(n12167) );
  XNOR U14346 ( .A(n14904), .B(n14905), .Z(n13118) );
  XNOR U14347 ( .A(n14906), .B(n14907), .Z(n9175) );
  AND U14348 ( .A(n12959), .B(n14908), .Z(n14906) );
  XOR U14349 ( .A(n14909), .B(n14910), .Z(n12959) );
  XOR U14350 ( .A(n10654), .B(n14911), .Z(n14900) );
  XOR U14351 ( .A(n13045), .B(n11985), .Z(n14911) );
  XNOR U14352 ( .A(n14912), .B(n14913), .Z(n11985) );
  ANDN U14353 ( .B(n13131), .A(n12950), .Z(n14912) );
  XOR U14354 ( .A(n14914), .B(n14915), .Z(n12950) );
  XNOR U14355 ( .A(n14916), .B(n14917), .Z(n13045) );
  ANDN U14356 ( .B(n13125), .A(n12955), .Z(n14916) );
  XNOR U14357 ( .A(n14918), .B(n14919), .Z(n12955) );
  XNOR U14358 ( .A(n14920), .B(n14921), .Z(n10654) );
  ANDN U14359 ( .B(n14922), .A(n12963), .Z(n14920) );
  XOR U14360 ( .A(n14923), .B(n14924), .Z(n12963) );
  XNOR U14361 ( .A(n14925), .B(n14926), .Z(n12780) );
  NOR U14362 ( .A(n14889), .B(n14927), .Z(n14925) );
  XNOR U14363 ( .A(n14928), .B(n8956), .Z(n5431) );
  ANDN U14364 ( .B(n8957), .A(n6538), .Z(n14928) );
  XNOR U14365 ( .A(n14929), .B(n13075), .Z(n6538) );
  XOR U14366 ( .A(n14930), .B(n11979), .Z(n8957) );
  XNOR U14367 ( .A(n4293), .B(n14931), .Z(n14881) );
  XOR U14368 ( .A(n5870), .B(n2123), .Z(n14931) );
  XOR U14369 ( .A(n14932), .B(n8953), .Z(n2123) );
  AND U14370 ( .A(n6535), .B(n6533), .Z(n14932) );
  XNOR U14371 ( .A(n14933), .B(n9659), .Z(n6533) );
  XOR U14372 ( .A(n14934), .B(n12223), .Z(n9659) );
  XOR U14373 ( .A(n14935), .B(n14936), .Z(n12223) );
  XNOR U14374 ( .A(n14495), .B(n12375), .Z(n14936) );
  XOR U14375 ( .A(n14937), .B(n14938), .Z(n12375) );
  ANDN U14376 ( .B(n13972), .A(n13974), .Z(n14937) );
  XOR U14377 ( .A(n14939), .B(n14535), .Z(n14495) );
  AND U14378 ( .A(n13970), .B(n13968), .Z(n14939) );
  XNOR U14379 ( .A(n14940), .B(n14941), .Z(n13968) );
  XNOR U14380 ( .A(n12041), .B(n14942), .Z(n14935) );
  XOR U14381 ( .A(n9926), .B(n12704), .Z(n14942) );
  XNOR U14382 ( .A(n14943), .B(n14523), .Z(n12704) );
  ANDN U14383 ( .B(n13985), .A(n13986), .Z(n14943) );
  XOR U14384 ( .A(n14944), .B(n14945), .Z(n13985) );
  XNOR U14385 ( .A(n14946), .B(n14532), .Z(n9926) );
  NOR U14386 ( .A(n13978), .B(n13977), .Z(n14946) );
  XOR U14387 ( .A(n14947), .B(n14948), .Z(n13977) );
  XNOR U14388 ( .A(n14949), .B(n14527), .Z(n12041) );
  AND U14389 ( .A(n13983), .B(n14526), .Z(n14949) );
  IV U14390 ( .A(n13981), .Z(n14526) );
  XOR U14391 ( .A(n14950), .B(n14951), .Z(n13981) );
  XNOR U14392 ( .A(n10359), .B(n14952), .Z(n6535) );
  XOR U14393 ( .A(n14953), .B(n8965), .Z(n5870) );
  ANDN U14394 ( .B(n8966), .A(n6526), .Z(n14953) );
  XNOR U14395 ( .A(n9526), .B(n14750), .Z(n6526) );
  XOR U14396 ( .A(n14954), .B(n14955), .Z(n14750) );
  NOR U14397 ( .A(n14956), .B(n14957), .Z(n14954) );
  XOR U14398 ( .A(n10374), .B(n14958), .Z(n8966) );
  XNOR U14399 ( .A(n14959), .B(n8962), .Z(n4293) );
  AND U14400 ( .A(n6541), .B(n6543), .Z(n14959) );
  XNOR U14401 ( .A(n14960), .B(n9704), .Z(n6543) );
  XNOR U14402 ( .A(n14961), .B(n14829), .Z(n9704) );
  XNOR U14403 ( .A(n14962), .B(n14963), .Z(n14829) );
  XNOR U14404 ( .A(n11516), .B(n12459), .Z(n14963) );
  XNOR U14405 ( .A(n14964), .B(n14965), .Z(n12459) );
  ANDN U14406 ( .B(n14826), .A(n14827), .Z(n14964) );
  XNOR U14407 ( .A(n14966), .B(n14967), .Z(n11516) );
  NOR U14408 ( .A(n14440), .B(n14439), .Z(n14966) );
  XNOR U14409 ( .A(n10696), .B(n14968), .Z(n14962) );
  XNOR U14410 ( .A(n11270), .B(n14969), .Z(n14968) );
  XOR U14411 ( .A(n14970), .B(n14971), .Z(n11270) );
  ANDN U14412 ( .B(n13435), .A(n13436), .Z(n14970) );
  XNOR U14413 ( .A(n14972), .B(n14973), .Z(n10696) );
  ANDN U14414 ( .B(n13431), .A(n13429), .Z(n14972) );
  XNOR U14415 ( .A(n14974), .B(n11192), .Z(n6541) );
  XNOR U14416 ( .A(n14975), .B(n11534), .Z(n11192) );
  XNOR U14417 ( .A(n14976), .B(n14977), .Z(n11534) );
  XNOR U14418 ( .A(n12698), .B(n11563), .Z(n14977) );
  XNOR U14419 ( .A(n14978), .B(n14979), .Z(n11563) );
  AND U14420 ( .A(n14980), .B(n14981), .Z(n14978) );
  XNOR U14421 ( .A(n14982), .B(n14983), .Z(n12698) );
  ANDN U14422 ( .B(n14984), .A(n14985), .Z(n14982) );
  XNOR U14423 ( .A(n9400), .B(n14986), .Z(n14976) );
  XOR U14424 ( .A(n14987), .B(n12668), .Z(n14986) );
  XNOR U14425 ( .A(n14988), .B(n14989), .Z(n12668) );
  ANDN U14426 ( .B(n14990), .A(n14991), .Z(n14988) );
  XNOR U14427 ( .A(n14992), .B(n14993), .Z(n9400) );
  AND U14428 ( .A(n14994), .B(n14995), .Z(n14992) );
  XOR U14429 ( .A(n14996), .B(n8945), .Z(n8897) );
  IV U14430 ( .A(n14820), .Z(n8945) );
  XNOR U14431 ( .A(n14997), .B(n12366), .Z(n14820) );
  NOR U14432 ( .A(n6507), .B(n13852), .Z(n14996) );
  XOR U14433 ( .A(n14998), .B(n11837), .Z(n13852) );
  XNOR U14434 ( .A(n14115), .B(n11464), .Z(n6507) );
  IV U14435 ( .A(n11544), .Z(n11464) );
  XOR U14436 ( .A(n14999), .B(n15000), .Z(n11544) );
  XNOR U14437 ( .A(n15001), .B(n15002), .Z(n14115) );
  ANDN U14438 ( .B(n15003), .A(n15004), .Z(n15001) );
  XOR U14439 ( .A(n15005), .B(n6178), .Z(out[1000]) );
  XOR U14440 ( .A(n9130), .B(n2307), .Z(n6178) );
  XNOR U14441 ( .A(n10085), .B(n6138), .Z(n2307) );
  XNOR U14442 ( .A(n15006), .B(n15007), .Z(n6138) );
  XOR U14443 ( .A(n2343), .B(n5447), .Z(n15007) );
  XOR U14444 ( .A(n15008), .B(n8002), .Z(n5447) );
  XOR U14445 ( .A(n11538), .B(n13527), .Z(n8002) );
  XNOR U14446 ( .A(n15009), .B(n14225), .Z(n13527) );
  NOR U14447 ( .A(n14177), .B(n14176), .Z(n15009) );
  AND U14448 ( .A(n9141), .B(n9139), .Z(n15008) );
  XOR U14449 ( .A(n10359), .B(n15010), .Z(n9139) );
  XOR U14450 ( .A(n13588), .B(n15011), .Z(n10359) );
  XOR U14451 ( .A(n15012), .B(n15013), .Z(n13588) );
  XNOR U14452 ( .A(n12350), .B(n10250), .Z(n15013) );
  XOR U14453 ( .A(n15014), .B(n15015), .Z(n10250) );
  NOR U14454 ( .A(n15016), .B(n15017), .Z(n15014) );
  XOR U14455 ( .A(n15018), .B(n15019), .Z(n12350) );
  NOR U14456 ( .A(n15020), .B(n15021), .Z(n15018) );
  XOR U14457 ( .A(n10365), .B(n15022), .Z(n15012) );
  XNOR U14458 ( .A(n15023), .B(n15024), .Z(n15022) );
  XNOR U14459 ( .A(n15025), .B(n15026), .Z(n10365) );
  XNOR U14460 ( .A(n15029), .B(n9994), .Z(n9141) );
  XOR U14461 ( .A(n13367), .B(n15030), .Z(n9994) );
  XOR U14462 ( .A(n15031), .B(n15032), .Z(n13367) );
  XNOR U14463 ( .A(n10202), .B(n10826), .Z(n15032) );
  XOR U14464 ( .A(n15033), .B(n15034), .Z(n10826) );
  ANDN U14465 ( .B(n15035), .A(n15036), .Z(n15033) );
  XNOR U14466 ( .A(n15037), .B(n15038), .Z(n10202) );
  ANDN U14467 ( .B(n15039), .A(n13207), .Z(n15037) );
  XOR U14468 ( .A(n9912), .B(n15040), .Z(n15031) );
  XOR U14469 ( .A(n15041), .B(n11731), .Z(n15040) );
  XOR U14470 ( .A(n15042), .B(n15043), .Z(n11731) );
  NOR U14471 ( .A(n13217), .B(n15044), .Z(n15042) );
  XOR U14472 ( .A(n15045), .B(n15046), .Z(n9912) );
  NOR U14473 ( .A(n13213), .B(n15047), .Z(n15045) );
  XNOR U14474 ( .A(n15048), .B(n8006), .Z(n2343) );
  XOR U14475 ( .A(n13839), .B(n10050), .Z(n8006) );
  XNOR U14476 ( .A(n15049), .B(n15050), .Z(n13839) );
  AND U14477 ( .A(n15051), .B(n15052), .Z(n15049) );
  AND U14478 ( .A(n8005), .B(n9135), .Z(n15048) );
  XOR U14479 ( .A(n15053), .B(n13856), .Z(n9135) );
  XOR U14480 ( .A(n15054), .B(n12986), .Z(n13856) );
  XNOR U14481 ( .A(n15055), .B(n15056), .Z(n12986) );
  XNOR U14482 ( .A(n10024), .B(n12237), .Z(n15056) );
  XOR U14483 ( .A(n15057), .B(n15058), .Z(n12237) );
  AND U14484 ( .A(n15059), .B(n14236), .Z(n15057) );
  XNOR U14485 ( .A(n15060), .B(n15061), .Z(n10024) );
  ANDN U14486 ( .B(n15062), .A(n15063), .Z(n15060) );
  XNOR U14487 ( .A(n11973), .B(n15064), .Z(n15055) );
  XNOR U14488 ( .A(n11824), .B(n15065), .Z(n15064) );
  XOR U14489 ( .A(n15066), .B(n15067), .Z(n11824) );
  AND U14490 ( .A(n14242), .B(n15068), .Z(n15066) );
  XNOR U14491 ( .A(n15069), .B(n15070), .Z(n11973) );
  AND U14492 ( .A(n15071), .B(n14246), .Z(n15069) );
  XOR U14493 ( .A(n14630), .B(n9573), .Z(n8005) );
  XNOR U14494 ( .A(n15072), .B(n15073), .Z(n14630) );
  AND U14495 ( .A(n15074), .B(n14070), .Z(n15072) );
  IV U14496 ( .A(n15075), .Z(n14070) );
  XOR U14497 ( .A(n3160), .B(n15076), .Z(n15006) );
  XOR U14498 ( .A(n6312), .B(n7995), .Z(n15076) );
  XNOR U14499 ( .A(n15077), .B(n8011), .Z(n7995) );
  XNOR U14500 ( .A(n9191), .B(n15078), .Z(n8011) );
  XNOR U14501 ( .A(n14961), .B(n11989), .Z(n9191) );
  XOR U14502 ( .A(n15079), .B(n15080), .Z(n11989) );
  XNOR U14503 ( .A(n12332), .B(n13156), .Z(n15080) );
  XOR U14504 ( .A(n15081), .B(n15082), .Z(n13156) );
  ANDN U14505 ( .B(n14662), .A(n15083), .Z(n15081) );
  XNOR U14506 ( .A(n15084), .B(n15085), .Z(n12332) );
  AND U14507 ( .A(n15086), .B(n15087), .Z(n15084) );
  XOR U14508 ( .A(n11760), .B(n15088), .Z(n15079) );
  XOR U14509 ( .A(n14641), .B(n13197), .Z(n15088) );
  XNOR U14510 ( .A(n15089), .B(n14648), .Z(n13197) );
  ANDN U14511 ( .B(n15090), .A(n14647), .Z(n15089) );
  XOR U14512 ( .A(n15091), .B(n15092), .Z(n14641) );
  ANDN U14513 ( .B(n15093), .A(n14651), .Z(n15091) );
  XOR U14514 ( .A(n15094), .B(n14658), .Z(n11760) );
  ANDN U14515 ( .B(n15095), .A(n14657), .Z(n15094) );
  XOR U14516 ( .A(n15096), .B(n15097), .Z(n14961) );
  XNOR U14517 ( .A(n9387), .B(n12179), .Z(n15097) );
  XNOR U14518 ( .A(n15098), .B(n15099), .Z(n12179) );
  NOR U14519 ( .A(n15100), .B(n15101), .Z(n15098) );
  XNOR U14520 ( .A(n15102), .B(n15103), .Z(n9387) );
  NOR U14521 ( .A(n15104), .B(n15105), .Z(n15102) );
  XOR U14522 ( .A(n12867), .B(n15106), .Z(n15096) );
  XNOR U14523 ( .A(n15107), .B(n12040), .Z(n15106) );
  XOR U14524 ( .A(n15108), .B(n15109), .Z(n12040) );
  XOR U14525 ( .A(n15112), .B(n15113), .Z(n12867) );
  ANDN U14526 ( .B(n15114), .A(n15115), .Z(n15112) );
  ANDN U14527 ( .B(n9137), .A(n8010), .Z(n15077) );
  XNOR U14528 ( .A(n15116), .B(n10997), .Z(n8010) );
  XOR U14529 ( .A(n12945), .B(n15117), .Z(n10997) );
  XOR U14530 ( .A(n15118), .B(n15119), .Z(n12945) );
  XOR U14531 ( .A(n12767), .B(n12002), .Z(n15119) );
  XOR U14532 ( .A(n15120), .B(n12773), .Z(n12002) );
  XOR U14533 ( .A(n15121), .B(n15122), .Z(n12773) );
  ANDN U14534 ( .B(n15123), .A(n12772), .Z(n15120) );
  XNOR U14535 ( .A(n15124), .B(n14798), .Z(n12767) );
  ANDN U14536 ( .B(n14799), .A(n15125), .Z(n15124) );
  XNOR U14537 ( .A(n11664), .B(n15126), .Z(n15118) );
  XOR U14538 ( .A(n9109), .B(n11840), .Z(n15126) );
  XNOR U14539 ( .A(n15127), .B(n14889), .Z(n11840) );
  XOR U14540 ( .A(n15128), .B(n15129), .Z(n14889) );
  XOR U14541 ( .A(n15131), .B(n12776), .Z(n9109) );
  XNOR U14542 ( .A(n15132), .B(n15133), .Z(n12776) );
  ANDN U14543 ( .B(n12777), .A(n15134), .Z(n15131) );
  XOR U14544 ( .A(n15135), .B(n12783), .Z(n11664) );
  IV U14545 ( .A(n14893), .Z(n12783) );
  XOR U14546 ( .A(n15136), .B(n15137), .Z(n14893) );
  AND U14547 ( .A(n15138), .B(n12784), .Z(n15135) );
  XOR U14548 ( .A(n12455), .B(n15139), .Z(n9137) );
  XOR U14549 ( .A(n12597), .B(n15140), .Z(n12455) );
  XOR U14550 ( .A(n15141), .B(n15142), .Z(n12597) );
  XOR U14551 ( .A(n11858), .B(n11665), .Z(n15142) );
  XOR U14552 ( .A(n15143), .B(n15144), .Z(n11665) );
  ANDN U14553 ( .B(n15145), .A(n15146), .Z(n15143) );
  XNOR U14554 ( .A(n15147), .B(n14587), .Z(n11858) );
  IV U14555 ( .A(n15148), .Z(n14587) );
  NOR U14556 ( .A(n15149), .B(n15150), .Z(n15147) );
  XNOR U14557 ( .A(n11997), .B(n15151), .Z(n15141) );
  XOR U14558 ( .A(n15152), .B(n15153), .Z(n15151) );
  XNOR U14559 ( .A(n15154), .B(n14574), .Z(n11997) );
  AND U14560 ( .A(n15155), .B(n15156), .Z(n15154) );
  XNOR U14561 ( .A(n15157), .B(n8015), .Z(n6312) );
  XNOR U14562 ( .A(n15158), .B(n12662), .Z(n8015) );
  AND U14563 ( .A(n14435), .B(n15159), .Z(n15157) );
  XOR U14564 ( .A(n15160), .B(n8018), .Z(n3160) );
  XNOR U14565 ( .A(n15161), .B(n10995), .Z(n8018) );
  XNOR U14566 ( .A(n14325), .B(n13226), .Z(n10995) );
  XNOR U14567 ( .A(n15162), .B(n15163), .Z(n13226) );
  XNOR U14568 ( .A(n12764), .B(n10558), .Z(n15163) );
  XOR U14569 ( .A(n15164), .B(n13782), .Z(n10558) );
  ANDN U14570 ( .B(n15165), .A(n15166), .Z(n15164) );
  XNOR U14571 ( .A(n15167), .B(n15168), .Z(n12764) );
  ANDN U14572 ( .B(n15169), .A(n15170), .Z(n15167) );
  XNOR U14573 ( .A(n10663), .B(n15171), .Z(n15162) );
  XOR U14574 ( .A(n12565), .B(n12535), .Z(n15171) );
  XNOR U14575 ( .A(n15172), .B(n13785), .Z(n12535) );
  ANDN U14576 ( .B(n15173), .A(n15174), .Z(n15172) );
  XOR U14577 ( .A(n15175), .B(n13776), .Z(n12565) );
  XNOR U14578 ( .A(n15178), .B(n13771), .Z(n10663) );
  ANDN U14579 ( .B(n15179), .A(n15180), .Z(n15178) );
  XOR U14580 ( .A(n15181), .B(n15182), .Z(n14325) );
  XNOR U14581 ( .A(n15183), .B(n10060), .Z(n15182) );
  XNOR U14582 ( .A(n15184), .B(n13800), .Z(n10060) );
  ANDN U14583 ( .B(n15185), .A(n15186), .Z(n15184) );
  XOR U14584 ( .A(n12146), .B(n15187), .Z(n15181) );
  XNOR U14585 ( .A(n11053), .B(n12134), .Z(n15187) );
  XNOR U14586 ( .A(n15188), .B(n13808), .Z(n12134) );
  AND U14587 ( .A(n15189), .B(n15190), .Z(n15188) );
  XOR U14588 ( .A(n15191), .B(n13805), .Z(n11053) );
  NOR U14589 ( .A(n15192), .B(n15193), .Z(n15191) );
  XOR U14590 ( .A(n15194), .B(n13791), .Z(n12146) );
  AND U14591 ( .A(n15195), .B(n15196), .Z(n15194) );
  AND U14592 ( .A(n9132), .B(n8019), .Z(n15160) );
  XOR U14593 ( .A(n15197), .B(n9067), .Z(n8019) );
  IV U14594 ( .A(n9274), .Z(n9067) );
  XOR U14595 ( .A(n14467), .B(n15198), .Z(n9274) );
  XOR U14596 ( .A(n15199), .B(n15200), .Z(n14467) );
  XOR U14597 ( .A(n10787), .B(n12717), .Z(n15200) );
  XNOR U14598 ( .A(n15201), .B(n15202), .Z(n12717) );
  NOR U14599 ( .A(n13097), .B(n13098), .Z(n15201) );
  XNOR U14600 ( .A(n15203), .B(n15204), .Z(n13098) );
  XOR U14601 ( .A(n15205), .B(n15206), .Z(n10787) );
  ANDN U14602 ( .B(n13105), .A(n13106), .Z(n15205) );
  XOR U14603 ( .A(n13599), .B(n15209), .Z(n15199) );
  XNOR U14604 ( .A(n11196), .B(n11536), .Z(n15209) );
  XOR U14605 ( .A(n15210), .B(n15211), .Z(n11536) );
  ANDN U14606 ( .B(n13092), .A(n13093), .Z(n15210) );
  XNOR U14607 ( .A(n15212), .B(n15213), .Z(n13093) );
  XNOR U14608 ( .A(n15214), .B(n15215), .Z(n11196) );
  AND U14609 ( .A(n13925), .B(n14466), .Z(n15214) );
  XOR U14610 ( .A(n15216), .B(n15217), .Z(n13925) );
  XOR U14611 ( .A(n15218), .B(n15219), .Z(n13599) );
  ANDN U14612 ( .B(n15220), .A(n13102), .Z(n15218) );
  XOR U14613 ( .A(n15221), .B(n15222), .Z(n13102) );
  XNOR U14614 ( .A(n15223), .B(n15224), .Z(n9132) );
  XOR U14615 ( .A(n15225), .B(n15226), .Z(n10085) );
  XNOR U14616 ( .A(n5062), .B(n1948), .Z(n15226) );
  XNOR U14617 ( .A(n15227), .B(n7931), .Z(n1948) );
  XNOR U14618 ( .A(n12304), .B(n10473), .Z(n7931) );
  XNOR U14619 ( .A(n15228), .B(n15229), .Z(n12304) );
  ANDN U14620 ( .B(n9158), .A(n9157), .Z(n15227) );
  XNOR U14621 ( .A(n13486), .B(n10712), .Z(n9157) );
  XNOR U14622 ( .A(n15232), .B(n14166), .Z(n13486) );
  ANDN U14623 ( .B(n14712), .A(n15233), .Z(n15232) );
  XNOR U14624 ( .A(n15234), .B(n12050), .Z(n9158) );
  XNOR U14625 ( .A(n15235), .B(n8067), .Z(n5062) );
  XOR U14626 ( .A(n9558), .B(n15236), .Z(n8067) );
  XOR U14627 ( .A(n12796), .B(n12999), .Z(n9558) );
  XNOR U14628 ( .A(n15237), .B(n15238), .Z(n12999) );
  XNOR U14629 ( .A(n12561), .B(n12741), .Z(n15238) );
  XOR U14630 ( .A(n15239), .B(n12755), .Z(n12741) );
  IV U14631 ( .A(n13460), .Z(n12755) );
  XOR U14632 ( .A(n15240), .B(n15217), .Z(n13460) );
  NOR U14633 ( .A(n12754), .B(n15241), .Z(n15239) );
  XNOR U14634 ( .A(n15242), .B(n13451), .Z(n12561) );
  IV U14635 ( .A(n13464), .Z(n13451) );
  XOR U14636 ( .A(n15243), .B(n15244), .Z(n13464) );
  AND U14637 ( .A(n13465), .B(n15245), .Z(n15242) );
  XNOR U14638 ( .A(n12527), .B(n15246), .Z(n15237) );
  XOR U14639 ( .A(n12057), .B(n11279), .Z(n15246) );
  XOR U14640 ( .A(n15247), .B(n12971), .Z(n11279) );
  XNOR U14641 ( .A(n15248), .B(n15249), .Z(n12971) );
  XNOR U14642 ( .A(n15251), .B(n12749), .Z(n12057) );
  XNOR U14643 ( .A(n15252), .B(n15253), .Z(n12749) );
  NOR U14644 ( .A(n12748), .B(n15254), .Z(n15251) );
  XNOR U14645 ( .A(n15255), .B(n12758), .Z(n12527) );
  XNOR U14646 ( .A(n15256), .B(n15257), .Z(n12758) );
  AND U14647 ( .A(n15258), .B(n12759), .Z(n15255) );
  XOR U14648 ( .A(n15259), .B(n15260), .Z(n12796) );
  XNOR U14649 ( .A(n10647), .B(n11984), .Z(n15260) );
  XNOR U14650 ( .A(n15261), .B(n15262), .Z(n11984) );
  AND U14651 ( .A(n15263), .B(n15264), .Z(n15261) );
  XOR U14652 ( .A(n15265), .B(n15266), .Z(n10647) );
  AND U14653 ( .A(n15267), .B(n15268), .Z(n15265) );
  XNOR U14654 ( .A(n12160), .B(n15269), .Z(n15259) );
  XOR U14655 ( .A(n9487), .B(n9355), .Z(n15269) );
  XOR U14656 ( .A(n15270), .B(n15271), .Z(n9355) );
  AND U14657 ( .A(n15272), .B(n15273), .Z(n15270) );
  XOR U14658 ( .A(n15274), .B(n15275), .Z(n9487) );
  NOR U14659 ( .A(n15276), .B(n15277), .Z(n15274) );
  XOR U14660 ( .A(n15278), .B(n15279), .Z(n12160) );
  ANDN U14661 ( .B(n15280), .A(n15281), .Z(n15278) );
  AND U14662 ( .A(n9153), .B(n9997), .Z(n15235) );
  XOR U14663 ( .A(n15282), .B(n13421), .Z(n9997) );
  XOR U14664 ( .A(n12891), .B(n14778), .Z(n13421) );
  XNOR U14665 ( .A(n15283), .B(n15284), .Z(n14778) );
  XNOR U14666 ( .A(n9569), .B(n14403), .Z(n15284) );
  XNOR U14667 ( .A(n15285), .B(n15286), .Z(n14403) );
  ANDN U14668 ( .B(n15287), .A(n14389), .Z(n15285) );
  XNOR U14669 ( .A(n15288), .B(n15289), .Z(n9569) );
  AND U14670 ( .A(n15290), .B(n14382), .Z(n15288) );
  XNOR U14671 ( .A(n9379), .B(n15291), .Z(n15283) );
  XOR U14672 ( .A(n10893), .B(n10221), .Z(n15291) );
  XOR U14673 ( .A(n15292), .B(n15293), .Z(n10221) );
  AND U14674 ( .A(n14386), .B(n15294), .Z(n15292) );
  XNOR U14675 ( .A(n15295), .B(n15296), .Z(n10893) );
  ANDN U14676 ( .B(n15297), .A(n14377), .Z(n15295) );
  XNOR U14677 ( .A(n15298), .B(n15299), .Z(n9379) );
  AND U14678 ( .A(n14373), .B(n15300), .Z(n15298) );
  XOR U14679 ( .A(n15301), .B(n15302), .Z(n12891) );
  XNOR U14680 ( .A(n12626), .B(n11403), .Z(n15302) );
  XOR U14681 ( .A(n15303), .B(n14413), .Z(n11403) );
  AND U14682 ( .A(n15304), .B(n14414), .Z(n15303) );
  XNOR U14683 ( .A(n15305), .B(n14419), .Z(n12626) );
  AND U14684 ( .A(n15306), .B(n15307), .Z(n15305) );
  XNOR U14685 ( .A(n12184), .B(n15308), .Z(n15301) );
  XOR U14686 ( .A(n11323), .B(n13908), .Z(n15308) );
  XNOR U14687 ( .A(n15309), .B(n14410), .Z(n13908) );
  AND U14688 ( .A(n14409), .B(n15310), .Z(n15309) );
  XNOR U14689 ( .A(n15311), .B(n14423), .Z(n11323) );
  ANDN U14690 ( .B(n14422), .A(n15312), .Z(n15311) );
  XNOR U14691 ( .A(n15313), .B(n14427), .Z(n12184) );
  NOR U14692 ( .A(n15314), .B(n14426), .Z(n15313) );
  XNOR U14693 ( .A(n9101), .B(n15315), .Z(n9153) );
  XNOR U14694 ( .A(n15316), .B(n13964), .Z(n9101) );
  XOR U14695 ( .A(n15317), .B(n15318), .Z(n13964) );
  XNOR U14696 ( .A(n12691), .B(n11047), .Z(n15318) );
  XOR U14697 ( .A(n15319), .B(n13897), .Z(n11047) );
  IV U14698 ( .A(n15320), .Z(n13897) );
  ANDN U14699 ( .B(n13871), .A(n13346), .Z(n15319) );
  XOR U14700 ( .A(n15321), .B(n15322), .Z(n13346) );
  XOR U14701 ( .A(n15323), .B(n13888), .Z(n12691) );
  ANDN U14702 ( .B(n13875), .A(n13354), .Z(n15323) );
  XOR U14703 ( .A(n15324), .B(n15325), .Z(n13354) );
  XOR U14704 ( .A(n9658), .B(n15326), .Z(n15317) );
  XOR U14705 ( .A(n10164), .B(n14933), .Z(n15326) );
  XNOR U14706 ( .A(n15327), .B(n13893), .Z(n14933) );
  AND U14707 ( .A(n13341), .B(n13868), .Z(n15327) );
  IV U14708 ( .A(n15328), .Z(n13868) );
  XOR U14709 ( .A(n15329), .B(n15330), .Z(n13341) );
  XNOR U14710 ( .A(n15331), .B(n13884), .Z(n10164) );
  AND U14711 ( .A(n13873), .B(n13350), .Z(n15331) );
  XOR U14712 ( .A(n15332), .B(n15333), .Z(n13350) );
  XNOR U14713 ( .A(n15334), .B(n13899), .Z(n9658) );
  NOR U14714 ( .A(n13337), .B(n13989), .Z(n15334) );
  XNOR U14715 ( .A(n15335), .B(n15336), .Z(n13337) );
  XNOR U14716 ( .A(n3703), .B(n15337), .Z(n15225) );
  XNOR U14717 ( .A(n9227), .B(n4172), .Z(n15337) );
  XNOR U14718 ( .A(n15338), .B(n7941), .Z(n4172) );
  XOR U14719 ( .A(n10094), .B(n15339), .Z(n7941) );
  NOR U14720 ( .A(n9234), .B(n9987), .Z(n15338) );
  XOR U14721 ( .A(n9513), .B(n15340), .Z(n9987) );
  XOR U14722 ( .A(n14999), .B(n12667), .Z(n9513) );
  XNOR U14723 ( .A(n15341), .B(n15342), .Z(n12667) );
  XNOR U14724 ( .A(n14930), .B(n14544), .Z(n15342) );
  XOR U14725 ( .A(n15343), .B(n15314), .Z(n14544) );
  ANDN U14726 ( .B(n15344), .A(n14425), .Z(n15343) );
  XNOR U14727 ( .A(n15345), .B(n15310), .Z(n14930) );
  ANDN U14728 ( .B(n15346), .A(n14408), .Z(n15345) );
  XNOR U14729 ( .A(n11054), .B(n15347), .Z(n15341) );
  XOR U14730 ( .A(n15348), .B(n11978), .Z(n15347) );
  XOR U14731 ( .A(n15349), .B(n15312), .Z(n11978) );
  AND U14732 ( .A(n15350), .B(n14421), .Z(n15349) );
  IV U14733 ( .A(n15351), .Z(n14421) );
  XNOR U14734 ( .A(n15352), .B(n15306), .Z(n11054) );
  AND U14735 ( .A(n14417), .B(n15353), .Z(n15352) );
  XOR U14736 ( .A(n15354), .B(n15355), .Z(n14999) );
  XOR U14737 ( .A(n12320), .B(n10372), .Z(n15355) );
  XNOR U14738 ( .A(n15356), .B(n15357), .Z(n10372) );
  AND U14739 ( .A(n15002), .B(n15358), .Z(n15356) );
  XNOR U14740 ( .A(n15359), .B(n12903), .Z(n12320) );
  AND U14741 ( .A(n15360), .B(n14109), .Z(n15359) );
  XNOR U14742 ( .A(n11271), .B(n15361), .Z(n15354) );
  XNOR U14743 ( .A(n14665), .B(n11925), .Z(n15361) );
  XOR U14744 ( .A(n15362), .B(n12900), .Z(n11925) );
  ANDN U14745 ( .B(n14112), .A(n14113), .Z(n15362) );
  XNOR U14746 ( .A(n15363), .B(n12908), .Z(n14665) );
  AND U14747 ( .A(n14117), .B(n15364), .Z(n15363) );
  XNOR U14748 ( .A(n15365), .B(n15366), .Z(n11271) );
  AND U14749 ( .A(n14120), .B(n15367), .Z(n15365) );
  XOR U14750 ( .A(n15368), .B(n10714), .Z(n9234) );
  XOR U14751 ( .A(n15369), .B(n13386), .Z(n10714) );
  XNOR U14752 ( .A(n15370), .B(n15371), .Z(n13386) );
  XNOR U14753 ( .A(n12798), .B(n12408), .Z(n15371) );
  XOR U14754 ( .A(n15372), .B(n14048), .Z(n12408) );
  ANDN U14755 ( .B(n15373), .A(n15374), .Z(n15372) );
  XOR U14756 ( .A(n15375), .B(n15376), .Z(n12798) );
  ANDN U14757 ( .B(n15377), .A(n15378), .Z(n15375) );
  XOR U14758 ( .A(n11314), .B(n15379), .Z(n15370) );
  XOR U14759 ( .A(n12842), .B(n12470), .Z(n15379) );
  XNOR U14760 ( .A(n15380), .B(n14037), .Z(n12470) );
  AND U14761 ( .A(n15381), .B(n15382), .Z(n15380) );
  XNOR U14762 ( .A(n15383), .B(n14044), .Z(n12842) );
  AND U14763 ( .A(n15384), .B(n15385), .Z(n15383) );
  XOR U14764 ( .A(n15386), .B(n15387), .Z(n11314) );
  NOR U14765 ( .A(n15388), .B(n15389), .Z(n15386) );
  XOR U14766 ( .A(n15390), .B(n7937), .Z(n9227) );
  XOR U14767 ( .A(n15391), .B(n12210), .Z(n7937) );
  IV U14768 ( .A(n13075), .Z(n12210) );
  XNOR U14769 ( .A(n15392), .B(n15393), .Z(n13075) );
  NOR U14770 ( .A(n9146), .B(n9147), .Z(n15390) );
  XOR U14771 ( .A(n14447), .B(n10590), .Z(n9147) );
  XOR U14772 ( .A(n11803), .B(n14471), .Z(n10590) );
  XOR U14773 ( .A(n15394), .B(n15395), .Z(n14471) );
  XNOR U14774 ( .A(n12049), .B(n15396), .Z(n15395) );
  XNOR U14775 ( .A(n15397), .B(n14214), .Z(n12049) );
  ANDN U14776 ( .B(n15398), .A(n15399), .Z(n15397) );
  XOR U14777 ( .A(n13936), .B(n15400), .Z(n15394) );
  XOR U14778 ( .A(n14128), .B(n15234), .Z(n15400) );
  XNOR U14779 ( .A(n15401), .B(n14203), .Z(n15234) );
  AND U14780 ( .A(n13946), .B(n15402), .Z(n15401) );
  XNOR U14781 ( .A(n15403), .B(n14210), .Z(n14128) );
  ANDN U14782 ( .B(n13955), .A(n15404), .Z(n15403) );
  IV U14783 ( .A(n15405), .Z(n13955) );
  XNOR U14784 ( .A(n15406), .B(n14200), .Z(n13936) );
  ANDN U14785 ( .B(n15407), .A(n13951), .Z(n15406) );
  XOR U14786 ( .A(n15408), .B(n15409), .Z(n11803) );
  XOR U14787 ( .A(n15410), .B(n9581), .Z(n15409) );
  XOR U14788 ( .A(n15411), .B(n13678), .Z(n9581) );
  ANDN U14789 ( .B(n15412), .A(n15413), .Z(n15411) );
  XOR U14790 ( .A(n12640), .B(n15414), .Z(n15408) );
  XOR U14791 ( .A(n12192), .B(n11034), .Z(n15414) );
  XOR U14792 ( .A(n15415), .B(n13665), .Z(n11034) );
  IV U14793 ( .A(n15416), .Z(n13665) );
  NOR U14794 ( .A(n14457), .B(n14456), .Z(n15415) );
  XNOR U14795 ( .A(n15417), .B(n13675), .Z(n12192) );
  NOR U14796 ( .A(n14454), .B(n14453), .Z(n15417) );
  ANDN U14797 ( .B(n14460), .A(n14459), .Z(n15418) );
  XNOR U14798 ( .A(n15419), .B(n15413), .Z(n14447) );
  XNOR U14799 ( .A(n10898), .B(n14570), .Z(n9146) );
  XNOR U14800 ( .A(n15420), .B(n15421), .Z(n14570) );
  AND U14801 ( .A(n15422), .B(n15144), .Z(n15420) );
  IV U14802 ( .A(n15423), .Z(n15144) );
  XNOR U14803 ( .A(n12161), .B(n14281), .Z(n10898) );
  XNOR U14804 ( .A(n15424), .B(n15425), .Z(n14281) );
  XNOR U14805 ( .A(n15426), .B(n12343), .Z(n15425) );
  XOR U14806 ( .A(n15427), .B(n15428), .Z(n12343) );
  NOR U14807 ( .A(n14581), .B(n14582), .Z(n15427) );
  XNOR U14808 ( .A(n11020), .B(n15429), .Z(n15424) );
  XNOR U14809 ( .A(n11577), .B(n15430), .Z(n15429) );
  XNOR U14810 ( .A(n15431), .B(n15150), .Z(n11577) );
  ANDN U14811 ( .B(n14585), .A(n14586), .Z(n15431) );
  XNOR U14812 ( .A(n15432), .B(n15155), .Z(n11020) );
  NOR U14813 ( .A(n14572), .B(n14573), .Z(n15432) );
  XOR U14814 ( .A(n15433), .B(n15434), .Z(n12161) );
  XOR U14815 ( .A(n12321), .B(n10276), .Z(n15434) );
  XOR U14816 ( .A(n15435), .B(n15436), .Z(n10276) );
  AND U14817 ( .A(n15275), .B(n15277), .Z(n15435) );
  XNOR U14818 ( .A(n15437), .B(n15438), .Z(n12321) );
  ANDN U14819 ( .B(n15279), .A(n15280), .Z(n15437) );
  XOR U14820 ( .A(n11499), .B(n15439), .Z(n15433) );
  XNOR U14821 ( .A(n13080), .B(n9823), .Z(n15439) );
  XNOR U14822 ( .A(n15440), .B(n15441), .Z(n9823) );
  ANDN U14823 ( .B(n15271), .A(n15272), .Z(n15440) );
  XNOR U14824 ( .A(n15442), .B(n15443), .Z(n13080) );
  NOR U14825 ( .A(n15262), .B(n15264), .Z(n15442) );
  XNOR U14826 ( .A(n15444), .B(n15445), .Z(n11499) );
  ANDN U14827 ( .B(n15266), .A(n15268), .Z(n15444) );
  XOR U14828 ( .A(n15446), .B(n7927), .Z(n3703) );
  XNOR U14829 ( .A(n14145), .B(n9768), .Z(n7927) );
  XNOR U14830 ( .A(n15447), .B(n15448), .Z(n14145) );
  ANDN U14831 ( .B(n15449), .A(n15450), .Z(n15447) );
  ANDN U14832 ( .B(n9151), .A(n9150), .Z(n15446) );
  XNOR U14833 ( .A(n15451), .B(n10235), .Z(n9150) );
  XNOR U14834 ( .A(n11524), .B(n12863), .Z(n10235) );
  XNOR U14835 ( .A(n15452), .B(n15453), .Z(n12863) );
  XNOR U14836 ( .A(n10360), .B(n14952), .Z(n15453) );
  XNOR U14837 ( .A(n15454), .B(n14490), .Z(n14952) );
  AND U14838 ( .A(n15455), .B(n15456), .Z(n15454) );
  XOR U14839 ( .A(n15457), .B(n14477), .Z(n10360) );
  AND U14840 ( .A(n15458), .B(n15459), .Z(n15457) );
  XNOR U14841 ( .A(n12642), .B(n15460), .Z(n15452) );
  XOR U14842 ( .A(n10818), .B(n15010), .Z(n15460) );
  XNOR U14843 ( .A(n15461), .B(n14481), .Z(n15010) );
  AND U14844 ( .A(n15462), .B(n15463), .Z(n15461) );
  XOR U14845 ( .A(n15464), .B(n14486), .Z(n10818) );
  AND U14846 ( .A(n15465), .B(n15466), .Z(n15464) );
  XOR U14847 ( .A(n15467), .B(n15468), .Z(n12642) );
  AND U14848 ( .A(n15469), .B(n15470), .Z(n15467) );
  XOR U14849 ( .A(n15471), .B(n15472), .Z(n11524) );
  XNOR U14850 ( .A(n13587), .B(n11454), .Z(n15472) );
  XNOR U14851 ( .A(n15473), .B(n15474), .Z(n11454) );
  AND U14852 ( .A(n15475), .B(n15476), .Z(n15473) );
  XNOR U14853 ( .A(n15477), .B(n15478), .Z(n13587) );
  NOR U14854 ( .A(n15479), .B(n15480), .Z(n15477) );
  XOR U14855 ( .A(n11831), .B(n15481), .Z(n15471) );
  XOR U14856 ( .A(n12552), .B(n10923), .Z(n15481) );
  XOR U14857 ( .A(n15482), .B(n15017), .Z(n10923) );
  ANDN U14858 ( .B(n15016), .A(n15483), .Z(n15482) );
  XNOR U14859 ( .A(n15484), .B(n15020), .Z(n12552) );
  ANDN U14860 ( .B(n15021), .A(n15485), .Z(n15484) );
  XOR U14861 ( .A(n15486), .B(n15028), .Z(n11831) );
  NOR U14862 ( .A(n15487), .B(n15027), .Z(n15486) );
  XOR U14863 ( .A(n15488), .B(n12191), .Z(n9151) );
  XNOR U14864 ( .A(n12541), .B(n14031), .Z(n12191) );
  XNOR U14865 ( .A(n15489), .B(n15490), .Z(n14031) );
  XNOR U14866 ( .A(n13083), .B(n12682), .Z(n15490) );
  XOR U14867 ( .A(n15491), .B(n15492), .Z(n12682) );
  ANDN U14868 ( .B(n15493), .A(n15494), .Z(n15491) );
  XNOR U14869 ( .A(n15495), .B(n15496), .Z(n13083) );
  XOR U14870 ( .A(n11455), .B(n15499), .Z(n15489) );
  XOR U14871 ( .A(n13157), .B(n12723), .Z(n15499) );
  XOR U14872 ( .A(n15500), .B(n15501), .Z(n12723) );
  ANDN U14873 ( .B(n15502), .A(n15503), .Z(n15500) );
  XNOR U14874 ( .A(n15504), .B(n15505), .Z(n13157) );
  NOR U14875 ( .A(n15506), .B(n15507), .Z(n15504) );
  XOR U14876 ( .A(n15508), .B(n15509), .Z(n11455) );
  NOR U14877 ( .A(n15510), .B(n15511), .Z(n15508) );
  XOR U14878 ( .A(n15512), .B(n15513), .Z(n12541) );
  XNOR U14879 ( .A(n10129), .B(n9793), .Z(n15513) );
  XOR U14880 ( .A(n15514), .B(n14620), .Z(n9793) );
  IV U14881 ( .A(n13327), .Z(n14620) );
  XOR U14882 ( .A(n15515), .B(n15516), .Z(n13327) );
  NOR U14883 ( .A(n15517), .B(n13326), .Z(n15514) );
  XOR U14884 ( .A(n15518), .B(n13174), .Z(n10129) );
  XNOR U14885 ( .A(n15519), .B(n15520), .Z(n13174) );
  XOR U14886 ( .A(n10989), .B(n15522), .Z(n15512) );
  XOR U14887 ( .A(n9397), .B(n11801), .Z(n15522) );
  XOR U14888 ( .A(n15523), .B(n13178), .Z(n11801) );
  XNOR U14889 ( .A(n15524), .B(n15525), .Z(n13178) );
  NOR U14890 ( .A(n13177), .B(n15526), .Z(n15523) );
  XOR U14891 ( .A(n15527), .B(n14611), .Z(n9397) );
  IV U14892 ( .A(n13170), .Z(n14611) );
  XNOR U14893 ( .A(n15528), .B(n15529), .Z(n13170) );
  NOR U14894 ( .A(n15530), .B(n13169), .Z(n15527) );
  XOR U14895 ( .A(n15531), .B(n14617), .Z(n10989) );
  IV U14896 ( .A(n13165), .Z(n14617) );
  XOR U14897 ( .A(n15532), .B(n15533), .Z(n13165) );
  NOR U14898 ( .A(n15534), .B(n13164), .Z(n15531) );
  XOR U14899 ( .A(n15535), .B(n8014), .Z(n9130) );
  IV U14900 ( .A(n15159), .Z(n8014) );
  XOR U14901 ( .A(n15536), .B(n11522), .Z(n15159) );
  NOR U14902 ( .A(n14435), .B(n9056), .Z(n15535) );
  XOR U14903 ( .A(n15396), .B(n12050), .Z(n9056) );
  XNOR U14904 ( .A(n15537), .B(n15538), .Z(n12050) );
  XOR U14905 ( .A(n15539), .B(n15540), .Z(n15396) );
  NOR U14906 ( .A(n13959), .B(n15541), .Z(n15539) );
  XNOR U14907 ( .A(n15542), .B(n9661), .Z(n14435) );
  NOR U14908 ( .A(n5661), .B(n5660), .Z(n15005) );
  XOR U14909 ( .A(n8959), .B(n5148), .Z(n5660) );
  XNOR U14910 ( .A(n15543), .B(n15544), .Z(n6494) );
  XNOR U14911 ( .A(n6306), .B(n2536), .Z(n15544) );
  XNOR U14912 ( .A(n15545), .B(n6525), .Z(n2536) );
  XNOR U14913 ( .A(n15546), .B(n9213), .Z(n6525) );
  XOR U14914 ( .A(n13373), .B(n11533), .Z(n9213) );
  XOR U14915 ( .A(n15547), .B(n15548), .Z(n11533) );
  XOR U14916 ( .A(n13397), .B(n12618), .Z(n15548) );
  XNOR U14917 ( .A(n15549), .B(n15550), .Z(n12618) );
  AND U14918 ( .A(n15551), .B(n15552), .Z(n15549) );
  XNOR U14919 ( .A(n15553), .B(n15554), .Z(n13397) );
  ANDN U14920 ( .B(n15555), .A(n15556), .Z(n15553) );
  XNOR U14921 ( .A(n12638), .B(n15557), .Z(n15547) );
  XOR U14922 ( .A(n10911), .B(n12004), .Z(n15557) );
  XOR U14923 ( .A(n15558), .B(n15559), .Z(n12004) );
  ANDN U14924 ( .B(n15560), .A(n14763), .Z(n15558) );
  XOR U14925 ( .A(n15561), .B(n15562), .Z(n10911) );
  XNOR U14926 ( .A(n15564), .B(n15565), .Z(n12638) );
  ANDN U14927 ( .B(n15566), .A(n14774), .Z(n15564) );
  XOR U14928 ( .A(n15567), .B(n15568), .Z(n13373) );
  XNOR U14929 ( .A(n9209), .B(n11878), .Z(n15568) );
  XNOR U14930 ( .A(n15569), .B(n14255), .Z(n11878) );
  AND U14931 ( .A(n14100), .B(n15570), .Z(n15569) );
  XNOR U14932 ( .A(n15571), .B(n15572), .Z(n9209) );
  AND U14933 ( .A(n15573), .B(n14093), .Z(n15571) );
  XOR U14934 ( .A(n11558), .B(n15574), .Z(n15567) );
  XOR U14935 ( .A(n12557), .B(n9217), .Z(n15574) );
  XOR U14936 ( .A(n15575), .B(n13410), .Z(n9217) );
  AND U14937 ( .A(n14089), .B(n15576), .Z(n15575) );
  XOR U14938 ( .A(n15577), .B(n13407), .Z(n12557) );
  IV U14939 ( .A(n15578), .Z(n13407) );
  ANDN U14940 ( .B(n14097), .A(n13406), .Z(n15577) );
  XNOR U14941 ( .A(n15579), .B(n13414), .Z(n11558) );
  AND U14942 ( .A(n13415), .B(n14085), .Z(n15579) );
  NOR U14943 ( .A(n8965), .B(n8964), .Z(n15545) );
  XOR U14944 ( .A(n10100), .B(n15580), .Z(n8964) );
  XOR U14945 ( .A(n15581), .B(n11656), .Z(n8965) );
  XNOR U14946 ( .A(n15582), .B(n14105), .Z(n11656) );
  XNOR U14947 ( .A(n15583), .B(n15584), .Z(n14105) );
  XNOR U14948 ( .A(n10432), .B(n11000), .Z(n15584) );
  XNOR U14949 ( .A(n15585), .B(n15350), .Z(n11000) );
  AND U14950 ( .A(n14423), .B(n15351), .Z(n15585) );
  XNOR U14951 ( .A(n15586), .B(n15529), .Z(n15351) );
  XOR U14952 ( .A(n15587), .B(n15588), .Z(n14423) );
  XNOR U14953 ( .A(n15589), .B(n15353), .Z(n10432) );
  ANDN U14954 ( .B(n14419), .A(n14417), .Z(n15589) );
  XNOR U14955 ( .A(n15592), .B(n15593), .Z(n14419) );
  XOR U14956 ( .A(n15340), .B(n15594), .Z(n15583) );
  XNOR U14957 ( .A(n9514), .B(n9680), .Z(n15594) );
  XNOR U14958 ( .A(n15595), .B(n15344), .Z(n9680) );
  AND U14959 ( .A(n14425), .B(n14427), .Z(n15595) );
  XOR U14960 ( .A(n15596), .B(n15597), .Z(n14427) );
  XNOR U14961 ( .A(n15598), .B(n15599), .Z(n14425) );
  XNOR U14962 ( .A(n15600), .B(n15601), .Z(n9514) );
  ANDN U14963 ( .B(n14412), .A(n14413), .Z(n15600) );
  XNOR U14964 ( .A(n15602), .B(n15603), .Z(n14413) );
  XNOR U14965 ( .A(n15604), .B(n15346), .Z(n15340) );
  AND U14966 ( .A(n14408), .B(n14410), .Z(n15604) );
  XNOR U14967 ( .A(n15605), .B(n15606), .Z(n14410) );
  XNOR U14968 ( .A(n15607), .B(n15608), .Z(n14408) );
  XOR U14969 ( .A(n15609), .B(n6530), .Z(n6306) );
  IV U14970 ( .A(n9013), .Z(n6530) );
  XOR U14971 ( .A(n14261), .B(n10431), .Z(n9013) );
  XNOR U14972 ( .A(n12835), .B(n11751), .Z(n10431) );
  XNOR U14973 ( .A(n15610), .B(n15611), .Z(n11751) );
  XOR U14974 ( .A(n15116), .B(n10996), .Z(n15611) );
  XOR U14975 ( .A(n15612), .B(n15613), .Z(n10996) );
  AND U14976 ( .A(n14263), .B(n14265), .Z(n15612) );
  XOR U14977 ( .A(n15614), .B(n15615), .Z(n14265) );
  XNOR U14978 ( .A(n15616), .B(n15617), .Z(n15116) );
  XOR U14979 ( .A(n13853), .B(n15619), .Z(n15610) );
  XNOR U14980 ( .A(n13685), .B(n11768), .Z(n15619) );
  XNOR U14981 ( .A(n15620), .B(n15621), .Z(n11768) );
  NOR U14982 ( .A(n14268), .B(n14269), .Z(n15620) );
  XOR U14983 ( .A(n15622), .B(n15623), .Z(n14269) );
  XNOR U14984 ( .A(n15624), .B(n15625), .Z(n13685) );
  XNOR U14985 ( .A(n15626), .B(n15627), .Z(n14273) );
  XNOR U14986 ( .A(n15628), .B(n15629), .Z(n13853) );
  AND U14987 ( .A(n14276), .B(n14818), .Z(n15628) );
  IV U14988 ( .A(n14277), .Z(n14818) );
  XOR U14989 ( .A(n15630), .B(n15631), .Z(n14277) );
  XOR U14990 ( .A(n15632), .B(n15633), .Z(n12835) );
  XOR U14991 ( .A(n12944), .B(n11561), .Z(n15633) );
  XOR U14992 ( .A(n15634), .B(n14799), .Z(n11561) );
  XOR U14993 ( .A(n15598), .B(n15635), .Z(n14799) );
  ANDN U14994 ( .B(n15125), .A(n15636), .Z(n15634) );
  XOR U14995 ( .A(n15637), .B(n12772), .Z(n12944) );
  XOR U14996 ( .A(n15638), .B(n15639), .Z(n12772) );
  IV U14997 ( .A(n15640), .Z(n14897) );
  XOR U14998 ( .A(n12930), .B(n15641), .Z(n15632) );
  XOR U14999 ( .A(n11048), .B(n10598), .Z(n15641) );
  XNOR U15000 ( .A(n15642), .B(n12784), .Z(n10598) );
  XOR U15001 ( .A(n15643), .B(n15644), .Z(n12784) );
  NOR U15002 ( .A(n15645), .B(n15138), .Z(n15642) );
  XNOR U15003 ( .A(n15646), .B(n12777), .Z(n11048) );
  XOR U15004 ( .A(n15647), .B(n15648), .Z(n12777) );
  AND U15005 ( .A(n14899), .B(n15134), .Z(n15646) );
  XNOR U15006 ( .A(n15649), .B(n14927), .Z(n12930) );
  XNOR U15007 ( .A(n15650), .B(n15651), .Z(n14927) );
  ANDN U15008 ( .B(n15130), .A(n14888), .Z(n15649) );
  XNOR U15009 ( .A(n15652), .B(n15618), .Z(n14261) );
  AND U15010 ( .A(n14814), .B(n15653), .Z(n15652) );
  XNOR U15011 ( .A(n15654), .B(n15655), .Z(n14814) );
  ANDN U15012 ( .B(n9014), .A(n14884), .Z(n15609) );
  XNOR U15013 ( .A(n3473), .B(n15656), .Z(n15543) );
  XNOR U15014 ( .A(n9003), .B(n4859), .Z(n15656) );
  XOR U15015 ( .A(n15657), .B(n6542), .Z(n4859) );
  IV U15016 ( .A(n9009), .Z(n6542) );
  XOR U15017 ( .A(n15658), .B(n9358), .Z(n9009) );
  IV U15018 ( .A(n10005), .Z(n9358) );
  XOR U15019 ( .A(n15659), .B(n13333), .Z(n10005) );
  XOR U15020 ( .A(n15660), .B(n15661), .Z(n13333) );
  XNOR U15021 ( .A(n12440), .B(n11704), .Z(n15661) );
  XOR U15022 ( .A(n15662), .B(n15663), .Z(n11704) );
  AND U15023 ( .A(n15664), .B(n15665), .Z(n15662) );
  XNOR U15024 ( .A(n15666), .B(n15667), .Z(n12440) );
  AND U15025 ( .A(n15668), .B(n15669), .Z(n15666) );
  XOR U15026 ( .A(n9550), .B(n15670), .Z(n15660) );
  XOR U15027 ( .A(n10057), .B(n13862), .Z(n15670) );
  XNOR U15028 ( .A(n15671), .B(n15672), .Z(n13862) );
  AND U15029 ( .A(n15673), .B(n15674), .Z(n15671) );
  XNOR U15030 ( .A(n15675), .B(n15676), .Z(n10057) );
  NOR U15031 ( .A(n15677), .B(n15678), .Z(n15675) );
  XNOR U15032 ( .A(n15679), .B(n15680), .Z(n9550) );
  ANDN U15033 ( .B(n15681), .A(n15682), .Z(n15679) );
  AND U15034 ( .A(n8962), .B(n9010), .Z(n15657) );
  XOR U15035 ( .A(n15683), .B(n11522), .Z(n9010) );
  XOR U15036 ( .A(n15684), .B(n14856), .Z(n11522) );
  XOR U15037 ( .A(n15685), .B(n15686), .Z(n14856) );
  XNOR U15038 ( .A(n9812), .B(n10442), .Z(n15686) );
  XNOR U15039 ( .A(n15687), .B(n14692), .Z(n10442) );
  AND U15040 ( .A(n13832), .B(n14693), .Z(n15687) );
  XOR U15041 ( .A(n14704), .B(n15688), .Z(n9812) );
  XOR U15042 ( .A(n15689), .B(n15690), .Z(n15688) );
  NAND U15043 ( .A(n15691), .B(n6455), .Z(n15690) );
  XNOR U15044 ( .A(n14442), .B(n15693), .Z(n15685) );
  XOR U15045 ( .A(n9554), .B(n14684), .Z(n15693) );
  XNOR U15046 ( .A(n15694), .B(n14689), .Z(n14684) );
  AND U15047 ( .A(n13824), .B(n15695), .Z(n15694) );
  XOR U15048 ( .A(n15696), .B(n15697), .Z(n9554) );
  ANDN U15049 ( .B(n13819), .A(n14699), .Z(n15696) );
  XOR U15050 ( .A(n15698), .B(n14696), .Z(n14442) );
  AND U15051 ( .A(n13828), .B(n15699), .Z(n15698) );
  XNOR U15052 ( .A(n10830), .B(n15700), .Z(n8962) );
  XOR U15053 ( .A(n15701), .B(n6539), .Z(n9003) );
  XOR U15054 ( .A(n11062), .B(n13777), .Z(n6539) );
  XNOR U15055 ( .A(n15702), .B(n15703), .Z(n13777) );
  AND U15056 ( .A(n15704), .B(n15168), .Z(n15702) );
  IV U15057 ( .A(n10044), .Z(n11062) );
  XNOR U15058 ( .A(n13049), .B(n14319), .Z(n10044) );
  XNOR U15059 ( .A(n15705), .B(n15706), .Z(n14319) );
  XNOR U15060 ( .A(n15707), .B(n15708), .Z(n15706) );
  XOR U15061 ( .A(n11981), .B(n15709), .Z(n15705) );
  XOR U15062 ( .A(n11708), .B(n11970), .Z(n15709) );
  XOR U15063 ( .A(n15710), .B(n15173), .Z(n11970) );
  NOR U15064 ( .A(n13786), .B(n13784), .Z(n15710) );
  XNOR U15065 ( .A(n15711), .B(n15176), .Z(n11708) );
  ANDN U15066 ( .B(n13774), .A(n13775), .Z(n15711) );
  XNOR U15067 ( .A(n15712), .B(n15166), .Z(n11981) );
  ANDN U15068 ( .B(n13780), .A(n13781), .Z(n15712) );
  XOR U15069 ( .A(n15713), .B(n15714), .Z(n13049) );
  XNOR U15070 ( .A(n15715), .B(n10894), .Z(n15714) );
  XOR U15071 ( .A(n15716), .B(n15186), .Z(n10894) );
  AND U15072 ( .A(n13801), .B(n13799), .Z(n15716) );
  XOR U15073 ( .A(n10447), .B(n15717), .Z(n15713) );
  XNOR U15074 ( .A(n11287), .B(n14852), .Z(n15717) );
  XNOR U15075 ( .A(n15718), .B(n15192), .Z(n14852) );
  NOR U15076 ( .A(n13804), .B(n13803), .Z(n15718) );
  XNOR U15077 ( .A(n15719), .B(n15196), .Z(n11287) );
  IV U15078 ( .A(n15720), .Z(n15196) );
  AND U15079 ( .A(n13792), .B(n13790), .Z(n15719) );
  XNOR U15080 ( .A(n15721), .B(n15722), .Z(n10447) );
  ANDN U15081 ( .B(n13794), .A(n13795), .Z(n15721) );
  AND U15082 ( .A(n8956), .B(n8955), .Z(n15701) );
  IV U15083 ( .A(n9007), .Z(n8955) );
  XOR U15084 ( .A(n11002), .B(n14334), .Z(n9007) );
  XOR U15085 ( .A(n15723), .B(n15724), .Z(n14334) );
  IV U15086 ( .A(n9502), .Z(n11002) );
  XOR U15087 ( .A(n15726), .B(n14802), .Z(n9502) );
  XOR U15088 ( .A(n15727), .B(n15728), .Z(n14802) );
  XOR U15089 ( .A(n14257), .B(n10919), .Z(n15728) );
  XOR U15090 ( .A(n15729), .B(n12380), .Z(n10919) );
  ANDN U15091 ( .B(n15730), .A(n15731), .Z(n15729) );
  XNOR U15092 ( .A(n15732), .B(n15733), .Z(n14257) );
  XOR U15093 ( .A(n13273), .B(n15736), .Z(n15727) );
  XOR U15094 ( .A(n13185), .B(n11006), .Z(n15736) );
  XOR U15095 ( .A(n15737), .B(n12301), .Z(n11006) );
  AND U15096 ( .A(n15738), .B(n15739), .Z(n15737) );
  XNOR U15097 ( .A(n15740), .B(n15230), .Z(n13185) );
  XOR U15098 ( .A(n15743), .B(n12308), .Z(n13273) );
  IV U15099 ( .A(n15744), .Z(n12308) );
  XOR U15100 ( .A(n15747), .B(n11448), .Z(n8956) );
  XOR U15101 ( .A(n15748), .B(n9016), .Z(n3473) );
  XOR U15102 ( .A(n15749), .B(n9805), .Z(n9016) );
  XNOR U15103 ( .A(n13468), .B(n14056), .Z(n9805) );
  XNOR U15104 ( .A(n15750), .B(n15751), .Z(n14056) );
  XOR U15105 ( .A(n14249), .B(n10169), .Z(n15751) );
  XNOR U15106 ( .A(n15752), .B(n15753), .Z(n10169) );
  AND U15107 ( .A(n15754), .B(n15755), .Z(n15752) );
  XNOR U15108 ( .A(n15756), .B(n14152), .Z(n14249) );
  AND U15109 ( .A(n15757), .B(n15758), .Z(n15756) );
  XOR U15110 ( .A(n10300), .B(n15759), .Z(n15750) );
  XOR U15111 ( .A(n9493), .B(n12869), .Z(n15759) );
  XOR U15112 ( .A(n15760), .B(n15450), .Z(n12869) );
  ANDN U15113 ( .B(n15761), .A(n15762), .Z(n15760) );
  XOR U15114 ( .A(n15763), .B(n14143), .Z(n9493) );
  AND U15115 ( .A(n15764), .B(n15765), .Z(n15763) );
  XNOR U15116 ( .A(n15766), .B(n14149), .Z(n10300) );
  ANDN U15117 ( .B(n15767), .A(n15768), .Z(n15766) );
  XOR U15118 ( .A(n15769), .B(n15770), .Z(n13468) );
  XNOR U15119 ( .A(n9935), .B(n11857), .Z(n15770) );
  NOR U15120 ( .A(n15773), .B(n15774), .Z(n15771) );
  XOR U15121 ( .A(n15775), .B(n15776), .Z(n9935) );
  NOR U15122 ( .A(n15777), .B(n14860), .Z(n15775) );
  XNOR U15123 ( .A(n9660), .B(n15778), .Z(n15769) );
  XOR U15124 ( .A(n15779), .B(n15542), .Z(n15778) );
  XNOR U15125 ( .A(n15780), .B(n15781), .Z(n15542) );
  ANDN U15126 ( .B(n15782), .A(n14870), .Z(n15780) );
  XNOR U15127 ( .A(n15783), .B(n15784), .Z(n9660) );
  ANDN U15128 ( .B(n8952), .A(n8953), .Z(n15748) );
  XOR U15129 ( .A(n15786), .B(n10226), .Z(n8953) );
  XNOR U15130 ( .A(n15041), .B(n9913), .Z(n8952) );
  IV U15131 ( .A(n10203), .Z(n9913) );
  XOR U15132 ( .A(n13382), .B(n15787), .Z(n10203) );
  XOR U15133 ( .A(n15788), .B(n15789), .Z(n13382) );
  XOR U15134 ( .A(n14001), .B(n12993), .Z(n15789) );
  XOR U15135 ( .A(n15790), .B(n15791), .Z(n12993) );
  XOR U15136 ( .A(n15792), .B(n15793), .Z(n14001) );
  NOR U15137 ( .A(n13729), .B(n13728), .Z(n15792) );
  XNOR U15138 ( .A(n12053), .B(n15794), .Z(n15788) );
  XNOR U15139 ( .A(n12670), .B(n11585), .Z(n15794) );
  XNOR U15140 ( .A(n15795), .B(n15796), .Z(n11585) );
  NOR U15141 ( .A(n13734), .B(n13733), .Z(n15795) );
  XNOR U15142 ( .A(n15797), .B(n15798), .Z(n12670) );
  ANDN U15143 ( .B(n13724), .A(n13725), .Z(n15797) );
  XNOR U15144 ( .A(n15799), .B(n15800), .Z(n12053) );
  ANDN U15145 ( .B(n15801), .A(n13738), .Z(n15799) );
  XNOR U15146 ( .A(n15802), .B(n15803), .Z(n15041) );
  AND U15147 ( .A(n13203), .B(n15804), .Z(n15802) );
  XNOR U15148 ( .A(n15805), .B(n15806), .Z(n6295) );
  XOR U15149 ( .A(n3685), .B(n5436), .Z(n15806) );
  XOR U15150 ( .A(n15807), .B(n9062), .Z(n5436) );
  IV U15151 ( .A(n9023), .Z(n9062) );
  XOR U15152 ( .A(n14772), .B(n15808), .Z(n9023) );
  XOR U15153 ( .A(n15809), .B(n15556), .Z(n14772) );
  ANDN U15154 ( .B(n15810), .A(n15811), .Z(n15809) );
  AND U15155 ( .A(n6564), .B(n9093), .Z(n15807) );
  IV U15156 ( .A(n6566), .Z(n9093) );
  XOR U15157 ( .A(n15812), .B(n10226), .Z(n6566) );
  XOR U15158 ( .A(n15813), .B(n15814), .Z(n10226) );
  XNOR U15159 ( .A(n12145), .B(n12894), .Z(n6564) );
  XNOR U15160 ( .A(n15815), .B(n15004), .Z(n12894) );
  AND U15161 ( .A(n15357), .B(n15816), .Z(n15815) );
  XOR U15162 ( .A(n15817), .B(n7037), .Z(n3685) );
  XNOR U15163 ( .A(n9684), .B(n13211), .Z(n7037) );
  XNOR U15164 ( .A(n15818), .B(n15035), .Z(n13211) );
  XOR U15165 ( .A(n10488), .B(n14879), .Z(n9684) );
  XNOR U15166 ( .A(n15821), .B(n15822), .Z(n14879) );
  XOR U15167 ( .A(n13366), .B(n12730), .Z(n15822) );
  XOR U15168 ( .A(n15823), .B(n15044), .Z(n12730) );
  ANDN U15169 ( .B(n13217), .A(n13218), .Z(n15823) );
  XNOR U15170 ( .A(n15824), .B(n15825), .Z(n13217) );
  XOR U15171 ( .A(n15826), .B(n15039), .Z(n13366) );
  ANDN U15172 ( .B(n13207), .A(n13208), .Z(n15826) );
  XOR U15173 ( .A(n15827), .B(n15828), .Z(n13207) );
  XOR U15174 ( .A(n11891), .B(n15829), .Z(n15821) );
  XOR U15175 ( .A(n12554), .B(n11434), .Z(n15829) );
  XOR U15176 ( .A(n15830), .B(n15036), .Z(n11434) );
  ANDN U15177 ( .B(n15820), .A(n15035), .Z(n15830) );
  XOR U15178 ( .A(n15831), .B(n15832), .Z(n15035) );
  XOR U15179 ( .A(n15833), .B(n15834), .Z(n12554) );
  XOR U15180 ( .A(n15835), .B(n15249), .Z(n13203) );
  XOR U15181 ( .A(n15836), .B(n15047), .Z(n11891) );
  XNOR U15182 ( .A(n15837), .B(n15838), .Z(n13213) );
  XOR U15183 ( .A(n15839), .B(n15840), .Z(n10488) );
  XOR U15184 ( .A(n10604), .B(n11242), .Z(n15840) );
  XOR U15185 ( .A(n15841), .B(n13738), .Z(n11242) );
  XOR U15186 ( .A(n15842), .B(n15843), .Z(n13738) );
  ANDN U15187 ( .B(n13739), .A(n15844), .Z(n15841) );
  XNOR U15188 ( .A(n15845), .B(n13742), .Z(n10604) );
  XOR U15189 ( .A(n15846), .B(n15591), .Z(n13742) );
  XOR U15190 ( .A(n10264), .B(n15848), .Z(n15839) );
  XNOR U15191 ( .A(n13700), .B(n11829), .Z(n15848) );
  XNOR U15192 ( .A(n15849), .B(n13725), .Z(n11829) );
  XOR U15193 ( .A(n15850), .B(n15851), .Z(n13725) );
  AND U15194 ( .A(n15852), .B(n15853), .Z(n15849) );
  XOR U15195 ( .A(n15854), .B(n13734), .Z(n13700) );
  XNOR U15196 ( .A(n15855), .B(n15856), .Z(n13734) );
  ANDN U15197 ( .B(n13735), .A(n15857), .Z(n15854) );
  XNOR U15198 ( .A(n15858), .B(n13729), .Z(n10264) );
  XNOR U15199 ( .A(n15831), .B(n15859), .Z(n13729) );
  ANDN U15200 ( .B(n15860), .A(n15861), .Z(n15858) );
  ANDN U15201 ( .B(n6557), .A(n6555), .Z(n15817) );
  XOR U15202 ( .A(n15862), .B(n11926), .Z(n6555) );
  XOR U15203 ( .A(n11789), .B(n15863), .Z(n11926) );
  XOR U15204 ( .A(n15864), .B(n15865), .Z(n11789) );
  XNOR U15205 ( .A(n10674), .B(n12713), .Z(n15865) );
  XNOR U15206 ( .A(n15866), .B(n15867), .Z(n12713) );
  AND U15207 ( .A(n15868), .B(n15869), .Z(n15866) );
  XNOR U15208 ( .A(n15870), .B(n15871), .Z(n10674) );
  NOR U15209 ( .A(n15872), .B(n15873), .Z(n15870) );
  XOR U15210 ( .A(n11551), .B(n15874), .Z(n15864) );
  XOR U15211 ( .A(n12230), .B(n12221), .Z(n15874) );
  XNOR U15212 ( .A(n15875), .B(n15876), .Z(n12221) );
  AND U15213 ( .A(n15877), .B(n15878), .Z(n15875) );
  XNOR U15214 ( .A(n15879), .B(n15880), .Z(n12230) );
  AND U15215 ( .A(n15881), .B(n15882), .Z(n15879) );
  XNOR U15216 ( .A(n15883), .B(n15884), .Z(n11551) );
  ANDN U15217 ( .B(n15885), .A(n15886), .Z(n15883) );
  XNOR U15218 ( .A(n11401), .B(n15887), .Z(n6557) );
  IV U15219 ( .A(n10100), .Z(n11401) );
  XOR U15220 ( .A(n12834), .B(n14014), .Z(n10100) );
  XNOR U15221 ( .A(n15888), .B(n15889), .Z(n14014) );
  XOR U15222 ( .A(n15890), .B(n12331), .Z(n15889) );
  XOR U15223 ( .A(n15891), .B(n13143), .Z(n12331) );
  NOR U15224 ( .A(n14012), .B(n14013), .Z(n15891) );
  XOR U15225 ( .A(n10782), .B(n15892), .Z(n15888) );
  XNOR U15226 ( .A(n13551), .B(n12151), .Z(n15892) );
  XNOR U15227 ( .A(n15893), .B(n13138), .Z(n12151) );
  AND U15228 ( .A(n13622), .B(n15894), .Z(n15893) );
  XNOR U15229 ( .A(n15895), .B(n15896), .Z(n13551) );
  ANDN U15230 ( .B(n13614), .A(n13615), .Z(n15895) );
  XNOR U15231 ( .A(n15897), .B(n15898), .Z(n10782) );
  XOR U15232 ( .A(n15899), .B(n15900), .Z(n12834) );
  XNOR U15233 ( .A(n11535), .B(n9903), .Z(n15900) );
  XOR U15234 ( .A(n15901), .B(n13363), .Z(n9903) );
  IV U15235 ( .A(n12965), .Z(n13363) );
  XNOR U15236 ( .A(n15902), .B(n15903), .Z(n12965) );
  NOR U15237 ( .A(n14921), .B(n12964), .Z(n15901) );
  XNOR U15238 ( .A(n12951), .B(n15904), .Z(n11535) );
  XOR U15239 ( .A(rc_i[1]), .B(n15905), .Z(n15904) );
  OR U15240 ( .A(n14913), .B(n12952), .Z(n15905) );
  XNOR U15241 ( .A(n15906), .B(n15907), .Z(n12951) );
  XOR U15242 ( .A(n11745), .B(n15908), .Z(n15899) );
  XNOR U15243 ( .A(n12199), .B(n9405), .Z(n15908) );
  XNOR U15244 ( .A(n15909), .B(n12956), .Z(n9405) );
  XNOR U15245 ( .A(n15910), .B(n15911), .Z(n12956) );
  NOR U15246 ( .A(n12957), .B(n14917), .Z(n15909) );
  XOR U15247 ( .A(n15912), .B(n13379), .Z(n12199) );
  IV U15248 ( .A(n13120), .Z(n13379) );
  XNOR U15249 ( .A(n15913), .B(n15914), .Z(n13120) );
  NOR U15250 ( .A(n13119), .B(n14903), .Z(n15912) );
  XNOR U15251 ( .A(n15915), .B(n12960), .Z(n11745) );
  XNOR U15252 ( .A(n15916), .B(n15917), .Z(n12960) );
  AND U15253 ( .A(n14907), .B(n12961), .Z(n15915) );
  XOR U15254 ( .A(n4295), .B(n15918), .Z(n15805) );
  XNOR U15255 ( .A(n5875), .B(n2127), .Z(n15918) );
  XNOR U15256 ( .A(n15919), .B(n7028), .Z(n2127) );
  XNOR U15257 ( .A(n12808), .B(n9163), .Z(n7028) );
  XOR U15258 ( .A(n13919), .B(n15920), .Z(n9163) );
  XOR U15259 ( .A(n15921), .B(n15922), .Z(n13919) );
  XOR U15260 ( .A(n12464), .B(n13086), .Z(n15922) );
  XNOR U15261 ( .A(n15923), .B(n15924), .Z(n13086) );
  AND U15262 ( .A(n15925), .B(n15926), .Z(n15923) );
  XNOR U15263 ( .A(n15927), .B(n15928), .Z(n12464) );
  ANDN U15264 ( .B(n15929), .A(n15930), .Z(n15927) );
  XOR U15265 ( .A(n11862), .B(n15931), .Z(n15921) );
  XOR U15266 ( .A(n11070), .B(n11397), .Z(n15931) );
  XOR U15267 ( .A(n15932), .B(n15933), .Z(n11397) );
  XNOR U15268 ( .A(n15936), .B(n15937), .Z(n11070) );
  ANDN U15269 ( .B(n15938), .A(n15939), .Z(n15936) );
  XOR U15270 ( .A(n15940), .B(n15941), .Z(n11862) );
  ANDN U15271 ( .B(n15942), .A(n15943), .Z(n15940) );
  XOR U15272 ( .A(n15944), .B(n15945), .Z(n12808) );
  ANDN U15273 ( .B(n15946), .A(n15947), .Z(n15944) );
  AND U15274 ( .A(n6560), .B(n6562), .Z(n15919) );
  XOR U15275 ( .A(n15948), .B(n10539), .Z(n6562) );
  IV U15276 ( .A(n9989), .Z(n10539) );
  XOR U15277 ( .A(n15949), .B(n14318), .Z(n9989) );
  XOR U15278 ( .A(n15950), .B(n15951), .Z(n14318) );
  XNOR U15279 ( .A(n12582), .B(n10381), .Z(n15951) );
  XOR U15280 ( .A(n15952), .B(n13238), .Z(n10381) );
  IV U15281 ( .A(n13755), .Z(n13238) );
  XOR U15282 ( .A(n15953), .B(n15954), .Z(n13755) );
  ANDN U15283 ( .B(n15955), .A(n15956), .Z(n15952) );
  XOR U15284 ( .A(n15957), .B(n13763), .Z(n12582) );
  XOR U15285 ( .A(n15958), .B(n15959), .Z(n13763) );
  AND U15286 ( .A(n13762), .B(n15960), .Z(n15957) );
  XOR U15287 ( .A(n12247), .B(n15961), .Z(n15950) );
  XOR U15288 ( .A(n12238), .B(n10546), .Z(n15961) );
  XNOR U15289 ( .A(n15962), .B(n13751), .Z(n10546) );
  ANDN U15290 ( .B(n13752), .A(n15963), .Z(n15962) );
  XNOR U15291 ( .A(n15964), .B(n13233), .Z(n12238) );
  XNOR U15292 ( .A(n15965), .B(n15533), .Z(n13233) );
  ANDN U15293 ( .B(n13765), .A(n15966), .Z(n15964) );
  XNOR U15294 ( .A(n15967), .B(n13243), .Z(n12247) );
  XOR U15295 ( .A(n15252), .B(n15968), .Z(n13243) );
  ANDN U15296 ( .B(n13759), .A(n15969), .Z(n15967) );
  XNOR U15297 ( .A(n14529), .B(n11177), .Z(n6560) );
  IV U15298 ( .A(n9766), .Z(n11177) );
  XNOR U15299 ( .A(n12390), .B(n12829), .Z(n9766) );
  XNOR U15300 ( .A(n15970), .B(n15971), .Z(n12829) );
  XOR U15301 ( .A(n14958), .B(n9670), .Z(n15971) );
  XNOR U15302 ( .A(n15972), .B(n13987), .Z(n9670) );
  AND U15303 ( .A(n14523), .B(n15973), .Z(n15972) );
  XNOR U15304 ( .A(n15974), .B(n15975), .Z(n14523) );
  XNOR U15305 ( .A(n15976), .B(n13973), .Z(n14958) );
  ANDN U15306 ( .B(n15977), .A(n15978), .Z(n15976) );
  XNOR U15307 ( .A(n10426), .B(n15979), .Z(n15970) );
  XOR U15308 ( .A(n10375), .B(n15980), .Z(n15979) );
  XOR U15309 ( .A(n15981), .B(n13979), .Z(n10375) );
  AND U15310 ( .A(n14532), .B(n15982), .Z(n15981) );
  XNOR U15311 ( .A(n15983), .B(n15984), .Z(n14532) );
  XOR U15312 ( .A(n15985), .B(n13969), .Z(n10426) );
  NOR U15313 ( .A(n14535), .B(n14534), .Z(n15985) );
  XOR U15314 ( .A(n15986), .B(n15987), .Z(n14535) );
  XOR U15315 ( .A(n15988), .B(n15989), .Z(n12390) );
  XOR U15316 ( .A(n15990), .B(n12613), .Z(n15989) );
  XNOR U15317 ( .A(n15991), .B(n15992), .Z(n12613) );
  NOR U15318 ( .A(n14504), .B(n14503), .Z(n15991) );
  XOR U15319 ( .A(n12175), .B(n15993), .Z(n15988) );
  XOR U15320 ( .A(n15994), .B(n12967), .Z(n15993) );
  XOR U15321 ( .A(n15995), .B(n15996), .Z(n12967) );
  XOR U15322 ( .A(n15997), .B(n15998), .Z(n12175) );
  NOR U15323 ( .A(n14512), .B(n14514), .Z(n15997) );
  XOR U15324 ( .A(n15999), .B(n15978), .Z(n14529) );
  ANDN U15325 ( .B(n14938), .A(n13972), .Z(n15999) );
  XNOR U15326 ( .A(n16000), .B(n16001), .Z(n13972) );
  IV U15327 ( .A(n15977), .Z(n14938) );
  XNOR U15328 ( .A(n16002), .B(n16003), .Z(n15977) );
  XOR U15329 ( .A(n16004), .B(n7034), .Z(n5875) );
  XOR U15330 ( .A(n15348), .B(n11979), .Z(n7034) );
  IV U15331 ( .A(n11055), .Z(n11979) );
  XOR U15332 ( .A(n13313), .B(n14683), .Z(n11055) );
  XNOR U15333 ( .A(n16005), .B(n16006), .Z(n14683) );
  XOR U15334 ( .A(n9583), .B(n11114), .Z(n16006) );
  XOR U15335 ( .A(n16007), .B(n12907), .Z(n11114) );
  XNOR U15336 ( .A(n16008), .B(n16009), .Z(n14117) );
  XOR U15337 ( .A(n16010), .B(n16011), .Z(n12908) );
  XOR U15338 ( .A(n16012), .B(n12904), .Z(n9583) );
  XOR U15339 ( .A(n16013), .B(n16014), .Z(n14109) );
  XNOR U15340 ( .A(n16015), .B(n16016), .Z(n12903) );
  XOR U15341 ( .A(n9786), .B(n16017), .Z(n16005) );
  XOR U15342 ( .A(n11843), .B(n10257), .Z(n16017) );
  XOR U15343 ( .A(n16018), .B(n16019), .Z(n10257) );
  NOR U15344 ( .A(n15002), .B(n15357), .Z(n16018) );
  XOR U15345 ( .A(n16020), .B(n16021), .Z(n15357) );
  XNOR U15346 ( .A(n16022), .B(n14910), .Z(n15002) );
  XNOR U15347 ( .A(n16023), .B(n12899), .Z(n11843) );
  NOR U15348 ( .A(n14112), .B(n12900), .Z(n16023) );
  XOR U15349 ( .A(n16024), .B(n16025), .Z(n12900) );
  XNOR U15350 ( .A(n16026), .B(n16027), .Z(n14112) );
  XNOR U15351 ( .A(n16028), .B(n16029), .Z(n9786) );
  NOR U15352 ( .A(n14120), .B(n15366), .Z(n16028) );
  XNOR U15353 ( .A(n16030), .B(n16031), .Z(n14120) );
  XOR U15354 ( .A(n16032), .B(n16033), .Z(n13313) );
  XOR U15355 ( .A(n12688), .B(n12865), .Z(n16033) );
  XOR U15356 ( .A(n16034), .B(n14414), .Z(n12865) );
  XNOR U15357 ( .A(n16035), .B(n16036), .Z(n14414) );
  ANDN U15358 ( .B(n15601), .A(n15304), .Z(n16034) );
  XOR U15359 ( .A(n16037), .B(n14418), .Z(n12688) );
  IV U15360 ( .A(n15307), .Z(n14418) );
  XNOR U15361 ( .A(n16038), .B(n16039), .Z(n15307) );
  NOR U15362 ( .A(n15306), .B(n15353), .Z(n16037) );
  XNOR U15363 ( .A(n16040), .B(n16041), .Z(n15353) );
  XNOR U15364 ( .A(n16042), .B(n16043), .Z(n15306) );
  XOR U15365 ( .A(n11706), .B(n16044), .Z(n16032) );
  XOR U15366 ( .A(n10793), .B(n12890), .Z(n16044) );
  XNOR U15367 ( .A(n16045), .B(n14409), .Z(n12890) );
  XNOR U15368 ( .A(n16046), .B(n16047), .Z(n14409) );
  NOR U15369 ( .A(n15310), .B(n15346), .Z(n16045) );
  XNOR U15370 ( .A(n16048), .B(n14948), .Z(n15346) );
  XNOR U15371 ( .A(n16049), .B(n16050), .Z(n15310) );
  XNOR U15372 ( .A(n16051), .B(n14422), .Z(n10793) );
  XNOR U15373 ( .A(n16052), .B(n16053), .Z(n14422) );
  ANDN U15374 ( .B(n15312), .A(n15350), .Z(n16051) );
  XNOR U15375 ( .A(n16056), .B(n16057), .Z(n15312) );
  XOR U15376 ( .A(n16058), .B(n14426), .Z(n11706) );
  XNOR U15377 ( .A(n16059), .B(n16060), .Z(n14426) );
  ANDN U15378 ( .B(n15314), .A(n15344), .Z(n16058) );
  XNOR U15379 ( .A(n16061), .B(n16062), .Z(n15344) );
  XOR U15380 ( .A(n16063), .B(n16064), .Z(n15314) );
  XNOR U15381 ( .A(n16065), .B(n15304), .Z(n15348) );
  XNOR U15382 ( .A(n16066), .B(n16067), .Z(n15304) );
  NOR U15383 ( .A(n14412), .B(n15601), .Z(n16065) );
  XOR U15384 ( .A(n16068), .B(n16069), .Z(n15601) );
  XOR U15385 ( .A(n16070), .B(n16071), .Z(n14412) );
  ANDN U15386 ( .B(n6553), .A(n6551), .Z(n16004) );
  XOR U15387 ( .A(n16072), .B(n9370), .Z(n6551) );
  XNOR U15388 ( .A(n12224), .B(n13385), .Z(n9370) );
  XNOR U15389 ( .A(n16073), .B(n16074), .Z(n13385) );
  XNOR U15390 ( .A(n13998), .B(n11443), .Z(n16074) );
  XNOR U15391 ( .A(n16075), .B(n16076), .Z(n11443) );
  AND U15392 ( .A(n16077), .B(n16078), .Z(n16075) );
  XNOR U15393 ( .A(n16079), .B(n12412), .Z(n13998) );
  ANDN U15394 ( .B(n16080), .A(n16081), .Z(n16079) );
  XOR U15395 ( .A(n9197), .B(n16082), .Z(n16073) );
  XOR U15396 ( .A(n10602), .B(n16083), .Z(n16082) );
  XNOR U15397 ( .A(n16084), .B(n14402), .Z(n10602) );
  AND U15398 ( .A(n16085), .B(n16086), .Z(n16084) );
  XNOR U15399 ( .A(n16087), .B(n13654), .Z(n9197) );
  AND U15400 ( .A(n16088), .B(n16089), .Z(n16087) );
  XOR U15401 ( .A(n16090), .B(n16091), .Z(n12224) );
  XOR U15402 ( .A(n12275), .B(n13605), .Z(n16091) );
  XOR U15403 ( .A(n16092), .B(n14510), .Z(n13605) );
  ANDN U15404 ( .B(n16093), .A(n14509), .Z(n16092) );
  XNOR U15405 ( .A(n16094), .B(n14514), .Z(n12275) );
  XNOR U15406 ( .A(n16095), .B(n15529), .Z(n14514) );
  ANDN U15407 ( .B(n16096), .A(n14513), .Z(n16094) );
  XOR U15408 ( .A(n11575), .B(n16097), .Z(n16090) );
  XOR U15409 ( .A(n10463), .B(n13154), .Z(n16097) );
  XNOR U15410 ( .A(n16098), .B(n14504), .Z(n13154) );
  XNOR U15411 ( .A(n16099), .B(n16100), .Z(n14504) );
  AND U15412 ( .A(n16101), .B(n16102), .Z(n16098) );
  XNOR U15413 ( .A(n16103), .B(n14517), .Z(n10463) );
  XNOR U15414 ( .A(n16104), .B(n15222), .Z(n14517) );
  ANDN U15415 ( .B(n16105), .A(n16106), .Z(n16103) );
  XNOR U15416 ( .A(n16107), .B(n14500), .Z(n11575) );
  XNOR U15417 ( .A(n11510), .B(n16109), .Z(n6553) );
  IV U15418 ( .A(n9597), .Z(n11510) );
  XOR U15419 ( .A(n16110), .B(n11757), .Z(n9597) );
  XNOR U15420 ( .A(n16111), .B(n16112), .Z(n11757) );
  XNOR U15421 ( .A(n11289), .B(n12281), .Z(n16112) );
  XOR U15422 ( .A(n16113), .B(n13585), .Z(n12281) );
  IV U15423 ( .A(n16115), .Z(n13581) );
  XNOR U15424 ( .A(n16116), .B(n12518), .Z(n11289) );
  ANDN U15425 ( .B(n16117), .A(n13577), .Z(n16116) );
  XOR U15426 ( .A(n11066), .B(n16118), .Z(n16111) );
  XOR U15427 ( .A(n16119), .B(n11527), .Z(n16118) );
  XNOR U15428 ( .A(n16120), .B(n12515), .Z(n11527) );
  ANDN U15429 ( .B(n16121), .A(n13579), .Z(n16120) );
  XNOR U15430 ( .A(n16122), .B(n13196), .Z(n11066) );
  XOR U15431 ( .A(n16124), .B(n7025), .Z(n4295) );
  XNOR U15432 ( .A(n16125), .B(n10691), .Z(n7025) );
  AND U15433 ( .A(n6568), .B(n9099), .Z(n16124) );
  IV U15434 ( .A(n6570), .Z(n9099) );
  XOR U15435 ( .A(n16128), .B(n9810), .Z(n6570) );
  XNOR U15436 ( .A(n16129), .B(n11448), .Z(n6568) );
  IV U15437 ( .A(n11320), .Z(n11448) );
  XNOR U15438 ( .A(n12715), .B(n16130), .Z(n11320) );
  XOR U15439 ( .A(n16131), .B(n16132), .Z(n12715) );
  XOR U15440 ( .A(n12159), .B(n13044), .Z(n16132) );
  XNOR U15441 ( .A(n16133), .B(n16134), .Z(n13044) );
  AND U15442 ( .A(n16135), .B(n14989), .Z(n16133) );
  XOR U15443 ( .A(n16136), .B(n16137), .Z(n12159) );
  ANDN U15444 ( .B(n14993), .A(n16138), .Z(n16136) );
  XOR U15445 ( .A(n12089), .B(n16139), .Z(n16131) );
  XOR U15446 ( .A(n9078), .B(n14758), .Z(n16139) );
  XOR U15447 ( .A(n16140), .B(n16141), .Z(n14758) );
  ANDN U15448 ( .B(n16142), .A(n14979), .Z(n16140) );
  XNOR U15449 ( .A(n16143), .B(n16144), .Z(n9078) );
  ANDN U15450 ( .B(n16145), .A(n16146), .Z(n16143) );
  XNOR U15451 ( .A(n16147), .B(n16148), .Z(n12089) );
  XNOR U15452 ( .A(n16150), .B(n9014), .Z(n8959) );
  XNOR U15453 ( .A(n16151), .B(n12604), .Z(n9014) );
  ANDN U15454 ( .B(n14884), .A(n6528), .Z(n16150) );
  XNOR U15455 ( .A(n14668), .B(n11602), .Z(n6528) );
  IV U15456 ( .A(n11675), .Z(n11602) );
  XNOR U15457 ( .A(n16152), .B(n11845), .Z(n11675) );
  XNOR U15458 ( .A(n16153), .B(n16154), .Z(n11845) );
  XNOR U15459 ( .A(n12462), .B(n10552), .Z(n16154) );
  XOR U15460 ( .A(n16155), .B(n16156), .Z(n10552) );
  AND U15461 ( .A(n16157), .B(n16158), .Z(n16155) );
  XNOR U15462 ( .A(n16159), .B(n16160), .Z(n12462) );
  ANDN U15463 ( .B(n14677), .A(n14678), .Z(n16159) );
  XNOR U15464 ( .A(n11411), .B(n16161), .Z(n16153) );
  XOR U15465 ( .A(n16162), .B(n12088), .Z(n16161) );
  XNOR U15466 ( .A(n16163), .B(n13299), .Z(n12088) );
  AND U15467 ( .A(n14682), .B(n16164), .Z(n16163) );
  XNOR U15468 ( .A(n16165), .B(n13294), .Z(n11411) );
  AND U15469 ( .A(n14670), .B(n14671), .Z(n16165) );
  XNOR U15470 ( .A(n16166), .B(n16157), .Z(n14668) );
  XOR U15471 ( .A(n10649), .B(n16167), .Z(n14884) );
  IV U15472 ( .A(n9574), .Z(n10649) );
  XOR U15473 ( .A(n16168), .B(n13836), .Z(n9574) );
  XOR U15474 ( .A(n16169), .B(n16170), .Z(n13836) );
  XNOR U15475 ( .A(n12933), .B(n12474), .Z(n16170) );
  XOR U15476 ( .A(n16171), .B(n16172), .Z(n12474) );
  ANDN U15477 ( .B(n16173), .A(n16174), .Z(n16171) );
  XOR U15478 ( .A(n16175), .B(n16176), .Z(n12933) );
  NOR U15479 ( .A(n16177), .B(n16178), .Z(n16175) );
  XOR U15480 ( .A(n11572), .B(n16179), .Z(n16169) );
  XOR U15481 ( .A(n12267), .B(n11292), .Z(n16179) );
  XNOR U15482 ( .A(n16180), .B(n16181), .Z(n11292) );
  NOR U15483 ( .A(n16182), .B(n16183), .Z(n16180) );
  XNOR U15484 ( .A(n16184), .B(n16185), .Z(n12267) );
  NOR U15485 ( .A(n16186), .B(n16187), .Z(n16184) );
  XOR U15486 ( .A(n16188), .B(n16189), .Z(n11572) );
  NOR U15487 ( .A(n16190), .B(n16191), .Z(n16188) );
  XOR U15488 ( .A(n12026), .B(n2092), .Z(n5661) );
  XNOR U15489 ( .A(n8345), .B(n9855), .Z(n2092) );
  XNOR U15490 ( .A(n16192), .B(n16193), .Z(n9855) );
  XOR U15491 ( .A(n5473), .B(n3597), .Z(n16193) );
  XOR U15492 ( .A(n16194), .B(n8438), .Z(n3597) );
  IV U15493 ( .A(n12117), .Z(n8438) );
  XOR U15494 ( .A(n16195), .B(n12857), .Z(n12117) );
  IV U15495 ( .A(n12604), .Z(n12857) );
  XOR U15496 ( .A(n16196), .B(n16197), .Z(n12604) );
  ANDN U15497 ( .B(n8490), .A(n8491), .Z(n16194) );
  XOR U15498 ( .A(n16198), .B(n11072), .Z(n8491) );
  XNOR U15499 ( .A(n16199), .B(n15582), .Z(n11072) );
  XOR U15500 ( .A(n16200), .B(n16201), .Z(n15582) );
  XNOR U15501 ( .A(n10693), .B(n12416), .Z(n16201) );
  XNOR U15502 ( .A(n16202), .B(n14388), .Z(n12416) );
  NOR U15503 ( .A(n14387), .B(n15293), .Z(n16202) );
  XNOR U15504 ( .A(n16203), .B(n14378), .Z(n10693) );
  AND U15505 ( .A(n15296), .B(n14379), .Z(n16203) );
  XOR U15506 ( .A(n12665), .B(n16204), .Z(n16200) );
  XNOR U15507 ( .A(n12641), .B(n11727), .Z(n16204) );
  XNOR U15508 ( .A(n16205), .B(n14383), .Z(n11727) );
  ANDN U15509 ( .B(n14384), .A(n15289), .Z(n16205) );
  XOR U15510 ( .A(n16206), .B(n14374), .Z(n12641) );
  AND U15511 ( .A(n15299), .B(n16207), .Z(n16206) );
  XNOR U15512 ( .A(n16208), .B(n14393), .Z(n12665) );
  ANDN U15513 ( .B(n16209), .A(n15286), .Z(n16208) );
  XOR U15514 ( .A(n16210), .B(n9496), .Z(n8490) );
  IV U15515 ( .A(n11837), .Z(n9496) );
  XNOR U15516 ( .A(n16212), .B(n16213), .Z(n15030) );
  XOR U15517 ( .A(n16214), .B(n11763), .Z(n16213) );
  XOR U15518 ( .A(n16215), .B(n16191), .Z(n11763) );
  AND U15519 ( .A(n16216), .B(n16217), .Z(n16215) );
  XNOR U15520 ( .A(n10018), .B(n16218), .Z(n16212) );
  XOR U15521 ( .A(n12858), .B(n10556), .Z(n16218) );
  XNOR U15522 ( .A(n16219), .B(n16186), .Z(n10556) );
  AND U15523 ( .A(n16220), .B(n16221), .Z(n16219) );
  XNOR U15524 ( .A(n16222), .B(n16183), .Z(n12858) );
  ANDN U15525 ( .B(n16223), .A(n16224), .Z(n16222) );
  XNOR U15526 ( .A(n16225), .B(n16226), .Z(n10018) );
  AND U15527 ( .A(n16227), .B(n16228), .Z(n16225) );
  XNOR U15528 ( .A(n16229), .B(n12110), .Z(n5473) );
  XNOR U15529 ( .A(n16230), .B(n10730), .Z(n12110) );
  XOR U15530 ( .A(n15814), .B(n16231), .Z(n10730) );
  XOR U15531 ( .A(n16232), .B(n16233), .Z(n15814) );
  XOR U15532 ( .A(n11787), .B(n12804), .Z(n16233) );
  XOR U15533 ( .A(n16234), .B(n12817), .Z(n12804) );
  AND U15534 ( .A(n12818), .B(n16235), .Z(n16234) );
  XNOR U15535 ( .A(n16236), .B(n15946), .Z(n11787) );
  AND U15536 ( .A(n15947), .B(n16237), .Z(n16236) );
  XNOR U15537 ( .A(n10564), .B(n16238), .Z(n16232) );
  XOR U15538 ( .A(n12323), .B(n11698), .Z(n16238) );
  XOR U15539 ( .A(n16239), .B(n14322), .Z(n11698) );
  ANDN U15540 ( .B(n14323), .A(n16240), .Z(n16239) );
  XNOR U15541 ( .A(n16241), .B(n12812), .Z(n12323) );
  ANDN U15542 ( .B(n12811), .A(n16242), .Z(n16241) );
  XNOR U15543 ( .A(n16243), .B(n12822), .Z(n10564) );
  ANDN U15544 ( .B(n12821), .A(n16244), .Z(n16243) );
  ANDN U15545 ( .B(n8488), .A(n8486), .Z(n16229) );
  XNOR U15546 ( .A(n15024), .B(n10251), .Z(n8486) );
  XOR U15547 ( .A(n16245), .B(n16246), .Z(n15024) );
  AND U15548 ( .A(n15480), .B(n15478), .Z(n16245) );
  XNOR U15549 ( .A(n16247), .B(n10679), .Z(n8488) );
  XNOR U15550 ( .A(n14196), .B(n13746), .Z(n10679) );
  XNOR U15551 ( .A(n16248), .B(n16249), .Z(n13746) );
  XOR U15552 ( .A(n10145), .B(n9816), .Z(n16249) );
  XNOR U15553 ( .A(n16250), .B(n15027), .Z(n9816) );
  XNOR U15554 ( .A(n16251), .B(n16252), .Z(n15027) );
  AND U15555 ( .A(n15487), .B(n16253), .Z(n16250) );
  XNOR U15556 ( .A(n16254), .B(n15021), .Z(n10145) );
  XNOR U15557 ( .A(n16255), .B(n16256), .Z(n15021) );
  AND U15558 ( .A(n15485), .B(n16257), .Z(n16254) );
  XOR U15559 ( .A(n11523), .B(n16258), .Z(n16248) );
  XOR U15560 ( .A(n10708), .B(n11512), .Z(n16258) );
  XNOR U15561 ( .A(n16259), .B(n15480), .Z(n11512) );
  XNOR U15562 ( .A(n16260), .B(n16261), .Z(n15480) );
  AND U15563 ( .A(n15479), .B(n16262), .Z(n16259) );
  XNOR U15564 ( .A(n16263), .B(n16264), .Z(n10708) );
  AND U15565 ( .A(n16265), .B(n16266), .Z(n16263) );
  XNOR U15566 ( .A(n16267), .B(n15016), .Z(n11523) );
  XNOR U15567 ( .A(n16268), .B(n16269), .Z(n15016) );
  ANDN U15568 ( .B(n15483), .A(n16270), .Z(n16267) );
  XOR U15569 ( .A(n16271), .B(n16272), .Z(n14196) );
  XNOR U15570 ( .A(n12186), .B(n15451), .Z(n16272) );
  XOR U15571 ( .A(n16273), .B(n16274), .Z(n15451) );
  NOR U15572 ( .A(n15465), .B(n14485), .Z(n16273) );
  XOR U15573 ( .A(n16275), .B(n16276), .Z(n12186) );
  XOR U15574 ( .A(n14492), .B(n16277), .Z(n16271) );
  XOR U15575 ( .A(n14707), .B(n10234), .Z(n16277) );
  XOR U15576 ( .A(n16278), .B(n16279), .Z(n10234) );
  XOR U15577 ( .A(n16280), .B(n16281), .Z(n14707) );
  NOR U15578 ( .A(n15469), .B(n16282), .Z(n16280) );
  XOR U15579 ( .A(n16283), .B(n16284), .Z(n14492) );
  NOR U15580 ( .A(n14489), .B(n15455), .Z(n16283) );
  XNOR U15581 ( .A(n6253), .B(n16285), .Z(n16192) );
  XOR U15582 ( .A(n2392), .B(n5676), .Z(n16285) );
  XNOR U15583 ( .A(n16286), .B(n8425), .Z(n5676) );
  XOR U15584 ( .A(n9526), .B(n14748), .Z(n8425) );
  XOR U15585 ( .A(n16287), .B(n16288), .Z(n14748) );
  ANDN U15586 ( .B(n16289), .A(n16290), .Z(n16287) );
  XOR U15587 ( .A(n11277), .B(n11074), .Z(n9526) );
  XOR U15588 ( .A(n16291), .B(n16292), .Z(n11074) );
  XOR U15589 ( .A(n11161), .B(n12131), .Z(n16292) );
  XOR U15590 ( .A(n16293), .B(n16294), .Z(n12131) );
  AND U15591 ( .A(n11964), .B(n11966), .Z(n16293) );
  XNOR U15592 ( .A(n16295), .B(n16296), .Z(n11161) );
  XOR U15593 ( .A(n11693), .B(n16297), .Z(n16291) );
  XOR U15594 ( .A(n16298), .B(n11390), .Z(n16297) );
  XNOR U15595 ( .A(n16299), .B(n16300), .Z(n11390) );
  XNOR U15596 ( .A(n16301), .B(n16302), .Z(n11693) );
  XOR U15597 ( .A(n16303), .B(n16304), .Z(n11277) );
  XOR U15598 ( .A(n12365), .B(n12787), .Z(n16304) );
  XOR U15599 ( .A(n16305), .B(n16306), .Z(n12787) );
  ANDN U15600 ( .B(n14956), .A(n14955), .Z(n16305) );
  XNOR U15601 ( .A(n16307), .B(n16308), .Z(n12365) );
  ANDN U15602 ( .B(n16309), .A(n14753), .Z(n16307) );
  XNOR U15603 ( .A(n12636), .B(n16310), .Z(n16303) );
  XNOR U15604 ( .A(n16311), .B(n14997), .Z(n16310) );
  XOR U15605 ( .A(n16312), .B(n16313), .Z(n14997) );
  NOR U15606 ( .A(n14742), .B(n14741), .Z(n16312) );
  XNOR U15607 ( .A(n16314), .B(n16315), .Z(n12636) );
  AND U15608 ( .A(n9858), .B(n12115), .Z(n16286) );
  XNOR U15609 ( .A(n15990), .B(n12176), .Z(n12115) );
  XNOR U15610 ( .A(n16316), .B(n16317), .Z(n15990) );
  ANDN U15611 ( .B(n14499), .A(n14500), .Z(n16316) );
  XNOR U15612 ( .A(n16318), .B(n16319), .Z(n14500) );
  XOR U15613 ( .A(n14770), .B(n9082), .Z(n9858) );
  IV U15614 ( .A(n15808), .Z(n9082) );
  XNOR U15615 ( .A(n12979), .B(n11990), .Z(n15808) );
  XNOR U15616 ( .A(n16320), .B(n16321), .Z(n11990) );
  XNOR U15617 ( .A(n12045), .B(n9523), .Z(n16321) );
  XNOR U15618 ( .A(n16322), .B(n15573), .Z(n9523) );
  NOR U15619 ( .A(n14094), .B(n14093), .Z(n16322) );
  XNOR U15620 ( .A(n16323), .B(n16324), .Z(n14093) );
  XOR U15621 ( .A(n16325), .B(n13406), .Z(n12045) );
  XNOR U15622 ( .A(n16326), .B(n15954), .Z(n13406) );
  NOR U15623 ( .A(n14098), .B(n14097), .Z(n16325) );
  XOR U15624 ( .A(n15607), .B(n16327), .Z(n14097) );
  XOR U15625 ( .A(n13285), .B(n16328), .Z(n16320) );
  XOR U15626 ( .A(n13372), .B(n9603), .Z(n16328) );
  XOR U15627 ( .A(n16329), .B(n13411), .Z(n9603) );
  IV U15628 ( .A(n15576), .Z(n13411) );
  XOR U15629 ( .A(n16330), .B(n16331), .Z(n15576) );
  NOR U15630 ( .A(n14090), .B(n14089), .Z(n16329) );
  XNOR U15631 ( .A(n15906), .B(n16332), .Z(n14089) );
  XNOR U15632 ( .A(n16333), .B(n13415), .Z(n13372) );
  XNOR U15633 ( .A(n16334), .B(n15525), .Z(n13415) );
  ANDN U15634 ( .B(n16335), .A(n14085), .Z(n16333) );
  XNOR U15635 ( .A(n16336), .B(n16337), .Z(n14085) );
  XOR U15636 ( .A(n16338), .B(n14256), .Z(n13285) );
  IV U15637 ( .A(n15570), .Z(n14256) );
  XNOR U15638 ( .A(n16339), .B(n16340), .Z(n15570) );
  ANDN U15639 ( .B(n16341), .A(n14100), .Z(n16338) );
  XOR U15640 ( .A(n16342), .B(n16343), .Z(n14100) );
  XOR U15641 ( .A(n16344), .B(n16345), .Z(n12979) );
  XOR U15642 ( .A(n9212), .B(n13550), .Z(n16345) );
  XOR U15643 ( .A(n16346), .B(n16347), .Z(n13550) );
  XOR U15644 ( .A(n16348), .B(n16349), .Z(n14763) );
  XNOR U15645 ( .A(n16350), .B(n15563), .Z(n9212) );
  XOR U15646 ( .A(n14904), .B(n16351), .Z(n14767) );
  XOR U15647 ( .A(n15546), .B(n16352), .Z(n16344) );
  XOR U15648 ( .A(n12324), .B(n12225), .Z(n16352) );
  XNOR U15649 ( .A(n16353), .B(n15566), .Z(n12225) );
  AND U15650 ( .A(n14774), .B(n14775), .Z(n16353) );
  XOR U15651 ( .A(n16354), .B(n16355), .Z(n14774) );
  XNOR U15652 ( .A(n16356), .B(n15555), .Z(n12324) );
  ANDN U15653 ( .B(n15556), .A(n15810), .Z(n16356) );
  XOR U15654 ( .A(n16357), .B(n16252), .Z(n15556) );
  XNOR U15655 ( .A(n16358), .B(n15551), .Z(n15546) );
  XNOR U15656 ( .A(n16360), .B(n15552), .Z(n14770) );
  XNOR U15657 ( .A(n16361), .B(n16362), .Z(n15552) );
  AND U15658 ( .A(n16363), .B(n16359), .Z(n16360) );
  XNOR U15659 ( .A(n16364), .B(n8429), .Z(n2392) );
  XOR U15660 ( .A(n10909), .B(n16365), .Z(n8429) );
  XOR U15661 ( .A(n14078), .B(n12601), .Z(n10909) );
  XOR U15662 ( .A(n16366), .B(n16367), .Z(n12601) );
  XNOR U15663 ( .A(n15786), .B(n10225), .Z(n16367) );
  XOR U15664 ( .A(n16368), .B(n16369), .Z(n10225) );
  ANDN U15665 ( .B(n16370), .A(n16371), .Z(n16368) );
  XNOR U15666 ( .A(n16372), .B(n16373), .Z(n15786) );
  ANDN U15667 ( .B(n16374), .A(n16375), .Z(n16372) );
  XNOR U15668 ( .A(n12372), .B(n16376), .Z(n16366) );
  XOR U15669 ( .A(n13591), .B(n15812), .Z(n16376) );
  XNOR U15670 ( .A(n16377), .B(n16378), .Z(n15812) );
  AND U15671 ( .A(n16379), .B(n16380), .Z(n16377) );
  XNOR U15672 ( .A(n16381), .B(n16382), .Z(n13591) );
  NOR U15673 ( .A(n16383), .B(n16384), .Z(n16381) );
  XNOR U15674 ( .A(n16385), .B(n16386), .Z(n12372) );
  AND U15675 ( .A(n16387), .B(n16388), .Z(n16385) );
  XOR U15676 ( .A(n16389), .B(n16390), .Z(n14078) );
  XOR U15677 ( .A(n11374), .B(n13390), .Z(n16390) );
  XOR U15678 ( .A(n16391), .B(n16392), .Z(n13390) );
  ANDN U15679 ( .B(n16393), .A(n16394), .Z(n16391) );
  XOR U15680 ( .A(n16395), .B(n16396), .Z(n11374) );
  ANDN U15681 ( .B(n16397), .A(n16398), .Z(n16395) );
  XOR U15682 ( .A(n10021), .B(n16399), .Z(n16389) );
  XNOR U15683 ( .A(n16400), .B(n14126), .Z(n16399) );
  XNOR U15684 ( .A(n16401), .B(n16402), .Z(n14126) );
  ANDN U15685 ( .B(n16403), .A(n16404), .Z(n16401) );
  XOR U15686 ( .A(n16405), .B(n16406), .Z(n10021) );
  AND U15687 ( .A(n16407), .B(n16408), .Z(n16405) );
  ANDN U15688 ( .B(n12112), .A(n8477), .Z(n16364) );
  XOR U15689 ( .A(n10118), .B(n16409), .Z(n8477) );
  XOR U15690 ( .A(n15369), .B(n13659), .Z(n10118) );
  XOR U15691 ( .A(n16410), .B(n16411), .Z(n13659) );
  XOR U15692 ( .A(n14429), .B(n12883), .Z(n16411) );
  XOR U15693 ( .A(n16412), .B(n15526), .Z(n12883) );
  ANDN U15694 ( .B(n14608), .A(n13176), .Z(n16412) );
  XNOR U15695 ( .A(n16413), .B(n16414), .Z(n13176) );
  ANDN U15696 ( .B(n13168), .A(n14610), .Z(n16415) );
  XNOR U15697 ( .A(n16416), .B(n16417), .Z(n13168) );
  XNOR U15698 ( .A(n13017), .B(n16418), .Z(n16410) );
  XNOR U15699 ( .A(n16419), .B(n16420), .Z(n16418) );
  XNOR U15700 ( .A(n16421), .B(n16422), .Z(n13017) );
  ANDN U15701 ( .B(n14619), .A(n13325), .Z(n16421) );
  XNOR U15702 ( .A(n16423), .B(n16252), .Z(n13325) );
  XOR U15703 ( .A(n16424), .B(n16425), .Z(n15369) );
  XNOR U15704 ( .A(n9686), .B(n16426), .Z(n16425) );
  XNOR U15705 ( .A(n16427), .B(n15510), .Z(n9686) );
  ANDN U15706 ( .B(n16428), .A(n16429), .Z(n16427) );
  XNOR U15707 ( .A(n10886), .B(n16430), .Z(n16424) );
  XOR U15708 ( .A(n16431), .B(n10913), .Z(n16430) );
  XNOR U15709 ( .A(n16432), .B(n15507), .Z(n10913) );
  AND U15710 ( .A(n16433), .B(n16434), .Z(n16432) );
  XOR U15711 ( .A(n16435), .B(n15493), .Z(n10886) );
  NOR U15712 ( .A(n16436), .B(n16437), .Z(n16435) );
  XOR U15713 ( .A(n15430), .B(n11021), .Z(n12112) );
  XNOR U15714 ( .A(n16438), .B(n16439), .Z(n15430) );
  NOR U15715 ( .A(n14578), .B(n14577), .Z(n16438) );
  XNOR U15716 ( .A(n16440), .B(n8435), .Z(n6253) );
  XOR U15717 ( .A(n16441), .B(n16442), .Z(n8435) );
  NOR U15718 ( .A(n8481), .B(n8480), .Z(n16440) );
  XOR U15719 ( .A(n12145), .B(n12895), .Z(n8480) );
  XNOR U15720 ( .A(n16443), .B(n14122), .Z(n12895) );
  AND U15721 ( .A(n16029), .B(n15366), .Z(n16443) );
  XOR U15722 ( .A(n16444), .B(n15603), .Z(n15366) );
  XOR U15723 ( .A(n13909), .B(n16445), .Z(n12145) );
  XOR U15724 ( .A(n16446), .B(n16447), .Z(n13909) );
  XNOR U15725 ( .A(n12928), .B(n13224), .Z(n16447) );
  XOR U15726 ( .A(n16448), .B(n15360), .Z(n13224) );
  IV U15727 ( .A(n14110), .Z(n15360) );
  XNOR U15728 ( .A(n16449), .B(n15529), .Z(n14110) );
  ANDN U15729 ( .B(n12904), .A(n12902), .Z(n16448) );
  XNOR U15730 ( .A(n16450), .B(n16451), .Z(n12902) );
  XOR U15731 ( .A(n16452), .B(n16453), .Z(n12904) );
  XNOR U15732 ( .A(n16454), .B(n14113), .Z(n12928) );
  XNOR U15733 ( .A(n16455), .B(n16456), .Z(n14113) );
  ANDN U15734 ( .B(n12898), .A(n12899), .Z(n16454) );
  XNOR U15735 ( .A(n16457), .B(n16458), .Z(n12899) );
  XNOR U15736 ( .A(n16459), .B(n16460), .Z(n12898) );
  XOR U15737 ( .A(n11051), .B(n16461), .Z(n16446) );
  XOR U15738 ( .A(n11694), .B(n13287), .Z(n16461) );
  XOR U15739 ( .A(n16462), .B(n15358), .Z(n13287) );
  IV U15740 ( .A(n15003), .Z(n15358) );
  XNOR U15741 ( .A(n16463), .B(n16062), .Z(n15003) );
  AND U15742 ( .A(n15004), .B(n16019), .Z(n16462) );
  IV U15743 ( .A(n15816), .Z(n16019) );
  XNOR U15744 ( .A(n16464), .B(n16465), .Z(n15816) );
  XOR U15745 ( .A(n16466), .B(n14924), .Z(n15004) );
  XOR U15746 ( .A(n16467), .B(n15364), .Z(n11694) );
  IV U15747 ( .A(n14118), .Z(n15364) );
  XOR U15748 ( .A(n16468), .B(n16469), .Z(n14118) );
  NOR U15749 ( .A(n12906), .B(n12907), .Z(n16467) );
  XOR U15750 ( .A(n16470), .B(n15856), .Z(n12907) );
  XNOR U15751 ( .A(n16471), .B(n16472), .Z(n12906) );
  XOR U15752 ( .A(n16473), .B(n15367), .Z(n11051) );
  IV U15753 ( .A(n14121), .Z(n15367) );
  XOR U15754 ( .A(n16474), .B(n15122), .Z(n14121) );
  ANDN U15755 ( .B(n14122), .A(n16029), .Z(n16473) );
  XNOR U15756 ( .A(n16475), .B(n16476), .Z(n16029) );
  XNOR U15757 ( .A(n16477), .B(n16478), .Z(n14122) );
  XNOR U15758 ( .A(n16479), .B(n12069), .Z(n8481) );
  XNOR U15759 ( .A(n16126), .B(n16480), .Z(n12069) );
  XOR U15760 ( .A(n16481), .B(n16482), .Z(n16126) );
  XNOR U15761 ( .A(n9394), .B(n16483), .Z(n16482) );
  XOR U15762 ( .A(n16484), .B(n14720), .Z(n9394) );
  AND U15763 ( .A(n16485), .B(n16486), .Z(n16484) );
  XOR U15764 ( .A(n16487), .B(n16488), .Z(n16481) );
  XNOR U15765 ( .A(n11248), .B(n13900), .Z(n16488) );
  XNOR U15766 ( .A(n16489), .B(n14737), .Z(n13900) );
  AND U15767 ( .A(n16490), .B(n16491), .Z(n16489) );
  XOR U15768 ( .A(n16492), .B(n14724), .Z(n11248) );
  AND U15769 ( .A(n16493), .B(n16494), .Z(n16492) );
  XOR U15770 ( .A(n16495), .B(n16496), .Z(n8345) );
  XOR U15771 ( .A(n3811), .B(n5121), .Z(n16496) );
  XOR U15772 ( .A(n16497), .B(n9760), .Z(n5121) );
  XNOR U15773 ( .A(n16498), .B(n9810), .Z(n9760) );
  XOR U15774 ( .A(n15684), .B(n16499), .Z(n9810) );
  XOR U15775 ( .A(n16500), .B(n16501), .Z(n15684) );
  XNOR U15776 ( .A(n11651), .B(n12709), .Z(n16501) );
  XNOR U15777 ( .A(n16502), .B(n13265), .Z(n12709) );
  NOR U15778 ( .A(n13266), .B(n14847), .Z(n16502) );
  XNOR U15779 ( .A(n16503), .B(n13255), .Z(n11651) );
  ANDN U15780 ( .B(n13256), .A(n14844), .Z(n16503) );
  XOR U15781 ( .A(n11732), .B(n16504), .Z(n16500) );
  XOR U15782 ( .A(n10593), .B(n11410), .Z(n16504) );
  XOR U15783 ( .A(n16505), .B(n13252), .Z(n11410) );
  NOR U15784 ( .A(n13251), .B(n14836), .Z(n16505) );
  XOR U15785 ( .A(n16506), .B(n16507), .Z(n10593) );
  NOR U15786 ( .A(n16508), .B(n14840), .Z(n16506) );
  XOR U15787 ( .A(n16509), .B(n16510), .Z(n11732) );
  NOR U15788 ( .A(n13261), .B(n14833), .Z(n16509) );
  ANDN U15789 ( .B(n12032), .A(n12033), .Z(n16497) );
  XNOR U15790 ( .A(n9393), .B(n16487), .Z(n12033) );
  XNOR U15791 ( .A(n16511), .B(n14729), .Z(n16487) );
  AND U15792 ( .A(n16512), .B(n16513), .Z(n16511) );
  IV U15793 ( .A(n11247), .Z(n9393) );
  XOR U15794 ( .A(n15426), .B(n11021), .Z(n12032) );
  IV U15795 ( .A(n12344), .Z(n11021) );
  XOR U15796 ( .A(n11677), .B(n13082), .Z(n12344) );
  XNOR U15797 ( .A(n16514), .B(n16515), .Z(n13082) );
  XNOR U15798 ( .A(n12735), .B(n11294), .Z(n16515) );
  XOR U15799 ( .A(n16516), .B(n16517), .Z(n11294) );
  ANDN U15800 ( .B(n15438), .A(n15279), .Z(n16516) );
  XNOR U15801 ( .A(n16518), .B(n16519), .Z(n15279) );
  XNOR U15802 ( .A(n16520), .B(n16521), .Z(n12735) );
  ANDN U15803 ( .B(n15436), .A(n15275), .Z(n16520) );
  XNOR U15804 ( .A(n16522), .B(n16523), .Z(n15275) );
  XOR U15805 ( .A(n16524), .B(n16525), .Z(n16514) );
  XOR U15806 ( .A(n10230), .B(n11005), .Z(n16525) );
  XNOR U15807 ( .A(n16526), .B(n16527), .Z(n11005) );
  ANDN U15808 ( .B(n15441), .A(n15271), .Z(n16526) );
  XOR U15809 ( .A(n16528), .B(n15639), .Z(n15271) );
  XOR U15810 ( .A(n16529), .B(n16530), .Z(n10230) );
  AND U15811 ( .A(n15262), .B(n15443), .Z(n16529) );
  XNOR U15812 ( .A(n16531), .B(n16532), .Z(n15262) );
  XOR U15813 ( .A(n16533), .B(n16534), .Z(n11677) );
  XOR U15814 ( .A(n15139), .B(n12727), .Z(n16534) );
  XOR U15815 ( .A(n16535), .B(n15146), .Z(n12727) );
  NOR U15816 ( .A(n15145), .B(n15421), .Z(n16535) );
  XOR U15817 ( .A(n16536), .B(n16537), .Z(n15139) );
  AND U15818 ( .A(n14581), .B(n15428), .Z(n16536) );
  XNOR U15819 ( .A(n16538), .B(n16539), .Z(n14581) );
  XNOR U15820 ( .A(n12456), .B(n16540), .Z(n16533) );
  XOR U15821 ( .A(n9489), .B(n11771), .Z(n16540) );
  XOR U15822 ( .A(n16541), .B(n16542), .Z(n11771) );
  XOR U15823 ( .A(n16543), .B(n16544), .Z(n14577) );
  XOR U15824 ( .A(n16545), .B(n15149), .Z(n9489) );
  XNOR U15825 ( .A(n16546), .B(n16478), .Z(n14585) );
  XOR U15826 ( .A(n16547), .B(n16548), .Z(n15150) );
  XOR U15827 ( .A(n16549), .B(n15156), .Z(n12456) );
  ANDN U15828 ( .B(n14572), .A(n15155), .Z(n16549) );
  XNOR U15829 ( .A(n15132), .B(n16550), .Z(n15155) );
  XNOR U15830 ( .A(n16551), .B(n16552), .Z(n14572) );
  XNOR U15831 ( .A(n16553), .B(n15145), .Z(n15426) );
  XOR U15832 ( .A(n16554), .B(n16555), .Z(n15145) );
  ANDN U15833 ( .B(n15421), .A(n15422), .Z(n16553) );
  XNOR U15834 ( .A(n16556), .B(n16557), .Z(n15421) );
  XNOR U15835 ( .A(n16558), .B(n12103), .Z(n3811) );
  IV U15836 ( .A(n8404), .Z(n12103) );
  XOR U15837 ( .A(n16420), .B(n12884), .Z(n8404) );
  XNOR U15838 ( .A(n16559), .B(n15521), .Z(n16420) );
  AND U15839 ( .A(n13172), .B(n14614), .Z(n16559) );
  XOR U15840 ( .A(n16560), .B(n16062), .Z(n13172) );
  AND U15841 ( .A(n12024), .B(n12025), .Z(n16558) );
  XOR U15842 ( .A(n15065), .B(n11825), .Z(n12025) );
  XOR U15843 ( .A(n13417), .B(n12368), .Z(n11825) );
  XOR U15844 ( .A(n16561), .B(n16562), .Z(n12368) );
  XNOR U15845 ( .A(n14880), .B(n15391), .Z(n16562) );
  XOR U15846 ( .A(n16563), .B(n16564), .Z(n15391) );
  XNOR U15847 ( .A(n16567), .B(n16394), .Z(n14880) );
  NOR U15848 ( .A(n16568), .B(n16569), .Z(n16567) );
  XOR U15849 ( .A(n14929), .B(n16570), .Z(n16561) );
  XOR U15850 ( .A(n13074), .B(n12209), .Z(n16570) );
  XNOR U15851 ( .A(n16571), .B(n16404), .Z(n12209) );
  ANDN U15852 ( .B(n16572), .A(n16573), .Z(n16571) );
  XNOR U15853 ( .A(n16574), .B(n16398), .Z(n13074) );
  ANDN U15854 ( .B(n16575), .A(n16576), .Z(n16574) );
  XOR U15855 ( .A(n16577), .B(n16407), .Z(n14929) );
  XOR U15856 ( .A(n16580), .B(n16581), .Z(n13417) );
  XNOR U15857 ( .A(n9893), .B(n12968), .Z(n16581) );
  XNOR U15858 ( .A(n16582), .B(n14238), .Z(n12968) );
  NOR U15859 ( .A(n15059), .B(n15058), .Z(n16582) );
  XOR U15860 ( .A(n16583), .B(n14244), .Z(n9893) );
  XOR U15861 ( .A(n16584), .B(n16585), .Z(n16580) );
  XNOR U15862 ( .A(n11243), .B(n13422), .Z(n16585) );
  XOR U15863 ( .A(n16586), .B(n14234), .Z(n13422) );
  ANDN U15864 ( .B(n16587), .A(n16588), .Z(n16586) );
  XOR U15865 ( .A(n16589), .B(n16590), .Z(n11243) );
  ANDN U15866 ( .B(n15061), .A(n15062), .Z(n16589) );
  XNOR U15867 ( .A(n16591), .B(n16588), .Z(n15065) );
  ANDN U15868 ( .B(n14232), .A(n16587), .Z(n16591) );
  XOR U15869 ( .A(n10266), .B(n16592), .Z(n12024) );
  IV U15870 ( .A(n16442), .Z(n10266) );
  XOR U15871 ( .A(n5805), .B(n16593), .Z(n16495) );
  XOR U15872 ( .A(n1746), .B(n12093), .Z(n16593) );
  XNOR U15873 ( .A(n16594), .B(n8415), .Z(n12093) );
  XNOR U15874 ( .A(n16595), .B(n11166), .Z(n8415) );
  XNOR U15875 ( .A(n16596), .B(n16597), .Z(n11166) );
  AND U15876 ( .A(n12022), .B(n12021), .Z(n16594) );
  IV U15877 ( .A(n12105), .Z(n12021) );
  XOR U15878 ( .A(n11257), .B(n16598), .Z(n12105) );
  XOR U15879 ( .A(n16599), .B(n16600), .Z(n13246) );
  XNOR U15880 ( .A(n9599), .B(n10099), .Z(n16600) );
  XOR U15881 ( .A(n16601), .B(n13431), .Z(n10099) );
  XNOR U15882 ( .A(n16602), .B(n16603), .Z(n13431) );
  ANDN U15883 ( .B(n16604), .A(n13430), .Z(n16601) );
  XNOR U15884 ( .A(n16605), .B(n13436), .Z(n9599) );
  XOR U15885 ( .A(n16606), .B(n16340), .Z(n13436) );
  AND U15886 ( .A(n16607), .B(n16608), .Z(n16605) );
  XOR U15887 ( .A(n9352), .B(n16609), .Z(n16599) );
  XOR U15888 ( .A(n13423), .B(n13179), .Z(n16609) );
  XNOR U15889 ( .A(n16610), .B(n14827), .Z(n13179) );
  XOR U15890 ( .A(n16611), .B(n16612), .Z(n14827) );
  ANDN U15891 ( .B(n16613), .A(n16614), .Z(n16610) );
  XOR U15892 ( .A(n16615), .B(n13441), .Z(n13423) );
  XNOR U15893 ( .A(n16617), .B(n14440), .Z(n9352) );
  XNOR U15894 ( .A(n16618), .B(n16057), .Z(n14440) );
  XNOR U15895 ( .A(n16620), .B(n16621), .Z(n14009) );
  XOR U15896 ( .A(n11381), .B(n12317), .Z(n16621) );
  XOR U15897 ( .A(n16622), .B(n15110), .Z(n12317) );
  NOR U15898 ( .A(n16623), .B(n16624), .Z(n16622) );
  XOR U15899 ( .A(n16625), .B(n15114), .Z(n11381) );
  ANDN U15900 ( .B(n16626), .A(n16627), .Z(n16625) );
  XOR U15901 ( .A(n10574), .B(n16628), .Z(n16620) );
  XOR U15902 ( .A(n10295), .B(n11744), .Z(n16628) );
  ANDN U15903 ( .B(n16630), .A(n16631), .Z(n16629) );
  XNOR U15904 ( .A(n16632), .B(n16633), .Z(n10295) );
  AND U15905 ( .A(n16634), .B(n16635), .Z(n16632) );
  NOR U15906 ( .A(n16637), .B(n16638), .Z(n16636) );
  XOR U15907 ( .A(n16639), .B(n16640), .Z(n12022) );
  XOR U15908 ( .A(n16641), .B(n8408), .Z(n1746) );
  XOR U15909 ( .A(n16162), .B(n11412), .Z(n8408) );
  IV U15910 ( .A(n10553), .Z(n11412) );
  XOR U15911 ( .A(n16445), .B(n14975), .Z(n10553) );
  XOR U15912 ( .A(n16642), .B(n16643), .Z(n14975) );
  XNOR U15913 ( .A(n11996), .B(n12763), .Z(n16643) );
  XOR U15914 ( .A(n16644), .B(n15886), .Z(n12763) );
  AND U15915 ( .A(n16645), .B(n16646), .Z(n16644) );
  XNOR U15916 ( .A(n16647), .B(n15868), .Z(n11996) );
  AND U15917 ( .A(n16648), .B(n16649), .Z(n16647) );
  XOR U15918 ( .A(n11927), .B(n16650), .Z(n16642) );
  XNOR U15919 ( .A(n15862), .B(n13684), .Z(n16650) );
  XNOR U15920 ( .A(n16651), .B(n15878), .Z(n13684) );
  ANDN U15921 ( .B(n16652), .A(n15877), .Z(n16651) );
  XNOR U15922 ( .A(n16653), .B(n15872), .Z(n15862) );
  ANDN U15923 ( .B(n15873), .A(n16654), .Z(n16653) );
  XNOR U15924 ( .A(n16655), .B(n15882), .Z(n11927) );
  ANDN U15925 ( .B(n16656), .A(n15881), .Z(n16655) );
  XOR U15926 ( .A(n16657), .B(n16658), .Z(n16445) );
  XNOR U15927 ( .A(n9693), .B(n11788), .Z(n16658) );
  XNOR U15928 ( .A(n16659), .B(n13308), .Z(n11788) );
  NOR U15929 ( .A(n16660), .B(n13307), .Z(n16659) );
  XOR U15930 ( .A(n16661), .B(n16662), .Z(n9693) );
  XNOR U15931 ( .A(n16663), .B(n16664), .Z(n14677) );
  XOR U15932 ( .A(n9910), .B(n16665), .Z(n16657) );
  XOR U15933 ( .A(n10655), .B(n10387), .Z(n16665) );
  XOR U15934 ( .A(n16666), .B(n13304), .Z(n10387) );
  ANDN U15935 ( .B(n16156), .A(n16157), .Z(n16666) );
  XNOR U15936 ( .A(n14944), .B(n16667), .Z(n16157) );
  IV U15937 ( .A(n13303), .Z(n16156) );
  XOR U15938 ( .A(n16668), .B(n16669), .Z(n13303) );
  XOR U15939 ( .A(n16670), .B(n13300), .Z(n10655) );
  NOR U15940 ( .A(n16164), .B(n13299), .Z(n16670) );
  XOR U15941 ( .A(n16671), .B(n16672), .Z(n13299) );
  IV U15942 ( .A(n14681), .Z(n16164) );
  XOR U15943 ( .A(n16673), .B(n16674), .Z(n14681) );
  XOR U15944 ( .A(n16675), .B(n13295), .Z(n9910) );
  NOR U15945 ( .A(n13294), .B(n14670), .Z(n16675) );
  XOR U15946 ( .A(n16676), .B(n16677), .Z(n14670) );
  XNOR U15947 ( .A(n16678), .B(n16014), .Z(n13294) );
  XNOR U15948 ( .A(n16679), .B(n13307), .Z(n16162) );
  XNOR U15949 ( .A(n16680), .B(n15987), .Z(n13307) );
  AND U15950 ( .A(n14675), .B(n16660), .Z(n16679) );
  IV U15951 ( .A(n14674), .Z(n16660) );
  XOR U15952 ( .A(n16681), .B(n16682), .Z(n14674) );
  ANDN U15953 ( .B(n12029), .A(n12030), .Z(n16641) );
  XNOR U15954 ( .A(n16683), .B(n10270), .Z(n12030) );
  XNOR U15955 ( .A(n15198), .B(n12602), .Z(n10270) );
  XNOR U15956 ( .A(n16684), .B(n16685), .Z(n12602) );
  XNOR U15957 ( .A(n11816), .B(n11312), .Z(n16685) );
  XNOR U15958 ( .A(n16686), .B(n12821), .Z(n11312) );
  XNOR U15959 ( .A(n16687), .B(n16688), .Z(n12821) );
  AND U15960 ( .A(n16244), .B(n16689), .Z(n16686) );
  XNOR U15961 ( .A(n16690), .B(n15947), .Z(n11816) );
  XOR U15962 ( .A(n16691), .B(n16692), .Z(n15947) );
  AND U15963 ( .A(n16693), .B(n16694), .Z(n16690) );
  XOR U15964 ( .A(n10731), .B(n16695), .Z(n16684) );
  XOR U15965 ( .A(n16230), .B(n13320), .Z(n16695) );
  XOR U15966 ( .A(n16696), .B(n14323), .Z(n13320) );
  XOR U15967 ( .A(n16697), .B(n16698), .Z(n14323) );
  AND U15968 ( .A(n16699), .B(n16240), .Z(n16696) );
  XOR U15969 ( .A(n16700), .B(n12818), .Z(n16230) );
  XOR U15970 ( .A(n16701), .B(n16702), .Z(n12818) );
  AND U15971 ( .A(n16703), .B(n16704), .Z(n16700) );
  XNOR U15972 ( .A(n16705), .B(n12811), .Z(n10731) );
  XNOR U15973 ( .A(n16706), .B(n16707), .Z(n12811) );
  AND U15974 ( .A(n16708), .B(n16242), .Z(n16705) );
  XOR U15975 ( .A(n16709), .B(n16710), .Z(n15198) );
  XNOR U15976 ( .A(n16711), .B(n13184), .Z(n16710) );
  XNOR U15977 ( .A(n16712), .B(n16713), .Z(n13184) );
  ANDN U15978 ( .B(n16714), .A(n16715), .Z(n16712) );
  XOR U15979 ( .A(n12694), .B(n16716), .Z(n16709) );
  XOR U15980 ( .A(n11781), .B(n12654), .Z(n16716) );
  XOR U15981 ( .A(n16717), .B(n16718), .Z(n12654) );
  ANDN U15982 ( .B(n15924), .A(n16719), .Z(n16717) );
  XNOR U15983 ( .A(n16720), .B(n16721), .Z(n11781) );
  AND U15984 ( .A(n15928), .B(n16722), .Z(n16720) );
  XNOR U15985 ( .A(n16723), .B(n16724), .Z(n12694) );
  AND U15986 ( .A(n16725), .B(n15941), .Z(n16723) );
  XOR U15987 ( .A(n15779), .B(n9661), .Z(n12029) );
  XNOR U15988 ( .A(n14251), .B(n12977), .Z(n9661) );
  XNOR U15989 ( .A(n16726), .B(n16727), .Z(n12977) );
  XNOR U15990 ( .A(n10105), .B(n14135), .Z(n16727) );
  XOR U15991 ( .A(n16728), .B(n16729), .Z(n14135) );
  AND U15992 ( .A(n15774), .B(n15772), .Z(n16728) );
  XNOR U15993 ( .A(n16730), .B(n14866), .Z(n10105) );
  AND U15994 ( .A(n15784), .B(n15785), .Z(n16730) );
  XOR U15995 ( .A(n12913), .B(n16731), .Z(n16726) );
  XNOR U15996 ( .A(n9171), .B(n11980), .Z(n16731) );
  XOR U15997 ( .A(n16732), .B(n14862), .Z(n11980) );
  ANDN U15998 ( .B(n15777), .A(n15776), .Z(n16732) );
  XNOR U15999 ( .A(n16733), .B(n14872), .Z(n9171) );
  ANDN U16000 ( .B(n15781), .A(n15782), .Z(n16733) );
  XNOR U16001 ( .A(n16734), .B(n14875), .Z(n12913) );
  AND U16002 ( .A(n16735), .B(n16736), .Z(n16734) );
  XOR U16003 ( .A(n16737), .B(n16738), .Z(n14251) );
  XNOR U16004 ( .A(n9928), .B(n13510), .Z(n16738) );
  XOR U16005 ( .A(n16739), .B(n14142), .Z(n13510) );
  ANDN U16006 ( .B(n14143), .A(n15765), .Z(n16739) );
  XNOR U16007 ( .A(n16268), .B(n16740), .Z(n14143) );
  XNOR U16008 ( .A(n16741), .B(n16742), .Z(n9928) );
  ANDN U16009 ( .B(n15753), .A(n15754), .Z(n16741) );
  XNOR U16010 ( .A(n9113), .B(n16743), .Z(n16737) );
  XOR U16011 ( .A(n9943), .B(n13019), .Z(n16743) );
  XOR U16012 ( .A(n16744), .B(n15449), .Z(n13019) );
  AND U16013 ( .A(n15762), .B(n15450), .Z(n16744) );
  XNOR U16014 ( .A(n16745), .B(n16746), .Z(n15450) );
  XOR U16015 ( .A(n16747), .B(n14148), .Z(n9943) );
  ANDN U16016 ( .B(n14149), .A(n15767), .Z(n16747) );
  XNOR U16017 ( .A(n16748), .B(n16749), .Z(n14149) );
  XNOR U16018 ( .A(n16750), .B(n14153), .Z(n9113) );
  NOR U16019 ( .A(n14152), .B(n15757), .Z(n16750) );
  XNOR U16020 ( .A(n16751), .B(n16752), .Z(n14152) );
  XNOR U16021 ( .A(n16753), .B(n16736), .Z(n15779) );
  NOR U16022 ( .A(n16735), .B(n14874), .Z(n16753) );
  XOR U16023 ( .A(n16754), .B(n8418), .Z(n5805) );
  IV U16024 ( .A(n12100), .Z(n8418) );
  XNOR U16025 ( .A(n15023), .B(n10251), .Z(n12100) );
  XOR U16026 ( .A(n11658), .B(n13222), .Z(n10251) );
  XOR U16027 ( .A(n16755), .B(n16756), .Z(n13222) );
  XNOR U16028 ( .A(n10934), .B(n10540), .Z(n16756) );
  XNOR U16029 ( .A(n16757), .B(n16253), .Z(n10540) );
  AND U16030 ( .A(n15026), .B(n15028), .Z(n16757) );
  XNOR U16031 ( .A(n16758), .B(n16759), .Z(n15028) );
  XOR U16032 ( .A(n16760), .B(n16270), .Z(n10934) );
  AND U16033 ( .A(n15017), .B(n16761), .Z(n16760) );
  XNOR U16034 ( .A(n12864), .B(n16763), .Z(n16755) );
  XOR U16035 ( .A(n15948), .B(n9990), .Z(n16763) );
  XNOR U16036 ( .A(n16764), .B(n16257), .Z(n9990) );
  AND U16037 ( .A(n15020), .B(n16765), .Z(n16764) );
  XNOR U16038 ( .A(n16766), .B(n16767), .Z(n15020) );
  XOR U16039 ( .A(n16768), .B(n16769), .Z(n15948) );
  ANDN U16040 ( .B(n16246), .A(n15478), .Z(n16768) );
  XNOR U16041 ( .A(n16770), .B(n16453), .Z(n15478) );
  XNOR U16042 ( .A(n16771), .B(n16265), .Z(n12864) );
  ANDN U16043 ( .B(n16772), .A(n15474), .Z(n16771) );
  XOR U16044 ( .A(n16773), .B(n16774), .Z(n11658) );
  XNOR U16045 ( .A(n12632), .B(n11012), .Z(n16774) );
  XNOR U16046 ( .A(n16775), .B(n15955), .Z(n11012) );
  IV U16047 ( .A(n13756), .Z(n15955) );
  XOR U16048 ( .A(n16776), .B(n16021), .Z(n13756) );
  ANDN U16049 ( .B(n15956), .A(n13237), .Z(n16775) );
  XNOR U16050 ( .A(n16777), .B(n13762), .Z(n12632) );
  XNOR U16051 ( .A(n16778), .B(n16779), .Z(n13762) );
  AND U16052 ( .A(n14851), .B(n16780), .Z(n16777) );
  XOR U16053 ( .A(n14317), .B(n16781), .Z(n16773) );
  XOR U16054 ( .A(n10918), .B(n11568), .Z(n16781) );
  XOR U16055 ( .A(n16782), .B(n13765), .Z(n11568) );
  XOR U16056 ( .A(n16783), .B(n16784), .Z(n13765) );
  AND U16057 ( .A(n15966), .B(n16785), .Z(n16782) );
  XOR U16058 ( .A(n16786), .B(n13752), .Z(n10918) );
  XOR U16059 ( .A(n16787), .B(n16788), .Z(n13752) );
  ANDN U16060 ( .B(n15963), .A(n16789), .Z(n16786) );
  XNOR U16061 ( .A(n16790), .B(n13759), .Z(n14317) );
  XNOR U16062 ( .A(n16791), .B(n16792), .Z(n13759) );
  ANDN U16063 ( .B(n15969), .A(n13241), .Z(n16790) );
  XNOR U16064 ( .A(n16793), .B(n16772), .Z(n15023) );
  AND U16065 ( .A(n15474), .B(n16264), .Z(n16793) );
  IV U16066 ( .A(n15476), .Z(n16264) );
  XNOR U16067 ( .A(n16794), .B(n16795), .Z(n15476) );
  XOR U16068 ( .A(n16796), .B(n16797), .Z(n15474) );
  XOR U16069 ( .A(n16798), .B(n12101), .Z(n12026) );
  XOR U16070 ( .A(n11649), .B(n14221), .Z(n12101) );
  XNOR U16071 ( .A(n16799), .B(n14186), .Z(n14221) );
  AND U16072 ( .A(n16800), .B(n16801), .Z(n16799) );
  AND U16073 ( .A(n8417), .B(n14464), .Z(n16798) );
  XOR U16074 ( .A(n16311), .B(n12366), .Z(n14464) );
  XNOR U16075 ( .A(n11866), .B(n16802), .Z(n12366) );
  XOR U16076 ( .A(n16803), .B(n16804), .Z(n11866) );
  XOR U16077 ( .A(n10877), .B(n11417), .Z(n16804) );
  XOR U16078 ( .A(n16805), .B(n16806), .Z(n11417) );
  IV U16079 ( .A(n16309), .Z(n14752) );
  XOR U16080 ( .A(n16807), .B(n16808), .Z(n16309) );
  XOR U16081 ( .A(n16809), .B(n16810), .Z(n10877) );
  NOR U16082 ( .A(n14745), .B(n16315), .Z(n16809) );
  XNOR U16083 ( .A(n16811), .B(n16812), .Z(n14745) );
  XOR U16084 ( .A(n11283), .B(n16813), .Z(n16803) );
  XNOR U16085 ( .A(n9504), .B(n16814), .Z(n16813) );
  XNOR U16086 ( .A(n16815), .B(n16816), .Z(n9504) );
  ANDN U16087 ( .B(n14741), .A(n16313), .Z(n16815) );
  XNOR U16088 ( .A(n16817), .B(n16818), .Z(n14741) );
  XNOR U16089 ( .A(n16819), .B(n16820), .Z(n11283) );
  ANDN U16090 ( .B(n16821), .A(n16288), .Z(n16819) );
  XNOR U16091 ( .A(n16822), .B(n16823), .Z(n16311) );
  ANDN U16092 ( .B(n16288), .A(n16289), .Z(n16822) );
  XNOR U16093 ( .A(n16824), .B(n16612), .Z(n16288) );
  XNOR U16094 ( .A(n14059), .B(n13912), .Z(n8417) );
  XOR U16095 ( .A(n14250), .B(n16825), .Z(n13912) );
  XOR U16096 ( .A(n16826), .B(n16827), .Z(n14250) );
  XNOR U16097 ( .A(n12443), .B(n14626), .Z(n16827) );
  XOR U16098 ( .A(n16828), .B(n14636), .Z(n14626) );
  ANDN U16099 ( .B(n14061), .A(n14062), .Z(n16828) );
  XNOR U16100 ( .A(n16829), .B(n16830), .Z(n14061) );
  XOR U16101 ( .A(n16831), .B(n15074), .Z(n12443) );
  AND U16102 ( .A(n14072), .B(n15075), .Z(n16831) );
  XOR U16103 ( .A(n16832), .B(n13991), .Z(n15075) );
  XNOR U16104 ( .A(n11298), .B(n16833), .Z(n16826) );
  XOR U16105 ( .A(n11036), .B(n12168), .Z(n16833) );
  XOR U16106 ( .A(n16834), .B(n16835), .Z(n12168) );
  ANDN U16107 ( .B(n14068), .A(n14066), .Z(n16834) );
  XNOR U16108 ( .A(n16836), .B(n16837), .Z(n11036) );
  ANDN U16109 ( .B(n14074), .A(n14075), .Z(n16836) );
  XOR U16110 ( .A(n16838), .B(n14639), .Z(n11298) );
  ANDN U16111 ( .B(n14640), .A(n16839), .Z(n16838) );
  XNOR U16112 ( .A(n16840), .B(n14640), .Z(n14059) );
  XNOR U16113 ( .A(n16841), .B(n16842), .Z(n14640) );
  ANDN U16114 ( .B(n16839), .A(n16843), .Z(n16840) );
  XOR U16115 ( .A(n16844), .B(n2598), .Z(out[0]) );
  XNOR U16116 ( .A(n2200), .B(n10452), .Z(n2598) );
  XNOR U16117 ( .A(n16845), .B(n8556), .Z(n10452) );
  ANDN U16118 ( .B(n10304), .A(n10486), .Z(n16845) );
  XNOR U16119 ( .A(n10544), .B(n16846), .Z(n10304) );
  XOR U16120 ( .A(n12628), .B(n15054), .Z(n10544) );
  XOR U16121 ( .A(n16847), .B(n16848), .Z(n15054) );
  XNOR U16122 ( .A(n11001), .B(n12367), .Z(n16848) );
  XOR U16123 ( .A(n16849), .B(n16572), .Z(n12367) );
  AND U16124 ( .A(n16573), .B(n16402), .Z(n16849) );
  XNOR U16125 ( .A(n16850), .B(n16569), .Z(n11001) );
  ANDN U16126 ( .B(n16568), .A(n16392), .Z(n16850) );
  XOR U16127 ( .A(n10255), .B(n16851), .Z(n16847) );
  XNOR U16128 ( .A(n11995), .B(n10729), .Z(n16851) );
  XOR U16129 ( .A(n16852), .B(n16853), .Z(n10729) );
  AND U16130 ( .A(n16576), .B(n16396), .Z(n16852) );
  IV U16131 ( .A(n16854), .Z(n16396) );
  XNOR U16132 ( .A(n16855), .B(n16566), .Z(n11995) );
  AND U16133 ( .A(n16565), .B(n16856), .Z(n16855) );
  XOR U16134 ( .A(n16857), .B(n16579), .Z(n10255) );
  NOR U16135 ( .A(n16578), .B(n16406), .Z(n16857) );
  XOR U16136 ( .A(n16858), .B(n16859), .Z(n12628) );
  XNOR U16137 ( .A(n11508), .B(n14052), .Z(n16859) );
  XNOR U16138 ( .A(n16860), .B(n16861), .Z(n14052) );
  ANDN U16139 ( .B(n16373), .A(n16862), .Z(n16860) );
  XNOR U16140 ( .A(n16863), .B(n16864), .Z(n11508) );
  AND U16141 ( .A(n16865), .B(n16382), .Z(n16863) );
  IV U16142 ( .A(n16866), .Z(n16382) );
  XOR U16143 ( .A(n10125), .B(n16867), .Z(n16858) );
  XOR U16144 ( .A(n16868), .B(n14705), .Z(n16867) );
  XNOR U16145 ( .A(n16869), .B(n16870), .Z(n14705) );
  AND U16146 ( .A(n16871), .B(n16386), .Z(n16869) );
  IV U16147 ( .A(n16872), .Z(n16386) );
  XOR U16148 ( .A(n16873), .B(n16874), .Z(n10125) );
  AND U16149 ( .A(n16875), .B(n16378), .Z(n16873) );
  IV U16150 ( .A(n16876), .Z(n16378) );
  XOR U16151 ( .A(n7992), .B(n5942), .Z(n2200) );
  XNOR U16152 ( .A(n16877), .B(n16878), .Z(n5942) );
  XNOR U16153 ( .A(n5251), .B(n3704), .Z(n16878) );
  XOR U16154 ( .A(n16879), .B(n8558), .Z(n3704) );
  IV U16155 ( .A(n10299), .Z(n8558) );
  XOR U16156 ( .A(n16880), .B(n10803), .Z(n10299) );
  XNOR U16157 ( .A(n11903), .B(n13554), .Z(n10803) );
  XNOR U16158 ( .A(n16881), .B(n16882), .Z(n13554) );
  XNOR U16159 ( .A(n14801), .B(n11548), .Z(n16882) );
  XOR U16160 ( .A(n16883), .B(n15730), .Z(n11548) );
  ANDN U16161 ( .B(n15731), .A(n12378), .Z(n16883) );
  XNOR U16162 ( .A(n16884), .B(n15735), .Z(n14801) );
  ANDN U16163 ( .B(n16885), .A(n16886), .Z(n16884) );
  XOR U16164 ( .A(n10218), .B(n16887), .Z(n16881) );
  XNOR U16165 ( .A(n12349), .B(n11391), .Z(n16887) );
  XNOR U16166 ( .A(n16888), .B(n15739), .Z(n11391) );
  NOR U16167 ( .A(n12300), .B(n15738), .Z(n16888) );
  XNOR U16168 ( .A(n16889), .B(n15742), .Z(n12349) );
  NOR U16169 ( .A(n15741), .B(n15229), .Z(n16889) );
  XNOR U16170 ( .A(n16890), .B(n15745), .Z(n10218) );
  AND U16171 ( .A(n12307), .B(n15746), .Z(n16890) );
  IV U16172 ( .A(n16891), .Z(n12307) );
  XOR U16173 ( .A(n16892), .B(n16893), .Z(n11903) );
  XOR U16174 ( .A(n12610), .B(n10595), .Z(n16893) );
  XOR U16175 ( .A(n16894), .B(n14270), .Z(n10595) );
  IV U16176 ( .A(n14812), .Z(n14270) );
  XNOR U16177 ( .A(n16895), .B(n16896), .Z(n14812) );
  NOR U16178 ( .A(n15621), .B(n14811), .Z(n16894) );
  XNOR U16179 ( .A(n16897), .B(n14264), .Z(n12610) );
  XOR U16180 ( .A(n16898), .B(n16899), .Z(n14264) );
  ANDN U16181 ( .B(n16900), .A(n15613), .Z(n16897) );
  XOR U16182 ( .A(n11556), .B(n16901), .Z(n16892) );
  XOR U16183 ( .A(n10232), .B(n9402), .Z(n16901) );
  XOR U16184 ( .A(n16902), .B(n15653), .Z(n9402) );
  IV U16185 ( .A(n14816), .Z(n15653) );
  XOR U16186 ( .A(n16903), .B(n16904), .Z(n14816) );
  NOR U16187 ( .A(n15617), .B(n14815), .Z(n16902) );
  XNOR U16188 ( .A(n16905), .B(n14274), .Z(n10232) );
  XNOR U16189 ( .A(n16906), .B(n16907), .Z(n14274) );
  ANDN U16190 ( .B(n15625), .A(n14806), .Z(n16905) );
  XNOR U16191 ( .A(n16908), .B(n14278), .Z(n11556) );
  XNOR U16192 ( .A(n16909), .B(n16910), .Z(n14278) );
  ANDN U16193 ( .B(n14819), .A(n15629), .Z(n16908) );
  AND U16194 ( .A(n7901), .B(n8559), .Z(n16879) );
  XOR U16195 ( .A(n15410), .B(n9582), .Z(n8559) );
  XNOR U16196 ( .A(n13322), .B(n15538), .Z(n9582) );
  XNOR U16197 ( .A(n16911), .B(n16912), .Z(n15538) );
  XOR U16198 ( .A(n11721), .B(n13860), .Z(n16912) );
  XOR U16199 ( .A(n16913), .B(n13952), .Z(n13860) );
  XOR U16200 ( .A(n16914), .B(n16779), .Z(n13952) );
  ANDN U16201 ( .B(n14200), .A(n15407), .Z(n16913) );
  XOR U16202 ( .A(n15974), .B(n16915), .Z(n14200) );
  XNOR U16203 ( .A(n16916), .B(n13960), .Z(n11721) );
  XNOR U16204 ( .A(n16917), .B(n15325), .Z(n13960) );
  AND U16205 ( .A(n15541), .B(n14207), .Z(n16916) );
  IV U16206 ( .A(n15540), .Z(n14207) );
  XOR U16207 ( .A(n16918), .B(n16919), .Z(n15540) );
  XOR U16208 ( .A(n14195), .B(n16920), .Z(n16911) );
  XOR U16209 ( .A(n12543), .B(n10228), .Z(n16920) );
  XOR U16210 ( .A(n16921), .B(n14202), .Z(n10228) );
  IV U16211 ( .A(n13947), .Z(n14202) );
  XOR U16212 ( .A(n16922), .B(n16469), .Z(n13947) );
  ANDN U16213 ( .B(n14203), .A(n15402), .Z(n16921) );
  XNOR U16214 ( .A(n16923), .B(n16924), .Z(n14203) );
  XNOR U16215 ( .A(n16925), .B(n13956), .Z(n12543) );
  XNOR U16216 ( .A(n16926), .B(n16552), .Z(n13956) );
  AND U16217 ( .A(n14210), .B(n15404), .Z(n16925) );
  XOR U16218 ( .A(n16927), .B(n16340), .Z(n14210) );
  XNOR U16219 ( .A(n16928), .B(n14213), .Z(n14195) );
  ANDN U16220 ( .B(n14214), .A(n15398), .Z(n16928) );
  XOR U16221 ( .A(n16049), .B(n16929), .Z(n14214) );
  XOR U16222 ( .A(n16930), .B(n16931), .Z(n13322) );
  XNOR U16223 ( .A(n9915), .B(n9533), .Z(n16931) );
  XOR U16224 ( .A(n16932), .B(n13679), .Z(n9533) );
  ANDN U16225 ( .B(n15413), .A(n13678), .Z(n16932) );
  XNOR U16226 ( .A(n16933), .B(n16934), .Z(n13678) );
  XOR U16227 ( .A(n16935), .B(n16053), .Z(n15413) );
  XOR U16228 ( .A(n16936), .B(n13940), .Z(n9915) );
  AND U16229 ( .A(n14459), .B(n13939), .Z(n16936) );
  XOR U16230 ( .A(n16937), .B(n16938), .Z(n13939) );
  XNOR U16231 ( .A(n16939), .B(n16940), .Z(n14459) );
  XOR U16232 ( .A(n11123), .B(n16941), .Z(n16930) );
  XOR U16233 ( .A(n11130), .B(n10271), .Z(n16941) );
  XNOR U16234 ( .A(n16942), .B(n13674), .Z(n10271) );
  AND U16235 ( .A(n13675), .B(n14453), .Z(n16942) );
  XNOR U16236 ( .A(n16943), .B(n16944), .Z(n14453) );
  XNOR U16237 ( .A(n16945), .B(n16919), .Z(n13675) );
  XOR U16238 ( .A(n16946), .B(n16947), .Z(n11130) );
  NOR U16239 ( .A(n13670), .B(n14449), .Z(n16946) );
  XOR U16240 ( .A(n16948), .B(n13666), .Z(n11123) );
  AND U16241 ( .A(n14456), .B(n15416), .Z(n16948) );
  XOR U16242 ( .A(n16949), .B(n16950), .Z(n15416) );
  XNOR U16243 ( .A(n16951), .B(n16952), .Z(n14456) );
  XNOR U16244 ( .A(n16953), .B(n13670), .Z(n15410) );
  XOR U16245 ( .A(n16954), .B(n16955), .Z(n13670) );
  ANDN U16246 ( .B(n14449), .A(n14450), .Z(n16953) );
  XNOR U16247 ( .A(n16956), .B(n16957), .Z(n14449) );
  XNOR U16248 ( .A(n16958), .B(n10916), .Z(n7901) );
  IV U16249 ( .A(n11373), .Z(n10916) );
  XNOR U16250 ( .A(n16959), .B(n14003), .Z(n11373) );
  XNOR U16251 ( .A(n16960), .B(n16961), .Z(n14003) );
  XOR U16252 ( .A(n11805), .B(n9916), .Z(n16961) );
  XOR U16253 ( .A(n16962), .B(n14559), .Z(n9916) );
  ANDN U16254 ( .B(n13714), .A(n16963), .Z(n16962) );
  XNOR U16255 ( .A(n16964), .B(n14554), .Z(n11805) );
  AND U16256 ( .A(n16965), .B(n13718), .Z(n16964) );
  XOR U16257 ( .A(n12888), .B(n16966), .Z(n16960) );
  XNOR U16258 ( .A(n16967), .B(n14010), .Z(n16966) );
  XNOR U16259 ( .A(n16968), .B(n14557), .Z(n14010) );
  ANDN U16260 ( .B(n13708), .A(n16969), .Z(n16968) );
  XNOR U16261 ( .A(n16970), .B(n14561), .Z(n12888) );
  AND U16262 ( .A(n16971), .B(n13704), .Z(n16970) );
  XNOR U16263 ( .A(n16972), .B(n8551), .Z(n5251) );
  XNOR U16264 ( .A(n16214), .B(n10019), .Z(n8551) );
  XNOR U16265 ( .A(n15787), .B(n16597), .Z(n10019) );
  XNOR U16266 ( .A(n16973), .B(n16974), .Z(n16597) );
  XOR U16267 ( .A(n12699), .B(n16167), .Z(n16974) );
  XOR U16268 ( .A(n16975), .B(n16182), .Z(n16167) );
  AND U16269 ( .A(n16183), .B(n16976), .Z(n16975) );
  XOR U16270 ( .A(n16416), .B(n16977), .Z(n16183) );
  XOR U16271 ( .A(n16978), .B(n16173), .Z(n12699) );
  AND U16272 ( .A(n16174), .B(n16979), .Z(n16978) );
  XNOR U16273 ( .A(n12258), .B(n16980), .Z(n16973) );
  XOR U16274 ( .A(n9575), .B(n10650), .Z(n16980) );
  XNOR U16275 ( .A(n16981), .B(n16178), .Z(n10650) );
  ANDN U16276 ( .B(n16177), .A(n16228), .Z(n16981) );
  IV U16277 ( .A(n16226), .Z(n16177) );
  XOR U16278 ( .A(n16982), .B(n16983), .Z(n16226) );
  XNOR U16279 ( .A(n16984), .B(n16187), .Z(n9575) );
  ANDN U16280 ( .B(n16186), .A(n16220), .Z(n16984) );
  XNOR U16281 ( .A(n16985), .B(n15516), .Z(n16186) );
  XNOR U16282 ( .A(n16986), .B(n16190), .Z(n12258) );
  ANDN U16283 ( .B(n16191), .A(n16216), .Z(n16986) );
  XNOR U16284 ( .A(n16987), .B(n16988), .Z(n16191) );
  XOR U16285 ( .A(n16989), .B(n16990), .Z(n15787) );
  XOR U16286 ( .A(n16991), .B(n10093), .Z(n16990) );
  XNOR U16287 ( .A(n16992), .B(n13215), .Z(n10093) );
  AND U16288 ( .A(n15047), .B(n16993), .Z(n16992) );
  XNOR U16289 ( .A(n16994), .B(n16995), .Z(n15047) );
  XNOR U16290 ( .A(n15339), .B(n16996), .Z(n16989) );
  XNOR U16291 ( .A(n9507), .B(n10308), .Z(n16996) );
  XNOR U16292 ( .A(n16997), .B(n15819), .Z(n10308) );
  ANDN U16293 ( .B(n15036), .A(n15034), .Z(n16997) );
  XNOR U16294 ( .A(n16998), .B(n16999), .Z(n15036) );
  XNOR U16295 ( .A(n17000), .B(n13209), .Z(n9507) );
  ANDN U16296 ( .B(n15038), .A(n15039), .Z(n17000) );
  XNOR U16297 ( .A(n17001), .B(n16348), .Z(n15039) );
  XOR U16298 ( .A(n17002), .B(n13205), .Z(n15339) );
  AND U16299 ( .A(n15803), .B(n15834), .Z(n17002) );
  IV U16300 ( .A(n15804), .Z(n15834) );
  XNOR U16301 ( .A(n17003), .B(n17004), .Z(n15804) );
  XNOR U16302 ( .A(n17005), .B(n16174), .Z(n16214) );
  XOR U16303 ( .A(n17006), .B(n17007), .Z(n16174) );
  AND U16304 ( .A(n8552), .B(n7893), .Z(n16972) );
  XOR U16305 ( .A(n11121), .B(n17009), .Z(n7893) );
  XNOR U16306 ( .A(n17010), .B(n13087), .Z(n11121) );
  XOR U16307 ( .A(n17011), .B(n17012), .Z(n13087) );
  XNOR U16308 ( .A(n15197), .B(n10538), .Z(n17012) );
  XOR U16309 ( .A(n17013), .B(n16722), .Z(n10538) );
  IV U16310 ( .A(n17014), .Z(n16722) );
  ANDN U16311 ( .B(n15930), .A(n15928), .Z(n17013) );
  XNOR U16312 ( .A(n17015), .B(n17016), .Z(n15928) );
  XNOR U16313 ( .A(n17017), .B(n17018), .Z(n15197) );
  ANDN U16314 ( .B(n15939), .A(n15937), .Z(n17017) );
  XNOR U16315 ( .A(n12826), .B(n17019), .Z(n17011) );
  XOR U16316 ( .A(n9273), .B(n9066), .Z(n17019) );
  XNOR U16317 ( .A(n17020), .B(n16715), .Z(n9066) );
  AND U16318 ( .A(n15934), .B(n15933), .Z(n17020) );
  IV U16319 ( .A(n16714), .Z(n15933) );
  XOR U16320 ( .A(n17021), .B(n16995), .Z(n16714) );
  XOR U16321 ( .A(n17022), .B(n16725), .Z(n9273) );
  XOR U16322 ( .A(n16691), .B(n17023), .Z(n15941) );
  XNOR U16323 ( .A(n17024), .B(n16719), .Z(n12826) );
  NOR U16324 ( .A(n15925), .B(n15924), .Z(n17024) );
  XOR U16325 ( .A(n15911), .B(n17025), .Z(n15924) );
  XNOR U16326 ( .A(n16442), .B(n17026), .Z(n8552) );
  XNOR U16327 ( .A(n17027), .B(n17028), .Z(n12805) );
  XOR U16328 ( .A(n10839), .B(n13918), .Z(n17028) );
  XOR U16329 ( .A(n17029), .B(n15939), .Z(n13918) );
  XNOR U16330 ( .A(n17030), .B(n17031), .Z(n15939) );
  NOR U16331 ( .A(n17032), .B(n15938), .Z(n17029) );
  XNOR U16332 ( .A(n17033), .B(n15930), .Z(n10839) );
  XNOR U16333 ( .A(n17034), .B(n17035), .Z(n15930) );
  NOR U16334 ( .A(n16721), .B(n15929), .Z(n17033) );
  XOR U16335 ( .A(n11453), .B(n17036), .Z(n17027) );
  XOR U16336 ( .A(n10901), .B(n12477), .Z(n17036) );
  XOR U16337 ( .A(n17037), .B(n15925), .Z(n12477) );
  XOR U16338 ( .A(n17038), .B(n17039), .Z(n15925) );
  XNOR U16339 ( .A(n17040), .B(n15934), .Z(n10901) );
  XOR U16340 ( .A(n17041), .B(n17042), .Z(n15934) );
  NOR U16341 ( .A(n15935), .B(n16713), .Z(n17040) );
  XNOR U16342 ( .A(n17043), .B(n15942), .Z(n11453) );
  XNOR U16343 ( .A(n17044), .B(n17045), .Z(n15942) );
  ANDN U16344 ( .B(n15943), .A(n16724), .Z(n17043) );
  XNOR U16345 ( .A(n6352), .B(n17047), .Z(n16877) );
  XOR U16346 ( .A(n2547), .B(n8539), .Z(n17047) );
  XOR U16347 ( .A(n17048), .B(n8544), .Z(n8539) );
  XOR U16348 ( .A(n17049), .B(n9216), .Z(n8544) );
  IV U16349 ( .A(n15224), .Z(n9216) );
  XOR U16350 ( .A(n14258), .B(n13189), .Z(n15224) );
  XNOR U16351 ( .A(n17050), .B(n17051), .Z(n13189) );
  XNOR U16352 ( .A(n12294), .B(n11181), .Z(n17051) );
  XOR U16353 ( .A(n17052), .B(n13056), .Z(n11181) );
  ANDN U16354 ( .B(n17053), .A(n15724), .Z(n17052) );
  XNOR U16355 ( .A(n17054), .B(n13061), .Z(n12294) );
  ANDN U16356 ( .B(n14332), .A(n13060), .Z(n17054) );
  XOR U16357 ( .A(n12284), .B(n17055), .Z(n17050) );
  XOR U16358 ( .A(n10702), .B(n10159), .Z(n17055) );
  XNOR U16359 ( .A(n17056), .B(n13064), .Z(n10159) );
  AND U16360 ( .A(n13065), .B(n14329), .Z(n17056) );
  XOR U16361 ( .A(n17057), .B(n17058), .Z(n10702) );
  NOR U16362 ( .A(n14337), .B(n13692), .Z(n17057) );
  XNOR U16363 ( .A(n17059), .B(n13068), .Z(n12284) );
  ANDN U16364 ( .B(n17060), .A(n14340), .Z(n17059) );
  XOR U16365 ( .A(n17061), .B(n17062), .Z(n14258) );
  XNOR U16366 ( .A(n11749), .B(n9563), .Z(n17062) );
  XNOR U16367 ( .A(n17063), .B(n12309), .Z(n9563) );
  ANDN U16368 ( .B(n15744), .A(n15745), .Z(n17063) );
  XNOR U16369 ( .A(n17064), .B(n17065), .Z(n15745) );
  XOR U16370 ( .A(n17066), .B(n16552), .Z(n15744) );
  XNOR U16371 ( .A(n17067), .B(n12302), .Z(n11749) );
  NOR U16372 ( .A(n12301), .B(n15739), .Z(n17067) );
  XNOR U16373 ( .A(n17068), .B(n17069), .Z(n15739) );
  XOR U16374 ( .A(n17070), .B(n16808), .Z(n12301) );
  XNOR U16375 ( .A(n11581), .B(n17071), .Z(n17061) );
  XOR U16376 ( .A(n9096), .B(n10640), .Z(n17071) );
  XOR U16377 ( .A(n17072), .B(n17073), .Z(n10640) );
  AND U16378 ( .A(n15733), .B(n15735), .Z(n17072) );
  XOR U16379 ( .A(n17074), .B(n17075), .Z(n15735) );
  XNOR U16380 ( .A(n17076), .B(n15231), .Z(n9096) );
  AND U16381 ( .A(n15230), .B(n15742), .Z(n17076) );
  XOR U16382 ( .A(n17077), .B(n17078), .Z(n15742) );
  XNOR U16383 ( .A(n16268), .B(n17079), .Z(n15230) );
  XNOR U16384 ( .A(n17080), .B(n12379), .Z(n11581) );
  ANDN U16385 ( .B(n12380), .A(n15730), .Z(n17080) );
  XNOR U16386 ( .A(n17081), .B(n17082), .Z(n15730) );
  XOR U16387 ( .A(n17083), .B(n17084), .Z(n12380) );
  ANDN U16388 ( .B(n8545), .A(n7897), .Z(n17048) );
  XNOR U16389 ( .A(n12429), .B(n11466), .Z(n7897) );
  IV U16390 ( .A(n11238), .Z(n11466) );
  XOR U16391 ( .A(n15659), .B(n17085), .Z(n11238) );
  XOR U16392 ( .A(n17086), .B(n17087), .Z(n15659) );
  XNOR U16393 ( .A(n11503), .B(n12373), .Z(n17087) );
  XNOR U16394 ( .A(n17088), .B(n17089), .Z(n12373) );
  XNOR U16395 ( .A(n17092), .B(n17093), .Z(n11503) );
  ANDN U16396 ( .B(n17094), .A(n17095), .Z(n17092) );
  XNOR U16397 ( .A(n12219), .B(n17096), .Z(n17086) );
  XOR U16398 ( .A(n11046), .B(n17097), .Z(n17096) );
  XOR U16399 ( .A(n17098), .B(n17099), .Z(n11046) );
  AND U16400 ( .A(n17100), .B(n17101), .Z(n17098) );
  XOR U16401 ( .A(n17102), .B(n17103), .Z(n12219) );
  ANDN U16402 ( .B(n17104), .A(n17105), .Z(n17102) );
  XNOR U16403 ( .A(n17106), .B(n14309), .Z(n12429) );
  ANDN U16404 ( .B(n17107), .A(n17108), .Z(n17106) );
  XNOR U16405 ( .A(n17109), .B(n12461), .Z(n8545) );
  IV U16406 ( .A(n9946), .Z(n12461) );
  XNOR U16407 ( .A(n12577), .B(n14132), .Z(n9946) );
  XNOR U16408 ( .A(n17110), .B(n17111), .Z(n14132) );
  XNOR U16409 ( .A(n10882), .B(n12313), .Z(n17111) );
  XOR U16410 ( .A(n17112), .B(n14347), .Z(n12313) );
  AND U16411 ( .A(n14134), .B(n13502), .Z(n17112) );
  XNOR U16412 ( .A(n17113), .B(n16003), .Z(n13502) );
  XNOR U16413 ( .A(n17114), .B(n16009), .Z(n14134) );
  XNOR U16414 ( .A(n17115), .B(n13016), .Z(n10882) );
  ANDN U16415 ( .B(n13029), .A(n13015), .Z(n17115) );
  XNOR U16416 ( .A(n17116), .B(n16818), .Z(n13015) );
  XOR U16417 ( .A(n14914), .B(n17117), .Z(n13029) );
  XOR U16418 ( .A(n12465), .B(n17118), .Z(n17110) );
  XNOR U16419 ( .A(n9553), .B(n9666), .Z(n17118) );
  XNOR U16420 ( .A(n17119), .B(n13004), .Z(n9666) );
  AND U16421 ( .A(n13005), .B(n13038), .Z(n17119) );
  XOR U16422 ( .A(n17120), .B(n17121), .Z(n13038) );
  XNOR U16423 ( .A(n17122), .B(n17123), .Z(n13005) );
  XOR U16424 ( .A(n17124), .B(n17125), .Z(n9553) );
  AND U16425 ( .A(n13033), .B(n13035), .Z(n17124) );
  XOR U16426 ( .A(n17126), .B(n17127), .Z(n13035) );
  XOR U16427 ( .A(n17128), .B(n17129), .Z(n12465) );
  ANDN U16428 ( .B(n13009), .A(n13388), .Z(n17128) );
  XNOR U16429 ( .A(n17130), .B(n17131), .Z(n13388) );
  XNOR U16430 ( .A(n17003), .B(n17132), .Z(n13009) );
  XOR U16431 ( .A(n17133), .B(n17134), .Z(n12577) );
  XNOR U16432 ( .A(n10361), .B(n11432), .Z(n17134) );
  XOR U16433 ( .A(n17135), .B(n12972), .Z(n11432) );
  XOR U16434 ( .A(n17136), .B(n17137), .Z(n12972) );
  ANDN U16435 ( .B(n13457), .A(n15250), .Z(n17135) );
  XNOR U16436 ( .A(n17138), .B(n13465), .Z(n10361) );
  XOR U16437 ( .A(n17139), .B(n17140), .Z(n13465) );
  XOR U16438 ( .A(n12998), .B(n17141), .Z(n17133) );
  XOR U16439 ( .A(n11118), .B(n10064), .Z(n17141) );
  XNOR U16440 ( .A(n17142), .B(n12748), .Z(n10064) );
  XOR U16441 ( .A(n17143), .B(n17144), .Z(n12748) );
  ANDN U16442 ( .B(n15254), .A(n13454), .Z(n17142) );
  XNOR U16443 ( .A(n17145), .B(n12754), .Z(n11118) );
  XNOR U16444 ( .A(n17146), .B(n16988), .Z(n12754) );
  AND U16445 ( .A(n13459), .B(n15241), .Z(n17145) );
  XNOR U16446 ( .A(n17147), .B(n12759), .Z(n12998) );
  XNOR U16447 ( .A(n17148), .B(n17149), .Z(n12759) );
  NOR U16448 ( .A(n13462), .B(n15258), .Z(n17147) );
  XOR U16449 ( .A(n17150), .B(n8555), .Z(n2547) );
  XOR U16450 ( .A(n14631), .B(n9573), .Z(n8555) );
  XOR U16451 ( .A(n17151), .B(n17152), .Z(n14631) );
  AND U16452 ( .A(n16835), .B(n14066), .Z(n17151) );
  XOR U16453 ( .A(n17153), .B(n16009), .Z(n14066) );
  IV U16454 ( .A(n17154), .Z(n16009) );
  ANDN U16455 ( .B(n10486), .A(n8556), .Z(n17150) );
  XOR U16456 ( .A(n10154), .B(n14653), .Z(n8556) );
  XNOR U16457 ( .A(n17155), .B(n17156), .Z(n14653) );
  ANDN U16458 ( .B(n15085), .A(n15086), .Z(n17155) );
  XNOR U16459 ( .A(n12558), .B(n17157), .Z(n10154) );
  XOR U16460 ( .A(n17158), .B(n17159), .Z(n12558) );
  XNOR U16461 ( .A(n12181), .B(n9594), .Z(n17159) );
  XOR U16462 ( .A(n17160), .B(n17161), .Z(n9594) );
  AND U16463 ( .A(n14658), .B(n14656), .Z(n17160) );
  XOR U16464 ( .A(n17162), .B(n17163), .Z(n14658) );
  XNOR U16465 ( .A(n17164), .B(n17165), .Z(n12181) );
  AND U16466 ( .A(n14660), .B(n15082), .Z(n17164) );
  IV U16467 ( .A(n14661), .Z(n15082) );
  XNOR U16468 ( .A(n17166), .B(n17167), .Z(n14661) );
  XNOR U16469 ( .A(n13902), .B(n17168), .Z(n17158) );
  XNOR U16470 ( .A(n14007), .B(n9712), .Z(n17168) );
  XNOR U16471 ( .A(n17169), .B(n17170), .Z(n9712) );
  AND U16472 ( .A(n14650), .B(n15092), .Z(n17169) );
  IV U16473 ( .A(n14652), .Z(n15092) );
  XNOR U16474 ( .A(n17171), .B(n15329), .Z(n14652) );
  XOR U16475 ( .A(n17172), .B(n17173), .Z(n14007) );
  ANDN U16476 ( .B(n14646), .A(n14648), .Z(n17172) );
  XNOR U16477 ( .A(n17174), .B(n17175), .Z(n14648) );
  XNOR U16478 ( .A(n17176), .B(n17177), .Z(n13902) );
  NOR U16479 ( .A(n17156), .B(n15085), .Z(n17176) );
  XNOR U16480 ( .A(n17126), .B(n17178), .Z(n15085) );
  XOR U16481 ( .A(n11538), .B(n13525), .Z(n10486) );
  XOR U16482 ( .A(n17179), .B(n17180), .Z(n13525) );
  AND U16483 ( .A(n14188), .B(n14190), .Z(n17179) );
  XOR U16484 ( .A(n17181), .B(n14709), .Z(n11538) );
  XOR U16485 ( .A(n17182), .B(n17183), .Z(n14709) );
  XOR U16486 ( .A(n13268), .B(n14217), .Z(n17183) );
  XOR U16487 ( .A(n17184), .B(n14228), .Z(n14217) );
  NOR U16488 ( .A(n13522), .B(n13523), .Z(n17184) );
  XNOR U16489 ( .A(n17185), .B(n17186), .Z(n13523) );
  XNOR U16490 ( .A(n17187), .B(n17188), .Z(n13522) );
  XNOR U16491 ( .A(n17189), .B(n16800), .Z(n13268) );
  ANDN U16492 ( .B(n13529), .A(n13530), .Z(n17189) );
  XNOR U16493 ( .A(n17190), .B(n17191), .Z(n13530) );
  IV U16494 ( .A(n16801), .Z(n13529) );
  XOR U16495 ( .A(n17192), .B(n17193), .Z(n16801) );
  XOR U16496 ( .A(n13276), .B(n17194), .Z(n17182) );
  XOR U16497 ( .A(n12590), .B(n11915), .Z(n17194) );
  XOR U16498 ( .A(n17195), .B(n14622), .Z(n11915) );
  ANDN U16499 ( .B(n13518), .A(n13519), .Z(n17195) );
  XNOR U16500 ( .A(n17196), .B(n17197), .Z(n13519) );
  XNOR U16501 ( .A(n17198), .B(n17199), .Z(n13518) );
  XNOR U16502 ( .A(n17200), .B(n17201), .Z(n12590) );
  ANDN U16503 ( .B(n17180), .A(n14188), .Z(n17200) );
  XOR U16504 ( .A(n17202), .B(n17203), .Z(n14188) );
  XOR U16505 ( .A(n17204), .B(n14226), .Z(n13276) );
  ANDN U16506 ( .B(n14176), .A(n14225), .Z(n17204) );
  XNOR U16507 ( .A(n17205), .B(n17206), .Z(n14225) );
  XNOR U16508 ( .A(n17207), .B(n17208), .Z(n14176) );
  XOR U16509 ( .A(n17209), .B(n8547), .Z(n6352) );
  XOR U16510 ( .A(n10094), .B(n16991), .Z(n8547) );
  XOR U16511 ( .A(n17210), .B(n17211), .Z(n16991) );
  AND U16512 ( .A(n15044), .B(n17212), .Z(n17210) );
  XOR U16513 ( .A(n16751), .B(n17213), .Z(n15044) );
  XOR U16514 ( .A(n14002), .B(n16168), .Z(n10094) );
  XOR U16515 ( .A(n17214), .B(n17215), .Z(n16168) );
  XOR U16516 ( .A(n10481), .B(n11139), .Z(n17215) );
  XOR U16517 ( .A(n17216), .B(n13214), .Z(n11139) );
  XNOR U16518 ( .A(n17217), .B(n17218), .Z(n13214) );
  AND U16519 ( .A(n13215), .B(n15046), .Z(n17216) );
  IV U16520 ( .A(n16993), .Z(n15046) );
  XNOR U16521 ( .A(n17219), .B(n16672), .Z(n16993) );
  XNOR U16522 ( .A(n17220), .B(n17221), .Z(n13215) );
  XNOR U16523 ( .A(n17222), .B(n13218), .Z(n10481) );
  XNOR U16524 ( .A(n17223), .B(n17224), .Z(n13218) );
  AND U16525 ( .A(n15043), .B(n17211), .Z(n17222) );
  IV U16526 ( .A(n13219), .Z(n17211) );
  XNOR U16527 ( .A(n17225), .B(n17031), .Z(n13219) );
  IV U16528 ( .A(n17212), .Z(n15043) );
  XOR U16529 ( .A(n17226), .B(n17227), .Z(n17212) );
  XOR U16530 ( .A(n10120), .B(n17228), .Z(n17214) );
  XNOR U16531 ( .A(n13198), .B(n11838), .Z(n17228) );
  XNOR U16532 ( .A(n17229), .B(n13204), .Z(n11838) );
  XNOR U16533 ( .A(n17230), .B(n17231), .Z(n13204) );
  ANDN U16534 ( .B(n13205), .A(n15803), .Z(n17229) );
  XNOR U16535 ( .A(n15650), .B(n17232), .Z(n15803) );
  XOR U16536 ( .A(n17233), .B(n17234), .Z(n13205) );
  XNOR U16537 ( .A(n17235), .B(n15820), .Z(n13198) );
  XOR U16538 ( .A(n17236), .B(n16055), .Z(n15820) );
  AND U16539 ( .A(n15034), .B(n15819), .Z(n17235) );
  XNOR U16540 ( .A(n17237), .B(n17238), .Z(n15819) );
  XOR U16541 ( .A(n17239), .B(n17240), .Z(n15034) );
  XNOR U16542 ( .A(n17241), .B(n13208), .Z(n10120) );
  XNOR U16543 ( .A(n17242), .B(n17243), .Z(n13208) );
  NOR U16544 ( .A(n15038), .B(n13209), .Z(n17241) );
  XNOR U16545 ( .A(n17245), .B(n16539), .Z(n15038) );
  XOR U16546 ( .A(n17246), .B(n17247), .Z(n14002) );
  XOR U16547 ( .A(n10438), .B(n10941), .Z(n17247) );
  XOR U16548 ( .A(n17248), .B(n15857), .Z(n10941) );
  AND U16549 ( .A(n15796), .B(n13733), .Z(n17248) );
  XNOR U16550 ( .A(n17249), .B(n16261), .Z(n13733) );
  XNOR U16551 ( .A(n17250), .B(n15861), .Z(n10438) );
  ANDN U16552 ( .B(n13728), .A(n15793), .Z(n17250) );
  XOR U16553 ( .A(n10835), .B(n17252), .Z(n17246) );
  XNOR U16554 ( .A(n9111), .B(n17253), .Z(n17252) );
  XNOR U16555 ( .A(n17254), .B(n15852), .Z(n9111) );
  IV U16556 ( .A(n17255), .Z(n15852) );
  NOR U16557 ( .A(n15798), .B(n13724), .Z(n17254) );
  XNOR U16558 ( .A(n17256), .B(n17131), .Z(n13724) );
  XNOR U16559 ( .A(n17257), .B(n15847), .Z(n10835) );
  AND U16560 ( .A(n15791), .B(n13741), .Z(n17257) );
  XOR U16561 ( .A(n17258), .B(n17259), .Z(n13741) );
  ANDN U16562 ( .B(n8548), .A(n7888), .Z(n17209) );
  XNOR U16563 ( .A(n15707), .B(n11971), .Z(n7888) );
  XNOR U16564 ( .A(n17260), .B(n15170), .Z(n15707) );
  ANDN U16565 ( .B(n15703), .A(n15704), .Z(n17260) );
  XOR U16566 ( .A(n16110), .B(n16127), .Z(n9505) );
  XNOR U16567 ( .A(n17261), .B(n17262), .Z(n16127) );
  XNOR U16568 ( .A(n10773), .B(n17263), .Z(n17262) );
  XNOR U16569 ( .A(n17264), .B(n14957), .Z(n10773) );
  AND U16570 ( .A(n17265), .B(n16306), .Z(n17264) );
  IV U16571 ( .A(n17266), .Z(n16306) );
  XNOR U16572 ( .A(n10933), .B(n17267), .Z(n17261) );
  XOR U16573 ( .A(n10952), .B(n11820), .Z(n17267) );
  XOR U16574 ( .A(n17268), .B(n14743), .Z(n11820) );
  ANDN U16575 ( .B(n16313), .A(n16816), .Z(n17268) );
  XNOR U16576 ( .A(n17269), .B(n17270), .Z(n16313) );
  XOR U16577 ( .A(n17271), .B(n14754), .Z(n10952) );
  AND U16578 ( .A(n16806), .B(n16308), .Z(n17271) );
  XOR U16579 ( .A(n17272), .B(n17273), .Z(n16308) );
  XOR U16580 ( .A(n17274), .B(n16290), .Z(n10933) );
  AND U16581 ( .A(n16820), .B(n16823), .Z(n17274) );
  IV U16582 ( .A(n16821), .Z(n16823) );
  XOR U16583 ( .A(n17275), .B(n17276), .Z(n16821) );
  XOR U16584 ( .A(n17277), .B(n17278), .Z(n16110) );
  XNOR U16585 ( .A(n12603), .B(n13071), .Z(n17278) );
  NOR U16586 ( .A(n16294), .B(n17280), .Z(n17279) );
  XNOR U16587 ( .A(n17281), .B(n11949), .Z(n12603) );
  ANDN U16588 ( .B(n17282), .A(n17283), .Z(n17281) );
  XOR U16589 ( .A(n12856), .B(n17284), .Z(n17277) );
  XOR U16590 ( .A(n16195), .B(n16151), .Z(n17284) );
  XOR U16591 ( .A(n17285), .B(n11962), .Z(n16151) );
  XNOR U16592 ( .A(n17287), .B(n11958), .Z(n16195) );
  ANDN U16593 ( .B(n17288), .A(n16296), .Z(n17287) );
  XNOR U16594 ( .A(n17289), .B(n11953), .Z(n12856) );
  ANDN U16595 ( .B(n17290), .A(n16302), .Z(n17289) );
  XNOR U16596 ( .A(n17291), .B(n17265), .Z(n16814) );
  AND U16597 ( .A(n14955), .B(n17266), .Z(n17291) );
  XOR U16598 ( .A(n17292), .B(n16016), .Z(n17266) );
  XOR U16599 ( .A(n17293), .B(n16788), .Z(n14955) );
  XOR U16600 ( .A(n17294), .B(n17295), .Z(n7992) );
  XNOR U16601 ( .A(n4912), .B(n10568), .Z(n17295) );
  XOR U16602 ( .A(n17296), .B(n6928), .Z(n10568) );
  XNOR U16603 ( .A(n14240), .B(n10896), .Z(n6928) );
  IV U16604 ( .A(n10113), .Z(n10896) );
  XNOR U16605 ( .A(n17299), .B(n15063), .Z(n14240) );
  AND U16606 ( .A(n17300), .B(n16590), .Z(n17299) );
  ANDN U16607 ( .B(n10483), .A(n9305), .Z(n17296) );
  XNOR U16608 ( .A(n13712), .B(n10436), .Z(n9305) );
  XNOR U16609 ( .A(n13381), .B(n16480), .Z(n10436) );
  XNOR U16610 ( .A(n17301), .B(n17302), .Z(n16480) );
  XOR U16611 ( .A(n17303), .B(n11150), .Z(n17302) );
  XNOR U16612 ( .A(n17304), .B(n17305), .Z(n11150) );
  AND U16613 ( .A(n17306), .B(n17307), .Z(n17304) );
  XOR U16614 ( .A(n11025), .B(n17308), .Z(n17301) );
  XOR U16615 ( .A(n10642), .B(n10143), .Z(n17308) );
  XOR U16616 ( .A(n17309), .B(n17310), .Z(n10143) );
  ANDN U16617 ( .B(n17311), .A(n17312), .Z(n17309) );
  XOR U16618 ( .A(n17313), .B(n17314), .Z(n10642) );
  ANDN U16619 ( .B(n17315), .A(n17316), .Z(n17313) );
  XNOR U16620 ( .A(n17317), .B(n17318), .Z(n11025) );
  AND U16621 ( .A(n17319), .B(n17320), .Z(n17317) );
  XOR U16622 ( .A(n17321), .B(n17322), .Z(n13381) );
  XNOR U16623 ( .A(n11728), .B(n11372), .Z(n17322) );
  XNOR U16624 ( .A(n17323), .B(n16971), .Z(n11372) );
  NOR U16625 ( .A(n13704), .B(n13705), .Z(n17323) );
  XNOR U16626 ( .A(n17324), .B(n15615), .Z(n13705) );
  XNOR U16627 ( .A(n17325), .B(n16067), .Z(n13704) );
  XOR U16628 ( .A(n17326), .B(n16969), .Z(n11728) );
  NOR U16629 ( .A(n13708), .B(n13709), .Z(n17326) );
  XNOR U16630 ( .A(n17327), .B(n15603), .Z(n13709) );
  XNOR U16631 ( .A(n17328), .B(n17329), .Z(n13708) );
  XOR U16632 ( .A(n16958), .B(n17330), .Z(n17321) );
  XNOR U16633 ( .A(n14824), .B(n10915), .Z(n17330) );
  XOR U16634 ( .A(n17331), .B(n16963), .Z(n10915) );
  NOR U16635 ( .A(n13714), .B(n13715), .Z(n17331) );
  XOR U16636 ( .A(n17332), .B(n17333), .Z(n13715) );
  XNOR U16637 ( .A(n17334), .B(n17197), .Z(n13714) );
  XNOR U16638 ( .A(n17335), .B(n17336), .Z(n14824) );
  NOR U16639 ( .A(n17337), .B(n14550), .Z(n17335) );
  XNOR U16640 ( .A(n17338), .B(n16965), .Z(n16958) );
  NOR U16641 ( .A(n13718), .B(n13719), .Z(n17338) );
  XOR U16642 ( .A(n17339), .B(n16988), .Z(n13719) );
  XOR U16643 ( .A(n17340), .B(n17341), .Z(n13718) );
  XNOR U16644 ( .A(n17342), .B(n17337), .Z(n13712) );
  ANDN U16645 ( .B(n14550), .A(n14551), .Z(n17342) );
  XOR U16646 ( .A(n16547), .B(n17343), .Z(n14550) );
  XNOR U16647 ( .A(n17344), .B(n10665), .Z(n10483) );
  IV U16648 ( .A(n16640), .Z(n10665) );
  XOR U16649 ( .A(n17010), .B(n15393), .Z(n16640) );
  XNOR U16650 ( .A(n17345), .B(n17346), .Z(n15393) );
  XOR U16651 ( .A(n11115), .B(n12600), .Z(n17346) );
  XOR U16652 ( .A(n17347), .B(n16387), .Z(n12600) );
  XNOR U16653 ( .A(n17348), .B(n16374), .Z(n11115) );
  ANDN U16654 ( .B(n16375), .A(n16861), .Z(n17348) );
  XOR U16655 ( .A(n10385), .B(n17349), .Z(n17345) );
  XOR U16656 ( .A(n12158), .B(n10837), .Z(n17349) );
  XOR U16657 ( .A(n17350), .B(n16384), .Z(n10837) );
  ANDN U16658 ( .B(n16383), .A(n16864), .Z(n17350) );
  IV U16659 ( .A(n17351), .Z(n16383) );
  XNOR U16660 ( .A(n17352), .B(n16370), .Z(n12158) );
  ANDN U16661 ( .B(n16371), .A(n17353), .Z(n17352) );
  XNOR U16662 ( .A(n17354), .B(n16379), .Z(n10385) );
  ANDN U16663 ( .B(n17355), .A(n16874), .Z(n17354) );
  XOR U16664 ( .A(n17356), .B(n17357), .Z(n17010) );
  XNOR U16665 ( .A(n11643), .B(n14623), .Z(n17357) );
  XOR U16666 ( .A(n17358), .B(n16237), .Z(n14623) );
  IV U16667 ( .A(n16694), .Z(n16237) );
  XNOR U16668 ( .A(n17359), .B(n17360), .Z(n16694) );
  ANDN U16669 ( .B(n15945), .A(n16693), .Z(n17358) );
  XNOR U16670 ( .A(n17361), .B(n16240), .Z(n11643) );
  XNOR U16671 ( .A(n17362), .B(n17363), .Z(n16240) );
  NOR U16672 ( .A(n16699), .B(n14321), .Z(n17361) );
  XOR U16673 ( .A(n10269), .B(n17364), .Z(n17356) );
  XOR U16674 ( .A(n10122), .B(n16683), .Z(n17364) );
  XOR U16675 ( .A(n17365), .B(n16235), .Z(n16683) );
  IV U16676 ( .A(n16704), .Z(n16235) );
  XNOR U16677 ( .A(n17366), .B(n13896), .Z(n16704) );
  ANDN U16678 ( .B(n12816), .A(n16703), .Z(n17365) );
  XNOR U16679 ( .A(n17367), .B(n16242), .Z(n10122) );
  XNOR U16680 ( .A(n17368), .B(n17369), .Z(n16242) );
  NOR U16681 ( .A(n12810), .B(n16708), .Z(n17367) );
  XNOR U16682 ( .A(n17370), .B(n16244), .Z(n10269) );
  XNOR U16683 ( .A(n17371), .B(n16021), .Z(n16244) );
  NOR U16684 ( .A(n12820), .B(n16689), .Z(n17370) );
  XOR U16685 ( .A(n17372), .B(n6933), .Z(n4912) );
  IV U16686 ( .A(n10579), .Z(n6933) );
  XOR U16687 ( .A(n15183), .B(n10061), .Z(n10579) );
  IV U16688 ( .A(n12135), .Z(n10061) );
  XOR U16689 ( .A(n15726), .B(n12765), .Z(n12135) );
  XNOR U16690 ( .A(n17373), .B(n17374), .Z(n12765) );
  XNOR U16691 ( .A(n13187), .B(n11798), .Z(n17374) );
  XOR U16692 ( .A(n17375), .B(n13792), .Z(n11798) );
  XNOR U16693 ( .A(n17376), .B(n15208), .Z(n13792) );
  XOR U16694 ( .A(n16024), .B(n17377), .Z(n13791) );
  XNOR U16695 ( .A(n17378), .B(n13795), .Z(n13187) );
  XNOR U16696 ( .A(n17379), .B(n17380), .Z(n13795) );
  ANDN U16697 ( .B(n13796), .A(n17381), .Z(n17378) );
  XOR U16698 ( .A(n10009), .B(n17382), .Z(n17373) );
  XOR U16699 ( .A(n12051), .B(n11765), .Z(n17382) );
  XOR U16700 ( .A(n17383), .B(n13801), .Z(n11765) );
  XNOR U16701 ( .A(n17384), .B(n16337), .Z(n13801) );
  NOR U16702 ( .A(n15185), .B(n13800), .Z(n17383) );
  XOR U16703 ( .A(n17174), .B(n17385), .Z(n13800) );
  XNOR U16704 ( .A(n17386), .B(n13804), .Z(n12051) );
  XNOR U16705 ( .A(n17387), .B(n17388), .Z(n13804) );
  ANDN U16706 ( .B(n15193), .A(n13805), .Z(n17386) );
  XNOR U16707 ( .A(n17389), .B(n17390), .Z(n13805) );
  XOR U16708 ( .A(n17391), .B(n17392), .Z(n10009) );
  NOR U16709 ( .A(n15189), .B(n13808), .Z(n17391) );
  XOR U16710 ( .A(n17393), .B(n16746), .Z(n13808) );
  XOR U16711 ( .A(n17394), .B(n17395), .Z(n15726) );
  XOR U16712 ( .A(n15223), .B(n17049), .Z(n17395) );
  XOR U16713 ( .A(n17396), .B(n13065), .Z(n17049) );
  XNOR U16714 ( .A(n17397), .B(n17398), .Z(n13065) );
  XOR U16715 ( .A(n17399), .B(n16792), .Z(n14329) );
  XOR U16716 ( .A(n17400), .B(n13055), .Z(n15223) );
  IV U16717 ( .A(n17053), .Z(n13055) );
  XOR U16718 ( .A(n17083), .B(n17401), .Z(n17053) );
  ANDN U16719 ( .B(n15724), .A(n15725), .Z(n17400) );
  XNOR U16720 ( .A(n17402), .B(n17403), .Z(n15724) );
  XNOR U16721 ( .A(n11317), .B(n17404), .Z(n17394) );
  XNOR U16722 ( .A(n12216), .B(n9215), .Z(n17404) );
  XNOR U16723 ( .A(n17405), .B(n13692), .Z(n9215) );
  XOR U16724 ( .A(n17406), .B(n17407), .Z(n13692) );
  AND U16725 ( .A(n14337), .B(n14338), .Z(n17405) );
  XNOR U16726 ( .A(n17408), .B(n16047), .Z(n14337) );
  XOR U16727 ( .A(n17409), .B(n13060), .Z(n12216) );
  XOR U16728 ( .A(n17410), .B(n16062), .Z(n13060) );
  XNOR U16729 ( .A(n17411), .B(n17412), .Z(n14332) );
  XNOR U16730 ( .A(n17413), .B(n13069), .Z(n11317) );
  IV U16731 ( .A(n17060), .Z(n13069) );
  XOR U16732 ( .A(n17414), .B(n17415), .Z(n17060) );
  AND U16733 ( .A(n14341), .B(n14340), .Z(n17413) );
  XOR U16734 ( .A(n17417), .B(n13796), .Z(n15183) );
  XNOR U16735 ( .A(n17418), .B(n14941), .Z(n13796) );
  ANDN U16736 ( .B(n17381), .A(n15722), .Z(n17417) );
  NOR U16737 ( .A(n9300), .B(n10468), .Z(n17372) );
  XNOR U16738 ( .A(n13558), .B(n9261), .Z(n10468) );
  XNOR U16739 ( .A(n11913), .B(n17085), .Z(n9261) );
  XNOR U16740 ( .A(n17419), .B(n17420), .Z(n17085) );
  XNOR U16741 ( .A(n11595), .B(n12685), .Z(n17420) );
  XNOR U16742 ( .A(n17421), .B(n17422), .Z(n12685) );
  ANDN U16743 ( .B(n12424), .A(n12422), .Z(n17421) );
  XNOR U16744 ( .A(n17423), .B(n14315), .Z(n11595) );
  AND U16745 ( .A(n12426), .B(n17424), .Z(n17423) );
  XOR U16746 ( .A(n17425), .B(n17426), .Z(n12426) );
  XNOR U16747 ( .A(n11983), .B(n17427), .Z(n17419) );
  XOR U16748 ( .A(n9517), .B(n11318), .Z(n17427) );
  XOR U16749 ( .A(n17428), .B(n14308), .Z(n11318) );
  AND U16750 ( .A(n17108), .B(n14309), .Z(n17428) );
  XNOR U16751 ( .A(n17003), .B(n17429), .Z(n14309) );
  XOR U16752 ( .A(n17430), .B(n17431), .Z(n9517) );
  AND U16753 ( .A(n12438), .B(n12436), .Z(n17430) );
  XNOR U16754 ( .A(n17432), .B(n14305), .Z(n11983) );
  AND U16755 ( .A(n12434), .B(n14304), .Z(n17432) );
  IV U16756 ( .A(n12432), .Z(n14304) );
  XOR U16757 ( .A(n17433), .B(n17434), .Z(n12432) );
  XOR U16758 ( .A(n17435), .B(n17436), .Z(n11913) );
  XOR U16759 ( .A(n13085), .B(n14283), .Z(n17436) );
  XNOR U16760 ( .A(n17437), .B(n14299), .Z(n14283) );
  AND U16761 ( .A(n13568), .B(n12490), .Z(n17437) );
  XOR U16762 ( .A(n17438), .B(n17439), .Z(n12490) );
  XNOR U16763 ( .A(n17440), .B(n17441), .Z(n13568) );
  XNOR U16764 ( .A(n17442), .B(n14288), .Z(n13085) );
  AND U16765 ( .A(n13566), .B(n12499), .Z(n17442) );
  XOR U16766 ( .A(n17443), .B(n17069), .Z(n12499) );
  XNOR U16767 ( .A(n15650), .B(n17444), .Z(n13566) );
  IV U16768 ( .A(n17445), .Z(n15650) );
  XNOR U16769 ( .A(n13698), .B(n17446), .Z(n17435) );
  XOR U16770 ( .A(n12523), .B(n9178), .Z(n17446) );
  XNOR U16771 ( .A(n17447), .B(n14295), .Z(n9178) );
  ANDN U16772 ( .B(n14296), .A(n12495), .Z(n17447) );
  XOR U16773 ( .A(n17448), .B(n14293), .Z(n12523) );
  XNOR U16774 ( .A(n17449), .B(n17167), .Z(n12486) );
  XOR U16775 ( .A(n17450), .B(n17451), .Z(n13564) );
  XNOR U16776 ( .A(n17452), .B(n14290), .Z(n13698) );
  ANDN U16777 ( .B(n12503), .A(n13560), .Z(n17452) );
  XOR U16778 ( .A(n17453), .B(n16792), .Z(n13560) );
  IV U16779 ( .A(n13561), .Z(n12503) );
  XOR U16780 ( .A(n17454), .B(n17455), .Z(n13561) );
  XOR U16781 ( .A(n17456), .B(n14296), .Z(n13558) );
  XOR U16782 ( .A(n17457), .B(n17458), .Z(n14296) );
  AND U16783 ( .A(n12497), .B(n12495), .Z(n17456) );
  XOR U16784 ( .A(n17459), .B(n16749), .Z(n12495) );
  XNOR U16785 ( .A(n16419), .B(n12884), .Z(n9300) );
  IV U16786 ( .A(n13018), .Z(n12884) );
  XOR U16787 ( .A(n13941), .B(n17460), .Z(n13018) );
  XOR U16788 ( .A(n17461), .B(n17462), .Z(n13941) );
  XNOR U16789 ( .A(n11887), .B(n14443), .Z(n17462) );
  XOR U16790 ( .A(n17463), .B(n14457), .Z(n14443) );
  XNOR U16791 ( .A(n17464), .B(n17465), .Z(n14457) );
  ANDN U16792 ( .B(n13666), .A(n13664), .Z(n17463) );
  XOR U16793 ( .A(n17468), .B(n17469), .Z(n13666) );
  XNOR U16794 ( .A(n17470), .B(n14460), .Z(n11887) );
  XNOR U16795 ( .A(n17471), .B(n16910), .Z(n14460) );
  IV U16796 ( .A(n17472), .Z(n16910) );
  ANDN U16797 ( .B(n13940), .A(n13938), .Z(n17470) );
  XOR U16798 ( .A(n17473), .B(n17474), .Z(n13938) );
  XNOR U16799 ( .A(n17475), .B(n17231), .Z(n13940) );
  XOR U16800 ( .A(n13328), .B(n17476), .Z(n17461) );
  XNOR U16801 ( .A(n13443), .B(n14345), .Z(n17476) );
  XNOR U16802 ( .A(n17477), .B(n15412), .Z(n14345) );
  XOR U16803 ( .A(n17478), .B(n15525), .Z(n15412) );
  AND U16804 ( .A(n13677), .B(n13679), .Z(n17477) );
  XOR U16805 ( .A(n17479), .B(n16011), .Z(n13679) );
  XNOR U16806 ( .A(n17480), .B(n16055), .Z(n13677) );
  XNOR U16807 ( .A(n17481), .B(n14454), .Z(n13443) );
  XOR U16808 ( .A(n17482), .B(n17483), .Z(n14454) );
  ANDN U16809 ( .B(n13673), .A(n13674), .Z(n17481) );
  XNOR U16810 ( .A(n17484), .B(n17485), .Z(n13674) );
  XNOR U16811 ( .A(n17486), .B(n16476), .Z(n13673) );
  XNOR U16812 ( .A(n17487), .B(n14450), .Z(n13328) );
  XOR U16813 ( .A(n17488), .B(n17489), .Z(n14450) );
  AND U16814 ( .A(n13669), .B(n16947), .Z(n17487) );
  IV U16815 ( .A(n13671), .Z(n16947) );
  XOR U16816 ( .A(n17490), .B(n16924), .Z(n13671) );
  XNOR U16817 ( .A(n17491), .B(n17492), .Z(n13669) );
  XNOR U16818 ( .A(n17493), .B(n15534), .Z(n16419) );
  XOR U16819 ( .A(n17494), .B(n17495), .Z(n13163) );
  XOR U16820 ( .A(n2644), .B(n17496), .Z(n17294) );
  XOR U16821 ( .A(n3522), .B(n5703), .Z(n17496) );
  XOR U16822 ( .A(n17497), .B(n6922), .Z(n5703) );
  XOR U16823 ( .A(n16711), .B(n11782), .Z(n6922) );
  XNOR U16824 ( .A(n13601), .B(n16231), .Z(n11782) );
  XNOR U16825 ( .A(n17498), .B(n17499), .Z(n16231) );
  XNOR U16826 ( .A(n11967), .B(n16592), .Z(n17499) );
  XOR U16827 ( .A(n17500), .B(n15935), .Z(n16592) );
  XOR U16828 ( .A(n17501), .B(n17502), .Z(n15935) );
  AND U16829 ( .A(n16713), .B(n16715), .Z(n17500) );
  XNOR U16830 ( .A(n17503), .B(n17504), .Z(n16715) );
  XNOR U16831 ( .A(n17505), .B(n17506), .Z(n16713) );
  XOR U16832 ( .A(n17507), .B(n15938), .Z(n11967) );
  XNOR U16833 ( .A(n17508), .B(n17509), .Z(n15938) );
  AND U16834 ( .A(n17032), .B(n17018), .Z(n17507) );
  IV U16835 ( .A(n17510), .Z(n17018) );
  XOR U16836 ( .A(n17026), .B(n17511), .Z(n17498) );
  XNOR U16837 ( .A(n16441), .B(n10267), .Z(n17511) );
  XOR U16838 ( .A(n17512), .B(n15929), .Z(n10267) );
  XOR U16839 ( .A(n17513), .B(n17514), .Z(n15929) );
  AND U16840 ( .A(n16721), .B(n17014), .Z(n17512) );
  XOR U16841 ( .A(n17515), .B(n16842), .Z(n17014) );
  IV U16842 ( .A(n16362), .Z(n16842) );
  XNOR U16843 ( .A(n17516), .B(n17517), .Z(n16721) );
  XNOR U16844 ( .A(n17518), .B(n15926), .Z(n16441) );
  XOR U16845 ( .A(n17519), .B(n17520), .Z(n15926) );
  ANDN U16846 ( .B(n16719), .A(n16718), .Z(n17518) );
  XNOR U16847 ( .A(n17521), .B(n17522), .Z(n16718) );
  XNOR U16848 ( .A(n17524), .B(n15943), .Z(n17026) );
  XNOR U16849 ( .A(n17525), .B(n16669), .Z(n15943) );
  ANDN U16850 ( .B(n16724), .A(n16725), .Z(n17524) );
  XOR U16851 ( .A(n17526), .B(n15222), .Z(n16725) );
  XNOR U16852 ( .A(n17272), .B(n17527), .Z(n16724) );
  IV U16853 ( .A(n16903), .Z(n17272) );
  XOR U16854 ( .A(n17528), .B(n17529), .Z(n13601) );
  XNOR U16855 ( .A(n17530), .B(n11854), .Z(n17529) );
  XOR U16856 ( .A(n17531), .B(n13932), .Z(n11854) );
  IV U16857 ( .A(n17532), .Z(n13932) );
  ANDN U16858 ( .B(n13097), .A(n15202), .Z(n17531) );
  XNOR U16859 ( .A(n17533), .B(n17534), .Z(n13097) );
  XOR U16860 ( .A(n13113), .B(n17535), .Z(n17528) );
  XOR U16861 ( .A(n10007), .B(n17536), .Z(n17535) );
  XNOR U16862 ( .A(n17537), .B(n13926), .Z(n10007) );
  XOR U16863 ( .A(n17538), .B(n16995), .Z(n14466) );
  XNOR U16864 ( .A(n17539), .B(n13930), .Z(n13113) );
  AND U16865 ( .A(n13101), .B(n17540), .Z(n17539) );
  IV U16866 ( .A(n15220), .Z(n13101) );
  XNOR U16867 ( .A(n17541), .B(n17407), .Z(n15220) );
  XNOR U16868 ( .A(n17542), .B(n17032), .Z(n16711) );
  XNOR U16869 ( .A(n17543), .B(n14948), .Z(n17032) );
  AND U16870 ( .A(n15937), .B(n17510), .Z(n17542) );
  XOR U16871 ( .A(n17544), .B(n13883), .Z(n17510) );
  XOR U16872 ( .A(n17545), .B(n17546), .Z(n15937) );
  NOR U16873 ( .A(n9303), .B(n10480), .Z(n17497) );
  XNOR U16874 ( .A(n11376), .B(n14483), .Z(n10480) );
  XNOR U16875 ( .A(n17547), .B(n16282), .Z(n14483) );
  ANDN U16876 ( .B(n17548), .A(n15468), .Z(n17547) );
  XOR U16877 ( .A(n15949), .B(n15537), .Z(n11376) );
  XOR U16878 ( .A(n17549), .B(n17550), .Z(n15537) );
  XNOR U16879 ( .A(n16247), .B(n11821), .Z(n17550) );
  XOR U16880 ( .A(n17551), .B(n15465), .Z(n11821) );
  AND U16881 ( .A(n14487), .B(n14485), .Z(n17551) );
  XOR U16882 ( .A(n17554), .B(n17555), .Z(n14485) );
  XNOR U16883 ( .A(n17556), .B(n15462), .Z(n16247) );
  XNOR U16884 ( .A(n17557), .B(n17558), .Z(n15462) );
  ANDN U16885 ( .B(n14479), .A(n14480), .Z(n17556) );
  XOR U16886 ( .A(n17559), .B(n17560), .Z(n14479) );
  XNOR U16887 ( .A(n13073), .B(n17561), .Z(n17549) );
  XOR U16888 ( .A(n11313), .B(n10678), .Z(n17561) );
  XNOR U16889 ( .A(n17562), .B(n15458), .Z(n10678) );
  NOR U16890 ( .A(n14476), .B(n14475), .Z(n17562) );
  XOR U16891 ( .A(n17565), .B(n17566), .Z(n14475) );
  XNOR U16892 ( .A(n17567), .B(n15469), .Z(n11313) );
  XOR U16893 ( .A(n15917), .B(n17568), .Z(n15469) );
  ANDN U16894 ( .B(n16282), .A(n17548), .Z(n17567) );
  XOR U16895 ( .A(n17569), .B(n17570), .Z(n16282) );
  XNOR U16896 ( .A(n17571), .B(n15455), .Z(n13073) );
  XOR U16897 ( .A(n17572), .B(n16069), .Z(n15455) );
  AND U16898 ( .A(n14491), .B(n14489), .Z(n17571) );
  XNOR U16899 ( .A(n15831), .B(n17573), .Z(n14489) );
  XOR U16900 ( .A(n17574), .B(n17575), .Z(n15949) );
  XNOR U16901 ( .A(n12790), .B(n9921), .Z(n17575) );
  XNOR U16902 ( .A(n17576), .B(n15487), .Z(n9921) );
  XNOR U16903 ( .A(n17577), .B(n15655), .Z(n15487) );
  NOR U16904 ( .A(n15026), .B(n16253), .Z(n17576) );
  XOR U16905 ( .A(n17491), .B(n17578), .Z(n16253) );
  XNOR U16906 ( .A(n15831), .B(n17579), .Z(n15026) );
  XOR U16907 ( .A(n17580), .B(n15475), .Z(n12790) );
  IV U16908 ( .A(n16266), .Z(n15475) );
  XOR U16909 ( .A(n17581), .B(n15954), .Z(n16266) );
  NOR U16910 ( .A(n16772), .B(n16265), .Z(n17580) );
  XOR U16911 ( .A(n17582), .B(n17583), .Z(n16265) );
  XOR U16912 ( .A(n17584), .B(n17585), .Z(n16772) );
  XOR U16913 ( .A(n11735), .B(n17586), .Z(n17574) );
  XOR U16914 ( .A(n11430), .B(n13745), .Z(n17586) );
  XNOR U16915 ( .A(n17587), .B(n15485), .Z(n13745) );
  XNOR U16916 ( .A(n17588), .B(n17589), .Z(n15485) );
  ANDN U16917 ( .B(n15019), .A(n16257), .Z(n17587) );
  XOR U16918 ( .A(n17590), .B(n17520), .Z(n16257) );
  IV U16919 ( .A(n16765), .Z(n15019) );
  XNOR U16920 ( .A(n15913), .B(n17591), .Z(n16765) );
  XNOR U16921 ( .A(n17592), .B(n15483), .Z(n11430) );
  XNOR U16922 ( .A(n17593), .B(n15222), .Z(n15483) );
  AND U16923 ( .A(n16270), .B(n15015), .Z(n17592) );
  IV U16924 ( .A(n16761), .Z(n15015) );
  XOR U16925 ( .A(n17594), .B(n17595), .Z(n16761) );
  XOR U16926 ( .A(n17596), .B(n17270), .Z(n16270) );
  XNOR U16927 ( .A(n17597), .B(n15479), .Z(n11735) );
  XOR U16928 ( .A(n17598), .B(n14951), .Z(n15479) );
  ANDN U16929 ( .B(n16769), .A(n16246), .Z(n17597) );
  XNOR U16930 ( .A(n17599), .B(n16896), .Z(n16246) );
  IV U16931 ( .A(n16262), .Z(n16769) );
  XOR U16932 ( .A(n17600), .B(n17380), .Z(n16262) );
  XOR U16933 ( .A(n13359), .B(n17601), .Z(n9303) );
  IV U16934 ( .A(n9069), .Z(n13359) );
  XOR U16935 ( .A(n13111), .B(n12622), .Z(n9069) );
  XNOR U16936 ( .A(n17602), .B(n17603), .Z(n12622) );
  XNOR U16937 ( .A(n12831), .B(n12254), .Z(n17603) );
  XOR U16938 ( .A(n17604), .B(n17605), .Z(n12254) );
  ANDN U16939 ( .B(n17606), .A(n12399), .Z(n17604) );
  XNOR U16940 ( .A(n17607), .B(n16088), .Z(n12831) );
  IV U16941 ( .A(n17608), .Z(n13653) );
  XOR U16942 ( .A(n12340), .B(n17609), .Z(n17602) );
  XNOR U16943 ( .A(n10047), .B(n13384), .Z(n17609) );
  XOR U16944 ( .A(n17610), .B(n17611), .Z(n13384) );
  NOR U16945 ( .A(n16077), .B(n17612), .Z(n17610) );
  XNOR U16946 ( .A(n17613), .B(n17614), .Z(n10047) );
  NOR U16947 ( .A(n16085), .B(n14400), .Z(n17613) );
  XNOR U16948 ( .A(n17615), .B(n16080), .Z(n12340) );
  AND U16949 ( .A(n16081), .B(n12410), .Z(n17615) );
  IV U16950 ( .A(n17616), .Z(n12410) );
  XOR U16951 ( .A(n17617), .B(n17618), .Z(n13111) );
  XNOR U16952 ( .A(n9369), .B(n16072), .Z(n17618) );
  XOR U16953 ( .A(n17619), .B(n14505), .Z(n16072) );
  IV U16954 ( .A(n16102), .Z(n14505) );
  XOR U16955 ( .A(n17620), .B(n15213), .Z(n16102) );
  AND U16956 ( .A(n15992), .B(n17621), .Z(n17619) );
  XOR U16957 ( .A(n17622), .B(n14513), .Z(n9369) );
  XNOR U16958 ( .A(n17623), .B(n16067), .Z(n14513) );
  IV U16959 ( .A(n17451), .Z(n16067) );
  IV U16960 ( .A(n17624), .Z(n15998) );
  XNOR U16961 ( .A(n11835), .B(n17625), .Z(n17617) );
  XNOR U16962 ( .A(n9774), .B(n10554), .Z(n17625) );
  XNOR U16963 ( .A(n17626), .B(n14509), .Z(n10554) );
  XNOR U16964 ( .A(n17627), .B(n17483), .Z(n14509) );
  ANDN U16965 ( .B(n17628), .A(n17629), .Z(n17626) );
  XOR U16966 ( .A(n17630), .B(n14518), .Z(n9774) );
  IV U16967 ( .A(n16105), .Z(n14518) );
  XOR U16968 ( .A(n15958), .B(n17631), .Z(n16105) );
  AND U16969 ( .A(n15996), .B(n16106), .Z(n17630) );
  XNOR U16970 ( .A(n17632), .B(n14501), .Z(n11835) );
  XOR U16971 ( .A(n17633), .B(n17634), .Z(n14501) );
  ANDN U16972 ( .B(n16108), .A(n16317), .Z(n17632) );
  XOR U16973 ( .A(n17635), .B(n9310), .Z(n3522) );
  IV U16974 ( .A(n10585), .Z(n9310) );
  XNOR U16975 ( .A(n17636), .B(n11369), .Z(n10585) );
  XNOR U16976 ( .A(n15316), .B(n17637), .Z(n11369) );
  XOR U16977 ( .A(n17638), .B(n17639), .Z(n15316) );
  XOR U16978 ( .A(n11637), .B(n12607), .Z(n17639) );
  XOR U16979 ( .A(n17640), .B(n17641), .Z(n12607) );
  ANDN U16980 ( .B(n17642), .A(n15676), .Z(n17640) );
  XNOR U16981 ( .A(n17643), .B(n17644), .Z(n11637) );
  ANDN U16982 ( .B(n15667), .A(n17645), .Z(n17643) );
  XOR U16983 ( .A(n11172), .B(n17646), .Z(n17638) );
  XOR U16984 ( .A(n17647), .B(n12384), .Z(n17646) );
  XOR U16985 ( .A(n17648), .B(n17649), .Z(n12384) );
  NOR U16986 ( .A(n15672), .B(n17650), .Z(n17648) );
  XNOR U16987 ( .A(n17651), .B(n17652), .Z(n11172) );
  NOR U16988 ( .A(n9296), .B(n10471), .Z(n17635) );
  XNOR U16989 ( .A(n12396), .B(n11894), .Z(n10471) );
  IV U16990 ( .A(n14398), .Z(n11894) );
  XOR U16991 ( .A(n17654), .B(n17655), .Z(n14398) );
  XNOR U16992 ( .A(n17656), .B(n17612), .Z(n12396) );
  NOR U16993 ( .A(n16076), .B(n17657), .Z(n17656) );
  XOR U16994 ( .A(n10695), .B(n14969), .Z(n9296) );
  XNOR U16995 ( .A(n17658), .B(n17659), .Z(n14969) );
  AND U16996 ( .A(n13439), .B(n13441), .Z(n17658) );
  XOR U16997 ( .A(n17660), .B(n17661), .Z(n13441) );
  XOR U16998 ( .A(n14125), .B(n17662), .Z(n10695) );
  XOR U16999 ( .A(n17663), .B(n17664), .Z(n14125) );
  XNOR U17000 ( .A(n12992), .B(n12555), .Z(n17664) );
  XNOR U17001 ( .A(n17665), .B(n16508), .Z(n12555) );
  ANDN U17002 ( .B(n14840), .A(n14841), .Z(n17665) );
  XNOR U17003 ( .A(n17666), .B(n17667), .Z(n14840) );
  XNOR U17004 ( .A(n17668), .B(n13261), .Z(n12992) );
  XNOR U17005 ( .A(n17669), .B(n17661), .Z(n13261) );
  AND U17006 ( .A(n14833), .B(n17670), .Z(n17668) );
  XOR U17007 ( .A(n16751), .B(n17671), .Z(n14833) );
  XNOR U17008 ( .A(n11521), .B(n17672), .Z(n17663) );
  XOR U17009 ( .A(n15536), .B(n15683), .Z(n17672) );
  XNOR U17010 ( .A(n17673), .B(n13266), .Z(n15683) );
  XNOR U17011 ( .A(n17674), .B(n15623), .Z(n13266) );
  ANDN U17012 ( .B(n14847), .A(n14848), .Z(n17673) );
  XNOR U17013 ( .A(n17220), .B(n17675), .Z(n14847) );
  XOR U17014 ( .A(n17676), .B(n13256), .Z(n15536) );
  XNOR U17015 ( .A(n17677), .B(n17678), .Z(n13256) );
  AND U17016 ( .A(n14844), .B(n14845), .Z(n17676) );
  XNOR U17017 ( .A(n17679), .B(n17680), .Z(n14844) );
  XNOR U17018 ( .A(n17681), .B(n13251), .Z(n11521) );
  XOR U17019 ( .A(n17682), .B(n17683), .Z(n13251) );
  ANDN U17020 ( .B(n14836), .A(n14837), .Z(n17681) );
  XOR U17021 ( .A(n17684), .B(n17685), .Z(n14836) );
  XOR U17022 ( .A(n17686), .B(n6918), .Z(n2644) );
  XOR U17023 ( .A(n10830), .B(n17687), .Z(n6918) );
  XNOR U17024 ( .A(n17688), .B(n17689), .Z(n14546) );
  XNOR U17025 ( .A(n11792), .B(n17690), .Z(n17689) );
  XOR U17026 ( .A(n17691), .B(n17316), .Z(n11792) );
  ANDN U17027 ( .B(n17692), .A(n17693), .Z(n17691) );
  XNOR U17028 ( .A(n13283), .B(n17694), .Z(n17688) );
  XOR U17029 ( .A(n17695), .B(n14566), .Z(n17694) );
  XNOR U17030 ( .A(n17696), .B(n17320), .Z(n14566) );
  ANDN U17031 ( .B(n17697), .A(n17698), .Z(n17696) );
  XOR U17032 ( .A(n17699), .B(n17312), .Z(n13283) );
  XNOR U17033 ( .A(n17702), .B(n17703), .Z(n11278) );
  XOR U17034 ( .A(n9905), .B(n11730), .Z(n17703) );
  XNOR U17035 ( .A(n17704), .B(n16485), .Z(n11730) );
  NOR U17036 ( .A(n14719), .B(n14718), .Z(n17704) );
  XOR U17037 ( .A(n17705), .B(n16493), .Z(n9905) );
  AND U17038 ( .A(n14723), .B(n14722), .Z(n17705) );
  XOR U17039 ( .A(n10643), .B(n17706), .Z(n17702) );
  XOR U17040 ( .A(n11864), .B(n10816), .Z(n17706) );
  XNOR U17041 ( .A(n17707), .B(n16512), .Z(n10816) );
  ANDN U17042 ( .B(n14727), .A(n14728), .Z(n17707) );
  XNOR U17043 ( .A(n17708), .B(n17709), .Z(n11864) );
  ANDN U17044 ( .B(n14731), .A(n14732), .Z(n17708) );
  XOR U17045 ( .A(n17710), .B(n16490), .Z(n10643) );
  ANDN U17046 ( .B(n14735), .A(n14736), .Z(n17710) );
  ANDN U17047 ( .B(n9308), .A(n10476), .Z(n17686) );
  XOR U17048 ( .A(n10704), .B(n14781), .Z(n10476) );
  XOR U17049 ( .A(n17711), .B(n17712), .Z(n14781) );
  ANDN U17050 ( .B(n17713), .A(n14354), .Z(n17711) );
  XOR U17051 ( .A(n13600), .B(n14404), .Z(n10704) );
  XOR U17052 ( .A(n17714), .B(n17715), .Z(n14404) );
  XOR U17053 ( .A(n13857), .B(n14000), .Z(n17715) );
  XOR U17054 ( .A(n17716), .B(n14384), .Z(n14000) );
  XOR U17055 ( .A(n14944), .B(n17717), .Z(n14384) );
  ANDN U17056 ( .B(n15289), .A(n15290), .Z(n17716) );
  XNOR U17057 ( .A(n17718), .B(n17719), .Z(n15289) );
  XOR U17058 ( .A(n17720), .B(n14394), .Z(n13857) );
  IV U17059 ( .A(n16209), .Z(n14394) );
  XOR U17060 ( .A(n17721), .B(n17472), .Z(n16209) );
  AND U17061 ( .A(n15286), .B(n17722), .Z(n17720) );
  XNOR U17062 ( .A(n17723), .B(n15333), .Z(n15286) );
  XOR U17063 ( .A(n11707), .B(n17724), .Z(n17714) );
  XNOR U17064 ( .A(n15581), .B(n11655), .Z(n17724) );
  XNOR U17065 ( .A(n17725), .B(n14379), .Z(n11655) );
  XNOR U17066 ( .A(n15329), .B(n17726), .Z(n14379) );
  NOR U17067 ( .A(n15296), .B(n15297), .Z(n17725) );
  XNOR U17068 ( .A(n16416), .B(n17727), .Z(n15296) );
  XNOR U17069 ( .A(n17728), .B(n14375), .Z(n15581) );
  IV U17070 ( .A(n16207), .Z(n14375) );
  XOR U17071 ( .A(n17729), .B(n17730), .Z(n16207) );
  NOR U17072 ( .A(n15300), .B(n15299), .Z(n17728) );
  XNOR U17073 ( .A(n17731), .B(n17732), .Z(n15299) );
  XOR U17074 ( .A(n17733), .B(n14387), .Z(n11707) );
  XNOR U17075 ( .A(n17734), .B(n17735), .Z(n14387) );
  AND U17076 ( .A(n15293), .B(n17736), .Z(n17733) );
  XNOR U17077 ( .A(n17737), .B(n16523), .Z(n15293) );
  XOR U17078 ( .A(n17738), .B(n17739), .Z(n13600) );
  XOR U17079 ( .A(n16198), .B(n11119), .Z(n17739) );
  XOR U17080 ( .A(n17740), .B(n17741), .Z(n11119) );
  NOR U17081 ( .A(n14790), .B(n14791), .Z(n17740) );
  XOR U17082 ( .A(n17742), .B(n14361), .Z(n16198) );
  AND U17083 ( .A(n14794), .B(n14795), .Z(n17742) );
  XOR U17084 ( .A(n11885), .B(n17743), .Z(n17738) );
  XOR U17085 ( .A(n11071), .B(n12912), .Z(n17743) );
  XOR U17086 ( .A(n17744), .B(n14369), .Z(n12912) );
  NOR U17087 ( .A(n14787), .B(n14788), .Z(n17744) );
  XNOR U17088 ( .A(n17745), .B(n14356), .Z(n11071) );
  ANDN U17089 ( .B(n17712), .A(n17713), .Z(n17745) );
  XNOR U17090 ( .A(n17746), .B(n14365), .Z(n11885) );
  AND U17091 ( .A(n14783), .B(n17747), .Z(n17746) );
  XOR U17092 ( .A(n14633), .B(n9573), .Z(n9308) );
  XNOR U17093 ( .A(n17748), .B(n16211), .Z(n9573) );
  XNOR U17094 ( .A(n17749), .B(n17750), .Z(n16211) );
  XNOR U17095 ( .A(n12693), .B(n12333), .Z(n17750) );
  XOR U17096 ( .A(n17751), .B(n13843), .Z(n12333) );
  AND U17097 ( .A(n17752), .B(n17753), .Z(n17751) );
  XNOR U17098 ( .A(n17754), .B(n17755), .Z(n12693) );
  XOR U17099 ( .A(n11438), .B(n17758), .Z(n17749) );
  XOR U17100 ( .A(n16595), .B(n11165), .Z(n17758) );
  XNOR U17101 ( .A(n17759), .B(n17760), .Z(n11165) );
  NOR U17102 ( .A(n17761), .B(n17762), .Z(n17759) );
  XOR U17103 ( .A(n17763), .B(n14193), .Z(n16595) );
  IV U17104 ( .A(n17764), .Z(n14193) );
  ANDN U17105 ( .B(n17765), .A(n17766), .Z(n17763) );
  XOR U17106 ( .A(n17767), .B(n15052), .Z(n11438) );
  XOR U17107 ( .A(n17770), .B(n17771), .Z(n14633) );
  NOR U17108 ( .A(n14074), .B(n16837), .Z(n17770) );
  AND U17109 ( .A(n4065), .B(n2597), .Z(n16844) );
  XNOR U17110 ( .A(n7589), .B(n2610), .Z(n2597) );
  XNOR U17111 ( .A(n5931), .B(n6348), .Z(n2610) );
  XNOR U17112 ( .A(n17773), .B(n17774), .Z(n6348) );
  XOR U17113 ( .A(n2646), .B(n5333), .Z(n17774) );
  XOR U17114 ( .A(n17775), .B(n7503), .Z(n5333) );
  IV U17115 ( .A(n6804), .Z(n7503) );
  XOR U17116 ( .A(n16083), .B(n10603), .Z(n6804) );
  XNOR U17117 ( .A(n13606), .B(n12844), .Z(n10603) );
  XNOR U17118 ( .A(n17776), .B(n17777), .Z(n12844) );
  XOR U17119 ( .A(n10150), .B(n13116), .Z(n17777) );
  XNOR U17120 ( .A(n17778), .B(n17779), .Z(n13116) );
  ANDN U17121 ( .B(n15378), .A(n15376), .Z(n17778) );
  XNOR U17122 ( .A(n17780), .B(n14043), .Z(n10150) );
  AND U17123 ( .A(n14044), .B(n17781), .Z(n17780) );
  XOR U17124 ( .A(n17782), .B(n17735), .Z(n14044) );
  IV U17125 ( .A(n17045), .Z(n17735) );
  XNOR U17126 ( .A(n14030), .B(n17783), .Z(n17776) );
  XOR U17127 ( .A(n12481), .B(n12572), .Z(n17783) );
  XNOR U17128 ( .A(n17784), .B(n14542), .Z(n12572) );
  AND U17129 ( .A(n15389), .B(n14541), .Z(n17784) );
  IV U17130 ( .A(n15387), .Z(n14541) );
  XOR U17131 ( .A(n17785), .B(n17786), .Z(n15387) );
  XNOR U17132 ( .A(n17787), .B(n14047), .Z(n12481) );
  AND U17133 ( .A(n15374), .B(n14048), .Z(n17787) );
  XNOR U17134 ( .A(n17788), .B(n15655), .Z(n14048) );
  XNOR U17135 ( .A(n17789), .B(n14038), .Z(n14030) );
  AND U17136 ( .A(n14037), .B(n17790), .Z(n17789) );
  XNOR U17137 ( .A(n17791), .B(n17792), .Z(n14037) );
  XOR U17138 ( .A(n17793), .B(n17794), .Z(n13606) );
  XNOR U17139 ( .A(n10671), .B(n9898), .Z(n17794) );
  XNOR U17140 ( .A(n17795), .B(n17657), .Z(n9898) );
  AND U17141 ( .A(n16076), .B(n17611), .Z(n17795) );
  IV U17142 ( .A(n16078), .Z(n17611) );
  XOR U17143 ( .A(n17796), .B(n16896), .Z(n16078) );
  XNOR U17144 ( .A(n17797), .B(n17045), .Z(n16076) );
  XOR U17145 ( .A(n17798), .B(n14401), .Z(n10671) );
  AND U17146 ( .A(n14402), .B(n17614), .Z(n17798) );
  IV U17147 ( .A(n16086), .Z(n17614) );
  XNOR U17148 ( .A(n17799), .B(n17800), .Z(n16086) );
  XOR U17149 ( .A(n17801), .B(n17802), .Z(n14402) );
  XNOR U17150 ( .A(n10652), .B(n17803), .Z(n17793) );
  XOR U17151 ( .A(n9497), .B(n9087), .Z(n17803) );
  XOR U17152 ( .A(n17804), .B(n13655), .Z(n9087) );
  NOR U17153 ( .A(n13654), .B(n16088), .Z(n17804) );
  XOR U17154 ( .A(n17805), .B(n13991), .Z(n16088) );
  XOR U17155 ( .A(n17806), .B(n17560), .Z(n13654) );
  XNOR U17156 ( .A(n17807), .B(n12411), .Z(n9497) );
  ANDN U17157 ( .B(n12412), .A(n16080), .Z(n17807) );
  XNOR U17158 ( .A(n17808), .B(n17809), .Z(n16080) );
  XNOR U17159 ( .A(n17810), .B(n17811), .Z(n12412) );
  XOR U17160 ( .A(n17812), .B(n12401), .Z(n10652) );
  AND U17161 ( .A(n12400), .B(n17605), .Z(n17812) );
  IV U17162 ( .A(n17813), .Z(n17605) );
  XNOR U17163 ( .A(n17814), .B(n12400), .Z(n16083) );
  XNOR U17164 ( .A(n17815), .B(n17816), .Z(n12400) );
  ANDN U17165 ( .B(n17813), .A(n17606), .Z(n17814) );
  XNOR U17166 ( .A(n17817), .B(n16252), .Z(n17813) );
  NOR U17167 ( .A(n7599), .B(n6803), .Z(n17775) );
  XOR U17168 ( .A(n10377), .B(n17818), .Z(n6803) );
  IV U17169 ( .A(n10162), .Z(n10377) );
  XOR U17170 ( .A(n14878), .B(n14627), .Z(n10162) );
  XOR U17171 ( .A(n17819), .B(n17820), .Z(n14627) );
  XOR U17172 ( .A(n11836), .B(n9495), .Z(n17820) );
  XOR U17173 ( .A(n17821), .B(n17766), .Z(n9495) );
  AND U17174 ( .A(n14192), .B(n17822), .Z(n17821) );
  XNOR U17175 ( .A(n17823), .B(n17757), .Z(n11836) );
  NOR U17176 ( .A(n17756), .B(n17824), .Z(n17823) );
  XNOR U17177 ( .A(n16210), .B(n17825), .Z(n17819) );
  XOR U17178 ( .A(n14998), .B(n12451), .Z(n17825) );
  XNOR U17179 ( .A(n17826), .B(n17827), .Z(n12451) );
  NOR U17180 ( .A(n17752), .B(n13841), .Z(n17826) );
  XNOR U17181 ( .A(n17828), .B(n17762), .Z(n14998) );
  AND U17182 ( .A(n17761), .B(n17829), .Z(n17828) );
  XNOR U17183 ( .A(n17830), .B(n17769), .Z(n16210) );
  ANDN U17184 ( .B(n17768), .A(n15050), .Z(n17830) );
  XOR U17185 ( .A(n17831), .B(n17832), .Z(n14878) );
  XOR U17186 ( .A(n10151), .B(n9993), .Z(n17832) );
  XOR U17187 ( .A(n17833), .B(n16216), .Z(n9993) );
  XNOR U17188 ( .A(n17834), .B(n17835), .Z(n16216) );
  IV U17189 ( .A(n17836), .Z(n16189) );
  XOR U17190 ( .A(n17837), .B(n16979), .Z(n10151) );
  XNOR U17191 ( .A(n17838), .B(n16698), .Z(n16979) );
  AND U17192 ( .A(n17008), .B(n16172), .Z(n17837) );
  XOR U17193 ( .A(n9365), .B(n17839), .Z(n17831) );
  XOR U17194 ( .A(n10175), .B(n15029), .Z(n17839) );
  XNOR U17195 ( .A(n17840), .B(n16220), .Z(n15029) );
  XNOR U17196 ( .A(n17841), .B(n17842), .Z(n16220) );
  NOR U17197 ( .A(n16185), .B(n16221), .Z(n17840) );
  XOR U17198 ( .A(n17843), .B(n16976), .Z(n10175) );
  IV U17199 ( .A(n16223), .Z(n16976) );
  XOR U17200 ( .A(n15132), .B(n17844), .Z(n16223) );
  ANDN U17201 ( .B(n16224), .A(n16181), .Z(n17843) );
  XNOR U17202 ( .A(n17845), .B(n16228), .Z(n9365) );
  XOR U17203 ( .A(n17846), .B(n17847), .Z(n16228) );
  ANDN U17204 ( .B(n16176), .A(n16227), .Z(n17845) );
  XNOR U17205 ( .A(n16400), .B(n10022), .Z(n7599) );
  IV U17206 ( .A(n13391), .Z(n10022) );
  XOR U17207 ( .A(n15813), .B(n17298), .Z(n13391) );
  XNOR U17208 ( .A(n17848), .B(n17849), .Z(n17298) );
  XNOR U17209 ( .A(n10545), .B(n14663), .Z(n17849) );
  XNOR U17210 ( .A(n17850), .B(n16573), .Z(n14663) );
  XNOR U17211 ( .A(n17851), .B(n17589), .Z(n16573) );
  NOR U17212 ( .A(n16403), .B(n16402), .Z(n17850) );
  XNOR U17213 ( .A(n17852), .B(n16940), .Z(n16402) );
  XNOR U17214 ( .A(n17853), .B(n16568), .Z(n10545) );
  XNOR U17215 ( .A(n17854), .B(n17855), .Z(n16568) );
  ANDN U17216 ( .B(n16392), .A(n16393), .Z(n17853) );
  XNOR U17217 ( .A(n17856), .B(n17857), .Z(n16392) );
  XOR U17218 ( .A(n16846), .B(n17858), .Z(n17848) );
  XOR U17219 ( .A(n11057), .B(n12679), .Z(n17858) );
  XNOR U17220 ( .A(n17859), .B(n16576), .Z(n12679) );
  XOR U17221 ( .A(n17860), .B(n17861), .Z(n16576) );
  ANDN U17222 ( .B(n16854), .A(n16397), .Z(n17859) );
  XOR U17223 ( .A(n17862), .B(n16014), .Z(n16854) );
  XOR U17224 ( .A(n17863), .B(n16578), .Z(n11057) );
  XNOR U17225 ( .A(n17864), .B(n14948), .Z(n16578) );
  AND U17226 ( .A(n16406), .B(n17865), .Z(n17863) );
  XNOR U17227 ( .A(n17553), .B(n17866), .Z(n16406) );
  XNOR U17228 ( .A(n17867), .B(n16565), .Z(n16846) );
  XNOR U17229 ( .A(n17868), .B(n17869), .Z(n16565) );
  XOR U17230 ( .A(n17871), .B(n17872), .Z(n15813) );
  XOR U17231 ( .A(n12288), .B(n10273), .Z(n17872) );
  XNOR U17232 ( .A(n17873), .B(n16865), .Z(n10273) );
  AND U17233 ( .A(n16384), .B(n16866), .Z(n17873) );
  XOR U17234 ( .A(n17874), .B(n17583), .Z(n16866) );
  XNOR U17235 ( .A(n17875), .B(n15533), .Z(n16384) );
  IV U17236 ( .A(n17876), .Z(n15533) );
  XOR U17237 ( .A(n17877), .B(n16875), .Z(n12288) );
  ANDN U17238 ( .B(n16876), .A(n16379), .Z(n17877) );
  XNOR U17239 ( .A(n17878), .B(n17879), .Z(n16379) );
  XNOR U17240 ( .A(n17880), .B(n13896), .Z(n16876) );
  XNOR U17241 ( .A(n12251), .B(n17881), .Z(n17871) );
  XOR U17242 ( .A(n12627), .B(n10988), .Z(n17881) );
  XOR U17243 ( .A(n17882), .B(n17883), .Z(n10988) );
  ANDN U17244 ( .B(n16369), .A(n16370), .Z(n17882) );
  XNOR U17245 ( .A(n17884), .B(n17360), .Z(n16370) );
  XNOR U17246 ( .A(n17885), .B(n16862), .Z(n12627) );
  XOR U17247 ( .A(n17886), .B(n16698), .Z(n16374) );
  XOR U17248 ( .A(n17887), .B(n17888), .Z(n16373) );
  XOR U17249 ( .A(n17889), .B(n16871), .Z(n12251) );
  ANDN U17250 ( .B(n16872), .A(n16387), .Z(n17889) );
  XNOR U17251 ( .A(n17890), .B(n16041), .Z(n16387) );
  XOR U17252 ( .A(n17891), .B(n17892), .Z(n16872) );
  XOR U17253 ( .A(n17893), .B(n16856), .Z(n16400) );
  XOR U17254 ( .A(n17894), .B(n17895), .Z(n16856) );
  AND U17255 ( .A(n17870), .B(n16564), .Z(n17893) );
  IV U17256 ( .A(n17896), .Z(n16564) );
  XNOR U17257 ( .A(n17897), .B(n6808), .Z(n2646) );
  XOR U17258 ( .A(n9892), .B(n16584), .Z(n6808) );
  XOR U17259 ( .A(n17898), .B(n14248), .Z(n16584) );
  NOR U17260 ( .A(n15071), .B(n15070), .Z(n17898) );
  XOR U17261 ( .A(n15392), .B(n17181), .Z(n9892) );
  XNOR U17262 ( .A(n17899), .B(n17900), .Z(n17181) );
  XNOR U17263 ( .A(n10364), .B(n14077), .Z(n17900) );
  XNOR U17264 ( .A(n17901), .B(n14233), .Z(n14077) );
  AND U17265 ( .A(n16588), .B(n14234), .Z(n17901) );
  XNOR U17266 ( .A(n17902), .B(n17903), .Z(n14234) );
  XNOR U17267 ( .A(n17904), .B(n15325), .Z(n16588) );
  XNOR U17268 ( .A(n17905), .B(n14237), .Z(n10364) );
  AND U17269 ( .A(n14238), .B(n15058), .Z(n17905) );
  XOR U17270 ( .A(n15824), .B(n17906), .Z(n15058) );
  XNOR U17271 ( .A(n17907), .B(n17908), .Z(n14238) );
  XOR U17272 ( .A(n10310), .B(n17909), .Z(n17899) );
  XOR U17273 ( .A(n11711), .B(n12406), .Z(n17909) );
  XNOR U17274 ( .A(n17910), .B(n17300), .Z(n12406) );
  XOR U17275 ( .A(n17911), .B(n17458), .Z(n15061) );
  XNOR U17276 ( .A(n17912), .B(n15603), .Z(n16590) );
  XOR U17277 ( .A(n17913), .B(n14247), .Z(n11711) );
  AND U17278 ( .A(n15070), .B(n14248), .Z(n17913) );
  XNOR U17279 ( .A(n17914), .B(n17915), .Z(n14248) );
  XNOR U17280 ( .A(n17916), .B(n16702), .Z(n15070) );
  IV U17281 ( .A(n17917), .Z(n16702) );
  XNOR U17282 ( .A(n17918), .B(n14243), .Z(n10310) );
  ANDN U17283 ( .B(n15067), .A(n14244), .Z(n17918) );
  XNOR U17284 ( .A(n17919), .B(n17678), .Z(n14244) );
  XNOR U17285 ( .A(n17920), .B(n16071), .Z(n15067) );
  XOR U17286 ( .A(n17921), .B(n17922), .Z(n15392) );
  XOR U17287 ( .A(n10910), .B(n10128), .Z(n17922) );
  XNOR U17288 ( .A(n17923), .B(n16397), .Z(n10128) );
  XOR U17289 ( .A(n17924), .B(n17925), .Z(n16397) );
  AND U17290 ( .A(n16398), .B(n16853), .Z(n17923) );
  IV U17291 ( .A(n16575), .Z(n16853) );
  XOR U17292 ( .A(n17926), .B(n17585), .Z(n16575) );
  XNOR U17293 ( .A(n17927), .B(n17928), .Z(n16398) );
  XOR U17294 ( .A(n17929), .B(n17870), .Z(n10910) );
  XOR U17295 ( .A(n17930), .B(n16016), .Z(n17870) );
  IV U17296 ( .A(n16674), .Z(n16016) );
  AND U17297 ( .A(n16566), .B(n17896), .Z(n17929) );
  XOR U17298 ( .A(n17931), .B(n17667), .Z(n17896) );
  XOR U17299 ( .A(n17932), .B(n17933), .Z(n16566) );
  XNOR U17300 ( .A(n16365), .B(n17934), .Z(n17921) );
  XOR U17301 ( .A(n12564), .B(n12139), .Z(n17934) );
  XOR U17302 ( .A(n17935), .B(n16408), .Z(n12139) );
  IV U17303 ( .A(n17865), .Z(n16408) );
  XOR U17304 ( .A(n17936), .B(n17937), .Z(n17865) );
  XNOR U17305 ( .A(n17938), .B(n16795), .Z(n16579) );
  XOR U17306 ( .A(n17939), .B(n17940), .Z(n16407) );
  XOR U17307 ( .A(n17941), .B(n16393), .Z(n12564) );
  XNOR U17308 ( .A(n17258), .B(n17942), .Z(n16393) );
  AND U17309 ( .A(n16569), .B(n16394), .Z(n17941) );
  XNOR U17310 ( .A(n16318), .B(n17943), .Z(n16394) );
  XOR U17311 ( .A(n17946), .B(n16403), .Z(n16365) );
  XOR U17312 ( .A(n17947), .B(n17948), .Z(n16403) );
  ANDN U17313 ( .B(n16404), .A(n16572), .Z(n17946) );
  XNOR U17314 ( .A(n17949), .B(n16523), .Z(n16572) );
  XNOR U17315 ( .A(n17950), .B(n16818), .Z(n16404) );
  IV U17316 ( .A(n17951), .Z(n16818) );
  ANDN U17317 ( .B(n9934), .A(n6807), .Z(n17897) );
  XNOR U17318 ( .A(n3312), .B(n17952), .Z(n17773) );
  XOR U17319 ( .A(n5315), .B(n6797), .Z(n17952) );
  XNOR U17320 ( .A(n17953), .B(n6812), .Z(n6797) );
  XNOR U17321 ( .A(n9537), .B(n13134), .Z(n6812) );
  XOR U17322 ( .A(n17954), .B(n13997), .Z(n13134) );
  ANDN U17323 ( .B(n17955), .A(n15898), .Z(n17954) );
  XOR U17324 ( .A(n14280), .B(n13375), .Z(n9537) );
  XOR U17325 ( .A(n17956), .B(n17957), .Z(n13375) );
  XOR U17326 ( .A(n13609), .B(n10936), .Z(n17957) );
  XOR U17327 ( .A(n17958), .B(n15894), .Z(n10936) );
  IV U17328 ( .A(n13623), .Z(n15894) );
  XNOR U17329 ( .A(n17959), .B(n17960), .Z(n13623) );
  NOR U17330 ( .A(n13137), .B(n13136), .Z(n17958) );
  XOR U17331 ( .A(n17961), .B(n17962), .Z(n13136) );
  XNOR U17332 ( .A(n17963), .B(n14013), .Z(n13609) );
  XNOR U17333 ( .A(n17964), .B(n17965), .Z(n14013) );
  XOR U17334 ( .A(n17966), .B(n15958), .Z(n13141) );
  XOR U17335 ( .A(n12174), .B(n17967), .Z(n17956) );
  XOR U17336 ( .A(n11841), .B(n9715), .Z(n17967) );
  XOR U17337 ( .A(n17968), .B(n17969), .Z(n9715) );
  NOR U17338 ( .A(n13150), .B(n13149), .Z(n17968) );
  XOR U17339 ( .A(n17970), .B(n16796), .Z(n13149) );
  XNOR U17340 ( .A(n17971), .B(n13615), .Z(n11841) );
  XNOR U17341 ( .A(n17972), .B(n17973), .Z(n13615) );
  XOR U17342 ( .A(n17974), .B(n17467), .Z(n13145) );
  XNOR U17343 ( .A(n17975), .B(n13996), .Z(n12174) );
  XNOR U17344 ( .A(n15913), .B(n17976), .Z(n13996) );
  XOR U17345 ( .A(n17977), .B(n17978), .Z(n13997) );
  XOR U17346 ( .A(n17979), .B(n17980), .Z(n14280) );
  XNOR U17347 ( .A(n10443), .B(n11529), .Z(n17980) );
  XOR U17348 ( .A(n17981), .B(n13637), .Z(n11529) );
  XOR U17349 ( .A(n17982), .B(n17972), .Z(n13637) );
  AND U17350 ( .A(n14592), .B(n14591), .Z(n17981) );
  XOR U17351 ( .A(n17983), .B(n17534), .Z(n14591) );
  XNOR U17352 ( .A(n17984), .B(n13646), .Z(n10443) );
  XOR U17353 ( .A(n17985), .B(n17879), .Z(n13646) );
  ANDN U17354 ( .B(n14594), .A(n13645), .Z(n17984) );
  XOR U17355 ( .A(n17986), .B(n17987), .Z(n13645) );
  XNOR U17356 ( .A(n9265), .B(n17988), .Z(n17979) );
  XOR U17357 ( .A(n9189), .B(n11676), .Z(n17988) );
  XNOR U17358 ( .A(n17989), .B(n13633), .Z(n11676) );
  XNOR U17359 ( .A(n17332), .B(n17990), .Z(n13633) );
  ANDN U17360 ( .B(n13632), .A(n14597), .Z(n17989) );
  XOR U17361 ( .A(n17991), .B(n15984), .Z(n13632) );
  XOR U17362 ( .A(n17992), .B(n13642), .Z(n9189) );
  IV U17363 ( .A(n14026), .Z(n13642) );
  XNOR U17364 ( .A(n17993), .B(n17994), .Z(n14026) );
  ANDN U17365 ( .B(n14599), .A(n13641), .Z(n17992) );
  XOR U17366 ( .A(n17995), .B(n17945), .Z(n13641) );
  XNOR U17367 ( .A(n17996), .B(n13629), .Z(n9265) );
  XNOR U17368 ( .A(n17997), .B(n17998), .Z(n13629) );
  ANDN U17369 ( .B(n13628), .A(n14601), .Z(n17996) );
  XNOR U17370 ( .A(n17841), .B(n17999), .Z(n13628) );
  AND U17371 ( .A(n7596), .B(n6813), .Z(n17953) );
  XOR U17372 ( .A(n10932), .B(n17263), .Z(n6813) );
  XOR U17373 ( .A(n18000), .B(n14746), .Z(n17263) );
  ANDN U17374 ( .B(n16315), .A(n16810), .Z(n18000) );
  XNOR U17375 ( .A(n18001), .B(n18002), .Z(n16315) );
  IV U17376 ( .A(n10772), .Z(n10932) );
  XOR U17377 ( .A(n18003), .B(n16197), .Z(n10772) );
  XNOR U17378 ( .A(n18004), .B(n18005), .Z(n16197) );
  XOR U17379 ( .A(n11752), .B(n11591), .Z(n18005) );
  XNOR U17380 ( .A(n18006), .B(n11948), .Z(n11591) );
  ANDN U17381 ( .B(n11949), .A(n17282), .Z(n18006) );
  XNOR U17382 ( .A(n18007), .B(n18008), .Z(n11949) );
  XNOR U17383 ( .A(n18009), .B(n11952), .Z(n11752) );
  XNOR U17384 ( .A(n18010), .B(n18011), .Z(n11952) );
  ANDN U17385 ( .B(n11953), .A(n17290), .Z(n18009) );
  XNOR U17386 ( .A(n15824), .B(n18012), .Z(n11953) );
  XNOR U17387 ( .A(n11422), .B(n18013), .Z(n18004) );
  XNOR U17388 ( .A(n9565), .B(n10578), .Z(n18013) );
  XOR U17389 ( .A(n18014), .B(n11966), .Z(n10578) );
  XNOR U17390 ( .A(n18015), .B(n18016), .Z(n11966) );
  AND U17391 ( .A(n17280), .B(n11965), .Z(n18014) );
  XNOR U17392 ( .A(n18017), .B(n18018), .Z(n11965) );
  XOR U17393 ( .A(n18019), .B(n11961), .Z(n9565) );
  XNOR U17394 ( .A(n18020), .B(n17809), .Z(n11961) );
  ANDN U17395 ( .B(n17286), .A(n11962), .Z(n18019) );
  XOR U17396 ( .A(n18021), .B(n18022), .Z(n11962) );
  XNOR U17397 ( .A(n18023), .B(n11957), .Z(n11422) );
  XNOR U17398 ( .A(n18024), .B(n17509), .Z(n11957) );
  ANDN U17399 ( .B(n11958), .A(n17288), .Z(n18023) );
  XOR U17400 ( .A(n18025), .B(n18026), .Z(n11958) );
  XNOR U17401 ( .A(n11045), .B(n17097), .Z(n7596) );
  XNOR U17402 ( .A(n18027), .B(n18028), .Z(n17097) );
  AND U17403 ( .A(n18029), .B(n18030), .Z(n18027) );
  XOR U17404 ( .A(n12686), .B(n13863), .Z(n11045) );
  XOR U17405 ( .A(n18031), .B(n18032), .Z(n13863) );
  XNOR U17406 ( .A(n9490), .B(n13282), .Z(n18032) );
  XNOR U17407 ( .A(n18033), .B(n17650), .Z(n13282) );
  ANDN U17408 ( .B(n15672), .A(n15673), .Z(n18033) );
  XNOR U17409 ( .A(n18034), .B(n18035), .Z(n15672) );
  XOR U17410 ( .A(n18036), .B(n18037), .Z(n9490) );
  ANDN U17411 ( .B(n15663), .A(n15664), .Z(n18036) );
  XNOR U17412 ( .A(n15315), .B(n18038), .Z(n18031) );
  XOR U17413 ( .A(n9100), .B(n10103), .Z(n18038) );
  XNOR U17414 ( .A(n18039), .B(n17653), .Z(n10103) );
  AND U17415 ( .A(n15680), .B(n18040), .Z(n18039) );
  XNOR U17416 ( .A(n18041), .B(n17341), .Z(n15680) );
  XNOR U17417 ( .A(n18042), .B(n17645), .Z(n9100) );
  NOR U17418 ( .A(n15669), .B(n15667), .Z(n18042) );
  XOR U17419 ( .A(n18045), .B(n17642), .Z(n15315) );
  AND U17420 ( .A(n15677), .B(n15676), .Z(n18045) );
  XOR U17421 ( .A(n18046), .B(n18047), .Z(n15676) );
  XOR U17422 ( .A(n18048), .B(n18049), .Z(n12686) );
  XNOR U17423 ( .A(n11582), .B(n11368), .Z(n18049) );
  XNOR U17424 ( .A(n18050), .B(n18051), .Z(n11368) );
  XOR U17425 ( .A(n18052), .B(n18053), .Z(n11582) );
  NOR U17426 ( .A(n18054), .B(n17104), .Z(n18052) );
  XOR U17427 ( .A(n17636), .B(n18055), .Z(n18048) );
  XNOR U17428 ( .A(n11603), .B(n11406), .Z(n18055) );
  XOR U17429 ( .A(n18056), .B(n18057), .Z(n11406) );
  ANDN U17430 ( .B(n18028), .A(n18029), .Z(n18056) );
  XNOR U17431 ( .A(n18058), .B(n18059), .Z(n11603) );
  ANDN U17432 ( .B(n17089), .A(n17090), .Z(n18058) );
  XOR U17433 ( .A(n18060), .B(n18061), .Z(n17636) );
  AND U17434 ( .A(n17095), .B(n17093), .Z(n18060) );
  XNOR U17435 ( .A(n18062), .B(n6817), .Z(n5315) );
  XNOR U17436 ( .A(n18063), .B(n10785), .Z(n6817) );
  XOR U17437 ( .A(n14759), .B(n13904), .Z(n10785) );
  XOR U17438 ( .A(n18064), .B(n18065), .Z(n13904) );
  XNOR U17439 ( .A(n11450), .B(n9202), .Z(n18065) );
  XOR U17440 ( .A(n18066), .B(n16654), .Z(n9202) );
  AND U17441 ( .A(n18067), .B(n15871), .Z(n18066) );
  XNOR U17442 ( .A(n18068), .B(n16652), .Z(n11450) );
  AND U17443 ( .A(n18069), .B(n15876), .Z(n18068) );
  XNOR U17444 ( .A(n18070), .B(n18071), .Z(n18064) );
  XNOR U17445 ( .A(n12530), .B(n12449), .Z(n18071) );
  XNOR U17446 ( .A(n18072), .B(n16656), .Z(n12449) );
  ANDN U17447 ( .B(n15880), .A(n18073), .Z(n18072) );
  XNOR U17448 ( .A(n18074), .B(n16645), .Z(n12530) );
  ANDN U17449 ( .B(n18075), .A(n15884), .Z(n18074) );
  XOR U17450 ( .A(n18076), .B(n18077), .Z(n14759) );
  XNOR U17451 ( .A(n12978), .B(n11685), .Z(n18077) );
  XNOR U17452 ( .A(n18078), .B(n14991), .Z(n11685) );
  ANDN U17453 ( .B(n16134), .A(n16135), .Z(n18078) );
  XOR U17454 ( .A(n18079), .B(n14994), .Z(n12978) );
  AND U17455 ( .A(n16138), .B(n16137), .Z(n18079) );
  XOR U17456 ( .A(n11827), .B(n18080), .Z(n18076) );
  XOR U17457 ( .A(n12549), .B(n12387), .Z(n18080) );
  XOR U17458 ( .A(n18081), .B(n18082), .Z(n12387) );
  ANDN U17459 ( .B(n16141), .A(n16142), .Z(n18081) );
  XNOR U17460 ( .A(n18083), .B(n14984), .Z(n12549) );
  IV U17461 ( .A(n18084), .Z(n14984) );
  AND U17462 ( .A(n16148), .B(n16149), .Z(n18083) );
  XOR U17463 ( .A(n18085), .B(n18086), .Z(n11827) );
  ANDN U17464 ( .B(n18087), .A(n16145), .Z(n18085) );
  ANDN U17465 ( .B(n9951), .A(n6816), .Z(n18062) );
  XNOR U17466 ( .A(n10229), .B(n16524), .Z(n6816) );
  XOR U17467 ( .A(n18088), .B(n18089), .Z(n16524) );
  ANDN U17468 ( .B(n15445), .A(n15266), .Z(n18088) );
  XOR U17469 ( .A(n18090), .B(n16691), .Z(n15266) );
  IV U17470 ( .A(n17389), .Z(n16691) );
  XOR U17471 ( .A(n15140), .B(n12327), .Z(n10229) );
  XNOR U17472 ( .A(n18091), .B(n18092), .Z(n12327) );
  XNOR U17473 ( .A(n12460), .B(n17109), .Z(n18092) );
  XNOR U17474 ( .A(n18093), .B(n15258), .Z(n17109) );
  XOR U17475 ( .A(n18094), .B(n18095), .Z(n15258) );
  AND U17476 ( .A(n13462), .B(n12757), .Z(n18093) );
  XOR U17477 ( .A(n18096), .B(n17197), .Z(n12757) );
  XNOR U17478 ( .A(n18097), .B(n16041), .Z(n13462) );
  XNOR U17479 ( .A(n18098), .B(n15250), .Z(n12460) );
  XNOR U17480 ( .A(n18099), .B(n18100), .Z(n15250) );
  ANDN U17481 ( .B(n12970), .A(n13457), .Z(n18098) );
  XNOR U17482 ( .A(n18101), .B(n18102), .Z(n13457) );
  XNOR U17483 ( .A(n18103), .B(n18104), .Z(n12970) );
  XOR U17484 ( .A(n11635), .B(n18105), .Z(n18091) );
  XNOR U17485 ( .A(n13595), .B(n9945), .Z(n18105) );
  XNOR U17486 ( .A(n18106), .B(n15241), .Z(n9945) );
  XNOR U17487 ( .A(n18107), .B(n16021), .Z(n15241) );
  ANDN U17488 ( .B(n12753), .A(n13459), .Z(n18106) );
  XOR U17489 ( .A(n18108), .B(n18109), .Z(n13459) );
  XOR U17490 ( .A(n18110), .B(n16995), .Z(n12753) );
  XNOR U17491 ( .A(n18111), .B(n15245), .Z(n13595) );
  XOR U17492 ( .A(n18112), .B(n18113), .Z(n15245) );
  ANDN U17493 ( .B(n13452), .A(n13450), .Z(n18111) );
  XOR U17494 ( .A(n18114), .B(n18115), .Z(n13450) );
  XNOR U17495 ( .A(n18116), .B(n15588), .Z(n13452) );
  XNOR U17496 ( .A(n18117), .B(n15254), .Z(n11635) );
  XNOR U17497 ( .A(n18118), .B(n18119), .Z(n15254) );
  AND U17498 ( .A(n13454), .B(n12747), .Z(n18117) );
  XOR U17499 ( .A(n18120), .B(n18121), .Z(n12747) );
  XNOR U17500 ( .A(n18122), .B(n17042), .Z(n13454) );
  XOR U17501 ( .A(n18123), .B(n18124), .Z(n15140) );
  XNOR U17502 ( .A(n12232), .B(n12576), .Z(n18124) );
  XOR U17503 ( .A(n18125), .B(n15273), .Z(n12576) );
  IV U17504 ( .A(n18126), .Z(n15273) );
  NOR U17505 ( .A(n16527), .B(n15441), .Z(n18125) );
  XNOR U17506 ( .A(n18127), .B(n15607), .Z(n15441) );
  XOR U17507 ( .A(n18128), .B(n15263), .Z(n12232) );
  ANDN U17508 ( .B(n16530), .A(n15443), .Z(n18128) );
  XNOR U17509 ( .A(n18129), .B(n18130), .Z(n15443) );
  IV U17510 ( .A(n18131), .Z(n16530) );
  XOR U17511 ( .A(n12250), .B(n18132), .Z(n18123) );
  XOR U17512 ( .A(n11895), .B(n11148), .Z(n18132) );
  XNOR U17513 ( .A(n18133), .B(n15281), .Z(n11148) );
  NOR U17514 ( .A(n16517), .B(n15438), .Z(n18133) );
  XOR U17515 ( .A(n18134), .B(n18135), .Z(n15438) );
  XOR U17516 ( .A(n18136), .B(n15267), .Z(n11895) );
  NOR U17517 ( .A(n18089), .B(n15445), .Z(n18136) );
  XNOR U17518 ( .A(n18137), .B(n17388), .Z(n15445) );
  ANDN U17519 ( .B(n16521), .A(n15436), .Z(n18138) );
  XNOR U17520 ( .A(n18139), .B(n18140), .Z(n15436) );
  XOR U17521 ( .A(n13012), .B(n11936), .Z(n9951) );
  XNOR U17522 ( .A(n12742), .B(n14710), .Z(n11936) );
  XNOR U17523 ( .A(n18141), .B(n18142), .Z(n14710) );
  XNOR U17524 ( .A(n11762), .B(n12454), .Z(n18142) );
  XOR U17525 ( .A(n18143), .B(n15233), .Z(n12454) );
  ANDN U17526 ( .B(n14165), .A(n14712), .Z(n18143) );
  XNOR U17527 ( .A(n18144), .B(n18145), .Z(n14712) );
  XNOR U17528 ( .A(n18146), .B(n17369), .Z(n14165) );
  XNOR U17529 ( .A(n18147), .B(n13490), .Z(n11762) );
  ANDN U17530 ( .B(n13536), .A(n13538), .Z(n18147) );
  XNOR U17531 ( .A(n17959), .B(n18148), .Z(n13538) );
  XOR U17532 ( .A(n18149), .B(n18140), .Z(n13536) );
  XNOR U17533 ( .A(n9772), .B(n18150), .Z(n18141) );
  XOR U17534 ( .A(n9662), .B(n12718), .Z(n18150) );
  XOR U17535 ( .A(n18151), .B(n13484), .Z(n12718) );
  NOR U17536 ( .A(n14050), .B(n13483), .Z(n18151) );
  XOR U17537 ( .A(n16954), .B(n18152), .Z(n13483) );
  XNOR U17538 ( .A(n15903), .B(n18153), .Z(n14050) );
  ANDN U17539 ( .B(n13544), .A(n13542), .Z(n18154) );
  XNOR U17540 ( .A(n18156), .B(n18157), .Z(n13544) );
  XNOR U17541 ( .A(n18158), .B(n13479), .Z(n9772) );
  NOR U17542 ( .A(n13546), .B(n13480), .Z(n18158) );
  XNOR U17543 ( .A(n18159), .B(n18160), .Z(n13480) );
  XNOR U17544 ( .A(n18161), .B(n18162), .Z(n13546) );
  XOR U17545 ( .A(n18163), .B(n18164), .Z(n12742) );
  XOR U17546 ( .A(n10541), .B(n11584), .Z(n18164) );
  XOR U17547 ( .A(n18165), .B(n13389), .Z(n11584) );
  IV U17548 ( .A(n13506), .Z(n13389) );
  XOR U17549 ( .A(n18166), .B(n18167), .Z(n13506) );
  AND U17550 ( .A(n13007), .B(n17129), .Z(n18165) );
  IV U17551 ( .A(n13008), .Z(n17129) );
  XOR U17552 ( .A(n18168), .B(n15257), .Z(n13008) );
  IV U17553 ( .A(n17809), .Z(n15257) );
  XOR U17554 ( .A(n17234), .B(n18169), .Z(n13007) );
  XNOR U17555 ( .A(n18170), .B(n13504), .Z(n10541) );
  XOR U17556 ( .A(n18171), .B(n18172), .Z(n13504) );
  XOR U17557 ( .A(n18173), .B(n17485), .Z(n13503) );
  XOR U17558 ( .A(n18174), .B(n18026), .Z(n14347) );
  IV U17559 ( .A(n16988), .Z(n18026) );
  XNOR U17560 ( .A(n18175), .B(n18176), .Z(n16988) );
  XOR U17561 ( .A(n13474), .B(n18177), .Z(n18163) );
  XOR U17562 ( .A(n11776), .B(n10171), .Z(n18177) );
  XOR U17563 ( .A(n18178), .B(n13028), .Z(n10171) );
  IV U17564 ( .A(n13498), .Z(n13028) );
  XNOR U17565 ( .A(n18179), .B(n18180), .Z(n13498) );
  NOR U17566 ( .A(n13014), .B(n13016), .Z(n18178) );
  XNOR U17567 ( .A(n18181), .B(n18182), .Z(n13016) );
  XNOR U17568 ( .A(n18183), .B(n17140), .Z(n13014) );
  XOR U17569 ( .A(n18184), .B(n13034), .Z(n11776) );
  IV U17570 ( .A(n13496), .Z(n13034) );
  XNOR U17571 ( .A(n18185), .B(n17218), .Z(n13496) );
  XOR U17572 ( .A(n18186), .B(n13037), .Z(n13474) );
  XNOR U17573 ( .A(n18187), .B(n15520), .Z(n13037) );
  IV U17574 ( .A(n18113), .Z(n15520) );
  NOR U17575 ( .A(n13003), .B(n13004), .Z(n18186) );
  XNOR U17576 ( .A(n18188), .B(n16458), .Z(n13004) );
  XNOR U17577 ( .A(n18189), .B(n17458), .Z(n13003) );
  XNOR U17578 ( .A(n18190), .B(n13495), .Z(n13012) );
  XNOR U17579 ( .A(n18191), .B(n18192), .Z(n13495) );
  ANDN U17580 ( .B(n17125), .A(n13033), .Z(n18190) );
  XNOR U17581 ( .A(n18193), .B(n18194), .Z(n13033) );
  XNOR U17582 ( .A(n18195), .B(n17167), .Z(n17125) );
  XNOR U17583 ( .A(n18196), .B(n6821), .Z(n3312) );
  XNOR U17584 ( .A(n17253), .B(n9112), .Z(n6821) );
  IV U17585 ( .A(n10439), .Z(n9112) );
  XOR U17586 ( .A(n18197), .B(n13199), .Z(n10439) );
  XOR U17587 ( .A(n18198), .B(n18199), .Z(n13199) );
  XNOR U17588 ( .A(n10469), .B(n10205), .Z(n18199) );
  XNOR U17589 ( .A(n18200), .B(n13739), .Z(n10205) );
  XOR U17590 ( .A(n18201), .B(n17730), .Z(n13739) );
  ANDN U17591 ( .B(n15844), .A(n15800), .Z(n18200) );
  XOR U17592 ( .A(n18202), .B(n13743), .Z(n10469) );
  XOR U17593 ( .A(n18203), .B(n16995), .Z(n13743) );
  XNOR U17594 ( .A(n18204), .B(n18205), .Z(n16995) );
  ANDN U17595 ( .B(n15847), .A(n15791), .Z(n18202) );
  XNOR U17596 ( .A(n15598), .B(n18207), .Z(n15847) );
  XOR U17597 ( .A(n10239), .B(n18208), .Z(n18198) );
  XNOR U17598 ( .A(n9566), .B(n10487), .Z(n18208) );
  XNOR U17599 ( .A(n18209), .B(n13735), .Z(n10487) );
  XNOR U17600 ( .A(n18210), .B(n15249), .Z(n13735) );
  ANDN U17601 ( .B(n15857), .A(n15796), .Z(n18209) );
  XNOR U17602 ( .A(n18211), .B(n17917), .Z(n15796) );
  XNOR U17603 ( .A(n17397), .B(n18212), .Z(n15857) );
  XNOR U17604 ( .A(n18213), .B(n13730), .Z(n9566) );
  IV U17605 ( .A(n15860), .Z(n13730) );
  XNOR U17606 ( .A(n18214), .B(n18215), .Z(n15860) );
  AND U17607 ( .A(n15793), .B(n15861), .Z(n18213) );
  XNOR U17608 ( .A(n18114), .B(n18216), .Z(n15861) );
  XOR U17609 ( .A(n18217), .B(n18218), .Z(n15793) );
  XOR U17610 ( .A(n18219), .B(n13726), .Z(n10239) );
  IV U17611 ( .A(n15853), .Z(n13726) );
  XOR U17612 ( .A(n18220), .B(n16938), .Z(n15853) );
  AND U17613 ( .A(n15798), .B(n17255), .Z(n18219) );
  XOR U17614 ( .A(n18221), .B(n18222), .Z(n17255) );
  XNOR U17615 ( .A(n16954), .B(n18223), .Z(n15798) );
  XNOR U17616 ( .A(n18224), .B(n15844), .Z(n17253) );
  XOR U17617 ( .A(n17993), .B(n18225), .Z(n15844) );
  AND U17618 ( .A(n15800), .B(n13737), .Z(n18224) );
  IV U17619 ( .A(n15801), .Z(n13737) );
  XOR U17620 ( .A(n18226), .B(n16055), .Z(n15801) );
  XNOR U17621 ( .A(n18193), .B(n18227), .Z(n15800) );
  AND U17622 ( .A(n6820), .B(n7592), .Z(n18196) );
  XNOR U17623 ( .A(n17690), .B(n11793), .Z(n7592) );
  XNOR U17624 ( .A(n18228), .B(n18229), .Z(n17690) );
  ANDN U17625 ( .B(n18230), .A(n18231), .Z(n18228) );
  XNOR U17626 ( .A(n13944), .B(n9602), .Z(n6820) );
  XNOR U17627 ( .A(n15011), .B(n14444), .Z(n9602) );
  XNOR U17628 ( .A(n18232), .B(n18233), .Z(n14444) );
  XNOR U17629 ( .A(n11186), .B(n14470), .Z(n18233) );
  XNOR U17630 ( .A(n18234), .B(n15398), .Z(n14470) );
  XOR U17631 ( .A(n18235), .B(n18236), .Z(n15398) );
  AND U17632 ( .A(n15399), .B(n14212), .Z(n18234) );
  IV U17633 ( .A(n18237), .Z(n14212) );
  XNOR U17634 ( .A(n18238), .B(n15404), .Z(n11186) );
  XNOR U17635 ( .A(n16898), .B(n18239), .Z(n15404) );
  AND U17636 ( .A(n14209), .B(n15405), .Z(n18238) );
  XOR U17637 ( .A(n17205), .B(n18240), .Z(n15405) );
  IV U17638 ( .A(n13957), .Z(n14209) );
  XOR U17639 ( .A(n18241), .B(n18242), .Z(n13957) );
  XOR U17640 ( .A(n12789), .B(n18243), .Z(n18232) );
  XOR U17641 ( .A(n10560), .B(n10683), .Z(n18243) );
  XOR U17642 ( .A(n18244), .B(n15541), .Z(n10683) );
  XNOR U17643 ( .A(n18245), .B(n18246), .Z(n15541) );
  AND U17644 ( .A(n13959), .B(n14206), .Z(n18244) );
  IV U17645 ( .A(n13961), .Z(n14206) );
  XNOR U17646 ( .A(n18247), .B(n13896), .Z(n13961) );
  XNOR U17647 ( .A(n18248), .B(n17546), .Z(n13959) );
  XOR U17648 ( .A(n18249), .B(n15402), .Z(n10560) );
  XNOR U17649 ( .A(n18250), .B(n15856), .Z(n15402) );
  ANDN U17650 ( .B(n13948), .A(n13946), .Z(n18249) );
  XOR U17651 ( .A(n18251), .B(n18252), .Z(n13946) );
  XNOR U17652 ( .A(n18253), .B(n18254), .Z(n13948) );
  XNOR U17653 ( .A(n18255), .B(n15407), .Z(n12789) );
  XNOR U17654 ( .A(n18256), .B(n16812), .Z(n15407) );
  AND U17655 ( .A(n13951), .B(n13953), .Z(n18255) );
  XOR U17656 ( .A(n18257), .B(n18258), .Z(n13953) );
  XNOR U17657 ( .A(n18259), .B(n17243), .Z(n13951) );
  XOR U17658 ( .A(n18260), .B(n18261), .Z(n15011) );
  XNOR U17659 ( .A(n9799), .B(n10689), .Z(n18261) );
  XOR U17660 ( .A(n18262), .B(n14491), .Z(n10689) );
  XNOR U17661 ( .A(n18263), .B(n15325), .Z(n14491) );
  ANDN U17662 ( .B(n16284), .A(n14490), .Z(n18262) );
  XNOR U17663 ( .A(n18264), .B(n15623), .Z(n14490) );
  IV U17664 ( .A(n15456), .Z(n16284) );
  XNOR U17665 ( .A(n16547), .B(n18265), .Z(n15456) );
  XNOR U17666 ( .A(n18266), .B(n14476), .Z(n9799) );
  XNOR U17667 ( .A(n18267), .B(n16749), .Z(n14476) );
  AND U17668 ( .A(n14477), .B(n16279), .Z(n18266) );
  IV U17669 ( .A(n15459), .Z(n16279) );
  XOR U17670 ( .A(n18268), .B(n17243), .Z(n15459) );
  XNOR U17671 ( .A(n18269), .B(n18270), .Z(n14477) );
  XOR U17672 ( .A(n13221), .B(n18271), .Z(n18260) );
  XNOR U17673 ( .A(n12591), .B(n11290), .Z(n18271) );
  XNOR U17674 ( .A(n18272), .B(n14487), .Z(n11290) );
  AND U17675 ( .A(n14486), .B(n16274), .Z(n18272) );
  IV U17676 ( .A(n15466), .Z(n16274) );
  XOR U17677 ( .A(n18274), .B(n18242), .Z(n15466) );
  XOR U17678 ( .A(n18275), .B(n17948), .Z(n14486) );
  XNOR U17679 ( .A(n18276), .B(n17548), .Z(n12591) );
  XNOR U17680 ( .A(n18277), .B(n17595), .Z(n17548) );
  AND U17681 ( .A(n15468), .B(n16281), .Z(n18276) );
  IV U17682 ( .A(n15470), .Z(n16281) );
  XOR U17683 ( .A(n18278), .B(n18279), .Z(n15470) );
  XOR U17684 ( .A(n18280), .B(n17928), .Z(n15468) );
  XNOR U17685 ( .A(n18281), .B(n14480), .Z(n13221) );
  XNOR U17686 ( .A(n18282), .B(n17123), .Z(n14480) );
  XNOR U17687 ( .A(n18283), .B(n13896), .Z(n14481) );
  IV U17688 ( .A(n15463), .Z(n16276) );
  XOR U17689 ( .A(n18286), .B(n14924), .Z(n15463) );
  XNOR U17690 ( .A(n18287), .B(n15399), .Z(n13944) );
  XNOR U17691 ( .A(n18288), .B(n16331), .Z(n15399) );
  ANDN U17692 ( .B(n18237), .A(n14213), .Z(n18287) );
  XOR U17693 ( .A(n16950), .B(n18289), .Z(n14213) );
  XOR U17694 ( .A(n18291), .B(n18292), .Z(n5931) );
  XNOR U17695 ( .A(n1842), .B(n5178), .Z(n18292) );
  XOR U17696 ( .A(n18293), .B(n7697), .Z(n5178) );
  XNOR U17697 ( .A(n17647), .B(n11173), .Z(n7697) );
  IV U17698 ( .A(n12385), .Z(n11173) );
  XOR U17699 ( .A(n14934), .B(n12927), .Z(n12385) );
  XNOR U17700 ( .A(n18294), .B(n18295), .Z(n12927) );
  XOR U17701 ( .A(n11904), .B(n11504), .Z(n18295) );
  XOR U17702 ( .A(n18296), .B(n15682), .Z(n11504) );
  AND U17703 ( .A(n17652), .B(n17653), .Z(n18296) );
  XOR U17704 ( .A(n15329), .B(n18297), .Z(n17653) );
  XOR U17705 ( .A(n18298), .B(n15674), .Z(n11904) );
  AND U17706 ( .A(n17650), .B(n18299), .Z(n18298) );
  XOR U17707 ( .A(n18300), .B(n17933), .Z(n17650) );
  XOR U17708 ( .A(n10715), .B(n18301), .Z(n18294) );
  XNOR U17709 ( .A(n11928), .B(n11546), .Z(n18301) );
  XNOR U17710 ( .A(n18302), .B(n15665), .Z(n11546) );
  ANDN U17711 ( .B(n18303), .A(n18037), .Z(n18302) );
  XNOR U17712 ( .A(n18304), .B(n15678), .Z(n11928) );
  ANDN U17713 ( .B(n17641), .A(n17642), .Z(n18304) );
  XNOR U17714 ( .A(n18305), .B(n18306), .Z(n17642) );
  XOR U17715 ( .A(n18307), .B(n15668), .Z(n10715) );
  AND U17716 ( .A(n17644), .B(n17645), .Z(n18307) );
  XOR U17717 ( .A(n18308), .B(n17835), .Z(n17645) );
  XOR U17718 ( .A(n18309), .B(n18310), .Z(n14934) );
  XNOR U17719 ( .A(n9169), .B(n13877), .Z(n18310) );
  XNOR U17720 ( .A(n18312), .B(n17360), .Z(n13343) );
  AND U17721 ( .A(n13893), .B(n15328), .Z(n18311) );
  XOR U17722 ( .A(n18313), .B(n17895), .Z(n15328) );
  XNOR U17723 ( .A(n18314), .B(n15516), .Z(n13893) );
  XNOR U17724 ( .A(n18315), .B(n13356), .Z(n9169) );
  XOR U17725 ( .A(n17220), .B(n18316), .Z(n13356) );
  NOR U17726 ( .A(n13875), .B(n13888), .Z(n18315) );
  XNOR U17727 ( .A(n15906), .B(n18317), .Z(n13888) );
  XOR U17728 ( .A(n18046), .B(n18318), .Z(n13875) );
  XNOR U17729 ( .A(n10243), .B(n18319), .Z(n18309) );
  XOR U17730 ( .A(n9560), .B(n10213), .Z(n18319) );
  XNOR U17731 ( .A(n18320), .B(n13339), .Z(n10213) );
  XNOR U17732 ( .A(n18321), .B(n16001), .Z(n13339) );
  AND U17733 ( .A(n13989), .B(n13899), .Z(n18320) );
  XNOR U17734 ( .A(n18322), .B(n18323), .Z(n13899) );
  XOR U17735 ( .A(n18324), .B(n16011), .Z(n13989) );
  XOR U17736 ( .A(n18325), .B(n13348), .Z(n9560) );
  XOR U17737 ( .A(n18326), .B(n14924), .Z(n13348) );
  ANDN U17738 ( .B(n15320), .A(n13871), .Z(n18325) );
  XOR U17739 ( .A(n18327), .B(n17489), .Z(n13871) );
  XNOR U17740 ( .A(n18328), .B(n14948), .Z(n15320) );
  XOR U17741 ( .A(n18331), .B(n13352), .Z(n10243) );
  XNOR U17742 ( .A(n18332), .B(n17144), .Z(n13352) );
  ANDN U17743 ( .B(n13884), .A(n13873), .Z(n18331) );
  XNOR U17744 ( .A(n18333), .B(n18334), .Z(n13873) );
  XNOR U17745 ( .A(n18335), .B(n16519), .Z(n13884) );
  XNOR U17746 ( .A(n18336), .B(n18303), .Z(n17647) );
  ANDN U17747 ( .B(n18037), .A(n15663), .Z(n18336) );
  XNOR U17748 ( .A(n18337), .B(n15333), .Z(n15663) );
  XNOR U17749 ( .A(n18338), .B(n18339), .Z(n18037) );
  AND U17750 ( .A(n6853), .B(n7577), .Z(n18293) );
  XOR U17751 ( .A(n18340), .B(n10139), .Z(n7577) );
  XNOR U17752 ( .A(n18341), .B(n16130), .Z(n10139) );
  XNOR U17753 ( .A(n18342), .B(n18343), .Z(n16130) );
  XNOR U17754 ( .A(n12940), .B(n11882), .Z(n18343) );
  XNOR U17755 ( .A(n18344), .B(n16359), .Z(n11882) );
  XOR U17756 ( .A(n18345), .B(n16677), .Z(n16359) );
  IV U17757 ( .A(n17595), .Z(n16677) );
  ANDN U17758 ( .B(n15550), .A(n16363), .Z(n18344) );
  XNOR U17759 ( .A(n18346), .B(n14775), .Z(n12940) );
  XOR U17760 ( .A(n18347), .B(n18348), .Z(n14775) );
  AND U17761 ( .A(n15565), .B(n14776), .Z(n18346) );
  XNOR U17762 ( .A(n12909), .B(n18349), .Z(n18342) );
  XOR U17763 ( .A(n9384), .B(n9531), .Z(n18349) );
  XOR U17764 ( .A(n18350), .B(n15810), .Z(n9531) );
  XOR U17765 ( .A(n18351), .B(n18352), .Z(n15810) );
  AND U17766 ( .A(n15554), .B(n15811), .Z(n18350) );
  XNOR U17767 ( .A(n18353), .B(n14769), .Z(n9384) );
  XNOR U17768 ( .A(n18354), .B(n18355), .Z(n14769) );
  NOR U17769 ( .A(n14768), .B(n15562), .Z(n18353) );
  XOR U17770 ( .A(n18356), .B(n14764), .Z(n12909) );
  XNOR U17771 ( .A(n18357), .B(n17483), .Z(n14764) );
  ANDN U17772 ( .B(n14765), .A(n15559), .Z(n18356) );
  XNOR U17773 ( .A(n11691), .B(n13229), .Z(n6853) );
  XNOR U17774 ( .A(n18358), .B(n16789), .Z(n13229) );
  ANDN U17775 ( .B(n13750), .A(n13751), .Z(n18358) );
  XNOR U17776 ( .A(n18359), .B(n16261), .Z(n13751) );
  XOR U17777 ( .A(n13589), .B(n12766), .Z(n11691) );
  XNOR U17778 ( .A(n18360), .B(n18361), .Z(n12766) );
  XNOR U17779 ( .A(n11813), .B(n9269), .Z(n18361) );
  XNOR U17780 ( .A(n18362), .B(n13786), .Z(n9269) );
  XNOR U17781 ( .A(n18363), .B(n17075), .Z(n13786) );
  ANDN U17782 ( .B(n15174), .A(n13785), .Z(n18362) );
  XOR U17783 ( .A(n14914), .B(n18364), .Z(n13785) );
  XOR U17784 ( .A(n18365), .B(n18366), .Z(n11813) );
  ANDN U17785 ( .B(n15180), .A(n13771), .Z(n18365) );
  XOR U17786 ( .A(n18367), .B(n18368), .Z(n13771) );
  XOR U17787 ( .A(n10199), .B(n18369), .Z(n18360) );
  XOR U17788 ( .A(n11158), .B(n13766), .Z(n18369) );
  XNOR U17789 ( .A(n18370), .B(n13775), .Z(n13766) );
  XNOR U17790 ( .A(n18371), .B(n13883), .Z(n13775) );
  AND U17791 ( .A(n13776), .B(n15177), .Z(n18370) );
  XNOR U17792 ( .A(n18372), .B(n17469), .Z(n13776) );
  XNOR U17793 ( .A(n18373), .B(n13781), .Z(n11158) );
  XNOR U17794 ( .A(n18374), .B(n17786), .Z(n13781) );
  ANDN U17795 ( .B(n13782), .A(n15165), .Z(n18373) );
  XOR U17796 ( .A(n18375), .B(n18376), .Z(n13782) );
  XNOR U17797 ( .A(n18377), .B(n15704), .Z(n10199) );
  XNOR U17798 ( .A(n18378), .B(n18379), .Z(n15704) );
  NOR U17799 ( .A(n15168), .B(n15169), .Z(n18377) );
  XOR U17800 ( .A(n16543), .B(n18380), .Z(n15168) );
  XOR U17801 ( .A(n18381), .B(n18382), .Z(n13589) );
  XOR U17802 ( .A(n10288), .B(n9937), .Z(n18382) );
  XOR U17803 ( .A(n18383), .B(n15963), .Z(n9937) );
  XNOR U17804 ( .A(n18384), .B(n17474), .Z(n15963) );
  ANDN U17805 ( .B(n16789), .A(n13750), .Z(n18383) );
  XNOR U17806 ( .A(n18385), .B(n17732), .Z(n13750) );
  XOR U17807 ( .A(n15647), .B(n18386), .Z(n16789) );
  XOR U17808 ( .A(n18387), .B(n15960), .Z(n10288) );
  IV U17809 ( .A(n16780), .Z(n15960) );
  XNOR U17810 ( .A(n18388), .B(n18389), .Z(n16780) );
  NOR U17811 ( .A(n14851), .B(n13761), .Z(n18387) );
  XNOR U17812 ( .A(n18390), .B(n15222), .Z(n13761) );
  XOR U17813 ( .A(n18391), .B(n18392), .Z(n15222) );
  XOR U17814 ( .A(n18393), .B(n18394), .Z(n14851) );
  XOR U17815 ( .A(n11657), .B(n18395), .Z(n18381) );
  XOR U17816 ( .A(n10807), .B(n11646), .Z(n18395) );
  XNOR U17817 ( .A(n18396), .B(n15969), .Z(n11646) );
  XNOR U17818 ( .A(n18397), .B(n18368), .Z(n15969) );
  ANDN U17819 ( .B(n13241), .A(n13242), .Z(n18396) );
  XOR U17820 ( .A(n18398), .B(n18399), .Z(n13242) );
  XNOR U17821 ( .A(n18400), .B(n17270), .Z(n13241) );
  XNOR U17822 ( .A(n18401), .B(n15966), .Z(n10807) );
  XNOR U17823 ( .A(n18402), .B(n17879), .Z(n15966) );
  ANDN U17824 ( .B(n13231), .A(n13232), .Z(n18401) );
  XNOR U17825 ( .A(n18403), .B(n18404), .Z(n13232) );
  IV U17826 ( .A(n16785), .Z(n13231) );
  XOR U17827 ( .A(n18405), .B(n18406), .Z(n16785) );
  XNOR U17828 ( .A(n18407), .B(n15956), .Z(n11657) );
  XNOR U17829 ( .A(n17223), .B(n18408), .Z(n15956) );
  AND U17830 ( .A(n13237), .B(n13754), .Z(n18407) );
  IV U17831 ( .A(n13239), .Z(n13754) );
  XNOR U17832 ( .A(n18409), .B(n18022), .Z(n13239) );
  XOR U17833 ( .A(n18410), .B(n18379), .Z(n13237) );
  XOR U17834 ( .A(n18411), .B(n7691), .Z(n1842) );
  XOR U17835 ( .A(n11247), .B(n16483), .Z(n7691) );
  XNOR U17836 ( .A(n18412), .B(n14733), .Z(n16483) );
  ANDN U17837 ( .B(n17709), .A(n18413), .Z(n18412) );
  XOR U17838 ( .A(n18003), .B(n18414), .Z(n11247) );
  XOR U17839 ( .A(n18415), .B(n18416), .Z(n18003) );
  XNOR U17840 ( .A(n11033), .B(n11942), .Z(n18416) );
  XOR U17841 ( .A(n18417), .B(n14956), .Z(n11942) );
  XOR U17842 ( .A(n18418), .B(n17360), .Z(n14956) );
  ANDN U17843 ( .B(n14957), .A(n17265), .Z(n18417) );
  XNOR U17844 ( .A(n18419), .B(n17167), .Z(n17265) );
  XNOR U17845 ( .A(n18034), .B(n18420), .Z(n14957) );
  XNOR U17846 ( .A(n18421), .B(n16289), .Z(n11033) );
  XNOR U17847 ( .A(n18422), .B(n18423), .Z(n16289) );
  ANDN U17848 ( .B(n16290), .A(n16820), .Z(n18421) );
  XOR U17849 ( .A(n18424), .B(n18425), .Z(n16820) );
  XNOR U17850 ( .A(n18426), .B(n16027), .Z(n16290) );
  XOR U17851 ( .A(n11794), .B(n18427), .Z(n18415) );
  XOR U17852 ( .A(n9084), .B(n10795), .Z(n18427) );
  XOR U17853 ( .A(n18428), .B(n14747), .Z(n10795) );
  XNOR U17854 ( .A(n18429), .B(n16746), .Z(n14747) );
  XNOR U17855 ( .A(n18430), .B(n15984), .Z(n14746) );
  XOR U17856 ( .A(n18431), .B(n17908), .Z(n16810) );
  XOR U17857 ( .A(n18432), .B(n14753), .Z(n9084) );
  XNOR U17858 ( .A(n18433), .B(n18434), .Z(n14753) );
  ANDN U17859 ( .B(n14754), .A(n16806), .Z(n18432) );
  XOR U17860 ( .A(n14914), .B(n18435), .Z(n16806) );
  XNOR U17861 ( .A(n18436), .B(n18121), .Z(n14754) );
  XNOR U17862 ( .A(n18437), .B(n14742), .Z(n11794) );
  XNOR U17863 ( .A(n18438), .B(n18439), .Z(n14742) );
  AND U17864 ( .A(n16816), .B(n14743), .Z(n18437) );
  XNOR U17865 ( .A(n18440), .B(n16999), .Z(n14743) );
  IV U17866 ( .A(n18394), .Z(n16999) );
  XNOR U17867 ( .A(n18441), .B(n18102), .Z(n16816) );
  ANDN U17868 ( .B(n7692), .A(n6846), .Z(n18411) );
  XOR U17869 ( .A(n18442), .B(n9183), .Z(n6846) );
  XOR U17870 ( .A(n18443), .B(n16596), .Z(n9183) );
  XOR U17871 ( .A(n18444), .B(n18445), .Z(n16596) );
  XOR U17872 ( .A(n13835), .B(n10600), .Z(n18445) );
  XNOR U17873 ( .A(n18446), .B(n18447), .Z(n10600) );
  AND U17874 ( .A(n17760), .B(n17762), .Z(n18446) );
  XNOR U17875 ( .A(n18448), .B(n16924), .Z(n17762) );
  XNOR U17876 ( .A(n18449), .B(n14194), .Z(n13835) );
  AND U17877 ( .A(n17766), .B(n17764), .Z(n18449) );
  XNOR U17878 ( .A(n18450), .B(n17800), .Z(n17764) );
  XNOR U17879 ( .A(n15132), .B(n18451), .Z(n17766) );
  XOR U17880 ( .A(n18452), .B(n18453), .Z(n15132) );
  XNOR U17881 ( .A(n10484), .B(n18454), .Z(n18444) );
  XOR U17882 ( .A(n9992), .B(n9683), .Z(n18454) );
  XOR U17883 ( .A(n18455), .B(n15051), .Z(n9683) );
  ANDN U17884 ( .B(n17769), .A(n15052), .Z(n18455) );
  XOR U17885 ( .A(n18456), .B(n16698), .Z(n15052) );
  XOR U17886 ( .A(n18457), .B(n18458), .Z(n17769) );
  XNOR U17887 ( .A(n18459), .B(n18460), .Z(n9992) );
  AND U17888 ( .A(n17755), .B(n17757), .Z(n18459) );
  XOR U17889 ( .A(n18461), .B(n18462), .Z(n17757) );
  XOR U17890 ( .A(n18463), .B(n13842), .Z(n10484) );
  ANDN U17891 ( .B(n17827), .A(n13843), .Z(n18463) );
  XOR U17892 ( .A(n18464), .B(n18465), .Z(n13843) );
  IV U17893 ( .A(n17753), .Z(n17827) );
  XOR U17894 ( .A(n18466), .B(n16682), .Z(n17753) );
  XNOR U17895 ( .A(n15994), .B(n12176), .Z(n7692) );
  XNOR U17896 ( .A(n18467), .B(n17655), .Z(n12176) );
  XNOR U17897 ( .A(n18468), .B(n18469), .Z(n17655) );
  XNOR U17898 ( .A(n12595), .B(n12276), .Z(n18469) );
  XOR U17899 ( .A(n18470), .B(n17606), .Z(n12276) );
  XNOR U17900 ( .A(n18471), .B(n16749), .Z(n17606) );
  AND U17901 ( .A(n12399), .B(n12401), .Z(n18470) );
  XNOR U17902 ( .A(n18472), .B(n18473), .Z(n12401) );
  XNOR U17903 ( .A(n17887), .B(n18474), .Z(n12399) );
  XNOR U17904 ( .A(n18475), .B(n16089), .Z(n12595) );
  XOR U17905 ( .A(n18476), .B(n17634), .Z(n16089) );
  ANDN U17906 ( .B(n17608), .A(n13655), .Z(n18475) );
  XOR U17907 ( .A(n18477), .B(n17439), .Z(n13655) );
  XOR U17908 ( .A(n18478), .B(n16362), .Z(n17608) );
  XOR U17909 ( .A(n11187), .B(n18479), .Z(n18468) );
  XOR U17910 ( .A(n12620), .B(n12329), .Z(n18479) );
  XNOR U17911 ( .A(n18480), .B(n16077), .Z(n12329) );
  XNOR U17912 ( .A(n18481), .B(n16478), .Z(n16077) );
  AND U17913 ( .A(n17612), .B(n17657), .Z(n18480) );
  XOR U17914 ( .A(n16543), .B(n18482), .Z(n17657) );
  XNOR U17915 ( .A(n18483), .B(n18379), .Z(n17612) );
  XNOR U17916 ( .A(n18484), .B(n16085), .Z(n12620) );
  XNOR U17917 ( .A(n18485), .B(n18486), .Z(n16085) );
  ANDN U17918 ( .B(n14400), .A(n14401), .Z(n18484) );
  XOR U17919 ( .A(n18487), .B(n16340), .Z(n14401) );
  XNOR U17920 ( .A(n18488), .B(n18489), .Z(n14400) );
  XNOR U17921 ( .A(n18490), .B(n16081), .Z(n11187) );
  XOR U17922 ( .A(n18491), .B(n18022), .Z(n16081) );
  AND U17923 ( .A(n12411), .B(n17616), .Z(n18490) );
  XNOR U17924 ( .A(n18492), .B(n16011), .Z(n17616) );
  XNOR U17925 ( .A(n18493), .B(n18494), .Z(n12411) );
  XNOR U17926 ( .A(n18495), .B(n17629), .Z(n15994) );
  AND U17927 ( .A(n14510), .B(n14508), .Z(n18495) );
  IV U17928 ( .A(n18496), .Z(n14508) );
  XOR U17929 ( .A(n17402), .B(n18497), .Z(n14510) );
  XNOR U17930 ( .A(n4092), .B(n18498), .Z(n18291) );
  XOR U17931 ( .A(n7671), .B(n3586), .Z(n18498) );
  XNOR U17932 ( .A(n18499), .B(n10033), .Z(n3586) );
  XNOR U17933 ( .A(n13487), .B(n10712), .Z(n10033) );
  XOR U17934 ( .A(n13023), .B(n18500), .Z(n10712) );
  XOR U17935 ( .A(n18501), .B(n18502), .Z(n13023) );
  XNOR U17936 ( .A(n11807), .B(n11909), .Z(n18502) );
  XNOR U17937 ( .A(n18503), .B(n14051), .Z(n11909) );
  XNOR U17938 ( .A(n18504), .B(n13883), .Z(n14051) );
  IV U17939 ( .A(n18505), .Z(n13883) );
  ANDN U17940 ( .B(n13484), .A(n13482), .Z(n18503) );
  XOR U17941 ( .A(n18506), .B(n16938), .Z(n13482) );
  XOR U17942 ( .A(n18507), .B(n17121), .Z(n13484) );
  XOR U17943 ( .A(n18508), .B(n14167), .Z(n11807) );
  XOR U17944 ( .A(n18509), .B(n18510), .Z(n14167) );
  AND U17945 ( .A(n15233), .B(n14166), .Z(n18508) );
  XOR U17946 ( .A(n17205), .B(n18511), .Z(n14166) );
  XNOR U17947 ( .A(n18512), .B(n17218), .Z(n15233) );
  XOR U17948 ( .A(n14159), .B(n18513), .Z(n18501) );
  XOR U17949 ( .A(n11400), .B(n10306), .Z(n18513) );
  XOR U17950 ( .A(n18514), .B(n13537), .Z(n10306) );
  XOR U17951 ( .A(n18515), .B(n17483), .Z(n13537) );
  NOR U17952 ( .A(n13489), .B(n13490), .Z(n18514) );
  XNOR U17953 ( .A(n15626), .B(n18516), .Z(n13490) );
  XNOR U17954 ( .A(n18517), .B(n18172), .Z(n13489) );
  XOR U17955 ( .A(n18518), .B(n13543), .Z(n11400) );
  XOR U17956 ( .A(n18519), .B(n15843), .Z(n13543) );
  NOR U17957 ( .A(n18155), .B(n14163), .Z(n18518) );
  XOR U17958 ( .A(n18520), .B(n13547), .Z(n14159) );
  IV U17959 ( .A(n14172), .Z(n13547) );
  XOR U17960 ( .A(n18521), .B(n17485), .Z(n14172) );
  ANDN U17961 ( .B(n13478), .A(n13479), .Z(n18520) );
  XNOR U17962 ( .A(n15911), .B(n18522), .Z(n13479) );
  XOR U17963 ( .A(n18523), .B(n17925), .Z(n13478) );
  XOR U17964 ( .A(n18524), .B(n14163), .Z(n13487) );
  XNOR U17965 ( .A(n18525), .B(n15208), .Z(n14163) );
  AND U17966 ( .A(n13542), .B(n18155), .Z(n18524) );
  XOR U17967 ( .A(n18015), .B(n18526), .Z(n18155) );
  XOR U17968 ( .A(n18527), .B(n18528), .Z(n13542) );
  ANDN U17969 ( .B(n10066), .A(n6842), .Z(n18499) );
  XOR U17970 ( .A(n13817), .B(n9278), .Z(n6842) );
  IV U17971 ( .A(n13040), .Z(n9278) );
  XOR U17972 ( .A(n14124), .B(n14136), .Z(n13040) );
  XNOR U17973 ( .A(n18529), .B(n18530), .Z(n14136) );
  XNOR U17974 ( .A(n12140), .B(n13394), .Z(n18530) );
  XNOR U17975 ( .A(n18531), .B(n14871), .Z(n13394) );
  NOR U17976 ( .A(n14872), .B(n15781), .Z(n18531) );
  XNOR U17977 ( .A(n18532), .B(n17451), .Z(n15781) );
  XNOR U17978 ( .A(n18533), .B(n18534), .Z(n17451) );
  XNOR U17979 ( .A(n18535), .B(n18399), .Z(n14872) );
  XNOR U17980 ( .A(n18536), .B(n14865), .Z(n12140) );
  ANDN U17981 ( .B(n14866), .A(n15784), .Z(n18536) );
  XOR U17982 ( .A(n18537), .B(n18473), .Z(n15784) );
  XOR U17983 ( .A(n18538), .B(n16003), .Z(n14866) );
  XOR U17984 ( .A(n11042), .B(n18539), .Z(n18529) );
  XOR U17985 ( .A(n10822), .B(n11683), .Z(n18539) );
  XNOR U17986 ( .A(n18540), .B(n14861), .Z(n11683) );
  XOR U17987 ( .A(n18217), .B(n18541), .Z(n14862) );
  XOR U17988 ( .A(n18542), .B(n17876), .Z(n15776) );
  XOR U17989 ( .A(n18543), .B(n14876), .Z(n10822) );
  NOR U17990 ( .A(n14875), .B(n16736), .Z(n18543) );
  XNOR U17991 ( .A(n18544), .B(n16100), .Z(n16736) );
  XOR U17992 ( .A(n18545), .B(n18546), .Z(n14875) );
  XNOR U17993 ( .A(n18547), .B(n18548), .Z(n11042) );
  NOR U17994 ( .A(n15772), .B(n16729), .Z(n18547) );
  XOR U17995 ( .A(n18549), .B(n18550), .Z(n15772) );
  XOR U17996 ( .A(n18551), .B(n18552), .Z(n14124) );
  XNOR U17997 ( .A(n9698), .B(n12739), .Z(n18552) );
  XOR U17998 ( .A(n18553), .B(n14693), .Z(n12739) );
  XNOR U17999 ( .A(n18554), .B(n15824), .Z(n14693) );
  NOR U18000 ( .A(n13834), .B(n13832), .Z(n18553) );
  XOR U18001 ( .A(n18555), .B(n17546), .Z(n13832) );
  XNOR U18002 ( .A(n18556), .B(n14703), .Z(n9698) );
  XNOR U18003 ( .A(n18557), .B(n18172), .Z(n14703) );
  AND U18004 ( .A(n18558), .B(n15692), .Z(n18556) );
  XNOR U18005 ( .A(n14855), .B(n18559), .Z(n18551) );
  XNOR U18006 ( .A(n9719), .B(n12571), .Z(n18559) );
  XOR U18007 ( .A(n18560), .B(n14697), .Z(n12571) );
  IV U18008 ( .A(n15699), .Z(n14697) );
  XOR U18009 ( .A(n15906), .B(n18561), .Z(n15699) );
  IV U18010 ( .A(n17064), .Z(n15906) );
  XOR U18011 ( .A(n18562), .B(n18563), .Z(n17064) );
  ANDN U18012 ( .B(n18564), .A(n13828), .Z(n18560) );
  XNOR U18013 ( .A(n18565), .B(n18566), .Z(n13828) );
  XNOR U18014 ( .A(n18567), .B(n14690), .Z(n9719) );
  IV U18015 ( .A(n15695), .Z(n14690) );
  XOR U18016 ( .A(n18568), .B(n15623), .Z(n15695) );
  XOR U18017 ( .A(n18569), .B(n14941), .Z(n13824) );
  IV U18018 ( .A(n16934), .Z(n14941) );
  XNOR U18019 ( .A(n18570), .B(n14699), .Z(n14855) );
  XOR U18020 ( .A(n18571), .B(n17564), .Z(n14699) );
  NOR U18021 ( .A(n13821), .B(n13819), .Z(n18570) );
  XOR U18022 ( .A(n18572), .B(n18464), .Z(n13819) );
  XOR U18023 ( .A(n18573), .B(n15692), .Z(n13817) );
  XNOR U18024 ( .A(n18574), .B(n16795), .Z(n15692) );
  ANDN U18025 ( .B(n18575), .A(n14702), .Z(n18573) );
  XNOR U18026 ( .A(n13846), .B(n10050), .Z(n10066) );
  XOR U18027 ( .A(n18576), .B(n17829), .Z(n13846) );
  ANDN U18028 ( .B(n18447), .A(n17760), .Z(n18576) );
  XNOR U18029 ( .A(n18577), .B(n17123), .Z(n17760) );
  IV U18030 ( .A(n18578), .Z(n17123) );
  XOR U18031 ( .A(n18579), .B(n7689), .Z(n7671) );
  IV U18032 ( .A(n10023), .Z(n7689) );
  XNOR U18033 ( .A(n16431), .B(n9687), .Z(n10023) );
  XOR U18034 ( .A(n18580), .B(n15502), .Z(n16431) );
  NOR U18035 ( .A(n18581), .B(n18582), .Z(n18580) );
  NOR U18036 ( .A(n7586), .B(n6831), .Z(n18579) );
  XNOR U18037 ( .A(n14139), .B(n9768), .Z(n6831) );
  XOR U18038 ( .A(n18583), .B(n18584), .Z(n17748) );
  XNOR U18039 ( .A(n18442), .B(n14216), .Z(n18584) );
  XNOR U18040 ( .A(n18585), .B(n16843), .Z(n14216) );
  NOR U18041 ( .A(n14639), .B(n14638), .Z(n18585) );
  XOR U18042 ( .A(n18586), .B(n17945), .Z(n14639) );
  XNOR U18043 ( .A(n18587), .B(n14067), .Z(n18442) );
  ANDN U18044 ( .B(n17152), .A(n16835), .Z(n18587) );
  XNOR U18045 ( .A(n18588), .B(n18589), .Z(n16835) );
  XOR U18046 ( .A(n9182), .B(n18590), .Z(n18583) );
  XNOR U18047 ( .A(n9949), .B(n13507), .Z(n18590) );
  XOR U18048 ( .A(n18591), .B(n14063), .Z(n13507) );
  IV U18049 ( .A(n18592), .Z(n14063) );
  NOR U18050 ( .A(n14636), .B(n14635), .Z(n18591) );
  XNOR U18051 ( .A(n18593), .B(n18594), .Z(n14636) );
  XNOR U18052 ( .A(n18595), .B(n14076), .Z(n9949) );
  IV U18053 ( .A(n18596), .Z(n14076) );
  ANDN U18054 ( .B(n16837), .A(n17771), .Z(n18595) );
  XOR U18055 ( .A(n18597), .B(n17197), .Z(n16837) );
  XNOR U18056 ( .A(n18598), .B(n18599), .Z(n17197) );
  XNOR U18057 ( .A(n18600), .B(n14071), .Z(n9182) );
  XOR U18058 ( .A(n18601), .B(n18602), .Z(n15074) );
  XNOR U18059 ( .A(n18603), .B(n18604), .Z(n13395) );
  XNOR U18060 ( .A(n14713), .B(n18605), .Z(n18604) );
  XOR U18061 ( .A(n18606), .B(n15764), .Z(n14713) );
  ANDN U18062 ( .B(n18607), .A(n14142), .Z(n18606) );
  XOR U18063 ( .A(n18608), .B(n18609), .Z(n14142) );
  XNOR U18064 ( .A(n12147), .B(n18610), .Z(n18603) );
  XOR U18065 ( .A(n10214), .B(n13314), .Z(n18610) );
  XOR U18066 ( .A(n18611), .B(n15768), .Z(n13314) );
  ANDN U18067 ( .B(n18612), .A(n14148), .Z(n18611) );
  XOR U18068 ( .A(n18613), .B(n18399), .Z(n14148) );
  XOR U18069 ( .A(n18614), .B(n15758), .Z(n10214) );
  ANDN U18070 ( .B(n14153), .A(n14151), .Z(n18614) );
  XNOR U18071 ( .A(n18615), .B(n18616), .Z(n14153) );
  XNOR U18072 ( .A(n18617), .B(n15755), .Z(n12147) );
  AND U18073 ( .A(n16742), .B(n18618), .Z(n18617) );
  XOR U18074 ( .A(n18619), .B(n18620), .Z(n14139) );
  XOR U18075 ( .A(n18621), .B(n18622), .Z(n18620) );
  OR U18076 ( .A(n15753), .B(n16742), .Z(n18622) );
  AND U18077 ( .A(n6835), .B(n15691), .Z(n18621) );
  XOR U18078 ( .A(n9480), .B(n18626), .Z(n7586) );
  IV U18079 ( .A(n12285), .Z(n9480) );
  XOR U18080 ( .A(n12212), .B(n11929), .Z(n12285) );
  XOR U18081 ( .A(n18627), .B(n18628), .Z(n11929) );
  XNOR U18082 ( .A(n12080), .B(n13332), .Z(n18628) );
  XOR U18083 ( .A(n18629), .B(n18040), .Z(n13332) );
  IV U18084 ( .A(n15681), .Z(n18040) );
  XNOR U18085 ( .A(n18630), .B(n15529), .Z(n15681) );
  XNOR U18086 ( .A(n18631), .B(n18632), .Z(n15529) );
  ANDN U18087 ( .B(n15682), .A(n17652), .Z(n18629) );
  XOR U18088 ( .A(n18633), .B(n17369), .Z(n17652) );
  XNOR U18089 ( .A(n18634), .B(n18389), .Z(n15682) );
  XNOR U18090 ( .A(n18635), .B(n15673), .Z(n12080) );
  XNOR U18091 ( .A(n18636), .B(n17678), .Z(n15673) );
  XOR U18092 ( .A(n18637), .B(n18638), .Z(n15674) );
  IV U18093 ( .A(n18299), .Z(n17649) );
  XOR U18094 ( .A(n18639), .B(n16456), .Z(n18299) );
  XOR U18095 ( .A(n11557), .B(n18640), .Z(n18627) );
  XOR U18096 ( .A(n9696), .B(n12312), .Z(n18640) );
  XNOR U18097 ( .A(n18641), .B(n15664), .Z(n12312) );
  XOR U18098 ( .A(n18642), .B(n18643), .Z(n15664) );
  XOR U18099 ( .A(n16950), .B(n18644), .Z(n18303) );
  IV U18100 ( .A(n17939), .Z(n16950) );
  XOR U18101 ( .A(n18645), .B(n18008), .Z(n15665) );
  XOR U18102 ( .A(n18646), .B(n15677), .Z(n9696) );
  XNOR U18103 ( .A(n18647), .B(n18648), .Z(n15677) );
  ANDN U18104 ( .B(n15678), .A(n17641), .Z(n18646) );
  XNOR U18105 ( .A(n18403), .B(n18649), .Z(n17641) );
  XOR U18106 ( .A(n18650), .B(n18651), .Z(n15678) );
  XOR U18107 ( .A(n17332), .B(n18653), .Z(n15669) );
  NOR U18108 ( .A(n17644), .B(n15668), .Z(n18652) );
  XNOR U18109 ( .A(n18654), .B(n16952), .Z(n15668) );
  IV U18110 ( .A(n18258), .Z(n16952) );
  XNOR U18111 ( .A(n18655), .B(n17439), .Z(n17644) );
  XOR U18112 ( .A(n18656), .B(n18657), .Z(n12212) );
  XNOR U18113 ( .A(n15658), .B(n12887), .Z(n18657) );
  XNOR U18114 ( .A(n18658), .B(n17104), .Z(n12887) );
  XNOR U18115 ( .A(n18659), .B(n17857), .Z(n17104) );
  ANDN U18116 ( .B(n17105), .A(n18660), .Z(n18658) );
  XOR U18117 ( .A(n18661), .B(n17095), .Z(n15658) );
  XNOR U18118 ( .A(n18662), .B(n18663), .Z(n17095) );
  XOR U18119 ( .A(n10004), .B(n18665), .Z(n18656) );
  XOR U18120 ( .A(n9357), .B(n14395), .Z(n18665) );
  XNOR U18121 ( .A(n18666), .B(n17090), .Z(n14395) );
  XNOR U18122 ( .A(n18667), .B(n16478), .Z(n17090) );
  ANDN U18123 ( .B(n17091), .A(n18668), .Z(n18666) );
  XNOR U18124 ( .A(n18669), .B(n18029), .Z(n9357) );
  XOR U18125 ( .A(n18670), .B(n17472), .Z(n18029) );
  XNOR U18126 ( .A(n18672), .B(n17100), .Z(n10004) );
  XNOR U18127 ( .A(n18637), .B(n18673), .Z(n17100) );
  ANDN U18128 ( .B(n18674), .A(n18675), .Z(n18672) );
  XOR U18129 ( .A(n18676), .B(n7699), .Z(n4092) );
  XNOR U18130 ( .A(n16868), .B(n10126), .Z(n7699) );
  XNOR U18131 ( .A(n15920), .B(n12369), .Z(n10126) );
  XNOR U18132 ( .A(n18677), .B(n18678), .Z(n12369) );
  XOR U18133 ( .A(n16639), .B(n11185), .Z(n18678) );
  XOR U18134 ( .A(n18679), .B(n16380), .Z(n11185) );
  IV U18135 ( .A(n17355), .Z(n16380) );
  XNOR U18136 ( .A(n18680), .B(n16465), .Z(n17355) );
  ANDN U18137 ( .B(n16874), .A(n16875), .Z(n18679) );
  XNOR U18138 ( .A(n18681), .B(n17407), .Z(n16875) );
  XNOR U18139 ( .A(n15607), .B(n18682), .Z(n16874) );
  XOR U18140 ( .A(n18683), .B(n18684), .Z(n15607) );
  XNOR U18141 ( .A(n18685), .B(n16388), .Z(n16639) );
  XOR U18142 ( .A(n18686), .B(n18394), .Z(n16388) );
  ANDN U18143 ( .B(n16870), .A(n16871), .Z(n18685) );
  XOR U18144 ( .A(n18687), .B(n17270), .Z(n16871) );
  XNOR U18145 ( .A(n17939), .B(n18688), .Z(n16870) );
  XOR U18146 ( .A(n18689), .B(n18690), .Z(n17939) );
  XNOR U18147 ( .A(n12918), .B(n18691), .Z(n18677) );
  XOR U18148 ( .A(n10664), .B(n17344), .Z(n18691) );
  XNOR U18149 ( .A(n18692), .B(n16371), .Z(n17344) );
  XOR U18150 ( .A(n18693), .B(n15122), .Z(n16371) );
  ANDN U18151 ( .B(n17353), .A(n17883), .Z(n18692) );
  XNOR U18152 ( .A(n18694), .B(n16375), .Z(n10664) );
  XOR U18153 ( .A(n18625), .B(n18695), .Z(n16375) );
  AND U18154 ( .A(n16861), .B(n16862), .Z(n18694) );
  XOR U18155 ( .A(n18696), .B(n18609), .Z(n16862) );
  XNOR U18156 ( .A(n18697), .B(n17933), .Z(n16861) );
  XNOR U18157 ( .A(n18698), .B(n17351), .Z(n12918) );
  XOR U18158 ( .A(n18699), .B(n17945), .Z(n17351) );
  ANDN U18159 ( .B(n16864), .A(n16865), .Z(n18698) );
  XOR U18160 ( .A(n18700), .B(n18651), .Z(n16865) );
  XOR U18161 ( .A(n18701), .B(n18702), .Z(n16864) );
  XOR U18162 ( .A(n18703), .B(n18704), .Z(n15920) );
  XNOR U18163 ( .A(n17009), .B(n12849), .Z(n18704) );
  XNOR U18164 ( .A(n18705), .B(n16693), .Z(n12849) );
  XOR U18165 ( .A(n18706), .B(n18707), .Z(n16693) );
  NOR U18166 ( .A(n15946), .B(n15945), .Z(n18705) );
  XOR U18167 ( .A(n18708), .B(n16053), .Z(n15945) );
  XOR U18168 ( .A(n18709), .B(n17031), .Z(n15946) );
  XNOR U18169 ( .A(n18710), .B(n16699), .Z(n17009) );
  XNOR U18170 ( .A(n18711), .B(n18712), .Z(n16699) );
  ANDN U18171 ( .B(n14321), .A(n14322), .Z(n18710) );
  XNOR U18172 ( .A(n18713), .B(n17469), .Z(n14322) );
  XNOR U18173 ( .A(n18403), .B(n18714), .Z(n14321) );
  XNOR U18174 ( .A(n12445), .B(n18715), .Z(n18703) );
  XOR U18175 ( .A(n12528), .B(n11122), .Z(n18715) );
  XNOR U18176 ( .A(n18716), .B(n16708), .Z(n11122) );
  XNOR U18177 ( .A(n18717), .B(n18718), .Z(n16708) );
  AND U18178 ( .A(n12812), .B(n12810), .Z(n18716) );
  XNOR U18179 ( .A(n18719), .B(n16100), .Z(n12810) );
  XNOR U18180 ( .A(n18720), .B(n18721), .Z(n12812) );
  XNOR U18181 ( .A(n18722), .B(n16703), .Z(n12528) );
  XOR U18182 ( .A(n18723), .B(n18022), .Z(n16703) );
  NOR U18183 ( .A(n12816), .B(n12817), .Z(n18722) );
  XNOR U18184 ( .A(n18724), .B(n18725), .Z(n12817) );
  XNOR U18185 ( .A(n18726), .B(n18727), .Z(n12816) );
  XNOR U18186 ( .A(n18728), .B(n16689), .Z(n12445) );
  XNOR U18187 ( .A(n18729), .B(n18730), .Z(n16689) );
  AND U18188 ( .A(n12820), .B(n12822), .Z(n18728) );
  XOR U18189 ( .A(n18625), .B(n18731), .Z(n12822) );
  XNOR U18190 ( .A(n18732), .B(n17520), .Z(n12820) );
  XNOR U18191 ( .A(n18733), .B(n17353), .Z(n16868) );
  XNOR U18192 ( .A(n18734), .B(n16003), .Z(n17353) );
  XNOR U18193 ( .A(n18735), .B(n18736), .Z(n16369) );
  XOR U18194 ( .A(n18737), .B(n18018), .Z(n17883) );
  ANDN U18195 ( .B(n7579), .A(n6828), .Z(n18676) );
  XNOR U18196 ( .A(n15708), .B(n11971), .Z(n6828) );
  IV U18197 ( .A(n11709), .Z(n11971) );
  XOR U18198 ( .A(n18738), .B(n12584), .Z(n11709) );
  XNOR U18199 ( .A(n18739), .B(n18740), .Z(n12584) );
  XOR U18200 ( .A(n12852), .B(n11143), .Z(n18740) );
  XOR U18201 ( .A(n18741), .B(n15165), .Z(n11143) );
  XNOR U18202 ( .A(n18742), .B(n16669), .Z(n15165) );
  IV U18203 ( .A(n18192), .Z(n16669) );
  ANDN U18204 ( .B(n15166), .A(n13780), .Z(n18741) );
  XOR U18205 ( .A(n18743), .B(n18744), .Z(n13780) );
  XOR U18206 ( .A(n18745), .B(n15591), .Z(n15166) );
  XNOR U18207 ( .A(n18746), .B(n15169), .Z(n12852) );
  ANDN U18208 ( .B(n15170), .A(n15703), .Z(n18746) );
  XNOR U18209 ( .A(n18750), .B(n17917), .Z(n15703) );
  XNOR U18210 ( .A(n18751), .B(n15336), .Z(n15170) );
  XNOR U18211 ( .A(n15161), .B(n18752), .Z(n18739) );
  XNOR U18212 ( .A(n11886), .B(n10994), .Z(n18752) );
  XOR U18213 ( .A(n18753), .B(n15180), .Z(n10994) );
  XNOR U18214 ( .A(n18755), .B(n15177), .Z(n11886) );
  XOR U18215 ( .A(n18756), .B(n18757), .Z(n15177) );
  ANDN U18216 ( .B(n15176), .A(n13774), .Z(n18755) );
  XNOR U18217 ( .A(n18758), .B(n18759), .Z(n13774) );
  XOR U18218 ( .A(n18625), .B(n18760), .Z(n15176) );
  XNOR U18219 ( .A(n18761), .B(n15174), .Z(n15161) );
  XNOR U18220 ( .A(n18762), .B(n18763), .Z(n15174) );
  ANDN U18221 ( .B(n13784), .A(n15173), .Z(n18761) );
  XNOR U18222 ( .A(n18764), .B(n18765), .Z(n15173) );
  XNOR U18223 ( .A(n18766), .B(n18022), .Z(n13784) );
  XOR U18224 ( .A(n18767), .B(n18533), .Z(n18022) );
  XOR U18225 ( .A(n18768), .B(n18769), .Z(n18533) );
  XNOR U18226 ( .A(n18770), .B(n18771), .Z(n18769) );
  XNOR U18227 ( .A(n14919), .B(n18772), .Z(n18768) );
  XNOR U18228 ( .A(n18773), .B(n18206), .Z(n18772) );
  XNOR U18229 ( .A(n18774), .B(n18775), .Z(n18206) );
  AND U18230 ( .A(n18776), .B(n18777), .Z(n18774) );
  XNOR U18231 ( .A(n18778), .B(n18779), .Z(n14919) );
  ANDN U18232 ( .B(n18780), .A(n18781), .Z(n18778) );
  XOR U18233 ( .A(n18782), .B(n15179), .Z(n15708) );
  XNOR U18234 ( .A(n18783), .B(n18236), .Z(n15179) );
  AND U18235 ( .A(n13770), .B(n18366), .Z(n18782) );
  IV U18236 ( .A(n13772), .Z(n18366) );
  XOR U18237 ( .A(n18784), .B(n16355), .Z(n13772) );
  XOR U18238 ( .A(n18785), .B(n18643), .Z(n13770) );
  XNOR U18239 ( .A(n12234), .B(n13257), .Z(n7579) );
  XOR U18240 ( .A(n18786), .B(n14842), .Z(n13257) );
  AND U18241 ( .A(n16508), .B(n18787), .Z(n18786) );
  XOR U18242 ( .A(n18788), .B(n17634), .Z(n16508) );
  IV U18243 ( .A(n18789), .Z(n17634) );
  XOR U18244 ( .A(n13467), .B(n13424), .Z(n12234) );
  XOR U18245 ( .A(n18790), .B(n18791), .Z(n13424) );
  XNOR U18246 ( .A(n9589), .B(n12574), .Z(n18791) );
  XOR U18247 ( .A(n18792), .B(n17670), .Z(n12574) );
  IV U18248 ( .A(n14834), .Z(n17670) );
  XOR U18249 ( .A(n18793), .B(n18002), .Z(n14834) );
  ANDN U18250 ( .B(n16510), .A(n13260), .Z(n18792) );
  XOR U18251 ( .A(n18794), .B(n17469), .Z(n13260) );
  IV U18252 ( .A(n13262), .Z(n16510) );
  XOR U18253 ( .A(n18795), .B(n18796), .Z(n13262) );
  XNOR U18254 ( .A(n18797), .B(n14837), .Z(n9589) );
  XNOR U18255 ( .A(n18798), .B(n17078), .Z(n14837) );
  AND U18256 ( .A(n13252), .B(n13250), .Z(n18797) );
  XOR U18257 ( .A(n17569), .B(n18799), .Z(n13250) );
  XOR U18258 ( .A(n18800), .B(n18801), .Z(n13252) );
  XOR U18259 ( .A(n12339), .B(n18802), .Z(n18790) );
  XOR U18260 ( .A(n9609), .B(n13813), .Z(n18802) );
  XOR U18261 ( .A(n18803), .B(n14845), .Z(n13813) );
  XNOR U18262 ( .A(n18804), .B(n18805), .Z(n14845) );
  ANDN U18263 ( .B(n13254), .A(n13255), .Z(n18803) );
  XOR U18264 ( .A(n18806), .B(n17186), .Z(n13255) );
  XNOR U18265 ( .A(n18588), .B(n18807), .Z(n13254) );
  XNOR U18266 ( .A(n18808), .B(n14841), .Z(n9609) );
  XNOR U18267 ( .A(n18809), .B(n16779), .Z(n14841) );
  XOR U18268 ( .A(n18810), .B(n18439), .Z(n14842) );
  IV U18269 ( .A(n18787), .Z(n16507) );
  XOR U18270 ( .A(n18811), .B(n18135), .Z(n18787) );
  XNOR U18271 ( .A(n18812), .B(n14848), .Z(n12339) );
  XNOR U18272 ( .A(n18044), .B(n18813), .Z(n14848) );
  ANDN U18273 ( .B(n13264), .A(n13265), .Z(n18812) );
  XNOR U18274 ( .A(n18814), .B(n15137), .Z(n13265) );
  XNOR U18275 ( .A(n18815), .B(n18816), .Z(n13264) );
  XOR U18276 ( .A(n18817), .B(n18818), .Z(n13467) );
  XOR U18277 ( .A(n11974), .B(n12975), .Z(n18818) );
  XOR U18278 ( .A(n18819), .B(n13830), .Z(n12975) );
  IV U18279 ( .A(n18564), .Z(n13830) );
  XOR U18280 ( .A(n18820), .B(n18323), .Z(n18564) );
  NOR U18281 ( .A(n13829), .B(n14696), .Z(n18819) );
  XOR U18282 ( .A(n18821), .B(n17730), .Z(n14696) );
  XNOR U18283 ( .A(n18822), .B(n17380), .Z(n13829) );
  XOR U18284 ( .A(n18824), .B(n18825), .Z(n13821) );
  ANDN U18285 ( .B(n15697), .A(n13820), .Z(n18823) );
  XOR U18286 ( .A(n18826), .B(n15244), .Z(n13820) );
  IV U18287 ( .A(n14700), .Z(n15697) );
  XOR U18288 ( .A(n18827), .B(n18789), .Z(n14700) );
  XOR U18289 ( .A(n11697), .B(n18828), .Z(n18817) );
  XOR U18290 ( .A(n11719), .B(n11549), .Z(n18828) );
  XOR U18291 ( .A(n18829), .B(n18558), .Z(n11549) );
  IV U18292 ( .A(n18575), .Z(n18558) );
  XOR U18293 ( .A(n18830), .B(n18376), .Z(n18575) );
  AND U18294 ( .A(n14702), .B(n14704), .Z(n18829) );
  XNOR U18295 ( .A(n18831), .B(n18832), .Z(n14704) );
  XOR U18296 ( .A(n16348), .B(n18833), .Z(n14702) );
  XOR U18297 ( .A(n18834), .B(n13826), .Z(n11719) );
  XOR U18298 ( .A(n17841), .B(n18835), .Z(n13826) );
  XNOR U18299 ( .A(n18836), .B(n18736), .Z(n14689) );
  XNOR U18300 ( .A(n18837), .B(n18473), .Z(n13825) );
  XOR U18301 ( .A(n18839), .B(n17203), .Z(n13834) );
  NOR U18302 ( .A(n13833), .B(n14692), .Z(n18838) );
  XNOR U18303 ( .A(n14918), .B(n18770), .Z(n14692) );
  XNOR U18304 ( .A(n18840), .B(n18841), .Z(n18770) );
  ANDN U18305 ( .B(n18842), .A(n18843), .Z(n18840) );
  XNOR U18306 ( .A(n18844), .B(n17667), .Z(n13833) );
  XOR U18307 ( .A(n18845), .B(n6807), .Z(n7589) );
  XNOR U18308 ( .A(n11649), .B(n14220), .Z(n6807) );
  XNOR U18309 ( .A(n18846), .B(n14189), .Z(n14220) );
  ANDN U18310 ( .B(n17201), .A(n17180), .Z(n18846) );
  XOR U18311 ( .A(n18847), .B(n16340), .Z(n17180) );
  XNOR U18312 ( .A(n18848), .B(n18849), .Z(n16340) );
  XOR U18313 ( .A(n17297), .B(n18500), .Z(n11649) );
  XNOR U18314 ( .A(n18850), .B(n18851), .Z(n18500) );
  XOR U18315 ( .A(n9770), .B(n12705), .Z(n18851) );
  XNOR U18316 ( .A(n18852), .B(n13531), .Z(n12705) );
  XNOR U18317 ( .A(n18853), .B(n15843), .Z(n13531) );
  ANDN U18318 ( .B(n14186), .A(n16800), .Z(n18852) );
  XOR U18319 ( .A(n18854), .B(n13991), .Z(n16800) );
  IV U18320 ( .A(n17514), .Z(n13991) );
  XOR U18321 ( .A(n18857), .B(n18002), .Z(n14186) );
  XOR U18322 ( .A(n18858), .B(n14184), .Z(n9770) );
  IV U18323 ( .A(n13524), .Z(n14184) );
  XNOR U18324 ( .A(n18859), .B(n16555), .Z(n13524) );
  NOR U18325 ( .A(n14183), .B(n14228), .Z(n18858) );
  XNOR U18326 ( .A(n18860), .B(n16039), .Z(n14228) );
  XNOR U18327 ( .A(n15592), .B(n18861), .Z(n14183) );
  XNOR U18328 ( .A(n12984), .B(n18862), .Z(n18850) );
  XNOR U18329 ( .A(n11780), .B(n9897), .Z(n18862) );
  XNOR U18330 ( .A(n18863), .B(n14177), .Z(n9897) );
  XOR U18331 ( .A(n18864), .B(n17467), .Z(n14177) );
  AND U18332 ( .A(n14226), .B(n14178), .Z(n18863) );
  XNOR U18333 ( .A(n18865), .B(n18394), .Z(n14178) );
  XNOR U18334 ( .A(n18866), .B(n18867), .Z(n18394) );
  XNOR U18335 ( .A(n18868), .B(n18869), .Z(n14226) );
  XNOR U18336 ( .A(n18870), .B(n14190), .Z(n11780) );
  XOR U18337 ( .A(n15598), .B(n18871), .Z(n14190) );
  ANDN U18338 ( .B(n14189), .A(n17201), .Z(n18870) );
  XNOR U18339 ( .A(n18872), .B(n16944), .Z(n17201) );
  XOR U18340 ( .A(n18873), .B(n18727), .Z(n14189) );
  XOR U18341 ( .A(n18874), .B(n13520), .Z(n12984) );
  XOR U18342 ( .A(n18875), .B(n18876), .Z(n13520) );
  AND U18343 ( .A(n14622), .B(n14180), .Z(n18874) );
  XNOR U18344 ( .A(n18877), .B(n18258), .Z(n14180) );
  XOR U18345 ( .A(n18878), .B(n18879), .Z(n14622) );
  XOR U18346 ( .A(n18880), .B(n18881), .Z(n17297) );
  XOR U18347 ( .A(n13848), .B(n15053), .Z(n18881) );
  XOR U18348 ( .A(n18882), .B(n15068), .Z(n15053) );
  XOR U18349 ( .A(n18883), .B(n17661), .Z(n15068) );
  IV U18350 ( .A(n16456), .Z(n17661) );
  XNOR U18351 ( .A(n18884), .B(n18885), .Z(n16456) );
  NOR U18352 ( .A(n14243), .B(n14242), .Z(n18882) );
  XNOR U18353 ( .A(n18886), .B(n18011), .Z(n14242) );
  XNOR U18354 ( .A(n17081), .B(n18887), .Z(n14243) );
  XNOR U18355 ( .A(n18888), .B(n15059), .Z(n13848) );
  XOR U18356 ( .A(n18889), .B(n18462), .Z(n15059) );
  NOR U18357 ( .A(n14237), .B(n14236), .Z(n18888) );
  XNOR U18358 ( .A(n17860), .B(n18890), .Z(n14236) );
  XNOR U18359 ( .A(n18891), .B(n16795), .Z(n14237) );
  XOR U18360 ( .A(n13855), .B(n18892), .Z(n18880) );
  XOR U18361 ( .A(n12791), .B(n12073), .Z(n18892) );
  XOR U18362 ( .A(n18893), .B(n16587), .Z(n12073) );
  XNOR U18363 ( .A(n18894), .B(n18895), .Z(n16587) );
  XOR U18364 ( .A(n17402), .B(n18896), .Z(n14232) );
  XOR U18365 ( .A(n18897), .B(n18578), .Z(n14233) );
  XNOR U18366 ( .A(n18898), .B(n15062), .Z(n12791) );
  XNOR U18367 ( .A(n18899), .B(n16552), .Z(n15062) );
  ANDN U18368 ( .B(n15063), .A(n17300), .Z(n18898) );
  XNOR U18369 ( .A(n17192), .B(n18900), .Z(n17300) );
  XNOR U18370 ( .A(n18901), .B(n18279), .Z(n15063) );
  XNOR U18371 ( .A(n18902), .B(n15071), .Z(n13855) );
  XNOR U18372 ( .A(n18903), .B(n18904), .Z(n15071) );
  XOR U18373 ( .A(n17190), .B(n18905), .Z(n14246) );
  XNOR U18374 ( .A(n18906), .B(n18712), .Z(n14247) );
  IV U18375 ( .A(n15333), .Z(n18712) );
  NOR U18376 ( .A(n9934), .B(n7510), .Z(n18845) );
  XOR U18377 ( .A(n14311), .B(n12137), .Z(n7510) );
  XOR U18378 ( .A(n18909), .B(n18910), .Z(n14311) );
  ANDN U18379 ( .B(n17431), .A(n12436), .Z(n18909) );
  XNOR U18380 ( .A(n18911), .B(n17458), .Z(n12436) );
  XOR U18381 ( .A(n18914), .B(n18915), .Z(n9934) );
  XNOR U18382 ( .A(n1800), .B(n9203), .Z(n4065) );
  XNOR U18383 ( .A(n18916), .B(n9262), .Z(n9203) );
  ANDN U18384 ( .B(n7076), .A(n6612), .Z(n18916) );
  XNOR U18385 ( .A(n9576), .B(n18917), .Z(n6612) );
  IV U18386 ( .A(n18914), .Z(n9576) );
  XOR U18387 ( .A(n12621), .B(n14604), .Z(n18914) );
  XOR U18388 ( .A(n18918), .B(n18919), .Z(n14604) );
  XNOR U18389 ( .A(n16409), .B(n11897), .Z(n18919) );
  XNOR U18390 ( .A(n18920), .B(n18581), .Z(n11897) );
  AND U18391 ( .A(n15501), .B(n18582), .Z(n18920) );
  XNOR U18392 ( .A(n18921), .B(n16429), .Z(n16409) );
  XNOR U18393 ( .A(n10119), .B(n18922), .Z(n18918) );
  XOR U18394 ( .A(n9376), .B(n10832), .Z(n18922) );
  XOR U18395 ( .A(n18923), .B(n16433), .Z(n10832) );
  ANDN U18396 ( .B(n18924), .A(n15505), .Z(n18923) );
  XNOR U18397 ( .A(n18925), .B(n18926), .Z(n9376) );
  ANDN U18398 ( .B(n18927), .A(n15496), .Z(n18925) );
  XNOR U18399 ( .A(n18928), .B(n16436), .Z(n10119) );
  ANDN U18400 ( .B(n16437), .A(n15492), .Z(n18928) );
  XOR U18401 ( .A(n18929), .B(n18930), .Z(n12621) );
  XNOR U18402 ( .A(n12681), .B(n15368), .Z(n18930) );
  XOR U18403 ( .A(n18931), .B(n15385), .Z(n15368) );
  IV U18404 ( .A(n17781), .Z(n15385) );
  XOR U18405 ( .A(n18932), .B(n16041), .Z(n17781) );
  NOR U18406 ( .A(n15384), .B(n14042), .Z(n18931) );
  IV U18407 ( .A(n18933), .Z(n15384) );
  XNOR U18408 ( .A(n18934), .B(n15389), .Z(n12681) );
  XNOR U18409 ( .A(n18935), .B(n18252), .Z(n15389) );
  AND U18410 ( .A(n15388), .B(n14540), .Z(n18934) );
  IV U18411 ( .A(n18936), .Z(n14540) );
  XOR U18412 ( .A(n12055), .B(n18937), .Z(n18929) );
  XNOR U18413 ( .A(n10713), .B(n14436), .Z(n18937) );
  XNOR U18414 ( .A(n18938), .B(n15378), .Z(n14436) );
  XNOR U18415 ( .A(n18939), .B(n18940), .Z(n15378) );
  NOR U18416 ( .A(n15377), .B(n18941), .Z(n18938) );
  IV U18417 ( .A(n18942), .Z(n15377) );
  XOR U18418 ( .A(n18943), .B(n17790), .Z(n10713) );
  IV U18419 ( .A(n15382), .Z(n17790) );
  XOR U18420 ( .A(n18743), .B(n18944), .Z(n15382) );
  XOR U18421 ( .A(n18945), .B(n15374), .Z(n12055) );
  XNOR U18422 ( .A(n18946), .B(n16053), .Z(n15374) );
  XOR U18423 ( .A(n18947), .B(n18948), .Z(n16053) );
  ANDN U18424 ( .B(n14046), .A(n15373), .Z(n18945) );
  IV U18425 ( .A(n18949), .Z(n14046) );
  IV U18426 ( .A(n3869), .Z(n1800) );
  XOR U18427 ( .A(n6580), .B(n6315), .Z(n3869) );
  XOR U18428 ( .A(n18950), .B(n18951), .Z(n6315) );
  XNOR U18429 ( .A(n5890), .B(n4301), .Z(n18951) );
  XNOR U18430 ( .A(n18952), .B(n7170), .Z(n4301) );
  XNOR U18431 ( .A(n16119), .B(n11067), .Z(n7170) );
  IV U18432 ( .A(n12282), .Z(n11067) );
  XOR U18433 ( .A(n16196), .B(n12077), .Z(n12282) );
  XNOR U18434 ( .A(n18953), .B(n18954), .Z(n12077) );
  XOR U18435 ( .A(n11286), .B(n11137), .Z(n18954) );
  XOR U18436 ( .A(n18955), .B(n12491), .Z(n11137) );
  XNOR U18437 ( .A(n18956), .B(n16331), .Z(n12491) );
  IV U18438 ( .A(n15851), .Z(n16331) );
  ANDN U18439 ( .B(n14298), .A(n14299), .Z(n18955) );
  XNOR U18440 ( .A(n18957), .B(n17517), .Z(n14299) );
  XNOR U18441 ( .A(n18958), .B(n17678), .Z(n14298) );
  XNOR U18442 ( .A(n18959), .B(n12487), .Z(n11286) );
  XOR U18443 ( .A(n18960), .B(n18718), .Z(n12487) );
  ANDN U18444 ( .B(n12488), .A(n14293), .Z(n18959) );
  XOR U18445 ( .A(n18961), .B(n15843), .Z(n14293) );
  XNOR U18446 ( .A(n17126), .B(n18962), .Z(n12488) );
  XOR U18447 ( .A(n10278), .B(n18963), .Z(n18953) );
  XNOR U18448 ( .A(n11325), .B(n11111), .Z(n18963) );
  XNOR U18449 ( .A(n18964), .B(n12497), .Z(n11111) );
  XOR U18450 ( .A(n18965), .B(n17407), .Z(n12497) );
  AND U18451 ( .A(n12496), .B(n14295), .Z(n18964) );
  XNOR U18452 ( .A(n18966), .B(n17415), .Z(n14295) );
  XNOR U18453 ( .A(n18967), .B(n18162), .Z(n12496) );
  XNOR U18454 ( .A(n18968), .B(n12500), .Z(n11325) );
  XNOR U18455 ( .A(n18969), .B(n18095), .Z(n12500) );
  AND U18456 ( .A(n14288), .B(n14287), .Z(n18968) );
  XOR U18457 ( .A(n18970), .B(n16552), .Z(n14287) );
  XNOR U18458 ( .A(n18971), .B(n18972), .Z(n16552) );
  XNOR U18459 ( .A(n14944), .B(n18973), .Z(n14288) );
  XNOR U18460 ( .A(n18974), .B(n12505), .Z(n10278) );
  XNOR U18461 ( .A(n18975), .B(n18976), .Z(n12505) );
  ANDN U18462 ( .B(n14290), .A(n12504), .Z(n18974) );
  XOR U18463 ( .A(n18977), .B(n17360), .Z(n12504) );
  XOR U18464 ( .A(n18980), .B(n18609), .Z(n14290) );
  XOR U18465 ( .A(n18981), .B(n18982), .Z(n16196) );
  XNOR U18466 ( .A(n11647), .B(n10458), .Z(n18982) );
  XNOR U18467 ( .A(n18983), .B(n12514), .Z(n10458) );
  XNOR U18468 ( .A(n18984), .B(n18095), .Z(n12514) );
  IV U18469 ( .A(n18727), .Z(n18095) );
  XNOR U18470 ( .A(n18985), .B(n18986), .Z(n18727) );
  ANDN U18471 ( .B(n12515), .A(n16121), .Z(n18983) );
  XOR U18472 ( .A(n18987), .B(n18254), .Z(n12515) );
  XNOR U18473 ( .A(n18988), .B(n13195), .Z(n11647) );
  XNOR U18474 ( .A(n18989), .B(n16453), .Z(n13195) );
  AND U18475 ( .A(n13196), .B(n16123), .Z(n18988) );
  XOR U18476 ( .A(n18990), .B(n18991), .Z(n13196) );
  XOR U18477 ( .A(n9188), .B(n18992), .Z(n18981) );
  XNOR U18478 ( .A(n12482), .B(n9708), .Z(n18992) );
  XNOR U18479 ( .A(n18993), .B(n12802), .Z(n9708) );
  XOR U18480 ( .A(n18994), .B(n15631), .Z(n12802) );
  ANDN U18481 ( .B(n12803), .A(n18995), .Z(n18993) );
  XNOR U18482 ( .A(n18996), .B(n12519), .Z(n12482) );
  XNOR U18483 ( .A(n18997), .B(n17730), .Z(n12519) );
  ANDN U18484 ( .B(n18998), .A(n12518), .Z(n18996) );
  XNOR U18485 ( .A(n18999), .B(n18109), .Z(n12518) );
  XNOR U18486 ( .A(n19000), .B(n13582), .Z(n9188) );
  XNOR U18487 ( .A(n19001), .B(n16337), .Z(n13582) );
  AND U18488 ( .A(n13585), .B(n16114), .Z(n19000) );
  XOR U18489 ( .A(n19002), .B(n17016), .Z(n13585) );
  IV U18490 ( .A(n15213), .Z(n17016) );
  XNOR U18491 ( .A(n19003), .B(n12803), .Z(n16119) );
  XNOR U18492 ( .A(n19004), .B(n17441), .Z(n12803) );
  AND U18493 ( .A(n18995), .B(n13572), .Z(n19003) );
  IV U18494 ( .A(n19005), .Z(n13572) );
  NOR U18495 ( .A(n6656), .B(n6657), .Z(n18952) );
  XNOR U18496 ( .A(n14868), .B(n10055), .Z(n6657) );
  XNOR U18497 ( .A(n14685), .B(n19006), .Z(n10055) );
  XOR U18498 ( .A(n19007), .B(n19008), .Z(n14685) );
  XNOR U18499 ( .A(n9804), .B(n13021), .Z(n19008) );
  XNOR U18500 ( .A(n19009), .B(n15774), .Z(n13021) );
  XOR U18501 ( .A(n17258), .B(n19010), .Z(n15774) );
  ANDN U18502 ( .B(n15773), .A(n18548), .Z(n19009) );
  XNOR U18503 ( .A(n19011), .B(n15777), .Z(n9804) );
  XOR U18504 ( .A(n19012), .B(n18510), .Z(n15777) );
  ANDN U18505 ( .B(n14860), .A(n14861), .Z(n19011) );
  XNOR U18506 ( .A(n19013), .B(n18759), .Z(n14861) );
  XOR U18507 ( .A(n19014), .B(n17879), .Z(n14860) );
  IV U18508 ( .A(n17855), .Z(n17879) );
  XNOR U18509 ( .A(n19015), .B(n19016), .Z(n17855) );
  XNOR U18510 ( .A(n15749), .B(n19017), .Z(n19007) );
  XNOR U18511 ( .A(n9821), .B(n12736), .Z(n19017) );
  XNOR U18512 ( .A(n19018), .B(n15782), .Z(n12736) );
  XNOR U18513 ( .A(n19019), .B(n19020), .Z(n15782) );
  ANDN U18514 ( .B(n14870), .A(n14871), .Z(n19018) );
  XNOR U18515 ( .A(n19021), .B(n18334), .Z(n14871) );
  XNOR U18516 ( .A(n19022), .B(n18765), .Z(n14870) );
  IV U18517 ( .A(n19023), .Z(n18765) );
  XNOR U18518 ( .A(n19024), .B(n16735), .Z(n9821) );
  XNOR U18519 ( .A(n19025), .B(n15644), .Z(n16735) );
  IV U18520 ( .A(n17380), .Z(n15644) );
  XNOR U18521 ( .A(n19026), .B(n19027), .Z(n17380) );
  AND U18522 ( .A(n14876), .B(n14874), .Z(n19024) );
  XNOR U18523 ( .A(n19028), .B(n19029), .Z(n14874) );
  XNOR U18524 ( .A(n17234), .B(n19030), .Z(n14876) );
  XNOR U18525 ( .A(n19031), .B(n15785), .Z(n15749) );
  XNOR U18526 ( .A(n16758), .B(n19032), .Z(n15785) );
  XNOR U18527 ( .A(n19033), .B(n16060), .Z(n14865) );
  IV U18528 ( .A(n17869), .Z(n16060) );
  XOR U18529 ( .A(n19034), .B(n16907), .Z(n14864) );
  IV U18530 ( .A(n16603), .Z(n16907) );
  XNOR U18531 ( .A(n19035), .B(n15773), .Z(n14868) );
  XOR U18532 ( .A(n19036), .B(n17555), .Z(n15773) );
  AND U18533 ( .A(n16729), .B(n18548), .Z(n19035) );
  XNOR U18534 ( .A(n17192), .B(n19037), .Z(n18548) );
  XOR U18535 ( .A(n19038), .B(n18736), .Z(n16729) );
  XNOR U18536 ( .A(n19039), .B(n11875), .Z(n6656) );
  XOR U18537 ( .A(n19040), .B(n7179), .Z(n5890) );
  XOR U18538 ( .A(n9201), .B(n18070), .Z(n7179) );
  XNOR U18539 ( .A(n19041), .B(n16648), .Z(n18070) );
  AND U18540 ( .A(n19042), .B(n15867), .Z(n19041) );
  IV U18541 ( .A(n11449), .Z(n9201) );
  XOR U18542 ( .A(n12980), .B(n16152), .Z(n11449) );
  XOR U18543 ( .A(n19043), .B(n19044), .Z(n16152) );
  XNOR U18544 ( .A(n13992), .B(n14853), .Z(n19044) );
  XOR U18545 ( .A(n19045), .B(n15869), .Z(n14853) );
  IV U18546 ( .A(n16649), .Z(n15869) );
  XOR U18547 ( .A(n19046), .B(n15987), .Z(n16649) );
  IV U18548 ( .A(n18252), .Z(n15987) );
  XOR U18549 ( .A(n19047), .B(n19048), .Z(n18252) );
  NOR U18550 ( .A(n19042), .B(n16648), .Z(n19045) );
  XNOR U18551 ( .A(n19049), .B(n19050), .Z(n16648) );
  XOR U18552 ( .A(n19051), .B(n15877), .Z(n13992) );
  XOR U18553 ( .A(n19052), .B(n18736), .Z(n15877) );
  NOR U18554 ( .A(n16652), .B(n18069), .Z(n19051) );
  XNOR U18555 ( .A(n19053), .B(n15597), .Z(n16652) );
  XOR U18556 ( .A(n11306), .B(n19054), .Z(n19043) );
  XOR U18557 ( .A(n11191), .B(n14974), .Z(n19054) );
  XOR U18558 ( .A(n19055), .B(n15873), .Z(n14974) );
  XNOR U18559 ( .A(n19056), .B(n19057), .Z(n15873) );
  ANDN U18560 ( .B(n16654), .A(n18067), .Z(n19055) );
  XNOR U18561 ( .A(n19058), .B(n19059), .Z(n16654) );
  XOR U18562 ( .A(n19060), .B(n15881), .Z(n11191) );
  XOR U18563 ( .A(n17491), .B(n19061), .Z(n15881) );
  ANDN U18564 ( .B(n18073), .A(n16656), .Z(n19060) );
  XNOR U18565 ( .A(n19062), .B(n18473), .Z(n16656) );
  XOR U18566 ( .A(n19063), .B(n15885), .Z(n11306) );
  IV U18567 ( .A(n16646), .Z(n15885) );
  XOR U18568 ( .A(n19064), .B(n17035), .Z(n16646) );
  ANDN U18569 ( .B(n19065), .A(n16645), .Z(n19063) );
  XOR U18570 ( .A(n19066), .B(n17144), .Z(n16645) );
  XOR U18571 ( .A(n19067), .B(n19068), .Z(n12980) );
  XNOR U18572 ( .A(n9923), .B(n11532), .Z(n19068) );
  XOR U18573 ( .A(n19069), .B(n14985), .Z(n11532) );
  ANDN U18574 ( .B(n18084), .A(n16148), .Z(n19069) );
  XNOR U18575 ( .A(n15824), .B(n19070), .Z(n16148) );
  XNOR U18576 ( .A(n19071), .B(n19072), .Z(n15824) );
  XNOR U18577 ( .A(n19073), .B(n16252), .Z(n18084) );
  XNOR U18578 ( .A(n19074), .B(n19075), .Z(n16252) );
  ANDN U18579 ( .B(n19077), .A(n14994), .Z(n19076) );
  XNOR U18580 ( .A(n19078), .B(n17426), .Z(n14994) );
  IV U18581 ( .A(n17517), .Z(n17426) );
  IV U18582 ( .A(n16137), .Z(n19077) );
  XOR U18583 ( .A(n19079), .B(n17509), .Z(n16137) );
  XOR U18584 ( .A(n10032), .B(n19080), .Z(n19067) );
  XNOR U18585 ( .A(n10888), .B(n10684), .Z(n19080) );
  XOR U18586 ( .A(n19081), .B(n19082), .Z(n10684) );
  ANDN U18587 ( .B(n16144), .A(n18086), .Z(n19081) );
  IV U18588 ( .A(n18087), .Z(n16144) );
  XNOR U18589 ( .A(n19083), .B(n16478), .Z(n18087) );
  XOR U18590 ( .A(n19084), .B(n19027), .Z(n16478) );
  XNOR U18591 ( .A(n19085), .B(n19086), .Z(n19027) );
  XOR U18592 ( .A(n13882), .B(n17544), .Z(n19086) );
  XOR U18593 ( .A(n19087), .B(n19088), .Z(n17544) );
  AND U18594 ( .A(n19089), .B(n19090), .Z(n19087) );
  XNOR U18595 ( .A(n19091), .B(n19092), .Z(n13882) );
  AND U18596 ( .A(n19093), .B(n19094), .Z(n19091) );
  XOR U18597 ( .A(n18371), .B(n19095), .Z(n19085) );
  XOR U18598 ( .A(n18504), .B(n19096), .Z(n19095) );
  XNOR U18599 ( .A(n19097), .B(n19098), .Z(n18504) );
  ANDN U18600 ( .B(n19099), .A(n19100), .Z(n19097) );
  XNOR U18601 ( .A(n19101), .B(n19102), .Z(n18371) );
  ANDN U18602 ( .B(n19103), .A(n19104), .Z(n19101) );
  XNOR U18603 ( .A(n19105), .B(n14980), .Z(n10888) );
  NOR U18604 ( .A(n14981), .B(n16141), .Z(n19105) );
  XNOR U18605 ( .A(n19106), .B(n19107), .Z(n16141) );
  IV U18606 ( .A(n18082), .Z(n14981) );
  XOR U18607 ( .A(n19108), .B(n18423), .Z(n18082) );
  XNOR U18608 ( .A(n19109), .B(n14990), .Z(n10032) );
  ANDN U18609 ( .B(n14991), .A(n16134), .Z(n19109) );
  XNOR U18610 ( .A(n19110), .B(n18406), .Z(n16134) );
  XOR U18611 ( .A(n19111), .B(n18425), .Z(n14991) );
  AND U18612 ( .A(n6641), .B(n6639), .Z(n19040) );
  XOR U18613 ( .A(n16426), .B(n9687), .Z(n6639) );
  XOR U18614 ( .A(n19112), .B(n19113), .Z(n12843) );
  XNOR U18615 ( .A(n12922), .B(n10253), .Z(n19113) );
  XNOR U18616 ( .A(n19114), .B(n15506), .Z(n10253) );
  ANDN U18617 ( .B(n15507), .A(n16433), .Z(n19114) );
  XNOR U18618 ( .A(n19115), .B(n17903), .Z(n16433) );
  XNOR U18619 ( .A(n19116), .B(n18832), .Z(n15507) );
  XNOR U18620 ( .A(n19117), .B(n15511), .Z(n12922) );
  AND U18621 ( .A(n15510), .B(n16429), .Z(n19117) );
  XOR U18622 ( .A(n17841), .B(n19118), .Z(n16429) );
  IV U18623 ( .A(n18099), .Z(n17841) );
  XOR U18624 ( .A(n19119), .B(n19120), .Z(n18099) );
  XNOR U18625 ( .A(n19121), .B(n18034), .Z(n15510) );
  XNOR U18626 ( .A(n12190), .B(n19122), .Z(n19112) );
  XOR U18627 ( .A(n10812), .B(n15488), .Z(n19122) );
  XNOR U18628 ( .A(n19123), .B(n15498), .Z(n15488) );
  AND U18629 ( .A(n18926), .B(n19124), .Z(n19123) );
  XNOR U18630 ( .A(n19125), .B(n15503), .Z(n10812) );
  ANDN U18631 ( .B(n18581), .A(n15502), .Z(n19125) );
  XNOR U18632 ( .A(n19126), .B(n17149), .Z(n15502) );
  XOR U18633 ( .A(n19127), .B(n16460), .Z(n18581) );
  XNOR U18634 ( .A(n19128), .B(n15494), .Z(n12190) );
  ANDN U18635 ( .B(n16436), .A(n15493), .Z(n19128) );
  XNOR U18636 ( .A(n19129), .B(n18347), .Z(n15493) );
  XOR U18637 ( .A(n19130), .B(n18976), .Z(n16436) );
  XNOR U18638 ( .A(n19131), .B(n19132), .Z(n17460) );
  XOR U18639 ( .A(n9512), .B(n10263), .Z(n19132) );
  XOR U18640 ( .A(n19133), .B(n13177), .Z(n10263) );
  XOR U18641 ( .A(n17003), .B(n19134), .Z(n13177) );
  ANDN U18642 ( .B(n15526), .A(n14608), .Z(n19133) );
  XOR U18643 ( .A(n19135), .B(n18643), .Z(n14608) );
  XOR U18644 ( .A(n17557), .B(n19136), .Z(n15526) );
  XNOR U18645 ( .A(n19137), .B(n13169), .Z(n9512) );
  XNOR U18646 ( .A(n19138), .B(n18439), .Z(n13169) );
  IV U18647 ( .A(n15336), .Z(n18439) );
  XNOR U18648 ( .A(n19139), .B(n19140), .Z(n15336) );
  AND U18649 ( .A(n14610), .B(n15530), .Z(n19137) );
  XOR U18650 ( .A(n17887), .B(n19141), .Z(n15530) );
  XNOR U18651 ( .A(n18347), .B(n19142), .Z(n14610) );
  XNOR U18652 ( .A(n10946), .B(n19143), .Z(n19131) );
  XNOR U18653 ( .A(n12539), .B(n12059), .Z(n19143) );
  XNOR U18654 ( .A(n19144), .B(n13173), .Z(n12059) );
  XNOR U18655 ( .A(n17464), .B(n19145), .Z(n13173) );
  IV U18656 ( .A(n16323), .Z(n17464) );
  ANDN U18657 ( .B(n15521), .A(n14614), .Z(n19144) );
  XOR U18658 ( .A(n19146), .B(n18180), .Z(n14614) );
  XNOR U18659 ( .A(n17959), .B(n19147), .Z(n15521) );
  XNOR U18660 ( .A(n19148), .B(n13326), .Z(n12539) );
  XNOR U18661 ( .A(n17234), .B(n19149), .Z(n13326) );
  ANDN U18662 ( .B(n15517), .A(n14619), .Z(n19148) );
  XNOR U18663 ( .A(n19150), .B(n19151), .Z(n14619) );
  IV U18664 ( .A(n16422), .Z(n15517) );
  XOR U18665 ( .A(n19152), .B(n17903), .Z(n16422) );
  IV U18666 ( .A(n18869), .Z(n17903) );
  XNOR U18667 ( .A(n19153), .B(n13164), .Z(n10946) );
  XNOR U18668 ( .A(n19154), .B(n16940), .Z(n13164) );
  ANDN U18669 ( .B(n15534), .A(n14616), .Z(n19153) );
  XNOR U18670 ( .A(n19155), .B(n19156), .Z(n14616) );
  XNOR U18671 ( .A(n19157), .B(n16954), .Z(n15534) );
  XOR U18672 ( .A(n19158), .B(n15497), .Z(n16426) );
  IV U18673 ( .A(n19124), .Z(n15497) );
  XOR U18674 ( .A(n19159), .B(n19160), .Z(n19124) );
  NOR U18675 ( .A(n18927), .B(n18926), .Z(n19158) );
  XOR U18676 ( .A(n19161), .B(n18389), .Z(n18926) );
  XNOR U18677 ( .A(n14312), .B(n12137), .Z(n6641) );
  XNOR U18678 ( .A(n12076), .B(n17637), .Z(n12137) );
  XNOR U18679 ( .A(n19162), .B(n19163), .Z(n17637) );
  XOR U18680 ( .A(n11919), .B(n12925), .Z(n19163) );
  XOR U18681 ( .A(n19164), .B(n18675), .Z(n12925) );
  AND U18682 ( .A(n18051), .B(n17099), .Z(n19164) );
  XNOR U18683 ( .A(n19165), .B(n16003), .Z(n17099) );
  XOR U18684 ( .A(n19166), .B(n19167), .Z(n16003) );
  XNOR U18685 ( .A(n19168), .B(n18660), .Z(n11919) );
  AND U18686 ( .A(n18054), .B(n18053), .Z(n19168) );
  IV U18687 ( .A(n19169), .Z(n18053) );
  IV U18688 ( .A(n17103), .Z(n18054) );
  XNOR U18689 ( .A(n19170), .B(n16039), .Z(n17103) );
  XOR U18690 ( .A(n11459), .B(n19171), .Z(n19162) );
  XOR U18691 ( .A(n9586), .B(n12149), .Z(n19171) );
  XNOR U18692 ( .A(n19172), .B(n18671), .Z(n12149) );
  ANDN U18693 ( .B(n19173), .A(n18028), .Z(n19172) );
  XOR U18694 ( .A(n19174), .B(n16940), .Z(n18028) );
  IV U18695 ( .A(n18904), .Z(n16940) );
  XNOR U18696 ( .A(n19177), .B(n18668), .Z(n9586) );
  XOR U18697 ( .A(n19178), .B(n17583), .Z(n17089) );
  XNOR U18698 ( .A(n19179), .B(n18664), .Z(n11459) );
  XOR U18699 ( .A(n19180), .B(n15213), .Z(n17093) );
  XOR U18700 ( .A(n19181), .B(n19182), .Z(n15213) );
  XOR U18701 ( .A(n19183), .B(n19184), .Z(n12076) );
  XNOR U18702 ( .A(n14823), .B(n12661), .Z(n19184) );
  XOR U18703 ( .A(n19185), .B(n19186), .Z(n12661) );
  ANDN U18704 ( .B(n14314), .A(n14315), .Z(n19185) );
  XNOR U18705 ( .A(n19187), .B(n19188), .Z(n14315) );
  XNOR U18706 ( .A(n19189), .B(n17107), .Z(n14823) );
  XOR U18707 ( .A(n17445), .B(n19190), .Z(n14308) );
  XOR U18708 ( .A(n15158), .B(n19191), .Z(n19183) );
  XOR U18709 ( .A(n19192), .B(n13598), .Z(n19191) );
  XNOR U18710 ( .A(n19193), .B(n12437), .Z(n13598) );
  NOR U18711 ( .A(n17431), .B(n18910), .Z(n19193) );
  XNOR U18712 ( .A(n19194), .B(n18215), .Z(n17431) );
  XOR U18713 ( .A(n19195), .B(n12423), .Z(n15158) );
  ANDN U18714 ( .B(n19196), .A(n17422), .Z(n19195) );
  XOR U18715 ( .A(n19197), .B(n19198), .Z(n14312) );
  AND U18716 ( .A(n12422), .B(n17422), .Z(n19197) );
  XNOR U18717 ( .A(n13886), .B(n19199), .Z(n17422) );
  XOR U18718 ( .A(n19200), .B(n17560), .Z(n12422) );
  XOR U18719 ( .A(n3701), .B(n19201), .Z(n18950) );
  XOR U18720 ( .A(n5449), .B(n2135), .Z(n19201) );
  XOR U18721 ( .A(n19202), .B(n9282), .Z(n2135) );
  IV U18722 ( .A(n7175), .Z(n9282) );
  XOR U18723 ( .A(n10110), .B(n14352), .Z(n7175) );
  XOR U18724 ( .A(n19203), .B(n14792), .Z(n14352) );
  NOR U18725 ( .A(n17741), .B(n19204), .Z(n19203) );
  XOR U18726 ( .A(n13312), .B(n12263), .Z(n10110) );
  XOR U18727 ( .A(n19205), .B(n19206), .Z(n12263) );
  XNOR U18728 ( .A(n13275), .B(n13365), .Z(n19206) );
  XOR U18729 ( .A(n19207), .B(n17747), .Z(n13365) );
  IV U18730 ( .A(n14784), .Z(n17747) );
  XOR U18731 ( .A(n19208), .B(n15322), .Z(n14784) );
  ANDN U18732 ( .B(n14363), .A(n14364), .Z(n19207) );
  XNOR U18733 ( .A(n19209), .B(n19210), .Z(n14363) );
  XNOR U18734 ( .A(n19211), .B(n14788), .Z(n13275) );
  XNOR U18735 ( .A(n19150), .B(n19212), .Z(n14788) );
  ANDN U18736 ( .B(n14367), .A(n14368), .Z(n19211) );
  XNOR U18737 ( .A(n19213), .B(n18651), .Z(n14367) );
  XNOR U18738 ( .A(n10805), .B(n19214), .Z(n19205) );
  XOR U18739 ( .A(n14777), .B(n11520), .Z(n19214) );
  XNOR U18740 ( .A(n19215), .B(n17713), .Z(n11520) );
  XNOR U18741 ( .A(n19216), .B(n18637), .Z(n17713) );
  ANDN U18742 ( .B(n14354), .A(n14355), .Z(n19215) );
  XOR U18743 ( .A(n19217), .B(n19218), .Z(n14354) );
  XNOR U18744 ( .A(n19219), .B(n14791), .Z(n14777) );
  AND U18745 ( .A(n19204), .B(n14792), .Z(n19219) );
  XOR U18746 ( .A(n19221), .B(n17491), .Z(n14792) );
  XNOR U18747 ( .A(n19222), .B(n14795), .Z(n10805) );
  XOR U18748 ( .A(n16687), .B(n19223), .Z(n14795) );
  NOR U18749 ( .A(n14360), .B(n14359), .Z(n19222) );
  XOR U18750 ( .A(n17402), .B(n19224), .Z(n14359) );
  IV U18751 ( .A(n19225), .Z(n14360) );
  XOR U18752 ( .A(n19226), .B(n19227), .Z(n13312) );
  XNOR U18753 ( .A(n11991), .B(n15282), .Z(n19227) );
  XOR U18754 ( .A(n19228), .B(n15287), .Z(n15282) );
  IV U18755 ( .A(n17722), .Z(n15287) );
  XOR U18756 ( .A(n17553), .B(n19229), .Z(n17722) );
  ANDN U18757 ( .B(n14389), .A(n14393), .Z(n19228) );
  XNOR U18758 ( .A(n19209), .B(n19230), .Z(n14393) );
  XNOR U18759 ( .A(n16903), .B(n19231), .Z(n14389) );
  XOR U18760 ( .A(n19233), .B(n19234), .Z(n15300) );
  NOR U18761 ( .A(n14373), .B(n14374), .Z(n19232) );
  XNOR U18762 ( .A(n13886), .B(n19235), .Z(n14374) );
  XOR U18763 ( .A(n19236), .B(n15598), .Z(n14373) );
  XOR U18764 ( .A(n19237), .B(n19238), .Z(n15598) );
  XOR U18765 ( .A(n11014), .B(n19239), .Z(n19226) );
  XOR U18766 ( .A(n13420), .B(n11462), .Z(n19239) );
  XOR U18767 ( .A(n19240), .B(n17736), .Z(n11462) );
  IV U18768 ( .A(n15294), .Z(n17736) );
  XNOR U18769 ( .A(n17223), .B(n19241), .Z(n15294) );
  NOR U18770 ( .A(n14388), .B(n14386), .Z(n19240) );
  XOR U18771 ( .A(n19242), .B(n18527), .Z(n14386) );
  XNOR U18772 ( .A(n19243), .B(n19244), .Z(n14388) );
  XNOR U18773 ( .A(n19245), .B(n15297), .Z(n13420) );
  XNOR U18774 ( .A(n16035), .B(n19246), .Z(n15297) );
  ANDN U18775 ( .B(n14377), .A(n14378), .Z(n19245) );
  XNOR U18776 ( .A(n19247), .B(n15827), .Z(n14378) );
  IV U18777 ( .A(n17887), .Z(n15827) );
  XOR U18778 ( .A(n19248), .B(n19249), .Z(n17887) );
  XNOR U18779 ( .A(n19250), .B(n18217), .Z(n14377) );
  XNOR U18780 ( .A(n19251), .B(n15290), .Z(n11014) );
  XNOR U18781 ( .A(n19252), .B(n15626), .Z(n15290) );
  NOR U18782 ( .A(n14383), .B(n14382), .Z(n19251) );
  XNOR U18783 ( .A(n16323), .B(n19253), .Z(n14382) );
  XNOR U18784 ( .A(n17081), .B(n19254), .Z(n14383) );
  IV U18785 ( .A(n18824), .Z(n17081) );
  NOR U18786 ( .A(n6649), .B(n6648), .Z(n19202) );
  XNOR U18787 ( .A(n14040), .B(n10017), .Z(n6648) );
  XNOR U18788 ( .A(n17654), .B(n13158), .Z(n10017) );
  XNOR U18789 ( .A(n19255), .B(n19256), .Z(n13158) );
  XNOR U18790 ( .A(n13647), .B(n12659), .Z(n19256) );
  XNOR U18791 ( .A(n19257), .B(n16437), .Z(n12659) );
  XOR U18792 ( .A(n19258), .B(n18236), .Z(n16437) );
  AND U18793 ( .A(n15494), .B(n15492), .Z(n19257) );
  XOR U18794 ( .A(n15647), .B(n19259), .Z(n15492) );
  XNOR U18795 ( .A(n19260), .B(n17504), .Z(n15494) );
  XNOR U18796 ( .A(n19261), .B(n18927), .Z(n13647) );
  XNOR U18797 ( .A(n19262), .B(n16318), .Z(n18927) );
  IV U18798 ( .A(n19263), .Z(n16318) );
  AND U18799 ( .A(n15496), .B(n15498), .Z(n19261) );
  XNOR U18800 ( .A(n19217), .B(n19264), .Z(n15498) );
  XNOR U18801 ( .A(n19265), .B(n18545), .Z(n15496) );
  XNOR U18802 ( .A(n12737), .B(n19266), .Z(n19255) );
  XNOR U18803 ( .A(n10292), .B(n14603), .Z(n19266) );
  XNOR U18804 ( .A(n19267), .B(n18582), .Z(n14603) );
  XNOR U18805 ( .A(n19268), .B(n14914), .Z(n18582) );
  XNOR U18806 ( .A(n19269), .B(n19270), .Z(n18204) );
  XNOR U18807 ( .A(n18729), .B(n19271), .Z(n19270) );
  XNOR U18808 ( .A(n19272), .B(n19273), .Z(n18729) );
  XOR U18809 ( .A(n17433), .B(n19276), .Z(n19269) );
  XNOR U18810 ( .A(n19277), .B(n19278), .Z(n19276) );
  XNOR U18811 ( .A(n19279), .B(n19280), .Z(n17433) );
  ANDN U18812 ( .B(n19281), .A(n19282), .Z(n19279) );
  ANDN U18813 ( .B(n15503), .A(n15501), .Z(n19267) );
  XOR U18814 ( .A(n19284), .B(n17144), .Z(n15501) );
  XNOR U18815 ( .A(n19285), .B(n17719), .Z(n15503) );
  XNOR U18816 ( .A(n19286), .B(n16434), .Z(n10292) );
  IV U18817 ( .A(n18924), .Z(n16434) );
  XNOR U18818 ( .A(n19287), .B(n17003), .Z(n18924) );
  XNOR U18819 ( .A(n19288), .B(n19289), .Z(n17003) );
  AND U18820 ( .A(n15506), .B(n15505), .Z(n19286) );
  XOR U18821 ( .A(n19290), .B(n19291), .Z(n15505) );
  XNOR U18822 ( .A(n19292), .B(n18725), .Z(n15506) );
  IV U18823 ( .A(n16458), .Z(n18725) );
  XNOR U18824 ( .A(n19293), .B(n16428), .Z(n12737) );
  XOR U18825 ( .A(n19294), .B(n18162), .Z(n16428) );
  ANDN U18826 ( .B(n15511), .A(n15509), .Z(n19293) );
  XNOR U18827 ( .A(n19295), .B(n17415), .Z(n15509) );
  IV U18828 ( .A(n19296), .Z(n17415) );
  XNOR U18829 ( .A(n19297), .B(n17566), .Z(n15511) );
  XOR U18830 ( .A(n19298), .B(n19299), .Z(n17654) );
  XNOR U18831 ( .A(n10780), .B(n18915), .Z(n19299) );
  XOR U18832 ( .A(n19300), .B(n15381), .Z(n18915) );
  XOR U18833 ( .A(n19301), .B(n18355), .Z(n15381) );
  AND U18834 ( .A(n14036), .B(n14038), .Z(n19300) );
  XNOR U18835 ( .A(n15252), .B(n19302), .Z(n14038) );
  XNOR U18836 ( .A(n19303), .B(n16043), .Z(n14036) );
  IV U18837 ( .A(n19291), .Z(n16043) );
  XNOR U18838 ( .A(n19304), .B(n15373), .Z(n10780) );
  XOR U18839 ( .A(n18545), .B(n19305), .Z(n15373) );
  AND U18840 ( .A(n14047), .B(n18949), .Z(n19304) );
  XOR U18841 ( .A(n19306), .B(n17800), .Z(n18949) );
  XNOR U18842 ( .A(n11826), .B(n19308), .Z(n19298) );
  XOR U18843 ( .A(n9577), .B(n18917), .Z(n19308) );
  XOR U18844 ( .A(n19309), .B(n18942), .Z(n18917) );
  XOR U18845 ( .A(n19310), .B(n19311), .Z(n18942) );
  ANDN U18846 ( .B(n18941), .A(n17779), .Z(n19309) );
  XOR U18847 ( .A(n19312), .B(n15388), .Z(n9577) );
  XOR U18848 ( .A(n19313), .B(n19314), .Z(n15388) );
  AND U18849 ( .A(n14542), .B(n18936), .Z(n19312) );
  XOR U18850 ( .A(n19315), .B(n18135), .Z(n18936) );
  XNOR U18851 ( .A(n19316), .B(n17802), .Z(n14542) );
  IV U18852 ( .A(n17121), .Z(n17802) );
  XOR U18853 ( .A(n19317), .B(n18933), .Z(n11826) );
  XOR U18854 ( .A(n19318), .B(n17685), .Z(n18933) );
  IV U18855 ( .A(n18279), .Z(n17685) );
  AND U18856 ( .A(n14042), .B(n14043), .Z(n19317) );
  XOR U18857 ( .A(n19319), .B(n18104), .Z(n14043) );
  IV U18858 ( .A(n18976), .Z(n18104) );
  XNOR U18859 ( .A(n19320), .B(n18162), .Z(n14042) );
  IV U18860 ( .A(n18876), .Z(n18162) );
  XOR U18861 ( .A(n19321), .B(n19322), .Z(n18876) );
  XNOR U18862 ( .A(n19323), .B(n18941), .Z(n14040) );
  XNOR U18863 ( .A(n19324), .B(n16256), .Z(n18941) );
  AND U18864 ( .A(n15376), .B(n17779), .Z(n19323) );
  XNOR U18865 ( .A(n19325), .B(n18462), .Z(n17779) );
  IV U18866 ( .A(n15204), .Z(n18462) );
  XOR U18867 ( .A(n19326), .B(n18473), .Z(n15376) );
  XOR U18868 ( .A(n15715), .B(n10448), .Z(n6649) );
  XOR U18869 ( .A(n13694), .B(n18738), .Z(n10448) );
  XOR U18870 ( .A(n19329), .B(n19330), .Z(n18738) );
  XNOR U18871 ( .A(n14324), .B(n10155), .Z(n19330) );
  XNOR U18872 ( .A(n19331), .B(n15185), .Z(n10155) );
  XOR U18873 ( .A(n19332), .B(n17240), .Z(n15185) );
  IV U18874 ( .A(n17489), .Z(n17240) );
  ANDN U18875 ( .B(n15186), .A(n13799), .Z(n19331) );
  XOR U18876 ( .A(n19333), .B(n19023), .Z(n13799) );
  XOR U18877 ( .A(n19334), .B(n16453), .Z(n15186) );
  XOR U18878 ( .A(n19335), .B(n15193), .Z(n14324) );
  AND U18879 ( .A(n13803), .B(n15192), .Z(n19335) );
  XNOR U18880 ( .A(n17198), .B(n19338), .Z(n15192) );
  XNOR U18881 ( .A(n19339), .B(n17546), .Z(n13803) );
  XOR U18882 ( .A(n11190), .B(n19340), .Z(n19329) );
  XNOR U18883 ( .A(n9095), .B(n12081), .Z(n19340) );
  XNOR U18884 ( .A(n19341), .B(n15195), .Z(n12081) );
  XOR U18885 ( .A(n19342), .B(n17719), .Z(n15195) );
  IV U18886 ( .A(n16047), .Z(n17719) );
  ANDN U18887 ( .B(n15720), .A(n13790), .Z(n19341) );
  XNOR U18888 ( .A(n19345), .B(n18759), .Z(n13790) );
  XOR U18889 ( .A(n19346), .B(n19296), .Z(n15720) );
  XOR U18890 ( .A(n19347), .B(n17381), .Z(n9095) );
  XNOR U18891 ( .A(n19348), .B(n17039), .Z(n17381) );
  ANDN U18892 ( .B(n15722), .A(n13794), .Z(n19347) );
  XNOR U18893 ( .A(n19349), .B(n19350), .Z(n13794) );
  XNOR U18894 ( .A(n19209), .B(n19351), .Z(n15722) );
  IV U18895 ( .A(n18743), .Z(n19209) );
  XOR U18896 ( .A(n18175), .B(n19352), .Z(n18743) );
  XOR U18897 ( .A(n19353), .B(n19354), .Z(n18175) );
  XNOR U18898 ( .A(n16466), .B(n14923), .Z(n19354) );
  XNOR U18899 ( .A(n19355), .B(n19356), .Z(n14923) );
  NOR U18900 ( .A(n19357), .B(n19358), .Z(n19355) );
  XNOR U18901 ( .A(n19359), .B(n19360), .Z(n16466) );
  XNOR U18902 ( .A(n18286), .B(n19363), .Z(n19353) );
  XOR U18903 ( .A(n18326), .B(n19364), .Z(n19363) );
  XOR U18904 ( .A(n19365), .B(n19366), .Z(n18326) );
  AND U18905 ( .A(n19367), .B(n19368), .Z(n19365) );
  XNOR U18906 ( .A(n19369), .B(n19370), .Z(n18286) );
  AND U18907 ( .A(n19371), .B(n19372), .Z(n19369) );
  XNOR U18908 ( .A(n19373), .B(n15189), .Z(n11190) );
  XNOR U18909 ( .A(n19374), .B(n17522), .Z(n15189) );
  XOR U18910 ( .A(n19375), .B(n19376), .Z(n13694) );
  XNOR U18911 ( .A(n13552), .B(n11830), .Z(n19376) );
  XOR U18912 ( .A(n19377), .B(n14333), .Z(n11830) );
  XOR U18913 ( .A(n19378), .B(n19337), .Z(n14333) );
  NOR U18914 ( .A(n13059), .B(n13061), .Z(n19377) );
  XNOR U18915 ( .A(n19379), .B(n16672), .Z(n13061) );
  XOR U18916 ( .A(n19380), .B(n17186), .Z(n13059) );
  XNOR U18917 ( .A(n19381), .B(n14338), .Z(n13552) );
  XOR U18918 ( .A(n19382), .B(n18130), .Z(n14338) );
  NOR U18919 ( .A(n13693), .B(n13691), .Z(n19381) );
  XNOR U18920 ( .A(n19383), .B(n18399), .Z(n13691) );
  IV U18921 ( .A(n17058), .Z(n13693) );
  XOR U18922 ( .A(n19384), .B(n19029), .Z(n17058) );
  IV U18923 ( .A(n18254), .Z(n19029) );
  XNOR U18924 ( .A(n12875), .B(n19385), .Z(n19375) );
  XNOR U18925 ( .A(n12850), .B(n10902), .Z(n19385) );
  XNOR U18926 ( .A(n19386), .B(n14330), .Z(n10902) );
  XOR U18927 ( .A(n19387), .B(n16746), .Z(n14330) );
  NOR U18928 ( .A(n13064), .B(n13063), .Z(n19386) );
  XNOR U18929 ( .A(n19388), .B(n17441), .Z(n13063) );
  XNOR U18930 ( .A(n19389), .B(n16767), .Z(n13064) );
  XNOR U18931 ( .A(n19390), .B(n15725), .Z(n12850) );
  XOR U18932 ( .A(n19391), .B(n17555), .Z(n15725) );
  AND U18933 ( .A(n13056), .B(n13054), .Z(n19390) );
  XNOR U18934 ( .A(n19392), .B(n18119), .Z(n13054) );
  XOR U18935 ( .A(n19393), .B(n17042), .Z(n13056) );
  XNOR U18936 ( .A(n19394), .B(n14341), .Z(n12875) );
  XNOR U18937 ( .A(n19395), .B(n16944), .Z(n14341) );
  ANDN U18938 ( .B(n13067), .A(n13068), .Z(n19394) );
  XNOR U18939 ( .A(n19396), .B(n16808), .Z(n13068) );
  XNOR U18940 ( .A(n18044), .B(n19397), .Z(n13067) );
  XNOR U18941 ( .A(n19398), .B(n15190), .Z(n15715) );
  XOR U18942 ( .A(n19399), .B(n19400), .Z(n15190) );
  ANDN U18943 ( .B(n17392), .A(n13807), .Z(n19398) );
  XOR U18944 ( .A(n17959), .B(n19401), .Z(n13807) );
  IV U18945 ( .A(n13809), .Z(n17392) );
  XOR U18946 ( .A(n19402), .B(n19403), .Z(n13809) );
  XOR U18947 ( .A(n19404), .B(n9404), .Z(n5449) );
  IV U18948 ( .A(n9285), .Z(n9404) );
  XNOR U18949 ( .A(n15107), .B(n9388), .Z(n9285) );
  XOR U18950 ( .A(n19405), .B(n19406), .Z(n14642) );
  XOR U18951 ( .A(n9528), .B(n9998), .Z(n19406) );
  XOR U18952 ( .A(n19407), .B(n16637), .Z(n9998) );
  ANDN U18953 ( .B(n15101), .A(n15099), .Z(n19407) );
  XOR U18954 ( .A(n19408), .B(n16630), .Z(n9528) );
  AND U18955 ( .A(n15105), .B(n19409), .Z(n19408) );
  XOR U18956 ( .A(n19410), .B(n19411), .Z(n19405) );
  XOR U18957 ( .A(n12987), .B(n12841), .Z(n19411) );
  XNOR U18958 ( .A(n19412), .B(n16624), .Z(n12841) );
  AND U18959 ( .A(n15111), .B(n19413), .Z(n19412) );
  XOR U18960 ( .A(n19414), .B(n16635), .Z(n12987) );
  IV U18961 ( .A(n19415), .Z(n16635) );
  NOR U18962 ( .A(n19416), .B(n19417), .Z(n19414) );
  XNOR U18963 ( .A(n19418), .B(n19419), .Z(n17662) );
  XNOR U18964 ( .A(n12575), .B(n9809), .Z(n19419) );
  XOR U18965 ( .A(n19420), .B(n19421), .Z(n9809) );
  ANDN U18966 ( .B(n14971), .A(n13435), .Z(n19420) );
  XOR U18967 ( .A(n19422), .B(n17035), .Z(n13435) );
  IV U18968 ( .A(n19423), .Z(n17035) );
  XOR U18969 ( .A(n19424), .B(n16619), .Z(n12575) );
  AND U18970 ( .A(n14439), .B(n14967), .Z(n19424) );
  XOR U18971 ( .A(n19425), .B(n16555), .Z(n14439) );
  XNOR U18972 ( .A(n16128), .B(n19426), .Z(n19418) );
  XOR U18973 ( .A(n16498), .B(n9939), .Z(n19426) );
  XOR U18974 ( .A(n19427), .B(n16616), .Z(n9939) );
  ANDN U18975 ( .B(n17659), .A(n13439), .Z(n19427) );
  XNOR U18976 ( .A(n17680), .B(n19428), .Z(n13439) );
  XOR U18977 ( .A(n19429), .B(n16614), .Z(n16498) );
  ANDN U18978 ( .B(n14965), .A(n14826), .Z(n19429) );
  XNOR U18979 ( .A(n19430), .B(n16779), .Z(n14826) );
  XNOR U18980 ( .A(n19431), .B(n16604), .Z(n16128) );
  ANDN U18981 ( .B(n13429), .A(n14973), .Z(n19431) );
  XOR U18982 ( .A(n19432), .B(n16039), .Z(n13429) );
  XNOR U18983 ( .A(n19433), .B(n19416), .Z(n15107) );
  ANDN U18984 ( .B(n19417), .A(n16633), .Z(n19433) );
  NOR U18985 ( .A(n6653), .B(n6652), .Z(n19404) );
  XNOR U18986 ( .A(n9399), .B(n14987), .Z(n6652) );
  XOR U18987 ( .A(n19434), .B(n16146), .Z(n14987) );
  AND U18988 ( .A(n18086), .B(n19435), .Z(n19434) );
  XOR U18989 ( .A(n19436), .B(n17186), .Z(n18086) );
  IV U18990 ( .A(n11562), .Z(n9399) );
  XNOR U18991 ( .A(n13398), .B(n15863), .Z(n11562) );
  XNOR U18992 ( .A(n19437), .B(n19438), .Z(n15863) );
  XNOR U18993 ( .A(n14536), .B(n15747), .Z(n19438) );
  XOR U18994 ( .A(n19439), .B(n16138), .Z(n15747) );
  XNOR U18995 ( .A(n19440), .B(n19441), .Z(n16138) );
  NOR U18996 ( .A(n14995), .B(n14993), .Z(n19439) );
  XNOR U18997 ( .A(n19442), .B(n19443), .Z(n14993) );
  XOR U18998 ( .A(n19444), .B(n19403), .Z(n14995) );
  XNOR U18999 ( .A(n19445), .B(n16142), .Z(n14536) );
  XNOR U19000 ( .A(n19446), .B(n16100), .Z(n16142) );
  ANDN U19001 ( .B(n14979), .A(n14980), .Z(n19445) );
  XOR U19002 ( .A(n18245), .B(n19447), .Z(n14980) );
  IV U19003 ( .A(n17914), .Z(n18245) );
  XNOR U19004 ( .A(n19448), .B(n16031), .Z(n14979) );
  XOR U19005 ( .A(n11447), .B(n19449), .Z(n19437) );
  XOR U19006 ( .A(n11319), .B(n16129), .Z(n19449) );
  XNOR U19007 ( .A(n19450), .B(n16145), .Z(n16129) );
  XNOR U19008 ( .A(n15917), .B(n19451), .Z(n16145) );
  AND U19009 ( .A(n16146), .B(n19082), .Z(n19450) );
  IV U19010 ( .A(n19435), .Z(n19082) );
  XOR U19011 ( .A(n19452), .B(n19291), .Z(n19435) );
  XNOR U19012 ( .A(n16543), .B(n19453), .Z(n16146) );
  XOR U19013 ( .A(n19454), .B(n16149), .Z(n11319) );
  XOR U19014 ( .A(n19455), .B(n16812), .Z(n16149) );
  IV U19015 ( .A(n17732), .Z(n16812) );
  XOR U19016 ( .A(n19456), .B(n19457), .Z(n17732) );
  ANDN U19017 ( .B(n14985), .A(n14983), .Z(n19454) );
  XOR U19018 ( .A(n18545), .B(n19458), .Z(n14983) );
  XNOR U19019 ( .A(n19459), .B(n18616), .Z(n14985) );
  IV U19020 ( .A(n16788), .Z(n18616) );
  XNOR U19021 ( .A(n19460), .B(n16135), .Z(n11447) );
  XNOR U19022 ( .A(n19461), .B(n17683), .Z(n16135) );
  NOR U19023 ( .A(n14989), .B(n14990), .Z(n19460) );
  XNOR U19024 ( .A(n14904), .B(n19462), .Z(n14990) );
  IV U19025 ( .A(n16796), .Z(n14904) );
  XOR U19026 ( .A(n19463), .B(n18979), .Z(n16796) );
  XOR U19027 ( .A(n19464), .B(n19465), .Z(n18979) );
  XNOR U19028 ( .A(n19466), .B(n18187), .Z(n19465) );
  XOR U19029 ( .A(n19467), .B(n19468), .Z(n18187) );
  ANDN U19030 ( .B(n19469), .A(n19470), .Z(n19467) );
  XOR U19031 ( .A(n19471), .B(n19472), .Z(n19464) );
  XOR U19032 ( .A(n15519), .B(n18112), .Z(n19472) );
  XOR U19033 ( .A(n19473), .B(n19474), .Z(n18112) );
  ANDN U19034 ( .B(n19475), .A(n19476), .Z(n19473) );
  XOR U19035 ( .A(n19477), .B(n19478), .Z(n15519) );
  ANDN U19036 ( .B(n19479), .A(n19480), .Z(n19477) );
  XNOR U19037 ( .A(n19481), .B(n18180), .Z(n14989) );
  XOR U19038 ( .A(n19482), .B(n19483), .Z(n13398) );
  XOR U19039 ( .A(n18340), .B(n11669), .Z(n19483) );
  XOR U19040 ( .A(n19484), .B(n14776), .Z(n11669) );
  XOR U19041 ( .A(n19485), .B(n18434), .Z(n14776) );
  NOR U19042 ( .A(n15565), .B(n15566), .Z(n19484) );
  XNOR U19043 ( .A(n17258), .B(n19486), .Z(n15566) );
  XNOR U19044 ( .A(n19487), .B(n17474), .Z(n15565) );
  XNOR U19045 ( .A(n19488), .B(n15811), .Z(n18340) );
  XOR U19046 ( .A(n18044), .B(n19489), .Z(n15811) );
  NOR U19047 ( .A(n15555), .B(n15554), .Z(n19488) );
  XNOR U19048 ( .A(n19490), .B(n19491), .Z(n15554) );
  XNOR U19049 ( .A(n19492), .B(n15217), .Z(n15555) );
  XOR U19050 ( .A(n10138), .B(n19493), .Z(n19482) );
  XOR U19051 ( .A(n11770), .B(n11822), .Z(n19493) );
  XNOR U19052 ( .A(n19494), .B(n14768), .Z(n11822) );
  XNOR U19053 ( .A(n19495), .B(n16460), .Z(n14768) );
  IV U19054 ( .A(n19156), .Z(n16460) );
  AND U19055 ( .A(n15562), .B(n15563), .Z(n19494) );
  XOR U19056 ( .A(n19496), .B(n18306), .Z(n15563) );
  XNOR U19057 ( .A(n18824), .B(n19497), .Z(n15562) );
  XOR U19058 ( .A(n19500), .B(n16363), .Z(n11770) );
  XOR U19059 ( .A(n17553), .B(n19501), .Z(n16363) );
  NOR U19060 ( .A(n15551), .B(n15550), .Z(n19500) );
  XNOR U19061 ( .A(n19502), .B(n19503), .Z(n15550) );
  XNOR U19062 ( .A(n19504), .B(n17517), .Z(n15551) );
  XNOR U19063 ( .A(n19505), .B(n19506), .Z(n18452) );
  XNOR U19064 ( .A(n18639), .B(n17660), .Z(n19506) );
  XOR U19065 ( .A(n19507), .B(n19508), .Z(n17660) );
  ANDN U19066 ( .B(n19509), .A(n19510), .Z(n19507) );
  XNOR U19067 ( .A(n19511), .B(n19512), .Z(n18639) );
  NOR U19068 ( .A(n19513), .B(n19514), .Z(n19511) );
  XOR U19069 ( .A(n16455), .B(n19515), .Z(n19505) );
  XOR U19070 ( .A(n18883), .B(n17669), .Z(n19515) );
  XNOR U19071 ( .A(n19516), .B(n19517), .Z(n17669) );
  ANDN U19072 ( .B(n19518), .A(n19519), .Z(n19516) );
  XNOR U19073 ( .A(n19520), .B(n19521), .Z(n18883) );
  ANDN U19074 ( .B(n19522), .A(n19523), .Z(n19520) );
  XNOR U19075 ( .A(n19524), .B(n19525), .Z(n16455) );
  ANDN U19076 ( .B(n19526), .A(n19527), .Z(n19524) );
  XNOR U19077 ( .A(n19529), .B(n14765), .Z(n10138) );
  XNOR U19078 ( .A(n17965), .B(n19530), .Z(n14765) );
  AND U19079 ( .A(n15559), .B(n16347), .Z(n19529) );
  IV U19080 ( .A(n15560), .Z(n16347) );
  XNOR U19081 ( .A(n19531), .B(n18759), .Z(n15560) );
  XNOR U19082 ( .A(n19532), .B(n17509), .Z(n15559) );
  XNOR U19083 ( .A(n17536), .B(n10008), .Z(n6653) );
  XNOR U19084 ( .A(n19533), .B(n13934), .Z(n17536) );
  ANDN U19085 ( .B(n19534), .A(n13105), .Z(n19533) );
  XNOR U19086 ( .A(n19535), .B(n19291), .Z(n13105) );
  XOR U19087 ( .A(n19538), .B(n7166), .Z(n3701) );
  IV U19088 ( .A(n9289), .Z(n7166) );
  XOR U19089 ( .A(n17695), .B(n11793), .Z(n9289) );
  XNOR U19090 ( .A(n11852), .B(n11865), .Z(n11793) );
  XNOR U19091 ( .A(n19539), .B(n19540), .Z(n11865) );
  XOR U19092 ( .A(n10945), .B(n11642), .Z(n19540) );
  XOR U19093 ( .A(n19541), .B(n16491), .Z(n11642) );
  NOR U19094 ( .A(n14735), .B(n16490), .Z(n19541) );
  XNOR U19095 ( .A(n19542), .B(n19314), .Z(n16490) );
  XNOR U19096 ( .A(n19543), .B(n19544), .Z(n14735) );
  XNOR U19097 ( .A(n19545), .B(n16513), .Z(n10945) );
  NOR U19098 ( .A(n16512), .B(n14727), .Z(n19545) );
  XNOR U19099 ( .A(n16663), .B(n19546), .Z(n14727) );
  XNOR U19100 ( .A(n15592), .B(n19547), .Z(n16512) );
  XOR U19101 ( .A(n10690), .B(n19548), .Z(n19539) );
  XOR U19102 ( .A(n16125), .B(n11804), .Z(n19548) );
  XOR U19103 ( .A(n19549), .B(n18413), .Z(n11804) );
  NOR U19104 ( .A(n14731), .B(n17709), .Z(n19549) );
  XOR U19105 ( .A(n19550), .B(n17589), .Z(n17709) );
  XNOR U19106 ( .A(n19551), .B(n16519), .Z(n14731) );
  XNOR U19107 ( .A(n19552), .B(n16486), .Z(n16125) );
  ANDN U19108 ( .B(n14718), .A(n16485), .Z(n19552) );
  XNOR U19109 ( .A(n19553), .B(n18879), .Z(n16485) );
  XNOR U19110 ( .A(n15252), .B(n19554), .Z(n14718) );
  XOR U19111 ( .A(n19555), .B(n19556), .Z(n10690) );
  NOR U19112 ( .A(n14722), .B(n16493), .Z(n19555) );
  XNOR U19113 ( .A(n19557), .B(n19558), .Z(n16493) );
  XNOR U19114 ( .A(n19559), .B(n15843), .Z(n14722) );
  XNOR U19115 ( .A(n18563), .B(n19560), .Z(n15843) );
  XOR U19116 ( .A(n19561), .B(n19562), .Z(n18563) );
  XOR U19117 ( .A(n19324), .B(n19563), .Z(n19562) );
  XNOR U19118 ( .A(n19564), .B(n19565), .Z(n19324) );
  AND U19119 ( .A(n19566), .B(n19567), .Z(n19564) );
  XOR U19120 ( .A(n19568), .B(n19569), .Z(n19561) );
  XOR U19121 ( .A(n16255), .B(n19570), .Z(n19569) );
  XNOR U19122 ( .A(n19571), .B(n19572), .Z(n16255) );
  ANDN U19123 ( .B(n19573), .A(n19574), .Z(n19571) );
  XOR U19124 ( .A(n19575), .B(n19576), .Z(n11852) );
  XNOR U19125 ( .A(n16479), .B(n14154), .Z(n19576) );
  XNOR U19126 ( .A(n19577), .B(n17319), .Z(n14154) );
  NOR U19127 ( .A(n17320), .B(n17697), .Z(n19577) );
  XOR U19128 ( .A(n19578), .B(n18707), .Z(n17320) );
  XNOR U19129 ( .A(n19579), .B(n17315), .Z(n16479) );
  ANDN U19130 ( .B(n17316), .A(n17692), .Z(n19579) );
  XNOR U19131 ( .A(n19580), .B(n16414), .Z(n17316) );
  XOR U19132 ( .A(n12352), .B(n19581), .Z(n19575) );
  XOR U19133 ( .A(n13310), .B(n12068), .Z(n19581) );
  XOR U19134 ( .A(n19582), .B(n19583), .Z(n12068) );
  NOR U19135 ( .A(n17306), .B(n19584), .Z(n19582) );
  XOR U19136 ( .A(n19585), .B(n19586), .Z(n13310) );
  NOR U19137 ( .A(n18229), .B(n18230), .Z(n19585) );
  XNOR U19138 ( .A(n19587), .B(n17311), .Z(n12352) );
  AND U19139 ( .A(n17312), .B(n17701), .Z(n19587) );
  XOR U19140 ( .A(n19588), .B(n17564), .Z(n17312) );
  XNOR U19141 ( .A(n19589), .B(n17306), .Z(n17695) );
  XNOR U19142 ( .A(n19590), .B(n19023), .Z(n17306) );
  ANDN U19143 ( .B(n19584), .A(n19591), .Z(n19589) );
  XNOR U19144 ( .A(n13401), .B(n9119), .Z(n6643) );
  XOR U19145 ( .A(n14008), .B(n18341), .Z(n9119) );
  XOR U19146 ( .A(n19592), .B(n19593), .Z(n18341) );
  XNOR U19147 ( .A(n12169), .B(n12840), .Z(n19593) );
  XNOR U19148 ( .A(n19594), .B(n14098), .Z(n12840) );
  XNOR U19149 ( .A(n19595), .B(n19544), .Z(n14098) );
  ANDN U19150 ( .B(n15578), .A(n13405), .Z(n19594) );
  XOR U19151 ( .A(n19596), .B(n19597), .Z(n13405) );
  XOR U19152 ( .A(n19598), .B(n18458), .Z(n15578) );
  XOR U19153 ( .A(n19599), .B(n16341), .Z(n12169) );
  IV U19154 ( .A(n14102), .Z(n16341) );
  XOR U19155 ( .A(n19600), .B(n15217), .Z(n14102) );
  NOR U19156 ( .A(n14101), .B(n14255), .Z(n19599) );
  XNOR U19157 ( .A(n18217), .B(n19601), .Z(n14255) );
  XNOR U19158 ( .A(n19602), .B(n19337), .Z(n14101) );
  XOR U19159 ( .A(n10990), .B(n19603), .Z(n19592) );
  XOR U19160 ( .A(n14080), .B(n12859), .Z(n19603) );
  XOR U19161 ( .A(n19604), .B(n16335), .Z(n12859) );
  IV U19162 ( .A(n14086), .Z(n16335) );
  XOR U19163 ( .A(n19605), .B(n18236), .Z(n14086) );
  ANDN U19164 ( .B(n14087), .A(n13414), .Z(n19604) );
  XNOR U19165 ( .A(n19606), .B(n16453), .Z(n13414) );
  XOR U19166 ( .A(n19607), .B(n19608), .Z(n16453) );
  XOR U19167 ( .A(n19609), .B(n18609), .Z(n14087) );
  XOR U19168 ( .A(n18637), .B(n19611), .Z(n14090) );
  NOR U19169 ( .A(n13410), .B(n13409), .Z(n19610) );
  XOR U19170 ( .A(n19612), .B(n19613), .Z(n13409) );
  XOR U19171 ( .A(n19614), .B(n17474), .Z(n13410) );
  XOR U19172 ( .A(n19615), .B(n19616), .Z(n17474) );
  XNOR U19173 ( .A(n19617), .B(n14094), .Z(n10990) );
  XNOR U19174 ( .A(n19618), .B(n17869), .Z(n14094) );
  NOR U19175 ( .A(n15572), .B(n14095), .Z(n19617) );
  XOR U19176 ( .A(n19619), .B(n19620), .Z(n14008) );
  XNOR U19177 ( .A(n19039), .B(n12043), .Z(n19620) );
  XOR U19178 ( .A(n19621), .B(n15087), .Z(n12043) );
  XNOR U19179 ( .A(n19622), .B(n16557), .Z(n17156) );
  XOR U19180 ( .A(n19623), .B(n15095), .Z(n19039) );
  ANDN U19181 ( .B(n17161), .A(n14656), .Z(n19623) );
  XNOR U19182 ( .A(n19624), .B(n16919), .Z(n14656) );
  IV U19183 ( .A(n15597), .Z(n16919) );
  XOR U19184 ( .A(n12644), .B(n19627), .Z(n19619) );
  XOR U19185 ( .A(n19628), .B(n11874), .Z(n19627) );
  XOR U19186 ( .A(n19629), .B(n15090), .Z(n11874) );
  ANDN U19187 ( .B(n17173), .A(n14646), .Z(n19629) );
  XOR U19188 ( .A(n19630), .B(n17441), .Z(n14646) );
  IV U19189 ( .A(n17847), .Z(n17441) );
  XNOR U19190 ( .A(n19631), .B(n19632), .Z(n17847) );
  XNOR U19191 ( .A(n19633), .B(n15083), .Z(n12644) );
  ANDN U19192 ( .B(n19634), .A(n14660), .Z(n19633) );
  XNOR U19193 ( .A(n19638), .B(n14095), .Z(n13401) );
  XNOR U19194 ( .A(n19639), .B(n17144), .Z(n14095) );
  XOR U19195 ( .A(n19640), .B(n18884), .Z(n17144) );
  XOR U19196 ( .A(n19641), .B(n19642), .Z(n18884) );
  XOR U19197 ( .A(n19596), .B(n19643), .Z(n19642) );
  XNOR U19198 ( .A(n19644), .B(n19645), .Z(n19596) );
  ANDN U19199 ( .B(n19508), .A(n19509), .Z(n19644) );
  XOR U19200 ( .A(n19646), .B(n19647), .Z(n19641) );
  XOR U19201 ( .A(n19490), .B(n19648), .Z(n19647) );
  XNOR U19202 ( .A(n19649), .B(n19650), .Z(n19490) );
  ANDN U19203 ( .B(n19517), .A(n19518), .Z(n19649) );
  ANDN U19204 ( .B(n15572), .A(n15573), .Z(n19638) );
  XNOR U19205 ( .A(n19651), .B(n18130), .Z(n15573) );
  IV U19206 ( .A(n17149), .Z(n18130) );
  XOR U19207 ( .A(n19652), .B(n19653), .Z(n17149) );
  XNOR U19208 ( .A(n17965), .B(n19654), .Z(n15572) );
  XOR U19209 ( .A(n15153), .B(n11859), .Z(n6644) );
  XOR U19210 ( .A(n19655), .B(n14579), .Z(n15153) );
  XOR U19211 ( .A(n19656), .B(n16519), .Z(n16439) );
  IV U19212 ( .A(n19657), .Z(n16519) );
  XOR U19213 ( .A(n19658), .B(n19659), .Z(n6580) );
  XNOR U19214 ( .A(n4868), .B(n4039), .Z(n19659) );
  XOR U19215 ( .A(n19660), .B(n6618), .Z(n4039) );
  IV U19216 ( .A(n9266), .Z(n6618) );
  XNOR U19217 ( .A(n15890), .B(n10783), .Z(n9266) );
  XNOR U19218 ( .A(n14431), .B(n12201), .Z(n10783) );
  XNOR U19219 ( .A(n19661), .B(n19662), .Z(n12201) );
  XNOR U19220 ( .A(n10210), .B(n11540), .Z(n19662) );
  XNOR U19221 ( .A(n19663), .B(n13137), .Z(n11540) );
  XOR U19222 ( .A(n19664), .B(n19665), .Z(n13137) );
  ANDN U19223 ( .B(n13138), .A(n13622), .Z(n19663) );
  XOR U19224 ( .A(n19666), .B(n17075), .Z(n13622) );
  XOR U19225 ( .A(n19667), .B(n19558), .Z(n13138) );
  XNOR U19226 ( .A(n19668), .B(n13150), .Z(n10210) );
  XNOR U19227 ( .A(n19669), .B(n16795), .Z(n13150) );
  XOR U19228 ( .A(n19670), .B(n19671), .Z(n16795) );
  ANDN U19229 ( .B(n13151), .A(n13619), .Z(n19668) );
  XNOR U19230 ( .A(n9174), .B(n19672), .Z(n19661) );
  XOR U19231 ( .A(n9117), .B(n11392), .Z(n19672) );
  XOR U19232 ( .A(n19673), .B(n13142), .Z(n11392) );
  XOR U19233 ( .A(n18773), .B(n14918), .Z(n13142) );
  XOR U19234 ( .A(n19674), .B(n19675), .Z(n18773) );
  ANDN U19235 ( .B(n19676), .A(n19677), .Z(n19674) );
  AND U19236 ( .A(n14012), .B(n13143), .Z(n19673) );
  XOR U19237 ( .A(n19678), .B(n19423), .Z(n13143) );
  XOR U19238 ( .A(n19679), .B(n17167), .Z(n14012) );
  XNOR U19239 ( .A(n19680), .B(n19681), .Z(n17167) );
  XNOR U19240 ( .A(n19682), .B(n13147), .Z(n9117) );
  XOR U19241 ( .A(n19683), .B(n16672), .Z(n13147) );
  ANDN U19242 ( .B(n13146), .A(n13614), .Z(n19682) );
  XOR U19243 ( .A(n19684), .B(n19685), .Z(n13614) );
  IV U19244 ( .A(n15896), .Z(n13146) );
  XOR U19245 ( .A(n19687), .B(n17955), .Z(n9174) );
  XOR U19246 ( .A(n19096), .B(n18505), .Z(n17955) );
  XNOR U19247 ( .A(n19690), .B(n19691), .Z(n19096) );
  ANDN U19248 ( .B(n19692), .A(n19693), .Z(n19690) );
  AND U19249 ( .A(n15898), .B(n13995), .Z(n19687) );
  XNOR U19250 ( .A(n17332), .B(n19694), .Z(n13995) );
  XOR U19251 ( .A(n19695), .B(n19696), .Z(n15898) );
  XOR U19252 ( .A(n19697), .B(n19698), .Z(n14431) );
  XNOR U19253 ( .A(n14567), .B(n12180), .Z(n19698) );
  XNOR U19254 ( .A(n19699), .B(n14599), .Z(n12180) );
  XNOR U19255 ( .A(n16663), .B(n19700), .Z(n14599) );
  ANDN U19256 ( .B(n14025), .A(n13640), .Z(n19699) );
  XNOR U19257 ( .A(n17914), .B(n19701), .Z(n13640) );
  XOR U19258 ( .A(n19702), .B(n19703), .Z(n14025) );
  XNOR U19259 ( .A(n19704), .B(n14592), .Z(n14567) );
  XNOR U19260 ( .A(n19705), .B(n18015), .Z(n14592) );
  IV U19261 ( .A(n19187), .Z(n18015) );
  AND U19262 ( .A(n14433), .B(n13636), .Z(n19704) );
  XOR U19263 ( .A(n16543), .B(n19706), .Z(n13636) );
  XOR U19264 ( .A(n19709), .B(n16343), .Z(n14433) );
  XOR U19265 ( .A(n14538), .B(n19710), .Z(n19697) );
  XNOR U19266 ( .A(n11444), .B(n10942), .Z(n19710) );
  XNOR U19267 ( .A(n19711), .B(n14597), .Z(n10942) );
  XOR U19268 ( .A(n19712), .B(n16830), .Z(n14597) );
  ANDN U19269 ( .B(n14019), .A(n13631), .Z(n19711) );
  XNOR U19270 ( .A(n19713), .B(n15129), .Z(n13631) );
  XNOR U19271 ( .A(n19715), .B(n14594), .Z(n11444) );
  XOR U19272 ( .A(n17397), .B(n19716), .Z(n14594) );
  IV U19273 ( .A(n15974), .Z(n17397) );
  XOR U19274 ( .A(n19717), .B(n19718), .Z(n15974) );
  AND U19275 ( .A(n14022), .B(n13644), .Z(n19715) );
  IV U19276 ( .A(n14023), .Z(n13644) );
  XOR U19277 ( .A(n16783), .B(n19719), .Z(n14023) );
  IV U19278 ( .A(n17965), .Z(n16783) );
  XNOR U19279 ( .A(n19139), .B(n19720), .Z(n17965) );
  XOR U19280 ( .A(n19721), .B(n19722), .Z(n19139) );
  XNOR U19281 ( .A(n19723), .B(n19724), .Z(n19722) );
  XOR U19282 ( .A(n19725), .B(n19726), .Z(n19721) );
  XOR U19283 ( .A(n19727), .B(n17811), .Z(n19726) );
  XNOR U19284 ( .A(n19728), .B(n19729), .Z(n17811) );
  XOR U19285 ( .A(n19731), .B(n19732), .Z(n14022) );
  XNOR U19286 ( .A(n19733), .B(n14601), .Z(n14538) );
  XOR U19287 ( .A(n18046), .B(n19734), .Z(n14601) );
  AND U19288 ( .A(n14028), .B(n13627), .Z(n19733) );
  XOR U19289 ( .A(n19735), .B(n18121), .Z(n13627) );
  XOR U19290 ( .A(n19058), .B(n19736), .Z(n14028) );
  IV U19291 ( .A(n15958), .Z(n19058) );
  XOR U19292 ( .A(n19737), .B(n19738), .Z(n15958) );
  XNOR U19293 ( .A(n19739), .B(n13151), .Z(n15890) );
  XOR U19294 ( .A(n19740), .B(n15249), .Z(n13151) );
  IV U19295 ( .A(n19741), .Z(n15249) );
  AND U19296 ( .A(n13619), .B(n17969), .Z(n19739) );
  IV U19297 ( .A(n13620), .Z(n17969) );
  XOR U19298 ( .A(n14944), .B(n19742), .Z(n13620) );
  XOR U19299 ( .A(n19743), .B(n19744), .Z(n14944) );
  XOR U19300 ( .A(n19745), .B(n17489), .Z(n13619) );
  XNOR U19301 ( .A(n19746), .B(n19747), .Z(n19016) );
  XNOR U19302 ( .A(n15586), .B(n15528), .Z(n19747) );
  XOR U19303 ( .A(n19748), .B(n19749), .Z(n15528) );
  ANDN U19304 ( .B(n19750), .A(n19751), .Z(n19748) );
  XOR U19305 ( .A(n19752), .B(n19753), .Z(n15586) );
  ANDN U19306 ( .B(n19754), .A(n19755), .Z(n19752) );
  XOR U19307 ( .A(n16449), .B(n19756), .Z(n19746) );
  XOR U19308 ( .A(n16095), .B(n18630), .Z(n19756) );
  XOR U19309 ( .A(n19757), .B(n19758), .Z(n18630) );
  ANDN U19310 ( .B(n19759), .A(n19760), .Z(n19757) );
  XOR U19311 ( .A(n19761), .B(n19762), .Z(n16095) );
  XNOR U19312 ( .A(n19765), .B(n19766), .Z(n16449) );
  NOR U19313 ( .A(n19767), .B(n19768), .Z(n19765) );
  ANDN U19314 ( .B(n9211), .A(n7078), .Z(n19660) );
  XNOR U19315 ( .A(n16967), .B(n9917), .Z(n7078) );
  XNOR U19316 ( .A(n18197), .B(n11850), .Z(n9917) );
  XNOR U19317 ( .A(n19770), .B(n19771), .Z(n11850) );
  XNOR U19318 ( .A(n15700), .B(n11507), .Z(n19771) );
  XOR U19319 ( .A(n19772), .B(n17701), .Z(n11507) );
  XOR U19320 ( .A(n19773), .B(n17857), .Z(n17701) );
  IV U19321 ( .A(n18011), .Z(n17857) );
  XOR U19322 ( .A(n19774), .B(n19775), .Z(n18011) );
  XNOR U19323 ( .A(n19776), .B(n19584), .Z(n15700) );
  XOR U19324 ( .A(n16758), .B(n19777), .Z(n19584) );
  ANDN U19325 ( .B(n19591), .A(n17305), .Z(n19776) );
  XOR U19326 ( .A(n10993), .B(n19778), .Z(n19770) );
  XOR U19327 ( .A(n10831), .B(n17687), .Z(n19778) );
  XOR U19328 ( .A(n19779), .B(n17692), .Z(n17687) );
  XNOR U19329 ( .A(n19780), .B(n18368), .Z(n17692) );
  AND U19330 ( .A(n17693), .B(n19781), .Z(n19779) );
  XOR U19331 ( .A(n19782), .B(n17697), .Z(n10831) );
  XNOR U19332 ( .A(n19783), .B(n16672), .Z(n17697) );
  XNOR U19333 ( .A(n19784), .B(n19785), .Z(n16672) );
  ANDN U19334 ( .B(n17698), .A(n17318), .Z(n19782) );
  XNOR U19335 ( .A(n19786), .B(n18230), .Z(n10993) );
  XNOR U19336 ( .A(n19563), .B(n19787), .Z(n18230) );
  XOR U19337 ( .A(n19788), .B(n19789), .Z(n19563) );
  NOR U19338 ( .A(n19790), .B(n19791), .Z(n19788) );
  XOR U19339 ( .A(n19793), .B(n19794), .Z(n18197) );
  XOR U19340 ( .A(n14545), .B(n13469), .Z(n19794) );
  XOR U19341 ( .A(n19795), .B(n13710), .Z(n13469) );
  XNOR U19342 ( .A(n17972), .B(n19796), .Z(n13710) );
  ANDN U19343 ( .B(n16969), .A(n14557), .Z(n19795) );
  XOR U19344 ( .A(n19797), .B(n18609), .Z(n14557) );
  XNOR U19345 ( .A(n19288), .B(n19798), .Z(n18609) );
  XOR U19346 ( .A(n19799), .B(n19800), .Z(n19288) );
  XNOR U19347 ( .A(n19013), .B(n19531), .Z(n19800) );
  XOR U19348 ( .A(n19801), .B(n19802), .Z(n19531) );
  NOR U19349 ( .A(n19803), .B(n19804), .Z(n19801) );
  XOR U19350 ( .A(n19805), .B(n19806), .Z(n19013) );
  XOR U19351 ( .A(n18758), .B(n19809), .Z(n19799) );
  XOR U19352 ( .A(n19345), .B(n19810), .Z(n19809) );
  XNOR U19353 ( .A(n19811), .B(n19812), .Z(n19345) );
  NOR U19354 ( .A(n19813), .B(n19814), .Z(n19811) );
  XNOR U19355 ( .A(n19815), .B(n19816), .Z(n18758) );
  ANDN U19356 ( .B(n19817), .A(n19818), .Z(n19815) );
  XOR U19357 ( .A(n16024), .B(n19819), .Z(n16969) );
  XNOR U19358 ( .A(n19820), .B(n13720), .Z(n14545) );
  XNOR U19359 ( .A(n19821), .B(n15588), .Z(n13720) );
  ANDN U19360 ( .B(n14554), .A(n16965), .Z(n19820) );
  XNOR U19361 ( .A(n19822), .B(n18816), .Z(n16965) );
  IV U19362 ( .A(n16261), .Z(n18816) );
  XOR U19363 ( .A(n19498), .B(n18330), .Z(n16261) );
  XOR U19364 ( .A(n19823), .B(n19824), .Z(n18330) );
  XOR U19365 ( .A(n17384), .B(n19001), .Z(n19824) );
  XOR U19366 ( .A(n19825), .B(n19826), .Z(n19001) );
  AND U19367 ( .A(n19827), .B(n19828), .Z(n19825) );
  XNOR U19368 ( .A(n19829), .B(n19830), .Z(n17384) );
  ANDN U19369 ( .B(n19831), .A(n19832), .Z(n19829) );
  XOR U19370 ( .A(n19833), .B(n19834), .Z(n19823) );
  XOR U19371 ( .A(n16336), .B(n19835), .Z(n19834) );
  XNOR U19372 ( .A(n19836), .B(n19837), .Z(n16336) );
  AND U19373 ( .A(n19838), .B(n19839), .Z(n19836) );
  XNOR U19374 ( .A(n19840), .B(n19841), .Z(n19498) );
  XNOR U19375 ( .A(n19783), .B(n19683), .Z(n19841) );
  XOR U19376 ( .A(n19842), .B(n19843), .Z(n19683) );
  ANDN U19377 ( .B(n19844), .A(n19845), .Z(n19842) );
  XNOR U19378 ( .A(n19846), .B(n19847), .Z(n19783) );
  ANDN U19379 ( .B(n19848), .A(n19849), .Z(n19846) );
  XOR U19380 ( .A(n17219), .B(n19850), .Z(n19840) );
  XOR U19381 ( .A(n16671), .B(n19379), .Z(n19850) );
  XNOR U19382 ( .A(n19851), .B(n19852), .Z(n19379) );
  AND U19383 ( .A(n19853), .B(n19854), .Z(n19851) );
  XNOR U19384 ( .A(n19855), .B(n19856), .Z(n16671) );
  ANDN U19385 ( .B(n19857), .A(n19858), .Z(n19855) );
  XNOR U19386 ( .A(n19859), .B(n19860), .Z(n17219) );
  AND U19387 ( .A(n19861), .B(n19862), .Z(n19859) );
  XOR U19388 ( .A(n19863), .B(n17504), .Z(n14554) );
  IV U19389 ( .A(n16469), .Z(n17504) );
  XNOR U19390 ( .A(n19864), .B(n18767), .Z(n16469) );
  XOR U19391 ( .A(n19865), .B(n19866), .Z(n18767) );
  XNOR U19392 ( .A(n18688), .B(n17940), .Z(n19866) );
  XOR U19393 ( .A(n19867), .B(n19868), .Z(n17940) );
  AND U19394 ( .A(n19869), .B(n19870), .Z(n19867) );
  XNOR U19395 ( .A(n19871), .B(n19872), .Z(n18688) );
  NOR U19396 ( .A(n19873), .B(n19874), .Z(n19871) );
  XNOR U19397 ( .A(n18289), .B(n19875), .Z(n19865) );
  XOR U19398 ( .A(n16949), .B(n18644), .Z(n19875) );
  XNOR U19399 ( .A(n19876), .B(n19877), .Z(n18644) );
  ANDN U19400 ( .B(n19878), .A(n19879), .Z(n19876) );
  XNOR U19401 ( .A(n19880), .B(n19881), .Z(n16949) );
  AND U19402 ( .A(n19882), .B(n19883), .Z(n19880) );
  XNOR U19403 ( .A(n19884), .B(n19885), .Z(n18289) );
  AND U19404 ( .A(n19886), .B(n19887), .Z(n19884) );
  XOR U19405 ( .A(n12188), .B(n19888), .Z(n19793) );
  XNOR U19406 ( .A(n12911), .B(n11907), .Z(n19888) );
  XNOR U19407 ( .A(n19889), .B(n14551), .Z(n11907) );
  XNOR U19408 ( .A(n19890), .B(n17937), .Z(n14551) );
  IV U19409 ( .A(n17039), .Z(n17937) );
  ANDN U19410 ( .B(n14552), .A(n17336), .Z(n19889) );
  XNOR U19411 ( .A(n19891), .B(n13716), .Z(n12911) );
  XOR U19412 ( .A(n19892), .B(n18258), .Z(n13716) );
  XNOR U19413 ( .A(n19893), .B(n19894), .Z(n18258) );
  AND U19414 ( .A(n16963), .B(n14559), .Z(n19891) );
  XNOR U19415 ( .A(n15903), .B(n19895), .Z(n14559) );
  XOR U19416 ( .A(n19896), .B(n17560), .Z(n16963) );
  XNOR U19417 ( .A(n19897), .B(n13706), .Z(n12188) );
  XNOR U19418 ( .A(n18527), .B(n19898), .Z(n13706) );
  ANDN U19419 ( .B(n14561), .A(n16971), .Z(n19897) );
  XNOR U19420 ( .A(n19899), .B(n17908), .Z(n16971) );
  XOR U19421 ( .A(n19900), .B(n18805), .Z(n14561) );
  IV U19422 ( .A(n15856), .Z(n18805) );
  XNOR U19423 ( .A(n19901), .B(n19902), .Z(n15856) );
  XNOR U19424 ( .A(n19903), .B(n14552), .Z(n16967) );
  XNOR U19425 ( .A(n19904), .B(n18566), .Z(n14552) );
  IV U19426 ( .A(n18368), .Z(n18566) );
  XNOR U19427 ( .A(n19905), .B(n19906), .Z(n18368) );
  AND U19428 ( .A(n17336), .B(n17337), .Z(n19903) );
  XOR U19429 ( .A(n19907), .B(n17131), .Z(n17337) );
  IV U19430 ( .A(n17987), .Z(n17131) );
  XNOR U19431 ( .A(n19908), .B(n17564), .Z(n17336) );
  XOR U19432 ( .A(n19192), .B(n12662), .Z(n9211) );
  XOR U19433 ( .A(n11327), .B(n12926), .Z(n12662) );
  XOR U19434 ( .A(n19909), .B(n19910), .Z(n12926) );
  XNOR U19435 ( .A(n12286), .B(n10801), .Z(n19910) );
  XOR U19436 ( .A(n19911), .B(n18030), .Z(n10801) );
  XOR U19437 ( .A(n19912), .B(n18651), .Z(n18030) );
  IV U19438 ( .A(n17208), .Z(n18651) );
  XNOR U19439 ( .A(n19913), .B(n19784), .Z(n17208) );
  XOR U19440 ( .A(n19914), .B(n19915), .Z(n19784) );
  XOR U19441 ( .A(n19916), .B(n19033), .Z(n19915) );
  XOR U19442 ( .A(n19917), .B(n19918), .Z(n19033) );
  ANDN U19443 ( .B(n19852), .A(n19853), .Z(n19917) );
  XOR U19444 ( .A(n16059), .B(n19919), .Z(n19914) );
  XOR U19445 ( .A(n19618), .B(n17868), .Z(n19919) );
  XOR U19446 ( .A(n19920), .B(n19921), .Z(n17868) );
  ANDN U19447 ( .B(n19847), .A(n19848), .Z(n19920) );
  XNOR U19448 ( .A(n19922), .B(n19923), .Z(n19618) );
  ANDN U19449 ( .B(n19856), .A(n19857), .Z(n19922) );
  XOR U19450 ( .A(n19924), .B(n19925), .Z(n16059) );
  AND U19451 ( .A(n18671), .B(n18057), .Z(n19911) );
  IV U19452 ( .A(n19173), .Z(n18057) );
  XOR U19453 ( .A(n16903), .B(n19926), .Z(n19173) );
  XOR U19454 ( .A(n19927), .B(n19928), .Z(n16903) );
  XOR U19455 ( .A(n15647), .B(n19929), .Z(n18671) );
  XOR U19456 ( .A(n19930), .B(n17094), .Z(n12286) );
  XOR U19457 ( .A(n19931), .B(n19932), .Z(n17094) );
  AND U19458 ( .A(n18664), .B(n18061), .Z(n19930) );
  XOR U19459 ( .A(n16954), .B(n19933), .Z(n18061) );
  XOR U19460 ( .A(n19934), .B(n18856), .Z(n16954) );
  XNOR U19461 ( .A(n19935), .B(n19936), .Z(n18856) );
  XNOR U19462 ( .A(n17808), .B(n18168), .Z(n19936) );
  XNOR U19463 ( .A(n19937), .B(n19938), .Z(n18168) );
  NOR U19464 ( .A(n19812), .B(n19939), .Z(n19937) );
  XOR U19465 ( .A(n19940), .B(n19941), .Z(n17808) );
  ANDN U19466 ( .B(n19802), .A(n19942), .Z(n19940) );
  XOR U19467 ( .A(n18020), .B(n19943), .Z(n19935) );
  XOR U19468 ( .A(n19944), .B(n15256), .Z(n19943) );
  XNOR U19469 ( .A(n19945), .B(n19946), .Z(n15256) );
  ANDN U19470 ( .B(n19806), .A(n19947), .Z(n19945) );
  XOR U19471 ( .A(n19948), .B(n19949), .Z(n18020) );
  NOR U19472 ( .A(n19950), .B(n19951), .Z(n19948) );
  XOR U19473 ( .A(n19952), .B(n18222), .Z(n18664) );
  XOR U19474 ( .A(n13279), .B(n19953), .Z(n19909) );
  XOR U19475 ( .A(n9481), .B(n18626), .Z(n19953) );
  XOR U19476 ( .A(n19954), .B(n17091), .Z(n18626) );
  XOR U19477 ( .A(n17332), .B(n19955), .Z(n17091) );
  XOR U19478 ( .A(n19956), .B(n19957), .Z(n17332) );
  AND U19479 ( .A(n18668), .B(n18059), .Z(n19954) );
  XOR U19480 ( .A(n19958), .B(n17925), .Z(n18059) );
  XNOR U19481 ( .A(n19959), .B(n15137), .Z(n18668) );
  IV U19482 ( .A(n17341), .Z(n15137) );
  XOR U19483 ( .A(n19960), .B(n19961), .Z(n17341) );
  XOR U19484 ( .A(n19962), .B(n18674), .Z(n9481) );
  IV U19485 ( .A(n17101), .Z(n18674) );
  XOR U19486 ( .A(n19963), .B(n18215), .Z(n17101) );
  ANDN U19487 ( .B(n18675), .A(n18051), .Z(n19962) );
  XNOR U19488 ( .A(n19568), .B(n16256), .Z(n18051) );
  XNOR U19489 ( .A(n19964), .B(n19965), .Z(n19568) );
  ANDN U19490 ( .B(n19966), .A(n19967), .Z(n19964) );
  XOR U19491 ( .A(n19159), .B(n19968), .Z(n18675) );
  XNOR U19492 ( .A(n19969), .B(n17105), .Z(n13279) );
  XNOR U19493 ( .A(n19970), .B(n19971), .Z(n17105) );
  AND U19494 ( .A(n18660), .B(n19169), .Z(n19969) );
  XOR U19495 ( .A(n19643), .B(n19491), .Z(n19169) );
  IV U19496 ( .A(n19597), .Z(n19491) );
  XOR U19497 ( .A(n19972), .B(n19973), .Z(n19643) );
  ANDN U19498 ( .B(n19525), .A(n19526), .Z(n19972) );
  XNOR U19499 ( .A(n19974), .B(n16555), .Z(n18660) );
  XOR U19500 ( .A(n19975), .B(n19976), .Z(n11327) );
  XOR U19501 ( .A(n11367), .B(n12211), .Z(n19976) );
  XOR U19502 ( .A(n19977), .B(n12438), .Z(n12211) );
  XOR U19503 ( .A(n19978), .B(n17928), .Z(n12438) );
  ANDN U19504 ( .B(n18910), .A(n12437), .Z(n19977) );
  XOR U19505 ( .A(n19979), .B(n19732), .Z(n12437) );
  XOR U19506 ( .A(n19980), .B(n19665), .Z(n18910) );
  IV U19507 ( .A(n18222), .Z(n19665) );
  XNOR U19508 ( .A(n19981), .B(n17108), .Z(n11367) );
  XNOR U19509 ( .A(n19982), .B(n18721), .Z(n17108) );
  NOR U19510 ( .A(n17107), .B(n14307), .Z(n19981) );
  XNOR U19511 ( .A(n19983), .B(n19984), .Z(n14307) );
  XNOR U19512 ( .A(n19985), .B(n18707), .Z(n17107) );
  XNOR U19513 ( .A(n12086), .B(n19986), .Z(n19975) );
  XOR U19514 ( .A(n11702), .B(n9908), .Z(n19986) );
  XOR U19515 ( .A(n19987), .B(n12434), .Z(n9908) );
  XNOR U19516 ( .A(n19988), .B(n18869), .Z(n12434) );
  XOR U19517 ( .A(n19989), .B(n19990), .Z(n18869) );
  AND U19518 ( .A(n12433), .B(n14303), .Z(n19987) );
  IV U19519 ( .A(n19991), .Z(n14303) );
  XOR U19520 ( .A(n19992), .B(n12424), .Z(n11702) );
  XNOR U19521 ( .A(n19993), .B(n15244), .Z(n12424) );
  IV U19522 ( .A(n17895), .Z(n15244) );
  XNOR U19523 ( .A(n19994), .B(n19995), .Z(n19625) );
  XOR U19524 ( .A(n18144), .B(n19996), .Z(n19995) );
  XNOR U19525 ( .A(n19997), .B(n19998), .Z(n18144) );
  ANDN U19526 ( .B(n19999), .A(n20000), .Z(n19997) );
  XOR U19527 ( .A(n20001), .B(n20002), .Z(n19994) );
  XNOR U19528 ( .A(n18466), .B(n16681), .Z(n20002) );
  XNOR U19529 ( .A(n20003), .B(n20004), .Z(n16681) );
  AND U19530 ( .A(n20005), .B(n20006), .Z(n20003) );
  XNOR U19531 ( .A(n20007), .B(n20008), .Z(n18466) );
  AND U19532 ( .A(n12423), .B(n19198), .Z(n19992) );
  IV U19533 ( .A(n19196), .Z(n19198) );
  XOR U19534 ( .A(n20012), .B(n17069), .Z(n19196) );
  XNOR U19535 ( .A(n19648), .B(n19597), .Z(n12423) );
  XNOR U19536 ( .A(n20013), .B(n20014), .Z(n19648) );
  ANDN U19537 ( .B(n19521), .A(n19522), .Z(n20013) );
  XOR U19538 ( .A(n20015), .B(n12428), .Z(n12086) );
  IV U19539 ( .A(n17424), .Z(n12428) );
  XOR U19540 ( .A(n19244), .B(n20016), .Z(n17424) );
  IV U19541 ( .A(n18156), .Z(n19244) );
  NOR U19542 ( .A(n12427), .B(n14314), .Z(n20015) );
  XNOR U19543 ( .A(n20017), .B(n18494), .Z(n14314) );
  IV U19544 ( .A(n19186), .Z(n12427) );
  XOR U19545 ( .A(n20018), .B(n17188), .Z(n19186) );
  IV U19546 ( .A(n17908), .Z(n17188) );
  XNOR U19547 ( .A(n20019), .B(n20020), .Z(n17908) );
  XOR U19548 ( .A(n20021), .B(n12433), .Z(n19192) );
  XNOR U19549 ( .A(n19150), .B(n20022), .Z(n12433) );
  AND U19550 ( .A(n14305), .B(n19991), .Z(n20021) );
  XNOR U19551 ( .A(n20023), .B(n17925), .Z(n19991) );
  XNOR U19552 ( .A(n20024), .B(n20025), .Z(n14305) );
  XNOR U19553 ( .A(n20026), .B(n6630), .Z(n4868) );
  XNOR U19554 ( .A(n9669), .B(n15980), .Z(n6630) );
  XOR U19555 ( .A(n20027), .B(n13982), .Z(n15980) );
  AND U19556 ( .A(n14527), .B(n14525), .Z(n20027) );
  XNOR U19557 ( .A(n20028), .B(n19657), .Z(n14527) );
  XOR U19558 ( .A(n20029), .B(n20030), .Z(n19657) );
  IV U19559 ( .A(n10374), .Z(n9669) );
  XOR U19560 ( .A(n12091), .B(n18467), .Z(n10374) );
  XOR U19561 ( .A(n20031), .B(n20032), .Z(n18467) );
  XNOR U19562 ( .A(n13360), .B(n11303), .Z(n20032) );
  XNOR U19563 ( .A(n20033), .B(n16106), .Z(n11303) );
  XNOR U19564 ( .A(n16687), .B(n20034), .Z(n16106) );
  IV U19565 ( .A(n18485), .Z(n16687) );
  ANDN U19566 ( .B(n14516), .A(n15996), .Z(n20033) );
  XOR U19567 ( .A(n16547), .B(n20035), .Z(n15996) );
  XOR U19568 ( .A(n20036), .B(n19732), .Z(n14516) );
  XOR U19569 ( .A(n20037), .B(n16096), .Z(n13360) );
  XOR U19570 ( .A(n20038), .B(n15129), .Z(n16096) );
  AND U19571 ( .A(n14512), .B(n17624), .Z(n20037) );
  XOR U19572 ( .A(n20039), .B(n18102), .Z(n17624) );
  XNOR U19573 ( .A(n20040), .B(n17270), .Z(n14512) );
  XOR U19574 ( .A(n18948), .B(n20041), .Z(n17270) );
  XNOR U19575 ( .A(n20042), .B(n20043), .Z(n18948) );
  XNOR U19576 ( .A(n18903), .B(n19174), .Z(n20043) );
  XOR U19577 ( .A(n20044), .B(n20045), .Z(n19174) );
  ANDN U19578 ( .B(n20046), .A(n20047), .Z(n20044) );
  XOR U19579 ( .A(n20048), .B(n20049), .Z(n18903) );
  AND U19580 ( .A(n20050), .B(n20051), .Z(n20048) );
  XOR U19581 ( .A(n16939), .B(n20052), .Z(n20042) );
  XOR U19582 ( .A(n17852), .B(n19154), .Z(n20052) );
  XNOR U19583 ( .A(n20053), .B(n20054), .Z(n19154) );
  ANDN U19584 ( .B(n20055), .A(n20056), .Z(n20053) );
  XOR U19585 ( .A(n20057), .B(n20058), .Z(n17852) );
  ANDN U19586 ( .B(n20059), .A(n20060), .Z(n20057) );
  XNOR U19587 ( .A(n20061), .B(n20062), .Z(n16939) );
  NOR U19588 ( .A(n20063), .B(n20064), .Z(n20061) );
  XOR U19589 ( .A(n9891), .B(n20065), .Z(n20031) );
  XOR U19590 ( .A(n9068), .B(n17601), .Z(n20065) );
  XOR U19591 ( .A(n20066), .B(n17628), .Z(n17601) );
  IV U19592 ( .A(n16093), .Z(n17628) );
  XOR U19593 ( .A(n19944), .B(n17809), .Z(n16093) );
  XNOR U19594 ( .A(n20067), .B(n20068), .Z(n17809) );
  XNOR U19595 ( .A(n20069), .B(n20070), .Z(n19944) );
  NOR U19596 ( .A(n19816), .B(n20071), .Z(n20069) );
  AND U19597 ( .A(n17629), .B(n18496), .Z(n20066) );
  XNOR U19598 ( .A(n20072), .B(n16465), .Z(n18496) );
  XNOR U19599 ( .A(n20073), .B(n18594), .Z(n17629) );
  XNOR U19600 ( .A(n20074), .B(n16101), .Z(n9068) );
  IV U19601 ( .A(n17621), .Z(n16101) );
  XOR U19602 ( .A(n20075), .B(n15851), .Z(n17621) );
  ANDN U19603 ( .B(n14503), .A(n15992), .Z(n20074) );
  XNOR U19604 ( .A(n20078), .B(n20079), .Z(n15992) );
  XOR U19605 ( .A(n17680), .B(n20080), .Z(n14503) );
  XNOR U19606 ( .A(n20081), .B(n16108), .Z(n9891) );
  XNOR U19607 ( .A(n20082), .B(n15984), .Z(n16108) );
  XOR U19608 ( .A(n20083), .B(n18254), .Z(n14499) );
  XOR U19609 ( .A(n20084), .B(n20085), .Z(n18254) );
  XNOR U19610 ( .A(n20086), .B(n17566), .Z(n16317) );
  IV U19611 ( .A(n19441), .Z(n17566) );
  XOR U19612 ( .A(n20087), .B(n20088), .Z(n12091) );
  XNOR U19613 ( .A(n12127), .B(n13110), .Z(n20088) );
  XOR U19614 ( .A(n20089), .B(n13978), .Z(n13110) );
  XOR U19615 ( .A(n17997), .B(n20090), .Z(n13978) );
  IV U19616 ( .A(n17198), .Z(n17997) );
  AND U19617 ( .A(n13979), .B(n14531), .Z(n20089) );
  IV U19618 ( .A(n15982), .Z(n14531) );
  XNOR U19619 ( .A(n20091), .B(n18102), .Z(n15982) );
  XOR U19620 ( .A(n20092), .B(n18180), .Z(n13979) );
  XNOR U19621 ( .A(n20093), .B(n13983), .Z(n12127) );
  XOR U19622 ( .A(n16035), .B(n20094), .Z(n13983) );
  IV U19623 ( .A(n19159), .Z(n16035) );
  XOR U19624 ( .A(n20095), .B(n20096), .Z(n19159) );
  ANDN U19625 ( .B(n13982), .A(n14525), .Z(n20093) );
  XNOR U19626 ( .A(n20097), .B(n17962), .Z(n14525) );
  XNOR U19627 ( .A(n20098), .B(n17730), .Z(n13982) );
  XOR U19628 ( .A(n18284), .B(n20041), .Z(n17730) );
  XNOR U19629 ( .A(n20099), .B(n20100), .Z(n20041) );
  XOR U19630 ( .A(n16752), .B(n17213), .Z(n20100) );
  XOR U19631 ( .A(n20101), .B(n19869), .Z(n17213) );
  ANDN U19632 ( .B(n20102), .A(n20103), .Z(n20101) );
  XOR U19633 ( .A(n20104), .B(n20105), .Z(n16752) );
  NOR U19634 ( .A(n20106), .B(n20107), .Z(n20104) );
  XNOR U19635 ( .A(n17671), .B(n20108), .Z(n20099) );
  XNOR U19636 ( .A(n20109), .B(n20110), .Z(n20108) );
  XNOR U19637 ( .A(n20111), .B(n19886), .Z(n17671) );
  NOR U19638 ( .A(n20112), .B(n20113), .Z(n20111) );
  XNOR U19639 ( .A(n20114), .B(n20115), .Z(n18284) );
  XNOR U19640 ( .A(n17578), .B(n19061), .Z(n20115) );
  XNOR U19641 ( .A(n20116), .B(n19677), .Z(n19061) );
  XNOR U19642 ( .A(n20119), .B(n18843), .Z(n17578) );
  ANDN U19643 ( .B(n20120), .A(n20121), .Z(n20119) );
  XOR U19644 ( .A(n17492), .B(n20122), .Z(n20114) );
  XNOR U19645 ( .A(n19221), .B(n20123), .Z(n20122) );
  XNOR U19646 ( .A(n20124), .B(n18776), .Z(n19221) );
  ANDN U19647 ( .B(n20125), .A(n20126), .Z(n20124) );
  XNOR U19648 ( .A(n20127), .B(n20128), .Z(n17492) );
  ANDN U19649 ( .B(n20129), .A(n20130), .Z(n20127) );
  XOR U19650 ( .A(n11441), .B(n20131), .Z(n20087) );
  XOR U19651 ( .A(n10280), .B(n12838), .Z(n20131) );
  XNOR U19652 ( .A(n20132), .B(n13974), .Z(n12838) );
  XNOR U19653 ( .A(n20133), .B(n18736), .Z(n13974) );
  XNOR U19654 ( .A(n20134), .B(n20135), .Z(n18736) );
  ANDN U19655 ( .B(n15978), .A(n13973), .Z(n20132) );
  XNOR U19656 ( .A(n20136), .B(n18721), .Z(n13973) );
  IV U19657 ( .A(n17502), .Z(n18721) );
  XNOR U19658 ( .A(n20137), .B(n17231), .Z(n15978) );
  XNOR U19659 ( .A(n20138), .B(n13986), .Z(n10280) );
  XNOR U19660 ( .A(n20139), .B(n17520), .Z(n13986) );
  XNOR U19661 ( .A(n20140), .B(n18534), .Z(n17520) );
  XNOR U19662 ( .A(n20141), .B(n20142), .Z(n18534) );
  XOR U19663 ( .A(n19455), .B(n18385), .Z(n20142) );
  XOR U19664 ( .A(n20143), .B(n20144), .Z(n18385) );
  AND U19665 ( .A(n20145), .B(n20146), .Z(n20143) );
  XNOR U19666 ( .A(n20147), .B(n20148), .Z(n19455) );
  ANDN U19667 ( .B(n20149), .A(n20150), .Z(n20147) );
  XOR U19668 ( .A(n18256), .B(n20151), .Z(n20141) );
  XOR U19669 ( .A(n16811), .B(n17731), .Z(n20151) );
  XNOR U19670 ( .A(n20152), .B(n20153), .Z(n17731) );
  AND U19671 ( .A(n20154), .B(n20155), .Z(n20152) );
  XNOR U19672 ( .A(n20156), .B(n20157), .Z(n16811) );
  AND U19673 ( .A(n20158), .B(n20159), .Z(n20156) );
  XNOR U19674 ( .A(n20160), .B(n20161), .Z(n18256) );
  AND U19675 ( .A(n20162), .B(n20163), .Z(n20160) );
  AND U19676 ( .A(n13987), .B(n14522), .Z(n20138) );
  IV U19677 ( .A(n15973), .Z(n14522) );
  XNOR U19678 ( .A(n20164), .B(n16465), .Z(n15973) );
  XOR U19679 ( .A(n15913), .B(n20165), .Z(n13987) );
  XOR U19680 ( .A(n20166), .B(n13970), .Z(n11441) );
  XOR U19681 ( .A(n20167), .B(n15204), .Z(n13970) );
  XOR U19682 ( .A(n19893), .B(n20168), .Z(n15204) );
  XOR U19683 ( .A(n20169), .B(n20170), .Z(n19893) );
  XNOR U19684 ( .A(n19316), .B(n18507), .Z(n20170) );
  XOR U19685 ( .A(n20171), .B(n20172), .Z(n18507) );
  AND U19686 ( .A(n20173), .B(n20174), .Z(n20171) );
  XNOR U19687 ( .A(n20175), .B(n20176), .Z(n19316) );
  ANDN U19688 ( .B(n20177), .A(n20178), .Z(n20175) );
  XNOR U19689 ( .A(n20179), .B(n20180), .Z(n20169) );
  XOR U19690 ( .A(n17801), .B(n17120), .Z(n20180) );
  XNOR U19691 ( .A(n20181), .B(n20182), .Z(n17120) );
  ANDN U19692 ( .B(n20183), .A(n20184), .Z(n20181) );
  XNOR U19693 ( .A(n20185), .B(n20186), .Z(n17801) );
  NOR U19694 ( .A(n20187), .B(n20188), .Z(n20185) );
  ANDN U19695 ( .B(n14534), .A(n13969), .Z(n20166) );
  XOR U19696 ( .A(n17680), .B(n20189), .Z(n13969) );
  IV U19697 ( .A(n16471), .Z(n17680) );
  XOR U19698 ( .A(n20192), .B(n19558), .Z(n14534) );
  IV U19699 ( .A(n18334), .Z(n19558) );
  XNOR U19700 ( .A(n20193), .B(n20194), .Z(n18334) );
  ANDN U19701 ( .B(n7069), .A(n9206), .Z(n20026) );
  XOR U19702 ( .A(n18605), .B(n13315), .Z(n9206) );
  XOR U19703 ( .A(n18443), .B(n19006), .Z(n13315) );
  XNOR U19704 ( .A(n20195), .B(n20196), .Z(n19006) );
  XNOR U19705 ( .A(n12289), .B(n14055), .Z(n20196) );
  XOR U19706 ( .A(n20197), .B(n15762), .Z(n14055) );
  XNOR U19707 ( .A(n20198), .B(n15984), .Z(n15762) );
  XOR U19708 ( .A(n20199), .B(n20200), .Z(n15984) );
  ANDN U19709 ( .B(n15448), .A(n15761), .Z(n20197) );
  XNOR U19710 ( .A(n20201), .B(n15757), .Z(n12289) );
  XNOR U19711 ( .A(n20202), .B(n17163), .Z(n15757) );
  IV U19712 ( .A(n15122), .Z(n17163) );
  XNOR U19713 ( .A(n20203), .B(n20204), .Z(n15122) );
  XOR U19714 ( .A(n20205), .B(n17369), .Z(n15758) );
  IV U19715 ( .A(n20079), .Z(n17369) );
  XOR U19716 ( .A(n19289), .B(n20206), .Z(n20079) );
  XNOR U19717 ( .A(n20207), .B(n20208), .Z(n19289) );
  XNOR U19718 ( .A(n20039), .B(n18101), .Z(n20208) );
  XOR U19719 ( .A(n20209), .B(n20210), .Z(n18101) );
  ANDN U19720 ( .B(n20211), .A(n20212), .Z(n20209) );
  XNOR U19721 ( .A(n20213), .B(n20214), .Z(n20039) );
  ANDN U19722 ( .B(n20215), .A(n20216), .Z(n20213) );
  XNOR U19723 ( .A(n18441), .B(n20217), .Z(n20207) );
  XNOR U19724 ( .A(n20091), .B(n20218), .Z(n20217) );
  XNOR U19725 ( .A(n20219), .B(n20220), .Z(n20091) );
  AND U19726 ( .A(n20221), .B(n20222), .Z(n20219) );
  XNOR U19727 ( .A(n20223), .B(n20224), .Z(n18441) );
  AND U19728 ( .A(n20225), .B(n20226), .Z(n20223) );
  XOR U19729 ( .A(n18545), .B(n20227), .Z(n14151) );
  XNOR U19730 ( .A(n20228), .B(n20229), .Z(n18545) );
  XOR U19731 ( .A(n11170), .B(n20230), .Z(n20195) );
  XOR U19732 ( .A(n10937), .B(n12003), .Z(n20230) );
  XNOR U19733 ( .A(n20231), .B(n15754), .Z(n12003) );
  XOR U19734 ( .A(n20232), .B(n19337), .Z(n15754) );
  XOR U19735 ( .A(n20233), .B(n15588), .Z(n15755) );
  IV U19736 ( .A(n20234), .Z(n15588) );
  IV U19737 ( .A(n18618), .Z(n18619) );
  XOR U19738 ( .A(n20235), .B(n17469), .Z(n18618) );
  XNOR U19739 ( .A(n20238), .B(n15767), .Z(n10937) );
  XOR U19740 ( .A(n20239), .B(n16938), .Z(n15767) );
  AND U19741 ( .A(n15768), .B(n14147), .Z(n20238) );
  IV U19742 ( .A(n18612), .Z(n14147) );
  XOR U19743 ( .A(n20240), .B(n16362), .Z(n18612) );
  XNOR U19744 ( .A(n20241), .B(n20242), .Z(n16362) );
  XNOR U19745 ( .A(n20243), .B(n20244), .Z(n15768) );
  XNOR U19746 ( .A(n20245), .B(n15765), .Z(n11170) );
  XOR U19747 ( .A(n17860), .B(n20246), .Z(n15765) );
  ANDN U19748 ( .B(n14141), .A(n15764), .Z(n20245) );
  XOR U19749 ( .A(n20247), .B(n16100), .Z(n15764) );
  XNOR U19750 ( .A(n20248), .B(n18849), .Z(n16100) );
  XNOR U19751 ( .A(n20249), .B(n20250), .Z(n18849) );
  XOR U19752 ( .A(n16618), .B(n16000), .Z(n20250) );
  XOR U19753 ( .A(n20251), .B(n20252), .Z(n16000) );
  XNOR U19754 ( .A(n20255), .B(n20256), .Z(n16618) );
  ANDN U19755 ( .B(n20257), .A(n20258), .Z(n20255) );
  XOR U19756 ( .A(n16056), .B(n20259), .Z(n20249) );
  XOR U19757 ( .A(n20260), .B(n18321), .Z(n20259) );
  XNOR U19758 ( .A(n20261), .B(n20262), .Z(n18321) );
  XNOR U19759 ( .A(n20265), .B(n20266), .Z(n16056) );
  ANDN U19760 ( .B(n20267), .A(n20268), .Z(n20265) );
  IV U19761 ( .A(n18607), .Z(n14141) );
  XOR U19762 ( .A(n20269), .B(n20270), .Z(n18607) );
  XOR U19763 ( .A(n20271), .B(n20272), .Z(n18443) );
  XNOR U19764 ( .A(n10058), .B(n10776), .Z(n20272) );
  XNOR U19765 ( .A(n20273), .B(n16839), .Z(n10776) );
  XNOR U19766 ( .A(n20274), .B(n16532), .Z(n16839) );
  IV U19767 ( .A(n16539), .Z(n16532) );
  AND U19768 ( .A(n16843), .B(n14638), .Z(n20273) );
  XOR U19769 ( .A(n17223), .B(n20275), .Z(n14638) );
  XOR U19770 ( .A(n14068), .B(n20277), .Z(n10058) );
  XOR U19771 ( .A(n20278), .B(n20279), .Z(n20277) );
  NAND U19772 ( .A(n15691), .B(n11363), .Z(n20279) );
  ANDN U19773 ( .B(n14067), .A(n17152), .Z(n20278) );
  XNOR U19774 ( .A(n17389), .B(n20280), .Z(n17152) );
  XOR U19775 ( .A(n17860), .B(n20283), .Z(n14067) );
  XOR U19776 ( .A(n19717), .B(n20284), .Z(n17860) );
  XOR U19777 ( .A(n20285), .B(n20286), .Z(n19717) );
  XOR U19778 ( .A(n18686), .B(n18440), .Z(n20286) );
  XOR U19779 ( .A(n20287), .B(n20288), .Z(n18440) );
  ANDN U19780 ( .B(n20289), .A(n20290), .Z(n20287) );
  XNOR U19781 ( .A(n20291), .B(n20292), .Z(n18686) );
  XOR U19782 ( .A(n18865), .B(n20295), .Z(n20285) );
  XOR U19783 ( .A(n18393), .B(n16998), .Z(n20295) );
  XNOR U19784 ( .A(n20296), .B(n20297), .Z(n16998) );
  XNOR U19785 ( .A(n20300), .B(n20301), .Z(n18393) );
  ANDN U19786 ( .B(n20302), .A(n20303), .Z(n20300) );
  XNOR U19787 ( .A(n20304), .B(n20305), .Z(n18865) );
  ANDN U19788 ( .B(n20306), .A(n20307), .Z(n20304) );
  XNOR U19789 ( .A(n20308), .B(n17546), .Z(n14068) );
  XNOR U19790 ( .A(n20309), .B(n20310), .Z(n17546) );
  XOR U19791 ( .A(n9895), .B(n20311), .Z(n20271) );
  XOR U19792 ( .A(n12546), .B(n10247), .Z(n20311) );
  XOR U19793 ( .A(n20312), .B(n14062), .Z(n10247) );
  XNOR U19794 ( .A(n20313), .B(n19314), .Z(n14062) );
  IV U19795 ( .A(n19971), .Z(n19314) );
  AND U19796 ( .A(n14635), .B(n18592), .Z(n20312) );
  XOR U19797 ( .A(n20314), .B(n19724), .Z(n18592) );
  XOR U19798 ( .A(n20315), .B(n20316), .Z(n19724) );
  ANDN U19799 ( .B(n20317), .A(n20318), .Z(n20315) );
  XNOR U19800 ( .A(n20319), .B(n20320), .Z(n14635) );
  XOR U19801 ( .A(n20321), .B(n14075), .Z(n12546) );
  XOR U19802 ( .A(n20322), .B(n18458), .Z(n14075) );
  IV U19803 ( .A(n18940), .Z(n18458) );
  AND U19804 ( .A(n17771), .B(n18596), .Z(n20321) );
  XOR U19805 ( .A(n20323), .B(n17075), .Z(n18596) );
  IV U19806 ( .A(n20324), .Z(n17075) );
  XOR U19807 ( .A(n20325), .B(n15655), .Z(n17771) );
  IV U19808 ( .A(n20025), .Z(n15655) );
  XNOR U19809 ( .A(n20328), .B(n14072), .Z(n9895) );
  XOR U19810 ( .A(n20243), .B(n20329), .Z(n14072) );
  IV U19811 ( .A(n18347), .Z(n20243) );
  XOR U19812 ( .A(n18684), .B(n18986), .Z(n18347) );
  XNOR U19813 ( .A(n20330), .B(n20331), .Z(n18986) );
  XNOR U19814 ( .A(n18250), .B(n19900), .Z(n20331) );
  XNOR U19815 ( .A(n20332), .B(n20333), .Z(n19900) );
  ANDN U19816 ( .B(n20334), .A(n20335), .Z(n20332) );
  XNOR U19817 ( .A(n20336), .B(n20337), .Z(n18250) );
  ANDN U19818 ( .B(n20338), .A(n20339), .Z(n20336) );
  XOR U19819 ( .A(n15855), .B(n20340), .Z(n20330) );
  XNOR U19820 ( .A(n16470), .B(n18804), .Z(n20340) );
  XNOR U19821 ( .A(n20341), .B(n20342), .Z(n18804) );
  ANDN U19822 ( .B(n20343), .A(n20344), .Z(n20341) );
  XNOR U19823 ( .A(n20345), .B(n20346), .Z(n16470) );
  NOR U19824 ( .A(n20347), .B(n20348), .Z(n20345) );
  XNOR U19825 ( .A(n20349), .B(n20350), .Z(n15855) );
  NOR U19826 ( .A(n20351), .B(n20352), .Z(n20349) );
  XNOR U19827 ( .A(n20353), .B(n20354), .Z(n18684) );
  XNOR U19828 ( .A(n20355), .B(n19391), .Z(n20354) );
  XNOR U19829 ( .A(n20356), .B(n20357), .Z(n19391) );
  ANDN U19830 ( .B(n20358), .A(n20359), .Z(n20356) );
  XOR U19831 ( .A(n19036), .B(n20360), .Z(n20353) );
  XOR U19832 ( .A(n20361), .B(n17554), .Z(n20360) );
  XNOR U19833 ( .A(n20362), .B(n20363), .Z(n17554) );
  ANDN U19834 ( .B(n20364), .A(n20365), .Z(n20362) );
  XNOR U19835 ( .A(n20366), .B(n20367), .Z(n19036) );
  ANDN U19836 ( .B(n20368), .A(n20369), .Z(n20366) );
  AND U19837 ( .A(n14071), .B(n15073), .Z(n20328) );
  XOR U19838 ( .A(n14918), .B(n18771), .Z(n15073) );
  XOR U19839 ( .A(n20370), .B(n20371), .Z(n18771) );
  ANDN U19840 ( .B(n20372), .A(n20128), .Z(n20370) );
  XNOR U19841 ( .A(n20373), .B(n20374), .Z(n18690) );
  XOR U19842 ( .A(n17521), .B(n19374), .Z(n20374) );
  XOR U19843 ( .A(n20375), .B(n20376), .Z(n19374) );
  NOR U19844 ( .A(n18780), .B(n18779), .Z(n20375) );
  XNOR U19845 ( .A(n20377), .B(n20130), .Z(n17521) );
  ANDN U19846 ( .B(n20371), .A(n20372), .Z(n20377) );
  XOR U19847 ( .A(n17785), .B(n20378), .Z(n20373) );
  XOR U19848 ( .A(n20379), .B(n18374), .Z(n20378) );
  XNOR U19849 ( .A(n20380), .B(n20121), .Z(n18374) );
  XNOR U19850 ( .A(n20381), .B(n20117), .Z(n17785) );
  XNOR U19851 ( .A(n20382), .B(n20383), .Z(n19457) );
  XOR U19852 ( .A(n20384), .B(n18493), .Z(n20383) );
  XOR U19853 ( .A(n20385), .B(n20386), .Z(n18493) );
  ANDN U19854 ( .B(n20153), .A(n20155), .Z(n20385) );
  XOR U19855 ( .A(n20387), .B(n20388), .Z(n20382) );
  XOR U19856 ( .A(n20017), .B(n16450), .Z(n20388) );
  XOR U19857 ( .A(n20389), .B(n20390), .Z(n16450) );
  ANDN U19858 ( .B(n20161), .A(n20163), .Z(n20389) );
  XOR U19859 ( .A(n20391), .B(n20392), .Z(n20017) );
  ANDN U19860 ( .B(n20157), .A(n20159), .Z(n20391) );
  XNOR U19861 ( .A(n20393), .B(n18434), .Z(n14071) );
  XOR U19862 ( .A(n20394), .B(n15761), .Z(n18605) );
  XOR U19863 ( .A(n20395), .B(n20324), .Z(n15761) );
  XOR U19864 ( .A(n19640), .B(n20396), .Z(n20324) );
  XOR U19865 ( .A(n20397), .B(n20398), .Z(n19640) );
  XNOR U19866 ( .A(n20399), .B(n18497), .Z(n20398) );
  XNOR U19867 ( .A(n20400), .B(n20401), .Z(n18497) );
  ANDN U19868 ( .B(n20402), .A(n20403), .Z(n20400) );
  XOR U19869 ( .A(n18896), .B(n20404), .Z(n20397) );
  XOR U19870 ( .A(n19224), .B(n17403), .Z(n20404) );
  XNOR U19871 ( .A(n20405), .B(n20406), .Z(n17403) );
  ANDN U19872 ( .B(n20407), .A(n20408), .Z(n20405) );
  XNOR U19873 ( .A(n20409), .B(n20410), .Z(n19224) );
  AND U19874 ( .A(n20411), .B(n20412), .Z(n20409) );
  XNOR U19875 ( .A(n20413), .B(n20414), .Z(n18896) );
  ANDN U19876 ( .B(n20415), .A(n20416), .Z(n20413) );
  XNOR U19877 ( .A(n20417), .B(n15129), .Z(n15449) );
  XOR U19878 ( .A(n20384), .B(n18494), .Z(n15448) );
  XOR U19879 ( .A(n20418), .B(n20419), .Z(n20384) );
  ANDN U19880 ( .B(n20144), .A(n20146), .Z(n20418) );
  IV U19881 ( .A(n9207), .Z(n7069) );
  XNOR U19882 ( .A(n16298), .B(n11162), .Z(n9207) );
  XNOR U19883 ( .A(n11914), .B(n16802), .Z(n11162) );
  XNOR U19884 ( .A(n20420), .B(n20421), .Z(n16802) );
  XNOR U19885 ( .A(n11511), .B(n10287), .Z(n20421) );
  XOR U19886 ( .A(n20422), .B(n17286), .Z(n10287) );
  XOR U19887 ( .A(n20423), .B(n17892), .Z(n17286) );
  AND U19888 ( .A(n16300), .B(n11960), .Z(n20422) );
  XOR U19889 ( .A(n20424), .B(n17917), .Z(n11960) );
  XNOR U19890 ( .A(n20425), .B(n19048), .Z(n17917) );
  XNOR U19891 ( .A(n20426), .B(n20427), .Z(n19048) );
  XOR U19892 ( .A(n16895), .B(n17796), .Z(n20427) );
  XOR U19893 ( .A(n20428), .B(n20429), .Z(n17796) );
  ANDN U19894 ( .B(n20430), .A(n20431), .Z(n20428) );
  XNOR U19895 ( .A(n20432), .B(n20433), .Z(n16895) );
  ANDN U19896 ( .B(n20434), .A(n20435), .Z(n20432) );
  XOR U19897 ( .A(n20436), .B(n20437), .Z(n20426) );
  XOR U19898 ( .A(n17599), .B(n20438), .Z(n20437) );
  XNOR U19899 ( .A(n20439), .B(n20440), .Z(n17599) );
  XOR U19900 ( .A(n20443), .B(n16934), .Z(n16300) );
  XNOR U19901 ( .A(n20445), .B(n20446), .Z(n19653) );
  XOR U19902 ( .A(n17884), .B(n18312), .Z(n20446) );
  XOR U19903 ( .A(n20447), .B(n19479), .Z(n18312) );
  ANDN U19904 ( .B(n19480), .A(n20448), .Z(n20447) );
  XNOR U19905 ( .A(n20449), .B(n19469), .Z(n17884) );
  ANDN U19906 ( .B(n19470), .A(n19729), .Z(n20449) );
  XOR U19907 ( .A(n17359), .B(n20450), .Z(n20445) );
  XOR U19908 ( .A(n18977), .B(n18418), .Z(n20450) );
  XNOR U19909 ( .A(n20451), .B(n19475), .Z(n18418) );
  ANDN U19910 ( .B(n19476), .A(n20452), .Z(n20451) );
  XNOR U19911 ( .A(n20453), .B(n20454), .Z(n18977) );
  ANDN U19912 ( .B(n20455), .A(n20456), .Z(n20453) );
  XNOR U19913 ( .A(n20457), .B(n20458), .Z(n17359) );
  AND U19914 ( .A(n20316), .B(n20459), .Z(n20457) );
  XNOR U19915 ( .A(n20460), .B(n17290), .Z(n11511) );
  XOR U19916 ( .A(n20461), .B(n16069), .Z(n17290) );
  IV U19917 ( .A(n16355), .Z(n16069) );
  XNOR U19918 ( .A(n20462), .B(n20463), .Z(n16355) );
  AND U19919 ( .A(n16302), .B(n11951), .Z(n20460) );
  XOR U19920 ( .A(n20464), .B(n18594), .Z(n11951) );
  XOR U19921 ( .A(n20465), .B(n20320), .Z(n16302) );
  IV U19922 ( .A(n16808), .Z(n20320) );
  XOR U19923 ( .A(n19536), .B(n20466), .Z(n16808) );
  XNOR U19924 ( .A(n20467), .B(n20468), .Z(n19536) );
  XOR U19925 ( .A(n15136), .B(n18041), .Z(n20468) );
  XOR U19926 ( .A(n20469), .B(n20470), .Z(n18041) );
  AND U19927 ( .A(n20471), .B(n20472), .Z(n20469) );
  XNOR U19928 ( .A(n20473), .B(n20474), .Z(n15136) );
  ANDN U19929 ( .B(n20475), .A(n20476), .Z(n20473) );
  XNOR U19930 ( .A(n17340), .B(n20477), .Z(n20467) );
  XOR U19931 ( .A(n18814), .B(n19959), .Z(n20477) );
  XNOR U19932 ( .A(n20478), .B(n20479), .Z(n19959) );
  AND U19933 ( .A(n20480), .B(n20481), .Z(n20478) );
  XNOR U19934 ( .A(n20482), .B(n20483), .Z(n18814) );
  XNOR U19935 ( .A(n20486), .B(n20487), .Z(n17340) );
  XNOR U19936 ( .A(n12255), .B(n20490), .Z(n20420) );
  XNOR U19937 ( .A(n16109), .B(n9598), .Z(n20490) );
  XNOR U19938 ( .A(n20491), .B(n17282), .Z(n9598) );
  XOR U19939 ( .A(n18990), .B(n20492), .Z(n17282) );
  ANDN U19940 ( .B(n17283), .A(n11947), .Z(n20491) );
  XNOR U19941 ( .A(n20493), .B(n17280), .Z(n16109) );
  XOR U19942 ( .A(n20494), .B(n18434), .Z(n17280) );
  XOR U19943 ( .A(n20495), .B(n20203), .Z(n18434) );
  XOR U19944 ( .A(n20496), .B(n20497), .Z(n20203) );
  XOR U19945 ( .A(n17543), .B(n17864), .Z(n20497) );
  XOR U19946 ( .A(n20498), .B(n20499), .Z(n17864) );
  ANDN U19947 ( .B(n20500), .A(n20501), .Z(n20498) );
  XNOR U19948 ( .A(n20502), .B(n19831), .Z(n17543) );
  AND U19949 ( .A(n20503), .B(n19832), .Z(n20502) );
  XOR U19950 ( .A(n14947), .B(n20504), .Z(n20496) );
  XOR U19951 ( .A(n16048), .B(n18328), .Z(n20504) );
  XNOR U19952 ( .A(n20505), .B(n19827), .Z(n18328) );
  XNOR U19953 ( .A(n20507), .B(n19839), .Z(n16048) );
  NOR U19954 ( .A(n20508), .B(n19838), .Z(n20507) );
  XNOR U19955 ( .A(n20509), .B(n20510), .Z(n14947) );
  ANDN U19956 ( .B(n16294), .A(n11964), .Z(n20493) );
  XNOR U19957 ( .A(n20513), .B(n15516), .Z(n11964) );
  IV U19958 ( .A(n19443), .Z(n15516) );
  XOR U19959 ( .A(n19343), .B(n20514), .Z(n19443) );
  XNOR U19960 ( .A(n20515), .B(n20516), .Z(n19343) );
  XNOR U19961 ( .A(n19983), .B(n20517), .Z(n20516) );
  XOR U19962 ( .A(n20518), .B(n20519), .Z(n19983) );
  AND U19963 ( .A(n19356), .B(n20520), .Z(n20518) );
  XOR U19964 ( .A(n20521), .B(n20522), .Z(n20515) );
  XOR U19965 ( .A(n18762), .B(n20523), .Z(n20522) );
  XOR U19966 ( .A(n20524), .B(n20525), .Z(n18762) );
  AND U19967 ( .A(n20526), .B(n19360), .Z(n20524) );
  IV U19968 ( .A(n20527), .Z(n19360) );
  XNOR U19969 ( .A(n20528), .B(n17502), .Z(n16294) );
  XNOR U19970 ( .A(n19120), .B(n19720), .Z(n17502) );
  XNOR U19971 ( .A(n20529), .B(n20530), .Z(n19720) );
  XOR U19972 ( .A(n20531), .B(n18521), .Z(n20530) );
  XOR U19973 ( .A(n20532), .B(n20533), .Z(n18521) );
  AND U19974 ( .A(n20534), .B(n20535), .Z(n20532) );
  XOR U19975 ( .A(n20536), .B(n20537), .Z(n20529) );
  XOR U19976 ( .A(n17484), .B(n18173), .Z(n20537) );
  XNOR U19977 ( .A(n20538), .B(n20539), .Z(n18173) );
  AND U19978 ( .A(n20540), .B(n20541), .Z(n20538) );
  XNOR U19979 ( .A(n20542), .B(n20543), .Z(n17484) );
  AND U19980 ( .A(n20544), .B(n20545), .Z(n20542) );
  XOR U19981 ( .A(n20546), .B(n20547), .Z(n19120) );
  XOR U19982 ( .A(n18267), .B(n17459), .Z(n20547) );
  XOR U19983 ( .A(n20548), .B(n20549), .Z(n17459) );
  ANDN U19984 ( .B(n20550), .A(n20551), .Z(n20548) );
  XNOR U19985 ( .A(n20552), .B(n20553), .Z(n18267) );
  ANDN U19986 ( .B(n20554), .A(n20555), .Z(n20552) );
  XOR U19987 ( .A(n18471), .B(n20556), .Z(n20546) );
  XOR U19988 ( .A(n20557), .B(n16748), .Z(n20556) );
  XNOR U19989 ( .A(n20558), .B(n20559), .Z(n16748) );
  ANDN U19990 ( .B(n20560), .A(n20561), .Z(n20558) );
  XNOR U19991 ( .A(n20562), .B(n20563), .Z(n18471) );
  ANDN U19992 ( .B(n20564), .A(n20565), .Z(n20562) );
  XOR U19993 ( .A(n20566), .B(n17288), .Z(n12255) );
  XNOR U19994 ( .A(n17220), .B(n20567), .Z(n17288) );
  XOR U19995 ( .A(n18689), .B(n20568), .Z(n17220) );
  XOR U19996 ( .A(n20569), .B(n20570), .Z(n18689) );
  XOR U19997 ( .A(n20571), .B(n18269), .Z(n20570) );
  XOR U19998 ( .A(n20572), .B(n20112), .Z(n18269) );
  XOR U19999 ( .A(n16413), .B(n20573), .Z(n20569) );
  XOR U20000 ( .A(n19580), .B(n20574), .Z(n20573) );
  XOR U20001 ( .A(n20575), .B(n20576), .Z(n19580) );
  XNOR U20002 ( .A(n20577), .B(n20106), .Z(n16413) );
  ANDN U20003 ( .B(n19879), .A(n19877), .Z(n20577) );
  AND U20004 ( .A(n16296), .B(n11956), .Z(n20566) );
  XOR U20005 ( .A(n20578), .B(n16674), .Z(n11956) );
  XOR U20006 ( .A(n20581), .B(n19503), .Z(n16296) );
  XOR U20007 ( .A(n20582), .B(n20583), .Z(n11914) );
  XNOR U20008 ( .A(n10133), .B(n11200), .Z(n20583) );
  XOR U20009 ( .A(n20584), .B(n18995), .Z(n11200) );
  XNOR U20010 ( .A(n20585), .B(n17892), .Z(n18995) );
  IV U20011 ( .A(n18140), .Z(n17892) );
  XNOR U20012 ( .A(n20586), .B(n20587), .Z(n20229) );
  XOR U20013 ( .A(n17480), .B(n18226), .Z(n20587) );
  XNOR U20014 ( .A(n20588), .B(n20589), .Z(n18226) );
  ANDN U20015 ( .B(n20590), .A(n20591), .Z(n20588) );
  XNOR U20016 ( .A(n20592), .B(n20369), .Z(n17480) );
  ANDN U20017 ( .B(n20593), .A(n20594), .Z(n20592) );
  XOR U20018 ( .A(n20595), .B(n20596), .Z(n20586) );
  XNOR U20019 ( .A(n16054), .B(n17236), .Z(n20596) );
  XOR U20020 ( .A(n20597), .B(n20598), .Z(n17236) );
  ANDN U20021 ( .B(n20599), .A(n20600), .Z(n20597) );
  XNOR U20022 ( .A(n20601), .B(n20364), .Z(n16054) );
  AND U20023 ( .A(n20602), .B(n20603), .Z(n20601) );
  AND U20024 ( .A(n12801), .B(n19005), .Z(n20584) );
  XOR U20025 ( .A(n20605), .B(n16944), .Z(n19005) );
  XNOR U20026 ( .A(n20606), .B(n20607), .Z(n16944) );
  XNOR U20027 ( .A(n20608), .B(n15322), .Z(n12801) );
  IV U20028 ( .A(n14910), .Z(n15322) );
  XOR U20029 ( .A(n20609), .B(n20610), .Z(n14910) );
  XNOR U20030 ( .A(n20611), .B(n16123), .Z(n10133) );
  XOR U20031 ( .A(n20612), .B(n17800), .Z(n16123) );
  AND U20032 ( .A(n13574), .B(n13194), .Z(n20611) );
  XOR U20033 ( .A(n17258), .B(n20613), .Z(n13194) );
  XOR U20034 ( .A(n20614), .B(n20067), .Z(n17258) );
  XOR U20035 ( .A(n20615), .B(n20616), .Z(n20067) );
  XOR U20036 ( .A(n19325), .B(n15203), .Z(n20616) );
  XOR U20037 ( .A(n20617), .B(n19813), .Z(n15203) );
  AND U20038 ( .A(n19939), .B(n19938), .Z(n20617) );
  XNOR U20039 ( .A(n20618), .B(n19803), .Z(n19325) );
  AND U20040 ( .A(n19942), .B(n20619), .Z(n20618) );
  XNOR U20041 ( .A(n20167), .B(n20620), .Z(n20615) );
  XNOR U20042 ( .A(n18461), .B(n18889), .Z(n20620) );
  XNOR U20043 ( .A(n20621), .B(n19807), .Z(n18889) );
  AND U20044 ( .A(n19947), .B(n19946), .Z(n20621) );
  XNOR U20045 ( .A(n20622), .B(n19818), .Z(n18461) );
  AND U20046 ( .A(n20071), .B(n20070), .Z(n20622) );
  XNOR U20047 ( .A(n20623), .B(n20624), .Z(n20167) );
  XOR U20048 ( .A(n20625), .B(n20626), .Z(n13574) );
  XNOR U20049 ( .A(n11755), .B(n20627), .Z(n20582) );
  XOR U20050 ( .A(n11010), .B(n11157), .Z(n20627) );
  XNOR U20051 ( .A(n20628), .B(n18998), .Z(n11157) );
  IV U20052 ( .A(n16117), .Z(n18998) );
  XNOR U20053 ( .A(n20629), .B(n18018), .Z(n16117) );
  ANDN U20054 ( .B(n13577), .A(n12517), .Z(n20628) );
  XNOR U20055 ( .A(n20630), .B(n17218), .Z(n12517) );
  XNOR U20056 ( .A(n20631), .B(n15217), .Z(n13577) );
  XNOR U20057 ( .A(n20632), .B(n20633), .Z(n19688) );
  XOR U20058 ( .A(n18535), .B(n20634), .Z(n20633) );
  XNOR U20059 ( .A(n20635), .B(n20636), .Z(n18535) );
  ANDN U20060 ( .B(n19098), .A(n19099), .Z(n20635) );
  XOR U20061 ( .A(n18613), .B(n20637), .Z(n20632) );
  XOR U20062 ( .A(n19383), .B(n18398), .Z(n20637) );
  XNOR U20063 ( .A(n20638), .B(n20639), .Z(n18398) );
  ANDN U20064 ( .B(n19102), .A(n19103), .Z(n20638) );
  XNOR U20065 ( .A(n20640), .B(n20641), .Z(n19383) );
  ANDN U20066 ( .B(n19092), .A(n19094), .Z(n20640) );
  XNOR U20067 ( .A(n20642), .B(n20643), .Z(n18613) );
  ANDN U20068 ( .B(n19691), .A(n19692), .Z(n20642) );
  XNOR U20069 ( .A(n20644), .B(n20645), .Z(n19744) );
  XOR U20070 ( .A(n17930), .B(n16015), .Z(n20645) );
  XOR U20071 ( .A(n20646), .B(n20647), .Z(n16015) );
  AND U20072 ( .A(n20648), .B(n20649), .Z(n20646) );
  XOR U20073 ( .A(n20650), .B(n20651), .Z(n17930) );
  XOR U20074 ( .A(n20578), .B(n20654), .Z(n20644) );
  XOR U20075 ( .A(n17292), .B(n16673), .Z(n20654) );
  XNOR U20076 ( .A(n20655), .B(n20656), .Z(n16673) );
  AND U20077 ( .A(n20657), .B(n20658), .Z(n20655) );
  XNOR U20078 ( .A(n20659), .B(n20660), .Z(n17292) );
  NOR U20079 ( .A(n20661), .B(n20662), .Z(n20659) );
  XNOR U20080 ( .A(n20663), .B(n20664), .Z(n20578) );
  NOR U20081 ( .A(n20665), .B(n20666), .Z(n20663) );
  XOR U20082 ( .A(n20667), .B(n16121), .Z(n11010) );
  XOR U20083 ( .A(n20668), .B(n17039), .Z(n16121) );
  XNOR U20084 ( .A(n19237), .B(n20669), .Z(n17039) );
  XOR U20085 ( .A(n20670), .B(n20671), .Z(n19237) );
  XNOR U20086 ( .A(n20672), .B(n18709), .Z(n20671) );
  XNOR U20087 ( .A(n20673), .B(n20674), .Z(n18709) );
  ANDN U20088 ( .B(n20675), .A(n20676), .Z(n20673) );
  XNOR U20089 ( .A(n17225), .B(n20677), .Z(n20670) );
  XNOR U20090 ( .A(n20678), .B(n17030), .Z(n20677) );
  XNOR U20091 ( .A(n20679), .B(n20680), .Z(n17030) );
  ANDN U20092 ( .B(n20681), .A(n20682), .Z(n20679) );
  XNOR U20093 ( .A(n20683), .B(n20684), .Z(n17225) );
  NOR U20094 ( .A(n20685), .B(n20686), .Z(n20683) );
  AND U20095 ( .A(n13579), .B(n12513), .Z(n20667) );
  XOR U20096 ( .A(n20379), .B(n17786), .Z(n12513) );
  IV U20097 ( .A(n17522), .Z(n17786) );
  XNOR U20098 ( .A(n20689), .B(n20126), .Z(n20379) );
  NOR U20099 ( .A(n18777), .B(n18775), .Z(n20689) );
  XNOR U20100 ( .A(n20179), .B(n17121), .Z(n13579) );
  XNOR U20101 ( .A(n20690), .B(n20691), .Z(n19798) );
  XNOR U20102 ( .A(n20692), .B(n20693), .Z(n20691) );
  XOR U20103 ( .A(n17943), .B(n20694), .Z(n20690) );
  XOR U20104 ( .A(n19262), .B(n16319), .Z(n20694) );
  XNOR U20105 ( .A(n20695), .B(n20696), .Z(n16319) );
  NOR U20106 ( .A(n20697), .B(n20698), .Z(n20695) );
  XOR U20107 ( .A(n20699), .B(n20700), .Z(n19262) );
  ANDN U20108 ( .B(n20178), .A(n20176), .Z(n20699) );
  XOR U20109 ( .A(n20701), .B(n20702), .Z(n17943) );
  ANDN U20110 ( .B(n20184), .A(n20182), .Z(n20701) );
  XNOR U20111 ( .A(n20704), .B(n20697), .Z(n20179) );
  AND U20112 ( .A(n20698), .B(n20705), .Z(n20704) );
  XNOR U20113 ( .A(n20706), .B(n16114), .Z(n11755) );
  XOR U20114 ( .A(n20707), .B(n18352), .Z(n16114) );
  IV U20115 ( .A(n17231), .Z(n18352) );
  XOR U20116 ( .A(n20708), .B(n20709), .Z(n17231) );
  AND U20117 ( .A(n13583), .B(n16115), .Z(n20706) );
  XNOR U20118 ( .A(n20710), .B(n16555), .Z(n16115) );
  XOR U20119 ( .A(n20711), .B(n20200), .Z(n16555) );
  XNOR U20120 ( .A(n20712), .B(n20713), .Z(n20200) );
  XOR U20121 ( .A(n19952), .B(n19664), .Z(n20713) );
  XOR U20122 ( .A(n20714), .B(n20715), .Z(n19664) );
  ANDN U20123 ( .B(n20716), .A(n20717), .Z(n20714) );
  XNOR U20124 ( .A(n20718), .B(n20719), .Z(n19952) );
  ANDN U20125 ( .B(n20720), .A(n20721), .Z(n20718) );
  XNOR U20126 ( .A(n18221), .B(n20722), .Z(n20712) );
  XOR U20127 ( .A(n19980), .B(n20723), .Z(n20722) );
  XNOR U20128 ( .A(n20724), .B(n20725), .Z(n19980) );
  ANDN U20129 ( .B(n20726), .A(n20727), .Z(n20724) );
  XNOR U20130 ( .A(n20728), .B(n20729), .Z(n18221) );
  AND U20131 ( .A(n20730), .B(n20731), .Z(n20728) );
  XOR U20132 ( .A(n20732), .B(n19107), .Z(n13583) );
  XNOR U20133 ( .A(n20733), .B(n17283), .Z(n16298) );
  XOR U20134 ( .A(n19835), .B(n16337), .Z(n17283) );
  IV U20135 ( .A(n20734), .Z(n16337) );
  XNOR U20136 ( .A(n20735), .B(n20736), .Z(n19835) );
  AND U20137 ( .A(n20501), .B(n20499), .Z(n20735) );
  AND U20138 ( .A(n11948), .B(n11947), .Z(n20733) );
  XNOR U20139 ( .A(n20737), .B(n17951), .Z(n11947) );
  XOR U20140 ( .A(n17959), .B(n20738), .Z(n11948) );
  XOR U20141 ( .A(n19238), .B(n20739), .Z(n17959) );
  XOR U20142 ( .A(n20740), .B(n20741), .Z(n19238) );
  XNOR U20143 ( .A(n19605), .B(n18783), .Z(n20741) );
  XOR U20144 ( .A(n20742), .B(n20743), .Z(n18783) );
  AND U20145 ( .A(n20744), .B(n20745), .Z(n20742) );
  XOR U20146 ( .A(n20746), .B(n20747), .Z(n19605) );
  AND U20147 ( .A(n20748), .B(n20749), .Z(n20746) );
  XNOR U20148 ( .A(n20750), .B(n20751), .Z(n20740) );
  XOR U20149 ( .A(n18235), .B(n19258), .Z(n20751) );
  XOR U20150 ( .A(n20752), .B(n20753), .Z(n19258) );
  AND U20151 ( .A(n20754), .B(n20755), .Z(n20752) );
  XOR U20152 ( .A(n20756), .B(n20757), .Z(n18235) );
  ANDN U20153 ( .B(n20758), .A(n19273), .Z(n20756) );
  XOR U20154 ( .A(n2558), .B(n20759), .Z(n19658) );
  XOR U20155 ( .A(n3483), .B(n9256), .Z(n20759) );
  XOR U20156 ( .A(n20760), .B(n6627), .Z(n9256) );
  IV U20157 ( .A(n9275), .Z(n6627) );
  XNOR U20158 ( .A(n12305), .B(n10473), .Z(n9275) );
  XNOR U20159 ( .A(n13695), .B(n15117), .Z(n10473) );
  XNOR U20160 ( .A(n20761), .B(n20762), .Z(n15117) );
  XNOR U20161 ( .A(n10769), .B(n11901), .Z(n20762) );
  XOR U20162 ( .A(n20763), .B(n16900), .Z(n11901) );
  IV U20163 ( .A(n14808), .Z(n16900) );
  XOR U20164 ( .A(n18338), .B(n20764), .Z(n14808) );
  ANDN U20165 ( .B(n15613), .A(n14263), .Z(n20763) );
  XNOR U20166 ( .A(n19916), .B(n17869), .Z(n14263) );
  XOR U20167 ( .A(n19905), .B(n20765), .Z(n17869) );
  XOR U20168 ( .A(n20766), .B(n20767), .Z(n19905) );
  XNOR U20169 ( .A(n20768), .B(n20769), .Z(n20767) );
  XOR U20170 ( .A(n20770), .B(n20771), .Z(n20766) );
  XOR U20171 ( .A(n17994), .B(n18225), .Z(n20771) );
  XOR U20172 ( .A(n20772), .B(n20503), .Z(n18225) );
  XOR U20173 ( .A(n20774), .B(n20511), .Z(n17994) );
  ANDN U20174 ( .B(n20775), .A(n20776), .Z(n20774) );
  XOR U20175 ( .A(n20777), .B(n20778), .Z(n19916) );
  ANDN U20176 ( .B(n19860), .A(n19861), .Z(n20777) );
  XNOR U20177 ( .A(n18464), .B(n20779), .Z(n15613) );
  XNOR U20178 ( .A(n20780), .B(n14815), .Z(n10769) );
  XOR U20179 ( .A(n20781), .B(n16476), .Z(n14815) );
  AND U20180 ( .A(n15617), .B(n15618), .Z(n20780) );
  XOR U20181 ( .A(n20782), .B(n16830), .Z(n15618) );
  XNOR U20182 ( .A(n20536), .B(n17485), .Z(n15617) );
  IV U20183 ( .A(n20783), .Z(n17485) );
  XNOR U20184 ( .A(n20784), .B(n20785), .Z(n20536) );
  AND U20185 ( .A(n20786), .B(n20787), .Z(n20784) );
  XNOR U20186 ( .A(n9674), .B(n20788), .Z(n20761) );
  XOR U20187 ( .A(n9218), .B(n11262), .Z(n20788) );
  XNOR U20188 ( .A(n20789), .B(n14811), .Z(n11262) );
  XOR U20189 ( .A(n20790), .B(n19932), .Z(n14811) );
  AND U20190 ( .A(n14268), .B(n15621), .Z(n20789) );
  XNOR U20191 ( .A(n20791), .B(n20792), .Z(n15621) );
  XNOR U20192 ( .A(n20793), .B(n18215), .Z(n14268) );
  XNOR U20193 ( .A(n20794), .B(n14806), .Z(n9218) );
  XOR U20194 ( .A(n20795), .B(n16041), .Z(n14806) );
  XNOR U20195 ( .A(n20796), .B(n20797), .Z(n18885) );
  XNOR U20196 ( .A(n20798), .B(n20799), .Z(n20797) );
  XOR U20197 ( .A(n20800), .B(n20801), .Z(n20796) );
  XNOR U20198 ( .A(n20802), .B(n17238), .Z(n20801) );
  XNOR U20199 ( .A(n20803), .B(n20804), .Z(n17238) );
  ANDN U20200 ( .B(n20805), .A(n20806), .Z(n20803) );
  XOR U20201 ( .A(n17223), .B(n20808), .Z(n15625) );
  XOR U20202 ( .A(n20809), .B(n18985), .Z(n17223) );
  XOR U20203 ( .A(n20810), .B(n20811), .Z(n18985) );
  XOR U20204 ( .A(n17376), .B(n20812), .Z(n20811) );
  XNOR U20205 ( .A(n20813), .B(n20814), .Z(n17376) );
  XOR U20206 ( .A(n15207), .B(n20817), .Z(n20810) );
  XOR U20207 ( .A(n20818), .B(n18525), .Z(n20817) );
  XNOR U20208 ( .A(n20819), .B(n20820), .Z(n18525) );
  ANDN U20209 ( .B(n20821), .A(n20822), .Z(n20819) );
  XNOR U20210 ( .A(n20823), .B(n20824), .Z(n15207) );
  AND U20211 ( .A(n20825), .B(n20826), .Z(n20823) );
  XOR U20212 ( .A(n20827), .B(n18796), .Z(n14272) );
  IV U20213 ( .A(n18172), .Z(n18796) );
  XOR U20214 ( .A(n20828), .B(n18631), .Z(n18172) );
  XOR U20215 ( .A(n20829), .B(n20830), .Z(n18631) );
  XOR U20216 ( .A(n18624), .B(n18731), .Z(n20830) );
  XOR U20217 ( .A(n20831), .B(n20832), .Z(n18731) );
  ANDN U20218 ( .B(n19755), .A(n19753), .Z(n20831) );
  XNOR U20219 ( .A(n20833), .B(n20834), .Z(n18624) );
  ANDN U20220 ( .B(n19764), .A(n19762), .Z(n20833) );
  XNOR U20221 ( .A(n18695), .B(n20835), .Z(n20829) );
  XOR U20222 ( .A(n20836), .B(n18760), .Z(n20835) );
  XNOR U20223 ( .A(n20837), .B(n20838), .Z(n18760) );
  ANDN U20224 ( .B(n19751), .A(n19749), .Z(n20837) );
  XOR U20225 ( .A(n20839), .B(n20840), .Z(n18695) );
  ANDN U20226 ( .B(n19760), .A(n19758), .Z(n20839) );
  XOR U20227 ( .A(n20841), .B(n14819), .Z(n9674) );
  XOR U20228 ( .A(n20842), .B(n19741), .Z(n14819) );
  XOR U20229 ( .A(n20843), .B(n20844), .Z(n19741) );
  ANDN U20230 ( .B(n15629), .A(n14276), .Z(n20841) );
  XNOR U20231 ( .A(n20845), .B(n19020), .Z(n14276) );
  XNOR U20232 ( .A(n20846), .B(n17928), .Z(n15629) );
  XOR U20233 ( .A(n20847), .B(n20848), .Z(n13695) );
  XNOR U20234 ( .A(n16880), .B(n12441), .Z(n20848) );
  XOR U20235 ( .A(n20849), .B(n15746), .Z(n12441) );
  XOR U20236 ( .A(n20850), .B(n18990), .Z(n15746) );
  AND U20237 ( .A(n12309), .B(n16891), .Z(n20849) );
  XOR U20238 ( .A(n17411), .B(n20851), .Z(n16891) );
  IV U20239 ( .A(n19150), .Z(n17411) );
  XNOR U20240 ( .A(n19456), .B(n20852), .Z(n19150) );
  XOR U20241 ( .A(n20853), .B(n20854), .Z(n19456) );
  XNOR U20242 ( .A(n16104), .B(n17593), .Z(n20854) );
  XOR U20243 ( .A(n20855), .B(n20856), .Z(n17593) );
  ANDN U20244 ( .B(n20857), .A(n20858), .Z(n20855) );
  XOR U20245 ( .A(n20859), .B(n20860), .Z(n16104) );
  ANDN U20246 ( .B(n20861), .A(n20862), .Z(n20859) );
  XNOR U20247 ( .A(n15221), .B(n20863), .Z(n20853) );
  XNOR U20248 ( .A(n17526), .B(n18390), .Z(n20863) );
  XNOR U20249 ( .A(n20864), .B(n20865), .Z(n18390) );
  AND U20250 ( .A(n20866), .B(n20867), .Z(n20864) );
  XNOR U20251 ( .A(n20868), .B(n20869), .Z(n17526) );
  ANDN U20252 ( .B(n20870), .A(n20871), .Z(n20868) );
  XNOR U20253 ( .A(n20872), .B(n20873), .Z(n15221) );
  ANDN U20254 ( .B(n20874), .A(n20875), .Z(n20872) );
  XNOR U20255 ( .A(n20876), .B(n20798), .Z(n12309) );
  XNOR U20256 ( .A(n20877), .B(n20878), .Z(n20798) );
  AND U20257 ( .A(n20879), .B(n20880), .Z(n20877) );
  XNOR U20258 ( .A(n20881), .B(n15738), .Z(n16880) );
  XNOR U20259 ( .A(n20882), .B(n16779), .Z(n15738) );
  XOR U20260 ( .A(n20883), .B(n19743), .Z(n16779) );
  XOR U20261 ( .A(n20884), .B(n20885), .Z(n19743) );
  XOR U20262 ( .A(n17136), .B(n17582), .Z(n20885) );
  XOR U20263 ( .A(n20886), .B(n20887), .Z(n17582) );
  AND U20264 ( .A(n20888), .B(n20889), .Z(n20886) );
  XNOR U20265 ( .A(n20890), .B(n20891), .Z(n17136) );
  ANDN U20266 ( .B(n20892), .A(n20893), .Z(n20890) );
  XNOR U20267 ( .A(n20894), .B(n20895), .Z(n20884) );
  XOR U20268 ( .A(n17874), .B(n19178), .Z(n20895) );
  XNOR U20269 ( .A(n20896), .B(n20897), .Z(n19178) );
  ANDN U20270 ( .B(n20898), .A(n20899), .Z(n20896) );
  XNOR U20271 ( .A(n20900), .B(n20901), .Z(n17874) );
  ANDN U20272 ( .B(n20902), .A(n20903), .Z(n20900) );
  AND U20273 ( .A(n12300), .B(n12302), .Z(n20881) );
  XOR U20274 ( .A(n20517), .B(n19984), .Z(n12302) );
  XNOR U20275 ( .A(n20904), .B(n20905), .Z(n20517) );
  XOR U20276 ( .A(n16547), .B(n20908), .Z(n12300) );
  XNOR U20277 ( .A(n20909), .B(n20281), .Z(n16547) );
  XNOR U20278 ( .A(n20910), .B(n20911), .Z(n20281) );
  XNOR U20279 ( .A(n16680), .B(n18251), .Z(n20911) );
  XOR U20280 ( .A(n20912), .B(n20913), .Z(n18251) );
  NOR U20281 ( .A(n20914), .B(n20297), .Z(n20912) );
  XNOR U20282 ( .A(n20915), .B(n20916), .Z(n16680) );
  NOR U20283 ( .A(n20917), .B(n20301), .Z(n20915) );
  XNOR U20284 ( .A(n15986), .B(n20918), .Z(n20910) );
  XNOR U20285 ( .A(n18935), .B(n19046), .Z(n20918) );
  XNOR U20286 ( .A(n20919), .B(n20920), .Z(n19046) );
  ANDN U20287 ( .B(n20921), .A(n20288), .Z(n20919) );
  XNOR U20288 ( .A(n20922), .B(n20923), .Z(n18935) );
  NOR U20289 ( .A(n20924), .B(n20305), .Z(n20922) );
  XNOR U20290 ( .A(n20925), .B(n20926), .Z(n15986) );
  NOR U20291 ( .A(n20927), .B(n20292), .Z(n20925) );
  XOR U20292 ( .A(n12450), .B(n20928), .Z(n20847) );
  XOR U20293 ( .A(n11310), .B(n10802), .Z(n20928) );
  XNOR U20294 ( .A(n20929), .B(n15734), .Z(n10802) );
  IV U20295 ( .A(n16885), .Z(n15734) );
  XNOR U20296 ( .A(n20557), .B(n16749), .Z(n16885) );
  XOR U20297 ( .A(n20930), .B(n20931), .Z(n16749) );
  XNOR U20298 ( .A(n20932), .B(n20933), .Z(n20557) );
  ANDN U20299 ( .B(n20934), .A(n20935), .Z(n20932) );
  XNOR U20300 ( .A(n20936), .B(n15741), .Z(n11310) );
  XOR U20301 ( .A(n18181), .B(n20937), .Z(n15741) );
  AND U20302 ( .A(n15229), .B(n15231), .Z(n20936) );
  XOR U20303 ( .A(n20938), .B(n16523), .Z(n15231) );
  IV U20304 ( .A(n18489), .Z(n16523) );
  XOR U20305 ( .A(n20939), .B(n20940), .Z(n18489) );
  XNOR U20306 ( .A(n18464), .B(n20941), .Z(n15229) );
  XNOR U20307 ( .A(n20942), .B(n15731), .Z(n12450) );
  XOR U20308 ( .A(n17993), .B(n20770), .Z(n15731) );
  ANDN U20309 ( .B(n20944), .A(n19837), .Z(n20943) );
  AND U20310 ( .A(n12379), .B(n12378), .Z(n20942) );
  XNOR U20311 ( .A(n20946), .B(n17472), .Z(n12379) );
  XNOR U20312 ( .A(n20947), .B(n20948), .Z(n20463) );
  XOR U20313 ( .A(n18483), .B(n18410), .Z(n20948) );
  XOR U20314 ( .A(n20949), .B(n20950), .Z(n18410) );
  AND U20315 ( .A(n20951), .B(n20952), .Z(n20949) );
  XNOR U20316 ( .A(n20953), .B(n20954), .Z(n18483) );
  NOR U20317 ( .A(n20955), .B(n20956), .Z(n20953) );
  XOR U20318 ( .A(n18378), .B(n20957), .Z(n20947) );
  XOR U20319 ( .A(n20958), .B(n20959), .Z(n20957) );
  XNOR U20320 ( .A(n20960), .B(n20961), .Z(n18378) );
  XOR U20321 ( .A(n20964), .B(n20965), .Z(n20514) );
  XNOR U20322 ( .A(n20966), .B(n17276), .Z(n20965) );
  XNOR U20323 ( .A(n20967), .B(n20968), .Z(n17276) );
  NOR U20324 ( .A(n20969), .B(n20970), .Z(n20967) );
  XOR U20325 ( .A(n18115), .B(n20971), .Z(n20964) );
  XOR U20326 ( .A(n18216), .B(n20972), .Z(n20971) );
  XNOR U20327 ( .A(n20973), .B(n20974), .Z(n18216) );
  ANDN U20328 ( .B(n20975), .A(n20976), .Z(n20973) );
  XNOR U20329 ( .A(n20977), .B(n20978), .Z(n18115) );
  AND U20330 ( .A(n20979), .B(n20980), .Z(n20977) );
  XNOR U20331 ( .A(n20981), .B(n16886), .Z(n12305) );
  XOR U20332 ( .A(n19271), .B(n18730), .Z(n16886) );
  XOR U20333 ( .A(n20982), .B(n20749), .Z(n19271) );
  IV U20334 ( .A(n20983), .Z(n20749) );
  NOR U20335 ( .A(n20984), .B(n20985), .Z(n20982) );
  ANDN U20336 ( .B(n17073), .A(n15733), .Z(n20981) );
  XNOR U20337 ( .A(n19471), .B(n18113), .Z(n15733) );
  XOR U20338 ( .A(n20986), .B(n20317), .Z(n19471) );
  ANDN U20339 ( .B(n20458), .A(n20459), .Z(n20986) );
  XOR U20340 ( .A(n20987), .B(n16062), .Z(n17073) );
  XNOR U20341 ( .A(n20988), .B(n20989), .Z(n19560) );
  XOR U20342 ( .A(n19059), .B(n19736), .Z(n20989) );
  XOR U20343 ( .A(n20990), .B(n20991), .Z(n19736) );
  ANDN U20344 ( .B(n20992), .A(n20993), .Z(n20990) );
  XNOR U20345 ( .A(n20994), .B(n20995), .Z(n19059) );
  AND U20346 ( .A(n20996), .B(n20997), .Z(n20994) );
  XNOR U20347 ( .A(n15959), .B(n20998), .Z(n20988) );
  XOR U20348 ( .A(n17966), .B(n17631), .Z(n20998) );
  XNOR U20349 ( .A(n20999), .B(n21000), .Z(n17631) );
  ANDN U20350 ( .B(n21001), .A(n21002), .Z(n20999) );
  XNOR U20351 ( .A(n21003), .B(n21004), .Z(n17966) );
  NOR U20352 ( .A(n21005), .B(n21006), .Z(n21003) );
  XOR U20353 ( .A(n21007), .B(n21008), .Z(n15959) );
  ANDN U20354 ( .B(n21009), .A(n21010), .Z(n21007) );
  XOR U20355 ( .A(n21011), .B(n21012), .Z(n20709) );
  XNOR U20356 ( .A(n19402), .B(n19931), .Z(n21012) );
  XOR U20357 ( .A(n21013), .B(n21014), .Z(n19931) );
  ANDN U20358 ( .B(n21015), .A(n21016), .Z(n21013) );
  XOR U20359 ( .A(n21017), .B(n21018), .Z(n19402) );
  ANDN U20360 ( .B(n21019), .A(n21020), .Z(n21017) );
  XNOR U20361 ( .A(n21021), .B(n21022), .Z(n21011) );
  XOR U20362 ( .A(n19444), .B(n20790), .Z(n21022) );
  XOR U20363 ( .A(n21023), .B(n21024), .Z(n20790) );
  ANDN U20364 ( .B(n21025), .A(n21026), .Z(n21023) );
  XOR U20365 ( .A(n21027), .B(n21028), .Z(n19444) );
  ANDN U20366 ( .B(n21029), .A(n21030), .Z(n21027) );
  ANDN U20367 ( .B(n9200), .A(n7071), .Z(n20760) );
  XNOR U20368 ( .A(n19628), .B(n12645), .Z(n7071) );
  IV U20369 ( .A(n11875), .Z(n12645) );
  XNOR U20370 ( .A(n21031), .B(n21032), .Z(n12319) );
  XNOR U20371 ( .A(n12345), .B(n9703), .Z(n21032) );
  XNOR U20372 ( .A(n21033), .B(n15105), .Z(n9703) );
  XNOR U20373 ( .A(n20531), .B(n20783), .Z(n15105) );
  XOR U20374 ( .A(n21034), .B(n20930), .Z(n20783) );
  XNOR U20375 ( .A(n21035), .B(n21036), .Z(n20930) );
  XOR U20376 ( .A(n17015), .B(n17620), .Z(n21036) );
  XOR U20377 ( .A(n21037), .B(n21038), .Z(n17620) );
  ANDN U20378 ( .B(n20933), .A(n20934), .Z(n21037) );
  XNOR U20379 ( .A(n21039), .B(n21040), .Z(n17015) );
  ANDN U20380 ( .B(n20553), .A(n20554), .Z(n21039) );
  XOR U20381 ( .A(n15212), .B(n21041), .Z(n21035) );
  XNOR U20382 ( .A(n19180), .B(n19002), .Z(n21041) );
  XNOR U20383 ( .A(n21042), .B(n21043), .Z(n19002) );
  ANDN U20384 ( .B(n20549), .A(n20550), .Z(n21042) );
  XNOR U20385 ( .A(n21044), .B(n21045), .Z(n19180) );
  ANDN U20386 ( .B(n20559), .A(n20560), .Z(n21044) );
  XNOR U20387 ( .A(n21046), .B(n21047), .Z(n15212) );
  AND U20388 ( .A(n20563), .B(n21048), .Z(n21046) );
  XOR U20389 ( .A(n21049), .B(n21050), .Z(n20531) );
  AND U20390 ( .A(n21051), .B(n21052), .Z(n21049) );
  AND U20391 ( .A(n16631), .B(n15104), .Z(n21033) );
  XOR U20392 ( .A(n21053), .B(n18242), .Z(n15104) );
  IV U20393 ( .A(n16031), .Z(n18242) );
  XOR U20394 ( .A(n21054), .B(n19167), .Z(n16031) );
  XNOR U20395 ( .A(n21055), .B(n21056), .Z(n19167) );
  XNOR U20396 ( .A(n18857), .B(n18001), .Z(n21056) );
  XOR U20397 ( .A(n21057), .B(n21058), .Z(n18001) );
  ANDN U20398 ( .B(n21059), .A(n21060), .Z(n21057) );
  XNOR U20399 ( .A(n21061), .B(n21062), .Z(n18857) );
  ANDN U20400 ( .B(n21063), .A(n21064), .Z(n21061) );
  XNOR U20401 ( .A(n18793), .B(n21065), .Z(n21055) );
  XOR U20402 ( .A(n21066), .B(n21067), .Z(n21065) );
  XNOR U20403 ( .A(n21068), .B(n21069), .Z(n18793) );
  ANDN U20404 ( .B(n21070), .A(n21071), .Z(n21068) );
  XNOR U20405 ( .A(n21072), .B(n15115), .Z(n12345) );
  NOR U20406 ( .A(n15114), .B(n16626), .Z(n21072) );
  XOR U20407 ( .A(n21073), .B(n18192), .Z(n15114) );
  XOR U20408 ( .A(n21074), .B(n21075), .Z(n18192) );
  XNOR U20409 ( .A(n14960), .B(n21076), .Z(n21031) );
  XNOR U20410 ( .A(n14565), .B(n9815), .Z(n21076) );
  XNOR U20411 ( .A(n21077), .B(n19417), .Z(n9815) );
  XNOR U20412 ( .A(n19570), .B(n16256), .Z(n19417) );
  IV U20413 ( .A(n19787), .Z(n16256) );
  XOR U20414 ( .A(n21078), .B(n19738), .Z(n19787) );
  XNOR U20415 ( .A(n21079), .B(n21080), .Z(n19738) );
  XNOR U20416 ( .A(n17187), .B(n20018), .Z(n21080) );
  XOR U20417 ( .A(n21081), .B(n21082), .Z(n20018) );
  ANDN U20418 ( .B(n19572), .A(n19573), .Z(n21081) );
  XNOR U20419 ( .A(n21083), .B(n21084), .Z(n17187) );
  ANDN U20420 ( .B(n19565), .A(n19567), .Z(n21083) );
  XOR U20421 ( .A(n17907), .B(n21085), .Z(n21079) );
  XOR U20422 ( .A(n18431), .B(n19899), .Z(n21085) );
  XOR U20423 ( .A(n21086), .B(n21087), .Z(n19899) );
  AND U20424 ( .A(n19789), .B(n19790), .Z(n21086) );
  XNOR U20425 ( .A(n21088), .B(n21089), .Z(n18431) );
  ANDN U20426 ( .B(n21090), .A(n21091), .Z(n21088) );
  XOR U20427 ( .A(n21092), .B(n21093), .Z(n17907) );
  AND U20428 ( .A(n19967), .B(n19965), .Z(n21092) );
  XNOR U20429 ( .A(n21094), .B(n21090), .Z(n19570) );
  ANDN U20430 ( .B(n21091), .A(n21095), .Z(n21094) );
  ANDN U20431 ( .B(n16633), .A(n16634), .Z(n21077) );
  XNOR U20432 ( .A(n21096), .B(n15129), .Z(n16633) );
  XNOR U20433 ( .A(n21097), .B(n19775), .Z(n15129) );
  XNOR U20434 ( .A(n21098), .B(n21099), .Z(n19775) );
  XOR U20435 ( .A(n19138), .B(n18438), .Z(n21099) );
  XOR U20436 ( .A(n21100), .B(n21101), .Z(n18438) );
  ANDN U20437 ( .B(n21102), .A(n21103), .Z(n21100) );
  XOR U20438 ( .A(n21104), .B(n21105), .Z(n19138) );
  ANDN U20439 ( .B(n21106), .A(n21107), .Z(n21104) );
  XOR U20440 ( .A(n15335), .B(n21108), .Z(n21098) );
  XNOR U20441 ( .A(n18751), .B(n18810), .Z(n21108) );
  XNOR U20442 ( .A(n21109), .B(n21110), .Z(n18810) );
  AND U20443 ( .A(n21111), .B(n21112), .Z(n21109) );
  XNOR U20444 ( .A(n21113), .B(n21114), .Z(n18751) );
  XNOR U20445 ( .A(n21117), .B(n21118), .Z(n15335) );
  XNOR U20446 ( .A(n21121), .B(n15111), .Z(n14565) );
  XOR U20447 ( .A(n21122), .B(n17243), .Z(n15111) );
  IV U20448 ( .A(n21123), .Z(n17243) );
  AND U20449 ( .A(n16623), .B(n15110), .Z(n21121) );
  XOR U20450 ( .A(n21124), .B(n17069), .Z(n15110) );
  XOR U20451 ( .A(n21125), .B(n21126), .Z(n17069) );
  XNOR U20452 ( .A(n21127), .B(n15101), .Z(n14960) );
  XNOR U20453 ( .A(n21128), .B(n17585), .Z(n15101) );
  IV U20454 ( .A(n18832), .Z(n17585) );
  AND U20455 ( .A(n16638), .B(n15100), .Z(n21127) );
  XNOR U20456 ( .A(n21131), .B(n18119), .Z(n15100) );
  XNOR U20457 ( .A(n21132), .B(n21133), .Z(n14081) );
  XNOR U20458 ( .A(n9192), .B(n12721), .Z(n21133) );
  XNOR U20459 ( .A(n21134), .B(n14651), .Z(n12721) );
  XNOR U20460 ( .A(n18156), .B(n21135), .Z(n14651) );
  AND U20461 ( .A(n17170), .B(n21136), .Z(n21134) );
  XOR U20462 ( .A(n21137), .B(n14662), .Z(n9192) );
  XOR U20463 ( .A(n18637), .B(n21138), .Z(n14662) );
  XOR U20464 ( .A(n20843), .B(n20939), .Z(n18637) );
  XOR U20465 ( .A(n21139), .B(n21140), .Z(n20939) );
  XNOR U20466 ( .A(n21141), .B(n17482), .Z(n21140) );
  XOR U20467 ( .A(n21142), .B(n20805), .Z(n17482) );
  NOR U20468 ( .A(n21143), .B(n21144), .Z(n21142) );
  XNOR U20469 ( .A(n18357), .B(n21145), .Z(n21139) );
  XNOR U20470 ( .A(n18515), .B(n17627), .Z(n21145) );
  XOR U20471 ( .A(n21146), .B(n21147), .Z(n17627) );
  ANDN U20472 ( .B(n21148), .A(n21149), .Z(n21146) );
  XNOR U20473 ( .A(n21150), .B(n21151), .Z(n18515) );
  ANDN U20474 ( .B(n21152), .A(n21153), .Z(n21150) );
  XNOR U20475 ( .A(n21154), .B(n21155), .Z(n18357) );
  ANDN U20476 ( .B(n21156), .A(n21157), .Z(n21154) );
  XOR U20477 ( .A(n21158), .B(n21159), .Z(n20843) );
  XNOR U20478 ( .A(n20133), .B(n18836), .Z(n21159) );
  XOR U20479 ( .A(n21160), .B(n21161), .Z(n18836) );
  NOR U20480 ( .A(n21162), .B(n21163), .Z(n21160) );
  XOR U20481 ( .A(n21164), .B(n21165), .Z(n20133) );
  NOR U20482 ( .A(n21166), .B(n21167), .Z(n21164) );
  XOR U20483 ( .A(n19052), .B(n21168), .Z(n21158) );
  XOR U20484 ( .A(n18735), .B(n19038), .Z(n21168) );
  XOR U20485 ( .A(n21169), .B(n21170), .Z(n19038) );
  NOR U20486 ( .A(n21171), .B(n21172), .Z(n21169) );
  XOR U20487 ( .A(n21173), .B(n21174), .Z(n18735) );
  ANDN U20488 ( .B(n21175), .A(n21176), .Z(n21173) );
  XOR U20489 ( .A(n21177), .B(n21178), .Z(n19052) );
  NOR U20490 ( .A(n21179), .B(n21180), .Z(n21177) );
  AND U20491 ( .A(n15083), .B(n17165), .Z(n21137) );
  IV U20492 ( .A(n19634), .Z(n17165) );
  XOR U20493 ( .A(n21181), .B(n18376), .Z(n19634) );
  IV U20494 ( .A(n18406), .Z(n18376) );
  XNOR U20495 ( .A(n21182), .B(n21183), .Z(n20168) );
  XNOR U20496 ( .A(n18696), .B(n18980), .Z(n21183) );
  XOR U20497 ( .A(n21184), .B(n19808), .Z(n18980) );
  XOR U20498 ( .A(round_reg[1225]), .B(n21185), .Z(n19946) );
  XNOR U20499 ( .A(round_reg[1298]), .B(n21186), .Z(n19807) );
  XNOR U20500 ( .A(n21187), .B(n21188), .Z(n18696) );
  XNOR U20501 ( .A(round_reg[1127]), .B(n21189), .Z(n19949) );
  XNOR U20502 ( .A(n18608), .B(n21190), .Z(n21182) );
  XNOR U20503 ( .A(n19797), .B(n19609), .Z(n21190) );
  XNOR U20504 ( .A(n21191), .B(n19804), .Z(n19609) );
  AND U20505 ( .A(n19803), .B(n19941), .Z(n21191) );
  IV U20506 ( .A(n20619), .Z(n19941) );
  XOR U20507 ( .A(round_reg[1153]), .B(n21192), .Z(n20619) );
  XOR U20508 ( .A(round_reg[1581]), .B(n21193), .Z(n19803) );
  XNOR U20509 ( .A(n21194), .B(n19817), .Z(n19797) );
  ANDN U20510 ( .B(n19818), .A(n20070), .Z(n21194) );
  XOR U20511 ( .A(round_reg[1078]), .B(n21195), .Z(n20070) );
  XOR U20512 ( .A(round_reg[1455]), .B(n21196), .Z(n19818) );
  XNOR U20513 ( .A(n21197), .B(n19814), .Z(n18608) );
  ANDN U20514 ( .B(n19813), .A(n19938), .Z(n21197) );
  XOR U20515 ( .A(round_reg[985]), .B(n21198), .Z(n19938) );
  XOR U20516 ( .A(round_reg[1361]), .B(n21199), .Z(n19813) );
  XNOR U20517 ( .A(n21200), .B(n21201), .Z(n20030) );
  XNOR U20518 ( .A(n17132), .B(n19134), .Z(n21201) );
  XNOR U20519 ( .A(n21202), .B(n20221), .Z(n19134) );
  XNOR U20520 ( .A(n21204), .B(n20226), .Z(n17132) );
  NOR U20521 ( .A(n21205), .B(n20225), .Z(n21204) );
  XOR U20522 ( .A(n17429), .B(n21206), .Z(n21200) );
  XOR U20523 ( .A(n19287), .B(n17004), .Z(n21206) );
  XNOR U20524 ( .A(n21207), .B(n21208), .Z(n17004) );
  NOR U20525 ( .A(n21209), .B(n21210), .Z(n21207) );
  XNOR U20526 ( .A(n21211), .B(n20215), .Z(n19287) );
  ANDN U20527 ( .B(n20216), .A(n21212), .Z(n21211) );
  XNOR U20528 ( .A(n21213), .B(n20211), .Z(n17429) );
  ANDN U20529 ( .B(n20212), .A(n21214), .Z(n21213) );
  XNOR U20530 ( .A(n19217), .B(n21215), .Z(n15083) );
  XNOR U20531 ( .A(n15078), .B(n21216), .Z(n21132) );
  XOR U20532 ( .A(n9392), .B(n12619), .Z(n21216) );
  XNOR U20533 ( .A(n21217), .B(n14647), .Z(n12619) );
  XNOR U20534 ( .A(n21218), .B(n18707), .Z(n14647) );
  XOR U20535 ( .A(n19321), .B(n19934), .Z(n18707) );
  XNOR U20536 ( .A(n21219), .B(n21220), .Z(n19934) );
  XNOR U20537 ( .A(n21221), .B(n19602), .Z(n21220) );
  XOR U20538 ( .A(n21222), .B(n21223), .Z(n19602) );
  AND U20539 ( .A(n21224), .B(n20700), .Z(n21222) );
  XNOR U20540 ( .A(n19378), .B(n21225), .Z(n21219) );
  XOR U20541 ( .A(n20232), .B(n19336), .Z(n21225) );
  XOR U20542 ( .A(n21226), .B(n20187), .Z(n19336) );
  XNOR U20543 ( .A(n21229), .B(n20183), .Z(n20232) );
  ANDN U20544 ( .B(n20702), .A(n21230), .Z(n21229) );
  XNOR U20545 ( .A(n21231), .B(n20174), .Z(n19378) );
  ANDN U20546 ( .B(n21232), .A(n21233), .Z(n21231) );
  XOR U20547 ( .A(n21234), .B(n21235), .Z(n19321) );
  XOR U20548 ( .A(n15828), .B(n19141), .Z(n21235) );
  XNOR U20549 ( .A(n21236), .B(n21237), .Z(n19141) );
  AND U20550 ( .A(n21238), .B(n21239), .Z(n21236) );
  XNOR U20551 ( .A(n21240), .B(n21241), .Z(n15828) );
  ANDN U20552 ( .B(n21242), .A(n21243), .Z(n21240) );
  XNOR U20553 ( .A(n17888), .B(n21244), .Z(n21234) );
  XNOR U20554 ( .A(n19247), .B(n18474), .Z(n21244) );
  XOR U20555 ( .A(n21245), .B(n21246), .Z(n18474) );
  AND U20556 ( .A(n21247), .B(n21248), .Z(n21245) );
  XNOR U20557 ( .A(n21249), .B(n21250), .Z(n19247) );
  ANDN U20558 ( .B(n21251), .A(n21252), .Z(n21249) );
  XNOR U20559 ( .A(n21253), .B(n21254), .Z(n17888) );
  ANDN U20560 ( .B(n21255), .A(n21256), .Z(n21253) );
  NOR U20561 ( .A(n17173), .B(n15090), .Z(n21217) );
  XNOR U20562 ( .A(n21257), .B(n16792), .Z(n15090) );
  XOR U20563 ( .A(n21258), .B(n16983), .Z(n17173) );
  IV U20564 ( .A(n16924), .Z(n16983) );
  XNOR U20565 ( .A(n21075), .B(n21259), .Z(n16924) );
  XNOR U20566 ( .A(n21260), .B(n21261), .Z(n21075) );
  XNOR U20567 ( .A(n18408), .B(n20808), .Z(n21261) );
  XNOR U20568 ( .A(n21262), .B(n20826), .Z(n20808) );
  IV U20569 ( .A(n21263), .Z(n20826) );
  NOR U20570 ( .A(n20825), .B(n21264), .Z(n21262) );
  XNOR U20571 ( .A(n21265), .B(n21266), .Z(n18408) );
  AND U20572 ( .A(n21267), .B(n21268), .Z(n21265) );
  XOR U20573 ( .A(n20275), .B(n21269), .Z(n21260) );
  XOR U20574 ( .A(n19241), .B(n17224), .Z(n21269) );
  XNOR U20575 ( .A(n21270), .B(n20821), .Z(n17224) );
  ANDN U20576 ( .B(n20822), .A(n21271), .Z(n21270) );
  XNOR U20577 ( .A(n21272), .B(n21273), .Z(n19241) );
  ANDN U20578 ( .B(n21274), .A(n21275), .Z(n21272) );
  XOR U20579 ( .A(n21276), .B(n20816), .Z(n20275) );
  XNOR U20580 ( .A(n14657), .B(n21278), .Z(n9392) );
  XOR U20581 ( .A(n21279), .B(n21280), .Z(n21278) );
  NAND U20582 ( .A(n4509), .B(n4365), .Z(n21280) );
  AND U20583 ( .A(n4510), .B(n15691), .Z(n4365) );
  AND U20584 ( .A(n6835), .B(n6455), .Z(n4509) );
  XNOR U20585 ( .A(n19466), .B(n18113), .Z(n17161) );
  XOR U20586 ( .A(n21097), .B(n20084), .Z(n18113) );
  XOR U20587 ( .A(n21281), .B(n21282), .Z(n20084) );
  XNOR U20588 ( .A(n18720), .B(n20136), .Z(n21282) );
  XOR U20589 ( .A(n21283), .B(n21284), .Z(n20136) );
  ANDN U20590 ( .B(n21285), .A(n21286), .Z(n21283) );
  XNOR U20591 ( .A(n21287), .B(n20534), .Z(n18720) );
  XOR U20592 ( .A(n17501), .B(n21289), .Z(n21281) );
  XOR U20593 ( .A(n19982), .B(n20528), .Z(n21289) );
  XOR U20594 ( .A(n21290), .B(n21291), .Z(n20528) );
  NOR U20595 ( .A(n20540), .B(n21292), .Z(n21290) );
  AND U20596 ( .A(n21294), .B(n21295), .Z(n21293) );
  XNOR U20597 ( .A(n21296), .B(n20786), .Z(n17501) );
  XOR U20598 ( .A(n21298), .B(n21299), .Z(n21097) );
  XNOR U20599 ( .A(n19530), .B(n16784), .Z(n21299) );
  XOR U20600 ( .A(n21300), .B(n21301), .Z(n16784) );
  XOR U20601 ( .A(n21303), .B(n21304), .Z(n19530) );
  ANDN U20602 ( .B(n21305), .A(n19479), .Z(n21303) );
  XOR U20603 ( .A(round_reg[461]), .B(n21306), .Z(n19479) );
  XOR U20604 ( .A(n19719), .B(n21307), .Z(n21298) );
  XOR U20605 ( .A(n17964), .B(n19654), .Z(n21307) );
  XOR U20606 ( .A(n21308), .B(n20318), .Z(n19654) );
  XOR U20607 ( .A(round_reg[559]), .B(n21309), .Z(n20458) );
  XOR U20608 ( .A(round_reg[921]), .B(n21310), .Z(n20317) );
  XOR U20609 ( .A(n21311), .B(n19730), .Z(n17964) );
  NOR U20610 ( .A(n19468), .B(n19469), .Z(n21311) );
  XOR U20611 ( .A(round_reg[627]), .B(n21312), .Z(n19469) );
  XOR U20612 ( .A(round_reg[693]), .B(n21313), .Z(n19468) );
  XOR U20613 ( .A(n21314), .B(n21315), .Z(n19719) );
  NOR U20614 ( .A(n19474), .B(n19475), .Z(n21314) );
  XOR U20615 ( .A(round_reg[391]), .B(n21316), .Z(n19475) );
  XOR U20616 ( .A(n21317), .B(n21302), .Z(n19466) );
  ANDN U20617 ( .B(n20454), .A(n20455), .Z(n21317) );
  XOR U20618 ( .A(round_reg[340]), .B(n21318), .Z(n20454) );
  XOR U20619 ( .A(n21319), .B(n18757), .Z(n15095) );
  XNOR U20620 ( .A(n21320), .B(n18180), .Z(n14657) );
  XOR U20621 ( .A(n21323), .B(n15086), .Z(n15078) );
  XOR U20622 ( .A(n17083), .B(n21324), .Z(n15086) );
  IV U20623 ( .A(n18588), .Z(n17083) );
  XOR U20624 ( .A(n18947), .B(n20703), .Z(n18588) );
  XNOR U20625 ( .A(n21325), .B(n21326), .Z(n20703) );
  XNOR U20626 ( .A(n17904), .B(n18263), .Z(n21326) );
  XOR U20627 ( .A(n21327), .B(n21243), .Z(n18263) );
  ANDN U20628 ( .B(n21328), .A(n21329), .Z(n21327) );
  XNOR U20629 ( .A(n21330), .B(n21247), .Z(n17904) );
  ANDN U20630 ( .B(n21331), .A(n21332), .Z(n21330) );
  XNOR U20631 ( .A(n15324), .B(n21333), .Z(n21325) );
  XOR U20632 ( .A(n21334), .B(n16917), .Z(n21333) );
  XNOR U20633 ( .A(n21335), .B(n21239), .Z(n16917) );
  ANDN U20634 ( .B(n21336), .A(n21337), .Z(n21335) );
  XNOR U20635 ( .A(n21338), .B(n21251), .Z(n15324) );
  ANDN U20636 ( .B(n21339), .A(n21340), .Z(n21338) );
  XOR U20637 ( .A(n21341), .B(n21342), .Z(n18947) );
  XNOR U20638 ( .A(n16611), .B(n17834), .Z(n21342) );
  XNOR U20639 ( .A(n21343), .B(n21344), .Z(n17834) );
  AND U20640 ( .A(n21345), .B(n21346), .Z(n21343) );
  XNOR U20641 ( .A(n21347), .B(n21348), .Z(n16611) );
  ANDN U20642 ( .B(n21349), .A(n21350), .Z(n21347) );
  XNOR U20643 ( .A(n21351), .B(n21352), .Z(n21341) );
  XNOR U20644 ( .A(n18308), .B(n16824), .Z(n21352) );
  XOR U20645 ( .A(n21353), .B(n21354), .Z(n16824) );
  ANDN U20646 ( .B(n21355), .A(n21356), .Z(n21353) );
  XNOR U20647 ( .A(n21357), .B(n21358), .Z(n18308) );
  ANDN U20648 ( .B(n17177), .A(n15087), .Z(n21323) );
  XOR U20649 ( .A(n21361), .B(n20234), .Z(n15087) );
  XNOR U20650 ( .A(n21362), .B(n21363), .Z(n20234) );
  XOR U20651 ( .A(n21364), .B(n18279), .Z(n17177) );
  XNOR U20652 ( .A(n20844), .B(n20242), .Z(n18279) );
  XNOR U20653 ( .A(n21365), .B(n21366), .Z(n20242) );
  XNOR U20654 ( .A(n19428), .B(n20080), .Z(n21366) );
  XNOR U20655 ( .A(n21367), .B(n21368), .Z(n20080) );
  AND U20656 ( .A(n21369), .B(n21370), .Z(n21367) );
  XNOR U20657 ( .A(n21371), .B(n21372), .Z(n19428) );
  ANDN U20658 ( .B(n21373), .A(n21374), .Z(n21371) );
  XOR U20659 ( .A(n20189), .B(n21375), .Z(n21365) );
  XOR U20660 ( .A(n17679), .B(n16472), .Z(n21375) );
  XNOR U20661 ( .A(n21376), .B(n21377), .Z(n16472) );
  ANDN U20662 ( .B(n21378), .A(n21379), .Z(n21376) );
  XNOR U20663 ( .A(n21380), .B(n21381), .Z(n17679) );
  ANDN U20664 ( .B(n21382), .A(n21383), .Z(n21380) );
  XNOR U20665 ( .A(n21384), .B(n21385), .Z(n20189) );
  ANDN U20666 ( .B(n21386), .A(n21387), .Z(n21384) );
  XOR U20667 ( .A(n21388), .B(n21389), .Z(n20844) );
  XNOR U20668 ( .A(n18522), .B(n17025), .Z(n21389) );
  XNOR U20669 ( .A(n21390), .B(n21391), .Z(n17025) );
  ANDN U20670 ( .B(n21392), .A(n21393), .Z(n21390) );
  XNOR U20671 ( .A(n21394), .B(n21395), .Z(n18522) );
  ANDN U20672 ( .B(n21396), .A(n20252), .Z(n21394) );
  XOR U20673 ( .A(n21397), .B(n21398), .Z(n21388) );
  XOR U20674 ( .A(n15910), .B(n17495), .Z(n21398) );
  XOR U20675 ( .A(n21399), .B(n21400), .Z(n17495) );
  ANDN U20676 ( .B(n21401), .A(n20266), .Z(n21399) );
  XOR U20677 ( .A(n21402), .B(n21403), .Z(n15910) );
  ANDN U20678 ( .B(n21404), .A(n20256), .Z(n21402) );
  XOR U20679 ( .A(n21405), .B(n15093), .Z(n19628) );
  IV U20680 ( .A(n21136), .Z(n15093) );
  XOR U20681 ( .A(n20750), .B(n18236), .Z(n21136) );
  XNOR U20682 ( .A(n19927), .B(n21406), .Z(n18236) );
  XOR U20683 ( .A(n21407), .B(n21408), .Z(n19927) );
  XOR U20684 ( .A(n19714), .B(n16943), .Z(n21408) );
  XOR U20685 ( .A(n21409), .B(n21410), .Z(n16943) );
  ANDN U20686 ( .B(n21411), .A(n21412), .Z(n21409) );
  XNOR U20687 ( .A(n21413), .B(n21414), .Z(n19714) );
  ANDN U20688 ( .B(n21415), .A(n21416), .Z(n21413) );
  XNOR U20689 ( .A(n19395), .B(n21417), .Z(n21407) );
  XNOR U20690 ( .A(n18872), .B(n20605), .Z(n21417) );
  XOR U20691 ( .A(n21418), .B(n21419), .Z(n20605) );
  ANDN U20692 ( .B(n21420), .A(n21421), .Z(n21418) );
  XNOR U20693 ( .A(n21422), .B(n21423), .Z(n18872) );
  ANDN U20694 ( .B(n21424), .A(n21425), .Z(n21422) );
  XNOR U20695 ( .A(n21426), .B(n21427), .Z(n19395) );
  ANDN U20696 ( .B(n21428), .A(n21429), .Z(n21426) );
  XNOR U20697 ( .A(n21430), .B(n21431), .Z(n20750) );
  ANDN U20698 ( .B(n21432), .A(n19280), .Z(n21430) );
  NOR U20699 ( .A(n14650), .B(n17170), .Z(n21405) );
  XNOR U20700 ( .A(n21433), .B(n17560), .Z(n17170) );
  XNOR U20701 ( .A(n21436), .B(n19020), .Z(n14650) );
  IV U20702 ( .A(n17962), .Z(n19020) );
  XOR U20703 ( .A(n19652), .B(n20019), .Z(n17962) );
  XOR U20704 ( .A(n21437), .B(n21438), .Z(n20019) );
  XOR U20705 ( .A(n19161), .B(n21439), .Z(n21438) );
  XNOR U20706 ( .A(n21440), .B(n21441), .Z(n19161) );
  ANDN U20707 ( .B(n21442), .A(n21443), .Z(n21440) );
  XOR U20708 ( .A(n18634), .B(n21444), .Z(n21437) );
  XOR U20709 ( .A(n18388), .B(n21445), .Z(n21444) );
  XNOR U20710 ( .A(n21446), .B(n21447), .Z(n18388) );
  ANDN U20711 ( .B(n21448), .A(n21449), .Z(n21446) );
  XNOR U20712 ( .A(n21450), .B(n21451), .Z(n18634) );
  NOR U20713 ( .A(n21452), .B(n21453), .Z(n21450) );
  XOR U20714 ( .A(n21454), .B(n21455), .Z(n19652) );
  XNOR U20715 ( .A(n16797), .B(n14905), .Z(n21455) );
  XOR U20716 ( .A(n21456), .B(n21107), .Z(n14905) );
  ANDN U20717 ( .B(n21457), .A(n21458), .Z(n21456) );
  XNOR U20718 ( .A(n21459), .B(n21112), .Z(n16797) );
  IV U20719 ( .A(n21460), .Z(n21112) );
  ANDN U20720 ( .B(n21461), .A(n21462), .Z(n21459) );
  XNOR U20721 ( .A(n16351), .B(n21463), .Z(n21454) );
  XNOR U20722 ( .A(n17970), .B(n19462), .Z(n21463) );
  XNOR U20723 ( .A(n21464), .B(n21115), .Z(n19462) );
  ANDN U20724 ( .B(n21465), .A(n21466), .Z(n21464) );
  XNOR U20725 ( .A(n21467), .B(n21103), .Z(n17970) );
  ANDN U20726 ( .B(n21468), .A(n21469), .Z(n21467) );
  XNOR U20727 ( .A(n21470), .B(n21119), .Z(n16351) );
  ANDN U20728 ( .B(n21471), .A(n21472), .Z(n21470) );
  XNOR U20729 ( .A(n14895), .B(n10875), .Z(n9200) );
  XNOR U20730 ( .A(n13046), .B(n12702), .Z(n10875) );
  XNOR U20731 ( .A(n21473), .B(n21474), .Z(n12702) );
  XNOR U20732 ( .A(n12833), .B(n11738), .Z(n21474) );
  XOR U20733 ( .A(n21475), .B(n15138), .Z(n11738) );
  XNOR U20734 ( .A(n15252), .B(n21476), .Z(n15138) );
  AND U20735 ( .A(n12782), .B(n15645), .Z(n21475) );
  IV U20736 ( .A(n14892), .Z(n15645) );
  XOR U20737 ( .A(n21479), .B(n18044), .Z(n14892) );
  XOR U20738 ( .A(n21480), .B(n19708), .Z(n18044) );
  XOR U20739 ( .A(n21481), .B(n21482), .Z(n19708) );
  XNOR U20740 ( .A(n18239), .B(n16899), .Z(n21482) );
  XOR U20741 ( .A(n21483), .B(n19566), .Z(n16899) );
  NOR U20742 ( .A(n21484), .B(n21084), .Z(n21483) );
  XNOR U20743 ( .A(n21485), .B(n21095), .Z(n18239) );
  ANDN U20744 ( .B(n21486), .A(n21089), .Z(n21485) );
  XOR U20745 ( .A(n19057), .B(n21487), .Z(n21481) );
  XOR U20746 ( .A(n21488), .B(n21489), .Z(n21487) );
  XOR U20747 ( .A(n21490), .B(n19966), .Z(n19057) );
  AND U20748 ( .A(n21491), .B(n21093), .Z(n21490) );
  XOR U20749 ( .A(n21492), .B(n17455), .Z(n12782) );
  XOR U20750 ( .A(n21493), .B(n15123), .Z(n12833) );
  XOR U20751 ( .A(n15917), .B(n21494), .Z(n15123) );
  AND U20752 ( .A(n12771), .B(n15640), .Z(n21493) );
  XOR U20753 ( .A(n19364), .B(n14924), .Z(n15640) );
  XOR U20754 ( .A(n21495), .B(n20077), .Z(n14924) );
  XOR U20755 ( .A(n21496), .B(n21497), .Z(n20077) );
  XNOR U20756 ( .A(n18185), .B(n20630), .Z(n21497) );
  XNOR U20757 ( .A(n21498), .B(n21499), .Z(n20630) );
  ANDN U20758 ( .B(n21500), .A(n21028), .Z(n21498) );
  XOR U20759 ( .A(n21501), .B(n21502), .Z(n18185) );
  AND U20760 ( .A(n21503), .B(n21504), .Z(n21501) );
  XNOR U20761 ( .A(n18512), .B(n21505), .Z(n21496) );
  XOR U20762 ( .A(n21506), .B(n17217), .Z(n21505) );
  XOR U20763 ( .A(n21507), .B(n21508), .Z(n17217) );
  ANDN U20764 ( .B(n21509), .A(n21024), .Z(n21507) );
  XNOR U20765 ( .A(n21510), .B(n21511), .Z(n18512) );
  ANDN U20766 ( .B(n21512), .A(n21513), .Z(n21510) );
  XNOR U20767 ( .A(n21514), .B(n20906), .Z(n19364) );
  ANDN U20768 ( .B(n21515), .A(n21516), .Z(n21514) );
  XNOR U20769 ( .A(n21517), .B(n16603), .Z(n12771) );
  XNOR U20770 ( .A(n11871), .B(n21518), .Z(n21473) );
  XOR U20771 ( .A(n9536), .B(n10363), .Z(n21518) );
  XOR U20772 ( .A(n21519), .B(n15125), .Z(n10363) );
  XOR U20773 ( .A(n16751), .B(n20110), .Z(n15125) );
  XNOR U20774 ( .A(n21520), .B(n19882), .Z(n20110) );
  ANDN U20775 ( .B(n20576), .A(n21521), .Z(n21520) );
  AND U20776 ( .A(n15636), .B(n14797), .Z(n21519) );
  XOR U20777 ( .A(n21522), .B(n15134), .Z(n9536) );
  XNOR U20778 ( .A(n21523), .B(n15606), .Z(n15134) );
  NOR U20779 ( .A(n12775), .B(n14899), .Z(n21522) );
  XNOR U20780 ( .A(n21488), .B(n16898), .Z(n14899) );
  XNOR U20781 ( .A(n21524), .B(n19791), .Z(n21488) );
  XOR U20782 ( .A(n21526), .B(n17205), .Z(n12775) );
  IV U20783 ( .A(n21527), .Z(n17205) );
  XOR U20784 ( .A(n21528), .B(n15130), .Z(n11871) );
  XOR U20785 ( .A(n21529), .B(n16049), .Z(n15130) );
  IV U20786 ( .A(n18338), .Z(n16049) );
  XOR U20787 ( .A(n19607), .B(n20708), .Z(n18338) );
  XNOR U20788 ( .A(n21530), .B(n21531), .Z(n20708) );
  XOR U20789 ( .A(n16987), .B(n18174), .Z(n21531) );
  XOR U20790 ( .A(n21532), .B(n19372), .Z(n18174) );
  ANDN U20791 ( .B(n21533), .A(n19371), .Z(n21532) );
  XNOR U20792 ( .A(n21534), .B(n21515), .Z(n16987) );
  ANDN U20793 ( .B(n21516), .A(n20905), .Z(n21534) );
  XNOR U20794 ( .A(n17146), .B(n21535), .Z(n21530) );
  XNOR U20795 ( .A(n18025), .B(n17339), .Z(n21535) );
  XNOR U20796 ( .A(n21536), .B(n19362), .Z(n17339) );
  ANDN U20797 ( .B(n20525), .A(n19361), .Z(n21536) );
  IV U20798 ( .A(n21537), .Z(n20525) );
  XNOR U20799 ( .A(n21538), .B(n19367), .Z(n18025) );
  AND U20800 ( .A(n21539), .B(n21540), .Z(n21538) );
  XNOR U20801 ( .A(n21541), .B(n19358), .Z(n17146) );
  AND U20802 ( .A(n20519), .B(n19357), .Z(n21541) );
  XOR U20803 ( .A(n21542), .B(n21543), .Z(n19607) );
  XNOR U20804 ( .A(n18944), .B(n18744), .Z(n21543) );
  XOR U20805 ( .A(n21544), .B(n21545), .Z(n18744) );
  ANDN U20806 ( .B(n21546), .A(n21547), .Z(n21544) );
  XOR U20807 ( .A(n21548), .B(n21549), .Z(n18944) );
  NOR U20808 ( .A(n21550), .B(n20974), .Z(n21548) );
  XOR U20809 ( .A(n19351), .B(n21551), .Z(n21542) );
  XOR U20810 ( .A(n19230), .B(n19210), .Z(n21551) );
  XNOR U20811 ( .A(n21552), .B(n21553), .Z(n19210) );
  NOR U20812 ( .A(n21554), .B(n20968), .Z(n21552) );
  XNOR U20813 ( .A(n21555), .B(n21556), .Z(n19230) );
  ANDN U20814 ( .B(n21557), .A(n20978), .Z(n21555) );
  XNOR U20815 ( .A(n21558), .B(n21559), .Z(n19351) );
  NOR U20816 ( .A(n21560), .B(n21561), .Z(n21558) );
  AND U20817 ( .A(n14888), .B(n14926), .Z(n21528) );
  IV U20818 ( .A(n14890), .Z(n14926) );
  XOR U20819 ( .A(n20894), .B(n17583), .Z(n14890) );
  IV U20820 ( .A(n17137), .Z(n17583) );
  XOR U20821 ( .A(n21562), .B(n21563), .Z(n20580) );
  XOR U20822 ( .A(n21564), .B(n20036), .Z(n21563) );
  XNOR U20823 ( .A(n21565), .B(n21566), .Z(n20036) );
  AND U20824 ( .A(n20665), .B(n20664), .Z(n21565) );
  XNOR U20825 ( .A(n16063), .B(n21567), .Z(n21562) );
  XNOR U20826 ( .A(n19731), .B(n19979), .Z(n21567) );
  XOR U20827 ( .A(n21568), .B(n21569), .Z(n19979) );
  AND U20828 ( .A(n20661), .B(n20660), .Z(n21568) );
  XNOR U20829 ( .A(n21570), .B(n21571), .Z(n19731) );
  ANDN U20830 ( .B(n20647), .A(n20648), .Z(n21570) );
  XNOR U20831 ( .A(n21572), .B(n21573), .Z(n16063) );
  ANDN U20832 ( .B(n20653), .A(n20651), .Z(n21572) );
  XNOR U20833 ( .A(n21575), .B(n21576), .Z(n20894) );
  AND U20834 ( .A(n21577), .B(n21578), .Z(n21575) );
  XOR U20835 ( .A(n21579), .B(n17987), .Z(n14888) );
  XOR U20836 ( .A(n21580), .B(n21130), .Z(n17987) );
  XOR U20837 ( .A(n21581), .B(n21582), .Z(n21130) );
  XNOR U20838 ( .A(n18864), .B(n21583), .Z(n21582) );
  XNOR U20839 ( .A(n21584), .B(n21585), .Z(n18864) );
  ANDN U20840 ( .B(n21586), .A(n21368), .Z(n21584) );
  XOR U20841 ( .A(n17974), .B(n21587), .Z(n21581) );
  XOR U20842 ( .A(n17466), .B(n21588), .Z(n21587) );
  XNOR U20843 ( .A(n21589), .B(n21590), .Z(n17466) );
  ANDN U20844 ( .B(n21591), .A(n21377), .Z(n21589) );
  XNOR U20845 ( .A(n21592), .B(n21593), .Z(n17974) );
  ANDN U20846 ( .B(n21594), .A(n21381), .Z(n21592) );
  XOR U20847 ( .A(n21595), .B(n21596), .Z(n13046) );
  XOR U20848 ( .A(n10101), .B(n11795), .Z(n21596) );
  XNOR U20849 ( .A(n21597), .B(n13119), .Z(n11795) );
  XOR U20850 ( .A(n21598), .B(n19176), .Z(n16751) );
  XOR U20851 ( .A(n21599), .B(n21600), .Z(n19176) );
  XOR U20852 ( .A(n18723), .B(n18766), .Z(n21600) );
  XOR U20853 ( .A(n21601), .B(n19883), .Z(n18766) );
  XOR U20854 ( .A(round_reg[641]), .B(n21602), .Z(n19883) );
  ANDN U20855 ( .B(n21521), .A(n19882), .Z(n21601) );
  XNOR U20856 ( .A(round_reg[639]), .B(n21603), .Z(n19882) );
  XOR U20857 ( .A(n21604), .B(n19879), .Z(n18723) );
  XNOR U20858 ( .A(round_reg[719]), .B(n21605), .Z(n19879) );
  AND U20859 ( .A(n20107), .B(n20105), .Z(n21604) );
  IV U20860 ( .A(n19878), .Z(n20105) );
  XNOR U20861 ( .A(round_reg[352]), .B(n21606), .Z(n19878) );
  XNOR U20862 ( .A(n18491), .B(n21607), .Z(n21599) );
  XOR U20863 ( .A(n18021), .B(n18409), .Z(n21607) );
  XNOR U20864 ( .A(n21608), .B(n19887), .Z(n18409) );
  XOR U20865 ( .A(round_reg[829]), .B(n21609), .Z(n19887) );
  ANDN U20866 ( .B(n20113), .A(n19886), .Z(n21608) );
  XNOR U20867 ( .A(round_reg[403]), .B(n21610), .Z(n19886) );
  XOR U20868 ( .A(n21611), .B(n21612), .Z(n18021) );
  NOR U20869 ( .A(n20102), .B(n19869), .Z(n21611) );
  XNOR U20870 ( .A(round_reg[473]), .B(n21613), .Z(n19869) );
  XNOR U20871 ( .A(n21614), .B(n19874), .Z(n18491) );
  ANDN U20872 ( .B(n19873), .A(n21615), .Z(n21614) );
  XNOR U20873 ( .A(n21616), .B(n19873), .Z(n20109) );
  XNOR U20874 ( .A(round_reg[571]), .B(n21617), .Z(n19873) );
  AND U20875 ( .A(n21615), .B(n21618), .Z(n21616) );
  AND U20876 ( .A(n14903), .B(n13378), .Z(n21597) );
  XOR U20877 ( .A(n21619), .B(n19544), .Z(n13378) );
  IV U20878 ( .A(n18109), .Z(n19544) );
  XNOR U20879 ( .A(n21620), .B(n21621), .Z(n19961) );
  XNOR U20880 ( .A(n18991), .B(n20792), .Z(n21621) );
  XOR U20881 ( .A(n21622), .B(n21623), .Z(n20792) );
  ANDN U20882 ( .B(n20489), .A(n20487), .Z(n21622) );
  XNOR U20883 ( .A(n21624), .B(n21625), .Z(n18991) );
  ANDN U20884 ( .B(n20479), .A(n20480), .Z(n21624) );
  XNOR U20885 ( .A(n21626), .B(n21627), .Z(n21620) );
  XOR U20886 ( .A(n20850), .B(n20492), .Z(n21627) );
  XNOR U20887 ( .A(n21628), .B(n21629), .Z(n20492) );
  ANDN U20888 ( .B(n20470), .A(n20471), .Z(n21628) );
  XNOR U20889 ( .A(n21630), .B(n21631), .Z(n20850) );
  AND U20890 ( .A(n20483), .B(n20485), .Z(n21630) );
  XNOR U20891 ( .A(n18601), .B(n21633), .Z(n14903) );
  XNOR U20892 ( .A(n21634), .B(n12961), .Z(n10101) );
  XOR U20893 ( .A(n21635), .B(n17569), .Z(n12961) );
  IV U20894 ( .A(n17190), .Z(n17569) );
  XOR U20895 ( .A(n19119), .B(n21636), .Z(n17190) );
  XOR U20896 ( .A(n21637), .B(n21638), .Z(n19119) );
  XOR U20897 ( .A(n19392), .B(n21639), .Z(n21638) );
  XNOR U20898 ( .A(n21640), .B(n21641), .Z(n19392) );
  ANDN U20899 ( .B(n21642), .A(n21643), .Z(n21640) );
  XOR U20900 ( .A(n21644), .B(n21645), .Z(n21637) );
  XOR U20901 ( .A(n21131), .B(n18118), .Z(n21645) );
  XNOR U20902 ( .A(n21646), .B(n21647), .Z(n18118) );
  ANDN U20903 ( .B(n21648), .A(n21649), .Z(n21646) );
  XNOR U20904 ( .A(n21650), .B(n21651), .Z(n21131) );
  ANDN U20905 ( .B(n21652), .A(n21653), .Z(n21650) );
  ANDN U20906 ( .B(n13129), .A(n14907), .Z(n21634) );
  XOR U20907 ( .A(n20802), .B(n20876), .Z(n14907) );
  XOR U20908 ( .A(n21654), .B(n21655), .Z(n20802) );
  ANDN U20909 ( .B(n21155), .A(n21656), .Z(n21654) );
  IV U20910 ( .A(n14908), .Z(n13129) );
  XOR U20911 ( .A(n21657), .B(n18643), .Z(n14908) );
  XNOR U20912 ( .A(n11402), .B(n21658), .Z(n21595) );
  XOR U20913 ( .A(n15887), .B(n15580), .Z(n21658) );
  XNOR U20914 ( .A(n21659), .B(n12957), .Z(n15580) );
  XOR U20915 ( .A(n21660), .B(n16024), .Z(n12957) );
  ANDN U20916 ( .B(n14917), .A(n13125), .Z(n21659) );
  XNOR U20917 ( .A(n21661), .B(n15603), .Z(n13125) );
  XOR U20918 ( .A(n21662), .B(n20607), .Z(n15603) );
  XNOR U20919 ( .A(n21663), .B(n21664), .Z(n20607) );
  XNOR U20920 ( .A(n17558), .B(n17385), .Z(n21664) );
  XNOR U20921 ( .A(n21665), .B(n21666), .Z(n17385) );
  ANDN U20922 ( .B(n21423), .A(n21424), .Z(n21665) );
  XNOR U20923 ( .A(n21667), .B(n21668), .Z(n17558) );
  ANDN U20924 ( .B(n21419), .A(n21420), .Z(n21667) );
  XOR U20925 ( .A(n17175), .B(n21669), .Z(n21663) );
  XOR U20926 ( .A(n19136), .B(n21670), .Z(n21669) );
  XNOR U20927 ( .A(n21671), .B(n21672), .Z(n19136) );
  ANDN U20928 ( .B(n21410), .A(n21411), .Z(n21671) );
  XNOR U20929 ( .A(n21673), .B(n21674), .Z(n17175) );
  ANDN U20930 ( .B(n21414), .A(n21415), .Z(n21673) );
  XNOR U20931 ( .A(n17192), .B(n21675), .Z(n14917) );
  XOR U20932 ( .A(n19047), .B(n19769), .Z(n17192) );
  XOR U20933 ( .A(n21676), .B(n21677), .Z(n19769) );
  XNOR U20934 ( .A(n17851), .B(n19550), .Z(n21677) );
  XOR U20935 ( .A(n21678), .B(n21679), .Z(n19550) );
  ANDN U20936 ( .B(n21680), .A(n21681), .Z(n21678) );
  XOR U20937 ( .A(n21682), .B(n21683), .Z(n17851) );
  XOR U20938 ( .A(n18159), .B(n21686), .Z(n21676) );
  XOR U20939 ( .A(n17588), .B(n21687), .Z(n21686) );
  XNOR U20940 ( .A(n21688), .B(n21689), .Z(n17588) );
  AND U20941 ( .A(n21690), .B(n21691), .Z(n21688) );
  XNOR U20942 ( .A(n21692), .B(n21693), .Z(n18159) );
  XOR U20943 ( .A(n21696), .B(n21697), .Z(n19047) );
  XOR U20944 ( .A(n21698), .B(n21699), .Z(n21697) );
  XOR U20945 ( .A(n18122), .B(n21700), .Z(n21696) );
  XOR U20946 ( .A(n19393), .B(n17041), .Z(n21700) );
  XNOR U20947 ( .A(n21701), .B(n20293), .Z(n17041) );
  AND U20948 ( .A(n20927), .B(n21702), .Z(n21701) );
  XNOR U20949 ( .A(n21703), .B(n20298), .Z(n19393) );
  AND U20950 ( .A(n20914), .B(n20913), .Z(n21703) );
  IV U20951 ( .A(n21704), .Z(n20913) );
  XNOR U20952 ( .A(n21705), .B(n20290), .Z(n18122) );
  XNOR U20953 ( .A(n21706), .B(n12964), .Z(n15887) );
  XNOR U20954 ( .A(n18166), .B(n21707), .Z(n12964) );
  IV U20955 ( .A(n18403), .Z(n18166) );
  XNOR U20956 ( .A(n21708), .B(n21709), .Z(n18403) );
  AND U20957 ( .A(n14921), .B(n13362), .Z(n21706) );
  IV U20958 ( .A(n14922), .Z(n13362) );
  XOR U20959 ( .A(n20723), .B(n18222), .Z(n14922) );
  XNOR U20960 ( .A(n21054), .B(n21363), .Z(n18222) );
  XNOR U20961 ( .A(n21710), .B(n21711), .Z(n21363) );
  XOR U20962 ( .A(n18636), .B(n17919), .Z(n21711) );
  XOR U20963 ( .A(n21712), .B(n21713), .Z(n17919) );
  ANDN U20964 ( .B(n21714), .A(n20716), .Z(n21712) );
  XNOR U20965 ( .A(n21715), .B(n21716), .Z(n18636) );
  XOR U20966 ( .A(n18958), .B(n21717), .Z(n21710) );
  XOR U20967 ( .A(n17677), .B(n21718), .Z(n21717) );
  XNOR U20968 ( .A(n21719), .B(n21720), .Z(n17677) );
  ANDN U20969 ( .B(n21721), .A(n20726), .Z(n21719) );
  XNOR U20970 ( .A(n21722), .B(n21723), .Z(n18958) );
  XOR U20971 ( .A(n21724), .B(n21725), .Z(n21054) );
  XOR U20972 ( .A(n21726), .B(n17815), .Z(n21725) );
  XOR U20973 ( .A(n21727), .B(n21728), .Z(n17815) );
  AND U20974 ( .A(n21729), .B(n20008), .Z(n21727) );
  XOR U20975 ( .A(n20464), .B(n21730), .Z(n21724) );
  XOR U20976 ( .A(n18593), .B(n20073), .Z(n21730) );
  XOR U20977 ( .A(n21731), .B(n21732), .Z(n20073) );
  NOR U20978 ( .A(n21733), .B(n20004), .Z(n21731) );
  XOR U20979 ( .A(n21734), .B(n21735), .Z(n18593) );
  NOR U20980 ( .A(n21736), .B(n21737), .Z(n21734) );
  XOR U20981 ( .A(n21738), .B(n21739), .Z(n20464) );
  NOR U20982 ( .A(n21740), .B(n21741), .Z(n21738) );
  XNOR U20983 ( .A(n21742), .B(n21743), .Z(n20723) );
  ANDN U20984 ( .B(n21744), .A(n21745), .Z(n21742) );
  XNOR U20985 ( .A(n19727), .B(n17810), .Z(n14921) );
  XNOR U20986 ( .A(n21746), .B(n20456), .Z(n19727) );
  ANDN U20987 ( .B(n21302), .A(n21301), .Z(n21746) );
  XOR U20988 ( .A(round_reg[707]), .B(n21747), .Z(n21302) );
  XNOR U20989 ( .A(n21748), .B(n12952), .Z(n11402) );
  XNOR U20990 ( .A(n21749), .B(n17445), .Z(n12952) );
  XOR U20991 ( .A(n21750), .B(n19626), .Z(n17445) );
  XNOR U20992 ( .A(n21751), .B(n21752), .Z(n19626) );
  XOR U20993 ( .A(n20198), .B(n20082), .Z(n21752) );
  XOR U20994 ( .A(n21753), .B(n20726), .Z(n20082) );
  XOR U20995 ( .A(round_reg[651]), .B(n21754), .Z(n20726) );
  ANDN U20996 ( .B(n20727), .A(n21755), .Z(n21753) );
  XNOR U20997 ( .A(n21756), .B(n21744), .Z(n20198) );
  ANDN U20998 ( .B(n21745), .A(n21757), .Z(n21756) );
  XOR U20999 ( .A(n15983), .B(n21758), .Z(n21751) );
  XOR U21000 ( .A(n18430), .B(n17991), .Z(n21758) );
  XNOR U21001 ( .A(n21759), .B(n20730), .Z(n17991) );
  XOR U21002 ( .A(round_reg[729]), .B(n21760), .Z(n20730) );
  XNOR U21003 ( .A(n21762), .B(n20716), .Z(n18430) );
  XOR U21004 ( .A(round_reg[943]), .B(n21763), .Z(n20716) );
  ANDN U21005 ( .B(n20717), .A(n21764), .Z(n21762) );
  XNOR U21006 ( .A(n21765), .B(n20720), .Z(n15983) );
  XOR U21007 ( .A(round_reg[775]), .B(n21766), .Z(n20720) );
  ANDN U21008 ( .B(n20721), .A(n21767), .Z(n21765) );
  ANDN U21009 ( .B(n14913), .A(n13131), .Z(n21748) );
  XNOR U21010 ( .A(n20634), .B(n18399), .Z(n13131) );
  XNOR U21011 ( .A(n21768), .B(n21769), .Z(n20579) );
  XOR U21012 ( .A(n18962), .B(n19613), .Z(n21769) );
  XOR U21013 ( .A(n21770), .B(n21771), .Z(n19613) );
  ANDN U21014 ( .B(n20639), .A(n19102), .Z(n21770) );
  XOR U21015 ( .A(round_reg[60]), .B(n21772), .Z(n19102) );
  XNOR U21016 ( .A(n21773), .B(n21774), .Z(n18962) );
  ANDN U21017 ( .B(n20641), .A(n19092), .Z(n21773) );
  XOR U21018 ( .A(round_reg[312]), .B(n21775), .Z(n19092) );
  XOR U21019 ( .A(n21776), .B(n21777), .Z(n21768) );
  XOR U21020 ( .A(n17178), .B(n17127), .Z(n21777) );
  XNOR U21021 ( .A(n21778), .B(n21779), .Z(n17127) );
  ANDN U21022 ( .B(n21780), .A(n19088), .Z(n21778) );
  XNOR U21023 ( .A(n21781), .B(n21782), .Z(n17178) );
  ANDN U21024 ( .B(n20636), .A(n19098), .Z(n21781) );
  XOR U21025 ( .A(round_reg[200]), .B(n21783), .Z(n19098) );
  XOR U21026 ( .A(n21785), .B(n21780), .Z(n20634) );
  ANDN U21027 ( .B(n19088), .A(n19089), .Z(n21785) );
  XOR U21028 ( .A(round_reg[82]), .B(n21786), .Z(n19088) );
  XNOR U21029 ( .A(n21787), .B(n18323), .Z(n14913) );
  XNOR U21030 ( .A(n21788), .B(n15636), .Z(n14895) );
  XNOR U21031 ( .A(n21789), .B(n16458), .Z(n15636) );
  XNOR U21032 ( .A(n21790), .B(n21791), .Z(n16458) );
  XOR U21033 ( .A(n21792), .B(n15591), .Z(n14797) );
  XNOR U21034 ( .A(n21793), .B(n17203), .Z(n14798) );
  IV U21035 ( .A(n18510), .Z(n17203) );
  XOR U21036 ( .A(n21796), .B(n6622), .Z(n3483) );
  IV U21037 ( .A(n9271), .Z(n6622) );
  XNOR U21038 ( .A(n13844), .B(n10050), .Z(n9271) );
  XNOR U21039 ( .A(n12935), .B(n16825), .Z(n10050) );
  XNOR U21040 ( .A(n21797), .B(n21798), .Z(n16825) );
  XOR U21041 ( .A(n10163), .B(n10881), .Z(n21798) );
  XNOR U21042 ( .A(n21799), .B(n17768), .Z(n10881) );
  XNOR U21043 ( .A(n18114), .B(n20966), .Z(n17768) );
  XNOR U21044 ( .A(n21800), .B(n21561), .Z(n20966) );
  ANDN U21045 ( .B(n21801), .A(n21802), .Z(n21800) );
  IV U21046 ( .A(n17275), .Z(n18114) );
  ANDN U21047 ( .B(n15050), .A(n15051), .Z(n21799) );
  XOR U21048 ( .A(n21803), .B(n15591), .Z(n15051) );
  XNOR U21049 ( .A(n21804), .B(n21805), .Z(n18912) );
  XOR U21050 ( .A(n19380), .B(n18806), .Z(n21805) );
  XOR U21051 ( .A(n21806), .B(n21807), .Z(n18806) );
  ANDN U21052 ( .B(n21808), .A(n21809), .Z(n21806) );
  XNOR U21053 ( .A(n21810), .B(n21811), .Z(n19380) );
  ANDN U21054 ( .B(n21812), .A(n21813), .Z(n21810) );
  XOR U21055 ( .A(n17185), .B(n21814), .Z(n21804) );
  XOR U21056 ( .A(n19436), .B(n21815), .Z(n21814) );
  XNOR U21057 ( .A(n21816), .B(n21817), .Z(n19436) );
  XNOR U21058 ( .A(n21820), .B(n21821), .Z(n17185) );
  ANDN U21059 ( .B(n21822), .A(n21823), .Z(n21820) );
  XOR U21060 ( .A(n21825), .B(n18663), .Z(n15050) );
  IV U21061 ( .A(n17506), .Z(n18663) );
  XNOR U21062 ( .A(n17752), .B(n21826), .Z(n10163) );
  XOR U21063 ( .A(n21827), .B(n21828), .Z(n21826) );
  NAND U21064 ( .A(n15691), .B(n4510), .Z(n21828) );
  ANDN U21065 ( .B(n13841), .A(n13842), .Z(n21827) );
  XNOR U21066 ( .A(n21698), .B(n17042), .Z(n13842) );
  XNOR U21067 ( .A(n21829), .B(n20307), .Z(n21698) );
  AND U21068 ( .A(n20924), .B(n20923), .Z(n21829) );
  XNOR U21069 ( .A(n21830), .B(n17945), .Z(n13841) );
  XOR U21070 ( .A(n19074), .B(n20909), .Z(n17945) );
  XOR U21071 ( .A(n21831), .B(n21832), .Z(n20909) );
  XNOR U21072 ( .A(n20424), .B(n16701), .Z(n21832) );
  XOR U21073 ( .A(n21833), .B(n21834), .Z(n16701) );
  ANDN U21074 ( .B(n20431), .A(n21835), .Z(n21833) );
  XOR U21075 ( .A(n21836), .B(n20442), .Z(n20424) );
  ANDN U21076 ( .B(n20441), .A(n21837), .Z(n21836) );
  XOR U21077 ( .A(n17916), .B(n21838), .Z(n21831) );
  XOR U21078 ( .A(n18750), .B(n18211), .Z(n21838) );
  XNOR U21079 ( .A(n21839), .B(n21840), .Z(n18211) );
  ANDN U21080 ( .B(n21841), .A(n21842), .Z(n21839) );
  XOR U21081 ( .A(n21843), .B(n21844), .Z(n18750) );
  ANDN U21082 ( .B(n20435), .A(n21845), .Z(n21843) );
  XOR U21083 ( .A(n21846), .B(n21847), .Z(n17916) );
  NOR U21084 ( .A(n21848), .B(n21849), .Z(n21846) );
  XOR U21085 ( .A(n21850), .B(n21851), .Z(n19074) );
  XNOR U21086 ( .A(n15627), .B(n17227), .Z(n21851) );
  XOR U21087 ( .A(n21852), .B(n21853), .Z(n17227) );
  ANDN U21088 ( .B(n21854), .A(n21855), .Z(n21852) );
  XNOR U21089 ( .A(n21856), .B(n21857), .Z(n15627) );
  AND U21090 ( .A(n21858), .B(n21859), .Z(n21856) );
  XOR U21091 ( .A(n21860), .B(n21861), .Z(n21850) );
  XOR U21092 ( .A(n19252), .B(n18516), .Z(n21861) );
  XNOR U21093 ( .A(n21862), .B(n21863), .Z(n18516) );
  NOR U21094 ( .A(n21864), .B(n21865), .Z(n21862) );
  XOR U21095 ( .A(n21866), .B(n21867), .Z(n19252) );
  ANDN U21096 ( .B(n21868), .A(n21869), .Z(n21866) );
  XOR U21097 ( .A(n20355), .B(n17555), .Z(n17752) );
  XOR U21098 ( .A(n21870), .B(n21871), .Z(n20355) );
  XOR U21099 ( .A(n21872), .B(n21873), .Z(n21871) );
  NAND U21100 ( .A(n6836), .B(n11365), .Z(n21873) );
  ANDN U21101 ( .B(n20598), .A(n21874), .Z(n21872) );
  IV U21102 ( .A(n21875), .Z(n20598) );
  XNOR U21103 ( .A(n17818), .B(n21876), .Z(n21797) );
  XOR U21104 ( .A(n12637), .B(n10378), .Z(n21876) );
  XOR U21105 ( .A(n21877), .B(n17822), .Z(n10378) );
  IV U21106 ( .A(n17765), .Z(n17822) );
  XOR U21107 ( .A(n18034), .B(n21878), .Z(n17765) );
  IV U21108 ( .A(n19049), .Z(n18034) );
  XNOR U21109 ( .A(n19352), .B(n20852), .Z(n19049) );
  XNOR U21110 ( .A(n21879), .B(n21880), .Z(n20852) );
  XOR U21111 ( .A(n17245), .B(n20274), .Z(n21880) );
  XNOR U21112 ( .A(n21881), .B(n20962), .Z(n20274) );
  ANDN U21113 ( .B(n21882), .A(n21883), .Z(n21881) );
  XNOR U21114 ( .A(n21884), .B(n20955), .Z(n17245) );
  ANDN U21115 ( .B(n21885), .A(n21886), .Z(n21884) );
  XNOR U21116 ( .A(n16538), .B(n21887), .Z(n21879) );
  XOR U21117 ( .A(n21888), .B(n16531), .Z(n21887) );
  XNOR U21118 ( .A(n21889), .B(n21890), .Z(n16531) );
  ANDN U21119 ( .B(n21891), .A(n21892), .Z(n21889) );
  XNOR U21120 ( .A(n21893), .B(n20951), .Z(n16538) );
  ANDN U21121 ( .B(n21894), .A(n21895), .Z(n21893) );
  XNOR U21122 ( .A(n21896), .B(n21897), .Z(n19352) );
  XOR U21123 ( .A(n17399), .B(n21257), .Z(n21897) );
  XNOR U21124 ( .A(n21898), .B(n20979), .Z(n21257) );
  AND U21125 ( .A(n21556), .B(n21899), .Z(n21898) );
  XNOR U21126 ( .A(n21900), .B(n21802), .Z(n17399) );
  AND U21127 ( .A(n21560), .B(n21559), .Z(n21900) );
  XOR U21128 ( .A(n16791), .B(n21901), .Z(n21896) );
  XOR U21129 ( .A(n17453), .B(n21902), .Z(n21901) );
  XNOR U21130 ( .A(n21903), .B(n21904), .Z(n17453) );
  ANDN U21131 ( .B(n21547), .A(n21545), .Z(n21903) );
  XNOR U21132 ( .A(n21905), .B(n20976), .Z(n16791) );
  ANDN U21133 ( .B(n21550), .A(n21549), .Z(n21905) );
  ANDN U21134 ( .B(n14194), .A(n14192), .Z(n21877) );
  XOR U21135 ( .A(n21906), .B(n19696), .Z(n14192) );
  IV U21136 ( .A(n18135), .Z(n19696) );
  XNOR U21137 ( .A(n21907), .B(n18978), .Z(n18135) );
  XNOR U21138 ( .A(n21908), .B(n21909), .Z(n18978) );
  XNOR U21139 ( .A(n18253), .B(n18987), .Z(n21909) );
  XOR U21140 ( .A(n21910), .B(n20540), .Z(n18987) );
  XOR U21141 ( .A(round_reg[13]), .B(n21911), .Z(n20540) );
  ANDN U21142 ( .B(n21292), .A(n21912), .Z(n21910) );
  XOR U21143 ( .A(n21913), .B(n20535), .Z(n18253) );
  XOR U21144 ( .A(round_reg[217]), .B(n21914), .Z(n20535) );
  ANDN U21145 ( .B(n21288), .A(n21915), .Z(n21913) );
  XOR U21146 ( .A(n20083), .B(n21916), .Z(n21908) );
  XOR U21147 ( .A(n19384), .B(n19028), .Z(n21916) );
  XOR U21148 ( .A(n21917), .B(n21051), .Z(n19028) );
  IV U21149 ( .A(n21295), .Z(n21051) );
  XOR U21150 ( .A(round_reg[265]), .B(n21185), .Z(n21295) );
  NOR U21151 ( .A(n21294), .B(n21918), .Z(n21917) );
  XOR U21152 ( .A(n21919), .B(n20544), .Z(n19384) );
  IV U21153 ( .A(n21285), .Z(n20544) );
  XOR U21154 ( .A(round_reg[99]), .B(n21920), .Z(n21285) );
  AND U21155 ( .A(n21286), .B(n21921), .Z(n21919) );
  XOR U21156 ( .A(n21922), .B(n20787), .Z(n20083) );
  NOR U21157 ( .A(n21297), .B(n21924), .Z(n21922) );
  XOR U21158 ( .A(n20791), .B(n21626), .Z(n14194) );
  XNOR U21159 ( .A(n21925), .B(n21926), .Z(n21626) );
  ANDN U21160 ( .B(n20474), .A(n20475), .Z(n21925) );
  IV U21161 ( .A(n18990), .Z(n20791) );
  XNOR U21162 ( .A(n21927), .B(n21928), .Z(n18990) );
  XOR U21163 ( .A(n21929), .B(n17761), .Z(n12637) );
  XOR U21164 ( .A(n19217), .B(n21930), .Z(n17761) );
  NOR U21165 ( .A(n18447), .B(n17829), .Z(n21929) );
  XNOR U21166 ( .A(n21931), .B(n16830), .Z(n17829) );
  IV U21167 ( .A(n19400), .Z(n16830) );
  XOR U21168 ( .A(n21932), .B(n21322), .Z(n19400) );
  XOR U21169 ( .A(n21933), .B(n21934), .Z(n21322) );
  XOR U21170 ( .A(n16522), .B(n18488), .Z(n21934) );
  XOR U21171 ( .A(n21935), .B(n19514), .Z(n18488) );
  NOR U21172 ( .A(n21936), .B(n21937), .Z(n21935) );
  XNOR U21173 ( .A(n21938), .B(n19527), .Z(n16522) );
  ANDN U21174 ( .B(n21939), .A(n19973), .Z(n21938) );
  XOR U21175 ( .A(n20938), .B(n21940), .Z(n21933) );
  XOR U21176 ( .A(n17949), .B(n17737), .Z(n21940) );
  XNOR U21177 ( .A(n21941), .B(n19523), .Z(n17737) );
  ANDN U21178 ( .B(n21942), .A(n20014), .Z(n21941) );
  XNOR U21179 ( .A(n21943), .B(n19519), .Z(n17949) );
  ANDN U21180 ( .B(n21944), .A(n19650), .Z(n21943) );
  XNOR U21181 ( .A(n21945), .B(n19510), .Z(n20938) );
  ANDN U21182 ( .B(n21946), .A(n19645), .Z(n21945) );
  XOR U21183 ( .A(n15647), .B(n21947), .Z(n18447) );
  XNOR U21184 ( .A(n21948), .B(n21949), .Z(n20828) );
  XOR U21185 ( .A(n17196), .B(n17334), .Z(n21949) );
  XOR U21186 ( .A(n21950), .B(n21951), .Z(n17334) );
  AND U21187 ( .A(n21952), .B(n21953), .Z(n21950) );
  XNOR U21188 ( .A(n21954), .B(n21955), .Z(n17196) );
  ANDN U21189 ( .B(n21956), .A(n21957), .Z(n21954) );
  XOR U21190 ( .A(n18096), .B(n21958), .Z(n21948) );
  XOR U21191 ( .A(n18290), .B(n18597), .Z(n21958) );
  XNOR U21192 ( .A(n21959), .B(n21960), .Z(n18597) );
  ANDN U21193 ( .B(n21961), .A(n21962), .Z(n21959) );
  XNOR U21194 ( .A(n21963), .B(n21964), .Z(n18290) );
  AND U21195 ( .A(n21965), .B(n21966), .Z(n21963) );
  XNOR U21196 ( .A(n21967), .B(n21968), .Z(n18096) );
  ANDN U21197 ( .B(n21969), .A(n21970), .Z(n21967) );
  XNOR U21198 ( .A(n21971), .B(n21972), .Z(n21636) );
  XNOR U21199 ( .A(n13887), .B(n19311), .Z(n21972) );
  XNOR U21200 ( .A(n21973), .B(n21974), .Z(n19311) );
  ANDN U21201 ( .B(n21975), .A(n21976), .Z(n21973) );
  XNOR U21202 ( .A(n21977), .B(n21978), .Z(n13887) );
  ANDN U21203 ( .B(n21979), .A(n21980), .Z(n21977) );
  XOR U21204 ( .A(n19199), .B(n21981), .Z(n21971) );
  XOR U21205 ( .A(n19235), .B(n21982), .Z(n21981) );
  XNOR U21206 ( .A(n21983), .B(n21984), .Z(n19235) );
  AND U21207 ( .A(n21985), .B(n21986), .Z(n21983) );
  XNOR U21208 ( .A(n21987), .B(n21988), .Z(n19199) );
  ANDN U21209 ( .B(n21989), .A(n21990), .Z(n21987) );
  XNOR U21210 ( .A(n21991), .B(n17756), .Z(n17818) );
  XNOR U21211 ( .A(n21992), .B(n15525), .Z(n17756) );
  XOR U21212 ( .A(n19636), .B(n18913), .Z(n15525) );
  XOR U21213 ( .A(n21993), .B(n21994), .Z(n18913) );
  XNOR U21214 ( .A(n17563), .B(n19588), .Z(n21994) );
  XOR U21215 ( .A(n21995), .B(n21275), .Z(n19588) );
  ANDN U21216 ( .B(n21996), .A(n21997), .Z(n21995) );
  XNOR U21217 ( .A(n21998), .B(n21277), .Z(n17563) );
  ANDN U21218 ( .B(n21999), .A(n20814), .Z(n21998) );
  XOR U21219 ( .A(n18571), .B(n22000), .Z(n21993) );
  XOR U21220 ( .A(n22001), .B(n19908), .Z(n22000) );
  XNOR U21221 ( .A(n22002), .B(n21271), .Z(n19908) );
  NOR U21222 ( .A(n22003), .B(n20820), .Z(n22002) );
  XNOR U21223 ( .A(n22004), .B(n21264), .Z(n18571) );
  ANDN U21224 ( .B(n22005), .A(n20824), .Z(n22004) );
  XOR U21225 ( .A(n22006), .B(n22007), .Z(n19636) );
  XNOR U21226 ( .A(n16269), .B(n17007), .Z(n22007) );
  XNOR U21227 ( .A(n22008), .B(n22009), .Z(n17007) );
  ANDN U21228 ( .B(n22010), .A(n20350), .Z(n22008) );
  XOR U21229 ( .A(n22011), .B(n22012), .Z(n16269) );
  ANDN U21230 ( .B(n20346), .A(n22013), .Z(n22011) );
  XOR U21231 ( .A(n16740), .B(n22014), .Z(n22006) );
  XOR U21232 ( .A(n22015), .B(n17079), .Z(n22014) );
  XOR U21233 ( .A(n22016), .B(n22017), .Z(n17079) );
  ANDN U21234 ( .B(n22018), .A(n20342), .Z(n22016) );
  XNOR U21235 ( .A(n22019), .B(n22020), .Z(n16740) );
  ANDN U21236 ( .B(n22021), .A(n20337), .Z(n22019) );
  AND U21237 ( .A(n18460), .B(n17824), .Z(n21991) );
  XOR U21238 ( .A(n22022), .B(n22023), .Z(n12935) );
  XNOR U21239 ( .A(n10095), .B(n11734), .Z(n22023) );
  XOR U21240 ( .A(n22024), .B(n16224), .Z(n11734) );
  XOR U21241 ( .A(n22025), .B(n18643), .Z(n16224) );
  XOR U21242 ( .A(n19671), .B(n21795), .Z(n18643) );
  XOR U21243 ( .A(n22026), .B(n22027), .Z(n21795) );
  XNOR U21244 ( .A(n18897), .B(n22028), .Z(n22027) );
  XOR U21245 ( .A(n22029), .B(n19759), .Z(n18897) );
  IV U21246 ( .A(n22030), .Z(n19759) );
  ANDN U21247 ( .B(n22031), .A(n22032), .Z(n22029) );
  XOR U21248 ( .A(n17122), .B(n22033), .Z(n22026) );
  XOR U21249 ( .A(n18282), .B(n18577), .Z(n22033) );
  XOR U21250 ( .A(n22034), .B(n19750), .Z(n18577) );
  ANDN U21251 ( .B(n20838), .A(n22035), .Z(n22034) );
  XOR U21252 ( .A(n22036), .B(n19754), .Z(n18282) );
  ANDN U21253 ( .B(n20832), .A(n22037), .Z(n22036) );
  XOR U21254 ( .A(n22038), .B(n19763), .Z(n17122) );
  ANDN U21255 ( .B(n20834), .A(n22039), .Z(n22038) );
  XOR U21256 ( .A(n22040), .B(n22041), .Z(n19671) );
  XNOR U21257 ( .A(n20094), .B(n19160), .Z(n22041) );
  XNOR U21258 ( .A(n22042), .B(n22043), .Z(n19160) );
  NOR U21259 ( .A(n21960), .B(n22044), .Z(n22042) );
  XNOR U21260 ( .A(n22045), .B(n22046), .Z(n20094) );
  NOR U21261 ( .A(n21968), .B(n22047), .Z(n22045) );
  XOR U21262 ( .A(n19968), .B(n22048), .Z(n22040) );
  XOR U21263 ( .A(n19246), .B(n16036), .Z(n22048) );
  XNOR U21264 ( .A(n22049), .B(n22050), .Z(n16036) );
  NOR U21265 ( .A(n21951), .B(n22051), .Z(n22049) );
  XNOR U21266 ( .A(n22052), .B(n22053), .Z(n19246) );
  NOR U21267 ( .A(n21964), .B(n22054), .Z(n22052) );
  XNOR U21268 ( .A(n22055), .B(n22056), .Z(n19968) );
  ANDN U21269 ( .B(n22057), .A(n21955), .Z(n22055) );
  AND U21270 ( .A(n16182), .B(n16181), .Z(n22024) );
  XNOR U21271 ( .A(n21687), .B(n17589), .Z(n16181) );
  IV U21272 ( .A(n18160), .Z(n17589) );
  XNOR U21273 ( .A(n18632), .B(n22058), .Z(n18160) );
  XNOR U21274 ( .A(n22059), .B(n22060), .Z(n18632) );
  XNOR U21275 ( .A(n16915), .B(n15975), .Z(n22060) );
  XOR U21276 ( .A(n22061), .B(n22062), .Z(n15975) );
  ANDN U21277 ( .B(n21684), .A(n21683), .Z(n22061) );
  XNOR U21278 ( .A(n22063), .B(n22064), .Z(n16915) );
  ANDN U21279 ( .B(n21681), .A(n21679), .Z(n22063) );
  XNOR U21280 ( .A(n17398), .B(n22065), .Z(n22059) );
  XOR U21281 ( .A(n19716), .B(n18212), .Z(n22065) );
  XOR U21282 ( .A(n22066), .B(n22067), .Z(n18212) );
  AND U21283 ( .A(n21693), .B(n21695), .Z(n22066) );
  XNOR U21284 ( .A(n22068), .B(n22069), .Z(n19716) );
  NOR U21285 ( .A(n22070), .B(n22071), .Z(n22068) );
  XNOR U21286 ( .A(n22072), .B(n22073), .Z(n17398) );
  ANDN U21287 ( .B(n21689), .A(n21690), .Z(n22072) );
  XOR U21288 ( .A(n22074), .B(n22071), .Z(n21687) );
  AND U21289 ( .A(n22070), .B(n22075), .Z(n22074) );
  XNOR U21290 ( .A(n22076), .B(n21123), .Z(n16182) );
  XOR U21291 ( .A(n19913), .B(n22077), .Z(n21123) );
  XOR U21292 ( .A(n22078), .B(n22079), .Z(n19913) );
  XOR U21293 ( .A(n16787), .B(n17293), .Z(n22079) );
  XOR U21294 ( .A(n22080), .B(n22081), .Z(n17293) );
  AND U21295 ( .A(n22082), .B(n22083), .Z(n22080) );
  XNOR U21296 ( .A(n22084), .B(n22085), .Z(n16787) );
  ANDN U21297 ( .B(n22086), .A(n22087), .Z(n22084) );
  XOR U21298 ( .A(n18615), .B(n22088), .Z(n22078) );
  XNOR U21299 ( .A(n19459), .B(n22089), .Z(n22088) );
  XNOR U21300 ( .A(n22090), .B(n22091), .Z(n19459) );
  ANDN U21301 ( .B(n22092), .A(n22093), .Z(n22090) );
  XOR U21302 ( .A(n22094), .B(n22095), .Z(n18615) );
  NOR U21303 ( .A(n22096), .B(n22097), .Z(n22094) );
  XNOR U21304 ( .A(n22098), .B(n16227), .Z(n10095) );
  XNOR U21305 ( .A(n22099), .B(n19703), .Z(n16227) );
  ANDN U21306 ( .B(n16178), .A(n16176), .Z(n22098) );
  XOR U21307 ( .A(n22100), .B(n17683), .Z(n16176) );
  IV U21308 ( .A(n17534), .Z(n17683) );
  XNOR U21309 ( .A(n21125), .B(n21928), .Z(n17534) );
  XNOR U21310 ( .A(n22101), .B(n22102), .Z(n21928) );
  XNOR U21311 ( .A(n17449), .B(n18195), .Z(n22102) );
  XNOR U21312 ( .A(n22103), .B(n22104), .Z(n18195) );
  AND U21313 ( .A(n20487), .B(n21623), .Z(n22103) );
  XNOR U21314 ( .A(round_reg[946]), .B(n22105), .Z(n20487) );
  XNOR U21315 ( .A(n22106), .B(n22107), .Z(n17449) );
  NOR U21316 ( .A(n21625), .B(n20479), .Z(n22106) );
  XOR U21317 ( .A(round_reg[778]), .B(n22108), .Z(n20479) );
  XOR U21318 ( .A(n18419), .B(n22109), .Z(n22101) );
  XOR U21319 ( .A(n17166), .B(n19679), .Z(n22109) );
  XNOR U21320 ( .A(n22110), .B(n22111), .Z(n19679) );
  XOR U21321 ( .A(round_reg[875]), .B(n22112), .Z(n20483) );
  XNOR U21322 ( .A(n22113), .B(n22114), .Z(n17166) );
  NOR U21323 ( .A(n21629), .B(n20470), .Z(n22113) );
  XOR U21324 ( .A(round_reg[654]), .B(n22115), .Z(n20470) );
  XNOR U21325 ( .A(n22116), .B(n22117), .Z(n18419) );
  ANDN U21326 ( .B(n22118), .A(n20474), .Z(n22116) );
  XOR U21327 ( .A(round_reg[732]), .B(n22119), .Z(n20474) );
  XOR U21328 ( .A(n22120), .B(n22121), .Z(n21125) );
  XNOR U21329 ( .A(n17797), .B(n17782), .Z(n22121) );
  XNOR U21330 ( .A(n22122), .B(n22123), .Z(n17782) );
  XNOR U21331 ( .A(n22126), .B(n22127), .Z(n17797) );
  ANDN U21332 ( .B(n22128), .A(n22129), .Z(n22126) );
  XOR U21333 ( .A(n17734), .B(n22130), .Z(n22120) );
  XOR U21334 ( .A(n17044), .B(n22131), .Z(n22130) );
  XNOR U21335 ( .A(n22132), .B(n22133), .Z(n17044) );
  XNOR U21336 ( .A(n22136), .B(n22137), .Z(n17734) );
  NOR U21337 ( .A(n22138), .B(n22139), .Z(n22136) );
  XNOR U21338 ( .A(n19263), .B(n20692), .Z(n16178) );
  XNOR U21339 ( .A(n22140), .B(n21227), .Z(n20692) );
  ANDN U21340 ( .B(n20188), .A(n20186), .Z(n22140) );
  XNOR U21341 ( .A(n9789), .B(n22141), .Z(n22022) );
  XOR U21342 ( .A(n14877), .B(n10607), .Z(n22141) );
  XOR U21343 ( .A(n22142), .B(n17008), .Z(n10607) );
  XOR U21344 ( .A(n22143), .B(n22144), .Z(n17008) );
  XNOR U21345 ( .A(n22145), .B(n16603), .Z(n16172) );
  XOR U21346 ( .A(n19990), .B(n22146), .Z(n16603) );
  XNOR U21347 ( .A(n22147), .B(n22148), .Z(n19990) );
  XOR U21348 ( .A(n18687), .B(n18400), .Z(n22148) );
  XOR U21349 ( .A(n22149), .B(n20056), .Z(n18400) );
  NOR U21350 ( .A(n20055), .B(n22150), .Z(n22149) );
  XNOR U21351 ( .A(n22151), .B(n20047), .Z(n18687) );
  NOR U21352 ( .A(n22152), .B(n20046), .Z(n22151) );
  XNOR U21353 ( .A(n20040), .B(n22153), .Z(n22147) );
  XOR U21354 ( .A(n17269), .B(n17596), .Z(n22153) );
  XNOR U21355 ( .A(n22154), .B(n20064), .Z(n17596) );
  AND U21356 ( .A(n20063), .B(n22155), .Z(n22154) );
  XNOR U21357 ( .A(n22156), .B(n22157), .Z(n17269) );
  ANDN U21358 ( .B(n22158), .A(n20050), .Z(n22156) );
  XNOR U21359 ( .A(n22159), .B(n20060), .Z(n20040) );
  NOR U21360 ( .A(n22160), .B(n20059), .Z(n22159) );
  XNOR U21361 ( .A(n21066), .B(n18002), .Z(n16173) );
  XOR U21362 ( .A(n22161), .B(n22162), .Z(n21066) );
  ANDN U21363 ( .B(n22163), .A(n22164), .Z(n22161) );
  XNOR U21364 ( .A(n22165), .B(n16221), .Z(n14877) );
  XNOR U21365 ( .A(n22166), .B(n15631), .Z(n16221) );
  IV U21366 ( .A(n17455), .Z(n15631) );
  XNOR U21367 ( .A(n22167), .B(n22168), .Z(n17455) );
  AND U21368 ( .A(n16185), .B(n16187), .Z(n22165) );
  XNOR U21369 ( .A(n20876), .B(n20799), .Z(n16187) );
  XNOR U21370 ( .A(n22169), .B(n22170), .Z(n20799) );
  AND U21371 ( .A(n21151), .B(n22171), .Z(n22169) );
  XNOR U21372 ( .A(n22172), .B(n18976), .Z(n16185) );
  XOR U21373 ( .A(n20614), .B(n19166), .Z(n18976) );
  XOR U21374 ( .A(n22173), .B(n22174), .Z(n19166) );
  XNOR U21375 ( .A(n18335), .B(n20028), .Z(n22174) );
  XOR U21376 ( .A(n22175), .B(n22176), .Z(n20028) );
  NOR U21377 ( .A(n22177), .B(n22178), .Z(n22175) );
  XOR U21378 ( .A(n22179), .B(n22180), .Z(n18335) );
  XOR U21379 ( .A(n19656), .B(n22183), .Z(n22173) );
  XOR U21380 ( .A(n19551), .B(n16518), .Z(n22183) );
  XOR U21381 ( .A(n22184), .B(n22185), .Z(n16518) );
  NOR U21382 ( .A(n22186), .B(n22187), .Z(n22184) );
  XOR U21383 ( .A(n22188), .B(n22189), .Z(n19551) );
  XOR U21384 ( .A(n22192), .B(n22193), .Z(n19656) );
  XOR U21385 ( .A(n22196), .B(n22197), .Z(n20614) );
  XNOR U21386 ( .A(n21181), .B(n19110), .Z(n22197) );
  XOR U21387 ( .A(n22198), .B(n20216), .Z(n19110) );
  ANDN U21388 ( .B(n21212), .A(n22199), .Z(n22198) );
  XNOR U21389 ( .A(n22200), .B(n20225), .Z(n21181) );
  XNOR U21390 ( .A(round_reg[358]), .B(n22201), .Z(n20225) );
  ANDN U21391 ( .B(n21205), .A(n22202), .Z(n22200) );
  IV U21392 ( .A(n22203), .Z(n21205) );
  XNOR U21393 ( .A(n18375), .B(n22204), .Z(n22196) );
  XOR U21394 ( .A(n18830), .B(n18405), .Z(n22204) );
  XNOR U21395 ( .A(n22205), .B(n20222), .Z(n18405) );
  XOR U21396 ( .A(round_reg[581]), .B(n22206), .Z(n20222) );
  ANDN U21397 ( .B(n21203), .A(n22207), .Z(n22205) );
  XNOR U21398 ( .A(n22208), .B(n21209), .Z(n18830) );
  AND U21399 ( .A(n21210), .B(n22209), .Z(n22208) );
  XOR U21400 ( .A(n22210), .B(n20212), .Z(n18375) );
  XNOR U21401 ( .A(round_reg[513]), .B(n22211), .Z(n20212) );
  ANDN U21402 ( .B(n21214), .A(n22212), .Z(n22210) );
  XNOR U21403 ( .A(n22213), .B(n16217), .Z(n9789) );
  XOR U21404 ( .A(n16024), .B(n22214), .Z(n16217) );
  XNOR U21405 ( .A(n20495), .B(n22215), .Z(n16024) );
  XOR U21406 ( .A(n22216), .B(n22217), .Z(n20495) );
  XOR U21407 ( .A(n19822), .B(n18359), .Z(n22217) );
  XOR U21408 ( .A(n22218), .B(n19844), .Z(n18359) );
  XOR U21409 ( .A(round_reg[998]), .B(n22201), .Z(n19844) );
  AND U21410 ( .A(n22219), .B(n19845), .Z(n22218) );
  XNOR U21411 ( .A(n22220), .B(n19848), .Z(n19822) );
  XOR U21412 ( .A(round_reg[1166]), .B(n22221), .Z(n19848) );
  AND U21413 ( .A(n22222), .B(n19849), .Z(n22220) );
  XOR U21414 ( .A(n18815), .B(n22223), .Z(n22216) );
  XOR U21415 ( .A(n17249), .B(n16260), .Z(n22223) );
  XNOR U21416 ( .A(n22224), .B(n19853), .Z(n16260) );
  XOR U21417 ( .A(round_reg[1238]), .B(n22225), .Z(n19853) );
  XNOR U21418 ( .A(n22227), .B(n19857), .Z(n17249) );
  XNOR U21419 ( .A(round_reg[1027]), .B(n21747), .Z(n19857) );
  ANDN U21420 ( .B(n19858), .A(n22228), .Z(n22227) );
  XNOR U21421 ( .A(n22229), .B(n19861), .Z(n18815) );
  XOR U21422 ( .A(round_reg[1140]), .B(n22230), .Z(n19861) );
  AND U21423 ( .A(n22231), .B(n22232), .Z(n22229) );
  AND U21424 ( .A(n16190), .B(n17836), .Z(n22213) );
  XNOR U21425 ( .A(n20678), .B(n17031), .Z(n17836) );
  XOR U21426 ( .A(n22233), .B(n22234), .Z(n20678) );
  ANDN U21427 ( .B(n22235), .A(n22236), .Z(n22233) );
  XNOR U21428 ( .A(n19217), .B(n22237), .Z(n16190) );
  XNOR U21429 ( .A(n18683), .B(n22238), .Z(n19217) );
  XOR U21430 ( .A(n22239), .B(n22240), .Z(n18683) );
  XOR U21431 ( .A(n17116), .B(n17950), .Z(n22240) );
  XOR U21432 ( .A(n22241), .B(n22242), .Z(n17950) );
  ANDN U21433 ( .B(n22243), .A(n22244), .Z(n22241) );
  XNOR U21434 ( .A(n22245), .B(n22246), .Z(n17116) );
  ANDN U21435 ( .B(n22247), .A(n22248), .Z(n22245) );
  XOR U21436 ( .A(n20737), .B(n22249), .Z(n22239) );
  XOR U21437 ( .A(n16817), .B(n22250), .Z(n22249) );
  XNOR U21438 ( .A(n22251), .B(n22252), .Z(n16817) );
  ANDN U21439 ( .B(n22253), .A(n22254), .Z(n22251) );
  XOR U21440 ( .A(n22255), .B(n22256), .Z(n20737) );
  NOR U21441 ( .A(n22257), .B(n22258), .Z(n22255) );
  XNOR U21442 ( .A(n22259), .B(n17824), .Z(n13844) );
  XNOR U21443 ( .A(n19833), .B(n20734), .Z(n17824) );
  XNOR U21444 ( .A(n22260), .B(n19785), .Z(n20734) );
  XNOR U21445 ( .A(n22261), .B(n22262), .Z(n19785) );
  XOR U21446 ( .A(n18565), .B(n19904), .Z(n22262) );
  XOR U21447 ( .A(n22263), .B(n22264), .Z(n19904) );
  ANDN U21448 ( .B(n19826), .A(n19827), .Z(n22263) );
  XOR U21449 ( .A(round_reg[592]), .B(n22265), .Z(n19827) );
  XOR U21450 ( .A(n22266), .B(n20773), .Z(n18565) );
  ANDN U21451 ( .B(n19830), .A(n19831), .Z(n22266) );
  XOR U21452 ( .A(round_reg[369]), .B(n22267), .Z(n19831) );
  XOR U21453 ( .A(round_reg[736]), .B(n22268), .Z(n19830) );
  XOR U21454 ( .A(n18367), .B(n22269), .Z(n22261) );
  XOR U21455 ( .A(n18397), .B(n19780), .Z(n22269) );
  XOR U21456 ( .A(n22270), .B(n22271), .Z(n19780) );
  ANDN U21457 ( .B(n20736), .A(n20499), .Z(n22270) );
  XOR U21458 ( .A(round_reg[420]), .B(n22272), .Z(n20499) );
  XNOR U21459 ( .A(n22273), .B(n20944), .Z(n18397) );
  ANDN U21460 ( .B(n19837), .A(n19839), .Z(n22273) );
  XOR U21461 ( .A(round_reg[490]), .B(n22274), .Z(n19839) );
  XOR U21462 ( .A(round_reg[879]), .B(n21309), .Z(n19837) );
  XOR U21463 ( .A(n22275), .B(n22276), .Z(n18367) );
  ANDN U21464 ( .B(n20776), .A(n20510), .Z(n22275) );
  XNOR U21465 ( .A(n22277), .B(n20776), .Z(n19833) );
  XOR U21466 ( .A(round_reg[950]), .B(n22278), .Z(n20776) );
  AND U21467 ( .A(n20510), .B(n20512), .Z(n22277) );
  XOR U21468 ( .A(round_reg[524]), .B(n22279), .Z(n20510) );
  NOR U21469 ( .A(n18460), .B(n17755), .Z(n22259) );
  XNOR U21470 ( .A(n22280), .B(n19423), .Z(n17755) );
  XNOR U21471 ( .A(n22281), .B(n22282), .Z(n19632) );
  XNOR U21472 ( .A(n20034), .B(n18486), .Z(n22282) );
  XNOR U21473 ( .A(n22283), .B(n22284), .Z(n18486) );
  ANDN U21474 ( .B(n22285), .A(n22286), .Z(n22283) );
  XNOR U21475 ( .A(n22287), .B(n22288), .Z(n20034) );
  ANDN U21476 ( .B(n22289), .A(n22290), .Z(n22287) );
  XOR U21477 ( .A(n22291), .B(n22292), .Z(n22281) );
  XOR U21478 ( .A(n19223), .B(n16688), .Z(n22292) );
  XNOR U21479 ( .A(n22293), .B(n22294), .Z(n16688) );
  ANDN U21480 ( .B(n22295), .A(n22296), .Z(n22293) );
  XNOR U21481 ( .A(n22297), .B(n22298), .Z(n19223) );
  XNOR U21482 ( .A(n22301), .B(n22302), .Z(n20466) );
  XOR U21483 ( .A(n18999), .B(n18108), .Z(n22302) );
  XOR U21484 ( .A(n22303), .B(n22124), .Z(n18108) );
  ANDN U21485 ( .B(n22304), .A(n22305), .Z(n22303) );
  XNOR U21486 ( .A(n22306), .B(n22134), .Z(n18999) );
  ANDN U21487 ( .B(n22307), .A(n22308), .Z(n22306) );
  XOR U21488 ( .A(n19543), .B(n22309), .Z(n22301) );
  XOR U21489 ( .A(n19595), .B(n21619), .Z(n22309) );
  XNOR U21490 ( .A(n22310), .B(n22311), .Z(n21619) );
  ANDN U21491 ( .B(n22312), .A(n22313), .Z(n22310) );
  XNOR U21492 ( .A(n22314), .B(n22129), .Z(n19595) );
  ANDN U21493 ( .B(n22315), .A(n22316), .Z(n22314) );
  XNOR U21494 ( .A(n22317), .B(n22138), .Z(n19543) );
  ANDN U21495 ( .B(n22318), .A(n22319), .Z(n22317) );
  XNOR U21496 ( .A(n18549), .B(n22320), .Z(n18460) );
  IV U21497 ( .A(n17972), .Z(n18549) );
  XOR U21498 ( .A(n20462), .B(n18285), .Z(n17972) );
  XOR U21499 ( .A(n22321), .B(n22322), .Z(n18285) );
  XNOR U21500 ( .A(n22323), .B(n17414), .Z(n22322) );
  XOR U21501 ( .A(n22324), .B(n20158), .Z(n17414) );
  ANDN U21502 ( .B(n20392), .A(n22325), .Z(n22324) );
  XNOR U21503 ( .A(n19346), .B(n22326), .Z(n22321) );
  XOR U21504 ( .A(n18966), .B(n19295), .Z(n22326) );
  XNOR U21505 ( .A(n22327), .B(n20150), .Z(n19295) );
  XOR U21506 ( .A(n22330), .B(n20154), .Z(n18966) );
  NOR U21507 ( .A(n20386), .B(n22331), .Z(n22330) );
  XNOR U21508 ( .A(n22332), .B(n20145), .Z(n19346) );
  XOR U21509 ( .A(n22334), .B(n22335), .Z(n20462) );
  XOR U21510 ( .A(n19313), .B(n20313), .Z(n22335) );
  XOR U21511 ( .A(n22336), .B(n22337), .Z(n20313) );
  ANDN U21512 ( .B(n22338), .A(n20865), .Z(n22336) );
  XNOR U21513 ( .A(n22339), .B(n22340), .Z(n19313) );
  AND U21514 ( .A(n20869), .B(n22341), .Z(n22339) );
  XOR U21515 ( .A(n19542), .B(n22342), .Z(n22334) );
  XOR U21516 ( .A(n19970), .B(n22343), .Z(n22342) );
  XNOR U21517 ( .A(n22344), .B(n22345), .Z(n19970) );
  AND U21518 ( .A(n20856), .B(n22346), .Z(n22344) );
  XNOR U21519 ( .A(n22347), .B(n22348), .Z(n19542) );
  AND U21520 ( .A(n20873), .B(n22349), .Z(n22347) );
  NOR U21521 ( .A(n9196), .B(n7074), .Z(n21796) );
  XNOR U21522 ( .A(n17530), .B(n10008), .Z(n7074) );
  IV U21523 ( .A(n11855), .Z(n10008) );
  XOR U21524 ( .A(n16199), .B(n17046), .Z(n11855) );
  XNOR U21525 ( .A(n22350), .B(n22351), .Z(n17046) );
  XOR U21526 ( .A(n12879), .B(n12936), .Z(n22351) );
  XNOR U21527 ( .A(n22352), .B(n13107), .Z(n12936) );
  XOR U21528 ( .A(n22353), .B(n15606), .Z(n13107) );
  IV U21529 ( .A(n18008), .Z(n15606) );
  XOR U21530 ( .A(n22354), .B(n22355), .Z(n18008) );
  AND U21531 ( .A(n13934), .B(n15206), .Z(n22352) );
  IV U21532 ( .A(n19534), .Z(n15206) );
  XOR U21533 ( .A(n21699), .B(n17042), .Z(n19534) );
  XNOR U21534 ( .A(n22356), .B(n22058), .Z(n17042) );
  XNOR U21535 ( .A(n22357), .B(n22358), .Z(n22058) );
  XNOR U21536 ( .A(n20283), .B(n18890), .Z(n22358) );
  XOR U21537 ( .A(n22359), .B(n20302), .Z(n18890) );
  AND U21538 ( .A(n20303), .B(n20916), .Z(n22359) );
  XOR U21539 ( .A(n22360), .B(n20289), .Z(n20283) );
  AND U21540 ( .A(n20290), .B(n20920), .Z(n22360) );
  XNOR U21541 ( .A(round_reg[551]), .B(n22361), .Z(n20920) );
  XOR U21542 ( .A(round_reg[913]), .B(n22362), .Z(n20290) );
  XNOR U21543 ( .A(n17861), .B(n22363), .Z(n22357) );
  XOR U21544 ( .A(n19686), .B(n20246), .Z(n22363) );
  XNOR U21545 ( .A(n22364), .B(n20299), .Z(n20246) );
  AND U21546 ( .A(n20298), .B(n21704), .Z(n22364) );
  XNOR U21547 ( .A(round_reg[453]), .B(n22365), .Z(n21704) );
  XOR U21548 ( .A(round_reg[842]), .B(n22366), .Z(n20298) );
  XOR U21549 ( .A(n22367), .B(n20306), .Z(n19686) );
  ANDN U21550 ( .B(n20307), .A(n20923), .Z(n22367) );
  XOR U21551 ( .A(round_reg[332]), .B(n22368), .Z(n20923) );
  XOR U21552 ( .A(round_reg[763]), .B(n22369), .Z(n20307) );
  XNOR U21553 ( .A(n22370), .B(n20294), .Z(n17861) );
  AND U21554 ( .A(n20293), .B(n20926), .Z(n22370) );
  IV U21555 ( .A(n21702), .Z(n20926) );
  XOR U21556 ( .A(round_reg[447]), .B(n22371), .Z(n21702) );
  XOR U21557 ( .A(round_reg[809]), .B(n22372), .Z(n20293) );
  XOR U21558 ( .A(n22373), .B(n20303), .Z(n21699) );
  XOR U21559 ( .A(round_reg[685]), .B(n22374), .Z(n20303) );
  XNOR U21560 ( .A(round_reg[619]), .B(n22375), .Z(n20916) );
  XNOR U21561 ( .A(n20958), .B(n18379), .Z(n13934) );
  XNOR U21562 ( .A(n22376), .B(n22377), .Z(n20958) );
  NOR U21563 ( .A(n22378), .B(n22379), .Z(n22376) );
  XOR U21564 ( .A(n22380), .B(n13103), .Z(n12879) );
  XNOR U21565 ( .A(n22323), .B(n19296), .Z(n13103) );
  XOR U21566 ( .A(n22381), .B(n22382), .Z(n19296) );
  XOR U21567 ( .A(n22383), .B(n20162), .Z(n22323) );
  ANDN U21568 ( .B(n20390), .A(n22384), .Z(n22383) );
  AND U21569 ( .A(n13930), .B(n15219), .Z(n22380) );
  IV U21570 ( .A(n17540), .Z(n15219) );
  XOR U21571 ( .A(n21583), .B(n17467), .Z(n17540) );
  XOR U21572 ( .A(n22385), .B(n22386), .Z(n21583) );
  ANDN U21573 ( .B(n22387), .A(n21372), .Z(n22385) );
  XNOR U21574 ( .A(n22388), .B(n17925), .Z(n13930) );
  XNOR U21575 ( .A(n22215), .B(n21259), .Z(n17925) );
  XNOR U21576 ( .A(n22389), .B(n22390), .Z(n21259) );
  XNOR U21577 ( .A(n16759), .B(n22391), .Z(n22390) );
  NOR U21578 ( .A(n22394), .B(n21811), .Z(n22392) );
  XOR U21579 ( .A(n19777), .B(n22395), .Z(n22389) );
  XOR U21580 ( .A(n19032), .B(n22396), .Z(n22395) );
  XOR U21581 ( .A(n22397), .B(n22398), .Z(n19032) );
  ANDN U21582 ( .B(n22399), .A(n22400), .Z(n22397) );
  XOR U21583 ( .A(n22401), .B(n22402), .Z(n19777) );
  ANDN U21584 ( .B(n22403), .A(n21821), .Z(n22401) );
  XOR U21585 ( .A(n22404), .B(n22405), .Z(n22215) );
  XNOR U21586 ( .A(n17082), .B(n18825), .Z(n22405) );
  XNOR U21587 ( .A(n22406), .B(n22093), .Z(n18825) );
  AND U21588 ( .A(n22407), .B(n22408), .Z(n22406) );
  XOR U21589 ( .A(n22409), .B(n22086), .Z(n17082) );
  ANDN U21590 ( .B(n22410), .A(n22411), .Z(n22409) );
  XOR U21591 ( .A(n18887), .B(n22412), .Z(n22404) );
  XNOR U21592 ( .A(n19254), .B(n19497), .Z(n22412) );
  XOR U21593 ( .A(n22413), .B(n22414), .Z(n19497) );
  NOR U21594 ( .A(n22415), .B(n22416), .Z(n22413) );
  XNOR U21595 ( .A(n22417), .B(n22096), .Z(n19254) );
  NOR U21596 ( .A(n22418), .B(n22419), .Z(n22417) );
  XOR U21597 ( .A(n22420), .B(n22421), .Z(n18887) );
  AND U21598 ( .A(n22422), .B(n22423), .Z(n22420) );
  XOR U21599 ( .A(n10707), .B(n22424), .Z(n22350) );
  XNOR U21600 ( .A(n11385), .B(n13686), .Z(n22424) );
  XNOR U21601 ( .A(n22425), .B(n13094), .Z(n13686) );
  XOR U21602 ( .A(n21351), .B(n16612), .Z(n13094) );
  IV U21603 ( .A(n17835), .Z(n16612) );
  XNOR U21604 ( .A(n19175), .B(n22426), .Z(n17835) );
  XNOR U21605 ( .A(n22427), .B(n22428), .Z(n19175) );
  XOR U21606 ( .A(n16922), .B(n16468), .Z(n22428) );
  XOR U21607 ( .A(n22429), .B(n22430), .Z(n16468) );
  AND U21608 ( .A(n20060), .B(n22431), .Z(n22429) );
  XOR U21609 ( .A(round_reg[934]), .B(n22432), .Z(n20060) );
  XNOR U21610 ( .A(n22433), .B(n22434), .Z(n16922) );
  AND U21611 ( .A(n20064), .B(n20062), .Z(n22433) );
  XNOR U21612 ( .A(round_reg[830]), .B(n22435), .Z(n20064) );
  XOR U21613 ( .A(n19260), .B(n22436), .Z(n22427) );
  XOR U21614 ( .A(n19863), .B(n17503), .Z(n22436) );
  XOR U21615 ( .A(n22437), .B(n22438), .Z(n17503) );
  NOR U21616 ( .A(n20051), .B(n20049), .Z(n22437) );
  IV U21617 ( .A(n22157), .Z(n20051) );
  XOR U21618 ( .A(round_reg[863]), .B(n22439), .Z(n22157) );
  XNOR U21619 ( .A(n22440), .B(n22441), .Z(n19863) );
  AND U21620 ( .A(n20056), .B(n20054), .Z(n22440) );
  XNOR U21621 ( .A(round_reg[642]), .B(n22442), .Z(n20056) );
  XNOR U21622 ( .A(n22443), .B(n22444), .Z(n19260) );
  XNOR U21623 ( .A(round_reg[720]), .B(n22445), .Z(n20047) );
  XNOR U21624 ( .A(n22446), .B(n22447), .Z(n21351) );
  AND U21625 ( .A(n22448), .B(n22449), .Z(n22446) );
  AND U21626 ( .A(n13923), .B(n22450), .Z(n22425) );
  XNOR U21627 ( .A(n22451), .B(n13099), .Z(n11385) );
  XNOR U21628 ( .A(n19646), .B(n19597), .Z(n13099) );
  XNOR U21629 ( .A(n22454), .B(n21937), .Z(n19646) );
  AND U21630 ( .A(n15202), .B(n17532), .Z(n22451) );
  XOR U21631 ( .A(n22455), .B(n18940), .Z(n17532) );
  XNOR U21632 ( .A(n22456), .B(n21129), .Z(n18940) );
  XNOR U21633 ( .A(n22457), .B(n22458), .Z(n21129) );
  XNOR U21634 ( .A(n18827), .B(n18476), .Z(n22458) );
  XOR U21635 ( .A(n22459), .B(n22460), .Z(n18476) );
  ANDN U21636 ( .B(n22461), .A(n22462), .Z(n22459) );
  XNOR U21637 ( .A(n22463), .B(n22464), .Z(n18827) );
  AND U21638 ( .A(n22465), .B(n22466), .Z(n22463) );
  XNOR U21639 ( .A(n22467), .B(n22468), .Z(n22457) );
  XOR U21640 ( .A(n18788), .B(n17633), .Z(n22468) );
  XOR U21641 ( .A(n22469), .B(n22470), .Z(n17633) );
  ANDN U21642 ( .B(n22471), .A(n22472), .Z(n22469) );
  XNOR U21643 ( .A(n22473), .B(n22474), .Z(n18788) );
  ANDN U21644 ( .B(n22475), .A(n22476), .Z(n22473) );
  XNOR U21645 ( .A(n22477), .B(n17439), .Z(n15202) );
  XOR U21646 ( .A(n22478), .B(n13927), .Z(n10707) );
  XOR U21647 ( .A(n22479), .B(n16465), .Z(n13927) );
  XNOR U21648 ( .A(n22480), .B(n22481), .Z(n19906) );
  XOR U21649 ( .A(n19388), .B(n17440), .Z(n22481) );
  XOR U21650 ( .A(n22482), .B(n22483), .Z(n17440) );
  ANDN U21651 ( .B(n22484), .A(n22485), .Z(n22482) );
  XNOR U21652 ( .A(n22486), .B(n22487), .Z(n19388) );
  ANDN U21653 ( .B(n22488), .A(n22489), .Z(n22486) );
  XNOR U21654 ( .A(n17846), .B(n22490), .Z(n22480) );
  XNOR U21655 ( .A(n19630), .B(n19004), .Z(n22490) );
  XNOR U21656 ( .A(n22491), .B(n22492), .Z(n19004) );
  XNOR U21657 ( .A(n22495), .B(n22496), .Z(n19630) );
  ANDN U21658 ( .B(n22497), .A(n22498), .Z(n22495) );
  XNOR U21659 ( .A(n22499), .B(n22500), .Z(n17846) );
  AND U21660 ( .A(n22501), .B(n22502), .Z(n22499) );
  AND U21661 ( .A(n13926), .B(n15215), .Z(n22478) );
  XNOR U21662 ( .A(n20361), .B(n17555), .Z(n15215) );
  XNOR U21663 ( .A(n19901), .B(n22504), .Z(n17555) );
  XOR U21664 ( .A(n22505), .B(n22506), .Z(n19901) );
  XOR U21665 ( .A(n17772), .B(n21992), .Z(n22506) );
  XOR U21666 ( .A(n22507), .B(n22010), .Z(n21992) );
  AND U21667 ( .A(n20352), .B(n20350), .Z(n22507) );
  XOR U21668 ( .A(round_reg[787]), .B(n22508), .Z(n20350) );
  XNOR U21669 ( .A(n22509), .B(n22510), .Z(n17772) );
  AND U21670 ( .A(n20335), .B(n20333), .Z(n22509) );
  XOR U21671 ( .A(n17478), .B(n22511), .Z(n22505) );
  XNOR U21672 ( .A(n16334), .B(n15524), .Z(n22511) );
  XNOR U21673 ( .A(n22512), .B(n22013), .Z(n15524) );
  ANDN U21674 ( .B(n20348), .A(n20346), .Z(n22512) );
  XNOR U21675 ( .A(round_reg[884]), .B(n22513), .Z(n20346) );
  XNOR U21676 ( .A(n22514), .B(n22021), .Z(n16334) );
  AND U21677 ( .A(n20339), .B(n20337), .Z(n22514) );
  XOR U21678 ( .A(round_reg[741]), .B(n22515), .Z(n20337) );
  XNOR U21679 ( .A(n22516), .B(n22018), .Z(n17478) );
  AND U21680 ( .A(n20344), .B(n20342), .Z(n22516) );
  XOR U21681 ( .A(round_reg[955]), .B(n22517), .Z(n20342) );
  XNOR U21682 ( .A(n22518), .B(n22519), .Z(n20361) );
  ANDN U21683 ( .B(n20589), .A(n22520), .Z(n22518) );
  XNOR U21684 ( .A(n17198), .B(n22521), .Z(n13926) );
  XOR U21685 ( .A(n22522), .B(n19528), .Z(n17198) );
  XOR U21686 ( .A(n22523), .B(n22524), .Z(n19528) );
  XOR U21687 ( .A(n19284), .B(n19639), .Z(n22524) );
  XOR U21688 ( .A(n22525), .B(n20407), .Z(n19639) );
  ANDN U21689 ( .B(n20408), .A(n22526), .Z(n22525) );
  XOR U21690 ( .A(n22527), .B(n22528), .Z(n19284) );
  ANDN U21691 ( .B(n22529), .A(n22530), .Z(n22527) );
  XOR U21692 ( .A(n19066), .B(n22531), .Z(n22523) );
  XOR U21693 ( .A(n17143), .B(n18332), .Z(n22531) );
  XNOR U21694 ( .A(n22532), .B(n20412), .Z(n18332) );
  NOR U21695 ( .A(n20411), .B(n22533), .Z(n22532) );
  XNOR U21696 ( .A(n22534), .B(n20415), .Z(n17143) );
  ANDN U21697 ( .B(n20416), .A(n22535), .Z(n22534) );
  XNOR U21698 ( .A(n22536), .B(n20402), .Z(n19066) );
  ANDN U21699 ( .B(n20403), .A(n22537), .Z(n22536) );
  XOR U21700 ( .A(n22538), .B(n22539), .Z(n16199) );
  XOR U21701 ( .A(n11670), .B(n14349), .Z(n22539) );
  XOR U21702 ( .A(n22540), .B(n14368), .Z(n14349) );
  XNOR U21703 ( .A(n17914), .B(n22541), .Z(n14368) );
  XOR U21704 ( .A(n20241), .B(n19328), .Z(n17914) );
  XNOR U21705 ( .A(n22542), .B(n22543), .Z(n19328) );
  XNOR U21706 ( .A(n20235), .B(n18372), .Z(n22543) );
  XNOR U21707 ( .A(n22544), .B(n22545), .Z(n18372) );
  XNOR U21708 ( .A(n22548), .B(n22549), .Z(n20235) );
  XOR U21709 ( .A(n22550), .B(n22551), .Z(n22549) );
  NAND U21710 ( .A(n4640), .B(n6454), .Z(n22551) );
  AND U21711 ( .A(n15691), .B(n6836), .Z(n6454) );
  AND U21712 ( .A(n22552), .B(n22553), .Z(n22550) );
  XOR U21713 ( .A(n18794), .B(n22554), .Z(n22542) );
  XOR U21714 ( .A(n18713), .B(n17468), .Z(n22554) );
  XNOR U21715 ( .A(n22555), .B(n22556), .Z(n17468) );
  ANDN U21716 ( .B(n22557), .A(n22558), .Z(n22555) );
  XNOR U21717 ( .A(n22559), .B(n22560), .Z(n18713) );
  ANDN U21718 ( .B(n22561), .A(n22562), .Z(n22559) );
  XNOR U21719 ( .A(n22563), .B(n22564), .Z(n18794) );
  ANDN U21720 ( .B(n22565), .A(n22566), .Z(n22563) );
  XOR U21721 ( .A(n22567), .B(n22568), .Z(n20241) );
  XOR U21722 ( .A(n22569), .B(n18878), .Z(n22568) );
  XOR U21723 ( .A(n22570), .B(n22472), .Z(n18878) );
  ANDN U21724 ( .B(n22571), .A(n22572), .Z(n22570) );
  XOR U21725 ( .A(n19553), .B(n22573), .Z(n22567) );
  XOR U21726 ( .A(n22574), .B(n17977), .Z(n22573) );
  XOR U21727 ( .A(n22575), .B(n22466), .Z(n17977) );
  IV U21728 ( .A(n22576), .Z(n22466) );
  ANDN U21729 ( .B(n22577), .A(n22578), .Z(n22575) );
  XNOR U21730 ( .A(n22579), .B(n22462), .Z(n19553) );
  ANDN U21731 ( .B(n22580), .A(n22581), .Z(n22579) );
  ANDN U21732 ( .B(n14787), .A(n14369), .Z(n22540) );
  XOR U21733 ( .A(n19278), .B(n18730), .Z(n14369) );
  IV U21734 ( .A(n17434), .Z(n18730) );
  XNOR U21735 ( .A(n22582), .B(n20754), .Z(n19278) );
  ANDN U21736 ( .B(n22583), .A(n22584), .Z(n22582) );
  XNOR U21737 ( .A(n22587), .B(n22588), .Z(n20959) );
  ANDN U21738 ( .B(n22589), .A(n21890), .Z(n22587) );
  XNOR U21739 ( .A(n22590), .B(n19204), .Z(n11670) );
  XOR U21740 ( .A(n18527), .B(n22591), .Z(n19204) );
  AND U21741 ( .A(n14790), .B(n17741), .Z(n22590) );
  XNOR U21742 ( .A(n15626), .B(n21860), .Z(n17741) );
  XOR U21743 ( .A(n22592), .B(n22593), .Z(n21860) );
  ANDN U21744 ( .B(n22594), .A(n22595), .Z(n22592) );
  IV U21745 ( .A(n17226), .Z(n15626) );
  XOR U21746 ( .A(n20425), .B(n19283), .Z(n17226) );
  XNOR U21747 ( .A(n22596), .B(n22597), .Z(n19283) );
  XOR U21748 ( .A(n19487), .B(n18384), .Z(n22597) );
  XNOR U21749 ( .A(n22598), .B(n22235), .Z(n18384) );
  AND U21750 ( .A(n22599), .B(n22600), .Z(n22598) );
  XNOR U21751 ( .A(n22601), .B(n20676), .Z(n19487) );
  AND U21752 ( .A(n22602), .B(n22603), .Z(n22601) );
  XOR U21753 ( .A(n19614), .B(n22604), .Z(n22596) );
  XNOR U21754 ( .A(n17473), .B(n19307), .Z(n22604) );
  XNOR U21755 ( .A(n22605), .B(n20682), .Z(n19307) );
  AND U21756 ( .A(n22606), .B(n22607), .Z(n22605) );
  XNOR U21757 ( .A(n22608), .B(n22609), .Z(n17473) );
  AND U21758 ( .A(n22610), .B(n22611), .Z(n22608) );
  XNOR U21759 ( .A(n22612), .B(n20685), .Z(n19614) );
  AND U21760 ( .A(n22613), .B(n22614), .Z(n22612) );
  XOR U21761 ( .A(n22615), .B(n22616), .Z(n20425) );
  XNOR U21762 ( .A(n22617), .B(n17886), .Z(n22616) );
  XOR U21763 ( .A(n22618), .B(n22619), .Z(n17886) );
  NOR U21764 ( .A(n21867), .B(n21868), .Z(n22618) );
  XOR U21765 ( .A(n17838), .B(n22620), .Z(n22615) );
  XNOR U21766 ( .A(n18456), .B(n16697), .Z(n22620) );
  XNOR U21767 ( .A(n22621), .B(n22622), .Z(n16697) );
  ANDN U21768 ( .B(n22623), .A(n22594), .Z(n22621) );
  XNOR U21769 ( .A(n22624), .B(n22625), .Z(n18456) );
  ANDN U21770 ( .B(n21857), .A(n21859), .Z(n22624) );
  XNOR U21771 ( .A(n22626), .B(n22627), .Z(n17838) );
  AND U21772 ( .A(n21864), .B(n21863), .Z(n22626) );
  XNOR U21773 ( .A(n22629), .B(n22630), .Z(n17439) );
  XOR U21774 ( .A(n10924), .B(n22631), .Z(n22538) );
  XOR U21775 ( .A(n12983), .B(n11322), .Z(n22631) );
  XOR U21776 ( .A(n22632), .B(n19225), .Z(n11322) );
  XOR U21777 ( .A(n16268), .B(n22015), .Z(n19225) );
  XOR U21778 ( .A(n22633), .B(n22634), .Z(n22015) );
  ANDN U21779 ( .B(n22510), .A(n20333), .Z(n22633) );
  XOR U21780 ( .A(round_reg[663]), .B(n22635), .Z(n20333) );
  IV U21781 ( .A(n17006), .Z(n16268) );
  XOR U21782 ( .A(n22636), .B(n20604), .Z(n17006) );
  XNOR U21783 ( .A(n22637), .B(n22638), .Z(n20604) );
  XOR U21784 ( .A(n18742), .B(n21073), .Z(n22638) );
  XOR U21785 ( .A(n22639), .B(n20347), .Z(n21073) );
  XNOR U21786 ( .A(round_reg[1242]), .B(n22640), .Z(n22013) );
  XOR U21787 ( .A(n22641), .B(n20338), .Z(n18742) );
  ANDN U21788 ( .B(n22020), .A(n22021), .Z(n22641) );
  XOR U21789 ( .A(round_reg[1144]), .B(n22642), .Z(n22021) );
  XOR U21790 ( .A(n17525), .B(n22643), .Z(n22637) );
  XOR U21791 ( .A(n16668), .B(n18191), .Z(n22643) );
  XNOR U21792 ( .A(n22644), .B(n20351), .Z(n18191) );
  ANDN U21793 ( .B(n22009), .A(n22010), .Z(n22644) );
  XOR U21794 ( .A(round_reg[1170]), .B(n22645), .Z(n22010) );
  XOR U21795 ( .A(n22646), .B(n20334), .Z(n16668) );
  ANDN U21796 ( .B(n22647), .A(n22510), .Z(n22646) );
  XOR U21797 ( .A(round_reg[1031]), .B(n21316), .Z(n22510) );
  XOR U21798 ( .A(n22648), .B(n20343), .Z(n17525) );
  NOR U21799 ( .A(n22018), .B(n22017), .Z(n22648) );
  XOR U21800 ( .A(round_reg[1002]), .B(n22649), .Z(n22018) );
  ANDN U21801 ( .B(n14361), .A(n14794), .Z(n22632) );
  XNOR U21802 ( .A(n17126), .B(n21776), .Z(n14794) );
  XNOR U21803 ( .A(n22650), .B(n22651), .Z(n21776) );
  ANDN U21804 ( .B(n20643), .A(n19691), .Z(n22650) );
  XNOR U21805 ( .A(round_reg[141]), .B(n22652), .Z(n19691) );
  IV U21806 ( .A(n19612), .Z(n17126) );
  XOR U21807 ( .A(n22522), .B(n22653), .Z(n19612) );
  XOR U21808 ( .A(n22654), .B(n22655), .Z(n22522) );
  XNOR U21809 ( .A(n20395), .B(n19666), .Z(n22655) );
  XOR U21810 ( .A(n22656), .B(n22657), .Z(n19666) );
  ANDN U21811 ( .B(n22658), .A(n22659), .Z(n22656) );
  XNOR U21812 ( .A(n22660), .B(n22661), .Z(n20395) );
  ANDN U21813 ( .B(n22662), .A(n22663), .Z(n22660) );
  XNOR U21814 ( .A(n20323), .B(n22664), .Z(n22654) );
  XOR U21815 ( .A(n17074), .B(n18363), .Z(n22664) );
  XOR U21816 ( .A(n22665), .B(n22666), .Z(n18363) );
  ANDN U21817 ( .B(n22667), .A(n22668), .Z(n22665) );
  XNOR U21818 ( .A(n22669), .B(n22670), .Z(n17074) );
  NOR U21819 ( .A(n22671), .B(n22672), .Z(n22669) );
  XNOR U21820 ( .A(n22673), .B(n22674), .Z(n20323) );
  ANDN U21821 ( .B(n22675), .A(n22676), .Z(n22673) );
  XOR U21822 ( .A(n17328), .B(n22677), .Z(n14361) );
  IV U21823 ( .A(n18193), .Z(n17328) );
  XNOR U21824 ( .A(n22678), .B(n14355), .Z(n12983) );
  XNOR U21825 ( .A(n13886), .B(n21982), .Z(n14355) );
  XNOR U21826 ( .A(n22679), .B(n22680), .Z(n21982) );
  ANDN U21827 ( .B(n22681), .A(n22682), .Z(n22679) );
  IV U21828 ( .A(n19310), .Z(n13886) );
  XOR U21829 ( .A(n18598), .B(n22683), .Z(n19310) );
  XOR U21830 ( .A(n22684), .B(n22685), .Z(n18598) );
  XNOR U21831 ( .A(n18785), .B(n18642), .Z(n22685) );
  XOR U21832 ( .A(n22686), .B(n22057), .Z(n18642) );
  AND U21833 ( .A(n21957), .B(n21955), .Z(n22686) );
  XOR U21834 ( .A(round_reg[1559]), .B(n22687), .Z(n21955) );
  XNOR U21835 ( .A(n22688), .B(n22054), .Z(n18785) );
  ANDN U21836 ( .B(n21964), .A(n21965), .Z(n22688) );
  XOR U21837 ( .A(round_reg[1433]), .B(n21613), .Z(n21964) );
  XNOR U21838 ( .A(n19135), .B(n22689), .Z(n22684) );
  XOR U21839 ( .A(n21657), .B(n22025), .Z(n22689) );
  XNOR U21840 ( .A(n22690), .B(n22047), .Z(n22025) );
  AND U21841 ( .A(n21970), .B(n21968), .Z(n22690) );
  XOR U21842 ( .A(round_reg[1494]), .B(n22691), .Z(n21968) );
  XNOR U21843 ( .A(n22692), .B(n22044), .Z(n21657) );
  AND U21844 ( .A(n21962), .B(n21960), .Z(n22692) );
  XOR U21845 ( .A(round_reg[1340]), .B(n21772), .Z(n21960) );
  XNOR U21846 ( .A(n22693), .B(n22051), .Z(n19135) );
  ANDN U21847 ( .B(n21951), .A(n21953), .Z(n22693) );
  XOR U21848 ( .A(round_reg[1403]), .B(n22369), .Z(n21951) );
  ANDN U21849 ( .B(n14356), .A(n17712), .Z(n22678) );
  XOR U21850 ( .A(n19263), .B(n20693), .Z(n17712) );
  XNOR U21851 ( .A(n22694), .B(n21233), .Z(n20693) );
  ANDN U21852 ( .B(n20172), .A(n20173), .Z(n22694) );
  XOR U21853 ( .A(n22695), .B(n22696), .Z(n19263) );
  XOR U21854 ( .A(n16348), .B(n22697), .Z(n14356) );
  XNOR U21855 ( .A(n22698), .B(n14364), .Z(n10924) );
  XNOR U21856 ( .A(n18181), .B(n22699), .Z(n14364) );
  ANDN U21857 ( .B(n14365), .A(n14783), .Z(n22698) );
  XNOR U21858 ( .A(n21815), .B(n17186), .Z(n14783) );
  XNOR U21859 ( .A(n22700), .B(n22701), .Z(n17186) );
  XNOR U21860 ( .A(n22702), .B(n22400), .Z(n21815) );
  AND U21861 ( .A(n22703), .B(n22704), .Z(n22702) );
  XOR U21862 ( .A(n22705), .B(n19156), .Z(n14365) );
  XOR U21863 ( .A(n21927), .B(n20711), .Z(n19156) );
  XNOR U21864 ( .A(n22706), .B(n22707), .Z(n20711) );
  XOR U21865 ( .A(n18116), .B(n19821), .Z(n22707) );
  XNOR U21866 ( .A(n22708), .B(n22709), .Z(n19821) );
  ANDN U21867 ( .B(n22710), .A(n22711), .Z(n22708) );
  XNOR U21868 ( .A(n22712), .B(n22713), .Z(n18116) );
  ANDN U21869 ( .B(n22714), .A(n22715), .Z(n22712) );
  XOR U21870 ( .A(n21361), .B(n22716), .Z(n22706) );
  XOR U21871 ( .A(n20233), .B(n15587), .Z(n22716) );
  XNOR U21872 ( .A(n22717), .B(n22718), .Z(n15587) );
  NOR U21873 ( .A(n22719), .B(n22720), .Z(n22717) );
  XNOR U21874 ( .A(n22721), .B(n22722), .Z(n20233) );
  ANDN U21875 ( .B(n22723), .A(n22724), .Z(n22721) );
  XOR U21876 ( .A(n22725), .B(n22726), .Z(n21361) );
  ANDN U21877 ( .B(n22727), .A(n22728), .Z(n22725) );
  XOR U21878 ( .A(n22729), .B(n22730), .Z(n21927) );
  XNOR U21879 ( .A(n21787), .B(n18322), .Z(n22730) );
  XOR U21880 ( .A(n22731), .B(n22732), .Z(n18322) );
  ANDN U21881 ( .B(n22733), .A(n22734), .Z(n22731) );
  XNOR U21882 ( .A(n22735), .B(n22736), .Z(n21787) );
  ANDN U21883 ( .B(n22737), .A(n22738), .Z(n22735) );
  XNOR U21884 ( .A(n22739), .B(n22740), .Z(n22729) );
  XOR U21885 ( .A(n18820), .B(n18647), .Z(n22740) );
  XOR U21886 ( .A(n22741), .B(n22742), .Z(n18647) );
  AND U21887 ( .A(n22743), .B(n22744), .Z(n22741) );
  XNOR U21888 ( .A(n22745), .B(n22746), .Z(n18820) );
  NOR U21889 ( .A(n22747), .B(n22748), .Z(n22745) );
  XNOR U21890 ( .A(n22749), .B(n13923), .Z(n17530) );
  XNOR U21891 ( .A(n20574), .B(n16414), .Z(n13923) );
  IV U21892 ( .A(n18270), .Z(n16414) );
  XNOR U21893 ( .A(n22750), .B(n20103), .Z(n20574) );
  AND U21894 ( .A(n19868), .B(n21612), .Z(n22750) );
  IV U21895 ( .A(n19870), .Z(n21612) );
  XOR U21896 ( .A(round_reg[862]), .B(n22751), .Z(n19870) );
  IV U21897 ( .A(n22752), .Z(n19868) );
  ANDN U21898 ( .B(n15211), .A(n13092), .Z(n22749) );
  XNOR U21899 ( .A(n18181), .B(n22753), .Z(n13092) );
  IV U21900 ( .A(n22143), .Z(n18181) );
  XOR U21901 ( .A(n18866), .B(n21478), .Z(n22143) );
  XNOR U21902 ( .A(n22754), .B(n22755), .Z(n21478) );
  XOR U21903 ( .A(n19073), .B(n16251), .Z(n22755) );
  XOR U21904 ( .A(n22756), .B(n21859), .Z(n16251) );
  XOR U21905 ( .A(round_reg[451]), .B(n22757), .Z(n21859) );
  ANDN U21906 ( .B(n22758), .A(n21858), .Z(n22756) );
  XNOR U21907 ( .A(n22759), .B(n21868), .Z(n19073) );
  XOR U21908 ( .A(round_reg[617]), .B(n22760), .Z(n21868) );
  ANDN U21909 ( .B(n21869), .A(n22761), .Z(n22759) );
  XNOR U21910 ( .A(n16357), .B(n22762), .Z(n22754) );
  XOR U21911 ( .A(n16423), .B(n17817), .Z(n22762) );
  XNOR U21912 ( .A(n22763), .B(n22594), .Z(n17817) );
  XNOR U21913 ( .A(round_reg[445]), .B(n22764), .Z(n22594) );
  ANDN U21914 ( .B(n22595), .A(n22765), .Z(n22763) );
  XNOR U21915 ( .A(n22766), .B(n21854), .Z(n16423) );
  ANDN U21916 ( .B(n21855), .A(n22767), .Z(n22766) );
  XNOR U21917 ( .A(n22768), .B(n21864), .Z(n16357) );
  XNOR U21918 ( .A(round_reg[549]), .B(n22769), .Z(n21864) );
  AND U21919 ( .A(n22770), .B(n21865), .Z(n22768) );
  XOR U21920 ( .A(n22771), .B(n22772), .Z(n18866) );
  XOR U21921 ( .A(n17995), .B(n17944), .Z(n22772) );
  XOR U21922 ( .A(n22773), .B(n20435), .Z(n17944) );
  XOR U21923 ( .A(round_reg[1052]), .B(n22119), .Z(n20435) );
  ANDN U21924 ( .B(n21845), .A(n22774), .Z(n22773) );
  XOR U21925 ( .A(n22775), .B(n21848), .Z(n17995) );
  ANDN U21926 ( .B(n21849), .A(n22776), .Z(n22775) );
  XOR U21927 ( .A(n21830), .B(n22777), .Z(n22771) );
  XNOR U21928 ( .A(n18586), .B(n18699), .Z(n22777) );
  XNOR U21929 ( .A(n22778), .B(n20431), .Z(n18699) );
  XOR U21930 ( .A(round_reg[1191]), .B(n22361), .Z(n20431) );
  AND U21931 ( .A(n22779), .B(n21835), .Z(n22778) );
  XOR U21932 ( .A(n22780), .B(n21841), .Z(n18586) );
  ANDN U21933 ( .B(n21842), .A(n22781), .Z(n22780) );
  XNOR U21934 ( .A(n22782), .B(n20441), .Z(n21830) );
  XOR U21935 ( .A(round_reg[1023]), .B(n22783), .Z(n20441) );
  AND U21936 ( .A(n22784), .B(n21837), .Z(n22782) );
  IV U21937 ( .A(n22450), .Z(n15211) );
  XOR U21938 ( .A(n18193), .B(n22785), .Z(n22450) );
  XNOR U21939 ( .A(n22787), .B(n22788), .Z(n20739) );
  XNOR U21940 ( .A(n17527), .B(n16904), .Z(n22788) );
  XNOR U21941 ( .A(n22789), .B(n21415), .Z(n16904) );
  XOR U21942 ( .A(round_reg[1425]), .B(n22790), .Z(n21415) );
  ANDN U21943 ( .B(n21416), .A(n22791), .Z(n22789) );
  XNOR U21944 ( .A(n22792), .B(n21420), .Z(n17527) );
  XOR U21945 ( .A(round_reg[1486]), .B(n22221), .Z(n21420) );
  ANDN U21946 ( .B(n21421), .A(n22793), .Z(n22792) );
  XOR U21947 ( .A(n19926), .B(n22794), .Z(n22787) );
  XOR U21948 ( .A(n19231), .B(n17273), .Z(n22794) );
  XNOR U21949 ( .A(n22795), .B(n21424), .Z(n17273) );
  XOR U21950 ( .A(round_reg[1332]), .B(n22796), .Z(n21424) );
  AND U21951 ( .A(n21425), .B(n22797), .Z(n22795) );
  XOR U21952 ( .A(n21411), .B(n22798), .Z(n19231) );
  XOR U21953 ( .A(n22799), .B(n22800), .Z(n22798) );
  NAND U21954 ( .A(n4656), .B(n4510), .Z(n22800) );
  AND U21955 ( .A(n6836), .B(n11365), .Z(n4510) );
  IV U21956 ( .A(rc_i[4]), .Z(n6836) );
  AND U21957 ( .A(n15691), .B(n11363), .Z(n4656) );
  ANDN U21958 ( .B(n21412), .A(n22801), .Z(n22799) );
  XOR U21959 ( .A(round_reg[1551]), .B(n22802), .Z(n21411) );
  XNOR U21960 ( .A(n22803), .B(n21428), .Z(n19926) );
  ANDN U21961 ( .B(n21429), .A(n22804), .Z(n22803) );
  XOR U21962 ( .A(n10142), .B(n17303), .Z(n9196) );
  XOR U21963 ( .A(n22805), .B(n19792), .Z(n17303) );
  AND U21964 ( .A(n18229), .B(n22806), .Z(n22805) );
  XNOR U21965 ( .A(n22574), .B(n18879), .Z(n18229) );
  XNOR U21966 ( .A(n22807), .B(n22476), .Z(n22574) );
  ANDN U21967 ( .B(n22808), .A(n22809), .Z(n22807) );
  XOR U21968 ( .A(n18414), .B(n16959), .Z(n10142) );
  XOR U21969 ( .A(n22810), .B(n22811), .Z(n16959) );
  XOR U21970 ( .A(n11723), .B(n11848), .Z(n22811) );
  XOR U21971 ( .A(n22812), .B(n17700), .Z(n11848) );
  XNOR U21972 ( .A(n20387), .B(n18494), .Z(n17700) );
  IV U21973 ( .A(n16451), .Z(n18494) );
  XNOR U21974 ( .A(n18392), .B(n20687), .Z(n16451) );
  XNOR U21975 ( .A(n22813), .B(n22814), .Z(n20687) );
  XNOR U21976 ( .A(n22320), .B(n18550), .Z(n22814) );
  XOR U21977 ( .A(n22815), .B(n22333), .Z(n18550) );
  XNOR U21978 ( .A(round_reg[1574]), .B(n22432), .Z(n20144) );
  XOR U21979 ( .A(round_reg[24]), .B(n22816), .Z(n20419) );
  XOR U21980 ( .A(n22817), .B(n22384), .Z(n22320) );
  XOR U21981 ( .A(round_reg[1509]), .B(n22769), .Z(n20161) );
  XOR U21982 ( .A(round_reg[276]), .B(n22818), .Z(n20390) );
  XOR U21983 ( .A(n19796), .B(n22819), .Z(n22813) );
  XNOR U21984 ( .A(n17982), .B(n17973), .Z(n22819) );
  XOR U21985 ( .A(n22820), .B(n22325), .Z(n17973) );
  NOR U21986 ( .A(n20392), .B(n20157), .Z(n22820) );
  XOR U21987 ( .A(round_reg[1448]), .B(n22821), .Z(n20157) );
  XOR U21988 ( .A(round_reg[228]), .B(n22822), .Z(n20392) );
  XNOR U21989 ( .A(n22823), .B(n22329), .Z(n17982) );
  ANDN U21990 ( .B(n22328), .A(n20148), .Z(n22823) );
  XOR U21991 ( .A(n22824), .B(n22331), .Z(n19796) );
  ANDN U21992 ( .B(n20386), .A(n20153), .Z(n22824) );
  XOR U21993 ( .A(round_reg[1291]), .B(n21754), .Z(n20153) );
  XOR U21994 ( .A(round_reg[110]), .B(n22825), .Z(n20386) );
  XNOR U21995 ( .A(n22826), .B(n22827), .Z(n18392) );
  XNOR U21996 ( .A(n18784), .B(n16354), .Z(n22827) );
  XOR U21997 ( .A(n22828), .B(n22349), .Z(n16354) );
  NOR U21998 ( .A(n20874), .B(n20873), .Z(n22828) );
  XNOR U21999 ( .A(round_reg[977]), .B(n22829), .Z(n20873) );
  XOR U22000 ( .A(n22830), .B(n22338), .Z(n18784) );
  ANDN U22001 ( .B(n20865), .A(n20866), .Z(n22830) );
  XOR U22002 ( .A(round_reg[1209]), .B(n22831), .Z(n20865) );
  XNOR U22003 ( .A(n17572), .B(n22832), .Z(n22826) );
  XNOR U22004 ( .A(n20461), .B(n16068), .Z(n22832) );
  XOR U22005 ( .A(n22833), .B(n22341), .Z(n16068) );
  NOR U22006 ( .A(n20870), .B(n20869), .Z(n22833) );
  XNOR U22007 ( .A(round_reg[1217]), .B(n22834), .Z(n20869) );
  XNOR U22008 ( .A(n22835), .B(n22346), .Z(n20461) );
  NOR U22009 ( .A(n20857), .B(n20856), .Z(n22835) );
  XNOR U22010 ( .A(round_reg[1070]), .B(n22825), .Z(n20856) );
  XNOR U22011 ( .A(n22836), .B(n22837), .Z(n17572) );
  NOR U22012 ( .A(n20860), .B(n20861), .Z(n22836) );
  XNOR U22013 ( .A(n22838), .B(n22328), .Z(n20387) );
  ANDN U22014 ( .B(n20148), .A(n20149), .Z(n22838) );
  XOR U22015 ( .A(round_reg[1354]), .B(n22839), .Z(n20148) );
  ANDN U22016 ( .B(n17310), .A(n17311), .Z(n22812) );
  XNOR U22017 ( .A(n19234), .B(n22840), .Z(n17311) );
  IV U22018 ( .A(n15592), .Z(n19234) );
  XOR U22019 ( .A(n18971), .B(n18749), .Z(n15592) );
  XNOR U22020 ( .A(n22841), .B(n22842), .Z(n18749) );
  XOR U22021 ( .A(n19532), .B(n17508), .Z(n22842) );
  XNOR U22022 ( .A(n22843), .B(n22844), .Z(n17508) );
  ANDN U22023 ( .B(n21576), .A(n22845), .Z(n22843) );
  XOR U22024 ( .A(n22846), .B(n22847), .Z(n19532) );
  XNOR U22025 ( .A(n18024), .B(n22849), .Z(n22841) );
  XOR U22026 ( .A(n19079), .B(n22850), .Z(n22849) );
  XNOR U22027 ( .A(n22851), .B(n22852), .Z(n19079) );
  ANDN U22028 ( .B(n20887), .A(n22853), .Z(n22851) );
  XNOR U22029 ( .A(n22854), .B(n22855), .Z(n18024) );
  ANDN U22030 ( .B(n20897), .A(n22856), .Z(n22854) );
  XOR U22031 ( .A(n22857), .B(n22858), .Z(n18971) );
  XNOR U22032 ( .A(n19208), .B(n14909), .Z(n22858) );
  XNOR U22033 ( .A(n22859), .B(n22860), .Z(n14909) );
  AND U22034 ( .A(n22861), .B(n22862), .Z(n22859) );
  XNOR U22035 ( .A(n22863), .B(n22864), .Z(n19208) );
  AND U22036 ( .A(n22865), .B(n22866), .Z(n22863) );
  XOR U22037 ( .A(n15321), .B(n22867), .Z(n22857) );
  XOR U22038 ( .A(n20608), .B(n16022), .Z(n22867) );
  XNOR U22039 ( .A(n22868), .B(n22869), .Z(n16022) );
  AND U22040 ( .A(n22870), .B(n22871), .Z(n22868) );
  XNOR U22041 ( .A(n22872), .B(n22873), .Z(n20608) );
  ANDN U22042 ( .B(n22874), .A(n22875), .Z(n22872) );
  XNOR U22043 ( .A(n22876), .B(n22877), .Z(n15321) );
  ANDN U22044 ( .B(n22878), .A(n22879), .Z(n22876) );
  XOR U22045 ( .A(n22880), .B(n19503), .Z(n17310) );
  IV U22046 ( .A(n15639), .Z(n19503) );
  XOR U22047 ( .A(n22881), .B(n22503), .Z(n15639) );
  XOR U22048 ( .A(n22882), .B(n22883), .Z(n22503) );
  XOR U22049 ( .A(n19678), .B(n22280), .Z(n22883) );
  XOR U22050 ( .A(n22884), .B(n22885), .Z(n22280) );
  ANDN U22051 ( .B(n22886), .A(n22887), .Z(n22884) );
  XOR U22052 ( .A(n22888), .B(n22300), .Z(n19678) );
  ANDN U22053 ( .B(n22299), .A(n22889), .Z(n22888) );
  XNOR U22054 ( .A(n17034), .B(n22890), .Z(n22882) );
  XOR U22055 ( .A(n19422), .B(n19064), .Z(n22890) );
  XOR U22056 ( .A(n22891), .B(n22285), .Z(n19064) );
  ANDN U22057 ( .B(n22286), .A(n22892), .Z(n22891) );
  XOR U22058 ( .A(n22893), .B(n22289), .Z(n19422) );
  XOR U22059 ( .A(n22895), .B(n22295), .Z(n17034) );
  ANDN U22060 ( .B(n22296), .A(n22896), .Z(n22895) );
  XNOR U22061 ( .A(n22897), .B(n17698), .Z(n11723) );
  XNOR U22062 ( .A(n18527), .B(n22898), .Z(n17698) );
  XOR U22063 ( .A(n20606), .B(n20883), .Z(n18527) );
  XOR U22064 ( .A(n22899), .B(n22900), .Z(n20883) );
  XNOR U22065 ( .A(n19111), .B(n17362), .Z(n22900) );
  XNOR U22066 ( .A(n22901), .B(n22878), .Z(n17362) );
  XNOR U22067 ( .A(n22904), .B(n22861), .Z(n19111) );
  IV U22068 ( .A(n22905), .Z(n22861) );
  ANDN U22069 ( .B(n22906), .A(n22907), .Z(n22904) );
  XNOR U22070 ( .A(n18424), .B(n22908), .Z(n22899) );
  XOR U22071 ( .A(n22909), .B(n22910), .Z(n22908) );
  XNOR U22072 ( .A(n22911), .B(n22865), .Z(n18424) );
  XOR U22073 ( .A(n22914), .B(n22915), .Z(n20606) );
  XOR U22074 ( .A(n22353), .B(n21523), .Z(n22915) );
  XOR U22075 ( .A(n22916), .B(n22917), .Z(n21523) );
  ANDN U22076 ( .B(n22918), .A(n22919), .Z(n22916) );
  XNOR U22077 ( .A(n22920), .B(n22921), .Z(n22353) );
  NOR U22078 ( .A(n22922), .B(n22923), .Z(n22920) );
  XOR U22079 ( .A(n18645), .B(n22924), .Z(n22914) );
  XOR U22080 ( .A(n18007), .B(n15605), .Z(n22924) );
  XNOR U22081 ( .A(n22925), .B(n22926), .Z(n15605) );
  ANDN U22082 ( .B(n22927), .A(n22928), .Z(n22925) );
  XNOR U22083 ( .A(n22929), .B(n22930), .Z(n18007) );
  ANDN U22084 ( .B(n22931), .A(n22932), .Z(n22929) );
  XNOR U22085 ( .A(n22933), .B(n22934), .Z(n18645) );
  ANDN U22086 ( .B(n22935), .A(n22936), .Z(n22933) );
  ANDN U22087 ( .B(n17318), .A(n17319), .Z(n22897) );
  XNOR U22088 ( .A(n22937), .B(n20270), .Z(n17319) );
  IV U22089 ( .A(n19703), .Z(n20270) );
  XOR U22090 ( .A(n22938), .B(n16014), .Z(n17318) );
  IV U22091 ( .A(n19685), .Z(n16014) );
  XNOR U22092 ( .A(n18972), .B(n22939), .Z(n19685) );
  XNOR U22093 ( .A(n22940), .B(n22941), .Z(n18972) );
  XOR U22094 ( .A(n22942), .B(n19389), .Z(n22941) );
  XOR U22095 ( .A(n22943), .B(n22944), .Z(n19389) );
  ANDN U22096 ( .B(n22945), .A(n22930), .Z(n22943) );
  XOR U22097 ( .A(n22946), .B(n22947), .Z(n22940) );
  XOR U22098 ( .A(n16766), .B(n16956), .Z(n22947) );
  XNOR U22099 ( .A(n22948), .B(n22949), .Z(n16956) );
  NOR U22100 ( .A(n22950), .B(n22926), .Z(n22948) );
  XNOR U22101 ( .A(n22951), .B(n22952), .Z(n16766) );
  ANDN U22102 ( .B(n22953), .A(n22921), .Z(n22951) );
  XOR U22103 ( .A(n9781), .B(n22954), .Z(n22810) );
  XOR U22104 ( .A(n10732), .B(n10549), .Z(n22954) );
  XNOR U22105 ( .A(n22955), .B(n18231), .Z(n10549) );
  XOR U22106 ( .A(n22028), .B(n18578), .Z(n18231) );
  XOR U22107 ( .A(n20095), .B(n20282), .Z(n18578) );
  XNOR U22108 ( .A(n22956), .B(n22957), .Z(n20282) );
  XNOR U22109 ( .A(n19037), .B(n17193), .Z(n22957) );
  XNOR U22110 ( .A(n22958), .B(n21690), .Z(n17193) );
  XNOR U22111 ( .A(round_reg[1054]), .B(n22959), .Z(n21690) );
  XNOR U22112 ( .A(n22961), .B(n22070), .Z(n19037) );
  XOR U22113 ( .A(round_reg[1265]), .B(n22962), .Z(n22070) );
  XOR U22114 ( .A(n18900), .B(n22964), .Z(n22956) );
  XOR U22115 ( .A(n21675), .B(n18623), .Z(n22964) );
  XOR U22116 ( .A(n22965), .B(n21681), .Z(n18623) );
  XOR U22117 ( .A(round_reg[961]), .B(n22966), .Z(n21681) );
  XOR U22118 ( .A(n22968), .B(n21695), .Z(n21675) );
  XOR U22119 ( .A(round_reg[1103]), .B(n22969), .Z(n21695) );
  NOR U22120 ( .A(n21694), .B(n22970), .Z(n22968) );
  XOR U22121 ( .A(n22971), .B(n21684), .Z(n18900) );
  XNOR U22122 ( .A(round_reg[1193]), .B(n22972), .Z(n21684) );
  ANDN U22123 ( .B(n21685), .A(n22973), .Z(n22971) );
  XOR U22124 ( .A(n22974), .B(n22975), .Z(n20095) );
  XOR U22125 ( .A(n19332), .B(n18327), .Z(n22975) );
  XNOR U22126 ( .A(n22976), .B(n19760), .Z(n18327) );
  XOR U22127 ( .A(round_reg[8]), .B(n22977), .Z(n19760) );
  AND U22128 ( .A(n22032), .B(n22030), .Z(n22976) );
  XOR U22129 ( .A(round_reg[1558]), .B(n22225), .Z(n22030) );
  XOR U22130 ( .A(n22978), .B(n19755), .Z(n19332) );
  XNOR U22131 ( .A(round_reg[212]), .B(n22979), .Z(n19755) );
  ANDN U22132 ( .B(n22037), .A(n19754), .Z(n22978) );
  XNOR U22133 ( .A(round_reg[1432]), .B(n22980), .Z(n19754) );
  XNOR U22134 ( .A(n17488), .B(n22981), .Z(n22974) );
  XOR U22135 ( .A(n19745), .B(n17239), .Z(n22981) );
  XNOR U22136 ( .A(n22982), .B(n19764), .Z(n17239) );
  XNOR U22137 ( .A(round_reg[260]), .B(n22983), .Z(n19764) );
  ANDN U22138 ( .B(n22039), .A(n19763), .Z(n22982) );
  XNOR U22139 ( .A(round_reg[1493]), .B(n22984), .Z(n19763) );
  XNOR U22140 ( .A(n22985), .B(n19751), .Z(n19745) );
  XOR U22141 ( .A(round_reg[94]), .B(n22959), .Z(n19751) );
  XNOR U22142 ( .A(round_reg[1339]), .B(n22986), .Z(n19750) );
  XNOR U22143 ( .A(n22987), .B(n19768), .Z(n17488) );
  AND U22144 ( .A(n22988), .B(n19767), .Z(n22987) );
  IV U22145 ( .A(n22989), .Z(n19767) );
  XOR U22146 ( .A(n22990), .B(n22989), .Z(n22028) );
  XNOR U22147 ( .A(round_reg[1402]), .B(n22991), .Z(n22989) );
  ANDN U22148 ( .B(n22992), .A(n22988), .Z(n22990) );
  AND U22149 ( .A(n19586), .B(n19792), .Z(n22955) );
  XOR U22150 ( .A(n18046), .B(n22993), .Z(n19792) );
  IV U22151 ( .A(n22806), .Z(n19586) );
  XOR U22152 ( .A(n21334), .B(n15325), .Z(n22806) );
  XOR U22153 ( .A(n22696), .B(n22426), .Z(n15325) );
  XNOR U22154 ( .A(n22994), .B(n22995), .Z(n22426) );
  XNOR U22155 ( .A(n20779), .B(n18465), .Z(n22995) );
  XNOR U22156 ( .A(n22996), .B(n22997), .Z(n18465) );
  ANDN U22157 ( .B(n21360), .A(n21358), .Z(n22996) );
  XOR U22158 ( .A(n22998), .B(n22999), .Z(n20779) );
  NOR U22159 ( .A(n21344), .B(n21345), .Z(n22998) );
  XOR U22160 ( .A(n20941), .B(n23000), .Z(n22994) );
  XOR U22161 ( .A(n18572), .B(n23001), .Z(n23000) );
  XOR U22162 ( .A(n23002), .B(n23003), .Z(n18572) );
  NOR U22163 ( .A(n22449), .B(n22447), .Z(n23002) );
  XOR U22164 ( .A(n23004), .B(n23005), .Z(n20941) );
  ANDN U22165 ( .B(n21356), .A(n21354), .Z(n23004) );
  XNOR U22166 ( .A(n23006), .B(n23007), .Z(n22696) );
  XNOR U22167 ( .A(n19294), .B(n18875), .Z(n23007) );
  XOR U22168 ( .A(n23008), .B(n21252), .Z(n18875) );
  ANDN U22169 ( .B(n21340), .A(n21251), .Z(n23008) );
  XOR U22170 ( .A(round_reg[936]), .B(n23009), .Z(n21251) );
  XNOR U22171 ( .A(n23010), .B(n21238), .Z(n19294) );
  XNOR U22172 ( .A(round_reg[768]), .B(n23011), .Z(n21239) );
  XOR U22173 ( .A(n18967), .B(n23012), .Z(n23006) );
  XOR U22174 ( .A(n19320), .B(n18161), .Z(n23012) );
  XOR U22175 ( .A(n23013), .B(n21256), .Z(n18161) );
  ANDN U22176 ( .B(n23014), .A(n21255), .Z(n23013) );
  XNOR U22177 ( .A(n23015), .B(n21242), .Z(n19320) );
  AND U22178 ( .A(n21329), .B(n21243), .Z(n23015) );
  XOR U22179 ( .A(round_reg[644]), .B(n23016), .Z(n21243) );
  XNOR U22180 ( .A(n23017), .B(n21248), .Z(n18967) );
  ANDN U22181 ( .B(n21332), .A(n21247), .Z(n23017) );
  XNOR U22182 ( .A(round_reg[722]), .B(n21786), .Z(n21247) );
  XNOR U22183 ( .A(n23018), .B(n21255), .Z(n21334) );
  XOR U22184 ( .A(round_reg[865]), .B(n23019), .Z(n21255) );
  ANDN U22185 ( .B(n23020), .A(n23014), .Z(n23018) );
  XNOR U22186 ( .A(n23021), .B(n19591), .Z(n10732) );
  XNOR U22187 ( .A(n15903), .B(n23022), .Z(n19591) );
  AND U22188 ( .A(n17305), .B(n19583), .Z(n23021) );
  IV U22189 ( .A(n17307), .Z(n19583) );
  XNOR U22190 ( .A(n23023), .B(n17407), .Z(n17307) );
  XOR U22191 ( .A(n19075), .B(n21662), .Z(n17407) );
  XNOR U22192 ( .A(n23024), .B(n23025), .Z(n21662) );
  XOR U22193 ( .A(n17538), .B(n18203), .Z(n23025) );
  XNOR U22194 ( .A(n23026), .B(n19282), .Z(n18203) );
  ANDN U22195 ( .B(n21431), .A(n19281), .Z(n23026) );
  XNOR U22196 ( .A(n23027), .B(n22583), .Z(n17538) );
  ANDN U22197 ( .B(n22584), .A(n20753), .Z(n23027) );
  XOR U22198 ( .A(n16994), .B(n23028), .Z(n23024) );
  XOR U22199 ( .A(n17021), .B(n18110), .Z(n23028) );
  XNOR U22200 ( .A(n23029), .B(n19275), .Z(n18110) );
  NOR U22201 ( .A(n19274), .B(n20757), .Z(n23029) );
  XNOR U22202 ( .A(n23030), .B(n20984), .Z(n17021) );
  ANDN U22203 ( .B(n20985), .A(n20747), .Z(n23030) );
  XNOR U22204 ( .A(n23031), .B(n23032), .Z(n16994) );
  ANDN U22205 ( .B(n23033), .A(n20743), .Z(n23031) );
  XNOR U22206 ( .A(n23034), .B(n23035), .Z(n19075) );
  XNOR U22207 ( .A(n18364), .B(n17117), .Z(n23035) );
  XNOR U22208 ( .A(n23036), .B(n22600), .Z(n17117) );
  ANDN U22209 ( .B(n22234), .A(n22599), .Z(n23036) );
  IV U22210 ( .A(n23037), .Z(n22234) );
  XNOR U22211 ( .A(n23038), .B(n22613), .Z(n18364) );
  AND U22212 ( .A(n20684), .B(n23039), .Z(n23038) );
  XNOR U22213 ( .A(n14915), .B(n23040), .Z(n23034) );
  XNOR U22214 ( .A(n19268), .B(n18435), .Z(n23040) );
  XOR U22215 ( .A(n23041), .B(n22611), .Z(n18435) );
  ANDN U22216 ( .B(n23042), .A(n22610), .Z(n23041) );
  XNOR U22217 ( .A(n23043), .B(n22607), .Z(n19268) );
  ANDN U22218 ( .B(n20680), .A(n22606), .Z(n23043) );
  XOR U22219 ( .A(n23044), .B(n22603), .Z(n14915) );
  ANDN U22220 ( .B(n20674), .A(n22602), .Z(n23044) );
  XNOR U22221 ( .A(n20436), .B(n16896), .Z(n17305) );
  XNOR U22222 ( .A(n23045), .B(n23046), .Z(n20436) );
  AND U22223 ( .A(n21848), .B(n23047), .Z(n23045) );
  XOR U22224 ( .A(round_reg[1101]), .B(n22652), .Z(n21848) );
  XNOR U22225 ( .A(n23048), .B(n17693), .Z(n9781) );
  XOR U22226 ( .A(n22739), .B(n18323), .Z(n17693) );
  IV U22227 ( .A(n18648), .Z(n18323) );
  XNOR U22228 ( .A(n21362), .B(n19680), .Z(n18648) );
  XOR U22229 ( .A(n23049), .B(n23050), .Z(n19680) );
  XOR U22230 ( .A(n17454), .B(n21492), .Z(n23050) );
  XNOR U22231 ( .A(n23051), .B(n23052), .Z(n21492) );
  ANDN U22232 ( .B(n23053), .A(n23054), .Z(n23051) );
  XNOR U22233 ( .A(n23055), .B(n23056), .Z(n17454) );
  NOR U22234 ( .A(n22742), .B(n22743), .Z(n23055) );
  XOR U22235 ( .A(n22166), .B(n23057), .Z(n23049) );
  XOR U22236 ( .A(n18994), .B(n15630), .Z(n23057) );
  XNOR U22237 ( .A(n23058), .B(n23059), .Z(n15630) );
  AND U22238 ( .A(n22748), .B(n22746), .Z(n23058) );
  XNOR U22239 ( .A(n23060), .B(n23061), .Z(n18994) );
  NOR U22240 ( .A(n22732), .B(n22733), .Z(n23060) );
  XNOR U22241 ( .A(n23062), .B(n23063), .Z(n22166) );
  AND U22242 ( .A(n22736), .B(n23064), .Z(n23062) );
  XOR U22243 ( .A(n23065), .B(n23066), .Z(n21362) );
  XNOR U22244 ( .A(n16324), .B(n23067), .Z(n23066) );
  XNOR U22245 ( .A(n23068), .B(n23069), .Z(n16324) );
  NOR U22246 ( .A(n22709), .B(n22710), .Z(n23068) );
  XOR U22247 ( .A(n19145), .B(n23070), .Z(n23065) );
  XOR U22248 ( .A(n19253), .B(n17465), .Z(n23070) );
  XNOR U22249 ( .A(n23071), .B(n23072), .Z(n17465) );
  XNOR U22250 ( .A(n23073), .B(n23074), .Z(n19253) );
  AND U22251 ( .A(n22719), .B(n23075), .Z(n23073) );
  XNOR U22252 ( .A(n23076), .B(n23077), .Z(n19145) );
  XNOR U22253 ( .A(n23078), .B(n23054), .Z(n22739) );
  NOR U22254 ( .A(n23079), .B(n23053), .Z(n23078) );
  ANDN U22255 ( .B(n17314), .A(n17315), .Z(n23048) );
  XNOR U22256 ( .A(n23080), .B(n17154), .Z(n17315) );
  IV U22257 ( .A(n19781), .Z(n17314) );
  XOR U22258 ( .A(n21506), .B(n17218), .Z(n19781) );
  XOR U22259 ( .A(n21480), .B(n19344), .Z(n17218) );
  XOR U22260 ( .A(n23081), .B(n23082), .Z(n19344) );
  XNOR U22261 ( .A(n20165), .B(n23083), .Z(n23082) );
  XNOR U22262 ( .A(n23084), .B(n21030), .Z(n20165) );
  ANDN U22263 ( .B(n21499), .A(n21500), .Z(n23084) );
  XNOR U22264 ( .A(n17591), .B(n23085), .Z(n23081) );
  XOR U22265 ( .A(n15914), .B(n17976), .Z(n23085) );
  XOR U22266 ( .A(n23086), .B(n23087), .Z(n17976) );
  NOR U22267 ( .A(n21502), .B(n21503), .Z(n23086) );
  XNOR U22268 ( .A(n23088), .B(n21025), .Z(n15914) );
  AND U22269 ( .A(n23089), .B(n23090), .Z(n23088) );
  XNOR U22270 ( .A(n23091), .B(n23092), .Z(n17591) );
  NOR U22271 ( .A(n21512), .B(n21511), .Z(n23091) );
  XOR U22272 ( .A(n23093), .B(n23094), .Z(n21480) );
  XNOR U22273 ( .A(n17806), .B(n19896), .Z(n23094) );
  XNOR U22274 ( .A(n23095), .B(n21005), .Z(n19896) );
  ANDN U22275 ( .B(n23096), .A(n23097), .Z(n23095) );
  XNOR U22276 ( .A(n23098), .B(n20993), .Z(n17806) );
  ANDN U22277 ( .B(n23099), .A(n23100), .Z(n23098) );
  XOR U22278 ( .A(n19200), .B(n23101), .Z(n23093) );
  XOR U22279 ( .A(n17559), .B(n21433), .Z(n23101) );
  XNOR U22280 ( .A(n23102), .B(n20996), .Z(n21433) );
  ANDN U22281 ( .B(n23103), .A(n23104), .Z(n23102) );
  XOR U22282 ( .A(n23105), .B(n21002), .Z(n17559) );
  ANDN U22283 ( .B(n23106), .A(n23107), .Z(n23105) );
  XNOR U22284 ( .A(n23108), .B(n21010), .Z(n19200) );
  ANDN U22285 ( .B(n23109), .A(n23110), .Z(n23108) );
  XOR U22286 ( .A(n23111), .B(n23112), .Z(n21506) );
  NOR U22287 ( .A(n21018), .B(n23113), .Z(n23111) );
  XNOR U22288 ( .A(n23114), .B(n23115), .Z(n18414) );
  XNOR U22289 ( .A(n13907), .B(n14714), .Z(n23115) );
  XOR U22290 ( .A(n23116), .B(n14728), .Z(n14714) );
  XNOR U22291 ( .A(n21888), .B(n16539), .Z(n14728) );
  XNOR U22292 ( .A(n23117), .B(n23118), .Z(n18391) );
  XNOR U22293 ( .A(n17721), .B(n16909), .Z(n23118) );
  XOR U22294 ( .A(n23119), .B(n20952), .Z(n16909) );
  NOR U22295 ( .A(n21894), .B(n20951), .Z(n23119) );
  XNOR U22296 ( .A(round_reg[635]), .B(n22517), .Z(n20951) );
  XNOR U22297 ( .A(n23120), .B(n20956), .Z(n17721) );
  ANDN U22298 ( .B(n20955), .A(n21885), .Z(n23120) );
  XOR U22299 ( .A(round_reg[348]), .B(n23121), .Z(n20955) );
  XOR U22300 ( .A(n17471), .B(n23122), .Z(n23117) );
  XOR U22301 ( .A(n18670), .B(n20946), .Z(n23122) );
  XNOR U22302 ( .A(n23123), .B(n20963), .Z(n20946) );
  NOR U22303 ( .A(n21882), .B(n20962), .Z(n23123) );
  XNOR U22304 ( .A(round_reg[399]), .B(n21605), .Z(n20962) );
  XNOR U22305 ( .A(n23124), .B(n22378), .Z(n18670) );
  ANDN U22306 ( .B(n22379), .A(n23125), .Z(n23124) );
  XNOR U22307 ( .A(n23126), .B(n22589), .Z(n17471) );
  ANDN U22308 ( .B(n21890), .A(n21891), .Z(n23126) );
  XOR U22309 ( .A(round_reg[567]), .B(n23127), .Z(n21890) );
  XNOR U22310 ( .A(n23129), .B(n22379), .Z(n21888) );
  XOR U22311 ( .A(round_reg[469]), .B(n23130), .Z(n22379) );
  AND U22312 ( .A(n23125), .B(n23131), .Z(n23129) );
  ANDN U22313 ( .B(n14729), .A(n16513), .Z(n23116) );
  XOR U22314 ( .A(n17993), .B(n20769), .Z(n16513) );
  XOR U22315 ( .A(n23132), .B(n20500), .Z(n20769) );
  ANDN U22316 ( .B(n23133), .A(n20736), .Z(n23132) );
  XOR U22317 ( .A(round_reg[782]), .B(n23134), .Z(n20736) );
  XNOR U22318 ( .A(n23135), .B(n17506), .Z(n14729) );
  XOR U22319 ( .A(n23136), .B(n14732), .Z(n13907) );
  XOR U22320 ( .A(n23137), .B(n17948), .Z(n14732) );
  IV U22321 ( .A(n14951), .Z(n17948) );
  XNOR U22322 ( .A(n23138), .B(n23139), .Z(n20568) );
  XNOR U22323 ( .A(n19034), .B(n16602), .Z(n23139) );
  XNOR U22324 ( .A(n23140), .B(n20063), .Z(n16602) );
  XNOR U22325 ( .A(round_reg[404]), .B(n23141), .Z(n20063) );
  ANDN U22326 ( .B(n23142), .A(n22434), .Z(n23140) );
  XOR U22327 ( .A(n23143), .B(n20046), .Z(n19034) );
  XNOR U22328 ( .A(round_reg[353]), .B(n23144), .Z(n20046) );
  ANDN U22329 ( .B(n22152), .A(n22444), .Z(n23143) );
  XOR U22330 ( .A(n16906), .B(n23145), .Z(n23138) );
  XOR U22331 ( .A(n22145), .B(n21517), .Z(n23145) );
  XOR U22332 ( .A(n23146), .B(n20059), .Z(n21517) );
  XNOR U22333 ( .A(round_reg[572]), .B(n23147), .Z(n20059) );
  ANDN U22334 ( .B(n22160), .A(n22430), .Z(n23146) );
  XOR U22335 ( .A(n23148), .B(n20050), .Z(n22145) );
  XNOR U22336 ( .A(round_reg[474]), .B(n23149), .Z(n20050) );
  ANDN U22337 ( .B(n22438), .A(n22158), .Z(n23148) );
  XOR U22338 ( .A(n23150), .B(n20055), .Z(n16906) );
  XNOR U22339 ( .A(round_reg[576]), .B(n23151), .Z(n20055) );
  ANDN U22340 ( .B(n22150), .A(n22441), .Z(n23150) );
  XNOR U22341 ( .A(n23152), .B(n23153), .Z(n19249) );
  XNOR U22342 ( .A(n19988), .B(n19115), .Z(n23153) );
  XOR U22343 ( .A(n23154), .B(n21355), .Z(n19115) );
  ANDN U22344 ( .B(n23005), .A(n23155), .Z(n23154) );
  XOR U22345 ( .A(n23156), .B(n22448), .Z(n19988) );
  ANDN U22346 ( .B(n23003), .A(n23157), .Z(n23156) );
  XOR U22347 ( .A(n17902), .B(n23158), .Z(n23152) );
  XOR U22348 ( .A(n18868), .B(n19152), .Z(n23158) );
  XOR U22349 ( .A(n23159), .B(n21349), .Z(n19152) );
  NOR U22350 ( .A(n23160), .B(n23161), .Z(n23159) );
  XOR U22351 ( .A(n23162), .B(n21359), .Z(n18868) );
  NOR U22352 ( .A(n22997), .B(n23163), .Z(n23162) );
  XOR U22353 ( .A(n23164), .B(n21346), .Z(n17902) );
  ANDN U22354 ( .B(n22999), .A(n23165), .Z(n23164) );
  IV U22355 ( .A(n23166), .Z(n22999) );
  AND U22356 ( .A(n18413), .B(n14733), .Z(n23136) );
  XOR U22357 ( .A(n23167), .B(n18895), .Z(n14733) );
  IV U22358 ( .A(n18121), .Z(n18895) );
  XNOR U22359 ( .A(n23168), .B(n23169), .Z(n20310) );
  XNOR U22360 ( .A(n18682), .B(n16327), .Z(n23169) );
  XNOR U22361 ( .A(n23170), .B(n22243), .Z(n16327) );
  AND U22362 ( .A(n22244), .B(n23171), .Z(n23170) );
  XOR U22363 ( .A(n23172), .B(n22258), .Z(n18682) );
  AND U22364 ( .A(n22257), .B(n23173), .Z(n23172) );
  XOR U22365 ( .A(n15608), .B(n23174), .Z(n23168) );
  XOR U22366 ( .A(n18127), .B(n16762), .Z(n23174) );
  XNOR U22367 ( .A(n23175), .B(n22247), .Z(n16762) );
  ANDN U22368 ( .B(n22248), .A(n23176), .Z(n23175) );
  XNOR U22369 ( .A(n23177), .B(n23178), .Z(n18127) );
  ANDN U22370 ( .B(n23179), .A(n23180), .Z(n23177) );
  XNOR U22371 ( .A(n23181), .B(n22253), .Z(n15608) );
  ANDN U22372 ( .B(n22254), .A(n23182), .Z(n23181) );
  XNOR U22373 ( .A(n21439), .B(n18389), .Z(n18413) );
  XOR U22374 ( .A(n23184), .B(n23185), .Z(n21439) );
  XNOR U22375 ( .A(n12206), .B(n23188), .Z(n23114) );
  XOR U22376 ( .A(n12545), .B(n12587), .Z(n23188) );
  XOR U22377 ( .A(n23189), .B(n14736), .Z(n12587) );
  XNOR U22378 ( .A(n23190), .B(n16027), .Z(n14736) );
  IV U22379 ( .A(n16071), .Z(n16027) );
  XOR U22380 ( .A(n19026), .B(n23191), .Z(n16071) );
  XOR U22381 ( .A(n23192), .B(n23193), .Z(n19026) );
  XNOR U22382 ( .A(n20631), .B(n19492), .Z(n23193) );
  XOR U22383 ( .A(n23194), .B(n20658), .Z(n19492) );
  NOR U22384 ( .A(n23195), .B(n20657), .Z(n23194) );
  XNOR U22385 ( .A(n23196), .B(n20653), .Z(n20631) );
  ANDN U22386 ( .B(n20652), .A(n23198), .Z(n23196) );
  XNOR U22387 ( .A(n15216), .B(n23199), .Z(n23192) );
  XNOR U22388 ( .A(n15240), .B(n19600), .Z(n23199) );
  XNOR U22389 ( .A(n23200), .B(n20648), .Z(n19600) );
  XOR U22390 ( .A(round_reg[676]), .B(n23201), .Z(n20648) );
  XNOR U22391 ( .A(n23203), .B(n20661), .Z(n15240) );
  XNOR U22392 ( .A(round_reg[833]), .B(n21192), .Z(n20661) );
  ANDN U22393 ( .B(n20662), .A(n23204), .Z(n23203) );
  XNOR U22394 ( .A(n23205), .B(n20665), .Z(n15216) );
  XNOR U22395 ( .A(round_reg[904]), .B(n23206), .Z(n20665) );
  ANDN U22396 ( .B(n20666), .A(n23207), .Z(n23205) );
  ANDN U22397 ( .B(n14737), .A(n16491), .Z(n23189) );
  XNOR U22398 ( .A(n23208), .B(n17933), .Z(n16491) );
  IV U22399 ( .A(n20626), .Z(n17933) );
  XNOR U22400 ( .A(n23209), .B(n23210), .Z(n20626) );
  XOR U22401 ( .A(n16758), .B(n22391), .Z(n14737) );
  XNOR U22402 ( .A(n23211), .B(n23212), .Z(n22391) );
  ANDN U22403 ( .B(n23213), .A(n21817), .Z(n23211) );
  XNOR U22404 ( .A(n23214), .B(n14723), .Z(n12545) );
  XNOR U22405 ( .A(n19996), .B(n16682), .Z(n14723) );
  IV U22406 ( .A(n18145), .Z(n16682) );
  XOR U22407 ( .A(n23215), .B(n21737), .Z(n19996) );
  ANDN U22408 ( .B(n23216), .A(n23217), .Z(n23215) );
  AND U22409 ( .A(n14724), .B(n19556), .Z(n23214) );
  IV U22410 ( .A(n16494), .Z(n19556) );
  XOR U22411 ( .A(n23218), .B(n19023), .Z(n16494) );
  XNOR U22412 ( .A(n23219), .B(n20204), .Z(n19023) );
  XNOR U22413 ( .A(n23220), .B(n23221), .Z(n20204) );
  XOR U22414 ( .A(n23222), .B(n18422), .Z(n23221) );
  XOR U22415 ( .A(n23223), .B(n23224), .Z(n18422) );
  ANDN U22416 ( .B(n22492), .A(n23225), .Z(n23223) );
  XOR U22417 ( .A(n17324), .B(n23226), .Z(n23220) );
  XOR U22418 ( .A(n19108), .B(n15614), .Z(n23226) );
  XOR U22419 ( .A(n23227), .B(n23228), .Z(n15614) );
  ANDN U22420 ( .B(n23229), .A(n22496), .Z(n23227) );
  XOR U22421 ( .A(n23230), .B(n23231), .Z(n19108) );
  ANDN U22422 ( .B(n23232), .A(n22483), .Z(n23230) );
  XNOR U22423 ( .A(n23233), .B(n23234), .Z(n17324) );
  XNOR U22424 ( .A(n17491), .B(n20123), .Z(n14724) );
  XNOR U22425 ( .A(n23236), .B(n18781), .Z(n20123) );
  NOR U22426 ( .A(n23237), .B(n20376), .Z(n23236) );
  XOR U22427 ( .A(n21598), .B(n22381), .Z(n17491) );
  XOR U22428 ( .A(n23238), .B(n23239), .Z(n22381) );
  XOR U22429 ( .A(n20139), .B(n18273), .Z(n23239) );
  XOR U22430 ( .A(n23240), .B(n20159), .Z(n18273) );
  XNOR U22431 ( .A(round_reg[1071]), .B(n23241), .Z(n20159) );
  ANDN U22432 ( .B(n22325), .A(n20158), .Z(n23240) );
  XNOR U22433 ( .A(round_reg[703]), .B(n22783), .Z(n20158) );
  XOR U22434 ( .A(round_reg[637]), .B(n23242), .Z(n22325) );
  XNOR U22435 ( .A(n23243), .B(n20163), .Z(n20139) );
  XOR U22436 ( .A(round_reg[1120]), .B(n23244), .Z(n20163) );
  ANDN U22437 ( .B(n22384), .A(n20162), .Z(n23243) );
  XNOR U22438 ( .A(round_reg[717]), .B(n23245), .Z(n20162) );
  XNOR U22439 ( .A(round_reg[350]), .B(n23246), .Z(n22384) );
  XOR U22440 ( .A(n17519), .B(n23247), .Z(n23238) );
  XOR U22441 ( .A(n18732), .B(n17590), .Z(n23247) );
  XNOR U22442 ( .A(n23248), .B(n20146), .Z(n17590) );
  XNOR U22443 ( .A(round_reg[1210]), .B(n23249), .Z(n20146) );
  ANDN U22444 ( .B(n22333), .A(n20145), .Z(n23248) );
  XNOR U22445 ( .A(round_reg[827]), .B(n23250), .Z(n20145) );
  XNOR U22446 ( .A(round_reg[401]), .B(n21199), .Z(n22333) );
  XNOR U22447 ( .A(n23251), .B(n20155), .Z(n18732) );
  XOR U22448 ( .A(round_reg[1218]), .B(n23252), .Z(n20155) );
  ANDN U22449 ( .B(n22331), .A(n20154), .Z(n23251) );
  XNOR U22450 ( .A(round_reg[860]), .B(n23253), .Z(n20154) );
  XNOR U22451 ( .A(round_reg[471]), .B(n23254), .Z(n22331) );
  XNOR U22452 ( .A(n23255), .B(n20149), .Z(n17519) );
  XOR U22453 ( .A(round_reg[978]), .B(n21186), .Z(n20149) );
  AND U22454 ( .A(n20150), .B(n22329), .Z(n23255) );
  XNOR U22455 ( .A(round_reg[569]), .B(n22831), .Z(n22329) );
  XOR U22456 ( .A(round_reg[931]), .B(n23256), .Z(n20150) );
  XOR U22457 ( .A(n23257), .B(n23258), .Z(n21598) );
  XNOR U22458 ( .A(n17623), .B(n18532), .Z(n23258) );
  XNOR U22459 ( .A(n23259), .B(n18842), .Z(n18532) );
  XOR U22460 ( .A(round_reg[25]), .B(n21198), .Z(n18842) );
  ANDN U22461 ( .B(n18843), .A(n20120), .Z(n23259) );
  XOR U22462 ( .A(round_reg[1575]), .B(n23260), .Z(n18843) );
  XNOR U22463 ( .A(n23261), .B(n18777), .Z(n17623) );
  XOR U22464 ( .A(round_reg[111]), .B(n23262), .Z(n18777) );
  ANDN U22465 ( .B(n23263), .A(n18776), .Z(n23261) );
  XNOR U22466 ( .A(round_reg[1292]), .B(n22368), .Z(n18776) );
  XOR U22467 ( .A(n17325), .B(n23264), .Z(n23257) );
  XOR U22468 ( .A(n17450), .B(n16066), .Z(n23264) );
  XNOR U22469 ( .A(n23265), .B(n20372), .Z(n16066) );
  XOR U22470 ( .A(round_reg[277]), .B(n23266), .Z(n20372) );
  ANDN U22471 ( .B(n20128), .A(n20129), .Z(n23265) );
  XOR U22472 ( .A(round_reg[1510]), .B(n23267), .Z(n20128) );
  XNOR U22473 ( .A(n23268), .B(n18780), .Z(n17450) );
  XOR U22474 ( .A(round_reg[229]), .B(n22769), .Z(n18780) );
  AND U22475 ( .A(n23237), .B(n18781), .Z(n23268) );
  XOR U22476 ( .A(round_reg[1449]), .B(n22372), .Z(n18781) );
  XNOR U22477 ( .A(n23269), .B(n19676), .Z(n17325) );
  XOR U22478 ( .A(round_reg[170]), .B(n22274), .Z(n19676) );
  AND U22479 ( .A(n19677), .B(n20118), .Z(n23269) );
  XOR U22480 ( .A(round_reg[1355]), .B(n23270), .Z(n19677) );
  XOR U22481 ( .A(n23271), .B(n14719), .Z(n12206) );
  XNOR U22482 ( .A(n19277), .B(n17434), .Z(n14719) );
  XNOR U22483 ( .A(n19616), .B(n22939), .Z(n17434) );
  XNOR U22484 ( .A(n23272), .B(n23273), .Z(n22939) );
  XNOR U22485 ( .A(n17329), .B(n22785), .Z(n23273) );
  XNOR U22486 ( .A(n23274), .B(n21416), .Z(n22785) );
  XOR U22487 ( .A(round_reg[1048]), .B(n23275), .Z(n21416) );
  ANDN U22488 ( .B(n22791), .A(n21674), .Z(n23274) );
  XNOR U22489 ( .A(n23276), .B(n21429), .Z(n17329) );
  XOR U22490 ( .A(round_reg[1019]), .B(n22986), .Z(n21429) );
  ANDN U22491 ( .B(n22804), .A(n23277), .Z(n23276) );
  XOR U22492 ( .A(n18194), .B(n23278), .Z(n23272) );
  XOR U22493 ( .A(n18227), .B(n22677), .Z(n23278) );
  XNOR U22494 ( .A(n23279), .B(n21412), .Z(n22677) );
  XOR U22495 ( .A(round_reg[1187]), .B(n23280), .Z(n21412) );
  ANDN U22496 ( .B(n22801), .A(n21672), .Z(n23279) );
  XNOR U22497 ( .A(n23281), .B(n21425), .Z(n18227) );
  XOR U22498 ( .A(round_reg[1259]), .B(n22375), .Z(n21425) );
  XNOR U22499 ( .A(n23282), .B(n21421), .Z(n18194) );
  XOR U22500 ( .A(round_reg[1097]), .B(n23283), .Z(n21421) );
  ANDN U22501 ( .B(n22793), .A(n21668), .Z(n23282) );
  XOR U22502 ( .A(n23284), .B(n23285), .Z(n19616) );
  XNOR U22503 ( .A(n19401), .B(n18148), .Z(n23285) );
  XNOR U22504 ( .A(n23286), .B(n20745), .Z(n18148) );
  IV U22505 ( .A(n23287), .Z(n20745) );
  NOR U22506 ( .A(n23032), .B(n20744), .Z(n23286) );
  XNOR U22507 ( .A(n23288), .B(n21432), .Z(n19401) );
  AND U22508 ( .A(n19282), .B(n19280), .Z(n23288) );
  XOR U22509 ( .A(round_reg[1396]), .B(n23289), .Z(n19280) );
  XNOR U22510 ( .A(round_reg[1020]), .B(n21772), .Z(n19282) );
  IV U22511 ( .A(n23290), .Z(n21772) );
  XOR U22512 ( .A(n20738), .B(n23291), .Z(n23284) );
  XOR U22513 ( .A(n17960), .B(n19147), .Z(n23291) );
  XNOR U22514 ( .A(n23292), .B(n20755), .Z(n19147) );
  NOR U22515 ( .A(n22583), .B(n20754), .Z(n23292) );
  XNOR U22516 ( .A(round_reg[1552]), .B(n22265), .Z(n20754) );
  XOR U22517 ( .A(round_reg[1188]), .B(n23293), .Z(n22583) );
  XNOR U22518 ( .A(n23294), .B(n20748), .Z(n17960) );
  AND U22519 ( .A(n20984), .B(n20983), .Z(n23294) );
  XOR U22520 ( .A(round_reg[1426]), .B(n23295), .Z(n20983) );
  XNOR U22521 ( .A(round_reg[1049]), .B(n21760), .Z(n20984) );
  XNOR U22522 ( .A(n23296), .B(n20758), .Z(n20738) );
  AND U22523 ( .A(n19273), .B(n19275), .Z(n23296) );
  XNOR U22524 ( .A(round_reg[1098]), .B(n22108), .Z(n19275) );
  XNOR U22525 ( .A(round_reg[1487]), .B(n23297), .Z(n19273) );
  XOR U22526 ( .A(n23298), .B(n20744), .Z(n19277) );
  AND U22527 ( .A(n23032), .B(n23299), .Z(n23298) );
  XOR U22528 ( .A(round_reg[1260]), .B(n23300), .Z(n23032) );
  XOR U22529 ( .A(n22089), .B(n16788), .Z(n16486) );
  XOR U22530 ( .A(n20765), .B(n21824), .Z(n16788) );
  XOR U22531 ( .A(n23301), .B(n23302), .Z(n21824) );
  XNOR U22532 ( .A(n15859), .B(n17579), .Z(n23302) );
  XNOR U22533 ( .A(n23303), .B(n22419), .Z(n17579) );
  AND U22534 ( .A(n22097), .B(n23304), .Z(n23303) );
  XOR U22535 ( .A(n23305), .B(n22423), .Z(n15859) );
  IV U22536 ( .A(n23306), .Z(n22423) );
  ANDN U22537 ( .B(n23307), .A(n23308), .Z(n23305) );
  XOR U22538 ( .A(n17573), .B(n23309), .Z(n23301) );
  XOR U22539 ( .A(n23310), .B(n15832), .Z(n23309) );
  XOR U22540 ( .A(n23311), .B(n23312), .Z(n15832) );
  NOR U22541 ( .A(n22082), .B(n22081), .Z(n23311) );
  XOR U22542 ( .A(n23313), .B(n22408), .Z(n17573) );
  IV U22543 ( .A(n23314), .Z(n22408) );
  ANDN U22544 ( .B(n22091), .A(n22092), .Z(n23313) );
  XOR U22545 ( .A(n23315), .B(n23316), .Z(n20765) );
  XNOR U22546 ( .A(n18711), .B(n18906), .Z(n23316) );
  XOR U22547 ( .A(n23317), .B(n22222), .Z(n18906) );
  NOR U22548 ( .A(n19921), .B(n19847), .Z(n23317) );
  XOR U22549 ( .A(round_reg[1594]), .B(n23318), .Z(n19847) );
  XOR U22550 ( .A(n23319), .B(n22231), .Z(n18711) );
  ANDN U22551 ( .B(n23320), .A(n19860), .Z(n23319) );
  XOR U22552 ( .A(round_reg[1529]), .B(n22831), .Z(n19860) );
  XOR U22553 ( .A(n15332), .B(n23321), .Z(n23315) );
  XOR U22554 ( .A(n17723), .B(n18337), .Z(n23321) );
  XNOR U22555 ( .A(n23322), .B(n22228), .Z(n18337) );
  ANDN U22556 ( .B(n19923), .A(n19856), .Z(n23322) );
  XOR U22557 ( .A(round_reg[1468]), .B(n23323), .Z(n19856) );
  XNOR U22558 ( .A(n23324), .B(n22226), .Z(n17723) );
  ANDN U22559 ( .B(n19918), .A(n19852), .Z(n23324) );
  XOR U22560 ( .A(round_reg[1311]), .B(n23325), .Z(n19852) );
  XOR U22561 ( .A(n23326), .B(n22219), .Z(n15332) );
  ANDN U22562 ( .B(n19843), .A(n19925), .Z(n23326) );
  XOR U22563 ( .A(round_reg[1374]), .B(n22959), .Z(n19843) );
  IV U22564 ( .A(n23327), .Z(n22959) );
  XNOR U22565 ( .A(n23328), .B(n23308), .Z(n22089) );
  ANDN U22566 ( .B(n22421), .A(n23307), .Z(n23328) );
  XNOR U22567 ( .A(n23329), .B(n16746), .Z(n14720) );
  XOR U22568 ( .A(n23332), .B(n6614), .Z(n2558) );
  IV U22569 ( .A(n9263), .Z(n6614) );
  XNOR U22570 ( .A(n19410), .B(n9529), .Z(n9263) );
  XNOR U22571 ( .A(n16499), .B(n17157), .Z(n9529) );
  XNOR U22572 ( .A(n23333), .B(n23334), .Z(n17157) );
  XNOR U22573 ( .A(n12475), .B(n13657), .Z(n23334) );
  XOR U22574 ( .A(n23335), .B(n16626), .Z(n13657) );
  XNOR U22575 ( .A(n19187), .B(n23336), .Z(n16626) );
  XOR U22576 ( .A(n20193), .B(n19537), .Z(n19187) );
  XOR U22577 ( .A(n23337), .B(n23338), .Z(n19537) );
  XNOR U22578 ( .A(n23339), .B(n18218), .Z(n23338) );
  XNOR U22579 ( .A(n23340), .B(n22747), .Z(n18218) );
  ANDN U22580 ( .B(n23341), .A(n23059), .Z(n23340) );
  XOR U22581 ( .A(n19601), .B(n23342), .Z(n23337) );
  XOR U22582 ( .A(n19250), .B(n18541), .Z(n23342) );
  XNOR U22583 ( .A(n23343), .B(n22734), .Z(n18541) );
  ANDN U22584 ( .B(n23344), .A(n23061), .Z(n23343) );
  XOR U22585 ( .A(n23345), .B(n22744), .Z(n19250) );
  AND U22586 ( .A(n23056), .B(n23346), .Z(n23345) );
  XNOR U22587 ( .A(n23347), .B(n23079), .Z(n19601) );
  ANDN U22588 ( .B(n23348), .A(n23052), .Z(n23347) );
  XOR U22589 ( .A(n23349), .B(n23350), .Z(n20193) );
  XNOR U22590 ( .A(n17232), .B(n19190), .Z(n23350) );
  XNOR U22591 ( .A(n23351), .B(n22720), .Z(n19190) );
  ANDN U22592 ( .B(n23352), .A(n23074), .Z(n23351) );
  XNOR U22593 ( .A(n23353), .B(n22715), .Z(n17232) );
  ANDN U22594 ( .B(n23354), .A(n23355), .Z(n23353) );
  XOR U22595 ( .A(n17444), .B(n23356), .Z(n23349) );
  XOR U22596 ( .A(n21749), .B(n15651), .Z(n23356) );
  XNOR U22597 ( .A(n23357), .B(n22711), .Z(n15651) );
  ANDN U22598 ( .B(n23358), .A(n23069), .Z(n23357) );
  XNOR U22599 ( .A(n23359), .B(n22728), .Z(n21749) );
  ANDN U22600 ( .B(n23360), .A(n23072), .Z(n23359) );
  XNOR U22601 ( .A(n23361), .B(n22724), .Z(n17444) );
  ANDN U22602 ( .B(n23362), .A(n23077), .Z(n23361) );
  AND U22603 ( .A(n16627), .B(n15113), .Z(n23335) );
  XNOR U22604 ( .A(n23363), .B(n16638), .Z(n12475) );
  XNOR U22605 ( .A(n18156), .B(n23364), .Z(n16638) );
  XOR U22606 ( .A(n23365), .B(n19084), .Z(n18156) );
  XNOR U22607 ( .A(n23366), .B(n23367), .Z(n19084) );
  XNOR U22608 ( .A(n19106), .B(n18960), .Z(n23367) );
  XNOR U22609 ( .A(n23368), .B(n23369), .Z(n18960) );
  AND U22610 ( .A(n23370), .B(n22674), .Z(n23368) );
  XNOR U22611 ( .A(n23371), .B(n23372), .Z(n19106) );
  AND U22612 ( .A(n23373), .B(n22666), .Z(n23371) );
  XOR U22613 ( .A(n18717), .B(n23374), .Z(n23366) );
  XOR U22614 ( .A(n23375), .B(n20732), .Z(n23374) );
  XNOR U22615 ( .A(n23376), .B(n23377), .Z(n20732) );
  ANDN U22616 ( .B(n23378), .A(n22657), .Z(n23376) );
  XNOR U22617 ( .A(n23379), .B(n23380), .Z(n18717) );
  ANDN U22618 ( .B(n23381), .A(n22670), .Z(n23379) );
  AND U22619 ( .A(n15099), .B(n16637), .Z(n23363) );
  XNOR U22620 ( .A(n18464), .B(n23001), .Z(n16637) );
  XNOR U22621 ( .A(n23382), .B(n23161), .Z(n23001) );
  ANDN U22622 ( .B(n21350), .A(n21348), .Z(n23382) );
  XNOR U22623 ( .A(n23383), .B(n23384), .Z(n19864) );
  XNOR U22624 ( .A(n20567), .B(n17675), .Z(n23384) );
  XOR U22625 ( .A(n23385), .B(n23142), .Z(n17675) );
  IV U22626 ( .A(n22155), .Z(n23142) );
  XNOR U22627 ( .A(round_reg[27]), .B(n23386), .Z(n22155) );
  ANDN U22628 ( .B(n22434), .A(n20062), .Z(n23385) );
  XOR U22629 ( .A(round_reg[1213]), .B(n23387), .Z(n20062) );
  XOR U22630 ( .A(round_reg[1577]), .B(n22760), .Z(n22434) );
  XOR U22631 ( .A(n23388), .B(n22150), .Z(n20567) );
  XOR U22632 ( .A(round_reg[231]), .B(n22361), .Z(n22150) );
  ANDN U22633 ( .B(n22441), .A(n20054), .Z(n23388) );
  XOR U22634 ( .A(round_reg[1074]), .B(n23197), .Z(n20054) );
  XOR U22635 ( .A(round_reg[1451]), .B(n23389), .Z(n22441) );
  XNOR U22636 ( .A(n18316), .B(n23390), .Z(n23383) );
  XOR U22637 ( .A(n19220), .B(n17221), .Z(n23390) );
  XOR U22638 ( .A(n23391), .B(n22160), .Z(n17221) );
  XNOR U22639 ( .A(round_reg[172]), .B(n23392), .Z(n22160) );
  AND U22640 ( .A(n22430), .B(n20058), .Z(n23391) );
  IV U22641 ( .A(n22431), .Z(n20058) );
  XOR U22642 ( .A(round_reg[981]), .B(n23393), .Z(n22431) );
  XOR U22643 ( .A(round_reg[1357]), .B(n23245), .Z(n22430) );
  XOR U22644 ( .A(n23394), .B(n22152), .Z(n19220) );
  XNOR U22645 ( .A(round_reg[279]), .B(n23395), .Z(n22152) );
  AND U22646 ( .A(n22444), .B(n20045), .Z(n23394) );
  XNOR U22647 ( .A(round_reg[1123]), .B(n23396), .Z(n20045) );
  XOR U22648 ( .A(round_reg[1512]), .B(n23397), .Z(n22444) );
  XNOR U22649 ( .A(n23398), .B(n22158), .Z(n18316) );
  XOR U22650 ( .A(round_reg[113]), .B(n23399), .Z(n22158) );
  ANDN U22651 ( .B(n20049), .A(n22438), .Z(n23398) );
  XNOR U22652 ( .A(round_reg[1294]), .B(n22115), .Z(n22438) );
  XNOR U22653 ( .A(round_reg[1221]), .B(n23400), .Z(n20049) );
  XNOR U22654 ( .A(n23401), .B(n23402), .Z(n19322) );
  XOR U22655 ( .A(n17947), .B(n17598), .Z(n23402) );
  XOR U22656 ( .A(n23403), .B(n23155), .Z(n17598) );
  ANDN U22657 ( .B(n21354), .A(n23005), .Z(n23403) );
  XNOR U22658 ( .A(round_reg[577]), .B(n22834), .Z(n23005) );
  XNOR U22659 ( .A(round_reg[232]), .B(n23397), .Z(n21354) );
  XNOR U22660 ( .A(n23404), .B(n23157), .Z(n17947) );
  XNOR U22661 ( .A(round_reg[354]), .B(n23405), .Z(n23003) );
  XNOR U22662 ( .A(round_reg[280]), .B(n23406), .Z(n22447) );
  XNOR U22663 ( .A(n14950), .B(n23407), .Z(n23401) );
  XOR U22664 ( .A(n23137), .B(n18275), .Z(n23407) );
  XNOR U22665 ( .A(n23408), .B(n23160), .Z(n18275) );
  AND U22666 ( .A(n21348), .B(n23161), .Z(n23408) );
  XOR U22667 ( .A(round_reg[405]), .B(n23409), .Z(n23161) );
  XNOR U22668 ( .A(round_reg[28]), .B(n23121), .Z(n21348) );
  XNOR U22669 ( .A(n23410), .B(n23163), .Z(n23137) );
  AND U22670 ( .A(n21358), .B(n22997), .Z(n23410) );
  XOR U22671 ( .A(round_reg[475]), .B(n23411), .Z(n22997) );
  XNOR U22672 ( .A(round_reg[114]), .B(n23197), .Z(n21358) );
  XNOR U22673 ( .A(n23412), .B(n23165), .Z(n14950) );
  AND U22674 ( .A(n21344), .B(n23166), .Z(n23412) );
  XOR U22675 ( .A(round_reg[573]), .B(n23387), .Z(n23166) );
  XNOR U22676 ( .A(round_reg[173]), .B(n23413), .Z(n21344) );
  XNOR U22677 ( .A(n23414), .B(n17154), .Z(n15099) );
  XNOR U22678 ( .A(n23415), .B(n23416), .Z(n20194) );
  XOR U22679 ( .A(n19053), .B(n15596), .Z(n23416) );
  XOR U22680 ( .A(n23417), .B(n20721), .Z(n15596) );
  XOR U22681 ( .A(round_reg[413]), .B(n23418), .Z(n20721) );
  ANDN U22682 ( .B(n21767), .A(n21716), .Z(n23417) );
  XOR U22683 ( .A(n23419), .B(n20731), .Z(n19053) );
  XOR U22684 ( .A(round_reg[362]), .B(n23420), .Z(n20731) );
  ANDN U22685 ( .B(n21761), .A(n21723), .Z(n23419) );
  XOR U22686 ( .A(n16918), .B(n23421), .Z(n23415) );
  XOR U22687 ( .A(n19624), .B(n16945), .Z(n23421) );
  XNOR U22688 ( .A(n23422), .B(n20727), .Z(n16945) );
  XOR U22689 ( .A(round_reg[585]), .B(n21185), .Z(n20727) );
  ANDN U22690 ( .B(n21755), .A(n21720), .Z(n23422) );
  XNOR U22691 ( .A(n23423), .B(n21745), .Z(n19624) );
  XOR U22692 ( .A(round_reg[483]), .B(n23396), .Z(n21745) );
  ANDN U22693 ( .B(n21757), .A(n23424), .Z(n23423) );
  XNOR U22694 ( .A(n23425), .B(n20717), .Z(n16918) );
  XOR U22695 ( .A(round_reg[517]), .B(n23426), .Z(n20717) );
  ANDN U22696 ( .B(n21764), .A(n21713), .Z(n23425) );
  XNOR U22697 ( .A(n23427), .B(n23428), .Z(n19957) );
  XNOR U22698 ( .A(n18313), .B(n17894), .Z(n23428) );
  XNOR U22699 ( .A(n23429), .B(n23430), .Z(n17894) );
  AND U22700 ( .A(n23431), .B(n21739), .Z(n23429) );
  XNOR U22701 ( .A(n23432), .B(n20006), .Z(n18313) );
  ANDN U22702 ( .B(n21732), .A(n20005), .Z(n23432) );
  XOR U22703 ( .A(n19993), .B(n23433), .Z(n23427) );
  XNOR U22704 ( .A(n18826), .B(n15243), .Z(n23433) );
  XNOR U22705 ( .A(n23434), .B(n23216), .Z(n15243) );
  AND U22706 ( .A(n23217), .B(n21735), .Z(n23434) );
  IV U22707 ( .A(n23435), .Z(n21735) );
  XNOR U22708 ( .A(n23436), .B(n20010), .Z(n18826) );
  NOR U22709 ( .A(n20009), .B(n21728), .Z(n23436) );
  XNOR U22710 ( .A(n23437), .B(n19999), .Z(n19993) );
  ANDN U22711 ( .B(n20000), .A(n23438), .Z(n23437) );
  XNOR U22712 ( .A(n13699), .B(n23439), .Z(n23333) );
  XOR U22713 ( .A(n11256), .B(n16598), .Z(n23439) );
  XOR U22714 ( .A(n23440), .B(n16634), .Z(n16598) );
  XNOR U22715 ( .A(n20260), .B(n16057), .Z(n16634) );
  IV U22716 ( .A(n16001), .Z(n16057) );
  XOR U22717 ( .A(n23441), .B(n21791), .Z(n16001) );
  XNOR U22718 ( .A(n23442), .B(n23443), .Z(n21791) );
  XOR U22719 ( .A(n17684), .B(n18278), .Z(n23443) );
  XOR U22720 ( .A(n23444), .B(n21396), .Z(n18278) );
  AND U22721 ( .A(n20252), .B(n20254), .Z(n23444) );
  XOR U22722 ( .A(round_reg[1008]), .B(n23445), .Z(n20252) );
  XNOR U22723 ( .A(n23446), .B(n21404), .Z(n17684) );
  ANDN U22724 ( .B(n20256), .A(n20257), .Z(n23446) );
  XNOR U22725 ( .A(round_reg[1176]), .B(n23447), .Z(n20256) );
  XOR U22726 ( .A(n21364), .B(n23448), .Z(n23442) );
  XOR U22727 ( .A(n18901), .B(n19318), .Z(n23448) );
  XNOR U22728 ( .A(n23449), .B(n23450), .Z(n19318) );
  AND U22729 ( .A(n20262), .B(n20264), .Z(n23449) );
  XNOR U22730 ( .A(n23451), .B(n21392), .Z(n18901) );
  AND U22731 ( .A(n21393), .B(n23452), .Z(n23451) );
  XNOR U22732 ( .A(n23453), .B(n21401), .Z(n21364) );
  ANDN U22733 ( .B(n20266), .A(n20267), .Z(n23453) );
  XOR U22734 ( .A(round_reg[1150]), .B(n22435), .Z(n20266) );
  XNOR U22735 ( .A(n23454), .B(n21393), .Z(n20260) );
  XOR U22736 ( .A(round_reg[1037]), .B(n23245), .Z(n21393) );
  ANDN U22737 ( .B(n23455), .A(n23456), .Z(n23454) );
  AND U22738 ( .A(n19416), .B(n19415), .Z(n23440) );
  XOR U22739 ( .A(n23457), .B(n16039), .Z(n19415) );
  XNOR U22740 ( .A(n23459), .B(n23460), .Z(n20940) );
  XNOR U22741 ( .A(n18451), .B(n16550), .Z(n23460) );
  XNOR U22742 ( .A(n23461), .B(n19522), .Z(n16550) );
  XOR U22743 ( .A(round_reg[504]), .B(n22642), .Z(n19522) );
  AND U22744 ( .A(n19523), .B(n23462), .Z(n23461) );
  XOR U22745 ( .A(round_reg[79]), .B(n21605), .Z(n19523) );
  XNOR U22746 ( .A(n23463), .B(n19518), .Z(n18451) );
  XOR U22747 ( .A(round_reg[606]), .B(n23464), .Z(n19518) );
  ANDN U22748 ( .B(n19519), .A(n21944), .Z(n23463) );
  XOR U22749 ( .A(round_reg[197]), .B(n23426), .Z(n19519) );
  XOR U22750 ( .A(n17844), .B(n23465), .Z(n23459) );
  XNOR U22751 ( .A(n17416), .B(n15133), .Z(n23465) );
  XNOR U22752 ( .A(n23466), .B(n19513), .Z(n15133) );
  XNOR U22753 ( .A(round_reg[383]), .B(n22783), .Z(n19513) );
  AND U22754 ( .A(n21936), .B(n19514), .Z(n23466) );
  XOR U22755 ( .A(round_reg[309]), .B(n23467), .Z(n19514) );
  XNOR U22756 ( .A(n23468), .B(n19509), .Z(n17416) );
  XOR U22757 ( .A(round_reg[434]), .B(n23197), .Z(n19509) );
  XOR U22758 ( .A(round_reg[57]), .B(n23469), .Z(n19510) );
  XNOR U22759 ( .A(n23470), .B(n19526), .Z(n17844) );
  XOR U22760 ( .A(round_reg[538]), .B(n23471), .Z(n19526) );
  AND U22761 ( .A(n19527), .B(n23472), .Z(n23470) );
  XOR U22762 ( .A(round_reg[138]), .B(n22108), .Z(n19527) );
  XOR U22763 ( .A(n17174), .B(n21670), .Z(n19416) );
  XNOR U22764 ( .A(n23473), .B(n23277), .Z(n21670) );
  ANDN U22765 ( .B(n23474), .A(n21428), .Z(n23473) );
  XOR U22766 ( .A(round_reg[1395]), .B(n23475), .Z(n21428) );
  IV U22767 ( .A(n17557), .Z(n17174) );
  XOR U22768 ( .A(n22354), .B(n18205), .Z(n17557) );
  XNOR U22769 ( .A(n23476), .B(n23477), .Z(n18205) );
  XNOR U22770 ( .A(n16013), .B(n17862), .Z(n23477) );
  XOR U22771 ( .A(n23478), .B(n22804), .Z(n17862) );
  XNOR U22772 ( .A(round_reg[908]), .B(n23479), .Z(n22804) );
  AND U22773 ( .A(n23277), .B(n21427), .Z(n23478) );
  IV U22774 ( .A(n23474), .Z(n21427) );
  XOR U22775 ( .A(round_reg[146]), .B(n23295), .Z(n23474) );
  XOR U22776 ( .A(round_reg[546]), .B(n23480), .Z(n23277) );
  XOR U22777 ( .A(n23481), .B(n22801), .Z(n16013) );
  ANDN U22778 ( .B(n21672), .A(n21410), .Z(n23481) );
  XNOR U22779 ( .A(round_reg[1]), .B(n22966), .Z(n21410) );
  XOR U22780 ( .A(round_reg[442]), .B(n22991), .Z(n21672) );
  XNOR U22781 ( .A(n22938), .B(n23483), .Z(n23476) );
  XNOR U22782 ( .A(n16678), .B(n19684), .Z(n23483) );
  XOR U22783 ( .A(n23484), .B(n22797), .Z(n19684) );
  XOR U22784 ( .A(round_reg[837]), .B(n23485), .Z(n22797) );
  ANDN U22785 ( .B(n21666), .A(n21423), .Z(n23484) );
  XOR U22786 ( .A(round_reg[87]), .B(n23486), .Z(n21423) );
  XOR U22787 ( .A(round_reg[448]), .B(n23011), .Z(n21666) );
  XOR U22788 ( .A(n23487), .B(n22791), .Z(n16678) );
  XNOR U22789 ( .A(round_reg[680]), .B(n23488), .Z(n22791) );
  ANDN U22790 ( .B(n21674), .A(n21414), .Z(n23487) );
  XNOR U22791 ( .A(round_reg[205]), .B(n23489), .Z(n21414) );
  XNOR U22792 ( .A(round_reg[614]), .B(n22432), .Z(n21674) );
  XOR U22793 ( .A(n23490), .B(n22793), .Z(n22938) );
  XNOR U22794 ( .A(round_reg[758]), .B(n23491), .Z(n22793) );
  ANDN U22795 ( .B(n21668), .A(n21419), .Z(n23490) );
  XNOR U22796 ( .A(round_reg[317]), .B(n23242), .Z(n21419) );
  XOR U22797 ( .A(round_reg[327]), .B(n23492), .Z(n21668) );
  XOR U22798 ( .A(n23493), .B(n23494), .Z(n22354) );
  XNOR U22799 ( .A(n16551), .B(n16926), .Z(n23494) );
  XNOR U22800 ( .A(n23495), .B(n22950), .Z(n16926) );
  AND U22801 ( .A(n22926), .B(n23496), .Z(n23495) );
  XNOR U22802 ( .A(round_reg[1550]), .B(n23497), .Z(n22926) );
  XOR U22803 ( .A(n23498), .B(n23499), .Z(n16551) );
  XNOR U22804 ( .A(n17066), .B(n23500), .Z(n23493) );
  XNOR U22805 ( .A(n18899), .B(n18970), .Z(n23500) );
  XOR U22806 ( .A(n23501), .B(n22953), .Z(n18970) );
  AND U22807 ( .A(n22923), .B(n22921), .Z(n23501) );
  XOR U22808 ( .A(round_reg[1485]), .B(n23502), .Z(n22921) );
  XNOR U22809 ( .A(n23503), .B(n22945), .Z(n18899) );
  ANDN U22810 ( .B(n22930), .A(n22931), .Z(n23503) );
  XOR U22811 ( .A(round_reg[1331]), .B(n23504), .Z(n22930) );
  XOR U22812 ( .A(n23505), .B(n23506), .Z(n17066) );
  AND U22813 ( .A(n22934), .B(n23507), .Z(n23505) );
  XNOR U22814 ( .A(n23508), .B(n16631), .Z(n11256) );
  XNOR U22815 ( .A(n18601), .B(n23509), .Z(n16631) );
  IV U22816 ( .A(n16706), .Z(n18601) );
  XNOR U22817 ( .A(n21141), .B(n17483), .Z(n16630) );
  XNOR U22818 ( .A(n23510), .B(n23511), .Z(n20135) );
  XNOR U22819 ( .A(n23512), .B(n15330), .Z(n23511) );
  XOR U22820 ( .A(n23513), .B(n23514), .Z(n15330) );
  XOR U22821 ( .A(n18297), .B(n23515), .Z(n23510) );
  XOR U22822 ( .A(n17171), .B(n17726), .Z(n23515) );
  XNOR U22823 ( .A(n23516), .B(n23517), .Z(n17726) );
  XNOR U22824 ( .A(n23518), .B(n23519), .Z(n17171) );
  AND U22825 ( .A(n21172), .B(n23520), .Z(n23518) );
  XOR U22826 ( .A(n23521), .B(n23522), .Z(n18297) );
  ANDN U22827 ( .B(n23523), .A(n21174), .Z(n23521) );
  XOR U22828 ( .A(n23524), .B(n23525), .Z(n18453) );
  XNOR U22829 ( .A(n18097), .B(n18932), .Z(n23525) );
  XOR U22830 ( .A(n23526), .B(n21656), .Z(n18932) );
  NOR U22831 ( .A(n21156), .B(n21155), .Z(n23526) );
  XOR U22832 ( .A(round_reg[1477]), .B(n23485), .Z(n21155) );
  XOR U22833 ( .A(n23527), .B(n20806), .Z(n18097) );
  ANDN U22834 ( .B(n21144), .A(n20805), .Z(n23527) );
  XNOR U22835 ( .A(round_reg[1386]), .B(n23528), .Z(n20805) );
  XOR U22836 ( .A(n20795), .B(n23529), .Z(n23524) );
  XOR U22837 ( .A(n17890), .B(n16040), .Z(n23529) );
  XNOR U22838 ( .A(n23530), .B(n23531), .Z(n16040) );
  XOR U22839 ( .A(n23532), .B(n23533), .Z(n17890) );
  NOR U22840 ( .A(n21152), .B(n21151), .Z(n23532) );
  XOR U22841 ( .A(round_reg[1416]), .B(n23534), .Z(n21151) );
  XNOR U22842 ( .A(n23535), .B(n20879), .Z(n20795) );
  XOR U22843 ( .A(n23537), .B(n20880), .Z(n21141) );
  XOR U22844 ( .A(round_reg[1542]), .B(n23538), .Z(n20880) );
  NOR U22845 ( .A(n23536), .B(n23539), .Z(n23537) );
  IV U22846 ( .A(n19409), .Z(n15103) );
  XOR U22847 ( .A(n23540), .B(n16557), .Z(n19409) );
  IV U22848 ( .A(n17388), .Z(n16557) );
  XOR U22849 ( .A(n23541), .B(n23542), .Z(n22629) );
  XNOR U22850 ( .A(n18799), .B(n18905), .Z(n23542) );
  XOR U22851 ( .A(n23543), .B(n23544), .Z(n18905) );
  NOR U22852 ( .A(n23545), .B(n23546), .Z(n23543) );
  XOR U22853 ( .A(n23547), .B(n21642), .Z(n18799) );
  ANDN U22854 ( .B(n21643), .A(n23548), .Z(n23547) );
  XNOR U22855 ( .A(n17191), .B(n23549), .Z(n23541) );
  XOR U22856 ( .A(n21635), .B(n17570), .Z(n23549) );
  XOR U22857 ( .A(n23550), .B(n21652), .Z(n17570) );
  AND U22858 ( .A(n23551), .B(n21653), .Z(n23550) );
  XOR U22859 ( .A(n23552), .B(n23553), .Z(n21635) );
  AND U22860 ( .A(n23554), .B(n23555), .Z(n23552) );
  XOR U22861 ( .A(n23556), .B(n21648), .Z(n17191) );
  AND U22862 ( .A(n23557), .B(n21649), .Z(n23556) );
  XNOR U22863 ( .A(n23558), .B(n23559), .Z(n20085) );
  XNOR U22864 ( .A(n18100), .B(n17842), .Z(n23559) );
  XOR U22865 ( .A(n23560), .B(n20564), .Z(n17842) );
  IV U22866 ( .A(n21048), .Z(n20564) );
  XOR U22867 ( .A(round_reg[1406]), .B(n23561), .Z(n21048) );
  ANDN U22868 ( .B(n20565), .A(n23562), .Z(n23560) );
  XOR U22869 ( .A(n23563), .B(n20550), .Z(n18100) );
  XNOR U22870 ( .A(round_reg[1562]), .B(n23564), .Z(n20550) );
  ANDN U22871 ( .B(n20551), .A(n23565), .Z(n23563) );
  XNOR U22872 ( .A(n18835), .B(n23566), .Z(n23558) );
  XOR U22873 ( .A(n17999), .B(n19118), .Z(n23566) );
  XOR U22874 ( .A(n23567), .B(n20554), .Z(n19118) );
  XOR U22875 ( .A(round_reg[1436]), .B(n23568), .Z(n20554) );
  ANDN U22876 ( .B(n20555), .A(n23569), .Z(n23567) );
  XOR U22877 ( .A(n23570), .B(n20560), .Z(n17999) );
  XNOR U22878 ( .A(round_reg[1497]), .B(n21914), .Z(n20560) );
  ANDN U22879 ( .B(n20561), .A(n23571), .Z(n23570) );
  XOR U22880 ( .A(n23572), .B(n20934), .Z(n18835) );
  XOR U22881 ( .A(round_reg[1343]), .B(n22783), .Z(n20934) );
  ANDN U22882 ( .B(n20935), .A(n23573), .Z(n23572) );
  XNOR U22883 ( .A(n23574), .B(n16623), .Z(n13699) );
  XNOR U22884 ( .A(n22942), .B(n16767), .Z(n16623) );
  XNOR U22885 ( .A(n23575), .B(n23576), .Z(n22942) );
  ANDN U22886 ( .B(n23499), .A(n22917), .Z(n23575) );
  XOR U22887 ( .A(round_reg[1424]), .B(n23577), .Z(n22917) );
  AND U22888 ( .A(n16624), .B(n15109), .Z(n23574) );
  IV U22889 ( .A(n19413), .Z(n15109) );
  XOR U22890 ( .A(n20523), .B(n18763), .Z(n19413) );
  XOR U22891 ( .A(n23578), .B(n21533), .Z(n20523) );
  AND U22892 ( .A(n19370), .B(n23579), .Z(n23578) );
  XNOR U22893 ( .A(n23580), .B(n17506), .Z(n16624) );
  XNOR U22894 ( .A(n19989), .B(n19894), .Z(n17506) );
  XNOR U22895 ( .A(n23581), .B(n23582), .Z(n19894) );
  XNOR U22896 ( .A(n18589), .B(n18807), .Z(n23582) );
  XNOR U22897 ( .A(n23583), .B(n21332), .Z(n18807) );
  XNOR U22898 ( .A(round_reg[355]), .B(n23584), .Z(n21332) );
  NOR U22899 ( .A(n21246), .B(n21331), .Z(n23583) );
  XNOR U22900 ( .A(n23585), .B(n23014), .Z(n18589) );
  XNOR U22901 ( .A(round_reg[476]), .B(n23568), .Z(n23014) );
  XNOR U22902 ( .A(n21324), .B(n23586), .Z(n23581) );
  XOR U22903 ( .A(n17401), .B(n17084), .Z(n23586) );
  XNOR U22904 ( .A(n23587), .B(n21340), .Z(n17084) );
  XNOR U22905 ( .A(round_reg[574]), .B(n23588), .Z(n21340) );
  NOR U22906 ( .A(n21250), .B(n21339), .Z(n23587) );
  XNOR U22907 ( .A(n23589), .B(n21329), .Z(n17401) );
  XNOR U22908 ( .A(round_reg[578]), .B(n23252), .Z(n21329) );
  XNOR U22909 ( .A(n23590), .B(n21337), .Z(n21324) );
  XNOR U22910 ( .A(round_reg[406]), .B(n23591), .Z(n21337) );
  NOR U22911 ( .A(n21237), .B(n21336), .Z(n23590) );
  XOR U22912 ( .A(n23592), .B(n23593), .Z(n19989) );
  XNOR U22913 ( .A(n17251), .B(n16052), .Z(n23593) );
  XOR U22914 ( .A(n23594), .B(n21345), .Z(n16052) );
  XOR U22915 ( .A(round_reg[1358]), .B(n23595), .Z(n21345) );
  XNOR U22916 ( .A(round_reg[982]), .B(n23596), .Z(n21346) );
  XNOR U22917 ( .A(round_reg[935]), .B(n23260), .Z(n23165) );
  XNOR U22918 ( .A(n23597), .B(n21356), .Z(n17251) );
  XNOR U22919 ( .A(round_reg[1452]), .B(n23598), .Z(n21356) );
  ANDN U22920 ( .B(n23155), .A(n21355), .Z(n23597) );
  XNOR U22921 ( .A(round_reg[1075]), .B(n23475), .Z(n21355) );
  XOR U22922 ( .A(round_reg[643]), .B(n23599), .Z(n23155) );
  XNOR U22923 ( .A(n18708), .B(n23600), .Z(n23592) );
  XNOR U22924 ( .A(n18946), .B(n16935), .Z(n23600) );
  XNOR U22925 ( .A(n23601), .B(n21350), .Z(n16935) );
  XNOR U22926 ( .A(round_reg[1578]), .B(n23602), .Z(n21350) );
  ANDN U22927 ( .B(n23160), .A(n21349), .Z(n23601) );
  XNOR U22928 ( .A(round_reg[1214]), .B(n23588), .Z(n21349) );
  XNOR U22929 ( .A(round_reg[831]), .B(n23603), .Z(n23160) );
  XNOR U22930 ( .A(n23604), .B(n22449), .Z(n18946) );
  XOR U22931 ( .A(round_reg[1513]), .B(n22972), .Z(n22449) );
  ANDN U22932 ( .B(n23157), .A(n22448), .Z(n23604) );
  XNOR U22933 ( .A(round_reg[1124]), .B(n23482), .Z(n22448) );
  XNOR U22934 ( .A(round_reg[721]), .B(n21199), .Z(n23157) );
  XNOR U22935 ( .A(n23605), .B(n21360), .Z(n18708) );
  XNOR U22936 ( .A(round_reg[1295]), .B(n23606), .Z(n21360) );
  ANDN U22937 ( .B(n23163), .A(n21359), .Z(n23605) );
  XNOR U22938 ( .A(round_reg[1222]), .B(n23607), .Z(n21359) );
  XOR U22939 ( .A(round_reg[864]), .B(n23608), .Z(n23163) );
  XOR U22940 ( .A(n23609), .B(n23610), .Z(n16499) );
  XNOR U22941 ( .A(n9518), .B(n12342), .Z(n23610) );
  XNOR U22942 ( .A(n23611), .B(n13430), .Z(n12342) );
  XNOR U22943 ( .A(n20001), .B(n18145), .Z(n13430) );
  XOR U22944 ( .A(n20199), .B(n23612), .Z(n18145) );
  XOR U22945 ( .A(n23613), .B(n23614), .Z(n20199) );
  XNOR U22946 ( .A(n19448), .B(n16030), .Z(n23614) );
  XNOR U22947 ( .A(n23615), .B(n21733), .Z(n16030) );
  ANDN U22948 ( .B(n20004), .A(n20006), .Z(n23615) );
  XOR U22949 ( .A(round_reg[1585]), .B(n22962), .Z(n20006) );
  XOR U22950 ( .A(round_reg[35]), .B(n23584), .Z(n20004) );
  XNOR U22951 ( .A(n23616), .B(n23617), .Z(n19448) );
  ANDN U22952 ( .B(n19998), .A(n19999), .Z(n23616) );
  XOR U22953 ( .A(round_reg[1520]), .B(n23618), .Z(n19999) );
  XNOR U22954 ( .A(n18274), .B(n23619), .Z(n23613) );
  XOR U22955 ( .A(n21053), .B(n18241), .Z(n23619) );
  XOR U22956 ( .A(n23620), .B(n21729), .Z(n18241) );
  XNOR U22957 ( .A(round_reg[239]), .B(n21309), .Z(n20008) );
  XNOR U22958 ( .A(round_reg[1459]), .B(n23621), .Z(n20010) );
  XNOR U22959 ( .A(n23622), .B(n21736), .Z(n21053) );
  ANDN U22960 ( .B(n21737), .A(n23216), .Z(n23622) );
  XOR U22961 ( .A(round_reg[1302]), .B(n23596), .Z(n23216) );
  XOR U22962 ( .A(round_reg[121]), .B(n23623), .Z(n21737) );
  XNOR U22963 ( .A(n23624), .B(n21740), .Z(n18274) );
  ANDN U22964 ( .B(n21741), .A(n23430), .Z(n23624) );
  XNOR U22965 ( .A(n23625), .B(n21741), .Z(n20001) );
  XOR U22966 ( .A(round_reg[180]), .B(n22230), .Z(n21741) );
  ANDN U22967 ( .B(n23430), .A(n23431), .Z(n23625) );
  XOR U22968 ( .A(round_reg[1365]), .B(n23409), .Z(n23430) );
  XOR U22969 ( .A(n23626), .B(n17876), .Z(n16604) );
  XOR U22970 ( .A(n23628), .B(n23629), .Z(n22238) );
  XOR U22971 ( .A(n18537), .B(n19326), .Z(n23629) );
  XOR U22972 ( .A(n23630), .B(n22546), .Z(n19326) );
  ANDN U22973 ( .B(n22547), .A(n23631), .Z(n23630) );
  XNOR U22974 ( .A(n23632), .B(n22552), .Z(n18537) );
  XOR U22975 ( .A(n19062), .B(n23634), .Z(n23628) );
  XOR U22976 ( .A(n18837), .B(n18472), .Z(n23634) );
  XNOR U22977 ( .A(n23635), .B(n22557), .Z(n18472) );
  AND U22978 ( .A(n23636), .B(n22558), .Z(n23635) );
  XNOR U22979 ( .A(n23637), .B(n22561), .Z(n18837) );
  ANDN U22980 ( .B(n22562), .A(n23638), .Z(n23637) );
  XNOR U22981 ( .A(n23639), .B(n22565), .Z(n19062) );
  ANDN U22982 ( .B(n22566), .A(n23640), .Z(n23639) );
  XNOR U22983 ( .A(n23641), .B(n17140), .Z(n14973) );
  IV U22984 ( .A(n17078), .Z(n17140) );
  XOR U22985 ( .A(n20096), .B(n20326), .Z(n17078) );
  XNOR U22986 ( .A(n23642), .B(n23643), .Z(n20326) );
  XOR U22987 ( .A(n18506), .B(n18220), .Z(n23643) );
  XNOR U22988 ( .A(n23644), .B(n21985), .Z(n18220) );
  AND U22989 ( .A(n23645), .B(n23646), .Z(n23644) );
  XOR U22990 ( .A(n23647), .B(n21989), .Z(n18506) );
  IV U22991 ( .A(n23648), .Z(n21989) );
  ANDN U22992 ( .B(n23649), .A(n23650), .Z(n23647) );
  XNOR U22993 ( .A(n20239), .B(n23651), .Z(n23642) );
  XOR U22994 ( .A(n16937), .B(n23652), .Z(n23651) );
  XNOR U22995 ( .A(n23653), .B(n22681), .Z(n16937) );
  IV U22996 ( .A(n23654), .Z(n22681) );
  NOR U22997 ( .A(n23655), .B(n23656), .Z(n23653) );
  XNOR U22998 ( .A(n23657), .B(n21975), .Z(n20239) );
  ANDN U22999 ( .B(n23658), .A(n23659), .Z(n23657) );
  XNOR U23000 ( .A(n23660), .B(n23661), .Z(n20096) );
  XOR U23001 ( .A(n19014), .B(n17878), .Z(n23661) );
  XOR U23002 ( .A(n23662), .B(n23663), .Z(n17878) );
  AND U23003 ( .A(n22054), .B(n22053), .Z(n23662) );
  XOR U23004 ( .A(round_reg[213]), .B(n23664), .Z(n22054) );
  XOR U23005 ( .A(n23665), .B(n21969), .Z(n19014) );
  AND U23006 ( .A(n22047), .B(n22046), .Z(n23665) );
  XOR U23007 ( .A(round_reg[261]), .B(n22206), .Z(n22047) );
  XNOR U23008 ( .A(n17985), .B(n23666), .Z(n23660) );
  XNOR U23009 ( .A(n18402), .B(n17854), .Z(n23666) );
  XOR U23010 ( .A(n23667), .B(n21956), .Z(n17854) );
  ANDN U23011 ( .B(n22056), .A(n22057), .Z(n23667) );
  XNOR U23012 ( .A(round_reg[9]), .B(n23668), .Z(n22057) );
  XNOR U23013 ( .A(n23669), .B(n21961), .Z(n18402) );
  AND U23014 ( .A(n22044), .B(n22043), .Z(n23669) );
  XOR U23015 ( .A(round_reg[95]), .B(n23670), .Z(n22044) );
  XNOR U23016 ( .A(n23671), .B(n21952), .Z(n17985) );
  AND U23017 ( .A(n22051), .B(n22050), .Z(n23671) );
  XOR U23018 ( .A(round_reg[154]), .B(n23672), .Z(n22051) );
  XNOR U23019 ( .A(n23673), .B(n13437), .Z(n9518) );
  IV U23020 ( .A(n16608), .Z(n13437) );
  XNOR U23021 ( .A(n21644), .B(n18119), .Z(n16608) );
  XNOR U23022 ( .A(n23674), .B(n23675), .Z(n21644) );
  ANDN U23023 ( .B(n23553), .A(n23555), .Z(n23674) );
  NOR U23024 ( .A(n16607), .B(n14971), .Z(n23673) );
  XNOR U23025 ( .A(n23676), .B(n17595), .Z(n14971) );
  XNOR U23026 ( .A(n19956), .B(n20206), .Z(n17595) );
  XNOR U23027 ( .A(n23677), .B(n23678), .Z(n20206) );
  XNOR U23028 ( .A(n17906), .B(n18012), .Z(n23678) );
  XNOR U23029 ( .A(n23679), .B(n23680), .Z(n18012) );
  AND U23030 ( .A(n22193), .B(n23681), .Z(n23679) );
  XNOR U23031 ( .A(n23682), .B(n23683), .Z(n17906) );
  AND U23032 ( .A(n22189), .B(n23684), .Z(n23682) );
  XOR U23033 ( .A(n19070), .B(n23685), .Z(n23677) );
  XOR U23034 ( .A(n18554), .B(n15825), .Z(n23685) );
  XNOR U23035 ( .A(n23686), .B(n23687), .Z(n15825) );
  ANDN U23036 ( .B(n22180), .A(n23688), .Z(n23686) );
  XNOR U23037 ( .A(n23689), .B(n23690), .Z(n18554) );
  AND U23038 ( .A(n22185), .B(n23691), .Z(n23689) );
  XNOR U23039 ( .A(n23692), .B(n23693), .Z(n19070) );
  ANDN U23040 ( .B(n22176), .A(n23694), .Z(n23692) );
  XOR U23041 ( .A(n23695), .B(n23696), .Z(n19956) );
  XOR U23042 ( .A(n23697), .B(n19306), .Z(n23696) );
  XOR U23043 ( .A(n23698), .B(n23699), .Z(n19306) );
  XOR U23044 ( .A(n17799), .B(n23701), .Z(n23695) );
  XOR U23045 ( .A(n18450), .B(n20612), .Z(n23701) );
  XNOR U23046 ( .A(n23702), .B(n23703), .Z(n20612) );
  ANDN U23047 ( .B(n21069), .A(n23704), .Z(n23702) );
  XNOR U23048 ( .A(n23705), .B(n23706), .Z(n18450) );
  XNOR U23049 ( .A(n23708), .B(n23709), .Z(n17799) );
  IV U23050 ( .A(n19421), .Z(n16607) );
  XOR U23051 ( .A(n21527), .B(n23712), .Z(n19421) );
  XOR U23052 ( .A(n21907), .B(n20327), .Z(n21527) );
  XNOR U23053 ( .A(n23713), .B(n23714), .Z(n20327) );
  XNOR U23054 ( .A(n22477), .B(n18477), .Z(n23714) );
  XOR U23055 ( .A(n23715), .B(n21653), .Z(n18477) );
  XOR U23056 ( .A(round_reg[458]), .B(n22108), .Z(n21653) );
  ANDN U23057 ( .B(n23716), .A(n23551), .Z(n23715) );
  XNOR U23058 ( .A(n23717), .B(n23545), .Z(n22477) );
  AND U23059 ( .A(n23546), .B(n23718), .Z(n23717) );
  XOR U23060 ( .A(n22628), .B(n23719), .Z(n23713) );
  XOR U23061 ( .A(n18655), .B(n17438), .Z(n23719) );
  XNOR U23062 ( .A(n23720), .B(n21649), .Z(n17438) );
  XOR U23063 ( .A(round_reg[388]), .B(n23721), .Z(n21649) );
  ANDN U23064 ( .B(n23722), .A(n23557), .Z(n23720) );
  XNOR U23065 ( .A(n23723), .B(n21643), .Z(n18655) );
  XOR U23066 ( .A(round_reg[337]), .B(n22829), .Z(n21643) );
  XNOR U23067 ( .A(n23725), .B(n23555), .Z(n22628) );
  XOR U23068 ( .A(round_reg[556]), .B(n23726), .Z(n23555) );
  NOR U23069 ( .A(n23554), .B(n23727), .Z(n23725) );
  XOR U23070 ( .A(n23728), .B(n23729), .Z(n21907) );
  XOR U23071 ( .A(n17387), .B(n16556), .Z(n23729) );
  XOR U23072 ( .A(n23730), .B(n20555), .Z(n16556) );
  XOR U23073 ( .A(round_reg[1059]), .B(n21920), .Z(n20555) );
  ANDN U23074 ( .B(n23569), .A(n21040), .Z(n23730) );
  XNOR U23075 ( .A(n23731), .B(n20561), .Z(n17387) );
  XOR U23076 ( .A(round_reg[1108]), .B(n23732), .Z(n20561) );
  AND U23077 ( .A(n23571), .B(n21045), .Z(n23731) );
  XOR U23078 ( .A(n23540), .B(n23733), .Z(n23728) );
  XOR U23079 ( .A(n19622), .B(n18137), .Z(n23733) );
  XNOR U23080 ( .A(n23734), .B(n20551), .Z(n18137) );
  XOR U23081 ( .A(round_reg[1198]), .B(n23735), .Z(n20551) );
  ANDN U23082 ( .B(n23565), .A(n21043), .Z(n23734) );
  XNOR U23083 ( .A(n23736), .B(n20935), .Z(n19622) );
  XOR U23084 ( .A(round_reg[1270]), .B(n22278), .Z(n20935) );
  ANDN U23085 ( .B(n23573), .A(n21038), .Z(n23736) );
  XNOR U23086 ( .A(n23737), .B(n20565), .Z(n23540) );
  XOR U23087 ( .A(round_reg[966]), .B(n23738), .Z(n20565) );
  ANDN U23088 ( .B(n23562), .A(n21047), .Z(n23737) );
  XNOR U23089 ( .A(n13245), .B(n23739), .Z(n23609) );
  XOR U23090 ( .A(n9539), .B(n12177), .Z(n23739) );
  XNOR U23091 ( .A(n23740), .B(n14828), .Z(n12177) );
  IV U23092 ( .A(n16613), .Z(n14828) );
  XOR U23093 ( .A(n21021), .B(n19403), .Z(n16613) );
  IV U23094 ( .A(n19932), .Z(n19403) );
  XOR U23095 ( .A(n19737), .B(n18176), .Z(n19932) );
  XNOR U23096 ( .A(n23741), .B(n23742), .Z(n18176) );
  XNOR U23097 ( .A(n20075), .B(n15850), .Z(n23742) );
  XOR U23098 ( .A(n23743), .B(n23090), .Z(n15850) );
  IV U23099 ( .A(n21509), .Z(n23090) );
  XOR U23100 ( .A(round_reg[19]), .B(n23744), .Z(n21509) );
  AND U23101 ( .A(n21026), .B(n21024), .Z(n23743) );
  XNOR U23102 ( .A(n23746), .B(n21503), .Z(n20075) );
  XNOR U23103 ( .A(round_reg[223]), .B(n22439), .Z(n21503) );
  AND U23104 ( .A(n21016), .B(n21014), .Z(n23746) );
  IV U23105 ( .A(n21504), .Z(n21014) );
  XNOR U23106 ( .A(round_reg[1443]), .B(n23396), .Z(n21504) );
  XOR U23107 ( .A(n18956), .B(n23747), .Z(n23741) );
  XNOR U23108 ( .A(n18288), .B(n16330), .Z(n23747) );
  XNOR U23109 ( .A(n23748), .B(n23113), .Z(n16330) );
  ANDN U23110 ( .B(n21018), .A(n21019), .Z(n23748) );
  XNOR U23111 ( .A(round_reg[1504]), .B(n23608), .Z(n21018) );
  XNOR U23112 ( .A(n23749), .B(n21500), .Z(n18288) );
  XNOR U23113 ( .A(round_reg[105]), .B(n23750), .Z(n21500) );
  ANDN U23114 ( .B(n21028), .A(n21029), .Z(n23749) );
  XNOR U23115 ( .A(n23751), .B(n21512), .Z(n18956) );
  XOR U23116 ( .A(round_reg[164]), .B(n23482), .Z(n21512) );
  ANDN U23117 ( .B(n21513), .A(n23752), .Z(n23751) );
  XOR U23118 ( .A(n23753), .B(n23754), .Z(n19737) );
  XOR U23119 ( .A(n17486), .B(n20945), .Z(n23754) );
  XOR U23120 ( .A(n23755), .B(n23100), .Z(n20945) );
  ANDN U23121 ( .B(n20991), .A(n20992), .Z(n23755) );
  XNOR U23122 ( .A(n23756), .B(n23104), .Z(n17486) );
  ANDN U23123 ( .B(n20995), .A(n20997), .Z(n23756) );
  XOR U23124 ( .A(n20781), .B(n23757), .Z(n23753) );
  XOR U23125 ( .A(n16475), .B(n23758), .Z(n23757) );
  XNOR U23126 ( .A(n23759), .B(n23107), .Z(n16475) );
  ANDN U23127 ( .B(n21000), .A(n21001), .Z(n23759) );
  XNOR U23128 ( .A(n23760), .B(n23097), .Z(n20781) );
  AND U23129 ( .A(n21006), .B(n21004), .Z(n23760) );
  XOR U23130 ( .A(n23761), .B(n21513), .Z(n21021) );
  XNOR U23131 ( .A(round_reg[1349]), .B(n23762), .Z(n21513) );
  AND U23132 ( .A(n23092), .B(n23752), .Z(n23761) );
  ANDN U23133 ( .B(n16614), .A(n14965), .Z(n23740) );
  XNOR U23134 ( .A(n23763), .B(n18215), .Z(n14965) );
  XOR U23135 ( .A(n22881), .B(n23764), .Z(n18215) );
  XOR U23136 ( .A(n23765), .B(n23766), .Z(n22881) );
  XOR U23137 ( .A(n20319), .B(n16807), .Z(n23766) );
  XOR U23138 ( .A(n23767), .B(n22315), .Z(n16807) );
  ANDN U23139 ( .B(n22316), .A(n22127), .Z(n23767) );
  XNOR U23140 ( .A(n23768), .B(n22318), .Z(n20319) );
  ANDN U23141 ( .B(n22319), .A(n22137), .Z(n23768) );
  XOR U23142 ( .A(n17070), .B(n23769), .Z(n23765) );
  XOR U23143 ( .A(n19396), .B(n20465), .Z(n23769) );
  XNOR U23144 ( .A(n23770), .B(n22307), .Z(n20465) );
  ANDN U23145 ( .B(n22308), .A(n22133), .Z(n23770) );
  XNOR U23146 ( .A(n23771), .B(n22312), .Z(n19396) );
  ANDN U23147 ( .B(n22313), .A(n23772), .Z(n23771) );
  XNOR U23148 ( .A(n23773), .B(n22304), .Z(n17070) );
  ANDN U23149 ( .B(n22305), .A(n22123), .Z(n23773) );
  XNOR U23150 ( .A(n23310), .B(n15831), .Z(n16614) );
  XOR U23151 ( .A(n22701), .B(n18907), .Z(n15831) );
  XNOR U23152 ( .A(n23774), .B(n23775), .Z(n18907) );
  XOR U23153 ( .A(n18754), .B(n20494), .Z(n23775) );
  XNOR U23154 ( .A(n23776), .B(n19858), .Z(n20494) );
  XOR U23155 ( .A(round_reg[659]), .B(n23744), .Z(n19858) );
  ANDN U23156 ( .B(n22228), .A(n19923), .Z(n23776) );
  XOR U23157 ( .A(round_reg[248]), .B(n23777), .Z(n19923) );
  XNOR U23158 ( .A(round_reg[593]), .B(n23778), .Z(n22228) );
  XNOR U23159 ( .A(n23779), .B(n19862), .Z(n18754) );
  IV U23160 ( .A(n22232), .Z(n19862) );
  XOR U23161 ( .A(round_reg[737]), .B(n23780), .Z(n22232) );
  NOR U23162 ( .A(n23320), .B(n22231), .Z(n23779) );
  XNOR U23163 ( .A(round_reg[370]), .B(n23781), .Z(n22231) );
  IV U23164 ( .A(n20778), .Z(n23320) );
  XOR U23165 ( .A(round_reg[296]), .B(n23009), .Z(n20778) );
  XOR U23166 ( .A(n20393), .B(n23782), .Z(n23774) );
  XNOR U23167 ( .A(n19485), .B(n18433), .Z(n23782) );
  XNOR U23168 ( .A(n23783), .B(n19849), .Z(n18433) );
  XOR U23169 ( .A(round_reg[783]), .B(n23784), .Z(n19849) );
  ANDN U23170 ( .B(n19921), .A(n22222), .Z(n23783) );
  XNOR U23171 ( .A(round_reg[421]), .B(n22515), .Z(n22222) );
  XNOR U23172 ( .A(round_reg[44]), .B(n23785), .Z(n19921) );
  XNOR U23173 ( .A(n23786), .B(n19854), .Z(n19485) );
  XNOR U23174 ( .A(round_reg[880]), .B(n23618), .Z(n19854) );
  ANDN U23175 ( .B(n22226), .A(n19918), .Z(n23786) );
  XNOR U23176 ( .A(round_reg[66]), .B(n23787), .Z(n19918) );
  XOR U23177 ( .A(round_reg[491]), .B(n23389), .Z(n22226) );
  XNOR U23178 ( .A(n23788), .B(n19845), .Z(n20393) );
  XOR U23179 ( .A(round_reg[951]), .B(n23789), .Z(n19845) );
  ANDN U23180 ( .B(n19925), .A(n22219), .Z(n23788) );
  XNOR U23181 ( .A(round_reg[525]), .B(n23502), .Z(n22219) );
  XNOR U23182 ( .A(n23790), .B(n23791), .Z(n22701) );
  XNOR U23183 ( .A(n16025), .B(n19819), .Z(n23791) );
  XOR U23184 ( .A(n23792), .B(n22422), .Z(n19819) );
  AND U23185 ( .A(n23308), .B(n23306), .Z(n23792) );
  XOR U23186 ( .A(round_reg[1167]), .B(n23793), .Z(n23306) );
  XNOR U23187 ( .A(round_reg[784]), .B(n23577), .Z(n23308) );
  XNOR U23188 ( .A(n23794), .B(n22416), .Z(n16025) );
  AND U23189 ( .A(n22081), .B(n22415), .Z(n23794) );
  IV U23190 ( .A(n23312), .Z(n22415) );
  XNOR U23191 ( .A(round_reg[1028]), .B(n23721), .Z(n23312) );
  XNOR U23192 ( .A(round_reg[660]), .B(n21318), .Z(n22081) );
  XNOR U23193 ( .A(n17377), .B(n23795), .Z(n23790) );
  XOR U23194 ( .A(n21660), .B(n22214), .Z(n23795) );
  XNOR U23195 ( .A(n23796), .B(n22411), .Z(n22214) );
  AND U23196 ( .A(n22085), .B(n23797), .Z(n23796) );
  XNOR U23197 ( .A(n23798), .B(n22418), .Z(n21660) );
  AND U23198 ( .A(n22419), .B(n22095), .Z(n23798) );
  IV U23199 ( .A(n23304), .Z(n22095) );
  XOR U23200 ( .A(round_reg[952]), .B(n21775), .Z(n23304) );
  XOR U23201 ( .A(round_reg[999]), .B(n23799), .Z(n22419) );
  XOR U23202 ( .A(n23800), .B(n22407), .Z(n17377) );
  ANDN U23203 ( .B(n23314), .A(n22091), .Z(n23800) );
  XOR U23204 ( .A(round_reg[881]), .B(n23801), .Z(n22091) );
  XOR U23205 ( .A(round_reg[1239]), .B(n22687), .Z(n23314) );
  XOR U23206 ( .A(n23802), .B(n22410), .Z(n23310) );
  IV U23207 ( .A(n23797), .Z(n22410) );
  XOR U23208 ( .A(round_reg[1141]), .B(n23803), .Z(n23797) );
  ANDN U23209 ( .B(n22087), .A(n22085), .Z(n23802) );
  XNOR U23210 ( .A(round_reg[738]), .B(n23804), .Z(n22085) );
  XNOR U23211 ( .A(n23805), .B(n13440), .Z(n9539) );
  XOR U23212 ( .A(n22946), .B(n16957), .Z(n13440) );
  IV U23213 ( .A(n16767), .Z(n16957) );
  XOR U23214 ( .A(n20609), .B(n22786), .Z(n16767) );
  XNOR U23215 ( .A(n23806), .B(n23807), .Z(n22786) );
  XNOR U23216 ( .A(n16664), .B(n18702), .Z(n23807) );
  XNOR U23217 ( .A(n23808), .B(n22936), .Z(n18702) );
  ANDN U23218 ( .B(n23809), .A(n23506), .Z(n23808) );
  XNOR U23219 ( .A(n23810), .B(n22928), .Z(n16664) );
  AND U23220 ( .A(n22950), .B(n22949), .Z(n23810) );
  XNOR U23221 ( .A(round_reg[0]), .B(n23811), .Z(n22950) );
  XOR U23222 ( .A(n19546), .B(n23812), .Z(n23806) );
  XNOR U23223 ( .A(n19700), .B(n23813), .Z(n23812) );
  XOR U23224 ( .A(n23814), .B(n22932), .Z(n19700) );
  ANDN U23225 ( .B(n22944), .A(n22945), .Z(n23814) );
  XOR U23226 ( .A(round_reg[86]), .B(n23591), .Z(n22945) );
  XNOR U23227 ( .A(n23815), .B(n22922), .Z(n19546) );
  ANDN U23228 ( .B(n22952), .A(n22953), .Z(n23815) );
  XNOR U23229 ( .A(round_reg[316]), .B(n23816), .Z(n22953) );
  XOR U23230 ( .A(n23817), .B(n23818), .Z(n20609) );
  XOR U23231 ( .A(n23819), .B(n18280), .Z(n23818) );
  XOR U23232 ( .A(n23820), .B(n23821), .Z(n18280) );
  ANDN U23233 ( .B(n22869), .A(n22871), .Z(n23820) );
  XOR U23234 ( .A(n20846), .B(n23822), .Z(n23817) );
  XOR U23235 ( .A(n17927), .B(n19978), .Z(n23822) );
  XNOR U23236 ( .A(n23823), .B(n22912), .Z(n19978) );
  ANDN U23237 ( .B(n22864), .A(n22866), .Z(n23823) );
  XNOR U23238 ( .A(n23824), .B(n23825), .Z(n17927) );
  ANDN U23239 ( .B(n22873), .A(n22874), .Z(n23824) );
  XNOR U23240 ( .A(n23826), .B(n22902), .Z(n20846) );
  AND U23241 ( .A(n22879), .B(n22877), .Z(n23826) );
  XNOR U23242 ( .A(n23827), .B(n23809), .Z(n22946) );
  ANDN U23243 ( .B(n23506), .A(n22934), .Z(n23827) );
  XOR U23244 ( .A(round_reg[1394]), .B(n23197), .Z(n22934) );
  XOR U23245 ( .A(n23828), .B(n23829), .Z(n23197) );
  ANDN U23246 ( .B(n16616), .A(n17659), .Z(n23805) );
  XNOR U23247 ( .A(n17810), .B(n19725), .Z(n17659) );
  XNOR U23248 ( .A(n23830), .B(n20448), .Z(n19725) );
  AND U23249 ( .A(n19478), .B(n23831), .Z(n23830) );
  IV U23250 ( .A(n21305), .Z(n19478) );
  XOR U23251 ( .A(round_reg[850]), .B(n22645), .Z(n21305) );
  IV U23252 ( .A(n20314), .Z(n17810) );
  XNOR U23253 ( .A(n21445), .B(n18389), .Z(n16616) );
  XNOR U23254 ( .A(n19463), .B(n19707), .Z(n18389) );
  XNOR U23255 ( .A(n23832), .B(n23833), .Z(n19707) );
  XNOR U23256 ( .A(n18010), .B(n18886), .Z(n23833) );
  XOR U23257 ( .A(n23834), .B(n23835), .Z(n18886) );
  ANDN U23258 ( .B(n21441), .A(n21442), .Z(n23834) );
  XOR U23259 ( .A(n23836), .B(n23837), .Z(n18010) );
  AND U23260 ( .A(n23838), .B(n23839), .Z(n23836) );
  XOR U23261 ( .A(n19773), .B(n23840), .Z(n23832) );
  XOR U23262 ( .A(n17856), .B(n18659), .Z(n23840) );
  XOR U23263 ( .A(n23841), .B(n23842), .Z(n18659) );
  ANDN U23264 ( .B(n21447), .A(n21448), .Z(n23841) );
  XOR U23265 ( .A(n23843), .B(n23844), .Z(n17856) );
  AND U23266 ( .A(n21453), .B(n21451), .Z(n23843) );
  XOR U23267 ( .A(n23845), .B(n23846), .Z(n19773) );
  AND U23268 ( .A(n23185), .B(n23187), .Z(n23845) );
  XOR U23269 ( .A(n23847), .B(n23848), .Z(n19463) );
  XNOR U23270 ( .A(n19713), .B(n20417), .Z(n23848) );
  XOR U23271 ( .A(n23849), .B(n21120), .Z(n20417) );
  NOR U23272 ( .A(n21471), .B(n21119), .Z(n23849) );
  XOR U23273 ( .A(round_reg[969]), .B(n23668), .Z(n21119) );
  XNOR U23274 ( .A(n23850), .B(n21102), .Z(n19713) );
  ANDN U23275 ( .B(n21103), .A(n21468), .Z(n23850) );
  XNOR U23276 ( .A(round_reg[1201]), .B(n23851), .Z(n21103) );
  XOR U23277 ( .A(n15128), .B(n23852), .Z(n23847) );
  XOR U23278 ( .A(n20038), .B(n21096), .Z(n23852) );
  XOR U23279 ( .A(n23853), .B(n21116), .Z(n21096) );
  NOR U23280 ( .A(n21115), .B(n21465), .Z(n23853) );
  XOR U23281 ( .A(round_reg[1273]), .B(n23854), .Z(n21115) );
  XNOR U23282 ( .A(n23855), .B(n21106), .Z(n20038) );
  ANDN U23283 ( .B(n21107), .A(n21457), .Z(n23855) );
  XNOR U23284 ( .A(round_reg[1062]), .B(n23856), .Z(n21107) );
  XNOR U23285 ( .A(n23857), .B(n21111), .Z(n15128) );
  ANDN U23286 ( .B(n21460), .A(n21461), .Z(n23857) );
  XOR U23287 ( .A(round_reg[1111]), .B(n23254), .Z(n21460) );
  XNOR U23288 ( .A(n23858), .B(n23839), .Z(n21445) );
  NOR U23289 ( .A(n23859), .B(n23838), .Z(n23858) );
  XNOR U23290 ( .A(n23860), .B(n14441), .Z(n13245) );
  XOR U23291 ( .A(n20595), .B(n16055), .Z(n14441) );
  XOR U23292 ( .A(n21074), .B(n20309), .Z(n16055) );
  XOR U23293 ( .A(n23861), .B(n23862), .Z(n20309) );
  XOR U23294 ( .A(n18348), .B(n20329), .Z(n23862) );
  XOR U23295 ( .A(n23863), .B(n21874), .Z(n20329) );
  ANDN U23296 ( .B(n21875), .A(n20599), .Z(n23863) );
  XOR U23297 ( .A(round_reg[788]), .B(n23732), .Z(n21875) );
  XOR U23298 ( .A(n23864), .B(n20368), .Z(n18348) );
  ANDN U23299 ( .B(n20369), .A(n20593), .Z(n23864) );
  XOR U23300 ( .A(round_reg[742]), .B(n23865), .Z(n20369) );
  XOR U23301 ( .A(n20244), .B(n23866), .Z(n23861) );
  XOR U23302 ( .A(n19129), .B(n19142), .Z(n23866) );
  XOR U23303 ( .A(n23867), .B(n20359), .Z(n19142) );
  XOR U23304 ( .A(n23869), .B(n20365), .Z(n19129) );
  ANDN U23305 ( .B(n23870), .A(n20364), .Z(n23869) );
  XOR U23306 ( .A(round_reg[885]), .B(n23871), .Z(n20364) );
  XOR U23307 ( .A(n23872), .B(n22520), .Z(n20244) );
  NOR U23308 ( .A(n20590), .B(n20589), .Z(n23872) );
  XOR U23309 ( .A(round_reg[664]), .B(n22816), .Z(n20589) );
  XOR U23310 ( .A(n23873), .B(n23874), .Z(n21074) );
  XNOR U23311 ( .A(n18873), .B(n18094), .Z(n23874) );
  XNOR U23312 ( .A(n23875), .B(n20352), .Z(n18094) );
  XNOR U23313 ( .A(round_reg[425]), .B(n23876), .Z(n20352) );
  XNOR U23314 ( .A(round_reg[1598]), .B(n23877), .Z(n22009) );
  XOR U23315 ( .A(round_reg[48]), .B(n23445), .Z(n20351) );
  XNOR U23316 ( .A(n23878), .B(n20339), .Z(n18873) );
  XNOR U23317 ( .A(round_reg[374]), .B(n23879), .Z(n20339) );
  XNOR U23318 ( .A(round_reg[300]), .B(n23300), .Z(n20338) );
  XNOR U23319 ( .A(n18969), .B(n23880), .Z(n23873) );
  XOR U23320 ( .A(n18726), .B(n18984), .Z(n23880) );
  XNOR U23321 ( .A(n23881), .B(n20335), .Z(n18984) );
  XNOR U23322 ( .A(round_reg[597]), .B(n23266), .Z(n20335) );
  NOR U23323 ( .A(n22647), .B(n20334), .Z(n23881) );
  XNOR U23324 ( .A(round_reg[252]), .B(n23147), .Z(n20334) );
  IV U23325 ( .A(n22634), .Z(n22647) );
  XNOR U23326 ( .A(round_reg[1408]), .B(n23011), .Z(n22634) );
  XNOR U23327 ( .A(n23882), .B(n20348), .Z(n18726) );
  XNOR U23328 ( .A(round_reg[495]), .B(n21196), .Z(n20348) );
  AND U23329 ( .A(n20347), .B(n22012), .Z(n23882) );
  XOR U23330 ( .A(round_reg[70]), .B(n23883), .Z(n20347) );
  XNOR U23331 ( .A(n23884), .B(n20344), .Z(n18969) );
  XNOR U23332 ( .A(round_reg[529]), .B(n23885), .Z(n20344) );
  ANDN U23333 ( .B(n22017), .A(n20343), .Z(n23884) );
  XNOR U23334 ( .A(round_reg[129]), .B(n23886), .Z(n20343) );
  XOR U23335 ( .A(round_reg[1378]), .B(n23887), .Z(n22017) );
  XOR U23336 ( .A(n23888), .B(n20358), .Z(n20595) );
  XOR U23337 ( .A(round_reg[956]), .B(n23816), .Z(n20358) );
  ANDN U23338 ( .B(n23868), .A(n23889), .Z(n23888) );
  ANDN U23339 ( .B(n16619), .A(n14967), .Z(n23860) );
  XNOR U23340 ( .A(n20812), .B(n15208), .Z(n14967) );
  XOR U23341 ( .A(n23890), .B(n23891), .Z(n20812) );
  ANDN U23342 ( .B(n21266), .A(n21268), .Z(n23890) );
  XOR U23343 ( .A(n21221), .B(n19337), .Z(n16619) );
  XNOR U23344 ( .A(n19248), .B(n20068), .Z(n19337) );
  XNOR U23345 ( .A(n23892), .B(n23893), .Z(n20068) );
  XNOR U23346 ( .A(n18877), .B(n18257), .Z(n23893) );
  XOR U23347 ( .A(n23894), .B(n20188), .Z(n18257) );
  XNOR U23348 ( .A(round_reg[645]), .B(n23895), .Z(n20188) );
  AND U23349 ( .A(n20187), .B(n21228), .Z(n23894) );
  XNOR U23350 ( .A(round_reg[579]), .B(n23896), .Z(n20187) );
  XNOR U23351 ( .A(n23897), .B(n20698), .Z(n18877) );
  XOR U23352 ( .A(round_reg[723]), .B(n21610), .Z(n20698) );
  XOR U23353 ( .A(n18654), .B(n23899), .Z(n23892) );
  XOR U23354 ( .A(n19892), .B(n16951), .Z(n23899) );
  XOR U23355 ( .A(n23900), .B(n20178), .Z(n16951) );
  XNOR U23356 ( .A(round_reg[769]), .B(n23886), .Z(n20178) );
  ANDN U23357 ( .B(n21223), .A(n21224), .Z(n23900) );
  IV U23358 ( .A(n20177), .Z(n21223) );
  XNOR U23359 ( .A(round_reg[407]), .B(n23486), .Z(n20177) );
  XOR U23360 ( .A(n23901), .B(n20184), .Z(n19892) );
  XNOR U23361 ( .A(round_reg[866]), .B(n23480), .Z(n20184) );
  ANDN U23362 ( .B(n21230), .A(n20183), .Z(n23901) );
  XNOR U23363 ( .A(round_reg[477]), .B(n23902), .Z(n20183) );
  XNOR U23364 ( .A(n23903), .B(n20173), .Z(n18654) );
  XOR U23365 ( .A(round_reg[937]), .B(n22760), .Z(n20173) );
  XNOR U23366 ( .A(round_reg[575]), .B(n23904), .Z(n20174) );
  XOR U23367 ( .A(n23905), .B(n23906), .Z(n19248) );
  XNOR U23368 ( .A(n23580), .B(n21825), .Z(n23906) );
  XOR U23369 ( .A(n23907), .B(n21339), .Z(n21825) );
  XNOR U23370 ( .A(round_reg[174]), .B(n23908), .Z(n21339) );
  AND U23371 ( .A(n21252), .B(n21250), .Z(n23907) );
  XOR U23372 ( .A(round_reg[1359]), .B(n21605), .Z(n21250) );
  XNOR U23373 ( .A(round_reg[983]), .B(n22635), .Z(n21252) );
  XOR U23374 ( .A(n23909), .B(n21336), .Z(n23580) );
  XNOR U23375 ( .A(round_reg[29]), .B(n23910), .Z(n21336) );
  ANDN U23376 ( .B(n21237), .A(n21238), .Z(n23909) );
  XOR U23377 ( .A(round_reg[1215]), .B(n23904), .Z(n21238) );
  XOR U23378 ( .A(round_reg[1579]), .B(n22375), .Z(n21237) );
  XOR U23379 ( .A(n17505), .B(n23911), .Z(n23905) );
  XOR U23380 ( .A(n18662), .B(n23135), .Z(n23911) );
  XOR U23381 ( .A(n23912), .B(n21328), .Z(n23135) );
  XNOR U23382 ( .A(round_reg[233]), .B(n22972), .Z(n21328) );
  NOR U23383 ( .A(n21241), .B(n21242), .Z(n23912) );
  XOR U23384 ( .A(round_reg[1076]), .B(n23289), .Z(n21242) );
  XNOR U23385 ( .A(round_reg[1453]), .B(n23413), .Z(n21241) );
  XOR U23386 ( .A(n23913), .B(n23020), .Z(n18662) );
  XOR U23387 ( .A(round_reg[115]), .B(n23914), .Z(n23020) );
  ANDN U23388 ( .B(n21256), .A(n21254), .Z(n23913) );
  XNOR U23389 ( .A(round_reg[1296]), .B(n23915), .Z(n21254) );
  XNOR U23390 ( .A(round_reg[1223]), .B(n23916), .Z(n21256) );
  XOR U23391 ( .A(n23917), .B(n21331), .Z(n17505) );
  XNOR U23392 ( .A(round_reg[281]), .B(n23918), .Z(n21331) );
  ANDN U23393 ( .B(n21246), .A(n21248), .Z(n23917) );
  XOR U23394 ( .A(round_reg[1125]), .B(n23919), .Z(n21248) );
  XOR U23395 ( .A(round_reg[1514]), .B(n23920), .Z(n21246) );
  XNOR U23396 ( .A(n23921), .B(n20705), .Z(n21221) );
  XNOR U23397 ( .A(round_reg[356]), .B(n23201), .Z(n20705) );
  NOR U23398 ( .A(n20696), .B(n23898), .Z(n23921) );
  XNOR U23399 ( .A(n23922), .B(n16627), .Z(n19410) );
  XNOR U23400 ( .A(n15329), .B(n23512), .Z(n16627) );
  XOR U23401 ( .A(n23923), .B(n23924), .Z(n23512) );
  AND U23402 ( .A(n21163), .B(n23925), .Z(n23923) );
  XOR U23403 ( .A(n21580), .B(n20807), .Z(n15329) );
  XOR U23404 ( .A(n23926), .B(n23927), .Z(n20807) );
  XNOR U23405 ( .A(n16606), .B(n16927), .Z(n23927) );
  XOR U23406 ( .A(n23928), .B(n23929), .Z(n16927) );
  ANDN U23407 ( .B(n21178), .A(n23514), .Z(n23928) );
  XOR U23408 ( .A(round_reg[898]), .B(n23930), .Z(n21178) );
  XNOR U23409 ( .A(n23931), .B(n23932), .Z(n16606) );
  NOR U23410 ( .A(n23925), .B(n23924), .Z(n23931) );
  IV U23411 ( .A(n21161), .Z(n23925) );
  XOR U23412 ( .A(round_reg[794]), .B(n23672), .Z(n21161) );
  XOR U23413 ( .A(n16339), .B(n23933), .Z(n23926) );
  XOR U23414 ( .A(n18847), .B(n18487), .Z(n23933) );
  XNOR U23415 ( .A(n23934), .B(n23935), .Z(n18487) );
  ANDN U23416 ( .B(n21174), .A(n23522), .Z(n23934) );
  XOR U23417 ( .A(round_reg[891]), .B(n21617), .Z(n21174) );
  XNOR U23418 ( .A(n23936), .B(n23937), .Z(n18847) );
  AND U23419 ( .A(n23519), .B(n21170), .Z(n23936) );
  IV U23420 ( .A(n23520), .Z(n21170) );
  XOR U23421 ( .A(round_reg[670]), .B(n23246), .Z(n23520) );
  XNOR U23422 ( .A(n23938), .B(n23939), .Z(n16339) );
  AND U23423 ( .A(n23517), .B(n21165), .Z(n23938) );
  XOR U23424 ( .A(round_reg[748]), .B(n23940), .Z(n21165) );
  XOR U23425 ( .A(n23941), .B(n23942), .Z(n21580) );
  XNOR U23426 ( .A(n16099), .B(n18544), .Z(n23942) );
  XNOR U23427 ( .A(n23943), .B(n20257), .Z(n18544) );
  XNOR U23428 ( .A(round_reg[793]), .B(n23944), .Z(n20257) );
  AND U23429 ( .A(n20258), .B(n21403), .Z(n23943) );
  XNOR U23430 ( .A(n23945), .B(n20267), .Z(n16099) );
  XOR U23431 ( .A(round_reg[747]), .B(n23946), .Z(n20267) );
  AND U23432 ( .A(n20268), .B(n21400), .Z(n23945) );
  XOR U23433 ( .A(n19446), .B(n23947), .Z(n23941) );
  XOR U23434 ( .A(n18719), .B(n20247), .Z(n23947) );
  XOR U23435 ( .A(n23948), .B(n23452), .Z(n20247) );
  IV U23436 ( .A(n23455), .Z(n23452) );
  XOR U23437 ( .A(round_reg[669]), .B(n23910), .Z(n23455) );
  ANDN U23438 ( .B(n23456), .A(n21391), .Z(n23948) );
  XOR U23439 ( .A(n23949), .B(n20264), .Z(n18719) );
  XOR U23440 ( .A(round_reg[890]), .B(n23249), .Z(n20264) );
  ANDN U23441 ( .B(n20263), .A(n23950), .Z(n23949) );
  XOR U23442 ( .A(n23951), .B(n20254), .Z(n19446) );
  XOR U23443 ( .A(round_reg[897]), .B(n23952), .Z(n20254) );
  ANDN U23444 ( .B(n20253), .A(n21395), .Z(n23951) );
  XOR U23445 ( .A(n15837), .B(n23953), .Z(n15113) );
  IV U23446 ( .A(n16416), .Z(n15837) );
  XOR U23447 ( .A(n20236), .B(n19637), .Z(n16416) );
  XNOR U23448 ( .A(n23954), .B(n23955), .Z(n19637) );
  XOR U23449 ( .A(n18149), .B(n18139), .Z(n23955) );
  XOR U23450 ( .A(n23956), .B(n20599), .Z(n18139) );
  XOR U23451 ( .A(round_reg[426]), .B(n23528), .Z(n20599) );
  AND U23452 ( .A(n20600), .B(n23957), .Z(n23956) );
  XNOR U23453 ( .A(n23958), .B(n20593), .Z(n18149) );
  XNOR U23454 ( .A(round_reg[375]), .B(n23959), .Z(n20593) );
  ANDN U23455 ( .B(n20594), .A(n20367), .Z(n23958) );
  XOR U23456 ( .A(n20423), .B(n23960), .Z(n23954) );
  XNOR U23457 ( .A(n17891), .B(n20585), .Z(n23960) );
  XNOR U23458 ( .A(n23961), .B(n23868), .Z(n20585) );
  XOR U23459 ( .A(round_reg[530]), .B(n22645), .Z(n23868) );
  ANDN U23460 ( .B(n23889), .A(n20357), .Z(n23961) );
  XNOR U23461 ( .A(n23962), .B(n23870), .Z(n17891) );
  IV U23462 ( .A(n20603), .Z(n23870) );
  XOR U23463 ( .A(round_reg[496]), .B(n23963), .Z(n20603) );
  NOR U23464 ( .A(n20602), .B(n20363), .Z(n23962) );
  XNOR U23465 ( .A(n23964), .B(n20590), .Z(n20423) );
  XNOR U23466 ( .A(round_reg[598]), .B(n23965), .Z(n20590) );
  ANDN U23467 ( .B(n20591), .A(n22519), .Z(n23964) );
  XOR U23468 ( .A(n23966), .B(n23967), .Z(n20236) );
  XNOR U23469 ( .A(n19458), .B(n20227), .Z(n23967) );
  XOR U23470 ( .A(n23968), .B(n23180), .Z(n20227) );
  XOR U23471 ( .A(n23971), .B(n23176), .Z(n19458) );
  XNOR U23472 ( .A(n19305), .B(n23973), .Z(n23966) );
  XOR U23473 ( .A(n19265), .B(n18546), .Z(n23973) );
  XOR U23474 ( .A(n23974), .B(n23182), .Z(n18546) );
  ANDN U23475 ( .B(n23975), .A(n22252), .Z(n23974) );
  XNOR U23476 ( .A(n23976), .B(n23173), .Z(n19265) );
  AND U23477 ( .A(n23977), .B(n22256), .Z(n23976) );
  IV U23478 ( .A(n23978), .Z(n22256) );
  XNOR U23479 ( .A(n23979), .B(n23171), .Z(n19305) );
  IV U23480 ( .A(n23980), .Z(n23171) );
  NOR U23481 ( .A(n23981), .B(n22242), .Z(n23979) );
  XOR U23482 ( .A(n19810), .B(n18759), .Z(n15115) );
  XOR U23483 ( .A(n22695), .B(n23982), .Z(n18759) );
  XOR U23484 ( .A(n23983), .B(n23984), .Z(n22695) );
  XOR U23485 ( .A(n18706), .B(n19985), .Z(n23984) );
  XOR U23486 ( .A(n23985), .B(n21230), .Z(n19985) );
  XNOR U23487 ( .A(round_reg[116]), .B(n23289), .Z(n21230) );
  XNOR U23488 ( .A(round_reg[1297]), .B(n22829), .Z(n20702) );
  XOR U23489 ( .A(round_reg[1224]), .B(n23986), .Z(n20182) );
  XNOR U23490 ( .A(n23987), .B(n23898), .Z(n18706) );
  XNOR U23491 ( .A(round_reg[282]), .B(n22640), .Z(n23898) );
  AND U23492 ( .A(n20697), .B(n20696), .Z(n23987) );
  XOR U23493 ( .A(round_reg[1515]), .B(n22112), .Z(n20696) );
  XOR U23494 ( .A(round_reg[1126]), .B(n23988), .Z(n20697) );
  XOR U23495 ( .A(n20276), .B(n23989), .Z(n23983) );
  XNOR U23496 ( .A(n19578), .B(n21218), .Z(n23989) );
  XNOR U23497 ( .A(n23990), .B(n21224), .Z(n21218) );
  XOR U23498 ( .A(round_reg[30]), .B(n23246), .Z(n21224) );
  XNOR U23499 ( .A(round_reg[1580]), .B(n23300), .Z(n20700) );
  XOR U23500 ( .A(round_reg[1152]), .B(n23991), .Z(n20176) );
  XNOR U23501 ( .A(n23992), .B(n21228), .Z(n19578) );
  XNOR U23502 ( .A(round_reg[234]), .B(n23920), .Z(n21228) );
  AND U23503 ( .A(n20186), .B(n21227), .Z(n23992) );
  XOR U23504 ( .A(round_reg[1454]), .B(n23908), .Z(n21227) );
  XNOR U23505 ( .A(round_reg[1077]), .B(n23993), .Z(n20186) );
  XNOR U23506 ( .A(n23994), .B(n21232), .Z(n20276) );
  XOR U23507 ( .A(round_reg[175]), .B(n21196), .Z(n21232) );
  ANDN U23508 ( .B(n21233), .A(n20172), .Z(n23994) );
  XNOR U23509 ( .A(round_reg[984]), .B(n22816), .Z(n20172) );
  IV U23510 ( .A(n23995), .Z(n22816) );
  XOR U23511 ( .A(round_reg[1360]), .B(n22445), .Z(n21233) );
  XNOR U23512 ( .A(n23996), .B(n19950), .Z(n19810) );
  AND U23513 ( .A(n21188), .B(n20624), .Z(n23996) );
  XNOR U23514 ( .A(round_reg[1516]), .B(n23726), .Z(n20624) );
  NOR U23515 ( .A(n7076), .B(n9262), .Z(n23332) );
  XNOR U23516 ( .A(n15152), .B(n11859), .Z(n9262) );
  IV U23517 ( .A(n11666), .Z(n11859) );
  XOR U23518 ( .A(n14430), .B(n12578), .Z(n11666) );
  XNOR U23519 ( .A(n23997), .B(n23998), .Z(n12578) );
  XNOR U23520 ( .A(n12706), .B(n12991), .Z(n23998) );
  XNOR U23521 ( .A(n23999), .B(n15264), .Z(n12991) );
  XNOR U23522 ( .A(n18217), .B(n23339), .Z(n15264) );
  XNOR U23523 ( .A(n24000), .B(n22738), .Z(n23339) );
  ANDN U23524 ( .B(n24001), .A(n23063), .Z(n24000) );
  XOR U23525 ( .A(n19960), .B(n21750), .Z(n18217) );
  XOR U23526 ( .A(n24002), .B(n24003), .Z(n21750) );
  XOR U23527 ( .A(n19974), .B(n18859), .Z(n24003) );
  XOR U23528 ( .A(n24004), .B(n22727), .Z(n18859) );
  XOR U23529 ( .A(round_reg[1367]), .B(n23486), .Z(n22727) );
  ANDN U23530 ( .B(n22728), .A(n23360), .Z(n24004) );
  XOR U23531 ( .A(round_reg[991]), .B(n23325), .Z(n22728) );
  XOR U23532 ( .A(n24005), .B(n22719), .Z(n19974) );
  XNOR U23533 ( .A(round_reg[1587]), .B(n21312), .Z(n22719) );
  ANDN U23534 ( .B(n22720), .A(n23352), .Z(n24005) );
  XNOR U23535 ( .A(round_reg[1159]), .B(n24006), .Z(n22720) );
  XOR U23536 ( .A(n20710), .B(n24007), .Z(n24002) );
  XOR U23537 ( .A(n19425), .B(n16554), .Z(n24007) );
  XNOR U23538 ( .A(n24008), .B(n22710), .Z(n16554) );
  XOR U23539 ( .A(round_reg[1304]), .B(n23995), .Z(n22710) );
  ANDN U23540 ( .B(n22711), .A(n23358), .Z(n24008) );
  XOR U23541 ( .A(round_reg[1231]), .B(n22802), .Z(n22711) );
  XNOR U23542 ( .A(n24009), .B(n22723), .Z(n19425) );
  XOR U23543 ( .A(round_reg[1461]), .B(n23803), .Z(n22723) );
  ANDN U23544 ( .B(n22724), .A(n23362), .Z(n24009) );
  XNOR U23545 ( .A(round_reg[1084]), .B(n24010), .Z(n22724) );
  XOR U23546 ( .A(n24011), .B(n24012), .Z(n20710) );
  ANDN U23547 ( .B(n22715), .A(n23354), .Z(n24011) );
  XNOR U23548 ( .A(round_reg[1133]), .B(n24013), .Z(n22715) );
  XOR U23549 ( .A(n24014), .B(n24015), .Z(n19960) );
  XNOR U23550 ( .A(n16459), .B(n22705), .Z(n24015) );
  XNOR U23551 ( .A(n24016), .B(n22743), .Z(n22705) );
  XNOR U23552 ( .A(round_reg[415]), .B(n23670), .Z(n22743) );
  XOR U23553 ( .A(round_reg[38]), .B(n24017), .Z(n22744) );
  XOR U23554 ( .A(n24018), .B(n23064), .Z(n16459) );
  IV U23555 ( .A(n22737), .Z(n23064) );
  XOR U23556 ( .A(round_reg[364]), .B(n23785), .Z(n22737) );
  ANDN U23557 ( .B(n22738), .A(n24001), .Z(n24018) );
  XOR U23558 ( .A(round_reg[290]), .B(n24019), .Z(n22738) );
  XNOR U23559 ( .A(n19155), .B(n24020), .Z(n24014) );
  XNOR U23560 ( .A(n19495), .B(n19127), .Z(n24020) );
  XNOR U23561 ( .A(n24021), .B(n22733), .Z(n19127) );
  XNOR U23562 ( .A(round_reg[587]), .B(n24022), .Z(n22733) );
  ANDN U23563 ( .B(n22734), .A(n23344), .Z(n24021) );
  XNOR U23564 ( .A(round_reg[242]), .B(n24023), .Z(n22734) );
  XNOR U23565 ( .A(n24024), .B(n22748), .Z(n19495) );
  XNOR U23566 ( .A(round_reg[485]), .B(n23919), .Z(n22748) );
  AND U23567 ( .A(n22747), .B(n24025), .Z(n24024) );
  XNOR U23568 ( .A(round_reg[124]), .B(n24010), .Z(n22747) );
  IV U23569 ( .A(n24026), .Z(n24010) );
  XNOR U23570 ( .A(n24027), .B(n23053), .Z(n19155) );
  XNOR U23571 ( .A(round_reg[519]), .B(n24028), .Z(n23053) );
  ANDN U23572 ( .B(n23079), .A(n23348), .Z(n24027) );
  XOR U23573 ( .A(round_reg[183]), .B(n24029), .Z(n23079) );
  ANDN U23574 ( .B(n18131), .A(n15263), .Z(n23999) );
  XOR U23575 ( .A(n21718), .B(n17678), .Z(n15263) );
  XOR U23576 ( .A(n24030), .B(n24031), .Z(n17678) );
  XNOR U23577 ( .A(n24032), .B(n23424), .Z(n21718) );
  XOR U23578 ( .A(round_reg[872]), .B(n23397), .Z(n21744) );
  XNOR U23579 ( .A(n21639), .B(n18119), .Z(n18131) );
  XOR U23580 ( .A(n22683), .B(n20931), .Z(n18119) );
  XNOR U23581 ( .A(n24033), .B(n24034), .Z(n20931) );
  XOR U23582 ( .A(n24035), .B(n18169), .Z(n24034) );
  XOR U23583 ( .A(n24036), .B(n23722), .Z(n18169) );
  ANDN U23584 ( .B(n21647), .A(n21648), .Z(n24036) );
  XOR U23585 ( .A(n19030), .B(n24037), .Z(n24033) );
  XOR U23586 ( .A(n17233), .B(n19149), .Z(n24037) );
  XOR U23587 ( .A(n24038), .B(n23718), .Z(n19149) );
  ANDN U23588 ( .B(n24039), .A(n23544), .Z(n24038) );
  XNOR U23589 ( .A(n24040), .B(n23727), .Z(n17233) );
  ANDN U23590 ( .B(n23675), .A(n23553), .Z(n24040) );
  XNOR U23591 ( .A(round_reg[918]), .B(n23965), .Z(n23553) );
  XOR U23592 ( .A(n24041), .B(n23716), .Z(n19030) );
  ANDN U23593 ( .B(n21651), .A(n21652), .Z(n24041) );
  XNOR U23594 ( .A(round_reg[847]), .B(n23297), .Z(n21652) );
  IV U23595 ( .A(n23793), .Z(n23297) );
  XNOR U23596 ( .A(n24042), .B(n24043), .Z(n22683) );
  XOR U23597 ( .A(n18574), .B(n17938), .Z(n24043) );
  XOR U23598 ( .A(n24044), .B(n23656), .Z(n17938) );
  AND U23599 ( .A(n22682), .B(n22680), .Z(n24044) );
  XNOR U23600 ( .A(n24045), .B(n24046), .Z(n18574) );
  AND U23601 ( .A(n21980), .B(n21978), .Z(n24045) );
  XOR U23602 ( .A(n19669), .B(n24047), .Z(n24042) );
  XOR U23603 ( .A(n16794), .B(n18891), .Z(n24047) );
  XNOR U23604 ( .A(n24048), .B(n23650), .Z(n18891) );
  AND U23605 ( .A(n21990), .B(n21988), .Z(n24048) );
  XNOR U23606 ( .A(n24049), .B(n23659), .Z(n16794) );
  AND U23607 ( .A(n21976), .B(n21974), .Z(n24049) );
  XOR U23608 ( .A(n24050), .B(n23645), .Z(n19669) );
  ANDN U23609 ( .B(n21984), .A(n21986), .Z(n24050) );
  XOR U23610 ( .A(n24051), .B(n24039), .Z(n21639) );
  AND U23611 ( .A(n23545), .B(n23544), .Z(n24051) );
  XNOR U23612 ( .A(round_reg[690]), .B(n24052), .Z(n23544) );
  XNOR U23613 ( .A(round_reg[624]), .B(n24053), .Z(n23545) );
  XNOR U23614 ( .A(n24054), .B(n15280), .Z(n12706) );
  XNOR U23615 ( .A(n23697), .B(n17800), .Z(n15280) );
  XOR U23616 ( .A(n19071), .B(n20011), .Z(n17800) );
  XOR U23617 ( .A(n24055), .B(n24056), .Z(n20011) );
  XNOR U23618 ( .A(n18318), .B(n24057), .Z(n24056) );
  XOR U23619 ( .A(n24058), .B(n24059), .Z(n18318) );
  AND U23620 ( .A(n23709), .B(n23711), .Z(n24058) );
  XNOR U23621 ( .A(n22993), .B(n24060), .Z(n24055) );
  XOR U23622 ( .A(n19734), .B(n18047), .Z(n24060) );
  XOR U23623 ( .A(n24061), .B(n22164), .Z(n18047) );
  AND U23624 ( .A(n23699), .B(n23700), .Z(n24061) );
  XOR U23625 ( .A(n24062), .B(n21060), .Z(n19734) );
  ANDN U23626 ( .B(n23706), .A(n23707), .Z(n24062) );
  XOR U23627 ( .A(n24063), .B(n21064), .Z(n22993) );
  ANDN U23628 ( .B(n24064), .A(n24065), .Z(n24063) );
  XOR U23629 ( .A(n24066), .B(n24067), .Z(n19071) );
  XNOR U23630 ( .A(n16326), .B(n24068), .Z(n24067) );
  XNOR U23631 ( .A(n24069), .B(n22190), .Z(n16326) );
  ANDN U23632 ( .B(n23683), .A(n23684), .Z(n24069) );
  XNOR U23633 ( .A(n15953), .B(n24070), .Z(n24066) );
  XOR U23634 ( .A(n18800), .B(n17581), .Z(n24070) );
  XNOR U23635 ( .A(n24071), .B(n22181), .Z(n17581) );
  AND U23636 ( .A(n23688), .B(n23687), .Z(n24071) );
  XNOR U23637 ( .A(n24072), .B(n22194), .Z(n18800) );
  ANDN U23638 ( .B(n23680), .A(n23681), .Z(n24072) );
  XNOR U23639 ( .A(n24073), .B(n24074), .Z(n15953) );
  XNOR U23640 ( .A(n24075), .B(n24064), .Z(n23697) );
  AND U23641 ( .A(n21062), .B(n24065), .Z(n24075) );
  AND U23642 ( .A(n16517), .B(n15281), .Z(n24054) );
  XNOR U23643 ( .A(n17237), .B(n20800), .Z(n15281) );
  XNOR U23644 ( .A(n24076), .B(n24077), .Z(n20800) );
  AND U23645 ( .A(n23531), .B(n21147), .Z(n24076) );
  XOR U23646 ( .A(round_reg[1323]), .B(n24078), .Z(n21147) );
  IV U23647 ( .A(n20876), .Z(n17237) );
  XOR U23648 ( .A(n18848), .B(n22452), .Z(n20876) );
  XNOR U23649 ( .A(n24079), .B(n24080), .Z(n22452) );
  XOR U23650 ( .A(n13891), .B(n17666), .Z(n24080) );
  XOR U23651 ( .A(n24081), .B(n23539), .Z(n17666) );
  ANDN U23652 ( .B(n20878), .A(n20879), .Z(n24081) );
  XOR U23653 ( .A(round_reg[56]), .B(n24082), .Z(n20879) );
  XNOR U23654 ( .A(n24083), .B(n21157), .Z(n13891) );
  AND U23655 ( .A(n21656), .B(n21655), .Z(n24083) );
  XNOR U23656 ( .A(round_reg[308]), .B(n24084), .Z(n21656) );
  XOR U23657 ( .A(n18844), .B(n24085), .Z(n24079) );
  XOR U23658 ( .A(n17931), .B(n24086), .Z(n24085) );
  XNOR U23659 ( .A(n24087), .B(n21149), .Z(n17931) );
  ANDN U23660 ( .B(n24077), .A(n23531), .Z(n24087) );
  XOR U23661 ( .A(round_reg[78]), .B(n23595), .Z(n23531) );
  XNOR U23662 ( .A(n24088), .B(n21153), .Z(n18844) );
  AND U23663 ( .A(n23533), .B(n22170), .Z(n24088) );
  IV U23664 ( .A(n22171), .Z(n23533) );
  XOR U23665 ( .A(round_reg[196]), .B(n24089), .Z(n22171) );
  XOR U23666 ( .A(n24090), .B(n24091), .Z(n18848) );
  XOR U23667 ( .A(n18188), .B(n18724), .Z(n24091) );
  XOR U23668 ( .A(n24092), .B(n21171), .Z(n18724) );
  NOR U23669 ( .A(n23519), .B(n23937), .Z(n24092) );
  XOR U23670 ( .A(round_reg[1038]), .B(n23595), .Z(n23519) );
  XNOR U23671 ( .A(n24093), .B(n21179), .Z(n18188) );
  AND U23672 ( .A(n23514), .B(n23929), .Z(n24093) );
  XNOR U23673 ( .A(round_reg[1009]), .B(n22267), .Z(n23514) );
  XOR U23674 ( .A(n21789), .B(n24094), .Z(n24090) );
  XOR U23675 ( .A(n19292), .B(n16457), .Z(n24094) );
  XNOR U23676 ( .A(n24095), .B(n21176), .Z(n16457) );
  ANDN U23677 ( .B(n23522), .A(n23935), .Z(n24095) );
  XNOR U23678 ( .A(round_reg[1249]), .B(n23745), .Z(n23522) );
  XNOR U23679 ( .A(n24096), .B(n21166), .Z(n19292) );
  ANDN U23680 ( .B(n23939), .A(n23517), .Z(n24096) );
  XOR U23681 ( .A(round_reg[1151]), .B(n23603), .Z(n23517) );
  XNOR U23682 ( .A(n24097), .B(n21162), .Z(n21789) );
  ANDN U23683 ( .B(n23924), .A(n23932), .Z(n24097) );
  XNOR U23684 ( .A(round_reg[1177]), .B(n24098), .Z(n23924) );
  XOR U23685 ( .A(n23819), .B(n17928), .Z(n16517) );
  XNOR U23686 ( .A(n24099), .B(n24100), .Z(n23191) );
  XOR U23687 ( .A(n16667), .B(n14945), .Z(n24100) );
  XNOR U23688 ( .A(n24101), .B(n21578), .Z(n14945) );
  ANDN U23689 ( .B(n22844), .A(n21577), .Z(n24101) );
  XOR U23690 ( .A(n24102), .B(n20889), .Z(n16667) );
  ANDN U23691 ( .B(n22852), .A(n20888), .Z(n24102) );
  XOR U23692 ( .A(n18973), .B(n24103), .Z(n24099) );
  XOR U23693 ( .A(n19742), .B(n17717), .Z(n24103) );
  XOR U23694 ( .A(n24104), .B(n20899), .Z(n17717) );
  ANDN U23695 ( .B(n22855), .A(n20898), .Z(n24104) );
  XOR U23696 ( .A(n24105), .B(n20893), .Z(n19742) );
  XOR U23697 ( .A(n24106), .B(n20903), .Z(n18973) );
  ANDN U23698 ( .B(n24107), .A(n20902), .Z(n24106) );
  XNOR U23699 ( .A(n24109), .B(n22907), .Z(n23819) );
  AND U23700 ( .A(n22860), .B(n24110), .Z(n24109) );
  XOR U23701 ( .A(n15236), .B(n24111), .Z(n23997) );
  XOR U23702 ( .A(n9559), .B(n11134), .Z(n24111) );
  XNOR U23703 ( .A(n24112), .B(n15277), .Z(n11134) );
  XNOR U23704 ( .A(n23652), .B(n16938), .Z(n15277) );
  XNOR U23705 ( .A(n19015), .B(n22630), .Z(n16938) );
  XNOR U23706 ( .A(n24113), .B(n24114), .Z(n22630) );
  XNOR U23707 ( .A(n18386), .B(n19929), .Z(n24114) );
  XOR U23708 ( .A(n24115), .B(n21990), .Z(n19929) );
  XNOR U23709 ( .A(round_reg[10]), .B(n24116), .Z(n21990) );
  ANDN U23710 ( .B(n23648), .A(n23649), .Z(n24115) );
  XOR U23711 ( .A(round_reg[1560]), .B(n23406), .Z(n23648) );
  XOR U23712 ( .A(n24117), .B(n22682), .Z(n18386) );
  XNOR U23713 ( .A(round_reg[214]), .B(n22691), .Z(n22682) );
  AND U23714 ( .A(n23655), .B(n23654), .Z(n24117) );
  XOR U23715 ( .A(round_reg[1434]), .B(n23149), .Z(n23654) );
  XOR U23716 ( .A(n21947), .B(n24118), .Z(n24113) );
  XOR U23717 ( .A(n15648), .B(n19259), .Z(n24118) );
  XNOR U23718 ( .A(n24119), .B(n21986), .Z(n19259) );
  XOR U23719 ( .A(round_reg[155]), .B(n23411), .Z(n21986) );
  NOR U23720 ( .A(n23646), .B(n21985), .Z(n24119) );
  XNOR U23721 ( .A(round_reg[1404]), .B(n24026), .Z(n21985) );
  XOR U23722 ( .A(n24120), .B(n21976), .Z(n15648) );
  XNOR U23723 ( .A(round_reg[96]), .B(n22268), .Z(n21976) );
  XOR U23724 ( .A(round_reg[1341]), .B(n24121), .Z(n21975) );
  XOR U23725 ( .A(n24122), .B(n21980), .Z(n21947) );
  XNOR U23726 ( .A(round_reg[262]), .B(n23607), .Z(n21980) );
  ANDN U23727 ( .B(n24123), .A(n24124), .Z(n24122) );
  XOR U23728 ( .A(n24125), .B(n24126), .Z(n19015) );
  XOR U23729 ( .A(n20827), .B(n18171), .Z(n24126) );
  XOR U23730 ( .A(n24127), .B(n21965), .Z(n18171) );
  XOR U23731 ( .A(round_reg[1056]), .B(n22268), .Z(n21965) );
  ANDN U23732 ( .B(n23663), .A(n22053), .Z(n24127) );
  XOR U23733 ( .A(round_reg[622]), .B(n24128), .Z(n22053) );
  IV U23734 ( .A(n21966), .Z(n23663) );
  XNOR U23735 ( .A(round_reg[688]), .B(n23445), .Z(n21966) );
  XOR U23736 ( .A(n24129), .B(n21970), .Z(n20827) );
  XNOR U23737 ( .A(round_reg[1105]), .B(n22790), .Z(n21970) );
  XOR U23738 ( .A(round_reg[335]), .B(n23606), .Z(n22046) );
  XOR U23739 ( .A(round_reg[766]), .B(n23561), .Z(n21969) );
  XOR U23740 ( .A(n18557), .B(n24130), .Z(n24125) );
  XNOR U23741 ( .A(n18795), .B(n18517), .Z(n24130) );
  XOR U23742 ( .A(n24131), .B(n21957), .Z(n18517) );
  XNOR U23743 ( .A(round_reg[1195]), .B(n22112), .Z(n21957) );
  NOR U23744 ( .A(n21956), .B(n22056), .Z(n24131) );
  XOR U23745 ( .A(round_reg[386]), .B(n24132), .Z(n22056) );
  XNOR U23746 ( .A(round_reg[812]), .B(n23598), .Z(n21956) );
  XNOR U23747 ( .A(n24133), .B(n21962), .Z(n18795) );
  XNOR U23748 ( .A(round_reg[1267]), .B(n21312), .Z(n21962) );
  NOR U23749 ( .A(n21961), .B(n22043), .Z(n24133) );
  XOR U23750 ( .A(round_reg[456]), .B(n24134), .Z(n22043) );
  XNOR U23751 ( .A(round_reg[845]), .B(n23502), .Z(n21961) );
  XNOR U23752 ( .A(n24135), .B(n21953), .Z(n18557) );
  XOR U23753 ( .A(round_reg[963]), .B(n24136), .Z(n21953) );
  NOR U23754 ( .A(n21952), .B(n22050), .Z(n24135) );
  XOR U23755 ( .A(round_reg[554]), .B(n23920), .Z(n22050) );
  XNOR U23756 ( .A(round_reg[916]), .B(n24137), .Z(n21952) );
  XNOR U23757 ( .A(n24138), .B(n21979), .Z(n23652) );
  IV U23758 ( .A(n24123), .Z(n21979) );
  XOR U23759 ( .A(round_reg[1495]), .B(n24139), .Z(n24123) );
  ANDN U23760 ( .B(n24124), .A(n24046), .Z(n24138) );
  ANDN U23761 ( .B(n15276), .A(n16521), .Z(n24112) );
  XOR U23762 ( .A(n24140), .B(n18355), .Z(n16521) );
  XOR U23763 ( .A(n20218), .B(n18102), .Z(n15276) );
  XNOR U23764 ( .A(n23982), .B(n19072), .Z(n18102) );
  XNOR U23765 ( .A(n24141), .B(n24142), .Z(n19072) );
  XNOR U23766 ( .A(n17805), .B(n17513), .Z(n24142) );
  XOR U23767 ( .A(n24143), .B(n22212), .Z(n17513) );
  ANDN U23768 ( .B(n20210), .A(n20211), .Z(n24143) );
  XOR U23769 ( .A(round_reg[939]), .B(n22375), .Z(n20211) );
  XOR U23770 ( .A(n24144), .B(n22199), .Z(n17805) );
  NOR U23771 ( .A(n20214), .B(n20215), .Z(n24144) );
  XOR U23772 ( .A(round_reg[771]), .B(n22757), .Z(n20215) );
  XOR U23773 ( .A(n13990), .B(n24145), .Z(n24141) );
  XOR U23774 ( .A(n16832), .B(n18854), .Z(n24145) );
  XNOR U23775 ( .A(n24146), .B(n22209), .Z(n18854) );
  IV U23776 ( .A(n24147), .Z(n22209) );
  NOR U23777 ( .A(n24148), .B(n21208), .Z(n24146) );
  XOR U23778 ( .A(n24149), .B(n22207), .Z(n16832) );
  ANDN U23779 ( .B(n20220), .A(n20221), .Z(n24149) );
  XOR U23780 ( .A(round_reg[647]), .B(n23492), .Z(n20221) );
  XNOR U23781 ( .A(n24150), .B(n22202), .Z(n13990) );
  NOR U23782 ( .A(n20226), .B(n20224), .Z(n24150) );
  XOR U23783 ( .A(round_reg[725]), .B(n23409), .Z(n20226) );
  XOR U23784 ( .A(n24151), .B(n24152), .Z(n23982) );
  XNOR U23785 ( .A(n18152), .B(n16955), .Z(n24152) );
  XOR U23786 ( .A(n24153), .B(n20071), .Z(n16955) );
  XNOR U23787 ( .A(round_reg[646]), .B(n23738), .Z(n20071) );
  ANDN U23788 ( .B(n19816), .A(n19817), .Z(n24153) );
  XOR U23789 ( .A(round_reg[580]), .B(n22983), .Z(n19816) );
  XOR U23790 ( .A(n24154), .B(n19951), .Z(n18152) );
  XNOR U23791 ( .A(round_reg[724]), .B(n24155), .Z(n19951) );
  ANDN U23792 ( .B(n19950), .A(n21188), .Z(n24154) );
  XNOR U23793 ( .A(round_reg[283]), .B(n24156), .Z(n21188) );
  XOR U23794 ( .A(round_reg[357]), .B(n24157), .Z(n19950) );
  XOR U23795 ( .A(n19933), .B(n24158), .Z(n24151) );
  XNOR U23796 ( .A(n19157), .B(n18223), .Z(n24158) );
  XNOR U23797 ( .A(n24159), .B(n19947), .Z(n18223) );
  XNOR U23798 ( .A(round_reg[867]), .B(n23280), .Z(n19947) );
  ANDN U23799 ( .B(n19808), .A(n19806), .Z(n24159) );
  XNOR U23800 ( .A(round_reg[478]), .B(n21923), .Z(n19806) );
  XOR U23801 ( .A(n24160), .B(n19942), .Z(n19157) );
  XNOR U23802 ( .A(round_reg[770]), .B(n24161), .Z(n19942) );
  XNOR U23803 ( .A(round_reg[408]), .B(n23275), .Z(n19802) );
  XNOR U23804 ( .A(round_reg[31]), .B(n23325), .Z(n19804) );
  XOR U23805 ( .A(n24162), .B(n19939), .Z(n19933) );
  XNOR U23806 ( .A(round_reg[938]), .B(n23602), .Z(n19939) );
  AND U23807 ( .A(n19814), .B(n19812), .Z(n24162) );
  XOR U23808 ( .A(round_reg[512]), .B(n24163), .Z(n19812) );
  XNOR U23809 ( .A(round_reg[176]), .B(n23963), .Z(n19814) );
  XNOR U23810 ( .A(n24164), .B(n24148), .Z(n20218) );
  AND U23811 ( .A(n21209), .B(n21208), .Z(n24164) );
  XOR U23812 ( .A(round_reg[868]), .B(n23293), .Z(n21208) );
  XNOR U23813 ( .A(round_reg[479]), .B(n24165), .Z(n21209) );
  XOR U23814 ( .A(n24166), .B(n15268), .Z(n9559) );
  XNOR U23815 ( .A(n22569), .B(n17978), .Z(n15268) );
  IV U23816 ( .A(n18879), .Z(n17978) );
  XOR U23817 ( .A(n20190), .B(n20237), .Z(n18879) );
  XOR U23818 ( .A(n24167), .B(n24168), .Z(n20237) );
  XNOR U23819 ( .A(n17866), .B(n19501), .Z(n24168) );
  XNOR U23820 ( .A(n24169), .B(n24170), .Z(n19501) );
  ANDN U23821 ( .B(n22556), .A(n22557), .Z(n24169) );
  XOR U23822 ( .A(round_reg[1245]), .B(n24171), .Z(n22557) );
  XOR U23823 ( .A(n24172), .B(n24173), .Z(n17866) );
  ANDN U23824 ( .B(n22545), .A(n22546), .Z(n24172) );
  XOR U23825 ( .A(round_reg[1005]), .B(n22374), .Z(n22546) );
  XOR U23826 ( .A(n24174), .B(n24175), .Z(n24167) );
  XOR U23827 ( .A(n19229), .B(n17552), .Z(n24175) );
  XOR U23828 ( .A(n24176), .B(n24177), .Z(n17552) );
  ANDN U23829 ( .B(n22564), .A(n22565), .Z(n24176) );
  XOR U23830 ( .A(round_reg[1147]), .B(n23250), .Z(n22565) );
  XOR U23831 ( .A(n24178), .B(n24179), .Z(n19229) );
  ANDN U23832 ( .B(n22560), .A(n22561), .Z(n24178) );
  XOR U23833 ( .A(round_reg[1034]), .B(n22839), .Z(n22561) );
  XNOR U23834 ( .A(n24180), .B(n24181), .Z(n20190) );
  XOR U23835 ( .A(n18939), .B(n20322), .Z(n24181) );
  XOR U23836 ( .A(n24182), .B(n22465), .Z(n20322) );
  ANDN U23837 ( .B(n22576), .A(n22577), .Z(n24182) );
  XOR U23838 ( .A(round_reg[429]), .B(n24183), .Z(n22576) );
  XNOR U23839 ( .A(n24184), .B(n24185), .Z(n18939) );
  ANDN U23840 ( .B(n24186), .A(n24187), .Z(n24184) );
  XOR U23841 ( .A(n19598), .B(n24188), .Z(n24180) );
  XOR U23842 ( .A(n22455), .B(n18457), .Z(n24188) );
  XNOR U23843 ( .A(n24189), .B(n22475), .Z(n18457) );
  ANDN U23844 ( .B(n22476), .A(n22808), .Z(n24189) );
  XOR U23845 ( .A(round_reg[601]), .B(n23918), .Z(n22476) );
  XNOR U23846 ( .A(n24190), .B(n22471), .Z(n22455) );
  ANDN U23847 ( .B(n22472), .A(n22571), .Z(n24190) );
  XOR U23848 ( .A(round_reg[499]), .B(n23621), .Z(n22472) );
  XNOR U23849 ( .A(n24191), .B(n22461), .Z(n19598) );
  ANDN U23850 ( .B(n22462), .A(n22580), .Z(n24191) );
  XOR U23851 ( .A(round_reg[533]), .B(n22984), .Z(n22462) );
  XNOR U23852 ( .A(n24192), .B(n24186), .Z(n22569) );
  ANDN U23853 ( .B(n24187), .A(n24193), .Z(n24192) );
  ANDN U23854 ( .B(n18089), .A(n15267), .Z(n24166) );
  XOR U23855 ( .A(n20438), .B(n16896), .Z(n15267) );
  XOR U23856 ( .A(n24194), .B(n22356), .Z(n16896) );
  XOR U23857 ( .A(n24195), .B(n24196), .Z(n22356) );
  XNOR U23858 ( .A(n24197), .B(n17565), .Z(n24196) );
  XOR U23859 ( .A(n24198), .B(n22781), .Z(n17565) );
  ANDN U23860 ( .B(n24199), .A(n21840), .Z(n24198) );
  XNOR U23861 ( .A(n19440), .B(n24200), .Z(n24195) );
  XNOR U23862 ( .A(n19297), .B(n20086), .Z(n24200) );
  XNOR U23863 ( .A(n24201), .B(n22779), .Z(n20086) );
  AND U23864 ( .A(n20429), .B(n21834), .Z(n24201) );
  IV U23865 ( .A(n20430), .Z(n21834) );
  XOR U23866 ( .A(round_reg[1555]), .B(n24202), .Z(n20430) );
  XNOR U23867 ( .A(n24203), .B(n22776), .Z(n19297) );
  AND U23868 ( .A(n23046), .B(n21847), .Z(n24203) );
  IV U23869 ( .A(n23047), .Z(n21847) );
  XOR U23870 ( .A(round_reg[1490]), .B(n22645), .Z(n23047) );
  XNOR U23871 ( .A(n24204), .B(n22784), .Z(n19440) );
  AND U23872 ( .A(n20440), .B(n20442), .Z(n24204) );
  XOR U23873 ( .A(round_reg[1399]), .B(n24205), .Z(n20442) );
  XNOR U23874 ( .A(n24206), .B(n24199), .Z(n20438) );
  ANDN U23875 ( .B(n21840), .A(n21841), .Z(n24206) );
  XNOR U23876 ( .A(round_reg[1263]), .B(n24207), .Z(n21841) );
  XNOR U23877 ( .A(round_reg[1336]), .B(n24208), .Z(n21840) );
  XNOR U23878 ( .A(n24209), .B(n17792), .Z(n18089) );
  XNOR U23879 ( .A(n24210), .B(n15272), .Z(n15236) );
  XOR U23880 ( .A(n20672), .B(n17031), .Z(n15272) );
  XNOR U23881 ( .A(n21477), .B(n21406), .Z(n17031) );
  XNOR U23882 ( .A(n24211), .B(n24212), .Z(n21406) );
  XOR U23883 ( .A(n15602), .B(n17912), .Z(n24212) );
  XNOR U23884 ( .A(n24213), .B(n19281), .Z(n17912) );
  XNOR U23885 ( .A(round_reg[909]), .B(n24214), .Z(n19281) );
  NOR U23886 ( .A(n21432), .B(n21431), .Z(n24213) );
  XNOR U23887 ( .A(round_reg[547]), .B(n23280), .Z(n21431) );
  XOR U23888 ( .A(round_reg[147]), .B(n22508), .Z(n21432) );
  XNOR U23889 ( .A(n24215), .B(n22584), .Z(n15602) );
  XOR U23890 ( .A(round_reg[805]), .B(n23919), .Z(n22584) );
  ANDN U23891 ( .B(n20753), .A(n20755), .Z(n24215) );
  XOR U23892 ( .A(round_reg[2]), .B(n22442), .Z(n20755) );
  XOR U23893 ( .A(round_reg[443]), .B(n22369), .Z(n20753) );
  XOR U23894 ( .A(n17327), .B(n24216), .Z(n24211) );
  XOR U23895 ( .A(n16444), .B(n21661), .Z(n24216) );
  XOR U23896 ( .A(n24217), .B(n23299), .Z(n21661) );
  IV U23897 ( .A(n23033), .Z(n23299) );
  XOR U23898 ( .A(round_reg[838]), .B(n24218), .Z(n23033) );
  AND U23899 ( .A(n20743), .B(n23287), .Z(n24217) );
  XNOR U23900 ( .A(round_reg[88]), .B(n23275), .Z(n23287) );
  XNOR U23901 ( .A(round_reg[449]), .B(n24219), .Z(n20743) );
  XNOR U23902 ( .A(n24220), .B(n20985), .Z(n16444) );
  XOR U23903 ( .A(round_reg[681]), .B(n24221), .Z(n20985) );
  ANDN U23904 ( .B(n20747), .A(n20748), .Z(n24220) );
  XOR U23905 ( .A(round_reg[206]), .B(n22221), .Z(n20748) );
  XOR U23906 ( .A(round_reg[615]), .B(n23260), .Z(n20747) );
  XOR U23907 ( .A(n24222), .B(n19274), .Z(n17327) );
  XNOR U23908 ( .A(round_reg[759]), .B(n24223), .Z(n19274) );
  ANDN U23909 ( .B(n20757), .A(n20758), .Z(n24222) );
  XNOR U23910 ( .A(round_reg[318]), .B(n23877), .Z(n20758) );
  XNOR U23911 ( .A(round_reg[328]), .B(n22977), .Z(n20757) );
  XOR U23912 ( .A(n24224), .B(n24225), .Z(n21477) );
  XNOR U23913 ( .A(n18681), .B(n17406), .Z(n24225) );
  XOR U23914 ( .A(n24226), .B(n22602), .Z(n17406) );
  XNOR U23915 ( .A(round_reg[1427]), .B(n22508), .Z(n22602) );
  NOR U23916 ( .A(n20675), .B(n20674), .Z(n24226) );
  XOR U23917 ( .A(round_reg[1050]), .B(n24227), .Z(n20674) );
  XOR U23918 ( .A(n24228), .B(n22610), .Z(n18681) );
  XNOR U23919 ( .A(round_reg[1488]), .B(n24229), .Z(n22610) );
  NOR U23920 ( .A(n24230), .B(n23042), .Z(n24228) );
  XOR U23921 ( .A(n18965), .B(n24231), .Z(n24224) );
  XOR U23922 ( .A(n23023), .B(n17541), .Z(n24231) );
  XOR U23923 ( .A(n24232), .B(n22606), .Z(n17541) );
  XNOR U23924 ( .A(round_reg[1553]), .B(n22362), .Z(n22606) );
  NOR U23925 ( .A(n20681), .B(n20680), .Z(n24232) );
  XOR U23926 ( .A(round_reg[1189]), .B(n24233), .Z(n20680) );
  XOR U23927 ( .A(n24234), .B(n22599), .Z(n23023) );
  XNOR U23928 ( .A(round_reg[1334]), .B(n23879), .Z(n22599) );
  AND U23929 ( .A(n22236), .B(n23037), .Z(n24234) );
  XOR U23930 ( .A(round_reg[1261]), .B(n21193), .Z(n23037) );
  XOR U23931 ( .A(n24235), .B(n22614), .Z(n18965) );
  IV U23932 ( .A(n23039), .Z(n22614) );
  XOR U23933 ( .A(round_reg[1397]), .B(n23993), .Z(n23039) );
  ANDN U23934 ( .B(n20686), .A(n20684), .Z(n24235) );
  XOR U23935 ( .A(round_reg[1021]), .B(n24121), .Z(n20684) );
  XNOR U23936 ( .A(n24236), .B(n23042), .Z(n20672) );
  XOR U23937 ( .A(round_reg[1099]), .B(n24237), .Z(n23042) );
  AND U23938 ( .A(n22609), .B(n24230), .Z(n24236) );
  AND U23939 ( .A(n16527), .B(n18126), .Z(n24210) );
  XOR U23940 ( .A(n22850), .B(n17509), .Z(n18126) );
  XNOR U23941 ( .A(n24238), .B(n24239), .Z(n21709) );
  XOR U23942 ( .A(n18822), .B(n15643), .Z(n24239) );
  XNOR U23943 ( .A(n24240), .B(n20662), .Z(n15643) );
  XOR U23944 ( .A(round_reg[508]), .B(n23323), .Z(n20662) );
  ANDN U23945 ( .B(n23204), .A(n21569), .Z(n24240) );
  XNOR U23946 ( .A(n24241), .B(n20649), .Z(n18822) );
  XNOR U23947 ( .A(round_reg[610]), .B(n24019), .Z(n20649) );
  ANDN U23948 ( .B(n23202), .A(n21571), .Z(n24241) );
  XOR U23949 ( .A(n19025), .B(n24242), .Z(n24238) );
  XOR U23950 ( .A(n17379), .B(n17600), .Z(n24242) );
  XOR U23951 ( .A(n24243), .B(n20657), .Z(n17600) );
  XNOR U23952 ( .A(round_reg[438]), .B(n21195), .Z(n20657) );
  ANDN U23953 ( .B(n23195), .A(n24244), .Z(n24243) );
  XNOR U23954 ( .A(n24245), .B(n20652), .Z(n17379) );
  XOR U23955 ( .A(round_reg[323]), .B(n24136), .Z(n20652) );
  AND U23956 ( .A(n21573), .B(n23198), .Z(n24245) );
  XNOR U23957 ( .A(n24246), .B(n20666), .Z(n19025) );
  XOR U23958 ( .A(round_reg[542]), .B(n22751), .Z(n20666) );
  AND U23959 ( .A(n21566), .B(n23207), .Z(n24246) );
  XOR U23960 ( .A(n24247), .B(n24248), .Z(n20610) );
  XNOR U23961 ( .A(n17920), .B(n16070), .Z(n24248) );
  XOR U23962 ( .A(n24249), .B(n20892), .Z(n16070) );
  XNOR U23963 ( .A(round_reg[1045]), .B(n23409), .Z(n20892) );
  ANDN U23964 ( .B(n22848), .A(n22847), .Z(n24249) );
  XNOR U23965 ( .A(round_reg[677]), .B(n24157), .Z(n22847) );
  XOR U23966 ( .A(n24250), .B(n20898), .Z(n17920) );
  XNOR U23967 ( .A(round_reg[1094]), .B(n24251), .Z(n20898) );
  ANDN U23968 ( .B(n22856), .A(n22855), .Z(n24250) );
  XOR U23969 ( .A(round_reg[755]), .B(n23914), .Z(n22855) );
  IV U23970 ( .A(n23475), .Z(n23914) );
  XOR U23971 ( .A(n18426), .B(n24252), .Z(n24247) );
  XOR U23972 ( .A(n23190), .B(n16026), .Z(n24252) );
  XOR U23973 ( .A(n24253), .B(n20888), .Z(n16026) );
  XNOR U23974 ( .A(round_reg[1184]), .B(n24254), .Z(n20888) );
  ANDN U23975 ( .B(n22853), .A(n22852), .Z(n24253) );
  XOR U23976 ( .A(round_reg[801]), .B(n24255), .Z(n22852) );
  XOR U23977 ( .A(n24256), .B(n20902), .Z(n23190) );
  XNOR U23978 ( .A(round_reg[1256]), .B(n24257), .Z(n20902) );
  ANDN U23979 ( .B(n24258), .A(n24107), .Z(n24256) );
  XOR U23980 ( .A(n24259), .B(n21577), .Z(n18426) );
  XNOR U23981 ( .A(round_reg[1016]), .B(n24082), .Z(n21577) );
  ANDN U23982 ( .B(n22845), .A(n22844), .Z(n24259) );
  XNOR U23983 ( .A(round_reg[905]), .B(n21185), .Z(n22844) );
  XNOR U23984 ( .A(n24260), .B(n24107), .Z(n22850) );
  XOR U23985 ( .A(round_reg[834]), .B(n24261), .Z(n24107) );
  ANDN U23986 ( .B(n20901), .A(n24258), .Z(n24260) );
  XNOR U23987 ( .A(n17275), .B(n20972), .Z(n16527) );
  XOR U23988 ( .A(n24262), .B(n21546), .Z(n20972) );
  NOR U23989 ( .A(n24263), .B(n21904), .Z(n24262) );
  XOR U23990 ( .A(n24264), .B(n22586), .Z(n17275) );
  XOR U23991 ( .A(n24265), .B(n24266), .Z(n22586) );
  XNOR U23992 ( .A(n18339), .B(n16050), .Z(n24266) );
  XNOR U23993 ( .A(n24267), .B(n21550), .Z(n16050) );
  XOR U23994 ( .A(round_reg[714]), .B(n24268), .Z(n21550) );
  ANDN U23995 ( .B(n20974), .A(n20975), .Z(n24267) );
  XOR U23996 ( .A(round_reg[347]), .B(n23386), .Z(n20974) );
  XNOR U23997 ( .A(n24269), .B(n21554), .Z(n18339) );
  AND U23998 ( .A(n20970), .B(n20968), .Z(n24269) );
  XOR U23999 ( .A(round_reg[468]), .B(n23732), .Z(n20968) );
  XNOR U24000 ( .A(n20764), .B(n24270), .Z(n24265) );
  XOR U24001 ( .A(n21529), .B(n16929), .Z(n24270) );
  XOR U24002 ( .A(n24271), .B(n21557), .Z(n16929) );
  IV U24003 ( .A(n21899), .Z(n21557) );
  XNOR U24004 ( .A(round_reg[928]), .B(n24272), .Z(n21899) );
  AND U24005 ( .A(n20978), .B(n24273), .Z(n24271) );
  XOR U24006 ( .A(round_reg[566]), .B(n24274), .Z(n20978) );
  XNOR U24007 ( .A(n24275), .B(n21547), .Z(n21529) );
  XOR U24008 ( .A(round_reg[700]), .B(n23290), .Z(n21547) );
  XNOR U24009 ( .A(round_reg[634]), .B(n23318), .Z(n21546) );
  XNOR U24010 ( .A(n24276), .B(n21560), .Z(n20764) );
  XNOR U24011 ( .A(round_reg[824]), .B(n22642), .Z(n21560) );
  ANDN U24012 ( .B(n21561), .A(n21801), .Z(n24276) );
  XOR U24013 ( .A(round_reg[398]), .B(n23595), .Z(n21561) );
  XOR U24014 ( .A(n24277), .B(n24278), .Z(n14430) );
  XOR U24015 ( .A(n12156), .B(n10132), .Z(n24278) );
  XOR U24016 ( .A(n24279), .B(n14578), .Z(n10132) );
  XNOR U24017 ( .A(n22250), .B(n17951), .Z(n14578) );
  XNOR U24018 ( .A(n24280), .B(n24281), .Z(n19327) );
  XNOR U24019 ( .A(n17727), .B(n16977), .Z(n24281) );
  XOR U24020 ( .A(n24282), .B(n23970), .Z(n16977) );
  ANDN U24021 ( .B(n23969), .A(n23178), .Z(n24282) );
  XOR U24022 ( .A(n24283), .B(n23981), .Z(n17727) );
  ANDN U24023 ( .B(n22242), .A(n22243), .Z(n24283) );
  XOR U24024 ( .A(round_reg[72]), .B(n24284), .Z(n22243) );
  XOR U24025 ( .A(round_reg[497]), .B(n24285), .Z(n22242) );
  XOR U24026 ( .A(n15838), .B(n24286), .Z(n24280) );
  XOR U24027 ( .A(n16417), .B(n23953), .Z(n24286) );
  XNOR U24028 ( .A(n24287), .B(n23977), .Z(n23953) );
  AND U24029 ( .A(n22258), .B(n23978), .Z(n24287) );
  XOR U24030 ( .A(round_reg[531]), .B(n24288), .Z(n23978) );
  XNOR U24031 ( .A(round_reg[131]), .B(n22757), .Z(n22258) );
  XOR U24032 ( .A(n24289), .B(n23972), .Z(n16417) );
  ANDN U24033 ( .B(n22246), .A(n22247), .Z(n24289) );
  XOR U24034 ( .A(round_reg[302]), .B(n24128), .Z(n22247) );
  XOR U24035 ( .A(round_reg[376]), .B(n24082), .Z(n22246) );
  XNOR U24036 ( .A(n24290), .B(n23975), .Z(n15838) );
  ANDN U24037 ( .B(n22252), .A(n22253), .Z(n24290) );
  XOR U24038 ( .A(round_reg[254]), .B(n23588), .Z(n22253) );
  XOR U24039 ( .A(round_reg[599]), .B(n22687), .Z(n22252) );
  XOR U24040 ( .A(n24291), .B(n24292), .Z(n22504) );
  XNOR U24041 ( .A(n16776), .B(n19635), .Z(n24292) );
  XOR U24042 ( .A(n24293), .B(n20602), .Z(n19635) );
  AND U24043 ( .A(n20365), .B(n20363), .Z(n24293) );
  XOR U24044 ( .A(round_reg[1316]), .B(n23201), .Z(n20363) );
  XNOR U24045 ( .A(round_reg[1243]), .B(n24294), .Z(n20365) );
  XNOR U24046 ( .A(n24295), .B(n20594), .Z(n16776) );
  XOR U24047 ( .A(round_reg[301]), .B(n21193), .Z(n20594) );
  XOR U24048 ( .A(round_reg[1145]), .B(n24296), .Z(n20368) );
  XOR U24049 ( .A(round_reg[1534]), .B(n23588), .Z(n20367) );
  XOR U24050 ( .A(n17371), .B(n24297), .Z(n24291) );
  XOR U24051 ( .A(n16020), .B(n18107), .Z(n24297) );
  XNOR U24052 ( .A(n24298), .B(n20600), .Z(n18107) );
  XOR U24053 ( .A(round_reg[49]), .B(n22267), .Z(n20600) );
  AND U24054 ( .A(n21874), .B(n21870), .Z(n24298) );
  IV U24055 ( .A(n23957), .Z(n21870) );
  XOR U24056 ( .A(round_reg[1599]), .B(n24299), .Z(n23957) );
  XNOR U24057 ( .A(round_reg[1171]), .B(n24288), .Z(n21874) );
  XNOR U24058 ( .A(n24300), .B(n20591), .Z(n16020) );
  XOR U24059 ( .A(round_reg[253]), .B(n23387), .Z(n20591) );
  AND U24060 ( .A(n22520), .B(n22519), .Z(n24300) );
  XOR U24061 ( .A(round_reg[1409]), .B(n23886), .Z(n22519) );
  XNOR U24062 ( .A(round_reg[1032]), .B(n24284), .Z(n22520) );
  XNOR U24063 ( .A(n24301), .B(n23889), .Z(n17371) );
  XOR U24064 ( .A(round_reg[130]), .B(n24161), .Z(n23889) );
  AND U24065 ( .A(n20359), .B(n20357), .Z(n24301) );
  XOR U24066 ( .A(round_reg[1379]), .B(n21920), .Z(n20357) );
  XNOR U24067 ( .A(round_reg[1003]), .B(n24302), .Z(n20359) );
  XNOR U24068 ( .A(n24303), .B(n23969), .Z(n22250) );
  XOR U24069 ( .A(round_reg[427]), .B(n23946), .Z(n23969) );
  ANDN U24070 ( .B(n23178), .A(n23179), .Z(n24303) );
  XOR U24071 ( .A(round_reg[50]), .B(n23781), .Z(n23178) );
  AND U24072 ( .A(n14579), .B(n16542), .Z(n24279) );
  XOR U24073 ( .A(n17234), .B(n24035), .Z(n16542) );
  XOR U24074 ( .A(n24304), .B(n23724), .Z(n24035) );
  ANDN U24075 ( .B(n21641), .A(n21642), .Z(n24304) );
  XNOR U24076 ( .A(round_reg[704]), .B(n24305), .Z(n21642) );
  XOR U24077 ( .A(n19670), .B(n19181), .Z(n17234) );
  XNOR U24078 ( .A(n24306), .B(n24307), .Z(n19181) );
  XNOR U24079 ( .A(n17577), .B(n20024), .Z(n24307) );
  XOR U24080 ( .A(n24308), .B(n23557), .Z(n20024) );
  XNOR U24081 ( .A(round_reg[11]), .B(n21754), .Z(n23557) );
  NOR U24082 ( .A(n23722), .B(n21647), .Z(n24308) );
  XOR U24083 ( .A(round_reg[1197]), .B(n24309), .Z(n21647) );
  XNOR U24084 ( .A(round_reg[1561]), .B(n23918), .Z(n23722) );
  XNOR U24085 ( .A(n24310), .B(n23546), .Z(n17577) );
  XOR U24086 ( .A(round_reg[215]), .B(n24139), .Z(n23546) );
  XOR U24087 ( .A(round_reg[1058]), .B(n23804), .Z(n24039) );
  XNOR U24088 ( .A(round_reg[1435]), .B(n23411), .Z(n23718) );
  XOR U24089 ( .A(n17788), .B(n24311), .Z(n24306) );
  XOR U24090 ( .A(n15654), .B(n20325), .Z(n24311) );
  XNOR U24091 ( .A(n24312), .B(n23548), .Z(n20325) );
  XOR U24092 ( .A(round_reg[263]), .B(n23916), .Z(n23548) );
  ANDN U24093 ( .B(n23724), .A(n21641), .Z(n24312) );
  XOR U24094 ( .A(round_reg[1107]), .B(n22508), .Z(n21641) );
  XOR U24095 ( .A(round_reg[1496]), .B(n24313), .Z(n23724) );
  XOR U24096 ( .A(n24314), .B(n23551), .Z(n15654) );
  XNOR U24097 ( .A(round_reg[97]), .B(n23780), .Z(n23551) );
  XOR U24098 ( .A(round_reg[1269]), .B(n23467), .Z(n21651) );
  XOR U24099 ( .A(round_reg[1342]), .B(n24315), .Z(n23716) );
  XOR U24100 ( .A(n24316), .B(n23554), .Z(n17788) );
  XNOR U24101 ( .A(round_reg[156]), .B(n23568), .Z(n23554) );
  ANDN U24102 ( .B(n23727), .A(n23675), .Z(n24316) );
  XOR U24103 ( .A(round_reg[965]), .B(n23895), .Z(n23675) );
  XNOR U24104 ( .A(round_reg[1405]), .B(n22764), .Z(n23727) );
  XOR U24105 ( .A(n24317), .B(n24318), .Z(n19670) );
  XNOR U24106 ( .A(n17077), .B(n17139), .Z(n24318) );
  XOR U24107 ( .A(n24319), .B(n23655), .Z(n17139) );
  XOR U24108 ( .A(round_reg[1057]), .B(n24320), .Z(n23655) );
  ANDN U24109 ( .B(n23656), .A(n22680), .Z(n24319) );
  XOR U24110 ( .A(round_reg[623]), .B(n21763), .Z(n22680) );
  XOR U24111 ( .A(round_reg[689]), .B(n22267), .Z(n23656) );
  XNOR U24112 ( .A(n24321), .B(n24124), .Z(n17077) );
  XOR U24113 ( .A(round_reg[1106]), .B(n23295), .Z(n24124) );
  ANDN U24114 ( .B(n24046), .A(n21978), .Z(n24321) );
  XOR U24115 ( .A(round_reg[336]), .B(n23915), .Z(n21978) );
  XOR U24116 ( .A(round_reg[767]), .B(n22371), .Z(n24046) );
  XOR U24117 ( .A(n18798), .B(n24322), .Z(n24317) );
  XOR U24118 ( .A(n23641), .B(n18183), .Z(n24322) );
  XNOR U24119 ( .A(n24323), .B(n23649), .Z(n18183) );
  XOR U24120 ( .A(round_reg[1196]), .B(n23726), .Z(n23649) );
  ANDN U24121 ( .B(n23650), .A(n21988), .Z(n24323) );
  XNOR U24122 ( .A(round_reg[387]), .B(n21747), .Z(n21988) );
  XOR U24123 ( .A(round_reg[813]), .B(n23413), .Z(n23650) );
  XNOR U24124 ( .A(n24324), .B(n23658), .Z(n23641) );
  XNOR U24125 ( .A(round_reg[1268]), .B(n24325), .Z(n23658) );
  ANDN U24126 ( .B(n23659), .A(n21974), .Z(n24324) );
  XOR U24127 ( .A(round_reg[457]), .B(n23283), .Z(n21974) );
  XOR U24128 ( .A(round_reg[846]), .B(n22221), .Z(n23659) );
  XNOR U24129 ( .A(n24326), .B(n23646), .Z(n18798) );
  XOR U24130 ( .A(round_reg[964]), .B(n23016), .Z(n23646) );
  NOR U24131 ( .A(n21984), .B(n23645), .Z(n24326) );
  XOR U24132 ( .A(round_reg[917]), .B(n24327), .Z(n23645) );
  XOR U24133 ( .A(round_reg[555]), .B(n22112), .Z(n21984) );
  XNOR U24134 ( .A(n24328), .B(n24329), .Z(n22112) );
  XNOR U24135 ( .A(n17402), .B(n20399), .Z(n14579) );
  XOR U24136 ( .A(n24330), .B(n24331), .Z(n20399) );
  ANDN U24137 ( .B(n22530), .A(n22528), .Z(n24330) );
  XOR U24138 ( .A(n23365), .B(n22453), .Z(n17402) );
  XNOR U24139 ( .A(n24332), .B(n24333), .Z(n22453) );
  XOR U24140 ( .A(n19481), .B(n18179), .Z(n24333) );
  XNOR U24141 ( .A(n24334), .B(n21944), .Z(n18179) );
  ANDN U24142 ( .B(n19650), .A(n19517), .Z(n24334) );
  XOR U24143 ( .A(round_reg[672]), .B(n21606), .Z(n19517) );
  XOR U24144 ( .A(round_reg[1040]), .B(n22445), .Z(n19650) );
  XNOR U24145 ( .A(n24335), .B(n21936), .Z(n19481) );
  XNOR U24146 ( .A(round_reg[1478]), .B(n24218), .Z(n21936) );
  AND U24147 ( .A(n21937), .B(n19512), .Z(n24335) );
  XNOR U24148 ( .A(round_reg[750]), .B(n22825), .Z(n19512) );
  XOR U24149 ( .A(round_reg[1089]), .B(n23886), .Z(n21937) );
  IV U24150 ( .A(n24219), .Z(n23886) );
  XNOR U24151 ( .A(n19146), .B(n24338), .Z(n24332) );
  XNOR U24152 ( .A(n20092), .B(n21320), .Z(n24338) );
  XOR U24153 ( .A(n21946), .B(n24339), .Z(n21320) );
  XOR U24154 ( .A(n24340), .B(n6870), .Z(n24339) );
  NAND U24155 ( .A(n4640), .B(n24341), .Z(n6870) );
  AND U24156 ( .A(n11363), .B(n6455), .Z(n4640) );
  ANDN U24157 ( .B(n19645), .A(n19508), .Z(n24340) );
  XOR U24158 ( .A(round_reg[796]), .B(n23568), .Z(n19508) );
  XOR U24159 ( .A(round_reg[1179]), .B(n24342), .Z(n19645) );
  XOR U24160 ( .A(round_reg[1543]), .B(n23916), .Z(n21946) );
  XNOR U24161 ( .A(n24343), .B(n23462), .Z(n20092) );
  IV U24162 ( .A(n21942), .Z(n23462) );
  XOR U24163 ( .A(round_reg[1324]), .B(n23785), .Z(n21942) );
  ANDN U24164 ( .B(n20014), .A(n19521), .Z(n24343) );
  XOR U24165 ( .A(round_reg[893]), .B(n23387), .Z(n19521) );
  XOR U24166 ( .A(n24344), .B(n24345), .Z(n23387) );
  XOR U24167 ( .A(round_reg[1251]), .B(n23256), .Z(n20014) );
  XNOR U24168 ( .A(n24346), .B(n23472), .Z(n19146) );
  IV U24169 ( .A(n21939), .Z(n23472) );
  XOR U24170 ( .A(round_reg[1387]), .B(n23946), .Z(n21939) );
  ANDN U24171 ( .B(n19973), .A(n19525), .Z(n24346) );
  XOR U24172 ( .A(round_reg[900]), .B(n22983), .Z(n19525) );
  XOR U24173 ( .A(round_reg[1011]), .B(n23504), .Z(n19973) );
  XOR U24174 ( .A(n24347), .B(n24348), .Z(n23365) );
  XOR U24175 ( .A(n16829), .B(n19712), .Z(n24348) );
  XNOR U24176 ( .A(n24349), .B(n24350), .Z(n19712) );
  ANDN U24177 ( .B(n20410), .A(n20412), .Z(n24349) );
  XOR U24178 ( .A(round_reg[1325]), .B(n22374), .Z(n20412) );
  XNOR U24179 ( .A(n24351), .B(n24352), .Z(n16829) );
  ANDN U24180 ( .B(n20414), .A(n20415), .Z(n24351) );
  XOR U24181 ( .A(round_reg[1418]), .B(n22108), .Z(n20415) );
  XNOR U24182 ( .A(n24353), .B(n24354), .Z(n22108) );
  XOR U24183 ( .A(n21931), .B(n24355), .Z(n24347) );
  XNOR U24184 ( .A(n20782), .B(n19399), .Z(n24355) );
  XNOR U24185 ( .A(n24356), .B(n24357), .Z(n19399) );
  ANDN U24186 ( .B(n20406), .A(n20407), .Z(n24356) );
  XNOR U24187 ( .A(round_reg[1544]), .B(n23986), .Z(n20407) );
  XNOR U24188 ( .A(n24358), .B(n24359), .Z(n20782) );
  ANDN U24189 ( .B(n20401), .A(n20402), .Z(n24358) );
  XNOR U24190 ( .A(round_reg[1479]), .B(n24006), .Z(n20402) );
  IV U24191 ( .A(n24360), .Z(n20401) );
  XNOR U24192 ( .A(n24361), .B(n24362), .Z(n21931) );
  AND U24193 ( .A(n22528), .B(n24363), .Z(n24361) );
  XNOR U24194 ( .A(round_reg[1388]), .B(n24364), .Z(n22528) );
  XNOR U24195 ( .A(n24365), .B(n14573), .Z(n12156) );
  XOR U24196 ( .A(n20314), .B(n19723), .Z(n14573) );
  XNOR U24197 ( .A(n24366), .B(n20452), .Z(n19723) );
  AND U24198 ( .A(n19474), .B(n24367), .Z(n24366) );
  XOR U24199 ( .A(round_reg[817]), .B(n24368), .Z(n19474) );
  XOR U24200 ( .A(n21034), .B(n23210), .Z(n20314) );
  XNOR U24201 ( .A(n24369), .B(n24370), .Z(n23210) );
  XNOR U24202 ( .A(n16933), .B(n20443), .Z(n24370) );
  XNOR U24203 ( .A(n24371), .B(n19476), .Z(n20443) );
  XOR U24204 ( .A(round_reg[14]), .B(n22115), .Z(n19476) );
  AND U24205 ( .A(n20452), .B(n21315), .Z(n24371) );
  IV U24206 ( .A(n24367), .Z(n21315) );
  XOR U24207 ( .A(round_reg[1200]), .B(n23618), .Z(n24367) );
  XNOR U24208 ( .A(round_reg[1564]), .B(n24372), .Z(n20452) );
  XNOR U24209 ( .A(n24373), .B(n19470), .Z(n16933) );
  XOR U24210 ( .A(round_reg[218]), .B(n23471), .Z(n19470) );
  AND U24211 ( .A(n19729), .B(n19730), .Z(n24373) );
  XOR U24212 ( .A(round_reg[1061]), .B(n24374), .Z(n19730) );
  XOR U24213 ( .A(round_reg[1438]), .B(n21923), .Z(n19729) );
  XOR U24214 ( .A(n14940), .B(n24375), .Z(n24369) );
  XOR U24215 ( .A(n17418), .B(n18569), .Z(n24375) );
  XNOR U24216 ( .A(n24376), .B(n20455), .Z(n18569) );
  XOR U24217 ( .A(round_reg[266]), .B(n24377), .Z(n20455) );
  AND U24218 ( .A(n21301), .B(n20456), .Z(n24376) );
  XOR U24219 ( .A(round_reg[1499]), .B(n24342), .Z(n20456) );
  XNOR U24220 ( .A(round_reg[1110]), .B(n24378), .Z(n21301) );
  XNOR U24221 ( .A(n24379), .B(n19480), .Z(n17418) );
  XOR U24222 ( .A(round_reg[100]), .B(n22272), .Z(n19480) );
  AND U24223 ( .A(n20448), .B(n21304), .Z(n24379) );
  IV U24224 ( .A(n23831), .Z(n21304) );
  XOR U24225 ( .A(round_reg[1272]), .B(n21775), .Z(n23831) );
  XOR U24226 ( .A(round_reg[1281]), .B(n21602), .Z(n20448) );
  XNOR U24227 ( .A(n24380), .B(n20459), .Z(n14940) );
  XOR U24228 ( .A(round_reg[159]), .B(n24165), .Z(n20459) );
  ANDN U24229 ( .B(n20318), .A(n20316), .Z(n24380) );
  XNOR U24230 ( .A(round_reg[1344]), .B(n24381), .Z(n20316) );
  XOR U24231 ( .A(round_reg[968]), .B(n22977), .Z(n20318) );
  XOR U24232 ( .A(n24382), .B(n24383), .Z(n21034) );
  XNOR U24233 ( .A(n18756), .B(n19709), .Z(n24383) );
  XNOR U24234 ( .A(n24384), .B(n21915), .Z(n19709) );
  ANDN U24235 ( .B(n20533), .A(n20534), .Z(n24384) );
  XOR U24236 ( .A(round_reg[626]), .B(n22105), .Z(n20534) );
  XNOR U24237 ( .A(n24385), .B(n21918), .Z(n18756) );
  NOR U24238 ( .A(n21052), .B(n21050), .Z(n24385) );
  XOR U24239 ( .A(round_reg[339]), .B(n23744), .Z(n21052) );
  XOR U24240 ( .A(n21319), .B(n24386), .Z(n24382) );
  XNOR U24241 ( .A(n16342), .B(n24387), .Z(n24386) );
  XNOR U24242 ( .A(n24388), .B(n21921), .Z(n16342) );
  AND U24243 ( .A(n20543), .B(n21284), .Z(n24388) );
  IV U24244 ( .A(n20545), .Z(n21284) );
  XOR U24245 ( .A(round_reg[460]), .B(n24389), .Z(n20545) );
  XNOR U24246 ( .A(n24390), .B(n21924), .Z(n21319) );
  ANDN U24247 ( .B(n20785), .A(n20786), .Z(n24390) );
  XOR U24248 ( .A(round_reg[558]), .B(n23735), .Z(n20786) );
  XNOR U24249 ( .A(n21726), .B(n18594), .Z(n15156) );
  IV U24250 ( .A(n17816), .Z(n18594) );
  XNOR U24251 ( .A(n24391), .B(n24031), .Z(n17816) );
  XNOR U24252 ( .A(n24392), .B(n24393), .Z(n24031) );
  XNOR U24253 ( .A(n19955), .B(n18653), .Z(n24393) );
  XOR U24254 ( .A(n24394), .B(n20005), .Z(n18653) );
  XNOR U24255 ( .A(round_reg[1157]), .B(n23426), .Z(n20005) );
  IV U24256 ( .A(n23485), .Z(n23426) );
  XNOR U24257 ( .A(n24395), .B(n24396), .Z(n23485) );
  XOR U24258 ( .A(round_reg[774]), .B(n24397), .Z(n21732) );
  XNOR U24259 ( .A(round_reg[412]), .B(n22119), .Z(n21733) );
  XOR U24260 ( .A(n24398), .B(n20009), .Z(n19955) );
  XNOR U24261 ( .A(round_reg[1082]), .B(n22991), .Z(n20009) );
  ANDN U24262 ( .B(n21728), .A(n21729), .Z(n24398) );
  XNOR U24263 ( .A(round_reg[584]), .B(n23986), .Z(n21729) );
  IV U24264 ( .A(n23206), .Z(n23986) );
  XNOR U24265 ( .A(round_reg[650]), .B(n24399), .Z(n21728) );
  XOR U24266 ( .A(n19694), .B(n24400), .Z(n24392) );
  XOR U24267 ( .A(n17990), .B(n17333), .Z(n24400) );
  XNOR U24268 ( .A(n24401), .B(n20000), .Z(n17333) );
  XOR U24269 ( .A(round_reg[1131]), .B(n23389), .Z(n20000) );
  AND U24270 ( .A(n23438), .B(n23617), .Z(n24401) );
  IV U24271 ( .A(n24402), .Z(n23617) );
  XNOR U24272 ( .A(n24403), .B(n23431), .Z(n17990) );
  XOR U24273 ( .A(round_reg[989]), .B(n23910), .Z(n23431) );
  XOR U24274 ( .A(round_reg[942]), .B(n24404), .Z(n21739) );
  XOR U24275 ( .A(round_reg[516]), .B(n24405), .Z(n21740) );
  XNOR U24276 ( .A(n24406), .B(n23217), .Z(n19694) );
  XOR U24277 ( .A(round_reg[1229]), .B(n24214), .Z(n23217) );
  AND U24278 ( .A(n21736), .B(n23435), .Z(n24406) );
  XOR U24279 ( .A(round_reg[871]), .B(n22361), .Z(n23435) );
  XOR U24280 ( .A(round_reg[482]), .B(n24407), .Z(n21736) );
  XNOR U24281 ( .A(n24408), .B(n23438), .Z(n21726) );
  XOR U24282 ( .A(round_reg[728]), .B(n23275), .Z(n23438) );
  ANDN U24283 ( .B(n24402), .A(n19998), .Z(n24408) );
  XOR U24284 ( .A(round_reg[287]), .B(n24409), .Z(n19998) );
  XOR U24285 ( .A(round_reg[361]), .B(n24221), .Z(n24402) );
  XNOR U24286 ( .A(n18046), .B(n24057), .Z(n14574) );
  XOR U24287 ( .A(n24410), .B(n21071), .Z(n24057) );
  AND U24288 ( .A(n23704), .B(n23703), .Z(n24410) );
  XNOR U24289 ( .A(n24411), .B(n23612), .Z(n18046) );
  XNOR U24290 ( .A(n24412), .B(n24413), .Z(n23612) );
  XOR U24291 ( .A(n16002), .B(n18734), .Z(n24413) );
  XOR U24292 ( .A(n24414), .B(n21070), .Z(n18734) );
  ANDN U24293 ( .B(n21071), .A(n23703), .Z(n24414) );
  XOR U24294 ( .A(round_reg[941]), .B(n21193), .Z(n23703) );
  XNOR U24295 ( .A(round_reg[988]), .B(n24415), .Z(n21071) );
  XOR U24296 ( .A(n24416), .B(n24417), .Z(n16002) );
  ANDN U24297 ( .B(n24059), .A(n23709), .Z(n24416) );
  XOR U24298 ( .A(round_reg[773]), .B(n22365), .Z(n23709) );
  XOR U24299 ( .A(n19165), .B(n24418), .Z(n24412) );
  XOR U24300 ( .A(n18538), .B(n17113), .Z(n24418) );
  XNOR U24301 ( .A(n24419), .B(n21059), .Z(n17113) );
  ANDN U24302 ( .B(n21060), .A(n23706), .Z(n24419) );
  XOR U24303 ( .A(round_reg[870]), .B(n23267), .Z(n23706) );
  XNOR U24304 ( .A(round_reg[1228]), .B(n23479), .Z(n21060) );
  XNOR U24305 ( .A(n24420), .B(n22163), .Z(n18538) );
  ANDN U24306 ( .B(n22164), .A(n23699), .Z(n24420) );
  XOR U24307 ( .A(round_reg[649]), .B(n24421), .Z(n23699) );
  XNOR U24308 ( .A(round_reg[1081]), .B(n24422), .Z(n22164) );
  XNOR U24309 ( .A(n24423), .B(n21063), .Z(n19165) );
  ANDN U24310 ( .B(n21064), .A(n24064), .Z(n24423) );
  XOR U24311 ( .A(round_reg[727]), .B(n23486), .Z(n24064) );
  XNOR U24312 ( .A(round_reg[1130]), .B(n24424), .Z(n21064) );
  XOR U24313 ( .A(n11359), .B(n24425), .Z(n24277) );
  XNOR U24314 ( .A(n12795), .B(n9717), .Z(n24425) );
  XNOR U24315 ( .A(n24426), .B(n14582), .Z(n9717) );
  XNOR U24316 ( .A(n17553), .B(n24174), .Z(n14582) );
  XOR U24317 ( .A(n24427), .B(n24428), .Z(n24174) );
  NOR U24318 ( .A(n22548), .B(n22552), .Z(n24427) );
  XOR U24319 ( .A(round_reg[1173]), .B(n22984), .Z(n22552) );
  XOR U24320 ( .A(n20228), .B(n22456), .Z(n17553) );
  XNOR U24321 ( .A(n24429), .B(n24430), .Z(n22456) );
  XNOR U24322 ( .A(n18120), .B(n18894), .Z(n24430) );
  XOR U24323 ( .A(n24431), .B(n23636), .Z(n18894) );
  ANDN U24324 ( .B(n24170), .A(n22556), .Z(n24431) );
  XOR U24325 ( .A(round_reg[1318]), .B(n22201), .Z(n22556) );
  XNOR U24326 ( .A(n24432), .B(n23640), .Z(n18120) );
  XOR U24327 ( .A(round_reg[1472]), .B(n24163), .Z(n22564) );
  XOR U24328 ( .A(n18436), .B(n24433), .Z(n24429) );
  XOR U24329 ( .A(n23167), .B(n19735), .Z(n24433) );
  XNOR U24330 ( .A(n24434), .B(n23633), .Z(n19735) );
  XNOR U24331 ( .A(round_reg[1537]), .B(n22834), .Z(n22548) );
  XNOR U24332 ( .A(n24435), .B(n23638), .Z(n23167) );
  XOR U24333 ( .A(round_reg[1411]), .B(n22757), .Z(n22560) );
  XNOR U24334 ( .A(n24436), .B(n23631), .Z(n18436) );
  XOR U24335 ( .A(round_reg[1381]), .B(n22515), .Z(n22545) );
  IV U24336 ( .A(n24374), .Z(n22515) );
  XOR U24337 ( .A(n24437), .B(n24438), .Z(n20228) );
  XOR U24338 ( .A(n20308), .B(n19339), .Z(n24438) );
  XOR U24339 ( .A(n24439), .B(n22257), .Z(n19339) );
  XOR U24340 ( .A(round_reg[1380]), .B(n22272), .Z(n22257) );
  XOR U24341 ( .A(round_reg[957]), .B(n24440), .Z(n23977) );
  XNOR U24342 ( .A(round_reg[1004]), .B(n23785), .Z(n23173) );
  XOR U24343 ( .A(n23179), .B(n24441), .Z(n20308) );
  XOR U24344 ( .A(n24442), .B(n4579), .Z(n24441) );
  NAND U24345 ( .A(n4364), .B(n24341), .Z(n4579) );
  AND U24346 ( .A(n6835), .B(n11363), .Z(n4364) );
  IV U24347 ( .A(rc_i[0]), .Z(n6835) );
  AND U24348 ( .A(n23180), .B(n23970), .Z(n24442) );
  XNOR U24349 ( .A(round_reg[789]), .B(n23130), .Z(n23970) );
  XOR U24350 ( .A(round_reg[1172]), .B(n22979), .Z(n23180) );
  XNOR U24351 ( .A(round_reg[1536]), .B(n24443), .Z(n23179) );
  XOR U24352 ( .A(n18555), .B(n24444), .Z(n24437) );
  XOR U24353 ( .A(n17545), .B(n18248), .Z(n24444) );
  XNOR U24354 ( .A(n24445), .B(n22244), .Z(n18248) );
  XOR U24355 ( .A(round_reg[1317]), .B(n24157), .Z(n22244) );
  AND U24356 ( .A(n23981), .B(n23980), .Z(n24445) );
  XOR U24357 ( .A(round_reg[1244]), .B(n24446), .Z(n23980) );
  XNOR U24358 ( .A(round_reg[886]), .B(n24274), .Z(n23981) );
  XNOR U24359 ( .A(n24447), .B(n22254), .Z(n17545) );
  XOR U24360 ( .A(round_reg[1410]), .B(n24161), .Z(n22254) );
  ANDN U24361 ( .B(n23182), .A(n23975), .Z(n24447) );
  XOR U24362 ( .A(round_reg[665]), .B(n21198), .Z(n23975) );
  XNOR U24363 ( .A(round_reg[1033]), .B(n24448), .Z(n23182) );
  XNOR U24364 ( .A(n24449), .B(n22248), .Z(n18555) );
  XOR U24365 ( .A(round_reg[1535]), .B(n23904), .Z(n22248) );
  AND U24366 ( .A(n23176), .B(n23972), .Z(n24449) );
  XNOR U24367 ( .A(round_reg[743]), .B(n24450), .Z(n23972) );
  XNOR U24368 ( .A(round_reg[1146]), .B(n24451), .Z(n23176) );
  ANDN U24369 ( .B(n24452), .A(n16537), .Z(n24426) );
  XNOR U24370 ( .A(n24453), .B(n15422), .Z(n12795) );
  XNOR U24371 ( .A(n24454), .B(n18355), .Z(n15422) );
  IV U24372 ( .A(n19350), .Z(n18355) );
  XOR U24373 ( .A(n18562), .B(n19140), .Z(n19350) );
  XNOR U24374 ( .A(n24455), .B(n24456), .Z(n19140) );
  XNOR U24375 ( .A(n17932), .B(n18300), .Z(n24456) );
  XNOR U24376 ( .A(n24457), .B(n21466), .Z(n18300) );
  AND U24377 ( .A(n21114), .B(n21116), .Z(n24457) );
  XOR U24378 ( .A(round_reg[1282]), .B(n24458), .Z(n21116) );
  XNOR U24379 ( .A(n24459), .B(n21458), .Z(n17932) );
  NOR U24380 ( .A(n21106), .B(n21105), .Z(n24459) );
  XNOR U24381 ( .A(round_reg[1439]), .B(n24460), .Z(n21106) );
  XOR U24382 ( .A(n18697), .B(n24461), .Z(n24455) );
  XOR U24383 ( .A(n20625), .B(n23208), .Z(n24461) );
  XNOR U24384 ( .A(n24462), .B(n21469), .Z(n23208) );
  ANDN U24385 ( .B(n21101), .A(n21102), .Z(n24462) );
  XNOR U24386 ( .A(round_reg[1565]), .B(n24463), .Z(n21102) );
  XNOR U24387 ( .A(n24464), .B(n21462), .Z(n20625) );
  NOR U24388 ( .A(n21111), .B(n21110), .Z(n24464) );
  XOR U24389 ( .A(round_reg[1500]), .B(n23253), .Z(n21111) );
  XNOR U24390 ( .A(n24465), .B(n21472), .Z(n18697) );
  AND U24391 ( .A(n21118), .B(n21120), .Z(n24465) );
  XOR U24392 ( .A(round_reg[1345]), .B(n24466), .Z(n21120) );
  XOR U24393 ( .A(n24467), .B(n24468), .Z(n18562) );
  XNOR U24394 ( .A(n17568), .B(n21494), .Z(n24468) );
  XNOR U24395 ( .A(n24469), .B(n21443), .Z(n21494) );
  ANDN U24396 ( .B(n23835), .A(n24470), .Z(n24469) );
  XNOR U24397 ( .A(n24471), .B(n23859), .Z(n17568) );
  AND U24398 ( .A(n23837), .B(n24472), .Z(n24471) );
  XOR U24399 ( .A(n19451), .B(n24473), .Z(n24467) );
  XOR U24400 ( .A(n15916), .B(n24474), .Z(n24473) );
  XNOR U24401 ( .A(n24475), .B(n23186), .Z(n15916) );
  AND U24402 ( .A(n24476), .B(n23846), .Z(n24475) );
  IV U24403 ( .A(n24477), .Z(n23846) );
  XNOR U24404 ( .A(n24478), .B(n21452), .Z(n19451) );
  AND U24405 ( .A(n23844), .B(n24479), .Z(n24478) );
  IV U24406 ( .A(n24480), .Z(n23844) );
  AND U24407 ( .A(n15146), .B(n15423), .Z(n24453) );
  XOR U24408 ( .A(n24481), .B(n19703), .Z(n15423) );
  XOR U24409 ( .A(n19608), .B(n20140), .Z(n19703) );
  XOR U24410 ( .A(n24482), .B(n24483), .Z(n20140) );
  XNOR U24411 ( .A(n20022), .B(n20851), .Z(n24483) );
  XNOR U24412 ( .A(n24484), .B(n20857), .Z(n20851) );
  XOR U24413 ( .A(round_reg[702]), .B(n24485), .Z(n20857) );
  ANDN U24414 ( .B(n20858), .A(n22345), .Z(n24484) );
  XNOR U24415 ( .A(n24486), .B(n20870), .Z(n20022) );
  XOR U24416 ( .A(round_reg[859]), .B(n24342), .Z(n20870) );
  ANDN U24417 ( .B(n20871), .A(n22340), .Z(n24486) );
  XOR U24418 ( .A(n17412), .B(n24487), .Z(n24482) );
  XOR U24419 ( .A(n19212), .B(n19151), .Z(n24487) );
  XNOR U24420 ( .A(n24488), .B(n20874), .Z(n19151) );
  XOR U24421 ( .A(round_reg[930]), .B(n24019), .Z(n20874) );
  ANDN U24422 ( .B(n20875), .A(n22348), .Z(n24488) );
  XNOR U24423 ( .A(n24489), .B(n20861), .Z(n19212) );
  XOR U24424 ( .A(round_reg[716]), .B(n24490), .Z(n20861) );
  ANDN U24425 ( .B(n20862), .A(n24491), .Z(n24489) );
  XNOR U24426 ( .A(n24492), .B(n20866), .Z(n17412) );
  XOR U24427 ( .A(round_reg[826]), .B(n24493), .Z(n20866) );
  ANDN U24428 ( .B(n24494), .A(n22337), .Z(n24492) );
  XNOR U24429 ( .A(n24495), .B(n24496), .Z(n19608) );
  XNOR U24430 ( .A(n18420), .B(n21878), .Z(n24496) );
  XNOR U24431 ( .A(n24497), .B(n21882), .Z(n21878) );
  XOR U24432 ( .A(round_reg[22]), .B(n23596), .Z(n21882) );
  ANDN U24433 ( .B(n21883), .A(n20961), .Z(n24497) );
  XNOR U24434 ( .A(n24498), .B(n21891), .Z(n18420) );
  XOR U24435 ( .A(round_reg[167]), .B(n21189), .Z(n21891) );
  ANDN U24436 ( .B(n21892), .A(n22588), .Z(n24498) );
  XOR U24437 ( .A(n19050), .B(n24499), .Z(n24495) );
  XOR U24438 ( .A(n19121), .B(n18035), .Z(n24499) );
  XNOR U24439 ( .A(n24500), .B(n21894), .Z(n18035) );
  XOR U24440 ( .A(round_reg[226]), .B(n23480), .Z(n21894) );
  ANDN U24441 ( .B(n21895), .A(n20950), .Z(n24500) );
  XNOR U24442 ( .A(n24501), .B(n23125), .Z(n19121) );
  XOR U24443 ( .A(round_reg[108]), .B(n24364), .Z(n23125) );
  ANDN U24444 ( .B(n24502), .A(n22377), .Z(n24501) );
  XNOR U24445 ( .A(n24503), .B(n21885), .Z(n19050) );
  XOR U24446 ( .A(round_reg[274]), .B(n24504), .Z(n21885) );
  ANDN U24447 ( .B(n21886), .A(n20954), .Z(n24503) );
  XOR U24448 ( .A(n16348), .B(n24505), .Z(n15146) );
  XNOR U24449 ( .A(n24506), .B(n24507), .Z(n22168) );
  XNOR U24450 ( .A(n19188), .B(n18526), .Z(n24507) );
  XNOR U24451 ( .A(n24508), .B(n23348), .Z(n18526) );
  XOR U24452 ( .A(round_reg[1368]), .B(n23275), .Z(n23348) );
  XOR U24453 ( .A(n24509), .B(n24510), .Z(n23275) );
  AND U24454 ( .A(n23054), .B(n23052), .Z(n24508) );
  XOR U24455 ( .A(round_reg[992]), .B(n21606), .Z(n23052) );
  XNOR U24456 ( .A(round_reg[945]), .B(n22962), .Z(n23054) );
  XNOR U24457 ( .A(n24511), .B(n23346), .Z(n19188) );
  XOR U24458 ( .A(round_reg[1588]), .B(n24084), .Z(n23346) );
  ANDN U24459 ( .B(n22742), .A(n23056), .Z(n24511) );
  XNOR U24460 ( .A(round_reg[1160]), .B(n21783), .Z(n23056) );
  XNOR U24461 ( .A(round_reg[777]), .B(n23283), .Z(n22742) );
  XOR U24462 ( .A(n18016), .B(n24512), .Z(n24506) );
  XOR U24463 ( .A(n19705), .B(n23336), .Z(n24512) );
  XNOR U24464 ( .A(n24513), .B(n23344), .Z(n23336) );
  XOR U24465 ( .A(round_reg[1462]), .B(n24514), .Z(n23344) );
  AND U24466 ( .A(n22732), .B(n23061), .Z(n24513) );
  XNOR U24467 ( .A(round_reg[1085]), .B(n22764), .Z(n23061) );
  XNOR U24468 ( .A(round_reg[653]), .B(n24515), .Z(n22732) );
  XOR U24469 ( .A(n24516), .B(n24025), .Z(n19705) );
  IV U24470 ( .A(n23341), .Z(n24025) );
  XOR U24471 ( .A(round_reg[1305]), .B(n21198), .Z(n23341) );
  ANDN U24472 ( .B(n23059), .A(n22746), .Z(n24516) );
  XOR U24473 ( .A(round_reg[874]), .B(n23920), .Z(n22746) );
  XOR U24474 ( .A(round_reg[1232]), .B(n22265), .Z(n23059) );
  XNOR U24475 ( .A(n24517), .B(n24001), .Z(n18016) );
  XOR U24476 ( .A(round_reg[1523]), .B(n24518), .Z(n24001) );
  ANDN U24477 ( .B(n23063), .A(n22736), .Z(n24517) );
  XOR U24478 ( .A(round_reg[731]), .B(n24519), .Z(n22736) );
  XOR U24479 ( .A(round_reg[1134]), .B(n23908), .Z(n23063) );
  XOR U24480 ( .A(n24520), .B(n24521), .Z(n23764) );
  XNOR U24481 ( .A(n19290), .B(n19303), .Z(n24521) );
  XOR U24482 ( .A(n24522), .B(n20471), .Z(n19303) );
  XOR U24483 ( .A(round_reg[588]), .B(n24523), .Z(n20471) );
  ANDN U24484 ( .B(n24524), .A(n22114), .Z(n24522) );
  XNOR U24485 ( .A(n24525), .B(n20489), .Z(n19290) );
  XNOR U24486 ( .A(round_reg[520]), .B(n21783), .Z(n20489) );
  NOR U24487 ( .A(n20488), .B(n22104), .Z(n24525) );
  XOR U24488 ( .A(n16042), .B(n24526), .Z(n24520) );
  XNOR U24489 ( .A(n19535), .B(n19452), .Z(n24526) );
  XNOR U24490 ( .A(n24527), .B(n20485), .Z(n19452) );
  XOR U24491 ( .A(round_reg[486]), .B(n23988), .Z(n20485) );
  ANDN U24492 ( .B(n20484), .A(n22111), .Z(n24527) );
  XNOR U24493 ( .A(n24528), .B(n20480), .Z(n19535) );
  XOR U24494 ( .A(round_reg[416]), .B(n22268), .Z(n20480) );
  ANDN U24495 ( .B(n24529), .A(n22107), .Z(n24528) );
  XNOR U24496 ( .A(n24530), .B(n20475), .Z(n16042) );
  XOR U24497 ( .A(round_reg[365]), .B(n22374), .Z(n20475) );
  ANDN U24498 ( .B(n20476), .A(n22117), .Z(n24530) );
  XNOR U24499 ( .A(n24531), .B(n14586), .Z(n11359) );
  XNOR U24500 ( .A(n24387), .B(n18757), .Z(n14586) );
  IV U24501 ( .A(n16343), .Z(n18757) );
  XNOR U24502 ( .A(n24532), .B(n24533), .Z(n20444) );
  XNOR U24503 ( .A(n18134), .B(n21906), .Z(n24533) );
  XNOR U24504 ( .A(n24534), .B(n21297), .Z(n21906) );
  XNOR U24505 ( .A(round_reg[1407]), .B(n22371), .Z(n21297) );
  ANDN U24506 ( .B(n21924), .A(n20785), .Z(n24534) );
  XOR U24507 ( .A(round_reg[920]), .B(n23406), .Z(n20785) );
  XOR U24508 ( .A(round_reg[967]), .B(n23492), .Z(n21924) );
  XOR U24509 ( .A(n24535), .B(n21292), .Z(n18134) );
  XNOR U24510 ( .A(round_reg[1563]), .B(n24156), .Z(n21292) );
  ANDN U24511 ( .B(n21912), .A(n20539), .Z(n24535) );
  XOR U24512 ( .A(n19695), .B(n24536), .Z(n24532) );
  XOR U24513 ( .A(n19315), .B(n18811), .Z(n24536) );
  XOR U24514 ( .A(n24537), .B(n21286), .Z(n18811) );
  XNOR U24515 ( .A(round_reg[1280]), .B(n24538), .Z(n21286) );
  XOR U24516 ( .A(round_reg[849]), .B(n23885), .Z(n20543) );
  XNOR U24517 ( .A(round_reg[1271]), .B(n23789), .Z(n21921) );
  XOR U24518 ( .A(n24539), .B(n21288), .Z(n19315) );
  XNOR U24519 ( .A(round_reg[1437]), .B(n24540), .Z(n21288) );
  ANDN U24520 ( .B(n21915), .A(n20533), .Z(n24539) );
  XOR U24521 ( .A(round_reg[692]), .B(n22796), .Z(n20533) );
  XOR U24522 ( .A(round_reg[1060]), .B(n22272), .Z(n21915) );
  XOR U24523 ( .A(n24541), .B(n21294), .Z(n19695) );
  AND U24524 ( .A(n21050), .B(n21918), .Z(n24541) );
  XOR U24525 ( .A(round_reg[1109]), .B(n23130), .Z(n21918) );
  XNOR U24526 ( .A(round_reg[706]), .B(n24132), .Z(n21050) );
  XNOR U24527 ( .A(n24542), .B(n24543), .Z(n19182) );
  XOR U24528 ( .A(n23712), .B(n17206), .Z(n24543) );
  XOR U24529 ( .A(n24544), .B(n23569), .Z(n17206) );
  XNOR U24530 ( .A(round_reg[691]), .B(n24545), .Z(n23569) );
  ANDN U24531 ( .B(n21040), .A(n20553), .Z(n24544) );
  XOR U24532 ( .A(round_reg[216]), .B(n24313), .Z(n20553) );
  XOR U24533 ( .A(round_reg[625]), .B(n22962), .Z(n21040) );
  XNOR U24534 ( .A(n24546), .B(n23571), .Z(n23712) );
  XOR U24535 ( .A(round_reg[705]), .B(n24547), .Z(n23571) );
  XOR U24536 ( .A(round_reg[264]), .B(n23206), .Z(n20559) );
  XOR U24537 ( .A(n24548), .B(n24549), .Z(n23206) );
  XNOR U24538 ( .A(round_reg[338]), .B(n21186), .Z(n21045) );
  XNOR U24539 ( .A(n18511), .B(n24550), .Z(n24542) );
  XOR U24540 ( .A(n21526), .B(n18240), .Z(n24550) );
  XOR U24541 ( .A(n24551), .B(n23573), .Z(n18240) );
  ANDN U24542 ( .B(n21038), .A(n20933), .Z(n24551) );
  XOR U24543 ( .A(round_reg[98]), .B(n23804), .Z(n20933) );
  IV U24544 ( .A(n23887), .Z(n23804) );
  XOR U24545 ( .A(round_reg[459]), .B(n24552), .Z(n21038) );
  XOR U24546 ( .A(n24553), .B(n23562), .Z(n21526) );
  XNOR U24547 ( .A(round_reg[919]), .B(n23395), .Z(n23562) );
  IV U24548 ( .A(n22687), .Z(n23395) );
  XNOR U24549 ( .A(n24555), .B(n24556), .Z(n24510) );
  XNOR U24550 ( .A(round_reg[23]), .B(round_reg[1303]), .Z(n24556) );
  XOR U24551 ( .A(round_reg[343]), .B(n24557), .Z(n24555) );
  XOR U24552 ( .A(round_reg[983]), .B(round_reg[663]), .Z(n24557) );
  ANDN U24553 ( .B(n21047), .A(n20563), .Z(n24553) );
  XOR U24554 ( .A(round_reg[157]), .B(n23902), .Z(n20563) );
  XOR U24555 ( .A(round_reg[557]), .B(n24309), .Z(n21047) );
  XOR U24556 ( .A(n24558), .B(n23565), .Z(n18511) );
  XOR U24557 ( .A(round_reg[815]), .B(n21196), .Z(n23565) );
  ANDN U24558 ( .B(n21043), .A(n20549), .Z(n24558) );
  XOR U24559 ( .A(round_reg[12]), .B(n22368), .Z(n20549) );
  XOR U24560 ( .A(round_reg[389]), .B(n24559), .Z(n21043) );
  XNOR U24561 ( .A(n24560), .B(n21912), .Z(n24387) );
  XOR U24562 ( .A(round_reg[1199]), .B(n21309), .Z(n21912) );
  AND U24563 ( .A(n20539), .B(n21291), .Z(n24560) );
  IV U24564 ( .A(n20541), .Z(n21291) );
  XOR U24565 ( .A(round_reg[390]), .B(n23883), .Z(n20541) );
  XOR U24566 ( .A(round_reg[816]), .B(n23963), .Z(n20539) );
  AND U24567 ( .A(n15149), .B(n15148), .Z(n24531) );
  XOR U24568 ( .A(n20836), .B(n18625), .Z(n15148) );
  XNOR U24569 ( .A(n24561), .B(n24562), .Z(n18599) );
  XNOR U24570 ( .A(n21793), .B(n18509), .Z(n24562) );
  XNOR U24571 ( .A(n24563), .B(n22037), .Z(n18509) );
  XOR U24572 ( .A(round_reg[1055]), .B(n23670), .Z(n22037) );
  XNOR U24573 ( .A(round_reg[687]), .B(n24564), .Z(n20832) );
  XNOR U24574 ( .A(round_reg[621]), .B(n21193), .Z(n19753) );
  XNOR U24575 ( .A(n24567), .B(n22039), .Z(n21793) );
  XOR U24576 ( .A(round_reg[1104]), .B(n24568), .Z(n22039) );
  ANDN U24577 ( .B(n19762), .A(n20834), .Z(n24567) );
  XOR U24578 ( .A(round_reg[765]), .B(n22764), .Z(n20834) );
  XNOR U24579 ( .A(round_reg[334]), .B(n22115), .Z(n19762) );
  XNOR U24580 ( .A(n19012), .B(n24569), .Z(n24561) );
  XOR U24581 ( .A(n18839), .B(n17202), .Z(n24569) );
  XNOR U24582 ( .A(n24570), .B(n22032), .Z(n17202) );
  XNOR U24583 ( .A(round_reg[1194]), .B(n23920), .Z(n22032) );
  XNOR U24584 ( .A(n24571), .B(n24572), .Z(n23920) );
  AND U24585 ( .A(n19758), .B(n20840), .Z(n24570) );
  IV U24586 ( .A(n22031), .Z(n20840) );
  XNOR U24587 ( .A(round_reg[811]), .B(n23389), .Z(n22031) );
  XNOR U24588 ( .A(round_reg[385]), .B(n24547), .Z(n19758) );
  XNOR U24589 ( .A(n24573), .B(n22035), .Z(n18839) );
  XNOR U24590 ( .A(round_reg[1266]), .B(n22105), .Z(n22035) );
  ANDN U24591 ( .B(n19749), .A(n20838), .Z(n24573) );
  XNOR U24592 ( .A(round_reg[844]), .B(n22279), .Z(n20838) );
  XNOR U24593 ( .A(round_reg[455]), .B(n21766), .Z(n19749) );
  XNOR U24594 ( .A(n24574), .B(n22988), .Z(n19012) );
  XOR U24595 ( .A(round_reg[962]), .B(n24458), .Z(n22988) );
  IV U24596 ( .A(n22442), .Z(n24458) );
  XOR U24597 ( .A(n24575), .B(n24576), .Z(n19718) );
  XNOR U24598 ( .A(n16010), .B(n17479), .Z(n24576) );
  XOR U24599 ( .A(n24577), .B(n22963), .Z(n17479) );
  ANDN U24600 ( .B(n22071), .A(n22069), .Z(n24577) );
  XNOR U24601 ( .A(round_reg[1338]), .B(n24578), .Z(n22071) );
  XNOR U24602 ( .A(n24579), .B(n22960), .Z(n16010) );
  XOR U24603 ( .A(round_reg[1431]), .B(n23254), .Z(n21689) );
  XOR U24604 ( .A(n18324), .B(n24580), .Z(n24575) );
  XOR U24605 ( .A(n18492), .B(n24581), .Z(n24580) );
  XNOR U24606 ( .A(n24582), .B(n22970), .Z(n18492) );
  ANDN U24607 ( .B(n22067), .A(n21693), .Z(n24582) );
  XOR U24608 ( .A(round_reg[1492]), .B(n22979), .Z(n21693) );
  XNOR U24609 ( .A(n24583), .B(n22973), .Z(n18324) );
  AND U24610 ( .A(n21683), .B(n22062), .Z(n24583) );
  IV U24611 ( .A(n24584), .Z(n22062) );
  XNOR U24612 ( .A(round_reg[1557]), .B(n23266), .Z(n21683) );
  XNOR U24613 ( .A(n24585), .B(n22992), .Z(n20836) );
  XNOR U24614 ( .A(round_reg[915]), .B(n24202), .Z(n22992) );
  AND U24615 ( .A(n19768), .B(n19766), .Z(n24585) );
  XOR U24616 ( .A(round_reg[553]), .B(n22972), .Z(n19766) );
  XNOR U24617 ( .A(round_reg[153]), .B(n21613), .Z(n19768) );
  XOR U24618 ( .A(n15903), .B(n24586), .Z(n15149) );
  XNOR U24619 ( .A(n23441), .B(n23627), .Z(n15903) );
  XNOR U24620 ( .A(n24587), .B(n24588), .Z(n23627) );
  XNOR U24621 ( .A(n17915), .B(n19447), .Z(n24588) );
  XNOR U24622 ( .A(n24589), .B(n22571), .Z(n19447) );
  XOR U24623 ( .A(round_reg[74]), .B(n22839), .Z(n22571) );
  ANDN U24624 ( .B(n22572), .A(n22470), .Z(n24589) );
  XNOR U24625 ( .A(n24590), .B(n22580), .Z(n17915) );
  XOR U24626 ( .A(round_reg[133]), .B(n22365), .Z(n22580) );
  XOR U24627 ( .A(n19701), .B(n24591), .Z(n24587) );
  XOR U24628 ( .A(n22541), .B(n18246), .Z(n24591) );
  XNOR U24629 ( .A(n24592), .B(n24187), .Z(n18246) );
  XOR U24630 ( .A(round_reg[304]), .B(n24053), .Z(n24187) );
  AND U24631 ( .A(n24193), .B(n24593), .Z(n24592) );
  XNOR U24632 ( .A(n24594), .B(n22808), .Z(n22541) );
  XOR U24633 ( .A(round_reg[192]), .B(n24163), .Z(n22808) );
  AND U24634 ( .A(n22809), .B(n22474), .Z(n24594) );
  XNOR U24635 ( .A(n24595), .B(n22577), .Z(n19701) );
  XOR U24636 ( .A(round_reg[52]), .B(n22796), .Z(n22577) );
  AND U24637 ( .A(n22578), .B(n22464), .Z(n24595) );
  XOR U24638 ( .A(n24596), .B(n24597), .Z(n23441) );
  XNOR U24639 ( .A(n18478), .B(n20240), .Z(n24597) );
  XOR U24640 ( .A(n24598), .B(n21382), .Z(n20240) );
  ANDN U24641 ( .B(n21383), .A(n21593), .Z(n24598) );
  XOR U24642 ( .A(n24599), .B(n21378), .Z(n18478) );
  AND U24643 ( .A(n21379), .B(n21590), .Z(n24599) );
  XNOR U24644 ( .A(n16361), .B(n24600), .Z(n24596) );
  XOR U24645 ( .A(n17515), .B(n16841), .Z(n24600) );
  XOR U24646 ( .A(n24601), .B(n21373), .Z(n16841) );
  ANDN U24647 ( .B(n21374), .A(n22386), .Z(n24601) );
  XOR U24648 ( .A(n24602), .B(n21386), .Z(n17515) );
  AND U24649 ( .A(n21387), .B(n24603), .Z(n24602) );
  XOR U24650 ( .A(n24604), .B(n21369), .Z(n16361) );
  XOR U24651 ( .A(n24605), .B(n14583), .Z(n15152) );
  IV U24652 ( .A(n24452), .Z(n14583) );
  XOR U24653 ( .A(n23222), .B(n18423), .Z(n24452) );
  IV U24654 ( .A(n15615), .Z(n18423) );
  XNOR U24655 ( .A(n24606), .B(n24607), .Z(n18329) );
  XNOR U24656 ( .A(n23509), .B(n18602), .Z(n24607) );
  XNOR U24657 ( .A(n24608), .B(n22498), .Z(n18602) );
  NOR U24658 ( .A(n23228), .B(n23229), .Z(n24608) );
  XNOR U24659 ( .A(n24609), .B(n22485), .Z(n23509) );
  NOR U24660 ( .A(n23231), .B(n23232), .Z(n24609) );
  XOR U24661 ( .A(n24610), .B(n24611), .Z(n24606) );
  XNOR U24662 ( .A(n21633), .B(n16707), .Z(n24611) );
  XOR U24663 ( .A(n24612), .B(n22493), .Z(n16707) );
  AND U24664 ( .A(n23225), .B(n23224), .Z(n24612) );
  XOR U24665 ( .A(n24613), .B(n22489), .Z(n21633) );
  AND U24666 ( .A(n23234), .B(n23235), .Z(n24613) );
  XOR U24667 ( .A(n24614), .B(n24615), .Z(n21126) );
  XOR U24668 ( .A(n16745), .B(n23329), .Z(n24615) );
  XOR U24669 ( .A(n24616), .B(n22894), .Z(n23329) );
  NOR U24670 ( .A(n22288), .B(n24617), .Z(n24616) );
  XNOR U24671 ( .A(n24618), .B(n22889), .Z(n16745) );
  ANDN U24672 ( .B(n24619), .A(n22298), .Z(n24618) );
  XOR U24673 ( .A(n19387), .B(n24620), .Z(n24614) );
  XOR U24674 ( .A(n17393), .B(n18429), .Z(n24620) );
  XNOR U24675 ( .A(n24621), .B(n22896), .Z(n18429) );
  ANDN U24676 ( .B(n24622), .A(n22294), .Z(n24621) );
  XNOR U24677 ( .A(n24623), .B(n22887), .Z(n17393) );
  XNOR U24678 ( .A(n24626), .B(n22892), .Z(n19387) );
  NOR U24679 ( .A(n22284), .B(n24627), .Z(n24626) );
  XNOR U24680 ( .A(n24628), .B(n24629), .Z(n23222) );
  XOR U24681 ( .A(n22910), .B(n18425), .Z(n15428) );
  XOR U24682 ( .A(n24631), .B(n22875), .Z(n22910) );
  ANDN U24683 ( .B(n24632), .A(n23825), .Z(n24631) );
  XOR U24684 ( .A(n22617), .B(n16698), .Z(n16537) );
  XOR U24685 ( .A(n24194), .B(n19615), .Z(n16698) );
  XNOR U24686 ( .A(n24633), .B(n24634), .Z(n19615) );
  XNOR U24687 ( .A(n15599), .B(n18871), .Z(n24634) );
  XOR U24688 ( .A(n24635), .B(n20686), .Z(n18871) );
  XNOR U24689 ( .A(round_reg[910]), .B(n24636), .Z(n20686) );
  ANDN U24690 ( .B(n20685), .A(n22613), .Z(n24635) );
  XOR U24691 ( .A(round_reg[148]), .B(n23732), .Z(n22613) );
  XNOR U24692 ( .A(round_reg[548]), .B(n22822), .Z(n20685) );
  XNOR U24693 ( .A(n24637), .B(n20675), .Z(n15599) );
  XNOR U24694 ( .A(round_reg[682]), .B(n23420), .Z(n20675) );
  IV U24695 ( .A(n22649), .Z(n23420) );
  ANDN U24696 ( .B(n20676), .A(n22603), .Z(n24637) );
  XOR U24697 ( .A(round_reg[207]), .B(n23793), .Z(n22603) );
  XOR U24698 ( .A(round_reg[616]), .B(n24257), .Z(n20676) );
  XOR U24699 ( .A(n18207), .B(n24638), .Z(n24633) );
  XNOR U24700 ( .A(n19236), .B(n15635), .Z(n24638) );
  XNOR U24701 ( .A(n24639), .B(n22236), .Z(n15635) );
  XNOR U24702 ( .A(round_reg[839]), .B(n24028), .Z(n22236) );
  NOR U24703 ( .A(n22235), .B(n22600), .Z(n24639) );
  XOR U24704 ( .A(round_reg[89]), .B(n21760), .Z(n22600) );
  XNOR U24705 ( .A(round_reg[450]), .B(n24161), .Z(n22235) );
  XNOR U24706 ( .A(n24640), .B(n20681), .Z(n19236) );
  XNOR U24707 ( .A(round_reg[806]), .B(n23988), .Z(n20681) );
  ANDN U24708 ( .B(n20682), .A(n22607), .Z(n24640) );
  XOR U24709 ( .A(round_reg[3]), .B(n24136), .Z(n22607) );
  IV U24710 ( .A(n23599), .Z(n24136) );
  XOR U24711 ( .A(round_reg[444]), .B(n24026), .Z(n20682) );
  XNOR U24712 ( .A(n24641), .B(n24230), .Z(n18207) );
  XNOR U24713 ( .A(round_reg[760]), .B(n24642), .Z(n24230) );
  XNOR U24714 ( .A(round_reg[329]), .B(n24421), .Z(n22609) );
  XOR U24715 ( .A(round_reg[319]), .B(n21603), .Z(n22611) );
  XOR U24716 ( .A(n24643), .B(n24644), .Z(n24194) );
  XOR U24717 ( .A(n17936), .B(n19348), .Z(n24644) );
  XNOR U24718 ( .A(n24645), .B(n22761), .Z(n19348) );
  XOR U24719 ( .A(round_reg[683]), .B(n24078), .Z(n21867) );
  IV U24720 ( .A(n24302), .Z(n24078) );
  XOR U24721 ( .A(n24646), .B(n22767), .Z(n17936) );
  XNOR U24722 ( .A(n20668), .B(n24648), .Z(n24643) );
  XOR U24723 ( .A(n19890), .B(n17038), .Z(n24648) );
  XOR U24724 ( .A(n24649), .B(n22765), .Z(n17038) );
  AND U24725 ( .A(n22622), .B(n22593), .Z(n24649) );
  IV U24726 ( .A(n22623), .Z(n22593) );
  XOR U24727 ( .A(round_reg[807]), .B(n21189), .Z(n22623) );
  XNOR U24728 ( .A(n24650), .B(n22758), .Z(n19890) );
  NOR U24729 ( .A(n21857), .B(n22625), .Z(n24650) );
  XOR U24730 ( .A(round_reg[840]), .B(n21783), .Z(n21857) );
  XNOR U24731 ( .A(n24651), .B(n22770), .Z(n20668) );
  ANDN U24732 ( .B(n22627), .A(n21863), .Z(n24651) );
  XOR U24733 ( .A(round_reg[911]), .B(n22802), .Z(n21863) );
  XOR U24734 ( .A(n24652), .B(n24647), .Z(n22617) );
  NOR U24735 ( .A(n21854), .B(n21853), .Z(n24652) );
  XNOR U24736 ( .A(round_reg[761]), .B(n23623), .Z(n21853) );
  XOR U24737 ( .A(round_reg[330]), .B(n24116), .Z(n21854) );
  XOR U24738 ( .A(n11309), .B(n13291), .Z(n7076) );
  XNOR U24739 ( .A(n24653), .B(n14679), .Z(n13291) );
  ANDN U24740 ( .B(n16160), .A(n16662), .Z(n24653) );
  XOR U24741 ( .A(n24654), .B(n18018), .Z(n16160) );
  XOR U24742 ( .A(n24655), .B(n24656), .Z(n12714) );
  XNOR U24743 ( .A(n9797), .B(n11395), .Z(n24656) );
  XOR U24744 ( .A(n24657), .B(n18073), .Z(n11395) );
  XNOR U24745 ( .A(n16758), .B(n22396), .Z(n18073) );
  XOR U24746 ( .A(n24658), .B(n24659), .Z(n22396) );
  ANDN U24747 ( .B(n24660), .A(n21807), .Z(n24658) );
  XOR U24748 ( .A(n20809), .B(n19499), .Z(n16758) );
  XNOR U24749 ( .A(n24661), .B(n24662), .Z(n19499) );
  XOR U24750 ( .A(n18700), .B(n17207), .Z(n24662) );
  XOR U24751 ( .A(n24663), .B(n23307), .Z(n17207) );
  XNOR U24752 ( .A(round_reg[422]), .B(n23865), .Z(n23307) );
  NOR U24753 ( .A(n22422), .B(n22421), .Z(n24663) );
  XNOR U24754 ( .A(round_reg[45]), .B(n22374), .Z(n22421) );
  XOR U24755 ( .A(n24664), .B(n24665), .Z(n22374) );
  XOR U24756 ( .A(round_reg[1595]), .B(n22517), .Z(n22422) );
  XNOR U24757 ( .A(n24666), .B(n22087), .Z(n18700) );
  XNOR U24758 ( .A(round_reg[371]), .B(n23504), .Z(n22087) );
  XNOR U24759 ( .A(round_reg[297]), .B(n22760), .Z(n22086) );
  XOR U24760 ( .A(round_reg[1530]), .B(n23249), .Z(n22411) );
  XNOR U24761 ( .A(n18650), .B(n24667), .Z(n24661) );
  XOR U24762 ( .A(n19213), .B(n19912), .Z(n24667) );
  XNOR U24763 ( .A(n24668), .B(n22082), .Z(n19912) );
  XOR U24764 ( .A(round_reg[594]), .B(n24504), .Z(n22082) );
  AND U24765 ( .A(n22416), .B(n22414), .Z(n24668) );
  IV U24766 ( .A(n22083), .Z(n22414) );
  XNOR U24767 ( .A(round_reg[249]), .B(n22831), .Z(n22083) );
  XNOR U24768 ( .A(round_reg[1469]), .B(n21609), .Z(n22416) );
  XNOR U24769 ( .A(n24669), .B(n22092), .Z(n19213) );
  XOR U24770 ( .A(round_reg[492]), .B(n23598), .Z(n22092) );
  ANDN U24771 ( .B(n22093), .A(n22407), .Z(n24669) );
  XOR U24772 ( .A(round_reg[1312]), .B(n21606), .Z(n22407) );
  XNOR U24773 ( .A(round_reg[67]), .B(n21747), .Z(n22093) );
  XNOR U24774 ( .A(n24670), .B(n22097), .Z(n18650) );
  XNOR U24775 ( .A(round_reg[526]), .B(n22221), .Z(n22097) );
  AND U24776 ( .A(n22418), .B(n22096), .Z(n24670) );
  XOR U24777 ( .A(round_reg[190]), .B(n22435), .Z(n22096) );
  XNOR U24778 ( .A(round_reg[1375]), .B(n24673), .Z(n22418) );
  XOR U24779 ( .A(n24674), .B(n24675), .Z(n20809) );
  XOR U24780 ( .A(n17242), .B(n18268), .Z(n24675) );
  XNOR U24781 ( .A(n24676), .B(n22703), .Z(n18268) );
  ANDN U24782 ( .B(n24677), .A(n22399), .Z(n24676) );
  XNOR U24783 ( .A(n24678), .B(n21823), .Z(n17242) );
  NOR U24784 ( .A(n22403), .B(n22402), .Z(n24678) );
  XOR U24785 ( .A(n21122), .B(n24679), .Z(n24674) );
  XOR U24786 ( .A(n22076), .B(n18259), .Z(n24679) );
  XNOR U24787 ( .A(n24680), .B(n21809), .Z(n18259) );
  NOR U24788 ( .A(n24660), .B(n24659), .Z(n24680) );
  XNOR U24789 ( .A(n24681), .B(n21818), .Z(n22076) );
  ANDN U24790 ( .B(n23212), .A(n23213), .Z(n24681) );
  XOR U24791 ( .A(n24682), .B(n21812), .Z(n21122) );
  AND U24792 ( .A(n22394), .B(n22393), .Z(n24682) );
  NOR U24793 ( .A(n15880), .B(n15882), .Z(n24657) );
  XNOR U24794 ( .A(n21067), .B(n18002), .Z(n15882) );
  XNOR U24795 ( .A(n20029), .B(n24391), .Z(n18002) );
  XNOR U24796 ( .A(n24683), .B(n24684), .Z(n24391) );
  XNOR U24797 ( .A(n18345), .B(n16676), .Z(n24684) );
  XOR U24798 ( .A(n24685), .B(n23711), .Z(n16676) );
  XNOR U24799 ( .A(round_reg[411]), .B(n24519), .Z(n23711) );
  ANDN U24800 ( .B(n24417), .A(n23710), .Z(n24685) );
  XNOR U24801 ( .A(n24686), .B(n24065), .Z(n18345) );
  XOR U24802 ( .A(round_reg[360]), .B(n24687), .Z(n24065) );
  NOR U24803 ( .A(n21063), .B(n21062), .Z(n24686) );
  XNOR U24804 ( .A(round_reg[286]), .B(n23464), .Z(n21062) );
  XOR U24805 ( .A(round_reg[1519]), .B(n21309), .Z(n21063) );
  XOR U24806 ( .A(n24688), .B(n24689), .Z(n21309) );
  XNOR U24807 ( .A(n17594), .B(n24690), .Z(n24683) );
  XOR U24808 ( .A(n23676), .B(n18277), .Z(n24690) );
  XOR U24809 ( .A(n24691), .B(n23700), .Z(n18277) );
  XNOR U24810 ( .A(round_reg[583]), .B(n23916), .Z(n23700) );
  NOR U24811 ( .A(n22163), .B(n22162), .Z(n24691) );
  XNOR U24812 ( .A(round_reg[238]), .B(n23735), .Z(n22162) );
  XOR U24813 ( .A(round_reg[1458]), .B(n24692), .Z(n22163) );
  XNOR U24814 ( .A(n24693), .B(n23707), .Z(n23676) );
  XOR U24815 ( .A(round_reg[481]), .B(n24694), .Z(n23707) );
  ANDN U24816 ( .B(n21058), .A(n21059), .Z(n24693) );
  XOR U24817 ( .A(round_reg[1301]), .B(n23393), .Z(n21059) );
  XOR U24818 ( .A(round_reg[120]), .B(n24695), .Z(n21058) );
  XNOR U24819 ( .A(n24696), .B(n23704), .Z(n17594) );
  XNOR U24820 ( .A(round_reg[515]), .B(n24697), .Z(n23704) );
  XOR U24821 ( .A(round_reg[1364]), .B(n24155), .Z(n21070) );
  XNOR U24822 ( .A(round_reg[179]), .B(n23621), .Z(n21069) );
  XOR U24823 ( .A(n24698), .B(n24699), .Z(n20029) );
  XNOR U24824 ( .A(n20078), .B(n17368), .Z(n24699) );
  XOR U24825 ( .A(n24700), .B(n23691), .Z(n17368) );
  XOR U24826 ( .A(round_reg[1363]), .B(n21610), .Z(n23691) );
  ANDN U24827 ( .B(n22187), .A(n22185), .Z(n24700) );
  XNOR U24828 ( .A(round_reg[987]), .B(n23386), .Z(n22185) );
  XNOR U24829 ( .A(n24701), .B(n23694), .Z(n20078) );
  ANDN U24830 ( .B(n22178), .A(n22176), .Z(n24701) );
  XNOR U24831 ( .A(round_reg[1155]), .B(n24697), .Z(n22176) );
  XOR U24832 ( .A(n18633), .B(n24702), .Z(n24698) );
  XNOR U24833 ( .A(n20205), .B(n18146), .Z(n24702) );
  XNOR U24834 ( .A(n24703), .B(n23681), .Z(n18146) );
  XOR U24835 ( .A(round_reg[1300]), .B(n21318), .Z(n23681) );
  ANDN U24836 ( .B(n22195), .A(n22193), .Z(n24703) );
  XNOR U24837 ( .A(round_reg[1227]), .B(n24704), .Z(n22193) );
  XNOR U24838 ( .A(n24705), .B(n23688), .Z(n20205) );
  XNOR U24839 ( .A(round_reg[1457]), .B(n24285), .Z(n23688) );
  ANDN U24840 ( .B(n22182), .A(n22180), .Z(n24705) );
  XNOR U24841 ( .A(round_reg[1080]), .B(n24695), .Z(n22180) );
  XNOR U24842 ( .A(n24706), .B(n23684), .Z(n18633) );
  XOR U24843 ( .A(round_reg[1518]), .B(n23735), .Z(n23684) );
  ANDN U24844 ( .B(n22191), .A(n22189), .Z(n24706) );
  XNOR U24845 ( .A(round_reg[1129]), .B(n22372), .Z(n22189) );
  XOR U24846 ( .A(n24707), .B(n23710), .Z(n21067) );
  XNOR U24847 ( .A(round_reg[34]), .B(n23405), .Z(n23710) );
  NOR U24848 ( .A(n24417), .B(n24059), .Z(n24707) );
  XNOR U24849 ( .A(round_reg[1156]), .B(n24405), .Z(n24059) );
  XNOR U24850 ( .A(round_reg[1584]), .B(n24053), .Z(n24417) );
  XNOR U24851 ( .A(n24197), .B(n19441), .Z(n15880) );
  XNOR U24852 ( .A(n20284), .B(n20669), .Z(n19441) );
  XNOR U24853 ( .A(n24708), .B(n24709), .Z(n20669) );
  XNOR U24854 ( .A(n19554), .B(n15968), .Z(n24709) );
  XNOR U24855 ( .A(n24710), .B(n21865), .Z(n15968) );
  XOR U24856 ( .A(round_reg[149]), .B(n23130), .Z(n21865) );
  NOR U24857 ( .A(n22770), .B(n22627), .Z(n24710) );
  XOR U24858 ( .A(round_reg[1022]), .B(n24485), .Z(n22627) );
  XNOR U24859 ( .A(round_reg[1398]), .B(n21195), .Z(n22770) );
  IV U24860 ( .A(n23491), .Z(n21195) );
  XNOR U24861 ( .A(n24711), .B(n21855), .Z(n19554) );
  XOR U24862 ( .A(round_reg[256]), .B(n23151), .Z(n21855) );
  AND U24863 ( .A(n22767), .B(n24647), .Z(n24711) );
  XNOR U24864 ( .A(round_reg[1100]), .B(n24389), .Z(n24647) );
  XOR U24865 ( .A(round_reg[1489]), .B(n23885), .Z(n22767) );
  XOR U24866 ( .A(n19302), .B(n24712), .Z(n24708) );
  XOR U24867 ( .A(n21476), .B(n15253), .Z(n24712) );
  XOR U24868 ( .A(n24713), .B(n21858), .Z(n15253) );
  XNOR U24869 ( .A(round_reg[90]), .B(n24714), .Z(n21858) );
  XOR U24870 ( .A(round_reg[1335]), .B(n23959), .Z(n22758) );
  IV U24871 ( .A(n24715), .Z(n23959) );
  XNOR U24872 ( .A(round_reg[1262]), .B(n24128), .Z(n22625) );
  IV U24873 ( .A(n24404), .Z(n24128) );
  XNOR U24874 ( .A(n24716), .B(n21869), .Z(n21476) );
  XOR U24875 ( .A(round_reg[208]), .B(n24229), .Z(n21869) );
  AND U24876 ( .A(n22761), .B(n22619), .Z(n24716) );
  XNOR U24877 ( .A(round_reg[1051]), .B(n24519), .Z(n22619) );
  XOR U24878 ( .A(round_reg[1428]), .B(n23732), .Z(n22761) );
  XOR U24879 ( .A(n24717), .B(n24718), .Z(n23732) );
  XNOR U24880 ( .A(n24719), .B(n22595), .Z(n19302) );
  XOR U24881 ( .A(round_reg[4]), .B(n23016), .Z(n22595) );
  ANDN U24882 ( .B(n22765), .A(n22622), .Z(n24719) );
  XNOR U24883 ( .A(round_reg[1190]), .B(n24720), .Z(n22622) );
  XOR U24884 ( .A(round_reg[1554]), .B(n24504), .Z(n22765) );
  XOR U24885 ( .A(n24721), .B(n24722), .Z(n20284) );
  XNOR U24886 ( .A(n20937), .B(n22144), .Z(n24722) );
  XNOR U24887 ( .A(n24723), .B(n21849), .Z(n22144) );
  XOR U24888 ( .A(round_reg[762]), .B(n22991), .Z(n21849) );
  ANDN U24889 ( .B(n22776), .A(n23046), .Z(n24723) );
  XOR U24890 ( .A(round_reg[257]), .B(n22834), .Z(n23046) );
  IV U24891 ( .A(n23952), .Z(n22834) );
  XOR U24892 ( .A(n24724), .B(n24725), .Z(n23952) );
  XOR U24893 ( .A(round_reg[331]), .B(n21754), .Z(n22776) );
  XNOR U24894 ( .A(n24726), .B(n21842), .Z(n20937) );
  XOR U24895 ( .A(round_reg[841]), .B(n24727), .Z(n21842) );
  ANDN U24896 ( .B(n22781), .A(n24199), .Z(n24726) );
  XOR U24897 ( .A(round_reg[91]), .B(n24519), .Z(n24199) );
  XOR U24898 ( .A(round_reg[452]), .B(n24728), .Z(n22781) );
  XOR U24899 ( .A(n22753), .B(n24729), .Z(n24721) );
  XOR U24900 ( .A(n22699), .B(n18182), .Z(n24729) );
  XNOR U24901 ( .A(n24730), .B(n21837), .Z(n18182) );
  XOR U24902 ( .A(round_reg[912]), .B(n22265), .Z(n21837) );
  NOR U24903 ( .A(n20440), .B(n22784), .Z(n24730) );
  XOR U24904 ( .A(round_reg[550]), .B(n24720), .Z(n22784) );
  XOR U24905 ( .A(round_reg[150]), .B(n24378), .Z(n20440) );
  XNOR U24906 ( .A(n24731), .B(n21845), .Z(n22699) );
  XOR U24907 ( .A(round_reg[684]), .B(n23785), .Z(n21845) );
  XNOR U24908 ( .A(n24732), .B(n24733), .Z(n24328) );
  XNOR U24909 ( .A(round_reg[1579]), .B(round_reg[1259]), .Z(n24733) );
  XOR U24910 ( .A(round_reg[299]), .B(n24734), .Z(n24732) );
  XOR U24911 ( .A(round_reg[939]), .B(round_reg[619]), .Z(n24734) );
  ANDN U24912 ( .B(n22774), .A(n20433), .Z(n24731) );
  XNOR U24913 ( .A(n24736), .B(n21835), .Z(n22753) );
  XOR U24914 ( .A(round_reg[808]), .B(n22821), .Z(n21835) );
  NOR U24915 ( .A(n20429), .B(n22779), .Z(n24736) );
  XOR U24916 ( .A(round_reg[446]), .B(n23561), .Z(n22779) );
  XOR U24917 ( .A(round_reg[5]), .B(n23895), .Z(n20429) );
  XOR U24918 ( .A(n24737), .B(n22774), .Z(n24197) );
  XNOR U24919 ( .A(round_reg[618]), .B(n24738), .Z(n22774) );
  AND U24920 ( .A(n20433), .B(n21844), .Z(n24737) );
  IV U24921 ( .A(n20434), .Z(n21844) );
  XOR U24922 ( .A(round_reg[1429]), .B(n23130), .Z(n20434) );
  XOR U24923 ( .A(round_reg[209]), .B(n23885), .Z(n20433) );
  XNOR U24924 ( .A(n24741), .B(n19042), .Z(n9797) );
  XNOR U24925 ( .A(n20521), .B(n19984), .Z(n19042) );
  IV U24926 ( .A(n18763), .Z(n19984) );
  XOR U24927 ( .A(n24742), .B(n24264), .Z(n18763) );
  XNOR U24928 ( .A(n24743), .B(n24744), .Z(n24264) );
  XOR U24929 ( .A(n20137), .B(n17230), .Z(n24744) );
  XOR U24930 ( .A(n24745), .B(n21516), .Z(n17230) );
  XOR U24931 ( .A(round_reg[20]), .B(n21318), .Z(n21516) );
  IV U24932 ( .A(n24746), .Z(n21318) );
  AND U24933 ( .A(n20905), .B(n20907), .Z(n24745) );
  XOR U24934 ( .A(round_reg[1570]), .B(n24019), .Z(n20905) );
  XNOR U24935 ( .A(n24747), .B(n19357), .Z(n20137) );
  XOR U24936 ( .A(round_reg[224]), .B(n24254), .Z(n19357) );
  NOR U24937 ( .A(n20520), .B(n20519), .Z(n24747) );
  XNOR U24938 ( .A(round_reg[1444]), .B(n23482), .Z(n20519) );
  XOR U24939 ( .A(n20707), .B(n24748), .Z(n24743) );
  XNOR U24940 ( .A(n17475), .B(n18351), .Z(n24748) );
  XNOR U24941 ( .A(n24749), .B(n19361), .Z(n18351) );
  XNOR U24942 ( .A(round_reg[272]), .B(n22265), .Z(n19361) );
  XNOR U24943 ( .A(n24750), .B(n24751), .Z(n22265) );
  ANDN U24944 ( .B(n21537), .A(n20526), .Z(n24749) );
  XOR U24945 ( .A(round_reg[1505]), .B(n24752), .Z(n21537) );
  XOR U24946 ( .A(n24753), .B(n19368), .Z(n17475) );
  IV U24947 ( .A(n21540), .Z(n19368) );
  XOR U24948 ( .A(round_reg[106]), .B(n23528), .Z(n21540) );
  ANDN U24949 ( .B(n24754), .A(n21539), .Z(n24753) );
  XOR U24950 ( .A(n24755), .B(n19371), .Z(n20707) );
  XNOR U24951 ( .A(round_reg[165]), .B(n23919), .Z(n19371) );
  XNOR U24952 ( .A(round_reg[1350]), .B(n23883), .Z(n21533) );
  XOR U24953 ( .A(n24756), .B(n21539), .Z(n20521) );
  XNOR U24954 ( .A(round_reg[1287]), .B(n23492), .Z(n21539) );
  IV U24955 ( .A(n24757), .Z(n23492) );
  NOR U24956 ( .A(n19366), .B(n24754), .Z(n24756) );
  NOR U24957 ( .A(n15867), .B(n15868), .Z(n24741) );
  XOR U24958 ( .A(n22909), .B(n18425), .Z(n15868) );
  IV U24959 ( .A(n17363), .Z(n18425) );
  XNOR U24960 ( .A(n24758), .B(n24759), .Z(n21574) );
  XNOR U24961 ( .A(n17674), .B(n15622), .Z(n24759) );
  XOR U24962 ( .A(n24760), .B(n24258), .Z(n15622) );
  XNOR U24963 ( .A(round_reg[509]), .B(n21609), .Z(n24258) );
  ANDN U24964 ( .B(n20903), .A(n20901), .Z(n24760) );
  XNOR U24965 ( .A(round_reg[84]), .B(n24155), .Z(n20901) );
  XNOR U24966 ( .A(round_reg[1329]), .B(n22267), .Z(n20903) );
  XOR U24967 ( .A(n24761), .B(n24762), .Z(n22267) );
  XOR U24968 ( .A(n24763), .B(n22848), .Z(n17674) );
  XNOR U24969 ( .A(round_reg[611]), .B(n23256), .Z(n22848) );
  ANDN U24970 ( .B(n20893), .A(n20891), .Z(n24763) );
  XNOR U24971 ( .A(round_reg[202]), .B(n22366), .Z(n20891) );
  XNOR U24972 ( .A(round_reg[1422]), .B(n23134), .Z(n20893) );
  XOR U24973 ( .A(n18568), .B(n24764), .Z(n24758) );
  XOR U24974 ( .A(n18747), .B(n18264), .Z(n24764) );
  XOR U24975 ( .A(n24765), .B(n22853), .Z(n18264) );
  XNOR U24976 ( .A(round_reg[439]), .B(n24223), .Z(n22853) );
  XNOR U24977 ( .A(round_reg[62]), .B(n24485), .Z(n20887) );
  IV U24978 ( .A(n24315), .Z(n24485) );
  XOR U24979 ( .A(round_reg[1548]), .B(n24523), .Z(n20889) );
  XOR U24980 ( .A(n24766), .B(n22856), .Z(n18747) );
  XNOR U24981 ( .A(round_reg[324]), .B(n23016), .Z(n22856) );
  XNOR U24982 ( .A(round_reg[314]), .B(n23318), .Z(n20897) );
  XNOR U24983 ( .A(round_reg[1483]), .B(n24767), .Z(n20899) );
  XOR U24984 ( .A(n24768), .B(n22845), .Z(n18568) );
  XNOR U24985 ( .A(round_reg[543]), .B(n24769), .Z(n22845) );
  XNOR U24986 ( .A(round_reg[143]), .B(n23784), .Z(n21576) );
  XOR U24987 ( .A(round_reg[1392]), .B(n24770), .Z(n21578) );
  XOR U24988 ( .A(n24771), .B(n24772), .Z(n22355) );
  XNOR U24989 ( .A(n22840), .B(n18861), .Z(n24772) );
  XNOR U24990 ( .A(n24773), .B(n22866), .Z(n18861) );
  XOR U24991 ( .A(round_reg[1095]), .B(n21766), .Z(n22866) );
  ANDN U24992 ( .B(n22913), .A(n22865), .Z(n24773) );
  XNOR U24993 ( .A(round_reg[756]), .B(n23289), .Z(n22865) );
  XNOR U24994 ( .A(n24774), .B(n22874), .Z(n22840) );
  XOR U24995 ( .A(round_reg[1257]), .B(n22760), .Z(n22874) );
  XOR U24996 ( .A(n24775), .B(n24776), .Z(n22760) );
  ANDN U24997 ( .B(n22875), .A(n24632), .Z(n24774) );
  XOR U24998 ( .A(n15593), .B(n24777), .Z(n24771) );
  XNOR U24999 ( .A(n19233), .B(n19547), .Z(n24777) );
  XOR U25000 ( .A(n24778), .B(n22879), .Z(n19547) );
  XNOR U25001 ( .A(round_reg[1017]), .B(n23469), .Z(n22879) );
  ANDN U25002 ( .B(n22903), .A(n22878), .Z(n24778) );
  XOR U25003 ( .A(round_reg[906]), .B(n24779), .Z(n22878) );
  XNOR U25004 ( .A(n24780), .B(n24110), .Z(n19233) );
  IV U25005 ( .A(n22862), .Z(n24110) );
  XOR U25006 ( .A(round_reg[1046]), .B(n23591), .Z(n22862) );
  AND U25007 ( .A(n22905), .B(n24781), .Z(n24780) );
  XOR U25008 ( .A(round_reg[678]), .B(n22201), .Z(n22905) );
  IV U25009 ( .A(n24017), .Z(n22201) );
  XNOR U25010 ( .A(n24782), .B(n24783), .Z(n24017) );
  XNOR U25011 ( .A(n24784), .B(n22871), .Z(n15593) );
  XOR U25012 ( .A(round_reg[1185]), .B(n24752), .Z(n22871) );
  ANDN U25013 ( .B(n24785), .A(n22870), .Z(n24784) );
  XNOR U25014 ( .A(n24786), .B(n22870), .Z(n22909) );
  XNOR U25015 ( .A(round_reg[802]), .B(n24787), .Z(n22870) );
  XOR U25016 ( .A(n23375), .B(n19107), .Z(n15867) );
  IV U25017 ( .A(n18718), .Z(n19107) );
  XOR U25018 ( .A(n21932), .B(n19689), .Z(n18718) );
  XNOR U25019 ( .A(n24788), .B(n24789), .Z(n19689) );
  XOR U25020 ( .A(n19496), .B(n17791), .Z(n24789) );
  XOR U25021 ( .A(n24790), .B(n22676), .Z(n17791) );
  ANDN U25022 ( .B(n23369), .A(n23370), .Z(n24790) );
  XNOR U25023 ( .A(n24791), .B(n22668), .Z(n19496) );
  ANDN U25024 ( .B(n23372), .A(n23373), .Z(n24791) );
  XOR U25025 ( .A(n24792), .B(n24793), .Z(n24788) );
  XOR U25026 ( .A(n24209), .B(n18305), .Z(n24793) );
  XNOR U25027 ( .A(n24794), .B(n22659), .Z(n18305) );
  ANDN U25028 ( .B(n23377), .A(n23378), .Z(n24794) );
  XNOR U25029 ( .A(n24795), .B(n22663), .Z(n24209) );
  ANDN U25030 ( .B(n24796), .A(n24797), .Z(n24795) );
  XOR U25031 ( .A(n24798), .B(n24799), .Z(n21932) );
  XOR U25032 ( .A(n19170), .B(n23457), .Z(n24799) );
  XOR U25033 ( .A(n24800), .B(n22526), .Z(n23457) );
  ANDN U25034 ( .B(n24357), .A(n20406), .Z(n24800) );
  XOR U25035 ( .A(round_reg[58]), .B(n24578), .Z(n20406) );
  XNOR U25036 ( .A(n24801), .B(n22537), .Z(n19170) );
  ANDN U25037 ( .B(n24360), .A(n24359), .Z(n24801) );
  XNOR U25038 ( .A(round_reg[310]), .B(n22278), .Z(n24360) );
  XOR U25039 ( .A(n16038), .B(n24802), .Z(n24798) );
  XOR U25040 ( .A(n18860), .B(n19432), .Z(n24802) );
  XNOR U25041 ( .A(n24803), .B(n22535), .Z(n19432) );
  NOR U25042 ( .A(n20414), .B(n24352), .Z(n24803) );
  XOR U25043 ( .A(round_reg[198]), .B(n24218), .Z(n20414) );
  XNOR U25044 ( .A(n24804), .B(n22533), .Z(n18860) );
  ANDN U25045 ( .B(n24350), .A(n20410), .Z(n24804) );
  XOR U25046 ( .A(round_reg[80]), .B(n22445), .Z(n20410) );
  XOR U25047 ( .A(n24805), .B(n22529), .Z(n16038) );
  AND U25048 ( .A(n24362), .B(n24331), .Z(n24805) );
  IV U25049 ( .A(n24363), .Z(n24331) );
  XOR U25050 ( .A(round_reg[139]), .B(n24552), .Z(n24363) );
  XNOR U25051 ( .A(n24806), .B(n24796), .Z(n23375) );
  AND U25052 ( .A(n24797), .B(n22661), .Z(n24806) );
  XOR U25053 ( .A(n18063), .B(n24807), .Z(n24655) );
  XOR U25054 ( .A(n10784), .B(n10566), .Z(n24807) );
  XNOR U25055 ( .A(n24808), .B(n18067), .Z(n10566) );
  XNOR U25056 ( .A(n22131), .B(n17045), .Z(n18067) );
  XNOR U25057 ( .A(n23330), .B(n19681), .Z(n17045) );
  XNOR U25058 ( .A(n24809), .B(n24810), .Z(n19681) );
  XOR U25059 ( .A(n16349), .B(n24505), .Z(n24810) );
  XNOR U25060 ( .A(n24811), .B(n20476), .Z(n24505) );
  XOR U25061 ( .A(round_reg[291]), .B(n23256), .Z(n20476) );
  AND U25062 ( .A(n22117), .B(n21926), .Z(n24811) );
  IV U25063 ( .A(n22118), .Z(n21926) );
  XOR U25064 ( .A(round_reg[1135]), .B(n21196), .Z(n22118) );
  XOR U25065 ( .A(n24812), .B(n24813), .Z(n21196) );
  XOR U25066 ( .A(round_reg[1524]), .B(n22513), .Z(n22117) );
  XNOR U25067 ( .A(n24814), .B(n20488), .Z(n16349) );
  XNOR U25068 ( .A(round_reg[184]), .B(n22642), .Z(n20488) );
  ANDN U25069 ( .B(n22104), .A(n21623), .Z(n24814) );
  XNOR U25070 ( .A(round_reg[993]), .B(n24815), .Z(n21623) );
  XOR U25071 ( .A(round_reg[1369]), .B(n21760), .Z(n22104) );
  XOR U25072 ( .A(n24816), .B(n24817), .Z(n21760) );
  XNOR U25073 ( .A(n22697), .B(n24818), .Z(n24809) );
  XNOR U25074 ( .A(n17001), .B(n18833), .Z(n24818) );
  XOR U25075 ( .A(n24819), .B(n24524), .Z(n18833) );
  IV U25076 ( .A(n20472), .Z(n24524) );
  XNOR U25077 ( .A(round_reg[243]), .B(n24518), .Z(n20472) );
  AND U25078 ( .A(n21629), .B(n22114), .Z(n24819) );
  XOR U25079 ( .A(round_reg[1463]), .B(n24029), .Z(n22114) );
  XOR U25080 ( .A(round_reg[1086]), .B(n23561), .Z(n21629) );
  XNOR U25081 ( .A(n24820), .B(n20484), .Z(n17001) );
  XNOR U25082 ( .A(round_reg[125]), .B(n22764), .Z(n20484) );
  AND U25083 ( .A(n22111), .B(n21631), .Z(n24820) );
  XOR U25084 ( .A(round_reg[1233]), .B(n23778), .Z(n21631) );
  XOR U25085 ( .A(round_reg[1306]), .B(n24823), .Z(n22111) );
  XOR U25086 ( .A(n24824), .B(n24529), .Z(n22697) );
  IV U25087 ( .A(n20481), .Z(n24529) );
  XNOR U25088 ( .A(round_reg[39]), .B(n23799), .Z(n20481) );
  AND U25089 ( .A(n21625), .B(n22107), .Z(n24824) );
  XOR U25090 ( .A(round_reg[1589]), .B(n23467), .Z(n22107) );
  XNOR U25091 ( .A(round_reg[1161]), .B(n24727), .Z(n21625) );
  XOR U25092 ( .A(n24825), .B(n24826), .Z(n23330) );
  XOR U25093 ( .A(n23763), .B(n20793), .Z(n24826) );
  XOR U25094 ( .A(n24827), .B(n22319), .Z(n20793) );
  XOR U25095 ( .A(round_reg[733]), .B(n23418), .Z(n22319) );
  AND U25096 ( .A(n22139), .B(n22137), .Z(n24827) );
  XOR U25097 ( .A(round_reg[366]), .B(n24828), .Z(n22137) );
  XNOR U25098 ( .A(n24829), .B(n22313), .Z(n23763) );
  XOR U25099 ( .A(round_reg[876]), .B(n23726), .Z(n22313) );
  XOR U25100 ( .A(n19194), .B(n24831), .Z(n24825) );
  XOR U25101 ( .A(n18214), .B(n19963), .Z(n24831) );
  XNOR U25102 ( .A(n24832), .B(n22316), .Z(n19963) );
  XOR U25103 ( .A(round_reg[655]), .B(n23606), .Z(n22316) );
  ANDN U25104 ( .B(n22127), .A(n22128), .Z(n24832) );
  XOR U25105 ( .A(round_reg[589]), .B(n24214), .Z(n22127) );
  XNOR U25106 ( .A(n24833), .B(n22305), .Z(n18214) );
  XOR U25107 ( .A(round_reg[947]), .B(n21312), .Z(n22305) );
  AND U25108 ( .A(n22123), .B(n22125), .Z(n24833) );
  XOR U25109 ( .A(round_reg[521]), .B(n24727), .Z(n22123) );
  XNOR U25110 ( .A(n24834), .B(n22308), .Z(n19194) );
  XOR U25111 ( .A(round_reg[779]), .B(n24552), .Z(n22308) );
  AND U25112 ( .A(n22133), .B(n22135), .Z(n24834) );
  XOR U25113 ( .A(round_reg[417]), .B(n23780), .Z(n22133) );
  IV U25114 ( .A(n24320), .Z(n23780) );
  XNOR U25115 ( .A(n24835), .B(n23772), .Z(n22131) );
  XOR U25116 ( .A(round_reg[487]), .B(n21189), .Z(n23772) );
  ANDN U25117 ( .B(n24830), .A(n22311), .Z(n24835) );
  ANDN U25118 ( .B(n15872), .A(n15871), .Z(n24808) );
  XNOR U25119 ( .A(n20818), .B(n15208), .Z(n15871) );
  XNOR U25120 ( .A(n24836), .B(n24837), .Z(n19902) );
  XNOR U25121 ( .A(n17911), .B(n18189), .Z(n24837) );
  XNOR U25122 ( .A(n24838), .B(n22003), .Z(n18189) );
  ANDN U25123 ( .B(n20820), .A(n20821), .Z(n24838) );
  XNOR U25124 ( .A(round_reg[1597]), .B(n23242), .Z(n20821) );
  IV U25125 ( .A(n24440), .Z(n23242) );
  XOR U25126 ( .A(round_reg[47]), .B(n24564), .Z(n20820) );
  XOR U25127 ( .A(n24839), .B(n21999), .Z(n17911) );
  AND U25128 ( .A(n20814), .B(n20816), .Z(n24839) );
  XOR U25129 ( .A(round_reg[1532]), .B(n24840), .Z(n20816) );
  XOR U25130 ( .A(round_reg[299]), .B(n22375), .Z(n20814) );
  XOR U25131 ( .A(n24841), .B(n24842), .Z(n22375) );
  XOR U25132 ( .A(n18911), .B(n24843), .Z(n24836) );
  XNOR U25133 ( .A(n17523), .B(n17457), .Z(n24843) );
  XNOR U25134 ( .A(n24844), .B(n24845), .Z(n17457) );
  ANDN U25135 ( .B(n21997), .A(n21273), .Z(n24844) );
  XOR U25136 ( .A(n24846), .B(n24847), .Z(n17523) );
  ANDN U25137 ( .B(n23891), .A(n21266), .Z(n24846) );
  XOR U25138 ( .A(round_reg[1314]), .B(n23405), .Z(n21266) );
  XNOR U25139 ( .A(n24848), .B(n22005), .Z(n18911) );
  AND U25140 ( .A(n20824), .B(n21263), .Z(n24848) );
  XOR U25141 ( .A(round_reg[1377]), .B(n24320), .Z(n21263) );
  XNOR U25142 ( .A(n24849), .B(n24850), .Z(n24320) );
  XOR U25143 ( .A(round_reg[128]), .B(n23011), .Z(n20824) );
  XNOR U25144 ( .A(n24851), .B(n24852), .Z(n22077) );
  XOR U25145 ( .A(n15846), .B(n21792), .Z(n24852) );
  XNOR U25146 ( .A(n24853), .B(n22704), .Z(n21792) );
  NOR U25147 ( .A(n24677), .B(n22703), .Z(n24853) );
  XNOR U25148 ( .A(round_reg[1000]), .B(n24687), .Z(n22703) );
  IV U25149 ( .A(n22398), .Z(n24677) );
  XOR U25150 ( .A(round_reg[953]), .B(n23854), .Z(n22398) );
  XNOR U25151 ( .A(n24854), .B(n24855), .Z(n15846) );
  AND U25152 ( .A(n22402), .B(n21823), .Z(n24854) );
  XOR U25153 ( .A(round_reg[1168]), .B(n24229), .Z(n21823) );
  XNOR U25154 ( .A(round_reg[785]), .B(n22790), .Z(n22402) );
  XNOR U25155 ( .A(n21803), .B(n24856), .Z(n24851) );
  XOR U25156 ( .A(n15590), .B(n18745), .Z(n24856) );
  XNOR U25157 ( .A(n24857), .B(n24858), .Z(n18745) );
  AND U25158 ( .A(n24659), .B(n21809), .Z(n24857) );
  XOR U25159 ( .A(round_reg[1240]), .B(n23406), .Z(n21809) );
  XNOR U25160 ( .A(round_reg[882]), .B(n24859), .Z(n24659) );
  XNOR U25161 ( .A(n24860), .B(n21819), .Z(n15590) );
  ANDN U25162 ( .B(n21818), .A(n23212), .Z(n24860) );
  XNOR U25163 ( .A(round_reg[661]), .B(n24861), .Z(n23212) );
  XOR U25164 ( .A(round_reg[1029]), .B(n24559), .Z(n21818) );
  XNOR U25165 ( .A(n24862), .B(n21813), .Z(n21803) );
  NOR U25166 ( .A(n22393), .B(n21812), .Z(n24862) );
  XNOR U25167 ( .A(round_reg[1142]), .B(n24514), .Z(n21812) );
  XOR U25168 ( .A(round_reg[739]), .B(n21920), .Z(n22393) );
  XNOR U25169 ( .A(n24863), .B(n21997), .Z(n20818) );
  XNOR U25170 ( .A(round_reg[251]), .B(n21617), .Z(n21997) );
  ANDN U25171 ( .B(n21273), .A(n21274), .Z(n24863) );
  XOR U25172 ( .A(round_reg[1471]), .B(n23603), .Z(n21273) );
  XOR U25173 ( .A(n21564), .B(n16064), .Z(n15872) );
  IV U25174 ( .A(n19732), .Z(n16064) );
  XNOR U25175 ( .A(n24864), .B(n24865), .Z(n18748) );
  XNOR U25176 ( .A(n18404), .B(n18167), .Z(n24865) );
  XNOR U25177 ( .A(n24866), .B(n23202), .Z(n18167) );
  XOR U25178 ( .A(round_reg[201]), .B(n24727), .Z(n23202) );
  ANDN U25179 ( .B(n21571), .A(n20647), .Z(n24866) );
  XOR U25180 ( .A(round_reg[1044]), .B(n24155), .Z(n20647) );
  IV U25181 ( .A(n23141), .Z(n24155) );
  XOR U25182 ( .A(n24867), .B(n24868), .Z(n23141) );
  XNOR U25183 ( .A(round_reg[1421]), .B(n22652), .Z(n21571) );
  IV U25184 ( .A(n21306), .Z(n22652) );
  XNOR U25185 ( .A(round_reg[61]), .B(n24121), .Z(n23195) );
  ANDN U25186 ( .B(n24244), .A(n20656), .Z(n24869) );
  XOR U25187 ( .A(n18649), .B(n24870), .Z(n24864) );
  XOR U25188 ( .A(n21707), .B(n18714), .Z(n24870) );
  XNOR U25189 ( .A(n24871), .B(n23204), .Z(n18714) );
  XOR U25190 ( .A(round_reg[83]), .B(n21610), .Z(n23204) );
  IV U25191 ( .A(n24872), .Z(n21610) );
  ANDN U25192 ( .B(n21569), .A(n20660), .Z(n24871) );
  XOR U25193 ( .A(round_reg[1255]), .B(n23260), .Z(n20660) );
  XOR U25194 ( .A(round_reg[1328]), .B(n23445), .Z(n21569) );
  XNOR U25195 ( .A(n24873), .B(n23207), .Z(n21707) );
  XOR U25196 ( .A(round_reg[142]), .B(n23134), .Z(n23207) );
  NOR U25197 ( .A(n21566), .B(n20664), .Z(n24873) );
  XOR U25198 ( .A(round_reg[1015]), .B(n24715), .Z(n20664) );
  XNOR U25199 ( .A(round_reg[1391]), .B(n23262), .Z(n21566) );
  IV U25200 ( .A(n23241), .Z(n23262) );
  XNOR U25201 ( .A(n24874), .B(n23198), .Z(n18649) );
  XOR U25202 ( .A(round_reg[313]), .B(n24875), .Z(n23198) );
  ANDN U25203 ( .B(n20651), .A(n21573), .Z(n24874) );
  XNOR U25204 ( .A(round_reg[1482]), .B(n22366), .Z(n21573) );
  XNOR U25205 ( .A(round_reg[1093]), .B(n22365), .Z(n20651) );
  XNOR U25206 ( .A(n24876), .B(n24877), .Z(n22653) );
  XOR U25207 ( .A(n18737), .B(n24654), .Z(n24877) );
  XNOR U25208 ( .A(n24878), .B(n19100), .Z(n24654) );
  ANDN U25209 ( .B(n21782), .A(n20636), .Z(n24878) );
  XOR U25210 ( .A(round_reg[609]), .B(n23745), .Z(n20636) );
  XNOR U25211 ( .A(n24879), .B(n19093), .Z(n18737) );
  ANDN U25212 ( .B(n21774), .A(n20641), .Z(n24879) );
  XOR U25213 ( .A(round_reg[322]), .B(n22442), .Z(n20641) );
  XOR U25214 ( .A(n24880), .B(n24881), .Z(n22442) );
  XOR U25215 ( .A(n20629), .B(n24882), .Z(n24876) );
  XOR U25216 ( .A(n18017), .B(n24883), .Z(n24882) );
  XOR U25217 ( .A(n24884), .B(n19090), .Z(n18017) );
  IV U25218 ( .A(n24885), .Z(n19090) );
  ANDN U25219 ( .B(n21779), .A(n21780), .Z(n24884) );
  XOR U25220 ( .A(round_reg[507]), .B(n23250), .Z(n21780) );
  XNOR U25221 ( .A(n24886), .B(n19693), .Z(n20629) );
  ANDN U25222 ( .B(n22651), .A(n20643), .Z(n24886) );
  XOR U25223 ( .A(round_reg[541]), .B(n24887), .Z(n20643) );
  XNOR U25224 ( .A(n24888), .B(n24244), .Z(n21564) );
  XOR U25225 ( .A(round_reg[1547]), .B(n24704), .Z(n24244) );
  XOR U25226 ( .A(round_reg[800]), .B(n23244), .Z(n20658) );
  XOR U25227 ( .A(round_reg[1183]), .B(n24769), .Z(n20656) );
  XNOR U25228 ( .A(n24889), .B(n18069), .Z(n10784) );
  XOR U25229 ( .A(n21588), .B(n17467), .Z(n18069) );
  XOR U25230 ( .A(n20248), .B(n24890), .Z(n17467) );
  XOR U25231 ( .A(n24891), .B(n24892), .Z(n20248) );
  XNOR U25232 ( .A(n24586), .B(n18153), .Z(n24892) );
  XNOR U25233 ( .A(n24893), .B(n21387), .Z(n18153) );
  XOR U25234 ( .A(round_reg[500]), .B(n22230), .Z(n21387) );
  XNOR U25235 ( .A(n24895), .B(n21379), .Z(n24586) );
  XOR U25236 ( .A(round_reg[379]), .B(n22986), .Z(n21379) );
  XNOR U25237 ( .A(n24897), .B(n24898), .Z(n23829) );
  XNOR U25238 ( .A(round_reg[1329]), .B(round_reg[1009]), .Z(n24898) );
  XOR U25239 ( .A(round_reg[369]), .B(n24899), .Z(n24897) );
  XOR U25240 ( .A(round_reg[689]), .B(round_reg[49]), .Z(n24899) );
  XOR U25241 ( .A(n23022), .B(n24900), .Z(n24891) );
  XOR U25242 ( .A(n15902), .B(n19895), .Z(n24900) );
  XNOR U25243 ( .A(n24901), .B(n21374), .Z(n19895) );
  XOR U25244 ( .A(round_reg[602]), .B(n22640), .Z(n21374) );
  ANDN U25245 ( .B(n22386), .A(n22387), .Z(n24901) );
  XNOR U25246 ( .A(round_reg[193]), .B(n22211), .Z(n22386) );
  XNOR U25247 ( .A(n24902), .B(n21383), .Z(n15902) );
  XOR U25248 ( .A(round_reg[430]), .B(n22825), .Z(n21383) );
  ANDN U25249 ( .B(n21593), .A(n21594), .Z(n24902) );
  XNOR U25250 ( .A(round_reg[53]), .B(n21313), .Z(n21593) );
  XOR U25251 ( .A(n24903), .B(n21370), .Z(n23022) );
  XOR U25252 ( .A(round_reg[534]), .B(n24904), .Z(n21370) );
  NOR U25253 ( .A(n21586), .B(n21585), .Z(n24903) );
  XOR U25254 ( .A(round_reg[134]), .B(n24397), .Z(n21585) );
  XNOR U25255 ( .A(n24905), .B(n24603), .Z(n21588) );
  XOR U25256 ( .A(round_reg[75]), .B(n24906), .Z(n24603) );
  ANDN U25257 ( .B(n24894), .A(n21385), .Z(n24905) );
  XNOR U25258 ( .A(n24883), .B(n18018), .Z(n15878) );
  XNOR U25259 ( .A(n21708), .B(n20396), .Z(n18018) );
  XNOR U25260 ( .A(n24907), .B(n24908), .Z(n20396) );
  XNOR U25261 ( .A(n18157), .B(n20016), .Z(n24908) );
  XNOR U25262 ( .A(n24909), .B(n23381), .Z(n20016) );
  AND U25263 ( .A(n22672), .B(n22670), .Z(n24909) );
  XNOR U25264 ( .A(round_reg[321]), .B(n22966), .Z(n22670) );
  IV U25265 ( .A(n21602), .Z(n22966) );
  XOR U25266 ( .A(n24910), .B(n24911), .Z(n21602) );
  XNOR U25267 ( .A(n24912), .B(n23378), .Z(n18157) );
  XOR U25268 ( .A(round_reg[895]), .B(n23904), .Z(n23378) );
  ANDN U25269 ( .B(n22657), .A(n22658), .Z(n24912) );
  XNOR U25270 ( .A(round_reg[506]), .B(n24451), .Z(n22657) );
  XOR U25271 ( .A(n21135), .B(n24913), .Z(n24907) );
  XOR U25272 ( .A(n19243), .B(n23364), .Z(n24913) );
  XNOR U25273 ( .A(n24914), .B(n24797), .Z(n23364) );
  XOR U25274 ( .A(round_reg[674]), .B(n23405), .Z(n24797) );
  XNOR U25275 ( .A(round_reg[608]), .B(n24272), .Z(n22661) );
  XNOR U25276 ( .A(n24915), .B(n23370), .Z(n19243) );
  XOR U25277 ( .A(round_reg[902]), .B(n23607), .Z(n23370) );
  XNOR U25278 ( .A(round_reg[540]), .B(n23253), .Z(n22674) );
  XNOR U25279 ( .A(n24916), .B(n23373), .Z(n21135) );
  XOR U25280 ( .A(round_reg[798]), .B(n21923), .Z(n23373) );
  XOR U25281 ( .A(n24917), .B(n24918), .Z(n23289) );
  XOR U25282 ( .A(n24919), .B(n24920), .Z(n21708) );
  XOR U25283 ( .A(n19083), .B(n18481), .Z(n24920) );
  XOR U25284 ( .A(n24921), .B(n19692), .Z(n18481) );
  XOR U25285 ( .A(round_reg[1390]), .B(n22825), .Z(n19692) );
  XNOR U25286 ( .A(n24565), .B(n24689), .Z(n22825) );
  XNOR U25287 ( .A(n24922), .B(n24923), .Z(n24689) );
  XNOR U25288 ( .A(round_reg[1454]), .B(round_reg[1134]), .Z(n24923) );
  XOR U25289 ( .A(round_reg[174]), .B(n24924), .Z(n24922) );
  XOR U25290 ( .A(round_reg[814]), .B(round_reg[494]), .Z(n24924) );
  XNOR U25291 ( .A(n24925), .B(n24926), .Z(n24565) );
  XNOR U25292 ( .A(round_reg[1325]), .B(round_reg[1005]), .Z(n24926) );
  XOR U25293 ( .A(round_reg[365]), .B(n24927), .Z(n24925) );
  XOR U25294 ( .A(round_reg[685]), .B(round_reg[45]), .Z(n24927) );
  ANDN U25295 ( .B(n19693), .A(n22651), .Z(n24921) );
  XOR U25296 ( .A(round_reg[903]), .B(n23916), .Z(n22651) );
  XOR U25297 ( .A(n24928), .B(n24929), .Z(n23916) );
  XOR U25298 ( .A(round_reg[1014]), .B(n23879), .Z(n19693) );
  XNOR U25299 ( .A(n24930), .B(n19103), .Z(n19083) );
  XOR U25300 ( .A(round_reg[1546]), .B(n24377), .Z(n19103) );
  ANDN U25301 ( .B(n19104), .A(n21771), .Z(n24930) );
  XOR U25302 ( .A(n16477), .B(n24931), .Z(n24919) );
  XOR U25303 ( .A(n16546), .B(n18667), .Z(n24931) );
  XNOR U25304 ( .A(n24932), .B(n19089), .Z(n18667) );
  XOR U25305 ( .A(round_reg[1327]), .B(n24564), .Z(n19089) );
  ANDN U25306 ( .B(n24885), .A(n21779), .Z(n24932) );
  XOR U25307 ( .A(round_reg[832]), .B(n24163), .Z(n21779) );
  IV U25308 ( .A(n23991), .Z(n24163) );
  XNOR U25309 ( .A(n24934), .B(n24935), .Z(n24911) );
  XNOR U25310 ( .A(round_reg[1536]), .B(round_reg[1216]), .Z(n24935) );
  XOR U25311 ( .A(round_reg[256]), .B(n24936), .Z(n24934) );
  XOR U25312 ( .A(round_reg[896]), .B(round_reg[576]), .Z(n24936) );
  XNOR U25313 ( .A(round_reg[1254]), .B(n22432), .Z(n24885) );
  XNOR U25314 ( .A(n24937), .B(n19099), .Z(n16546) );
  XOR U25315 ( .A(round_reg[1420]), .B(n24389), .Z(n19099) );
  ANDN U25316 ( .B(n19100), .A(n21782), .Z(n24937) );
  XOR U25317 ( .A(round_reg[675]), .B(n23584), .Z(n21782) );
  XNOR U25318 ( .A(round_reg[1043]), .B(n24872), .Z(n19100) );
  XNOR U25319 ( .A(n24940), .B(n19094), .Z(n16477) );
  XOR U25320 ( .A(round_reg[1481]), .B(n24727), .Z(n19094) );
  NOR U25321 ( .A(n21774), .B(n19093), .Z(n24940) );
  XNOR U25322 ( .A(round_reg[1092]), .B(n24728), .Z(n19093) );
  XOR U25323 ( .A(round_reg[753]), .B(n24943), .Z(n21774) );
  XNOR U25324 ( .A(n24944), .B(n19104), .Z(n24883) );
  ANDN U25325 ( .B(n21771), .A(n20639), .Z(n24944) );
  XOR U25326 ( .A(round_reg[437]), .B(n23993), .Z(n20639) );
  XNOR U25327 ( .A(round_reg[799]), .B(n24460), .Z(n21771) );
  XNOR U25328 ( .A(n17993), .B(n20768), .Z(n15876) );
  XNOR U25329 ( .A(n24945), .B(n20506), .Z(n20768) );
  ANDN U25330 ( .B(n22264), .A(n19826), .Z(n24945) );
  XOR U25331 ( .A(round_reg[658]), .B(n21186), .Z(n19826) );
  XNOR U25332 ( .A(n19631), .B(n18908), .Z(n17993) );
  XOR U25333 ( .A(n24946), .B(n24947), .Z(n18908) );
  XOR U25334 ( .A(n15121), .B(n20202), .Z(n24947) );
  XNOR U25335 ( .A(n24948), .B(n19838), .Z(n20202) );
  XNOR U25336 ( .A(round_reg[65]), .B(n24547), .Z(n19838) );
  IV U25337 ( .A(n24466), .Z(n24547) );
  ANDN U25338 ( .B(n20508), .A(n20944), .Z(n24948) );
  XNOR U25339 ( .A(round_reg[1237]), .B(n24327), .Z(n20944) );
  IV U25340 ( .A(n23266), .Z(n24327) );
  XOR U25341 ( .A(n24718), .B(n24949), .Z(n23266) );
  XNOR U25342 ( .A(n24950), .B(n24951), .Z(n24718) );
  XNOR U25343 ( .A(round_reg[1492]), .B(round_reg[1172]), .Z(n24951) );
  XOR U25344 ( .A(round_reg[212]), .B(n24952), .Z(n24950) );
  XOR U25345 ( .A(round_reg[852]), .B(round_reg[532]), .Z(n24952) );
  XOR U25346 ( .A(round_reg[1310]), .B(n23246), .Z(n20508) );
  XNOR U25347 ( .A(n24953), .B(n19832), .Z(n15121) );
  XOR U25348 ( .A(round_reg[295]), .B(n23260), .Z(n19832) );
  XOR U25349 ( .A(n24954), .B(n24955), .Z(n23260) );
  ANDN U25350 ( .B(n20773), .A(n20503), .Z(n24953) );
  XNOR U25351 ( .A(round_reg[1528]), .B(n23777), .Z(n20503) );
  XNOR U25352 ( .A(round_reg[1139]), .B(n23621), .Z(n20773) );
  XNOR U25353 ( .A(n16474), .B(n24956), .Z(n24946) );
  XOR U25354 ( .A(n17162), .B(n18693), .Z(n24956) );
  XNOR U25355 ( .A(n24957), .B(n20501), .Z(n18693) );
  XNOR U25356 ( .A(round_reg[43]), .B(n24302), .Z(n20501) );
  NOR U25357 ( .A(n23133), .B(n20500), .Z(n24957) );
  XNOR U25358 ( .A(round_reg[1593]), .B(n24875), .Z(n20500) );
  IV U25359 ( .A(n22271), .Z(n23133) );
  XOR U25360 ( .A(round_reg[1165]), .B(n23489), .Z(n22271) );
  IV U25361 ( .A(n23502), .Z(n23489) );
  XOR U25362 ( .A(n24958), .B(n24959), .Z(n23502) );
  XNOR U25363 ( .A(n24960), .B(n19828), .Z(n17162) );
  XNOR U25364 ( .A(round_reg[247]), .B(n23127), .Z(n19828) );
  ANDN U25365 ( .B(n20506), .A(n22264), .Z(n24960) );
  XNOR U25366 ( .A(round_reg[1026]), .B(n23787), .Z(n22264) );
  XOR U25367 ( .A(round_reg[1467]), .B(n23250), .Z(n20506) );
  XNOR U25368 ( .A(n24961), .B(n20512), .Z(n16474) );
  XNOR U25369 ( .A(round_reg[188]), .B(n23323), .Z(n20512) );
  ANDN U25370 ( .B(n22276), .A(n20511), .Z(n24961) );
  XNOR U25371 ( .A(round_reg[1373]), .B(n23418), .Z(n20511) );
  IV U25372 ( .A(n24962), .Z(n23418) );
  IV U25373 ( .A(n20775), .Z(n22276) );
  XOR U25374 ( .A(round_reg[997]), .B(n24157), .Z(n20775) );
  XOR U25375 ( .A(n24963), .B(n24964), .Z(n19631) );
  XNOR U25376 ( .A(n19022), .B(n19590), .Z(n24964) );
  XOR U25377 ( .A(n24965), .B(n23232), .Z(n19590) );
  XNOR U25378 ( .A(round_reg[1025]), .B(n24466), .Z(n23232) );
  XNOR U25379 ( .A(n24966), .B(n24967), .Z(n24466) );
  ANDN U25380 ( .B(n22483), .A(n22484), .Z(n24965) );
  XOR U25381 ( .A(round_reg[657]), .B(n22829), .Z(n22483) );
  XNOR U25382 ( .A(n24968), .B(n23235), .Z(n19022) );
  XNOR U25383 ( .A(round_reg[1138]), .B(n24692), .Z(n23235) );
  ANDN U25384 ( .B(n22487), .A(n22488), .Z(n24968) );
  XOR U25385 ( .A(round_reg[735]), .B(n24673), .Z(n22487) );
  IV U25386 ( .A(n23670), .Z(n24673) );
  XOR U25387 ( .A(n24969), .B(n24970), .Z(n23670) );
  XNOR U25388 ( .A(n19333), .B(n24971), .Z(n24963) );
  XNOR U25389 ( .A(n18764), .B(n23218), .Z(n24971) );
  XNOR U25390 ( .A(n24972), .B(n23225), .Z(n23218) );
  XNOR U25391 ( .A(round_reg[1164]), .B(n22279), .Z(n23225) );
  ANDN U25392 ( .B(n22494), .A(n22492), .Z(n24972) );
  XNOR U25393 ( .A(round_reg[781]), .B(n21306), .Z(n22492) );
  XNOR U25394 ( .A(n24975), .B(n23229), .Z(n18764) );
  XNOR U25395 ( .A(round_reg[1236]), .B(n22818), .Z(n23229) );
  ANDN U25396 ( .B(n22496), .A(n22497), .Z(n24975) );
  XOR U25397 ( .A(n24976), .B(n24977), .Z(n23735) );
  XNOR U25398 ( .A(n24978), .B(n24630), .Z(n19333) );
  NOR U25399 ( .A(n22502), .B(n22500), .Z(n24978) );
  XNOR U25400 ( .A(round_reg[949]), .B(n23467), .Z(n22500) );
  XOR U25401 ( .A(n24979), .B(n19065), .Z(n18063) );
  IV U25402 ( .A(n18075), .Z(n19065) );
  XNOR U25403 ( .A(n15917), .B(n24474), .Z(n18075) );
  XNOR U25404 ( .A(n24980), .B(n21449), .Z(n24474) );
  AND U25405 ( .A(n24981), .B(n23842), .Z(n24980) );
  IV U25406 ( .A(n24982), .Z(n23842) );
  XNOR U25407 ( .A(n21078), .B(n23209), .Z(n15917) );
  XNOR U25408 ( .A(n24983), .B(n24984), .Z(n23209) );
  XOR U25409 ( .A(n19651), .B(n17148), .Z(n24984) );
  XOR U25410 ( .A(n24985), .B(n21457), .Z(n17148) );
  XOR U25411 ( .A(round_reg[694]), .B(n23879), .Z(n21457) );
  IV U25412 ( .A(n24986), .Z(n23879) );
  AND U25413 ( .A(n21105), .B(n21458), .Z(n24985) );
  XOR U25414 ( .A(round_reg[628]), .B(n24084), .Z(n21458) );
  XNOR U25415 ( .A(round_reg[219]), .B(n24342), .Z(n21105) );
  XNOR U25416 ( .A(n24987), .B(n21461), .Z(n19651) );
  XOR U25417 ( .A(round_reg[708]), .B(n23721), .Z(n21461) );
  AND U25418 ( .A(n21110), .B(n21462), .Z(n24987) );
  XOR U25419 ( .A(round_reg[341]), .B(n23393), .Z(n21462) );
  XNOR U25420 ( .A(round_reg[267]), .B(n24704), .Z(n21110) );
  XOR U25421 ( .A(n19382), .B(n24988), .Z(n24983) );
  XOR U25422 ( .A(n19126), .B(n18129), .Z(n24988) );
  XNOR U25423 ( .A(n24989), .B(n21468), .Z(n18129) );
  XOR U25424 ( .A(round_reg[818]), .B(n24692), .Z(n21468) );
  ANDN U25425 ( .B(n21469), .A(n21101), .Z(n24989) );
  XOR U25426 ( .A(round_reg[15]), .B(n23606), .Z(n21101) );
  XOR U25427 ( .A(round_reg[392]), .B(n24284), .Z(n21469) );
  XNOR U25428 ( .A(n24990), .B(n21465), .Z(n19126) );
  XOR U25429 ( .A(round_reg[851]), .B(n24288), .Z(n21465) );
  ANDN U25430 ( .B(n21466), .A(n21114), .Z(n24990) );
  XNOR U25431 ( .A(round_reg[101]), .B(n24374), .Z(n21114) );
  XNOR U25432 ( .A(n24991), .B(n24992), .Z(n24374) );
  XOR U25433 ( .A(round_reg[462]), .B(n23134), .Z(n21466) );
  XNOR U25434 ( .A(n24993), .B(n21471), .Z(n19382) );
  XOR U25435 ( .A(round_reg[922]), .B(n22640), .Z(n21471) );
  IV U25436 ( .A(n23564), .Z(n22640) );
  XNOR U25437 ( .A(n24994), .B(n24995), .Z(n23564) );
  ANDN U25438 ( .B(n21472), .A(n21118), .Z(n24993) );
  XNOR U25439 ( .A(round_reg[160]), .B(n24996), .Z(n21118) );
  XOR U25440 ( .A(round_reg[560]), .B(n23618), .Z(n21472) );
  XOR U25441 ( .A(n24997), .B(n24998), .Z(n21078) );
  XOR U25442 ( .A(n20097), .B(n19019), .Z(n24998) );
  XNOR U25443 ( .A(n24999), .B(n21453), .Z(n19019) );
  XNOR U25444 ( .A(round_reg[1346]), .B(n24132), .Z(n21453) );
  IV U25445 ( .A(n23787), .Z(n24132) );
  XOR U25446 ( .A(n25000), .B(n24724), .Z(n23787) );
  XOR U25447 ( .A(n25001), .B(n25002), .Z(n24724) );
  XNOR U25448 ( .A(round_reg[1]), .B(round_reg[1281]), .Z(n25002) );
  XOR U25449 ( .A(round_reg[321]), .B(n25003), .Z(n25001) );
  XOR U25450 ( .A(round_reg[961]), .B(round_reg[641]), .Z(n25003) );
  AND U25451 ( .A(n21452), .B(n25004), .Z(n24999) );
  XOR U25452 ( .A(round_reg[970]), .B(n24116), .Z(n21452) );
  XNOR U25453 ( .A(n25005), .B(n21442), .Z(n20097) );
  XOR U25454 ( .A(round_reg[1440]), .B(n23244), .Z(n21442) );
  IV U25455 ( .A(n24996), .Z(n23244) );
  AND U25456 ( .A(n24470), .B(n21443), .Z(n25005) );
  XOR U25457 ( .A(round_reg[1063]), .B(n24450), .Z(n21443) );
  XNOR U25458 ( .A(n21436), .B(n25006), .Z(n24997) );
  XNOR U25459 ( .A(n20845), .B(n17961), .Z(n25006) );
  XOR U25460 ( .A(n25007), .B(n23187), .Z(n17961) );
  XOR U25461 ( .A(round_reg[1566]), .B(n25008), .Z(n23187) );
  ANDN U25462 ( .B(n23186), .A(n24476), .Z(n25007) );
  XOR U25463 ( .A(round_reg[1202]), .B(n24859), .Z(n23186) );
  XNOR U25464 ( .A(n25009), .B(n23838), .Z(n20845) );
  XNOR U25465 ( .A(round_reg[1501]), .B(n24887), .Z(n23838) );
  AND U25466 ( .A(n23859), .B(n25010), .Z(n25009) );
  XOR U25467 ( .A(round_reg[1112]), .B(n22980), .Z(n23859) );
  IV U25468 ( .A(n25011), .Z(n22980) );
  XOR U25469 ( .A(n25012), .B(n21448), .Z(n21436) );
  XNOR U25470 ( .A(round_reg[1283]), .B(n23599), .Z(n21448) );
  ANDN U25471 ( .B(n21449), .A(n24981), .Z(n25012) );
  XOR U25472 ( .A(round_reg[1274]), .B(n23318), .Z(n21449) );
  AND U25473 ( .A(n15886), .B(n15884), .Z(n24979) );
  XNOR U25474 ( .A(n16663), .B(n23813), .Z(n15884) );
  XNOR U25475 ( .A(n25015), .B(n22919), .Z(n23813) );
  ANDN U25476 ( .B(n23576), .A(n23499), .Z(n25015) );
  XNOR U25477 ( .A(round_reg[204]), .B(n25016), .Z(n23499) );
  IV U25478 ( .A(n18701), .Z(n16663) );
  XOR U25479 ( .A(n19928), .B(n24108), .Z(n18701) );
  XOR U25480 ( .A(n25017), .B(n25018), .Z(n24108) );
  XOR U25481 ( .A(n19430), .B(n20882), .Z(n25018) );
  XOR U25482 ( .A(n25019), .B(n24632), .Z(n20882) );
  XOR U25483 ( .A(round_reg[510]), .B(n22435), .Z(n24632) );
  ANDN U25484 ( .B(n23825), .A(n22873), .Z(n25019) );
  XOR U25485 ( .A(round_reg[1330]), .B(n23781), .Z(n22873) );
  XOR U25486 ( .A(round_reg[85]), .B(n23409), .Z(n23825) );
  XOR U25487 ( .A(n25020), .B(n25021), .Z(n23409) );
  XOR U25488 ( .A(n25022), .B(n24781), .Z(n19430) );
  IV U25489 ( .A(n22906), .Z(n24781) );
  XOR U25490 ( .A(round_reg[612]), .B(n25023), .Z(n22906) );
  ANDN U25491 ( .B(n22907), .A(n22860), .Z(n25022) );
  XOR U25492 ( .A(round_reg[1423]), .B(n23784), .Z(n22860) );
  XOR U25493 ( .A(round_reg[203]), .B(n24767), .Z(n22907) );
  XOR U25494 ( .A(n18809), .B(n25024), .Z(n25017) );
  XOR U25495 ( .A(n16778), .B(n16914), .Z(n25024) );
  XOR U25496 ( .A(n25025), .B(n24785), .Z(n16914) );
  XOR U25497 ( .A(round_reg[440]), .B(n24642), .Z(n24785) );
  ANDN U25498 ( .B(n23821), .A(n22869), .Z(n25025) );
  XOR U25499 ( .A(round_reg[1549]), .B(n24214), .Z(n22869) );
  XOR U25500 ( .A(round_reg[63]), .B(n22783), .Z(n23821) );
  XOR U25501 ( .A(n25026), .B(n25027), .Z(n22783) );
  XOR U25502 ( .A(n25028), .B(n22913), .Z(n16778) );
  XOR U25503 ( .A(round_reg[325]), .B(n25029), .Z(n22913) );
  ANDN U25504 ( .B(n22912), .A(n22864), .Z(n25028) );
  XOR U25505 ( .A(round_reg[1484]), .B(n22279), .Z(n22864) );
  IV U25506 ( .A(n25016), .Z(n22279) );
  XNOR U25507 ( .A(n25030), .B(n25031), .Z(n25016) );
  XOR U25508 ( .A(round_reg[315]), .B(n22517), .Z(n22912) );
  XOR U25509 ( .A(n25032), .B(n22903), .Z(n18809) );
  XOR U25510 ( .A(round_reg[544]), .B(n23608), .Z(n22903) );
  IV U25511 ( .A(n24254), .Z(n23608) );
  XOR U25512 ( .A(n24969), .B(n25033), .Z(n24254) );
  XOR U25513 ( .A(n25034), .B(n25035), .Z(n24969) );
  XNOR U25514 ( .A(round_reg[1439]), .B(round_reg[1119]), .Z(n25035) );
  XOR U25515 ( .A(round_reg[159]), .B(n25036), .Z(n25034) );
  XOR U25516 ( .A(round_reg[799]), .B(round_reg[479]), .Z(n25036) );
  ANDN U25517 ( .B(n22902), .A(n22877), .Z(n25032) );
  XOR U25518 ( .A(round_reg[1393]), .B(n24943), .Z(n22877) );
  XOR U25519 ( .A(round_reg[144]), .B(n23577), .Z(n22902) );
  XNOR U25520 ( .A(n25037), .B(n25038), .Z(n19928) );
  XNOR U25521 ( .A(n18528), .B(n22591), .Z(n25038) );
  XNOR U25522 ( .A(n25039), .B(n22918), .Z(n22591) );
  XOR U25523 ( .A(round_reg[1047]), .B(n23486), .Z(n22918) );
  XOR U25524 ( .A(n25040), .B(n25041), .Z(n23486) );
  ANDN U25525 ( .B(n22919), .A(n23576), .Z(n25039) );
  XOR U25526 ( .A(round_reg[613]), .B(n25042), .Z(n23576) );
  XOR U25527 ( .A(round_reg[679]), .B(n23799), .Z(n22919) );
  XOR U25528 ( .A(n25043), .B(n22923), .Z(n18528) );
  XNOR U25529 ( .A(round_reg[1096]), .B(n24134), .Z(n22923) );
  ANDN U25530 ( .B(n22922), .A(n22952), .Z(n25043) );
  XOR U25531 ( .A(round_reg[326]), .B(n23738), .Z(n22952) );
  XOR U25532 ( .A(round_reg[757]), .B(n23993), .Z(n22922) );
  XOR U25533 ( .A(n25044), .B(n25045), .Z(n23993) );
  XOR U25534 ( .A(n22898), .B(n25046), .Z(n25037) );
  XOR U25535 ( .A(n19242), .B(n19898), .Z(n25046) );
  XNOR U25536 ( .A(n25047), .B(n22931), .Z(n19898) );
  XNOR U25537 ( .A(round_reg[1258]), .B(n24738), .Z(n22931) );
  ANDN U25538 ( .B(n22932), .A(n22944), .Z(n25047) );
  XOR U25539 ( .A(round_reg[511]), .B(n23603), .Z(n22944) );
  XNOR U25540 ( .A(round_reg[836]), .B(n24405), .Z(n22932) );
  XOR U25541 ( .A(n25048), .B(n23496), .Z(n19242) );
  IV U25542 ( .A(n22927), .Z(n23496) );
  XOR U25543 ( .A(round_reg[1186]), .B(n23480), .Z(n22927) );
  ANDN U25544 ( .B(n22928), .A(n22949), .Z(n25048) );
  XOR U25545 ( .A(round_reg[441]), .B(n23623), .Z(n22949) );
  XOR U25546 ( .A(round_reg[803]), .B(n23396), .Z(n22928) );
  XOR U25547 ( .A(n25049), .B(n23507), .Z(n22898) );
  IV U25548 ( .A(n22935), .Z(n23507) );
  XOR U25549 ( .A(round_reg[1018]), .B(n24578), .Z(n22935) );
  ANDN U25550 ( .B(n22936), .A(n23809), .Z(n25049) );
  XOR U25551 ( .A(round_reg[545]), .B(n24752), .Z(n23809) );
  IV U25552 ( .A(n23019), .Z(n24752) );
  XOR U25553 ( .A(round_reg[907]), .B(n24704), .Z(n22936) );
  IV U25554 ( .A(n24022), .Z(n24704) );
  XNOR U25555 ( .A(n24354), .B(n25050), .Z(n24022) );
  XOR U25556 ( .A(n25051), .B(n25052), .Z(n24354) );
  XNOR U25557 ( .A(round_reg[1482]), .B(round_reg[1162]), .Z(n25052) );
  XOR U25558 ( .A(round_reg[202]), .B(n25053), .Z(n25051) );
  XOR U25559 ( .A(round_reg[842]), .B(round_reg[522]), .Z(n25053) );
  XOR U25560 ( .A(n24068), .B(n18801), .Z(n15886) );
  IV U25561 ( .A(n15954), .Z(n18801) );
  XNOR U25562 ( .A(n24411), .B(n18855), .Z(n15954) );
  XNOR U25563 ( .A(n25054), .B(n25055), .Z(n18855) );
  XNOR U25564 ( .A(n17942), .B(n20613), .Z(n25055) );
  XNOR U25565 ( .A(n25056), .B(n21210), .Z(n20613) );
  XNOR U25566 ( .A(round_reg[118]), .B(n23491), .Z(n21210) );
  XNOR U25567 ( .A(n25057), .B(n25058), .Z(n23491) );
  AND U25568 ( .A(n24148), .B(n24147), .Z(n25056) );
  XOR U25569 ( .A(round_reg[1299]), .B(n23744), .Z(n24147) );
  XNOR U25570 ( .A(round_reg[1226]), .B(n24377), .Z(n24148) );
  XOR U25571 ( .A(n25059), .B(n22203), .Z(n17942) );
  XOR U25572 ( .A(round_reg[284]), .B(n24372), .Z(n22203) );
  AND U25573 ( .A(n20224), .B(n22202), .Z(n25059) );
  XOR U25574 ( .A(round_reg[1517]), .B(n24309), .Z(n22202) );
  XNOR U25575 ( .A(round_reg[1128]), .B(n22821), .Z(n20224) );
  XOR U25576 ( .A(n19486), .B(n25060), .Z(n25054) );
  XOR U25577 ( .A(n17259), .B(n19010), .Z(n25060) );
  XNOR U25578 ( .A(n25061), .B(n21214), .Z(n19010) );
  XOR U25579 ( .A(round_reg[177]), .B(n24285), .Z(n21214) );
  ANDN U25580 ( .B(n22212), .A(n20210), .Z(n25061) );
  XOR U25581 ( .A(round_reg[986]), .B(n24823), .Z(n20210) );
  XNOR U25582 ( .A(round_reg[1362]), .B(n25062), .Z(n22212) );
  XNOR U25583 ( .A(n25063), .B(n21203), .Z(n17259) );
  XOR U25584 ( .A(round_reg[236]), .B(n23726), .Z(n21203) );
  XNOR U25585 ( .A(n25065), .B(n25066), .Z(n24665) );
  XNOR U25586 ( .A(round_reg[1580]), .B(round_reg[1260]), .Z(n25066) );
  XOR U25587 ( .A(round_reg[300]), .B(n25067), .Z(n25065) );
  XOR U25588 ( .A(round_reg[940]), .B(round_reg[620]), .Z(n25067) );
  ANDN U25589 ( .B(n22207), .A(n20220), .Z(n25063) );
  XOR U25590 ( .A(round_reg[1079]), .B(n24223), .Z(n20220) );
  XNOR U25591 ( .A(round_reg[1456]), .B(n25068), .Z(n22207) );
  XNOR U25592 ( .A(n25069), .B(n21212), .Z(n19486) );
  XOR U25593 ( .A(round_reg[32]), .B(n21606), .Z(n21212) );
  XOR U25594 ( .A(n25070), .B(n25071), .Z(n21606) );
  AND U25595 ( .A(n20214), .B(n22199), .Z(n25069) );
  XNOR U25596 ( .A(round_reg[1582]), .B(n24404), .Z(n22199) );
  XOR U25597 ( .A(n25072), .B(n25073), .Z(n24404) );
  XNOR U25598 ( .A(round_reg[1154]), .B(n25074), .Z(n20214) );
  XOR U25599 ( .A(n25075), .B(n25076), .Z(n24411) );
  XNOR U25600 ( .A(n18103), .B(n19130), .Z(n25076) );
  XOR U25601 ( .A(n25077), .B(n22182), .Z(n19130) );
  XOR U25602 ( .A(round_reg[648]), .B(n22977), .Z(n22182) );
  IV U25603 ( .A(n25078), .Z(n22977) );
  NOR U25604 ( .A(n22181), .B(n23687), .Z(n25077) );
  XOR U25605 ( .A(round_reg[237]), .B(n24309), .Z(n23687) );
  XOR U25606 ( .A(round_reg[582]), .B(n23538), .Z(n22181) );
  IV U25607 ( .A(n23607), .Z(n23538) );
  XOR U25608 ( .A(n25079), .B(n25080), .Z(n23607) );
  XOR U25609 ( .A(n25081), .B(n22191), .Z(n18103) );
  XOR U25610 ( .A(round_reg[726]), .B(n25082), .Z(n22191) );
  NOR U25611 ( .A(n22190), .B(n23683), .Z(n25081) );
  XOR U25612 ( .A(round_reg[285]), .B(n24171), .Z(n23683) );
  XNOR U25613 ( .A(round_reg[359]), .B(n23799), .Z(n22190) );
  XOR U25614 ( .A(n18975), .B(n25083), .Z(n25075) );
  XNOR U25615 ( .A(n22172), .B(n19319), .Z(n25083) );
  XNOR U25616 ( .A(n25084), .B(n22178), .Z(n19319) );
  XOR U25617 ( .A(round_reg[772]), .B(n25085), .Z(n22178) );
  ANDN U25618 ( .B(n22177), .A(n23693), .Z(n25084) );
  XOR U25619 ( .A(n25086), .B(n22195), .Z(n22172) );
  XOR U25620 ( .A(round_reg[869]), .B(n24233), .Z(n22195) );
  IV U25621 ( .A(n22769), .Z(n24233) );
  XOR U25622 ( .A(n24782), .B(n25087), .Z(n22769) );
  XOR U25623 ( .A(n25088), .B(n25089), .Z(n24782) );
  XNOR U25624 ( .A(round_reg[1573]), .B(round_reg[1253]), .Z(n25089) );
  XOR U25625 ( .A(round_reg[293]), .B(n25090), .Z(n25088) );
  XOR U25626 ( .A(round_reg[933]), .B(round_reg[613]), .Z(n25090) );
  NOR U25627 ( .A(n22194), .B(n23680), .Z(n25086) );
  XOR U25628 ( .A(round_reg[119]), .B(n24223), .Z(n23680) );
  IV U25629 ( .A(n24205), .Z(n24223) );
  XNOR U25630 ( .A(n25091), .B(n25092), .Z(n24205) );
  XOR U25631 ( .A(round_reg[480]), .B(n24996), .Z(n22194) );
  XOR U25632 ( .A(n25095), .B(n22187), .Z(n18975) );
  XNOR U25633 ( .A(round_reg[940]), .B(n23300), .Z(n22187) );
  ANDN U25634 ( .B(n22186), .A(n23690), .Z(n25095) );
  XOR U25635 ( .A(round_reg[178]), .B(n24692), .Z(n23690) );
  IV U25636 ( .A(n24074), .Z(n22186) );
  XOR U25637 ( .A(round_reg[514]), .B(n24261), .Z(n24074) );
  IV U25638 ( .A(n25074), .Z(n24261) );
  XOR U25639 ( .A(n25096), .B(n22177), .Z(n24068) );
  XNOR U25640 ( .A(round_reg[410]), .B(n24227), .Z(n22177) );
  AND U25641 ( .A(n23694), .B(n23693), .Z(n25096) );
  XOR U25642 ( .A(round_reg[33]), .B(n23144), .Z(n23693) );
  XNOR U25643 ( .A(round_reg[1583]), .B(n21763), .Z(n23694) );
  XNOR U25644 ( .A(n25097), .B(n25098), .Z(n15000) );
  XNOR U25645 ( .A(n13357), .B(n13810), .Z(n25098) );
  XOR U25646 ( .A(n25099), .B(n14678), .Z(n13810) );
  XNOR U25647 ( .A(n24581), .B(n16011), .Z(n14678) );
  XNOR U25648 ( .A(n21794), .B(n18867), .Z(n16011) );
  XNOR U25649 ( .A(n25100), .B(n25101), .Z(n18867) );
  XOR U25650 ( .A(n20908), .B(n20035), .Z(n25101) );
  XOR U25651 ( .A(n25102), .B(n20927), .Z(n20035) );
  XNOR U25652 ( .A(round_reg[6]), .B(n23738), .Z(n20927) );
  XNOR U25653 ( .A(n25103), .B(n24395), .Z(n23738) );
  XOR U25654 ( .A(n25104), .B(n25105), .Z(n24395) );
  XNOR U25655 ( .A(round_reg[1541]), .B(round_reg[1221]), .Z(n25105) );
  XOR U25656 ( .A(round_reg[261]), .B(n25106), .Z(n25104) );
  XOR U25657 ( .A(round_reg[901]), .B(round_reg[581]), .Z(n25106) );
  AND U25658 ( .A(n20292), .B(n20294), .Z(n25102) );
  XOR U25659 ( .A(round_reg[1192]), .B(n25107), .Z(n20294) );
  XOR U25660 ( .A(round_reg[1556]), .B(n24137), .Z(n20292) );
  XNOR U25661 ( .A(n25108), .B(n20917), .Z(n20908) );
  XNOR U25662 ( .A(round_reg[210]), .B(n22645), .Z(n20917) );
  XNOR U25663 ( .A(n25109), .B(n25110), .Z(n22645) );
  ANDN U25664 ( .B(n20301), .A(n20302), .Z(n25108) );
  XNOR U25665 ( .A(round_reg[1053]), .B(n24962), .Z(n20302) );
  XOR U25666 ( .A(round_reg[1430]), .B(n24378), .Z(n20301) );
  XNOR U25667 ( .A(n17343), .B(n25111), .Z(n25100) );
  XNOR U25668 ( .A(n16548), .B(n18265), .Z(n25111) );
  XNOR U25669 ( .A(n25112), .B(n20921), .Z(n18265) );
  XOR U25670 ( .A(round_reg[151]), .B(n23254), .Z(n20921) );
  ANDN U25671 ( .B(n20288), .A(n20289), .Z(n25112) );
  XNOR U25672 ( .A(round_reg[960]), .B(n24538), .Z(n20289) );
  XOR U25673 ( .A(round_reg[1400]), .B(n24695), .Z(n20288) );
  IV U25674 ( .A(n24642), .Z(n24695) );
  XNOR U25675 ( .A(n25113), .B(n25114), .Z(n24642) );
  XNOR U25676 ( .A(n25115), .B(n20914), .Z(n16548) );
  XNOR U25677 ( .A(round_reg[92]), .B(n22119), .Z(n20914) );
  AND U25678 ( .A(n20297), .B(n20299), .Z(n25115) );
  XOR U25679 ( .A(round_reg[1264]), .B(n25116), .Z(n20299) );
  XOR U25680 ( .A(round_reg[1337]), .B(n23469), .Z(n20297) );
  XNOR U25681 ( .A(n25117), .B(n20924), .Z(n17343) );
  XNOR U25682 ( .A(round_reg[258]), .B(n23252), .Z(n20924) );
  XOR U25683 ( .A(round_reg[1102]), .B(n23134), .Z(n20306) );
  XOR U25684 ( .A(round_reg[1491]), .B(n24288), .Z(n20305) );
  IV U25685 ( .A(n25120), .Z(n24288) );
  XOR U25686 ( .A(n25121), .B(n25122), .Z(n21794) );
  XOR U25687 ( .A(n20280), .B(n17023), .Z(n25122) );
  XOR U25688 ( .A(n25123), .B(n21691), .Z(n17023) );
  XNOR U25689 ( .A(round_reg[686]), .B(n24828), .Z(n21691) );
  AND U25690 ( .A(n22960), .B(n22073), .Z(n25123) );
  XOR U25691 ( .A(round_reg[211]), .B(n25120), .Z(n22073) );
  XNOR U25692 ( .A(n25124), .B(n25125), .Z(n25120) );
  XOR U25693 ( .A(round_reg[620]), .B(n23300), .Z(n22960) );
  XNOR U25694 ( .A(n25128), .B(n21694), .Z(n20280) );
  XNOR U25695 ( .A(round_reg[764]), .B(n24026), .Z(n21694) );
  XNOR U25696 ( .A(n24345), .B(n25129), .Z(n24026) );
  XNOR U25697 ( .A(n25130), .B(n25131), .Z(n24345) );
  XNOR U25698 ( .A(round_reg[1468]), .B(round_reg[1148]), .Z(n25131) );
  XOR U25699 ( .A(round_reg[188]), .B(n25132), .Z(n25130) );
  XOR U25700 ( .A(round_reg[828]), .B(round_reg[508]), .Z(n25132) );
  ANDN U25701 ( .B(n22970), .A(n22067), .Z(n25128) );
  XOR U25702 ( .A(round_reg[259]), .B(n25133), .Z(n22067) );
  XNOR U25703 ( .A(round_reg[333]), .B(n21911), .Z(n22970) );
  IV U25704 ( .A(n24515), .Z(n21911) );
  XNOR U25705 ( .A(n16692), .B(n25134), .Z(n25121) );
  XNOR U25706 ( .A(n18090), .B(n17390), .Z(n25134) );
  XOR U25707 ( .A(n25135), .B(n22075), .Z(n17390) );
  XNOR U25708 ( .A(round_reg[843]), .B(n24767), .Z(n22075) );
  ANDN U25709 ( .B(n22069), .A(n22963), .Z(n25135) );
  XNOR U25710 ( .A(round_reg[454]), .B(n24251), .Z(n22963) );
  XOR U25711 ( .A(round_reg[93]), .B(n24962), .Z(n22069) );
  XNOR U25712 ( .A(n25136), .B(n25137), .Z(n24962) );
  XNOR U25713 ( .A(n25138), .B(n21680), .Z(n18090) );
  XNOR U25714 ( .A(round_reg[914]), .B(n24504), .Z(n21680) );
  AND U25715 ( .A(n22967), .B(n22064), .Z(n25138) );
  XOR U25716 ( .A(n25139), .B(n21685), .Z(n16692) );
  XOR U25717 ( .A(round_reg[810]), .B(n22274), .Z(n21685) );
  AND U25718 ( .A(n22973), .B(n24584), .Z(n25139) );
  XOR U25719 ( .A(round_reg[7]), .B(n24757), .Z(n24584) );
  XOR U25720 ( .A(round_reg[384]), .B(n24381), .Z(n22973) );
  XNOR U25721 ( .A(n25142), .B(n22967), .Z(n24581) );
  XOR U25722 ( .A(round_reg[552]), .B(n23397), .Z(n22967) );
  IV U25723 ( .A(n25107), .Z(n23397) );
  XOR U25724 ( .A(n25143), .B(n25144), .Z(n25107) );
  XOR U25725 ( .A(round_reg[152]), .B(n25011), .Z(n22064) );
  XNOR U25726 ( .A(round_reg[1401]), .B(n23623), .Z(n21679) );
  IV U25727 ( .A(n24422), .Z(n23623) );
  XNOR U25728 ( .A(n25145), .B(n25146), .Z(n24422) );
  XOR U25729 ( .A(n22343), .B(n19971), .Z(n14679) );
  XNOR U25730 ( .A(n25147), .B(n25148), .Z(n22585) );
  XOR U25731 ( .A(n19334), .B(n19606), .Z(n25148) );
  XOR U25732 ( .A(n25149), .B(n21892), .Z(n19606) );
  ANDN U25733 ( .B(n22588), .A(n22589), .Z(n25149) );
  XOR U25734 ( .A(round_reg[929]), .B(n23745), .Z(n22589) );
  XOR U25735 ( .A(round_reg[976]), .B(n23915), .Z(n22588) );
  XNOR U25736 ( .A(n25150), .B(n21883), .Z(n19334) );
  XOR U25737 ( .A(round_reg[1572]), .B(n25023), .Z(n21883) );
  AND U25738 ( .A(n20961), .B(n20963), .Z(n25150) );
  XOR U25739 ( .A(round_reg[825]), .B(n25151), .Z(n20963) );
  XOR U25740 ( .A(round_reg[1208]), .B(n23777), .Z(n20961) );
  XNOR U25741 ( .A(n16770), .B(n25152), .Z(n25147) );
  XOR U25742 ( .A(n18989), .B(n16452), .Z(n25152) );
  XNOR U25743 ( .A(n25153), .B(n23131), .Z(n16452) );
  IV U25744 ( .A(n24502), .Z(n23131) );
  XOR U25745 ( .A(round_reg[1289]), .B(n24421), .Z(n24502) );
  IV U25746 ( .A(n23668), .Z(n24421) );
  XOR U25747 ( .A(n24353), .B(n25154), .Z(n23668) );
  XOR U25748 ( .A(n25155), .B(n25156), .Z(n24353) );
  XNOR U25749 ( .A(round_reg[1353]), .B(round_reg[1033]), .Z(n25156) );
  XOR U25750 ( .A(round_reg[393]), .B(n25157), .Z(n25155) );
  XOR U25751 ( .A(round_reg[73]), .B(round_reg[713]), .Z(n25157) );
  AND U25752 ( .A(n22378), .B(n22377), .Z(n25153) );
  XOR U25753 ( .A(round_reg[1216]), .B(n23151), .Z(n22377) );
  IV U25754 ( .A(n24443), .Z(n23151) );
  XNOR U25755 ( .A(round_reg[858]), .B(n23471), .Z(n22378) );
  XOR U25756 ( .A(n25158), .B(n21895), .Z(n18989) );
  XNOR U25757 ( .A(round_reg[1446]), .B(n23988), .Z(n21895) );
  XNOR U25758 ( .A(round_reg[701]), .B(n24121), .Z(n20952) );
  XOR U25759 ( .A(round_reg[1069]), .B(n24183), .Z(n20950) );
  XOR U25760 ( .A(n25159), .B(n21886), .Z(n16770) );
  XOR U25761 ( .A(round_reg[1507]), .B(n23280), .Z(n21886) );
  AND U25762 ( .A(n20956), .B(n20954), .Z(n25159) );
  XOR U25763 ( .A(round_reg[1118]), .B(n21923), .Z(n20954) );
  XNOR U25764 ( .A(round_reg[715]), .B(n23270), .Z(n20956) );
  XOR U25765 ( .A(n25162), .B(n25163), .Z(n22382) );
  XOR U25766 ( .A(n22099), .B(n20269), .Z(n25163) );
  XNOR U25767 ( .A(n25164), .B(n20867), .Z(n20269) );
  IV U25768 ( .A(n24494), .Z(n20867) );
  XOR U25769 ( .A(round_reg[400]), .B(n22445), .Z(n24494) );
  XOR U25770 ( .A(n25165), .B(n25166), .Z(n22445) );
  ANDN U25771 ( .B(n22337), .A(n22338), .Z(n25164) );
  XNOR U25772 ( .A(round_reg[1573]), .B(n25167), .Z(n22338) );
  XOR U25773 ( .A(round_reg[23]), .B(n22635), .Z(n22337) );
  XNOR U25774 ( .A(n25168), .B(n20862), .Z(n22099) );
  XOR U25775 ( .A(round_reg[349]), .B(n23910), .Z(n20862) );
  AND U25776 ( .A(n22837), .B(n24491), .Z(n25168) );
  XOR U25777 ( .A(n19702), .B(n25169), .Z(n25162) );
  XOR U25778 ( .A(n22937), .B(n24481), .Z(n25169) );
  XNOR U25779 ( .A(n25170), .B(n20875), .Z(n24481) );
  XOR U25780 ( .A(round_reg[568]), .B(n23777), .Z(n20875) );
  ANDN U25781 ( .B(n22348), .A(n22349), .Z(n25170) );
  XNOR U25782 ( .A(round_reg[1353]), .B(n24448), .Z(n22349) );
  XOR U25783 ( .A(round_reg[168]), .B(n22821), .Z(n22348) );
  XNOR U25784 ( .A(n25171), .B(n20871), .Z(n22937) );
  XOR U25785 ( .A(round_reg[470]), .B(n24378), .Z(n20871) );
  ANDN U25786 ( .B(n22340), .A(n22341), .Z(n25171) );
  XNOR U25787 ( .A(round_reg[1290]), .B(n24399), .Z(n22341) );
  IV U25788 ( .A(n24116), .Z(n24399) );
  XOR U25789 ( .A(n25172), .B(n24942), .Z(n24116) );
  XNOR U25790 ( .A(n25173), .B(n25174), .Z(n24942) );
  XNOR U25791 ( .A(round_reg[1545]), .B(round_reg[1225]), .Z(n25174) );
  XOR U25792 ( .A(round_reg[265]), .B(n25175), .Z(n25173) );
  XOR U25793 ( .A(round_reg[905]), .B(round_reg[585]), .Z(n25175) );
  XOR U25794 ( .A(round_reg[109]), .B(n24183), .Z(n22340) );
  XNOR U25795 ( .A(n25176), .B(n20858), .Z(n19702) );
  XNOR U25796 ( .A(round_reg[636]), .B(n23816), .Z(n20858) );
  IV U25797 ( .A(n25177), .Z(n23816) );
  ANDN U25798 ( .B(n22345), .A(n22346), .Z(n25176) );
  XOR U25799 ( .A(round_reg[1447]), .B(n21189), .Z(n22346) );
  XOR U25800 ( .A(n25178), .B(n24783), .Z(n21189) );
  XNOR U25801 ( .A(n25179), .B(n25180), .Z(n24783) );
  XNOR U25802 ( .A(round_reg[1062]), .B(round_reg[102]), .Z(n25180) );
  XOR U25803 ( .A(round_reg[1382]), .B(n25181), .Z(n25179) );
  XOR U25804 ( .A(round_reg[742]), .B(round_reg[422]), .Z(n25181) );
  XOR U25805 ( .A(round_reg[227]), .B(n23280), .Z(n22345) );
  XOR U25806 ( .A(n25182), .B(n25183), .Z(n23280) );
  XNOR U25807 ( .A(n25184), .B(n24491), .Z(n22343) );
  XOR U25808 ( .A(round_reg[275]), .B(n24202), .Z(n24491) );
  ANDN U25809 ( .B(n20860), .A(n22837), .Z(n25184) );
  XNOR U25810 ( .A(round_reg[1508]), .B(n23293), .Z(n22837) );
  IV U25811 ( .A(n22822), .Z(n23293) );
  XNOR U25812 ( .A(round_reg[1119]), .B(n24165), .Z(n20860) );
  IV U25813 ( .A(n24460), .Z(n24165) );
  XNOR U25814 ( .A(n25187), .B(n25188), .Z(n24460) );
  XOR U25815 ( .A(n21902), .B(n16792), .Z(n16662) );
  XOR U25816 ( .A(n21495), .B(n23128), .Z(n16792) );
  XOR U25817 ( .A(n25189), .B(n25190), .Z(n23128) );
  XOR U25818 ( .A(n15515), .B(n16985), .Z(n25190) );
  XNOR U25819 ( .A(n25191), .B(n21801), .Z(n16985) );
  XNOR U25820 ( .A(round_reg[21]), .B(n24861), .Z(n21801) );
  IV U25821 ( .A(n23393), .Z(n24861) );
  XOR U25822 ( .A(n25192), .B(n25193), .Z(n23393) );
  ANDN U25823 ( .B(n21802), .A(n21559), .Z(n25191) );
  XOR U25824 ( .A(round_reg[1207]), .B(n23127), .Z(n21559) );
  XOR U25825 ( .A(round_reg[1571]), .B(n23256), .Z(n21802) );
  XOR U25826 ( .A(n25194), .B(n25195), .Z(n23256) );
  XNOR U25827 ( .A(n25196), .B(n20970), .Z(n15515) );
  XNOR U25828 ( .A(round_reg[107]), .B(n23946), .Z(n20970) );
  ANDN U25829 ( .B(n20969), .A(n21553), .Z(n25196) );
  XOR U25830 ( .A(n20513), .B(n25197), .Z(n25189) );
  XOR U25831 ( .A(n18314), .B(n19442), .Z(n25197) );
  XNOR U25832 ( .A(n25198), .B(n20975), .Z(n19442) );
  XNOR U25833 ( .A(round_reg[273]), .B(n23778), .Z(n20975) );
  IV U25834 ( .A(n22362), .Z(n23778) );
  XNOR U25835 ( .A(n25199), .B(n25200), .Z(n22362) );
  AND U25836 ( .A(n21549), .B(n20976), .Z(n25198) );
  XOR U25837 ( .A(round_reg[1506]), .B(n23480), .Z(n20976) );
  XOR U25838 ( .A(n24849), .B(n25201), .Z(n23480) );
  XOR U25839 ( .A(n25202), .B(n25203), .Z(n24849) );
  XNOR U25840 ( .A(round_reg[1441]), .B(round_reg[1121]), .Z(n25203) );
  XOR U25841 ( .A(round_reg[161]), .B(n25204), .Z(n25202) );
  XOR U25842 ( .A(round_reg[801]), .B(round_reg[481]), .Z(n25204) );
  XNOR U25843 ( .A(round_reg[1117]), .B(n23902), .Z(n21549) );
  XOR U25844 ( .A(n25205), .B(n24263), .Z(n18314) );
  XOR U25845 ( .A(round_reg[225]), .B(n23019), .Z(n24263) );
  AND U25846 ( .A(n21545), .B(n21904), .Z(n25205) );
  XOR U25847 ( .A(round_reg[1445]), .B(n23919), .Z(n21904) );
  XOR U25848 ( .A(n25208), .B(n25209), .Z(n23919) );
  XNOR U25849 ( .A(round_reg[1068]), .B(n24364), .Z(n21545) );
  XOR U25850 ( .A(n25210), .B(n24273), .Z(n20513) );
  IV U25851 ( .A(n20980), .Z(n24273) );
  XNOR U25852 ( .A(round_reg[166]), .B(n23988), .Z(n20980) );
  XOR U25853 ( .A(n24955), .B(n25211), .Z(n23988) );
  XNOR U25854 ( .A(n25212), .B(n25213), .Z(n24955) );
  XNOR U25855 ( .A(round_reg[1510]), .B(round_reg[1190]), .Z(n25213) );
  XOR U25856 ( .A(round_reg[230]), .B(n25214), .Z(n25212) );
  XOR U25857 ( .A(round_reg[870]), .B(round_reg[550]), .Z(n25214) );
  NOR U25858 ( .A(n20979), .B(n21556), .Z(n25210) );
  XOR U25859 ( .A(round_reg[975]), .B(n23606), .Z(n21556) );
  XOR U25860 ( .A(n25215), .B(n24672), .Z(n23606) );
  XNOR U25861 ( .A(n25216), .B(n25217), .Z(n24672) );
  XNOR U25862 ( .A(round_reg[1550]), .B(round_reg[1230]), .Z(n25217) );
  XOR U25863 ( .A(round_reg[270]), .B(n25218), .Z(n25216) );
  XOR U25864 ( .A(round_reg[910]), .B(round_reg[590]), .Z(n25218) );
  XNOR U25865 ( .A(round_reg[1351]), .B(n21316), .Z(n20979) );
  XOR U25866 ( .A(n25219), .B(n25220), .Z(n21495) );
  XNOR U25867 ( .A(n19285), .B(n19342), .Z(n25220) );
  XOR U25868 ( .A(round_reg[1067]), .B(n23946), .Z(n20520) );
  XOR U25869 ( .A(n25222), .B(n25064), .Z(n23946) );
  XNOR U25870 ( .A(n25223), .B(n25224), .Z(n25064) );
  XNOR U25871 ( .A(round_reg[1451]), .B(round_reg[1131]), .Z(n25224) );
  XOR U25872 ( .A(round_reg[171]), .B(n25225), .Z(n25223) );
  XOR U25873 ( .A(round_reg[811]), .B(round_reg[491]), .Z(n25225) );
  ANDN U25874 ( .B(n19358), .A(n19356), .Z(n25221) );
  XNOR U25875 ( .A(round_reg[699]), .B(n22986), .Z(n19356) );
  XNOR U25876 ( .A(round_reg[633]), .B(n24875), .Z(n19358) );
  IV U25877 ( .A(n23854), .Z(n24875) );
  XOR U25878 ( .A(n25226), .B(n25227), .Z(n23854) );
  XNOR U25879 ( .A(n25228), .B(n20526), .Z(n19285) );
  XOR U25880 ( .A(round_reg[1116]), .B(n23568), .Z(n20526) );
  XOR U25881 ( .A(n25229), .B(n25230), .Z(n23568) );
  AND U25882 ( .A(n19362), .B(n20527), .Z(n25228) );
  XNOR U25883 ( .A(round_reg[713]), .B(n24448), .Z(n20527) );
  XNOR U25884 ( .A(round_reg[346]), .B(n24823), .Z(n19362) );
  XOR U25885 ( .A(n16046), .B(n25231), .Z(n25219) );
  XNOR U25886 ( .A(n17718), .B(n17408), .Z(n25231) );
  XOR U25887 ( .A(n25232), .B(n20907), .Z(n17408) );
  XOR U25888 ( .A(round_reg[1206]), .B(n25233), .Z(n20907) );
  NOR U25889 ( .A(n20906), .B(n21515), .Z(n25232) );
  XOR U25890 ( .A(round_reg[397]), .B(n23245), .Z(n21515) );
  XNOR U25891 ( .A(round_reg[823]), .B(n24029), .Z(n20906) );
  XNOR U25892 ( .A(n25234), .B(n24754), .Z(n17718) );
  XOR U25893 ( .A(round_reg[1278]), .B(n23877), .Z(n24754) );
  ANDN U25894 ( .B(n19366), .A(n19367), .Z(n25234) );
  XOR U25895 ( .A(round_reg[467]), .B(n22508), .Z(n19367) );
  XOR U25896 ( .A(n25235), .B(n25236), .Z(n22508) );
  XNOR U25897 ( .A(round_reg[856]), .B(n23447), .Z(n19366) );
  XNOR U25898 ( .A(n25237), .B(n23579), .Z(n16046) );
  XOR U25899 ( .A(round_reg[974]), .B(n22115), .Z(n23579) );
  XOR U25900 ( .A(n24958), .B(n25238), .Z(n22115) );
  XOR U25901 ( .A(n25239), .B(n25240), .Z(n24958) );
  XNOR U25902 ( .A(round_reg[1549]), .B(round_reg[1229]), .Z(n25240) );
  XOR U25903 ( .A(round_reg[269]), .B(n25241), .Z(n25239) );
  XOR U25904 ( .A(round_reg[909]), .B(round_reg[589]), .Z(n25241) );
  NOR U25905 ( .A(n19370), .B(n19372), .Z(n25237) );
  XOR U25906 ( .A(round_reg[565]), .B(n25242), .Z(n19372) );
  XNOR U25907 ( .A(round_reg[927]), .B(n24409), .Z(n19370) );
  XNOR U25908 ( .A(n25243), .B(n20969), .Z(n21902) );
  XOR U25909 ( .A(round_reg[1288]), .B(n25078), .Z(n20969) );
  XOR U25910 ( .A(n25244), .B(n25245), .Z(n25078) );
  AND U25911 ( .A(n21554), .B(n21553), .Z(n25243) );
  XOR U25912 ( .A(round_reg[1279]), .B(n21603), .Z(n21553) );
  XNOR U25913 ( .A(round_reg[857]), .B(n24098), .Z(n21554) );
  XNOR U25914 ( .A(n25246), .B(n14682), .Z(n13357) );
  XNOR U25915 ( .A(n24086), .B(n17667), .Z(n14682) );
  IV U25916 ( .A(n13892), .Z(n17667) );
  XNOR U25917 ( .A(n21790), .B(n21321), .Z(n13892) );
  XNOR U25918 ( .A(n25247), .B(n25248), .Z(n21321) );
  XOR U25919 ( .A(n21138), .B(n18638), .Z(n25248) );
  XOR U25920 ( .A(n25249), .B(n21144), .Z(n18638) );
  XNOR U25921 ( .A(round_reg[1010]), .B(n23781), .Z(n21144) );
  IV U25922 ( .A(n24052), .Z(n23781) );
  XNOR U25923 ( .A(n25250), .B(n25251), .Z(n24052) );
  ANDN U25924 ( .B(n21143), .A(n20804), .Z(n25249) );
  XNOR U25925 ( .A(n25252), .B(n23536), .Z(n21138) );
  XNOR U25926 ( .A(round_reg[1178]), .B(n23471), .Z(n23536) );
  XNOR U25927 ( .A(n25254), .B(n25255), .Z(n24817) );
  XNOR U25928 ( .A(round_reg[1433]), .B(round_reg[1113]), .Z(n25255) );
  XOR U25929 ( .A(round_reg[153]), .B(n25256), .Z(n25254) );
  XOR U25930 ( .A(round_reg[793]), .B(round_reg[473]), .Z(n25256) );
  ANDN U25931 ( .B(n23539), .A(n20878), .Z(n25252) );
  XOR U25932 ( .A(round_reg[433]), .B(n24943), .Z(n20878) );
  XOR U25933 ( .A(round_reg[795]), .B(n23411), .Z(n23539) );
  XOR U25934 ( .A(n18673), .B(n25257), .Z(n25247) );
  XNOR U25935 ( .A(n19216), .B(n19611), .Z(n25257) );
  XOR U25936 ( .A(n25258), .B(n21152), .Z(n19611) );
  XOR U25937 ( .A(round_reg[1039]), .B(n21605), .Z(n21152) );
  XOR U25938 ( .A(n25259), .B(n25260), .Z(n21605) );
  XOR U25939 ( .A(round_reg[605]), .B(n24171), .Z(n22170) );
  XOR U25940 ( .A(round_reg[671]), .B(n23325), .Z(n21153) );
  XNOR U25941 ( .A(n25261), .B(n21156), .Z(n19216) );
  XOR U25942 ( .A(round_reg[1088]), .B(n23011), .Z(n21156) );
  XNOR U25943 ( .A(n25262), .B(n25263), .Z(n25027) );
  XNOR U25944 ( .A(round_reg[127]), .B(round_reg[1087]), .Z(n25263) );
  XOR U25945 ( .A(round_reg[1407]), .B(n25264), .Z(n25262) );
  XOR U25946 ( .A(round_reg[767]), .B(round_reg[447]), .Z(n25264) );
  XOR U25947 ( .A(n25265), .B(n25266), .Z(n24725) );
  XNOR U25948 ( .A(round_reg[1472]), .B(round_reg[1152]), .Z(n25266) );
  XOR U25949 ( .A(round_reg[192]), .B(n25267), .Z(n25265) );
  XOR U25950 ( .A(round_reg[832]), .B(round_reg[512]), .Z(n25267) );
  ANDN U25951 ( .B(n21157), .A(n21655), .Z(n25261) );
  XNOR U25952 ( .A(round_reg[382]), .B(n24315), .Z(n21655) );
  XOR U25953 ( .A(n25268), .B(n24344), .Z(n24315) );
  XOR U25954 ( .A(n25269), .B(n25270), .Z(n24344) );
  XNOR U25955 ( .A(round_reg[1597]), .B(round_reg[1277]), .Z(n25270) );
  XOR U25956 ( .A(round_reg[317]), .B(n25271), .Z(n25269) );
  XOR U25957 ( .A(round_reg[957]), .B(round_reg[637]), .Z(n25271) );
  XOR U25958 ( .A(round_reg[749]), .B(n24183), .Z(n21157) );
  XNOR U25959 ( .A(n25272), .B(n21148), .Z(n18673) );
  XOR U25960 ( .A(round_reg[1250]), .B(n24019), .Z(n21148) );
  XOR U25961 ( .A(n25273), .B(n25274), .Z(n24019) );
  ANDN U25962 ( .B(n21149), .A(n24077), .Z(n25272) );
  XOR U25963 ( .A(round_reg[503]), .B(n24029), .Z(n24077) );
  XOR U25964 ( .A(round_reg[892]), .B(n23147), .Z(n21149) );
  XOR U25965 ( .A(n25275), .B(n25276), .Z(n21790) );
  XOR U25966 ( .A(n19740), .B(n15248), .Z(n25276) );
  XOR U25967 ( .A(n25277), .B(n21175), .Z(n15248) );
  IV U25968 ( .A(n23523), .Z(n21175) );
  XOR U25969 ( .A(round_reg[502]), .B(n25278), .Z(n23523) );
  AND U25970 ( .A(n23935), .B(n21176), .Z(n25277) );
  XOR U25971 ( .A(round_reg[77]), .B(n23245), .Z(n21176) );
  XOR U25972 ( .A(n24671), .B(n25279), .Z(n23245) );
  XOR U25973 ( .A(n25280), .B(n25281), .Z(n24671) );
  XNOR U25974 ( .A(round_reg[141]), .B(round_reg[1101]), .Z(n25281) );
  XOR U25975 ( .A(round_reg[1421]), .B(n25282), .Z(n25280) );
  XOR U25976 ( .A(round_reg[781]), .B(round_reg[461]), .Z(n25282) );
  XNOR U25977 ( .A(round_reg[1322]), .B(n22649), .Z(n23935) );
  XOR U25978 ( .A(n25283), .B(n21167), .Z(n19740) );
  XOR U25979 ( .A(round_reg[381]), .B(n24121), .Z(n21167) );
  XOR U25980 ( .A(n25284), .B(n25285), .Z(n24121) );
  ANDN U25981 ( .B(n21166), .A(n23939), .Z(n25283) );
  XOR U25982 ( .A(round_reg[1476]), .B(n24089), .Z(n23939) );
  IV U25983 ( .A(n24405), .Z(n24089) );
  XOR U25984 ( .A(n25286), .B(n25287), .Z(n24405) );
  XOR U25985 ( .A(round_reg[307]), .B(n21312), .Z(n21166) );
  XOR U25986 ( .A(n24918), .B(n25288), .Z(n21312) );
  XNOR U25987 ( .A(n25289), .B(n25290), .Z(n24918) );
  XNOR U25988 ( .A(round_reg[1331]), .B(round_reg[1011]), .Z(n25290) );
  XOR U25989 ( .A(round_reg[371]), .B(n25291), .Z(n25289) );
  XOR U25990 ( .A(round_reg[691]), .B(round_reg[51]), .Z(n25291) );
  XNOR U25991 ( .A(n18210), .B(n25292), .Z(n25275) );
  XOR U25992 ( .A(n15835), .B(n20842), .Z(n25292) );
  XNOR U25993 ( .A(n25293), .B(n21163), .Z(n20842) );
  XOR U25994 ( .A(round_reg[432]), .B(n25294), .Z(n21163) );
  AND U25995 ( .A(n23932), .B(n21162), .Z(n25293) );
  XOR U25996 ( .A(round_reg[55]), .B(n24715), .Z(n21162) );
  XNOR U25997 ( .A(round_reg[1541]), .B(n23400), .Z(n23932) );
  IV U25998 ( .A(n22206), .Z(n23400) );
  XNOR U25999 ( .A(n25295), .B(n21172), .Z(n15835) );
  XOR U26000 ( .A(round_reg[604]), .B(n24372), .Z(n21172) );
  AND U26001 ( .A(n23937), .B(n21171), .Z(n25295) );
  XOR U26002 ( .A(round_reg[195]), .B(n24697), .Z(n21171) );
  XNOR U26003 ( .A(round_reg[1415]), .B(n21766), .Z(n23937) );
  XNOR U26004 ( .A(n25296), .B(n21180), .Z(n18210) );
  XOR U26005 ( .A(round_reg[536]), .B(n23447), .Z(n21180) );
  IV U26006 ( .A(n24313), .Z(n23447) );
  XNOR U26007 ( .A(n25297), .B(n25041), .Z(n24313) );
  XNOR U26008 ( .A(n25298), .B(n25299), .Z(n25041) );
  XNOR U26009 ( .A(round_reg[1431]), .B(round_reg[1111]), .Z(n25299) );
  XOR U26010 ( .A(round_reg[151]), .B(n25300), .Z(n25298) );
  XOR U26011 ( .A(round_reg[791]), .B(round_reg[471]), .Z(n25300) );
  XOR U26012 ( .A(round_reg[1385]), .B(n23876), .Z(n23929) );
  XOR U26013 ( .A(round_reg[136]), .B(n24134), .Z(n21179) );
  XNOR U26014 ( .A(n25301), .B(n21143), .Z(n24086) );
  XOR U26015 ( .A(round_reg[899]), .B(n25133), .Z(n21143) );
  AND U26016 ( .A(n20806), .B(n20804), .Z(n25301) );
  XOR U26017 ( .A(round_reg[537]), .B(n24098), .Z(n20804) );
  IV U26018 ( .A(n21914), .Z(n24098) );
  XNOR U26019 ( .A(n24509), .B(n25302), .Z(n21914) );
  XOR U26020 ( .A(n25303), .B(n25304), .Z(n24509) );
  XNOR U26021 ( .A(round_reg[1432]), .B(round_reg[1112]), .Z(n25304) );
  XOR U26022 ( .A(round_reg[152]), .B(n25305), .Z(n25303) );
  XOR U26023 ( .A(round_reg[792]), .B(round_reg[472]), .Z(n25305) );
  XNOR U26024 ( .A(round_reg[137]), .B(n23283), .Z(n20806) );
  XOR U26025 ( .A(n25245), .B(n25306), .Z(n23283) );
  XNOR U26026 ( .A(n25307), .B(n25308), .Z(n25245) );
  XNOR U26027 ( .A(round_reg[1352]), .B(round_reg[1032]), .Z(n25308) );
  XOR U26028 ( .A(round_reg[392]), .B(n25309), .Z(n25307) );
  XOR U26029 ( .A(round_reg[72]), .B(round_reg[712]), .Z(n25309) );
  NOR U26030 ( .A(n13298), .B(n13300), .Z(n25246) );
  XNOR U26031 ( .A(n15911), .B(n21397), .Z(n13300) );
  XNOR U26032 ( .A(n25310), .B(n23950), .Z(n21397) );
  ANDN U26033 ( .B(n23450), .A(n20262), .Z(n25310) );
  XOR U26034 ( .A(round_reg[1248]), .B(n24272), .Z(n20262) );
  IV U26035 ( .A(n17494), .Z(n15911) );
  XOR U26036 ( .A(n20134), .B(n20191), .Z(n17494) );
  XOR U26037 ( .A(n25311), .B(n25312), .Z(n20191) );
  XNOR U26038 ( .A(n18831), .B(n17584), .Z(n25312) );
  XNOR U26039 ( .A(n25313), .B(n21586), .Z(n17584) );
  XOR U26040 ( .A(round_reg[1383]), .B(n24450), .Z(n21586) );
  ANDN U26041 ( .B(n21368), .A(n21369), .Z(n25313) );
  XNOR U26042 ( .A(round_reg[896]), .B(n24443), .Z(n21369) );
  XNOR U26043 ( .A(n25314), .B(n25315), .Z(n24967) );
  XNOR U26044 ( .A(round_reg[1280]), .B(round_reg[0]), .Z(n25315) );
  XOR U26045 ( .A(round_reg[320]), .B(n25316), .Z(n25314) );
  XOR U26046 ( .A(round_reg[960]), .B(round_reg[640]), .Z(n25316) );
  XOR U26047 ( .A(round_reg[1007]), .B(n24564), .Z(n21368) );
  XOR U26048 ( .A(n21594), .B(n25318), .Z(n18831) );
  XOR U26049 ( .A(n25319), .B(n25320), .Z(n25318) );
  NAND U26050 ( .A(n11363), .B(n25321), .Z(n25320) );
  AND U26051 ( .A(n6455), .B(n15691), .Z(n25321) );
  IV U26052 ( .A(rc_i[2]), .Z(n6455) );
  IV U26053 ( .A(rc_i[1]), .Z(n11363) );
  ANDN U26054 ( .B(n21381), .A(n21382), .Z(n25319) );
  XNOR U26055 ( .A(round_reg[792]), .B(n25011), .Z(n21382) );
  XOR U26056 ( .A(round_reg[1175]), .B(n24139), .Z(n21381) );
  XNOR U26057 ( .A(round_reg[1539]), .B(n23896), .Z(n21594) );
  IV U26058 ( .A(n25133), .Z(n23896) );
  XOR U26059 ( .A(n21128), .B(n25322), .Z(n25311) );
  XOR U26060 ( .A(n17926), .B(n19116), .Z(n25322) );
  XNOR U26061 ( .A(n25323), .B(n24894), .Z(n19116) );
  XOR U26062 ( .A(round_reg[1320]), .B(n24687), .Z(n24894) );
  ANDN U26063 ( .B(n21385), .A(n21386), .Z(n25323) );
  XOR U26064 ( .A(round_reg[889]), .B(n22831), .Z(n21386) );
  XOR U26065 ( .A(n25324), .B(n25325), .Z(n25113) );
  XNOR U26066 ( .A(round_reg[1464]), .B(round_reg[1144]), .Z(n25325) );
  XOR U26067 ( .A(round_reg[184]), .B(n25326), .Z(n25324) );
  XOR U26068 ( .A(round_reg[824]), .B(round_reg[504]), .Z(n25326) );
  XOR U26069 ( .A(round_reg[1247]), .B(n24409), .Z(n21385) );
  IV U26070 ( .A(n25328), .Z(n24409) );
  XNOR U26071 ( .A(n25329), .B(n22387), .Z(n17926) );
  XOR U26072 ( .A(round_reg[1413]), .B(n22365), .Z(n22387) );
  XOR U26073 ( .A(n25079), .B(n25330), .Z(n22365) );
  XOR U26074 ( .A(n25331), .B(n25332), .Z(n25079) );
  XNOR U26075 ( .A(round_reg[1477]), .B(round_reg[1157]), .Z(n25332) );
  XOR U26076 ( .A(round_reg[197]), .B(n25333), .Z(n25331) );
  XOR U26077 ( .A(round_reg[837]), .B(round_reg[517]), .Z(n25333) );
  ANDN U26078 ( .B(n21372), .A(n21373), .Z(n25329) );
  XNOR U26079 ( .A(round_reg[668]), .B(n24415), .Z(n21373) );
  IV U26080 ( .A(n23121), .Z(n24415) );
  XOR U26081 ( .A(round_reg[1036]), .B(n24490), .Z(n21372) );
  XNOR U26082 ( .A(n25334), .B(n21591), .Z(n21128) );
  XOR U26083 ( .A(round_reg[1474]), .B(n25074), .Z(n21591) );
  ANDN U26084 ( .B(n21377), .A(n21378), .Z(n25334) );
  XOR U26085 ( .A(round_reg[746]), .B(n23528), .Z(n21378) );
  XOR U26086 ( .A(round_reg[1149]), .B(n21609), .Z(n21377) );
  XOR U26087 ( .A(n25337), .B(n25338), .Z(n20134) );
  XNOR U26088 ( .A(n17256), .B(n17130), .Z(n25338) );
  XOR U26089 ( .A(n25339), .B(n20263), .Z(n17130) );
  XNOR U26090 ( .A(round_reg[501]), .B(n25340), .Z(n20263) );
  ANDN U26091 ( .B(n23950), .A(n23450), .Z(n25339) );
  XOR U26092 ( .A(round_reg[1321]), .B(n24221), .Z(n23450) );
  XOR U26093 ( .A(round_reg[76]), .B(n24490), .Z(n23950) );
  XOR U26094 ( .A(n25341), .B(n23456), .Z(n17256) );
  XNOR U26095 ( .A(round_reg[603]), .B(n24156), .Z(n23456) );
  ANDN U26096 ( .B(n21391), .A(n21392), .Z(n25341) );
  XOR U26097 ( .A(round_reg[1414]), .B(n24251), .Z(n21392) );
  IV U26098 ( .A(n24397), .Z(n24251) );
  XNOR U26099 ( .A(n24928), .B(n25342), .Z(n24397) );
  XOR U26100 ( .A(n25343), .B(n25344), .Z(n24928) );
  XNOR U26101 ( .A(round_reg[1478]), .B(round_reg[1158]), .Z(n25344) );
  XOR U26102 ( .A(round_reg[198]), .B(n25345), .Z(n25343) );
  XOR U26103 ( .A(round_reg[838]), .B(round_reg[518]), .Z(n25345) );
  XOR U26104 ( .A(round_reg[194]), .B(n25074), .Z(n21391) );
  XOR U26105 ( .A(n25013), .B(n24966), .Z(n25074) );
  XOR U26106 ( .A(n25346), .B(n25347), .Z(n24966) );
  XNOR U26107 ( .A(round_reg[129]), .B(round_reg[1089]), .Z(n25347) );
  XOR U26108 ( .A(round_reg[1409]), .B(n25348), .Z(n25346) );
  XOR U26109 ( .A(round_reg[769]), .B(round_reg[449]), .Z(n25348) );
  XNOR U26110 ( .A(n25349), .B(n25350), .Z(n25013) );
  XNOR U26111 ( .A(round_reg[1538]), .B(round_reg[1218]), .Z(n25350) );
  XOR U26112 ( .A(round_reg[258]), .B(n25351), .Z(n25349) );
  XOR U26113 ( .A(round_reg[898]), .B(round_reg[578]), .Z(n25351) );
  XNOR U26114 ( .A(n21579), .B(n25352), .Z(n25337) );
  XNOR U26115 ( .A(n19907), .B(n17986), .Z(n25352) );
  XNOR U26116 ( .A(n25353), .B(n20268), .Z(n17986) );
  XNOR U26117 ( .A(round_reg[380]), .B(n23290), .Z(n20268) );
  XOR U26118 ( .A(n25354), .B(n25336), .Z(n23290) );
  XOR U26119 ( .A(n25355), .B(n25356), .Z(n25336) );
  XNOR U26120 ( .A(round_reg[124]), .B(round_reg[1084]), .Z(n25356) );
  XOR U26121 ( .A(round_reg[1404]), .B(n25357), .Z(n25355) );
  XOR U26122 ( .A(round_reg[764]), .B(round_reg[444]), .Z(n25357) );
  XOR U26123 ( .A(round_reg[1475]), .B(n24697), .Z(n21401) );
  XOR U26124 ( .A(n25000), .B(n25358), .Z(n24697) );
  XOR U26125 ( .A(n25359), .B(n25360), .Z(n25000) );
  XNOR U26126 ( .A(round_reg[130]), .B(round_reg[1090]), .Z(n25360) );
  XOR U26127 ( .A(round_reg[1410]), .B(n25361), .Z(n25359) );
  XOR U26128 ( .A(round_reg[770]), .B(round_reg[450]), .Z(n25361) );
  XOR U26129 ( .A(round_reg[306]), .B(n25362), .Z(n21400) );
  XOR U26130 ( .A(n25363), .B(n20253), .Z(n19907) );
  ANDN U26131 ( .B(n21395), .A(n21396), .Z(n25363) );
  XOR U26132 ( .A(round_reg[1384]), .B(n25364), .Z(n21396) );
  XOR U26133 ( .A(round_reg[135]), .B(n21766), .Z(n21395) );
  XNOR U26134 ( .A(n24548), .B(n25103), .Z(n21766) );
  XOR U26135 ( .A(n25365), .B(n25366), .Z(n25103) );
  XNOR U26136 ( .A(round_reg[1350]), .B(round_reg[1030]), .Z(n25366) );
  XOR U26137 ( .A(round_reg[390]), .B(n25367), .Z(n25365) );
  XOR U26138 ( .A(round_reg[710]), .B(round_reg[70]), .Z(n25367) );
  XOR U26139 ( .A(n25368), .B(n25369), .Z(n24548) );
  XNOR U26140 ( .A(round_reg[1479]), .B(round_reg[1159]), .Z(n25369) );
  XOR U26141 ( .A(round_reg[199]), .B(n25370), .Z(n25368) );
  XOR U26142 ( .A(round_reg[839]), .B(round_reg[519]), .Z(n25370) );
  XOR U26143 ( .A(n25371), .B(n20258), .Z(n21579) );
  XNOR U26144 ( .A(round_reg[431]), .B(n23241), .Z(n20258) );
  XOR U26145 ( .A(round_reg[1540]), .B(n22983), .Z(n21404) );
  XOR U26146 ( .A(round_reg[54]), .B(n24986), .Z(n21403) );
  XNOR U26147 ( .A(n25372), .B(n25373), .Z(n24986) );
  XNOR U26148 ( .A(n16323), .B(n23067), .Z(n13298) );
  XNOR U26149 ( .A(n25374), .B(n23355), .Z(n23067) );
  AND U26150 ( .A(n22713), .B(n24012), .Z(n25374) );
  IV U26151 ( .A(n22714), .Z(n24012) );
  XOR U26152 ( .A(round_reg[1522]), .B(n24859), .Z(n22714) );
  IV U26153 ( .A(n24023), .Z(n24859) );
  XOR U26154 ( .A(n22167), .B(n24030), .Z(n16323) );
  XNOR U26155 ( .A(n25375), .B(n25376), .Z(n24030) );
  XOR U26156 ( .A(n17114), .B(n23080), .Z(n25376) );
  XOR U26157 ( .A(n25377), .B(n21757), .Z(n23080) );
  XOR U26158 ( .A(round_reg[122]), .B(n22991), .Z(n21757) );
  XOR U26159 ( .A(n25226), .B(n25378), .Z(n22991) );
  XOR U26160 ( .A(n25379), .B(n25380), .Z(n25226) );
  XNOR U26161 ( .A(round_reg[1337]), .B(round_reg[1017]), .Z(n25380) );
  XOR U26162 ( .A(round_reg[377]), .B(n25381), .Z(n25379) );
  XOR U26163 ( .A(round_reg[697]), .B(round_reg[57]), .Z(n25381) );
  AND U26164 ( .A(n23424), .B(n21743), .Z(n25377) );
  XOR U26165 ( .A(round_reg[1230]), .B(n23497), .Z(n21743) );
  XOR U26166 ( .A(round_reg[1303]), .B(n22635), .Z(n23424) );
  XNOR U26167 ( .A(n25382), .B(n21761), .Z(n17114) );
  XOR U26168 ( .A(round_reg[288]), .B(n24272), .Z(n21761) );
  AND U26169 ( .A(n21723), .B(n20729), .Z(n25382) );
  XOR U26170 ( .A(round_reg[1132]), .B(n23392), .Z(n20729) );
  IV U26171 ( .A(n23598), .Z(n23392) );
  XOR U26172 ( .A(n25383), .B(n24566), .Z(n23598) );
  XOR U26173 ( .A(n25384), .B(n25385), .Z(n24566) );
  XNOR U26174 ( .A(round_reg[1516]), .B(round_reg[1196]), .Z(n25385) );
  XOR U26175 ( .A(round_reg[236]), .B(n25386), .Z(n25384) );
  XOR U26176 ( .A(round_reg[876]), .B(round_reg[556]), .Z(n25386) );
  XOR U26177 ( .A(round_reg[1521]), .B(n23801), .Z(n21723) );
  XOR U26178 ( .A(n23414), .B(n25387), .Z(n25375) );
  XOR U26179 ( .A(n17153), .B(n16008), .Z(n25387) );
  XNOR U26180 ( .A(n25388), .B(n21767), .Z(n16008) );
  XOR U26181 ( .A(round_reg[36]), .B(n23201), .Z(n21767) );
  AND U26182 ( .A(n21716), .B(n20719), .Z(n25388) );
  XOR U26183 ( .A(round_reg[1158]), .B(n25389), .Z(n20719) );
  XOR U26184 ( .A(round_reg[1586]), .B(n22105), .Z(n21716) );
  IV U26185 ( .A(n25362), .Z(n22105) );
  XOR U26186 ( .A(n25390), .B(n25391), .Z(n25362) );
  XNOR U26187 ( .A(n25392), .B(n21755), .Z(n17153) );
  XOR U26188 ( .A(round_reg[240]), .B(n23618), .Z(n21755) );
  XOR U26189 ( .A(n24761), .B(n25393), .Z(n23618) );
  XOR U26190 ( .A(n25394), .B(n25395), .Z(n24761) );
  XNOR U26191 ( .A(round_reg[1584]), .B(round_reg[1264]), .Z(n25395) );
  XOR U26192 ( .A(round_reg[304]), .B(n25396), .Z(n25394) );
  XOR U26193 ( .A(round_reg[944]), .B(round_reg[624]), .Z(n25396) );
  AND U26194 ( .A(n21720), .B(n20725), .Z(n25392) );
  IV U26195 ( .A(n21721), .Z(n20725) );
  XOR U26196 ( .A(round_reg[1083]), .B(n22369), .Z(n21721) );
  XOR U26197 ( .A(round_reg[1460]), .B(n22230), .Z(n21720) );
  XNOR U26198 ( .A(n25397), .B(n21764), .Z(n23414) );
  XOR U26199 ( .A(round_reg[181]), .B(n23803), .Z(n21764) );
  IV U26200 ( .A(n25340), .Z(n23803) );
  AND U26201 ( .A(n21713), .B(n20715), .Z(n25397) );
  IV U26202 ( .A(n21714), .Z(n20715) );
  XOR U26203 ( .A(round_reg[990]), .B(n23246), .Z(n21714) );
  XNOR U26204 ( .A(n25398), .B(n25188), .Z(n23246) );
  XNOR U26205 ( .A(n25399), .B(n25400), .Z(n25188) );
  XNOR U26206 ( .A(round_reg[1374]), .B(round_reg[1054]), .Z(n25400) );
  XOR U26207 ( .A(round_reg[414]), .B(n25401), .Z(n25399) );
  XOR U26208 ( .A(round_reg[94]), .B(round_reg[734]), .Z(n25401) );
  XOR U26209 ( .A(round_reg[1366]), .B(n23591), .Z(n21713) );
  IV U26210 ( .A(n25082), .Z(n23591) );
  XNOR U26211 ( .A(n24949), .B(n25402), .Z(n25082) );
  XOR U26212 ( .A(n25403), .B(n25404), .Z(n24949) );
  XNOR U26213 ( .A(round_reg[21]), .B(round_reg[1301]), .Z(n25404) );
  XOR U26214 ( .A(round_reg[341]), .B(n25405), .Z(n25403) );
  XOR U26215 ( .A(round_reg[981]), .B(round_reg[661]), .Z(n25405) );
  XOR U26216 ( .A(n25406), .B(n25407), .Z(n22167) );
  XOR U26217 ( .A(n19667), .B(n20192), .Z(n25407) );
  XOR U26218 ( .A(n25408), .B(n23362), .Z(n20192) );
  XOR U26219 ( .A(round_reg[652]), .B(n22368), .Z(n23362) );
  AND U26220 ( .A(n23077), .B(n22722), .Z(n25408) );
  XOR U26221 ( .A(round_reg[241]), .B(n23851), .Z(n22722) );
  XOR U26222 ( .A(round_reg[586]), .B(n24377), .Z(n23077) );
  IV U26223 ( .A(n24779), .Z(n24377) );
  XOR U26224 ( .A(n25410), .B(n25411), .Z(n25306) );
  XNOR U26225 ( .A(round_reg[1481]), .B(round_reg[1161]), .Z(n25411) );
  XOR U26226 ( .A(round_reg[201]), .B(n25412), .Z(n25410) );
  XOR U26227 ( .A(round_reg[841]), .B(round_reg[521]), .Z(n25412) );
  XNOR U26228 ( .A(n25413), .B(n23354), .Z(n19667) );
  XNOR U26229 ( .A(round_reg[730]), .B(n24227), .Z(n23354) );
  ANDN U26230 ( .B(n23355), .A(n22713), .Z(n25413) );
  XOR U26231 ( .A(round_reg[289]), .B(n23745), .Z(n22713) );
  XOR U26232 ( .A(n25414), .B(n25093), .Z(n23745) );
  XNOR U26233 ( .A(n25415), .B(n25416), .Z(n25093) );
  XNOR U26234 ( .A(round_reg[1504]), .B(round_reg[1184]), .Z(n25416) );
  XOR U26235 ( .A(round_reg[224]), .B(n25417), .Z(n25415) );
  XOR U26236 ( .A(round_reg[864]), .B(round_reg[544]), .Z(n25417) );
  XOR U26237 ( .A(round_reg[363]), .B(n24302), .Z(n23355) );
  XOR U26238 ( .A(n24571), .B(n25383), .Z(n24302) );
  XNOR U26239 ( .A(n25418), .B(n25419), .Z(n25383) );
  XNOR U26240 ( .A(round_reg[107]), .B(round_reg[1067]), .Z(n25419) );
  XOR U26241 ( .A(round_reg[1387]), .B(n25420), .Z(n25418) );
  XOR U26242 ( .A(round_reg[747]), .B(round_reg[427]), .Z(n25420) );
  XOR U26243 ( .A(n25421), .B(n25422), .Z(n24571) );
  XNOR U26244 ( .A(round_reg[1578]), .B(round_reg[1258]), .Z(n25422) );
  XOR U26245 ( .A(round_reg[298]), .B(n25423), .Z(n25421) );
  XOR U26246 ( .A(round_reg[938]), .B(round_reg[618]), .Z(n25423) );
  XOR U26247 ( .A(n19557), .B(n25424), .Z(n25406) );
  XOR U26248 ( .A(n19021), .B(n18333), .Z(n25424) );
  XNOR U26249 ( .A(n25425), .B(n23352), .Z(n18333) );
  XOR U26250 ( .A(round_reg[776]), .B(n24134), .Z(n23352) );
  IV U26251 ( .A(n23534), .Z(n24134) );
  XOR U26252 ( .A(n25426), .B(n25141), .Z(n23534) );
  XOR U26253 ( .A(n25427), .B(n25428), .Z(n25141) );
  XNOR U26254 ( .A(round_reg[1351]), .B(round_reg[1031]), .Z(n25428) );
  XOR U26255 ( .A(round_reg[391]), .B(n25429), .Z(n25427) );
  XOR U26256 ( .A(round_reg[71]), .B(round_reg[711]), .Z(n25429) );
  AND U26257 ( .A(n23074), .B(n22718), .Z(n25425) );
  IV U26258 ( .A(n23075), .Z(n22718) );
  XOR U26259 ( .A(round_reg[37]), .B(n24157), .Z(n23075) );
  XNOR U26260 ( .A(n25430), .B(n25431), .Z(n25211) );
  XNOR U26261 ( .A(round_reg[1061]), .B(round_reg[101]), .Z(n25431) );
  XOR U26262 ( .A(round_reg[1381]), .B(n25432), .Z(n25430) );
  XOR U26263 ( .A(round_reg[741]), .B(round_reg[421]), .Z(n25432) );
  XNOR U26264 ( .A(n25433), .B(n25434), .Z(n25185) );
  XNOR U26265 ( .A(round_reg[1572]), .B(round_reg[1252]), .Z(n25434) );
  XOR U26266 ( .A(round_reg[292]), .B(n25435), .Z(n25433) );
  XOR U26267 ( .A(round_reg[932]), .B(round_reg[612]), .Z(n25435) );
  XOR U26268 ( .A(round_reg[414]), .B(n23327), .Z(n23074) );
  XNOR U26269 ( .A(n25436), .B(n23358), .Z(n19021) );
  XOR U26270 ( .A(round_reg[873]), .B(n22972), .Z(n23358) );
  XNOR U26271 ( .A(n25437), .B(n25438), .Z(n22972) );
  AND U26272 ( .A(n22709), .B(n23069), .Z(n25436) );
  XOR U26273 ( .A(round_reg[484]), .B(n23482), .Z(n23069) );
  XOR U26274 ( .A(n25439), .B(n25440), .Z(n23482) );
  XNOR U26275 ( .A(round_reg[123]), .B(n22369), .Z(n22709) );
  XNOR U26276 ( .A(n25441), .B(n25442), .Z(n22369) );
  XNOR U26277 ( .A(n25443), .B(n23360), .Z(n19557) );
  XOR U26278 ( .A(round_reg[944]), .B(n24053), .Z(n23360) );
  IV U26279 ( .A(n25116), .Z(n24053) );
  XNOR U26280 ( .A(n24812), .B(n25444), .Z(n25116) );
  XOR U26281 ( .A(n25445), .B(n25446), .Z(n24812) );
  XNOR U26282 ( .A(round_reg[1519]), .B(round_reg[1199]), .Z(n25446) );
  XOR U26283 ( .A(round_reg[239]), .B(n25447), .Z(n25445) );
  XOR U26284 ( .A(round_reg[879]), .B(round_reg[559]), .Z(n25447) );
  AND U26285 ( .A(n23072), .B(n22726), .Z(n25443) );
  XOR U26286 ( .A(round_reg[182]), .B(n25278), .Z(n22726) );
  XOR U26287 ( .A(round_reg[518]), .B(n24218), .Z(n23072) );
  IV U26288 ( .A(n25389), .Z(n24218) );
  XNOR U26289 ( .A(n25448), .B(n25140), .Z(n25389) );
  XNOR U26290 ( .A(n25449), .B(n25450), .Z(n25140) );
  XNOR U26291 ( .A(round_reg[1542]), .B(round_reg[1222]), .Z(n25450) );
  XOR U26292 ( .A(round_reg[262]), .B(n25451), .Z(n25449) );
  XOR U26293 ( .A(round_reg[902]), .B(round_reg[582]), .Z(n25451) );
  XOR U26294 ( .A(n11180), .B(n25452), .Z(n25097) );
  XOR U26295 ( .A(n11064), .B(n13903), .Z(n25452) );
  XNOR U26296 ( .A(n25453), .B(n16158), .Z(n13903) );
  XOR U26297 ( .A(n23758), .B(n16476), .Z(n16158) );
  XNOR U26298 ( .A(n20076), .B(n20020), .Z(n16476) );
  XNOR U26299 ( .A(n25454), .B(n25455), .Z(n20020) );
  XNOR U26300 ( .A(n19453), .B(n16544), .Z(n25455) );
  XNOR U26301 ( .A(n25456), .B(n25457), .Z(n16544) );
  ANDN U26302 ( .B(n21084), .A(n19565), .Z(n25456) );
  XOR U26303 ( .A(round_reg[221]), .B(n24887), .Z(n19565) );
  XOR U26304 ( .A(round_reg[630]), .B(n22278), .Z(n21084) );
  XNOR U26305 ( .A(n25458), .B(n21486), .Z(n19453) );
  ANDN U26306 ( .B(n21089), .A(n21090), .Z(n25458) );
  XOR U26307 ( .A(round_reg[269]), .B(n24214), .Z(n21090) );
  XOR U26308 ( .A(n25459), .B(n25460), .Z(n24214) );
  XOR U26309 ( .A(round_reg[343]), .B(n22635), .Z(n21089) );
  XOR U26310 ( .A(n18380), .B(n25463), .Z(n25454) );
  XOR U26311 ( .A(n18482), .B(n19706), .Z(n25463) );
  XOR U26312 ( .A(n25464), .B(n21525), .Z(n19706) );
  NOR U26313 ( .A(n21087), .B(n19789), .Z(n25464) );
  XOR U26314 ( .A(round_reg[17]), .B(n22829), .Z(n19789) );
  XNOR U26315 ( .A(n25465), .B(n25466), .Z(n22829) );
  XOR U26316 ( .A(round_reg[394]), .B(n24268), .Z(n21087) );
  IV U26317 ( .A(n22839), .Z(n24268) );
  XOR U26318 ( .A(n25469), .B(n25470), .Z(n18482) );
  ANDN U26319 ( .B(n25471), .A(n19572), .Z(n25469) );
  XOR U26320 ( .A(round_reg[103]), .B(n24450), .Z(n19572) );
  XNOR U26321 ( .A(n25472), .B(n21491), .Z(n18380) );
  XOR U26322 ( .A(round_reg[162]), .B(n24787), .Z(n19965) );
  XOR U26323 ( .A(round_reg[562]), .B(n24023), .Z(n21093) );
  XOR U26324 ( .A(n25473), .B(n25474), .Z(n24023) );
  XOR U26325 ( .A(n25475), .B(n25476), .Z(n20076) );
  XOR U26326 ( .A(n19489), .B(n18043), .Z(n25476) );
  XNOR U26327 ( .A(n25477), .B(n23099), .Z(n18043) );
  ANDN U26328 ( .B(n23100), .A(n20991), .Z(n25477) );
  XOR U26329 ( .A(round_reg[1065]), .B(n23876), .Z(n23100) );
  XOR U26330 ( .A(n25478), .B(n23106), .Z(n19489) );
  ANDN U26331 ( .B(n23107), .A(n21000), .Z(n25478) );
  XOR U26332 ( .A(round_reg[854]), .B(n22691), .Z(n21000) );
  XOR U26333 ( .A(round_reg[1276]), .B(n25177), .Z(n23107) );
  XOR U26334 ( .A(n18813), .B(n25479), .Z(n25475) );
  XOR U26335 ( .A(n21479), .B(n19397), .Z(n25479) );
  XNOR U26336 ( .A(n25480), .B(n23103), .Z(n19397) );
  ANDN U26337 ( .B(n23104), .A(n20995), .Z(n25480) );
  XOR U26338 ( .A(round_reg[711]), .B(n21316), .Z(n20995) );
  XNOR U26339 ( .A(n25080), .B(n25481), .Z(n21316) );
  XNOR U26340 ( .A(n25482), .B(n25483), .Z(n25080) );
  XNOR U26341 ( .A(round_reg[326]), .B(round_reg[1286]), .Z(n25483) );
  XOR U26342 ( .A(round_reg[646]), .B(n25484), .Z(n25482) );
  XOR U26343 ( .A(round_reg[966]), .B(round_reg[6]), .Z(n25484) );
  XOR U26344 ( .A(round_reg[1114]), .B(n23149), .Z(n23104) );
  IV U26345 ( .A(n23672), .Z(n23149) );
  XOR U26346 ( .A(n25485), .B(n25486), .Z(n23672) );
  XNOR U26347 ( .A(n25487), .B(n23096), .Z(n21479) );
  ANDN U26348 ( .B(n23097), .A(n21004), .Z(n25487) );
  XNOR U26349 ( .A(round_reg[821]), .B(n25340), .Z(n21004) );
  XOR U26350 ( .A(n25488), .B(n25489), .Z(n25340) );
  XOR U26351 ( .A(round_reg[1204]), .B(n22513), .Z(n23097) );
  XNOR U26352 ( .A(n25490), .B(n23109), .Z(n18813) );
  ANDN U26353 ( .B(n23110), .A(n21008), .Z(n25490) );
  XNOR U26354 ( .A(n25491), .B(n23110), .Z(n23758) );
  XOR U26355 ( .A(round_reg[972]), .B(n22368), .Z(n23110) );
  XOR U26356 ( .A(n25492), .B(n24974), .Z(n22368) );
  XNOR U26357 ( .A(n25493), .B(n25494), .Z(n24974) );
  XNOR U26358 ( .A(round_reg[1356]), .B(round_reg[1036]), .Z(n25494) );
  XOR U26359 ( .A(round_reg[396]), .B(n25495), .Z(n25493) );
  XOR U26360 ( .A(round_reg[76]), .B(round_reg[716]), .Z(n25495) );
  ANDN U26361 ( .B(n21008), .A(n21009), .Z(n25491) );
  XNOR U26362 ( .A(round_reg[925]), .B(n24463), .Z(n21008) );
  IV U26363 ( .A(n24171), .Z(n24463) );
  XNOR U26364 ( .A(n25496), .B(n25497), .Z(n25230) );
  XNOR U26365 ( .A(round_reg[1500]), .B(round_reg[1180]), .Z(n25497) );
  XOR U26366 ( .A(round_reg[220]), .B(n25498), .Z(n25496) );
  XOR U26367 ( .A(round_reg[860]), .B(round_reg[540]), .Z(n25498) );
  ANDN U26368 ( .B(n13304), .A(n13302), .Z(n25453) );
  XNOR U26369 ( .A(n15913), .B(n23083), .Z(n13302) );
  XNOR U26370 ( .A(n25500), .B(n21020), .Z(n23083) );
  XNOR U26371 ( .A(round_reg[271]), .B(n22802), .Z(n23113) );
  XOR U26372 ( .A(n24742), .B(n21435), .Z(n15913) );
  XNOR U26373 ( .A(n25501), .B(n25502), .Z(n21435) );
  XOR U26374 ( .A(n18519), .B(n18961), .Z(n25502) );
  XOR U26375 ( .A(n25503), .B(n21001), .Z(n18961) );
  XOR U26376 ( .A(round_reg[465]), .B(n22790), .Z(n21001) );
  XOR U26377 ( .A(n25504), .B(n25505), .Z(n22790) );
  XOR U26378 ( .A(round_reg[1285]), .B(n23895), .Z(n23106) );
  IV U26379 ( .A(n25029), .Z(n23895) );
  XNOR U26380 ( .A(n25506), .B(n25507), .Z(n25342) );
  XNOR U26381 ( .A(round_reg[1349]), .B(round_reg[1029]), .Z(n25507) );
  XOR U26382 ( .A(round_reg[389]), .B(n25508), .Z(n25506) );
  XOR U26383 ( .A(round_reg[709]), .B(round_reg[69]), .Z(n25508) );
  XOR U26384 ( .A(n25509), .B(n25510), .Z(n25287) );
  XNOR U26385 ( .A(round_reg[1540]), .B(round_reg[1220]), .Z(n25510) );
  XOR U26386 ( .A(round_reg[260]), .B(n25511), .Z(n25509) );
  XOR U26387 ( .A(round_reg[900]), .B(round_reg[580]), .Z(n25511) );
  XNOR U26388 ( .A(round_reg[104]), .B(n25512), .Z(n21002) );
  XNOR U26389 ( .A(n25513), .B(n20992), .Z(n18519) );
  XOR U26390 ( .A(round_reg[631]), .B(n23789), .Z(n20992) );
  ANDN U26391 ( .B(n20993), .A(n23099), .Z(n25513) );
  XOR U26392 ( .A(round_reg[1442]), .B(n24787), .Z(n23099) );
  XOR U26393 ( .A(round_reg[222]), .B(n22751), .Z(n20993) );
  XOR U26394 ( .A(n18853), .B(n25514), .Z(n25501) );
  XNOR U26395 ( .A(n19559), .B(n15842), .Z(n25514) );
  XNOR U26396 ( .A(n25515), .B(n21006), .Z(n15842) );
  XNOR U26397 ( .A(round_reg[395]), .B(n23270), .Z(n21006) );
  IV U26398 ( .A(n24906), .Z(n23270) );
  ANDN U26399 ( .B(n21005), .A(n23096), .Z(n25515) );
  XOR U26400 ( .A(round_reg[1568]), .B(n24272), .Z(n23096) );
  XOR U26401 ( .A(n24850), .B(n25187), .Z(n24272) );
  XOR U26402 ( .A(n25516), .B(n25517), .Z(n25187) );
  XNOR U26403 ( .A(round_reg[1503]), .B(round_reg[1183]), .Z(n25517) );
  XOR U26404 ( .A(round_reg[223]), .B(n25518), .Z(n25516) );
  XOR U26405 ( .A(round_reg[863]), .B(round_reg[543]), .Z(n25518) );
  XNOR U26406 ( .A(n25519), .B(n25520), .Z(n24850) );
  XNOR U26407 ( .A(round_reg[32]), .B(round_reg[1312]), .Z(n25520) );
  XOR U26408 ( .A(round_reg[352]), .B(n25521), .Z(n25519) );
  XOR U26409 ( .A(round_reg[992]), .B(round_reg[672]), .Z(n25521) );
  XOR U26410 ( .A(round_reg[18]), .B(n21186), .Z(n21005) );
  XOR U26411 ( .A(n25522), .B(n25236), .Z(n21186) );
  XNOR U26412 ( .A(n25523), .B(n25524), .Z(n25236) );
  XNOR U26413 ( .A(round_reg[1362]), .B(round_reg[1042]), .Z(n25524) );
  XOR U26414 ( .A(round_reg[402]), .B(n25525), .Z(n25523) );
  XOR U26415 ( .A(round_reg[82]), .B(round_reg[722]), .Z(n25525) );
  XNOR U26416 ( .A(n25526), .B(n20997), .Z(n19559) );
  XOR U26417 ( .A(round_reg[344]), .B(n23995), .Z(n20997) );
  XOR U26418 ( .A(n25527), .B(n25528), .Z(n23995) );
  NOR U26419 ( .A(n23103), .B(n20996), .Z(n25526) );
  XNOR U26420 ( .A(round_reg[270]), .B(n24636), .Z(n20996) );
  XOR U26421 ( .A(round_reg[1503]), .B(n24769), .Z(n23103) );
  IV U26422 ( .A(n22439), .Z(n24769) );
  XOR U26423 ( .A(n25529), .B(n25070), .Z(n22439) );
  XOR U26424 ( .A(n25530), .B(n25531), .Z(n25070) );
  XNOR U26425 ( .A(round_reg[1567]), .B(round_reg[1247]), .Z(n25531) );
  XOR U26426 ( .A(round_reg[287]), .B(n25532), .Z(n25530) );
  XOR U26427 ( .A(round_reg[927]), .B(round_reg[607]), .Z(n25532) );
  XNOR U26428 ( .A(n25533), .B(n21009), .Z(n18853) );
  XOR U26429 ( .A(round_reg[563]), .B(n24518), .Z(n21009) );
  ANDN U26430 ( .B(n21010), .A(n23109), .Z(n25533) );
  XOR U26431 ( .A(round_reg[1348]), .B(n23721), .Z(n23109) );
  XOR U26432 ( .A(round_reg[163]), .B(n23396), .Z(n21010) );
  XOR U26433 ( .A(n25534), .B(n25535), .Z(n23396) );
  XOR U26434 ( .A(n25536), .B(n25537), .Z(n24742) );
  XNOR U26435 ( .A(n16560), .B(n17410), .Z(n25537) );
  XOR U26436 ( .A(n25538), .B(n21016), .Z(n17410) );
  XNOR U26437 ( .A(round_reg[1066]), .B(n23528), .Z(n21016) );
  XOR U26438 ( .A(n24775), .B(n24329), .Z(n23528) );
  XNOR U26439 ( .A(n25539), .B(n25540), .Z(n24329) );
  XNOR U26440 ( .A(round_reg[1450]), .B(round_reg[1130]), .Z(n25540) );
  XOR U26441 ( .A(round_reg[170]), .B(n25541), .Z(n25539) );
  XOR U26442 ( .A(round_reg[810]), .B(round_reg[490]), .Z(n25541) );
  XOR U26443 ( .A(n25542), .B(n25543), .Z(n24775) );
  XNOR U26444 ( .A(round_reg[1321]), .B(round_reg[1001]), .Z(n25543) );
  XOR U26445 ( .A(round_reg[361]), .B(n25544), .Z(n25542) );
  XOR U26446 ( .A(round_reg[681]), .B(round_reg[41]), .Z(n25544) );
  AND U26447 ( .A(n21502), .B(n23087), .Z(n25538) );
  IV U26448 ( .A(n21015), .Z(n23087) );
  XNOR U26449 ( .A(round_reg[698]), .B(n24578), .Z(n21015) );
  XNOR U26450 ( .A(round_reg[632]), .B(n21775), .Z(n21502) );
  XNOR U26451 ( .A(n25545), .B(n21019), .Z(n16560) );
  XOR U26452 ( .A(round_reg[1115]), .B(n23411), .Z(n21019) );
  XNOR U26453 ( .A(n25546), .B(n25547), .Z(n23411) );
  AND U26454 ( .A(n21020), .B(n23112), .Z(n25545) );
  XNOR U26455 ( .A(round_reg[345]), .B(n21198), .Z(n23112) );
  XNOR U26456 ( .A(n25548), .B(n25549), .Z(n25297) );
  XNOR U26457 ( .A(round_reg[1560]), .B(round_reg[1240]), .Z(n25549) );
  XOR U26458 ( .A(round_reg[280]), .B(n25550), .Z(n25548) );
  XOR U26459 ( .A(round_reg[920]), .B(round_reg[600]), .Z(n25550) );
  XOR U26460 ( .A(n25551), .B(n25552), .Z(n25486) );
  XNOR U26461 ( .A(round_reg[1369]), .B(round_reg[1049]), .Z(n25552) );
  XOR U26462 ( .A(round_reg[409]), .B(n25553), .Z(n25551) );
  XOR U26463 ( .A(round_reg[89]), .B(round_reg[729]), .Z(n25553) );
  XOR U26464 ( .A(round_reg[712]), .B(n24284), .Z(n21020) );
  XNOR U26465 ( .A(n25554), .B(n25555), .Z(n24941) );
  XNOR U26466 ( .A(round_reg[136]), .B(round_reg[1096]), .Z(n25555) );
  XOR U26467 ( .A(round_reg[1416]), .B(n25556), .Z(n25554) );
  XOR U26468 ( .A(round_reg[776]), .B(round_reg[456]), .Z(n25556) );
  XNOR U26469 ( .A(n25557), .B(n25558), .Z(n24929) );
  XNOR U26470 ( .A(round_reg[327]), .B(round_reg[1287]), .Z(n25558) );
  XOR U26471 ( .A(round_reg[647]), .B(n25559), .Z(n25557) );
  XOR U26472 ( .A(round_reg[967]), .B(round_reg[7]), .Z(n25559) );
  XOR U26473 ( .A(n16463), .B(n25560), .Z(n25536) );
  XNOR U26474 ( .A(n16061), .B(n20987), .Z(n25560) );
  XNOR U26475 ( .A(n25561), .B(n21026), .Z(n20987) );
  XNOR U26476 ( .A(round_reg[1205]), .B(n25242), .Z(n21026) );
  IV U26477 ( .A(n23871), .Z(n25242) );
  NOR U26478 ( .A(n23089), .B(n21025), .Z(n25561) );
  XNOR U26479 ( .A(round_reg[822]), .B(n24514), .Z(n21025) );
  IV U26480 ( .A(n25278), .Z(n24514) );
  XNOR U26481 ( .A(n25562), .B(n25563), .Z(n25278) );
  IV U26482 ( .A(n21508), .Z(n23089) );
  XNOR U26483 ( .A(round_reg[396]), .B(n24490), .Z(n21508) );
  XNOR U26484 ( .A(n25564), .B(n21029), .Z(n16061) );
  XOR U26485 ( .A(round_reg[1277]), .B(n24440), .Z(n21029) );
  XOR U26486 ( .A(n25565), .B(n25566), .Z(n24440) );
  ANDN U26487 ( .B(n21030), .A(n21499), .Z(n25564) );
  XOR U26488 ( .A(round_reg[466]), .B(n23295), .Z(n21499) );
  XOR U26489 ( .A(round_reg[855]), .B(n24139), .Z(n21030) );
  XNOR U26490 ( .A(n25528), .B(n25402), .Z(n24139) );
  XNOR U26491 ( .A(n25567), .B(n25568), .Z(n25402) );
  XNOR U26492 ( .A(round_reg[1430]), .B(round_reg[1110]), .Z(n25568) );
  XOR U26493 ( .A(round_reg[150]), .B(n25569), .Z(n25567) );
  XOR U26494 ( .A(round_reg[790]), .B(round_reg[470]), .Z(n25569) );
  XNOR U26495 ( .A(n25570), .B(n25571), .Z(n25528) );
  XNOR U26496 ( .A(round_reg[1559]), .B(round_reg[1239]), .Z(n25571) );
  XOR U26497 ( .A(round_reg[279]), .B(n25572), .Z(n25570) );
  XOR U26498 ( .A(round_reg[919]), .B(round_reg[599]), .Z(n25572) );
  XNOR U26499 ( .A(n25573), .B(n23752), .Z(n16463) );
  XOR U26500 ( .A(round_reg[973]), .B(n24515), .Z(n23752) );
  ANDN U26501 ( .B(n21511), .A(n23092), .Z(n25573) );
  XNOR U26502 ( .A(round_reg[926]), .B(n23464), .Z(n23092) );
  XNOR U26503 ( .A(round_reg[564]), .B(n22513), .Z(n21511) );
  IV U26504 ( .A(n25574), .Z(n22513) );
  XNOR U26505 ( .A(n18485), .B(n22291), .Z(n13304) );
  XNOR U26506 ( .A(n25575), .B(n24624), .Z(n22291) );
  ANDN U26507 ( .B(n22885), .A(n22886), .Z(n25575) );
  IV U26508 ( .A(n25576), .Z(n22885) );
  XOR U26509 ( .A(n23219), .B(n21632), .Z(n18485) );
  XNOR U26510 ( .A(n25577), .B(n25578), .Z(n21632) );
  XNOR U26511 ( .A(n17983), .B(n22100), .Z(n25578) );
  XOR U26512 ( .A(n25579), .B(n24830), .Z(n22100) );
  XNOR U26513 ( .A(round_reg[126]), .B(n23561), .Z(n24830) );
  XOR U26514 ( .A(n25565), .B(n25580), .Z(n23561) );
  XOR U26515 ( .A(n25581), .B(n25582), .Z(n25565) );
  XNOR U26516 ( .A(round_reg[1341]), .B(round_reg[1021]), .Z(n25582) );
  XOR U26517 ( .A(round_reg[381]), .B(n25583), .Z(n25581) );
  XOR U26518 ( .A(round_reg[701]), .B(round_reg[61]), .Z(n25583) );
  ANDN U26519 ( .B(n22311), .A(n22312), .Z(n25579) );
  XOR U26520 ( .A(round_reg[1234]), .B(n24504), .Z(n22312) );
  XNOR U26521 ( .A(n25505), .B(n24938), .Z(n24504) );
  XNOR U26522 ( .A(n25584), .B(n25585), .Z(n24938) );
  XNOR U26523 ( .A(round_reg[18]), .B(round_reg[1298]), .Z(n25585) );
  XOR U26524 ( .A(round_reg[338]), .B(n25586), .Z(n25584) );
  XOR U26525 ( .A(round_reg[978]), .B(round_reg[658]), .Z(n25586) );
  XNOR U26526 ( .A(n25587), .B(n25588), .Z(n25505) );
  XNOR U26527 ( .A(round_reg[1489]), .B(round_reg[1169]), .Z(n25588) );
  XOR U26528 ( .A(round_reg[209]), .B(n25589), .Z(n25587) );
  XOR U26529 ( .A(round_reg[849]), .B(round_reg[529]), .Z(n25589) );
  XOR U26530 ( .A(round_reg[1307]), .B(n23386), .Z(n22311) );
  XNOR U26531 ( .A(n25590), .B(n22139), .Z(n17983) );
  XNOR U26532 ( .A(round_reg[292]), .B(n25023), .Z(n22139) );
  ANDN U26533 ( .B(n22138), .A(n22318), .Z(n25590) );
  XOR U26534 ( .A(round_reg[1136]), .B(n23963), .Z(n22318) );
  IV U26535 ( .A(n25068), .Z(n23963) );
  XNOR U26536 ( .A(n25591), .B(n24896), .Z(n25068) );
  XNOR U26537 ( .A(n25592), .B(n25593), .Z(n24896) );
  XNOR U26538 ( .A(round_reg[1520]), .B(round_reg[1200]), .Z(n25593) );
  XOR U26539 ( .A(round_reg[240]), .B(n25594), .Z(n25592) );
  XOR U26540 ( .A(round_reg[880]), .B(round_reg[560]), .Z(n25594) );
  XNOR U26541 ( .A(round_reg[1525]), .B(n23871), .Z(n22138) );
  XNOR U26542 ( .A(n19461), .B(n25595), .Z(n25577) );
  XOR U26543 ( .A(n17682), .B(n17533), .Z(n25595) );
  XNOR U26544 ( .A(n25596), .B(n22135), .Z(n17533) );
  XOR U26545 ( .A(round_reg[40]), .B(n23488), .Z(n22135) );
  IV U26546 ( .A(n24687), .Z(n23488) );
  XOR U26547 ( .A(n25597), .B(n25598), .Z(n24687) );
  ANDN U26548 ( .B(n22134), .A(n22307), .Z(n25596) );
  XOR U26549 ( .A(round_reg[1162]), .B(n22366), .Z(n22307) );
  XOR U26550 ( .A(round_reg[1590]), .B(n22278), .Z(n22134) );
  XOR U26551 ( .A(n25599), .B(n25600), .Z(n25091) );
  XNOR U26552 ( .A(round_reg[1334]), .B(round_reg[1014]), .Z(n25600) );
  XOR U26553 ( .A(round_reg[374]), .B(n25601), .Z(n25599) );
  XOR U26554 ( .A(round_reg[694]), .B(round_reg[54]), .Z(n25601) );
  XNOR U26555 ( .A(n25602), .B(n25603), .Z(n25489) );
  XNOR U26556 ( .A(round_reg[1525]), .B(round_reg[1205]), .Z(n25603) );
  XOR U26557 ( .A(round_reg[245]), .B(n25604), .Z(n25602) );
  XOR U26558 ( .A(round_reg[885]), .B(round_reg[565]), .Z(n25604) );
  XOR U26559 ( .A(n25605), .B(n22128), .Z(n17682) );
  XNOR U26560 ( .A(round_reg[244]), .B(n25574), .Z(n22128) );
  XOR U26561 ( .A(n25606), .B(n25607), .Z(n25574) );
  ANDN U26562 ( .B(n22129), .A(n22315), .Z(n25605) );
  XNOR U26563 ( .A(round_reg[1087]), .B(n25608), .Z(n22315) );
  XOR U26564 ( .A(round_reg[1464]), .B(n22642), .Z(n22129) );
  XOR U26565 ( .A(n25227), .B(n25609), .Z(n22642) );
  XOR U26566 ( .A(n25610), .B(n25611), .Z(n25227) );
  XNOR U26567 ( .A(round_reg[1528]), .B(round_reg[1208]), .Z(n25611) );
  XOR U26568 ( .A(round_reg[248]), .B(n25612), .Z(n25610) );
  XOR U26569 ( .A(round_reg[888]), .B(round_reg[568]), .Z(n25612) );
  XNOR U26570 ( .A(n25613), .B(n22125), .Z(n19461) );
  XOR U26571 ( .A(round_reg[185]), .B(n25151), .Z(n22125) );
  ANDN U26572 ( .B(n22124), .A(n22304), .Z(n25613) );
  XOR U26573 ( .A(round_reg[994]), .B(n23405), .Z(n22304) );
  XNOR U26574 ( .A(n25534), .B(n25207), .Z(n23405) );
  XOR U26575 ( .A(n25614), .B(n25615), .Z(n25207) );
  XNOR U26576 ( .A(round_reg[1569]), .B(round_reg[1249]), .Z(n25615) );
  XOR U26577 ( .A(round_reg[289]), .B(n25616), .Z(n25614) );
  XOR U26578 ( .A(round_reg[929]), .B(round_reg[609]), .Z(n25616) );
  XOR U26579 ( .A(n25617), .B(n25618), .Z(n25534) );
  XNOR U26580 ( .A(round_reg[1378]), .B(round_reg[1058]), .Z(n25618) );
  XOR U26581 ( .A(round_reg[418]), .B(n25619), .Z(n25617) );
  XOR U26582 ( .A(round_reg[98]), .B(round_reg[738]), .Z(n25619) );
  XOR U26583 ( .A(round_reg[1370]), .B(n24714), .Z(n22124) );
  IV U26584 ( .A(n24227), .Z(n24714) );
  XOR U26585 ( .A(n25620), .B(n25621), .Z(n24227) );
  XOR U26586 ( .A(n25622), .B(n25623), .Z(n23219) );
  XOR U26587 ( .A(n17068), .B(n20012), .Z(n25623) );
  XNOR U26588 ( .A(n25624), .B(n24617), .Z(n20012) );
  ANDN U26589 ( .B(n22288), .A(n22289), .Z(n25624) );
  XNOR U26590 ( .A(round_reg[245]), .B(n23871), .Z(n22289) );
  XNOR U26591 ( .A(n24917), .B(n25373), .Z(n23871) );
  XNOR U26592 ( .A(n25625), .B(n25626), .Z(n25373) );
  XNOR U26593 ( .A(round_reg[1589]), .B(round_reg[1269]), .Z(n25626) );
  XOR U26594 ( .A(round_reg[309]), .B(n25627), .Z(n25625) );
  XOR U26595 ( .A(round_reg[949]), .B(round_reg[629]), .Z(n25627) );
  XOR U26596 ( .A(n25628), .B(n25629), .Z(n24917) );
  XNOR U26597 ( .A(round_reg[1460]), .B(round_reg[1140]), .Z(n25629) );
  XOR U26598 ( .A(round_reg[180]), .B(n25630), .Z(n25628) );
  XOR U26599 ( .A(round_reg[820]), .B(round_reg[500]), .Z(n25630) );
  XOR U26600 ( .A(round_reg[590]), .B(n24636), .Z(n22288) );
  IV U26601 ( .A(n23497), .Z(n24636) );
  XOR U26602 ( .A(n25260), .B(n24973), .Z(n23497) );
  XNOR U26603 ( .A(n25631), .B(n25632), .Z(n24973) );
  XNOR U26604 ( .A(round_reg[1485]), .B(round_reg[1165]), .Z(n25632) );
  XOR U26605 ( .A(round_reg[205]), .B(n25633), .Z(n25631) );
  XOR U26606 ( .A(round_reg[845]), .B(round_reg[525]), .Z(n25633) );
  XNOR U26607 ( .A(n25634), .B(n25635), .Z(n25260) );
  XNOR U26608 ( .A(round_reg[14]), .B(round_reg[1294]), .Z(n25635) );
  XOR U26609 ( .A(round_reg[334]), .B(n25636), .Z(n25634) );
  XOR U26610 ( .A(round_reg[974]), .B(round_reg[654]), .Z(n25636) );
  XNOR U26611 ( .A(n25637), .B(n24619), .Z(n17068) );
  AND U26612 ( .A(n22298), .B(n22300), .Z(n25637) );
  XOR U26613 ( .A(round_reg[293]), .B(n25167), .Z(n22300) );
  IV U26614 ( .A(n25042), .Z(n25167) );
  XOR U26615 ( .A(round_reg[367]), .B(n24564), .Z(n22298) );
  XNOR U26616 ( .A(n25591), .B(n24976), .Z(n24564) );
  XOR U26617 ( .A(n25638), .B(n25639), .Z(n24976) );
  XNOR U26618 ( .A(round_reg[1582]), .B(round_reg[1262]), .Z(n25639) );
  XOR U26619 ( .A(round_reg[302]), .B(n25640), .Z(n25638) );
  XOR U26620 ( .A(round_reg[942]), .B(round_reg[622]), .Z(n25640) );
  XOR U26621 ( .A(n25641), .B(n25642), .Z(n25591) );
  XNOR U26622 ( .A(round_reg[111]), .B(round_reg[1071]), .Z(n25642) );
  XOR U26623 ( .A(round_reg[1391]), .B(n25643), .Z(n25641) );
  XOR U26624 ( .A(round_reg[751]), .B(round_reg[431]), .Z(n25643) );
  XNOR U26625 ( .A(n17244), .B(n25644), .Z(n25622) );
  XNOR U26626 ( .A(n21124), .B(n17443), .Z(n25644) );
  XNOR U26627 ( .A(n25645), .B(n24622), .Z(n17443) );
  ANDN U26628 ( .B(n22294), .A(n22295), .Z(n25645) );
  XOR U26629 ( .A(round_reg[41]), .B(n24221), .Z(n22295) );
  XNOR U26630 ( .A(round_reg[418]), .B(n23887), .Z(n22294) );
  XNOR U26631 ( .A(n25414), .B(n25183), .Z(n23887) );
  XNOR U26632 ( .A(n25646), .B(n25647), .Z(n25183) );
  XNOR U26633 ( .A(round_reg[1442]), .B(round_reg[1122]), .Z(n25647) );
  XOR U26634 ( .A(round_reg[162]), .B(n25648), .Z(n25646) );
  XOR U26635 ( .A(round_reg[802]), .B(round_reg[482]), .Z(n25648) );
  XOR U26636 ( .A(n25649), .B(n25650), .Z(n25414) );
  XNOR U26637 ( .A(round_reg[33]), .B(round_reg[1313]), .Z(n25650) );
  XOR U26638 ( .A(round_reg[353]), .B(n25651), .Z(n25649) );
  XOR U26639 ( .A(round_reg[993]), .B(round_reg[673]), .Z(n25651) );
  XNOR U26640 ( .A(n25652), .B(n24625), .Z(n21124) );
  AND U26641 ( .A(n24624), .B(n25576), .Z(n25652) );
  XOR U26642 ( .A(round_reg[127]), .B(n25608), .Z(n25576) );
  IV U26643 ( .A(n22371), .Z(n25608) );
  XNOR U26644 ( .A(n25654), .B(n25655), .Z(n24933) );
  XNOR U26645 ( .A(round_reg[1471]), .B(round_reg[1151]), .Z(n25655) );
  XOR U26646 ( .A(round_reg[191]), .B(n25656), .Z(n25654) );
  XOR U26647 ( .A(round_reg[831]), .B(round_reg[511]), .Z(n25656) );
  XOR U26648 ( .A(round_reg[488]), .B(n22821), .Z(n24624) );
  XNOR U26649 ( .A(n25657), .B(n25658), .Z(n24776) );
  XNOR U26650 ( .A(round_reg[1512]), .B(round_reg[1192]), .Z(n25658) );
  XOR U26651 ( .A(round_reg[232]), .B(n25659), .Z(n25657) );
  XOR U26652 ( .A(round_reg[872]), .B(round_reg[552]), .Z(n25659) );
  XNOR U26653 ( .A(n25661), .B(n24627), .Z(n17244) );
  ANDN U26654 ( .B(n22284), .A(n22285), .Z(n25661) );
  XNOR U26655 ( .A(round_reg[186]), .B(n24451), .Z(n22285) );
  XOR U26656 ( .A(round_reg[522]), .B(n22366), .Z(n22284) );
  XNOR U26657 ( .A(n25662), .B(n25663), .Z(n22366) );
  XNOR U26658 ( .A(n25664), .B(n14675), .Z(n11064) );
  XNOR U26659 ( .A(n20571), .B(n18270), .Z(n14675) );
  XOR U26660 ( .A(n22146), .B(n20688), .Z(n18270) );
  XNOR U26661 ( .A(n25665), .B(n25666), .Z(n20688) );
  XOR U26662 ( .A(n13895), .B(n18247), .Z(n25666) );
  XNOR U26663 ( .A(n25667), .B(n23237), .Z(n18247) );
  XNOR U26664 ( .A(round_reg[1072]), .B(n24770), .Z(n23237) );
  AND U26665 ( .A(n18779), .B(n20376), .Z(n25667) );
  XOR U26666 ( .A(round_reg[640]), .B(n23811), .Z(n20376) );
  XOR U26667 ( .A(round_reg[638]), .B(n23877), .Z(n18779) );
  XNOR U26668 ( .A(n25668), .B(n20129), .Z(n13895) );
  XOR U26669 ( .A(round_reg[1121]), .B(n24694), .Z(n20129) );
  ANDN U26670 ( .B(n20130), .A(n20371), .Z(n25668) );
  XOR U26671 ( .A(round_reg[351]), .B(n23325), .Z(n20371) );
  XNOR U26672 ( .A(n25669), .B(n25094), .Z(n23325) );
  XOR U26673 ( .A(n25670), .B(n25671), .Z(n25094) );
  XNOR U26674 ( .A(round_reg[1375]), .B(round_reg[1055]), .Z(n25671) );
  XOR U26675 ( .A(round_reg[415]), .B(n25672), .Z(n25670) );
  XOR U26676 ( .A(round_reg[95]), .B(round_reg[735]), .Z(n25672) );
  XOR U26677 ( .A(round_reg[718]), .B(n23595), .Z(n20130) );
  XNOR U26678 ( .A(n25673), .B(n25674), .Z(n25460) );
  XNOR U26679 ( .A(round_reg[13]), .B(round_reg[1293]), .Z(n25674) );
  XOR U26680 ( .A(round_reg[333]), .B(n25675), .Z(n25673) );
  XOR U26681 ( .A(round_reg[973]), .B(round_reg[653]), .Z(n25675) );
  XNOR U26682 ( .A(n17366), .B(n25677), .Z(n25665) );
  XNOR U26683 ( .A(n17880), .B(n18283), .Z(n25677) );
  XNOR U26684 ( .A(n25678), .B(n20120), .Z(n18283) );
  XNOR U26685 ( .A(round_reg[1211]), .B(n21617), .Z(n20120) );
  AND U26686 ( .A(n20121), .B(n18841), .Z(n25678) );
  XOR U26687 ( .A(round_reg[402]), .B(n25062), .Z(n18841) );
  IV U26688 ( .A(n21786), .Z(n25062) );
  XOR U26689 ( .A(round_reg[828]), .B(n23323), .Z(n20121) );
  XNOR U26690 ( .A(n25679), .B(n23263), .Z(n17880) );
  IV U26691 ( .A(n20125), .Z(n23263) );
  XOR U26692 ( .A(round_reg[1219]), .B(n25133), .Z(n20125) );
  AND U26693 ( .A(n18775), .B(n20126), .Z(n25679) );
  XOR U26694 ( .A(round_reg[861]), .B(n24887), .Z(n20126) );
  XOR U26695 ( .A(round_reg[472]), .B(n25011), .Z(n18775) );
  XOR U26696 ( .A(n25682), .B(n25462), .Z(n25011) );
  XOR U26697 ( .A(n25683), .B(n25684), .Z(n25462) );
  XNOR U26698 ( .A(round_reg[1367]), .B(round_reg[1047]), .Z(n25684) );
  XOR U26699 ( .A(round_reg[407]), .B(n25685), .Z(n25683) );
  XOR U26700 ( .A(round_reg[87]), .B(round_reg[727]), .Z(n25685) );
  XNOR U26701 ( .A(n25686), .B(n20118), .Z(n17366) );
  XNOR U26702 ( .A(round_reg[979]), .B(n23744), .Z(n20118) );
  XOR U26703 ( .A(n24717), .B(n25110), .Z(n23744) );
  XNOR U26704 ( .A(n25687), .B(n25688), .Z(n25110) );
  XNOR U26705 ( .A(round_reg[1554]), .B(round_reg[1234]), .Z(n25688) );
  XOR U26706 ( .A(round_reg[274]), .B(n25689), .Z(n25687) );
  XOR U26707 ( .A(round_reg[914]), .B(round_reg[594]), .Z(n25689) );
  XOR U26708 ( .A(n25690), .B(n25691), .Z(n24717) );
  XNOR U26709 ( .A(round_reg[1363]), .B(round_reg[1043]), .Z(n25691) );
  XOR U26710 ( .A(round_reg[403]), .B(n25692), .Z(n25690) );
  XOR U26711 ( .A(round_reg[83]), .B(round_reg[723]), .Z(n25692) );
  AND U26712 ( .A(n20117), .B(n19675), .Z(n25686) );
  XOR U26713 ( .A(round_reg[570]), .B(n23249), .Z(n19675) );
  XOR U26714 ( .A(round_reg[932]), .B(n25023), .Z(n20117) );
  XOR U26715 ( .A(n25693), .B(n25694), .Z(n22146) );
  XNOR U26716 ( .A(n18821), .B(n18201), .Z(n25694) );
  XOR U26717 ( .A(n25695), .B(n21615), .Z(n18201) );
  XOR U26718 ( .A(round_reg[171]), .B(n23389), .Z(n21615) );
  XOR U26719 ( .A(n25696), .B(n25127), .Z(n23389) );
  XNOR U26720 ( .A(n25697), .B(n25698), .Z(n25127) );
  XNOR U26721 ( .A(round_reg[1515]), .B(round_reg[1195]), .Z(n25698) );
  XOR U26722 ( .A(round_reg[235]), .B(n25699), .Z(n25697) );
  XOR U26723 ( .A(round_reg[875]), .B(round_reg[555]), .Z(n25699) );
  AND U26724 ( .A(n19872), .B(n25700), .Z(n25695) );
  XNOR U26725 ( .A(n25701), .B(n20113), .Z(n18821) );
  XNOR U26726 ( .A(round_reg[26]), .B(n24823), .Z(n20113) );
  AND U26727 ( .A(n20112), .B(n19885), .Z(n25701) );
  XOR U26728 ( .A(round_reg[1212]), .B(n24840), .Z(n19885) );
  IV U26729 ( .A(n23147), .Z(n24840) );
  XOR U26730 ( .A(n25284), .B(n25441), .Z(n23147) );
  XNOR U26731 ( .A(n25702), .B(n25703), .Z(n25441) );
  XNOR U26732 ( .A(round_reg[1467]), .B(round_reg[1147]), .Z(n25703) );
  XOR U26733 ( .A(round_reg[187]), .B(n25704), .Z(n25702) );
  XOR U26734 ( .A(round_reg[827]), .B(round_reg[507]), .Z(n25704) );
  XOR U26735 ( .A(n25705), .B(n25706), .Z(n25284) );
  XNOR U26736 ( .A(round_reg[1596]), .B(round_reg[1276]), .Z(n25706) );
  XOR U26737 ( .A(round_reg[316]), .B(n25707), .Z(n25705) );
  XOR U26738 ( .A(round_reg[956]), .B(round_reg[636]), .Z(n25707) );
  XOR U26739 ( .A(round_reg[1576]), .B(n24257), .Z(n20112) );
  IV U26740 ( .A(n23009), .Z(n24257) );
  XNOR U26741 ( .A(n25178), .B(n25708), .Z(n23009) );
  XOR U26742 ( .A(n25709), .B(n25710), .Z(n25178) );
  XNOR U26743 ( .A(round_reg[1511]), .B(round_reg[1191]), .Z(n25710) );
  XOR U26744 ( .A(round_reg[231]), .B(n25711), .Z(n25709) );
  XOR U26745 ( .A(round_reg[871]), .B(round_reg[551]), .Z(n25711) );
  XNOR U26746 ( .A(n17729), .B(n25712), .Z(n25693) );
  XNOR U26747 ( .A(n20098), .B(n18997), .Z(n25712) );
  XNOR U26748 ( .A(n25713), .B(n21521), .Z(n18997) );
  XNOR U26749 ( .A(round_reg[230]), .B(n23267), .Z(n21521) );
  IV U26750 ( .A(n24720), .Z(n23267) );
  XNOR U26751 ( .A(n25714), .B(n24992), .Z(n24720) );
  XNOR U26752 ( .A(n25715), .B(n25716), .Z(n24992) );
  XNOR U26753 ( .A(round_reg[1445]), .B(round_reg[1125]), .Z(n25716) );
  XOR U26754 ( .A(round_reg[165]), .B(n25717), .Z(n25715) );
  XOR U26755 ( .A(round_reg[805]), .B(round_reg[485]), .Z(n25717) );
  ANDN U26756 ( .B(n19881), .A(n20576), .Z(n25713) );
  XNOR U26757 ( .A(round_reg[1450]), .B(n22274), .Z(n20576) );
  IV U26758 ( .A(n24424), .Z(n22274) );
  XOR U26759 ( .A(n24842), .B(n25718), .Z(n24424) );
  XNOR U26760 ( .A(n25719), .B(n25720), .Z(n24842) );
  XNOR U26761 ( .A(round_reg[1514]), .B(round_reg[1194]), .Z(n25720) );
  XOR U26762 ( .A(round_reg[234]), .B(n25721), .Z(n25719) );
  XOR U26763 ( .A(round_reg[874]), .B(round_reg[554]), .Z(n25721) );
  XOR U26764 ( .A(round_reg[1073]), .B(n23399), .Z(n19881) );
  IV U26765 ( .A(n24943), .Z(n23399) );
  XOR U26766 ( .A(n25473), .B(n25444), .Z(n24943) );
  XNOR U26767 ( .A(n25722), .B(n25723), .Z(n25444) );
  XNOR U26768 ( .A(round_reg[1328]), .B(round_reg[1008]), .Z(n25723) );
  XOR U26769 ( .A(round_reg[368]), .B(n25724), .Z(n25722) );
  XOR U26770 ( .A(round_reg[688]), .B(round_reg[48]), .Z(n25724) );
  XOR U26771 ( .A(n25725), .B(n25726), .Z(n25473) );
  XNOR U26772 ( .A(round_reg[1457]), .B(round_reg[1137]), .Z(n25726) );
  XOR U26773 ( .A(round_reg[177]), .B(n25727), .Z(n25725) );
  XOR U26774 ( .A(round_reg[817]), .B(round_reg[497]), .Z(n25727) );
  XNOR U26775 ( .A(n25728), .B(n20102), .Z(n20098) );
  XOR U26776 ( .A(round_reg[112]), .B(n24770), .Z(n20102) );
  AND U26777 ( .A(n20103), .B(n22752), .Z(n25728) );
  XNOR U26778 ( .A(round_reg[1220]), .B(n22983), .Z(n22752) );
  XNOR U26779 ( .A(n25729), .B(n25730), .Z(n22983) );
  XOR U26780 ( .A(round_reg[1293]), .B(n24515), .Z(n20103) );
  XOR U26781 ( .A(n25030), .B(n25118), .Z(n24515) );
  XNOR U26782 ( .A(n25731), .B(n25732), .Z(n25118) );
  XNOR U26783 ( .A(round_reg[1357]), .B(round_reg[1037]), .Z(n25732) );
  XOR U26784 ( .A(round_reg[397]), .B(n25733), .Z(n25731) );
  XOR U26785 ( .A(round_reg[77]), .B(round_reg[717]), .Z(n25733) );
  XOR U26786 ( .A(n25734), .B(n25735), .Z(n25030) );
  XNOR U26787 ( .A(round_reg[1548]), .B(round_reg[1228]), .Z(n25735) );
  XOR U26788 ( .A(round_reg[268]), .B(n25736), .Z(n25734) );
  XOR U26789 ( .A(round_reg[908]), .B(round_reg[588]), .Z(n25736) );
  XNOR U26790 ( .A(n25737), .B(n20107), .Z(n17729) );
  XNOR U26791 ( .A(round_reg[278]), .B(n22225), .Z(n20107) );
  IV U26792 ( .A(n23965), .Z(n22225) );
  XOR U26793 ( .A(n25040), .B(n24740), .Z(n23965) );
  XOR U26794 ( .A(n25738), .B(n25739), .Z(n24740) );
  XNOR U26795 ( .A(round_reg[1493]), .B(round_reg[1173]), .Z(n25739) );
  XOR U26796 ( .A(round_reg[213]), .B(n25740), .Z(n25738) );
  XOR U26797 ( .A(round_reg[853]), .B(round_reg[533]), .Z(n25740) );
  XOR U26798 ( .A(n25741), .B(n25742), .Z(n25040) );
  XNOR U26799 ( .A(round_reg[22]), .B(round_reg[1302]), .Z(n25742) );
  XOR U26800 ( .A(round_reg[342]), .B(n25743), .Z(n25741) );
  XOR U26801 ( .A(round_reg[982]), .B(round_reg[662]), .Z(n25743) );
  AND U26802 ( .A(n19877), .B(n20106), .Z(n25737) );
  XOR U26803 ( .A(round_reg[1511]), .B(n22361), .Z(n20106) );
  XOR U26804 ( .A(n25597), .B(n25744), .Z(n22361) );
  XOR U26805 ( .A(n25745), .B(n25746), .Z(n25597) );
  XNOR U26806 ( .A(round_reg[1575]), .B(round_reg[1255]), .Z(n25746) );
  XOR U26807 ( .A(round_reg[295]), .B(n25747), .Z(n25745) );
  XOR U26808 ( .A(round_reg[935]), .B(round_reg[615]), .Z(n25747) );
  XNOR U26809 ( .A(round_reg[1122]), .B(n24787), .Z(n19877) );
  IV U26810 ( .A(n24407), .Z(n24787) );
  XNOR U26811 ( .A(n25194), .B(n25748), .Z(n24407) );
  XOR U26812 ( .A(n25749), .B(n25750), .Z(n25194) );
  XNOR U26813 ( .A(round_reg[1506]), .B(round_reg[1186]), .Z(n25750) );
  XOR U26814 ( .A(round_reg[226]), .B(n25751), .Z(n25749) );
  XOR U26815 ( .A(round_reg[866]), .B(round_reg[546]), .Z(n25751) );
  XOR U26816 ( .A(n25752), .B(n21618), .Z(n20571) );
  IV U26817 ( .A(n25700), .Z(n21618) );
  XOR U26818 ( .A(round_reg[1356]), .B(n24490), .Z(n25700) );
  XNOR U26819 ( .A(n24959), .B(n25050), .Z(n24490) );
  XNOR U26820 ( .A(n25753), .B(n25754), .Z(n25050) );
  XNOR U26821 ( .A(round_reg[1291]), .B(round_reg[11]), .Z(n25754) );
  XOR U26822 ( .A(round_reg[331]), .B(n25755), .Z(n25753) );
  XOR U26823 ( .A(round_reg[971]), .B(round_reg[651]), .Z(n25755) );
  XNOR U26824 ( .A(n25756), .B(n25757), .Z(n24959) );
  XNOR U26825 ( .A(round_reg[140]), .B(round_reg[1100]), .Z(n25757) );
  XOR U26826 ( .A(round_reg[1420]), .B(n25758), .Z(n25756) );
  XOR U26827 ( .A(round_reg[780]), .B(round_reg[460]), .Z(n25758) );
  XOR U26828 ( .A(round_reg[980]), .B(n24746), .Z(n19872) );
  XOR U26829 ( .A(n24739), .B(n25125), .Z(n24746) );
  XNOR U26830 ( .A(n25759), .B(n25760), .Z(n25125) );
  XNOR U26831 ( .A(round_reg[1555]), .B(round_reg[1235]), .Z(n25760) );
  XOR U26832 ( .A(round_reg[275]), .B(n25761), .Z(n25759) );
  XOR U26833 ( .A(round_reg[915]), .B(round_reg[595]), .Z(n25761) );
  XNOR U26834 ( .A(n25762), .B(n25763), .Z(n24739) );
  XNOR U26835 ( .A(round_reg[1364]), .B(round_reg[1044]), .Z(n25763) );
  XOR U26836 ( .A(round_reg[404]), .B(n25764), .Z(n25762) );
  XOR U26837 ( .A(round_reg[84]), .B(round_reg[724]), .Z(n25764) );
  XNOR U26838 ( .A(round_reg[933]), .B(n25042), .Z(n19874) );
  NOR U26839 ( .A(n13306), .B(n13308), .Z(n25664) );
  XNOR U26840 ( .A(n22001), .B(n17564), .Z(n13308) );
  XOR U26841 ( .A(n22636), .B(n22700), .Z(n17564) );
  XOR U26842 ( .A(n25765), .B(n25766), .Z(n22700) );
  XNOR U26843 ( .A(n17924), .B(n18523), .Z(n25766) );
  XOR U26844 ( .A(n25767), .B(n22403), .Z(n18523) );
  XOR U26845 ( .A(round_reg[423]), .B(n24450), .Z(n22403) );
  XNOR U26846 ( .A(n25768), .B(n25143), .Z(n24450) );
  XNOR U26847 ( .A(n25769), .B(n25770), .Z(n25143) );
  XNOR U26848 ( .A(round_reg[1447]), .B(round_reg[1127]), .Z(n25770) );
  XOR U26849 ( .A(round_reg[167]), .B(n25771), .Z(n25769) );
  XOR U26850 ( .A(round_reg[807]), .B(round_reg[487]), .Z(n25771) );
  AND U26851 ( .A(n21821), .B(n24855), .Z(n25767) );
  IV U26852 ( .A(n21822), .Z(n24855) );
  XOR U26853 ( .A(round_reg[1596]), .B(n25177), .Z(n21822) );
  XOR U26854 ( .A(n24821), .B(n25772), .Z(n25177) );
  XOR U26855 ( .A(n25773), .B(n25774), .Z(n24821) );
  XNOR U26856 ( .A(round_reg[1340]), .B(round_reg[1020]), .Z(n25774) );
  XOR U26857 ( .A(round_reg[380]), .B(n25775), .Z(n25773) );
  XOR U26858 ( .A(round_reg[700]), .B(round_reg[60]), .Z(n25775) );
  XOR U26859 ( .A(round_reg[46]), .B(n24828), .Z(n21821) );
  XNOR U26860 ( .A(n25776), .B(n22394), .Z(n17924) );
  XNOR U26861 ( .A(round_reg[372]), .B(n22796), .Z(n22394) );
  AND U26862 ( .A(n21813), .B(n21811), .Z(n25776) );
  XOR U26863 ( .A(round_reg[298]), .B(n23602), .Z(n21811) );
  IV U26864 ( .A(n24738), .Z(n23602) );
  XNOR U26865 ( .A(n25222), .B(n25777), .Z(n24738) );
  XOR U26866 ( .A(n25778), .B(n25779), .Z(n25222) );
  XNOR U26867 ( .A(round_reg[1322]), .B(round_reg[1002]), .Z(n25779) );
  XOR U26868 ( .A(round_reg[362]), .B(n25780), .Z(n25778) );
  XOR U26869 ( .A(round_reg[682]), .B(round_reg[42]), .Z(n25780) );
  XOR U26870 ( .A(round_reg[1531]), .B(n21617), .Z(n21813) );
  XOR U26871 ( .A(n25781), .B(n25782), .Z(n25354) );
  XNOR U26872 ( .A(round_reg[1595]), .B(round_reg[1275]), .Z(n25782) );
  XOR U26873 ( .A(round_reg[315]), .B(n25783), .Z(n25781) );
  XOR U26874 ( .A(round_reg[955]), .B(round_reg[635]), .Z(n25783) );
  XNOR U26875 ( .A(n25784), .B(n25785), .Z(n25378) );
  XNOR U26876 ( .A(round_reg[1466]), .B(round_reg[1146]), .Z(n25785) );
  XOR U26877 ( .A(round_reg[186]), .B(n25786), .Z(n25784) );
  XOR U26878 ( .A(round_reg[826]), .B(round_reg[506]), .Z(n25786) );
  XOR U26879 ( .A(n19958), .B(n25787), .Z(n25765) );
  XOR U26880 ( .A(n22388), .B(n20023), .Z(n25787) );
  XNOR U26881 ( .A(n25788), .B(n23213), .Z(n20023) );
  XOR U26882 ( .A(round_reg[595]), .B(n24202), .Z(n23213) );
  AND U26883 ( .A(n21817), .B(n21819), .Z(n25788) );
  XNOR U26884 ( .A(round_reg[1470]), .B(n22435), .Z(n21819) );
  XNOR U26885 ( .A(n25285), .B(n25789), .Z(n22435) );
  XOR U26886 ( .A(n25790), .B(n25791), .Z(n25285) );
  XNOR U26887 ( .A(round_reg[125]), .B(round_reg[1085]), .Z(n25791) );
  XOR U26888 ( .A(round_reg[1405]), .B(n25792), .Z(n25790) );
  XOR U26889 ( .A(round_reg[765]), .B(round_reg[445]), .Z(n25792) );
  XOR U26890 ( .A(n25793), .B(n25145), .Z(n23249) );
  XOR U26891 ( .A(n25794), .B(n25795), .Z(n25145) );
  XNOR U26892 ( .A(round_reg[1465]), .B(round_reg[1145]), .Z(n25795) );
  XOR U26893 ( .A(round_reg[185]), .B(n25796), .Z(n25794) );
  XOR U26894 ( .A(round_reg[825]), .B(round_reg[505]), .Z(n25796) );
  XNOR U26895 ( .A(n25797), .B(n24660), .Z(n22388) );
  XOR U26896 ( .A(round_reg[493]), .B(n23413), .Z(n24660) );
  IV U26897 ( .A(n24013), .Z(n23413) );
  XOR U26898 ( .A(n25072), .B(n24735), .Z(n24013) );
  XOR U26899 ( .A(n25798), .B(n25799), .Z(n24735) );
  XNOR U26900 ( .A(round_reg[108]), .B(round_reg[1068]), .Z(n25799) );
  XOR U26901 ( .A(round_reg[1388]), .B(n25800), .Z(n25798) );
  XOR U26902 ( .A(round_reg[748]), .B(round_reg[428]), .Z(n25800) );
  XOR U26903 ( .A(n25801), .B(n25802), .Z(n25072) );
  XNOR U26904 ( .A(round_reg[1517]), .B(round_reg[1197]), .Z(n25802) );
  XOR U26905 ( .A(round_reg[237]), .B(n25803), .Z(n25801) );
  XOR U26906 ( .A(round_reg[877]), .B(round_reg[557]), .Z(n25803) );
  AND U26907 ( .A(n21807), .B(n24858), .Z(n25797) );
  IV U26908 ( .A(n21808), .Z(n24858) );
  XOR U26909 ( .A(round_reg[1313]), .B(n23144), .Z(n21808) );
  IV U26910 ( .A(n24815), .Z(n23144) );
  XOR U26911 ( .A(round_reg[68]), .B(n23721), .Z(n21807) );
  XNOR U26912 ( .A(n25680), .B(n24396), .Z(n23721) );
  XNOR U26913 ( .A(n25804), .B(n25805), .Z(n24396) );
  XNOR U26914 ( .A(round_reg[132]), .B(round_reg[1092]), .Z(n25805) );
  XOR U26915 ( .A(round_reg[1412]), .B(n25806), .Z(n25804) );
  XOR U26916 ( .A(round_reg[772]), .B(round_reg[452]), .Z(n25806) );
  XNOR U26917 ( .A(n25807), .B(n25808), .Z(n25680) );
  XNOR U26918 ( .A(round_reg[323]), .B(round_reg[1283]), .Z(n25808) );
  XOR U26919 ( .A(round_reg[3]), .B(n25809), .Z(n25807) );
  XOR U26920 ( .A(round_reg[963]), .B(round_reg[643]), .Z(n25809) );
  XNOR U26921 ( .A(n25810), .B(n22399), .Z(n19958) );
  XOR U26922 ( .A(round_reg[527]), .B(n23793), .Z(n22399) );
  XOR U26923 ( .A(n25811), .B(n25676), .Z(n23793) );
  XNOR U26924 ( .A(n25812), .B(n25813), .Z(n25676) );
  XNOR U26925 ( .A(round_reg[1422]), .B(round_reg[1102]), .Z(n25813) );
  XOR U26926 ( .A(round_reg[142]), .B(n25814), .Z(n25812) );
  XOR U26927 ( .A(round_reg[782]), .B(round_reg[462]), .Z(n25814) );
  ANDN U26928 ( .B(n22400), .A(n22704), .Z(n25810) );
  XOR U26929 ( .A(round_reg[1376]), .B(n22268), .Z(n22704) );
  XNOR U26930 ( .A(n25815), .B(n25816), .Z(n25206) );
  XNOR U26931 ( .A(round_reg[1440]), .B(round_reg[1120]), .Z(n25816) );
  XOR U26932 ( .A(round_reg[160]), .B(n25817), .Z(n25815) );
  XOR U26933 ( .A(round_reg[800]), .B(round_reg[480]), .Z(n25817) );
  XOR U26934 ( .A(round_reg[191]), .B(n23603), .Z(n22400) );
  XNOR U26935 ( .A(n25268), .B(n25317), .Z(n23603) );
  XOR U26936 ( .A(n25819), .B(n25820), .Z(n25317) );
  XNOR U26937 ( .A(round_reg[1535]), .B(round_reg[1215]), .Z(n25820) );
  XOR U26938 ( .A(round_reg[255]), .B(n25821), .Z(n25819) );
  XOR U26939 ( .A(round_reg[895]), .B(round_reg[575]), .Z(n25821) );
  XOR U26940 ( .A(n25822), .B(n25823), .Z(n25268) );
  XNOR U26941 ( .A(round_reg[126]), .B(round_reg[1086]), .Z(n25823) );
  XOR U26942 ( .A(round_reg[1406]), .B(n25824), .Z(n25822) );
  XOR U26943 ( .A(round_reg[766]), .B(round_reg[446]), .Z(n25824) );
  XOR U26944 ( .A(n25825), .B(n25826), .Z(n22636) );
  XOR U26945 ( .A(n16982), .B(n16923), .Z(n25826) );
  XNOR U26946 ( .A(n25827), .B(n20825), .Z(n16923) );
  XNOR U26947 ( .A(round_reg[1001]), .B(n24221), .Z(n20825) );
  XNOR U26948 ( .A(n25828), .B(n25829), .Z(n25718) );
  XNOR U26949 ( .A(round_reg[1065]), .B(round_reg[105]), .Z(n25829) );
  XOR U26950 ( .A(round_reg[1385]), .B(n25830), .Z(n25828) );
  XOR U26951 ( .A(round_reg[745]), .B(round_reg[425]), .Z(n25830) );
  XNOR U26952 ( .A(n25831), .B(n25832), .Z(n25144) );
  XNOR U26953 ( .A(round_reg[1576]), .B(round_reg[1256]), .Z(n25832) );
  XOR U26954 ( .A(round_reg[296]), .B(n25833), .Z(n25831) );
  XOR U26955 ( .A(round_reg[936]), .B(round_reg[616]), .Z(n25833) );
  ANDN U26956 ( .B(n21264), .A(n22005), .Z(n25827) );
  XOR U26957 ( .A(round_reg[528]), .B(n24229), .Z(n22005) );
  XOR U26958 ( .A(n25259), .B(n25465), .Z(n24229) );
  XNOR U26959 ( .A(n25834), .B(n25835), .Z(n25465) );
  XNOR U26960 ( .A(round_reg[1552]), .B(round_reg[1232]), .Z(n25835) );
  XOR U26961 ( .A(round_reg[272]), .B(n25836), .Z(n25834) );
  XOR U26962 ( .A(round_reg[912]), .B(round_reg[592]), .Z(n25836) );
  XOR U26963 ( .A(n25837), .B(n25838), .Z(n25259) );
  XNOR U26964 ( .A(round_reg[1423]), .B(round_reg[1103]), .Z(n25838) );
  XOR U26965 ( .A(round_reg[143]), .B(n25839), .Z(n25837) );
  XOR U26966 ( .A(round_reg[783]), .B(round_reg[463]), .Z(n25839) );
  XOR U26967 ( .A(round_reg[954]), .B(n23318), .Z(n21264) );
  XNOR U26968 ( .A(n25840), .B(n25841), .Z(n25442) );
  XNOR U26969 ( .A(round_reg[1338]), .B(round_reg[1018]), .Z(n25841) );
  XOR U26970 ( .A(round_reg[378]), .B(n25842), .Z(n25840) );
  XOR U26971 ( .A(round_reg[698]), .B(round_reg[58]), .Z(n25842) );
  XNOR U26972 ( .A(n25844), .B(n20822), .Z(n16982) );
  XOR U26973 ( .A(round_reg[1169]), .B(n23885), .Z(n20822) );
  XOR U26974 ( .A(n25522), .B(n25166), .Z(n23885) );
  XNOR U26975 ( .A(n25845), .B(n25846), .Z(n25166) );
  XNOR U26976 ( .A(round_reg[1424]), .B(round_reg[1104]), .Z(n25846) );
  XOR U26977 ( .A(round_reg[144]), .B(n25847), .Z(n25845) );
  XOR U26978 ( .A(round_reg[784]), .B(round_reg[464]), .Z(n25847) );
  XOR U26979 ( .A(n25848), .B(n25849), .Z(n25522) );
  XNOR U26980 ( .A(round_reg[1553]), .B(round_reg[1233]), .Z(n25849) );
  XOR U26981 ( .A(round_reg[273]), .B(n25850), .Z(n25848) );
  XOR U26982 ( .A(round_reg[913]), .B(round_reg[593]), .Z(n25850) );
  AND U26983 ( .A(n22003), .B(n21271), .Z(n25844) );
  XOR U26984 ( .A(round_reg[786]), .B(n23295), .Z(n21271) );
  XNOR U26985 ( .A(n25851), .B(n25852), .Z(n25466) );
  XNOR U26986 ( .A(round_reg[1361]), .B(round_reg[1041]), .Z(n25852) );
  XOR U26987 ( .A(round_reg[401]), .B(n25853), .Z(n25851) );
  XOR U26988 ( .A(round_reg[81]), .B(round_reg[721]), .Z(n25853) );
  XNOR U26989 ( .A(round_reg[424]), .B(n25364), .Z(n22003) );
  XNOR U26990 ( .A(n21258), .B(n25855), .Z(n25825) );
  XOR U26991 ( .A(n18448), .B(n17490), .Z(n25855) );
  XNOR U26992 ( .A(n25856), .B(n21268), .Z(n17490) );
  XOR U26993 ( .A(round_reg[1241]), .B(n23918), .Z(n21268) );
  IV U26994 ( .A(n21310), .Z(n23918) );
  XOR U26995 ( .A(n25682), .B(n25620), .Z(n21310) );
  XOR U26996 ( .A(n25857), .B(n25858), .Z(n25620) );
  XNOR U26997 ( .A(round_reg[25]), .B(round_reg[1305]), .Z(n25858) );
  XOR U26998 ( .A(round_reg[345]), .B(n25859), .Z(n25857) );
  XOR U26999 ( .A(round_reg[985]), .B(round_reg[665]), .Z(n25859) );
  XOR U27000 ( .A(n25860), .B(n25861), .Z(n25682) );
  XNOR U27001 ( .A(round_reg[1496]), .B(round_reg[1176]), .Z(n25861) );
  XOR U27002 ( .A(round_reg[216]), .B(n25862), .Z(n25860) );
  XOR U27003 ( .A(round_reg[856]), .B(round_reg[536]), .Z(n25862) );
  ANDN U27004 ( .B(n24847), .A(n21267), .Z(n25856) );
  XNOR U27005 ( .A(n25863), .B(n21274), .Z(n18448) );
  XOR U27006 ( .A(round_reg[1030]), .B(n23883), .Z(n21274) );
  AND U27007 ( .A(n21275), .B(n24845), .Z(n25863) );
  IV U27008 ( .A(n21996), .Z(n24845) );
  XOR U27009 ( .A(round_reg[596]), .B(n24137), .Z(n21996) );
  IV U27010 ( .A(n22818), .Z(n24137) );
  XOR U27011 ( .A(n25020), .B(n25235), .Z(n22818) );
  XOR U27012 ( .A(n25864), .B(n25865), .Z(n25235) );
  XNOR U27013 ( .A(round_reg[1491]), .B(round_reg[1171]), .Z(n25865) );
  XOR U27014 ( .A(round_reg[211]), .B(n25866), .Z(n25864) );
  XOR U27015 ( .A(round_reg[851]), .B(round_reg[531]), .Z(n25866) );
  XOR U27016 ( .A(n25867), .B(n25868), .Z(n25020) );
  XNOR U27017 ( .A(round_reg[20]), .B(round_reg[1300]), .Z(n25868) );
  XOR U27018 ( .A(round_reg[340]), .B(n25869), .Z(n25867) );
  XOR U27019 ( .A(round_reg[980]), .B(round_reg[660]), .Z(n25869) );
  XOR U27020 ( .A(round_reg[662]), .B(n23596), .Z(n21275) );
  XNOR U27021 ( .A(n25870), .B(n20815), .Z(n21258) );
  XNOR U27022 ( .A(round_reg[1143]), .B(n24029), .Z(n20815) );
  XOR U27023 ( .A(n25372), .B(n25871), .Z(n24029) );
  XOR U27024 ( .A(n25872), .B(n25873), .Z(n25372) );
  XNOR U27025 ( .A(round_reg[118]), .B(round_reg[1078]), .Z(n25873) );
  XOR U27026 ( .A(round_reg[1398]), .B(n25874), .Z(n25872) );
  XOR U27027 ( .A(round_reg[758]), .B(round_reg[438]), .Z(n25874) );
  NOR U27028 ( .A(n21999), .B(n21277), .Z(n25870) );
  XNOR U27029 ( .A(round_reg[740]), .B(n22272), .Z(n21277) );
  XNOR U27030 ( .A(n25875), .B(n25876), .Z(n25195) );
  XNOR U27031 ( .A(round_reg[355]), .B(round_reg[1315]), .Z(n25876) );
  XOR U27032 ( .A(round_reg[35]), .B(n25877), .Z(n25875) );
  XOR U27033 ( .A(round_reg[995]), .B(round_reg[675]), .Z(n25877) );
  XNOR U27034 ( .A(n25878), .B(n25879), .Z(n25087) );
  XNOR U27035 ( .A(round_reg[1444]), .B(round_reg[1124]), .Z(n25879) );
  XOR U27036 ( .A(round_reg[164]), .B(n25880), .Z(n25878) );
  XOR U27037 ( .A(round_reg[804]), .B(round_reg[484]), .Z(n25880) );
  XNOR U27038 ( .A(round_reg[373]), .B(n21313), .Z(n21999) );
  XOR U27039 ( .A(n25881), .B(n21267), .Z(n22001) );
  XNOR U27040 ( .A(round_reg[883]), .B(n24518), .Z(n21267) );
  NOR U27041 ( .A(n23891), .B(n24847), .Z(n25881) );
  XNOR U27042 ( .A(round_reg[494]), .B(n23908), .Z(n24847) );
  XOR U27043 ( .A(n24664), .B(n25882), .Z(n23908) );
  XOR U27044 ( .A(n25883), .B(n25884), .Z(n24664) );
  XNOR U27045 ( .A(round_reg[109]), .B(round_reg[1069]), .Z(n25884) );
  XOR U27046 ( .A(round_reg[1389]), .B(n25885), .Z(n25883) );
  XOR U27047 ( .A(round_reg[749]), .B(round_reg[429]), .Z(n25885) );
  XOR U27048 ( .A(round_reg[69]), .B(n24559), .Z(n23891) );
  XNOR U27049 ( .A(n22467), .B(n18789), .Z(n13306) );
  XOR U27050 ( .A(n25886), .B(n25887), .Z(n23183) );
  XNOR U27051 ( .A(n19264), .B(n21930), .Z(n25887) );
  XOR U27052 ( .A(n25888), .B(n22553), .Z(n21930) );
  XNOR U27053 ( .A(round_reg[790]), .B(n24378), .Z(n22553) );
  XNOR U27054 ( .A(n25193), .B(n24554), .Z(n24378) );
  XNOR U27055 ( .A(n25889), .B(n25890), .Z(n24554) );
  XNOR U27056 ( .A(round_reg[1494]), .B(round_reg[1174]), .Z(n25890) );
  XOR U27057 ( .A(round_reg[214]), .B(n25891), .Z(n25889) );
  XOR U27058 ( .A(round_reg[854]), .B(round_reg[534]), .Z(n25891) );
  XNOR U27059 ( .A(n25892), .B(n25893), .Z(n25193) );
  XNOR U27060 ( .A(round_reg[1365]), .B(round_reg[1045]), .Z(n25893) );
  XOR U27061 ( .A(round_reg[405]), .B(n25894), .Z(n25892) );
  XOR U27062 ( .A(round_reg[85]), .B(round_reg[725]), .Z(n25894) );
  AND U27063 ( .A(n23633), .B(n24428), .Z(n25888) );
  XOR U27064 ( .A(round_reg[51]), .B(n24545), .Z(n24428) );
  IV U27065 ( .A(n23504), .Z(n24545) );
  XOR U27066 ( .A(n25474), .B(n25895), .Z(n23504) );
  XOR U27067 ( .A(n25896), .B(n25897), .Z(n25474) );
  XNOR U27068 ( .A(round_reg[1586]), .B(round_reg[1266]), .Z(n25897) );
  XOR U27069 ( .A(round_reg[306]), .B(n25898), .Z(n25896) );
  XOR U27070 ( .A(round_reg[946]), .B(round_reg[626]), .Z(n25898) );
  XOR U27071 ( .A(round_reg[428]), .B(n24364), .Z(n23633) );
  IV U27072 ( .A(n23940), .Z(n24364) );
  XOR U27073 ( .A(n24841), .B(n25899), .Z(n23940) );
  XOR U27074 ( .A(n25900), .B(n25901), .Z(n24841) );
  XNOR U27075 ( .A(round_reg[1323]), .B(round_reg[1003]), .Z(n25901) );
  XOR U27076 ( .A(round_reg[363]), .B(n25902), .Z(n25900) );
  XOR U27077 ( .A(round_reg[683]), .B(round_reg[43]), .Z(n25902) );
  XNOR U27078 ( .A(n25903), .B(n22566), .Z(n19264) );
  XOR U27079 ( .A(round_reg[744]), .B(n25364), .Z(n22566) );
  AND U27080 ( .A(n23640), .B(n24177), .Z(n25903) );
  XOR U27081 ( .A(round_reg[303]), .B(n24207), .Z(n24177) );
  IV U27082 ( .A(n21763), .Z(n24207) );
  XNOR U27083 ( .A(n25905), .B(n25906), .Z(n25882) );
  XNOR U27084 ( .A(round_reg[1518]), .B(round_reg[1198]), .Z(n25906) );
  XOR U27085 ( .A(round_reg[238]), .B(n25907), .Z(n25905) );
  XOR U27086 ( .A(round_reg[878]), .B(round_reg[558]), .Z(n25907) );
  XOR U27087 ( .A(round_reg[377]), .B(n23469), .Z(n23640) );
  XOR U27088 ( .A(n25908), .B(n25909), .Z(n23469) );
  XOR U27089 ( .A(n22237), .B(n25910), .Z(n25886) );
  XNOR U27090 ( .A(n19218), .B(n21215), .Z(n25910) );
  XOR U27091 ( .A(n25911), .B(n22547), .Z(n21215) );
  XNOR U27092 ( .A(round_reg[958]), .B(n23877), .Z(n22547) );
  XNOR U27093 ( .A(n25335), .B(n25653), .Z(n23877) );
  XNOR U27094 ( .A(n25912), .B(n25913), .Z(n25653) );
  XNOR U27095 ( .A(round_reg[1342]), .B(round_reg[1022]), .Z(n25913) );
  XOR U27096 ( .A(round_reg[382]), .B(n25914), .Z(n25912) );
  XOR U27097 ( .A(round_reg[702]), .B(round_reg[62]), .Z(n25914) );
  XOR U27098 ( .A(n25915), .B(n25916), .Z(n25335) );
  XNOR U27099 ( .A(round_reg[1533]), .B(round_reg[1213]), .Z(n25916) );
  XOR U27100 ( .A(round_reg[253]), .B(n25917), .Z(n25915) );
  XOR U27101 ( .A(round_reg[893]), .B(round_reg[573]), .Z(n25917) );
  AND U27102 ( .A(n23631), .B(n24173), .Z(n25911) );
  XOR U27103 ( .A(round_reg[132]), .B(n25085), .Z(n24173) );
  XOR U27104 ( .A(round_reg[532]), .B(n22979), .Z(n23631) );
  XNOR U27105 ( .A(n25918), .B(n22558), .Z(n19218) );
  XOR U27106 ( .A(round_reg[887]), .B(n23127), .Z(n22558) );
  NOR U27107 ( .A(n23636), .B(n24170), .Z(n25918) );
  XNOR U27108 ( .A(round_reg[73]), .B(n24448), .Z(n24170) );
  XNOR U27109 ( .A(round_reg[498]), .B(n24692), .Z(n23636) );
  XOR U27110 ( .A(n25288), .B(n24762), .Z(n24692) );
  XNOR U27111 ( .A(n25919), .B(n25920), .Z(n24762) );
  XNOR U27112 ( .A(round_reg[113]), .B(round_reg[1073]), .Z(n25920) );
  XOR U27113 ( .A(round_reg[1393]), .B(n25921), .Z(n25919) );
  XOR U27114 ( .A(round_reg[753]), .B(round_reg[433]), .Z(n25921) );
  XOR U27115 ( .A(n25922), .B(n25923), .Z(n25288) );
  XNOR U27116 ( .A(round_reg[1522]), .B(round_reg[1202]), .Z(n25923) );
  XOR U27117 ( .A(round_reg[242]), .B(n25924), .Z(n25922) );
  XOR U27118 ( .A(round_reg[882]), .B(round_reg[562]), .Z(n25924) );
  XNOR U27119 ( .A(n25925), .B(n22562), .Z(n22237) );
  XOR U27120 ( .A(round_reg[666]), .B(n24823), .Z(n22562) );
  XOR U27121 ( .A(n25547), .B(n25302), .Z(n24823) );
  XNOR U27122 ( .A(n25926), .B(n25927), .Z(n25302) );
  XNOR U27123 ( .A(round_reg[1561]), .B(round_reg[1241]), .Z(n25927) );
  XOR U27124 ( .A(round_reg[281]), .B(n25928), .Z(n25926) );
  XOR U27125 ( .A(round_reg[921]), .B(round_reg[601]), .Z(n25928) );
  XOR U27126 ( .A(n25929), .B(n25930), .Z(n25547) );
  XNOR U27127 ( .A(round_reg[1370]), .B(round_reg[1050]), .Z(n25930) );
  XOR U27128 ( .A(round_reg[410]), .B(n25931), .Z(n25929) );
  XOR U27129 ( .A(round_reg[90]), .B(round_reg[730]), .Z(n25931) );
  AND U27130 ( .A(n23638), .B(n24179), .Z(n25925) );
  XNOR U27131 ( .A(round_reg[255]), .B(n23904), .Z(n24179) );
  XOR U27132 ( .A(n25933), .B(n25934), .Z(n25580) );
  XNOR U27133 ( .A(round_reg[1470]), .B(round_reg[1150]), .Z(n25934) );
  XOR U27134 ( .A(round_reg[190]), .B(n25935), .Z(n25933) );
  XOR U27135 ( .A(round_reg[830]), .B(round_reg[510]), .Z(n25935) );
  XOR U27136 ( .A(round_reg[600]), .B(n23406), .Z(n23638) );
  XOR U27137 ( .A(n24816), .B(n25936), .Z(n23406) );
  XOR U27138 ( .A(n25937), .B(n25938), .Z(n24816) );
  XNOR U27139 ( .A(round_reg[24]), .B(round_reg[1304]), .Z(n25938) );
  XOR U27140 ( .A(round_reg[344]), .B(n25939), .Z(n25937) );
  XOR U27141 ( .A(round_reg[984]), .B(round_reg[664]), .Z(n25939) );
  XOR U27142 ( .A(n25940), .B(n25941), .Z(n24890) );
  XOR U27143 ( .A(n18542), .B(n15965), .Z(n25941) );
  XOR U27144 ( .A(n25942), .B(n22581), .Z(n15965) );
  XOR U27145 ( .A(round_reg[1382]), .B(n23865), .Z(n22581) );
  ANDN U27146 ( .B(n22460), .A(n22461), .Z(n25942) );
  XOR U27147 ( .A(round_reg[959]), .B(n21603), .Z(n22461) );
  IV U27148 ( .A(n24299), .Z(n21603) );
  XOR U27149 ( .A(n25789), .B(n25943), .Z(n24299) );
  XOR U27150 ( .A(n25944), .B(n25945), .Z(n25789) );
  XNOR U27151 ( .A(round_reg[1534]), .B(round_reg[1214]), .Z(n25945) );
  XOR U27152 ( .A(round_reg[254]), .B(n25946), .Z(n25944) );
  XOR U27153 ( .A(round_reg[894]), .B(round_reg[574]), .Z(n25946) );
  XOR U27154 ( .A(round_reg[1006]), .B(n24828), .Z(n22460) );
  XNOR U27155 ( .A(n25947), .B(n22578), .Z(n18542) );
  XOR U27156 ( .A(round_reg[1538]), .B(n23252), .Z(n22578) );
  IV U27157 ( .A(n23930), .Z(n23252) );
  XNOR U27158 ( .A(n25948), .B(n24336), .Z(n23930) );
  XNOR U27159 ( .A(n25949), .B(n25950), .Z(n24336) );
  XNOR U27160 ( .A(round_reg[1473]), .B(round_reg[1153]), .Z(n25950) );
  XOR U27161 ( .A(round_reg[193]), .B(n25951), .Z(n25949) );
  XOR U27162 ( .A(round_reg[833]), .B(round_reg[513]), .Z(n25951) );
  XOR U27163 ( .A(round_reg[791]), .B(n23254), .Z(n22465) );
  XNOR U27164 ( .A(n25952), .B(n25936), .Z(n23254) );
  XNOR U27165 ( .A(n25953), .B(n25954), .Z(n25936) );
  XNOR U27166 ( .A(round_reg[1495]), .B(round_reg[1175]), .Z(n25954) );
  XOR U27167 ( .A(round_reg[215]), .B(n25955), .Z(n25953) );
  XOR U27168 ( .A(round_reg[855]), .B(round_reg[535]), .Z(n25955) );
  XOR U27169 ( .A(round_reg[1174]), .B(n24904), .Z(n22464) );
  IV U27170 ( .A(n22691), .Z(n24904) );
  XNOR U27171 ( .A(n25461), .B(n25021), .Z(n22691) );
  XNOR U27172 ( .A(n25956), .B(n25957), .Z(n25021) );
  XNOR U27173 ( .A(round_reg[1429]), .B(round_reg[1109]), .Z(n25957) );
  XOR U27174 ( .A(round_reg[149]), .B(n25958), .Z(n25956) );
  XOR U27175 ( .A(round_reg[789]), .B(round_reg[469]), .Z(n25958) );
  XNOR U27176 ( .A(n25959), .B(n25960), .Z(n25461) );
  XNOR U27177 ( .A(round_reg[1558]), .B(round_reg[1238]), .Z(n25960) );
  XOR U27178 ( .A(round_reg[278]), .B(n25961), .Z(n25959) );
  XOR U27179 ( .A(round_reg[918]), .B(round_reg[598]), .Z(n25961) );
  XOR U27180 ( .A(n23626), .B(n25962), .Z(n25940) );
  XOR U27181 ( .A(n17875), .B(n15532), .Z(n25962) );
  XNOR U27182 ( .A(n25963), .B(n22572), .Z(n15532) );
  XOR U27183 ( .A(round_reg[1319]), .B(n23799), .Z(n22572) );
  XOR U27184 ( .A(n25714), .B(n25660), .Z(n23799) );
  XNOR U27185 ( .A(n25964), .B(n25965), .Z(n25660) );
  XNOR U27186 ( .A(round_reg[1063]), .B(round_reg[103]), .Z(n25965) );
  XOR U27187 ( .A(round_reg[1383]), .B(n25966), .Z(n25964) );
  XOR U27188 ( .A(round_reg[743]), .B(round_reg[423]), .Z(n25966) );
  XOR U27189 ( .A(n25967), .B(n25968), .Z(n25714) );
  XNOR U27190 ( .A(round_reg[1574]), .B(round_reg[1254]), .Z(n25968) );
  XOR U27191 ( .A(round_reg[294]), .B(n25969), .Z(n25967) );
  XOR U27192 ( .A(round_reg[934]), .B(round_reg[614]), .Z(n25969) );
  ANDN U27193 ( .B(n22470), .A(n22471), .Z(n25963) );
  XOR U27194 ( .A(round_reg[888]), .B(n23777), .Z(n22471) );
  XNOR U27195 ( .A(n25970), .B(n25971), .Z(n25092) );
  XNOR U27196 ( .A(round_reg[1463]), .B(round_reg[1143]), .Z(n25971) );
  XOR U27197 ( .A(round_reg[183]), .B(n25972), .Z(n25970) );
  XOR U27198 ( .A(round_reg[823]), .B(round_reg[503]), .Z(n25972) );
  XNOR U27199 ( .A(n25973), .B(n25974), .Z(n25909) );
  XNOR U27200 ( .A(round_reg[1592]), .B(round_reg[1272]), .Z(n25974) );
  XOR U27201 ( .A(round_reg[312]), .B(n25975), .Z(n25973) );
  XOR U27202 ( .A(round_reg[952]), .B(round_reg[632]), .Z(n25975) );
  XNOR U27203 ( .A(round_reg[1246]), .B(n25008), .Z(n22470) );
  IV U27204 ( .A(n23464), .Z(n25008) );
  XOR U27205 ( .A(n25977), .B(n25978), .Z(n24970) );
  XNOR U27206 ( .A(round_reg[30]), .B(round_reg[1310]), .Z(n25978) );
  XOR U27207 ( .A(round_reg[350]), .B(n25979), .Z(n25977) );
  XOR U27208 ( .A(round_reg[990]), .B(round_reg[670]), .Z(n25979) );
  XNOR U27209 ( .A(n25980), .B(n22809), .Z(n17875) );
  XOR U27210 ( .A(round_reg[1412]), .B(n24728), .Z(n22809) );
  IV U27211 ( .A(n25085), .Z(n24728) );
  XOR U27212 ( .A(n25981), .B(n25014), .Z(n25085) );
  XOR U27213 ( .A(n25982), .B(n25983), .Z(n25014) );
  XNOR U27214 ( .A(round_reg[1347]), .B(round_reg[1027]), .Z(n25983) );
  XOR U27215 ( .A(round_reg[387]), .B(n25984), .Z(n25982) );
  XOR U27216 ( .A(round_reg[707]), .B(round_reg[67]), .Z(n25984) );
  XOR U27217 ( .A(round_reg[667]), .B(n23386), .Z(n22475) );
  XOR U27218 ( .A(n25253), .B(n25229), .Z(n23386) );
  XOR U27219 ( .A(n25985), .B(n25986), .Z(n25229) );
  XNOR U27220 ( .A(round_reg[1371]), .B(round_reg[1051]), .Z(n25986) );
  XOR U27221 ( .A(round_reg[411]), .B(n25987), .Z(n25985) );
  XOR U27222 ( .A(round_reg[91]), .B(round_reg[731]), .Z(n25987) );
  XNOR U27223 ( .A(n25988), .B(n25989), .Z(n25253) );
  XNOR U27224 ( .A(round_reg[1562]), .B(round_reg[1242]), .Z(n25989) );
  XOR U27225 ( .A(round_reg[282]), .B(n25990), .Z(n25988) );
  XOR U27226 ( .A(round_reg[922]), .B(round_reg[602]), .Z(n25990) );
  XOR U27227 ( .A(round_reg[1035]), .B(n24906), .Z(n22474) );
  XNOR U27228 ( .A(n25991), .B(n25992), .Z(n25031) );
  XNOR U27229 ( .A(round_reg[139]), .B(round_reg[1099]), .Z(n25992) );
  XOR U27230 ( .A(round_reg[1419]), .B(n25993), .Z(n25991) );
  XOR U27231 ( .A(round_reg[779]), .B(round_reg[459]), .Z(n25993) );
  XOR U27232 ( .A(n25994), .B(n25995), .Z(n25409) );
  XNOR U27233 ( .A(round_reg[1290]), .B(round_reg[10]), .Z(n25995) );
  XOR U27234 ( .A(round_reg[330]), .B(n25996), .Z(n25994) );
  XOR U27235 ( .A(round_reg[970]), .B(round_reg[650]), .Z(n25996) );
  XNOR U27236 ( .A(n25997), .B(n24193), .Z(n23626) );
  XOR U27237 ( .A(round_reg[1473]), .B(n21192), .Z(n24193) );
  IV U27238 ( .A(n22211), .Z(n21192) );
  XOR U27239 ( .A(n25999), .B(n26000), .Z(n24881) );
  XNOR U27240 ( .A(round_reg[1537]), .B(round_reg[1217]), .Z(n26000) );
  XOR U27241 ( .A(round_reg[257]), .B(n26001), .Z(n25999) );
  XOR U27242 ( .A(round_reg[897]), .B(round_reg[577]), .Z(n26001) );
  ANDN U27243 ( .B(n26002), .A(n24185), .Z(n25997) );
  XNOR U27244 ( .A(n26003), .B(n24593), .Z(n22467) );
  IV U27245 ( .A(n26002), .Z(n24593) );
  XOR U27246 ( .A(round_reg[1148]), .B(n23323), .Z(n26002) );
  XNOR U27247 ( .A(n26004), .B(n26005), .Z(n25566) );
  XNOR U27248 ( .A(round_reg[1532]), .B(round_reg[1212]), .Z(n26005) );
  XOR U27249 ( .A(round_reg[252]), .B(n26006), .Z(n26004) );
  XOR U27250 ( .A(round_reg[892]), .B(round_reg[572]), .Z(n26006) );
  ANDN U27251 ( .B(n24185), .A(n24186), .Z(n26003) );
  XOR U27252 ( .A(round_reg[378]), .B(n24578), .Z(n24186) );
  XOR U27253 ( .A(n26008), .B(n25327), .Z(n24578) );
  XNOR U27254 ( .A(n26009), .B(n26010), .Z(n25327) );
  XNOR U27255 ( .A(round_reg[1593]), .B(round_reg[1273]), .Z(n26010) );
  XOR U27256 ( .A(round_reg[313]), .B(n26011), .Z(n26009) );
  XOR U27257 ( .A(round_reg[953]), .B(round_reg[633]), .Z(n26011) );
  XOR U27258 ( .A(round_reg[745]), .B(n23876), .Z(n24185) );
  IV U27259 ( .A(n23750), .Z(n23876) );
  XNOR U27260 ( .A(n24572), .B(n25708), .Z(n23750) );
  XNOR U27261 ( .A(n26012), .B(n26013), .Z(n25708) );
  XNOR U27262 ( .A(round_reg[1320]), .B(round_reg[1000]), .Z(n26013) );
  XOR U27263 ( .A(round_reg[360]), .B(n26014), .Z(n26012) );
  XOR U27264 ( .A(round_reg[680]), .B(round_reg[40]), .Z(n26014) );
  XOR U27265 ( .A(n26015), .B(n26016), .Z(n24572) );
  XNOR U27266 ( .A(round_reg[1449]), .B(round_reg[1129]), .Z(n26016) );
  XOR U27267 ( .A(round_reg[169]), .B(n26017), .Z(n26015) );
  XOR U27268 ( .A(round_reg[809]), .B(round_reg[489]), .Z(n26017) );
  XOR U27269 ( .A(n26018), .B(n14671), .Z(n11180) );
  XOR U27270 ( .A(n16706), .B(n24610), .Z(n14671) );
  XOR U27271 ( .A(n26019), .B(n22501), .Z(n24610) );
  AND U27272 ( .A(n24629), .B(n24630), .Z(n26019) );
  XNOR U27273 ( .A(round_reg[996]), .B(n23201), .Z(n24630) );
  XNOR U27274 ( .A(n25208), .B(n25182), .Z(n23201) );
  XOR U27275 ( .A(n26020), .B(n26021), .Z(n25182) );
  XNOR U27276 ( .A(round_reg[1571]), .B(round_reg[1251]), .Z(n26021) );
  XOR U27277 ( .A(round_reg[291]), .B(n26022), .Z(n26020) );
  XOR U27278 ( .A(round_reg[931]), .B(round_reg[611]), .Z(n26022) );
  XOR U27279 ( .A(n26023), .B(n26024), .Z(n25208) );
  XNOR U27280 ( .A(round_reg[1060]), .B(round_reg[100]), .Z(n26024) );
  XOR U27281 ( .A(round_reg[1380]), .B(n26025), .Z(n26023) );
  XOR U27282 ( .A(round_reg[740]), .B(round_reg[420]), .Z(n26025) );
  XOR U27283 ( .A(n22260), .B(n23331), .Z(n16706) );
  XOR U27284 ( .A(n26026), .B(n26027), .Z(n23331) );
  XOR U27285 ( .A(n20581), .B(n16528), .Z(n26027) );
  XOR U27286 ( .A(n26028), .B(n22286), .Z(n16528) );
  XOR U27287 ( .A(round_reg[1371]), .B(n24519), .Z(n22286) );
  XOR U27288 ( .A(n26029), .B(n24995), .Z(n24519) );
  XNOR U27289 ( .A(n26030), .B(n26031), .Z(n24995) );
  XNOR U27290 ( .A(round_reg[26]), .B(round_reg[1306]), .Z(n26031) );
  XOR U27291 ( .A(round_reg[346]), .B(n26032), .Z(n26030) );
  XOR U27292 ( .A(round_reg[986]), .B(round_reg[666]), .Z(n26032) );
  AND U27293 ( .A(n24627), .B(n22892), .Z(n26028) );
  XOR U27294 ( .A(round_reg[995]), .B(n23584), .Z(n22892) );
  XNOR U27295 ( .A(n26033), .B(n26034), .Z(n25201) );
  XNOR U27296 ( .A(round_reg[1570]), .B(round_reg[1250]), .Z(n26034) );
  XOR U27297 ( .A(round_reg[290]), .B(n26035), .Z(n26033) );
  XOR U27298 ( .A(round_reg[930]), .B(round_reg[610]), .Z(n26035) );
  XNOR U27299 ( .A(n26036), .B(n26037), .Z(n25440) );
  XNOR U27300 ( .A(round_reg[1379]), .B(round_reg[1059]), .Z(n26037) );
  XOR U27301 ( .A(round_reg[419]), .B(n26038), .Z(n26036) );
  XOR U27302 ( .A(round_reg[99]), .B(round_reg[739]), .Z(n26038) );
  XNOR U27303 ( .A(round_reg[948]), .B(n24084), .Z(n24627) );
  IV U27304 ( .A(n24325), .Z(n24084) );
  XOR U27305 ( .A(n25044), .B(n26039), .Z(n24325) );
  XOR U27306 ( .A(n26040), .B(n26041), .Z(n25044) );
  XNOR U27307 ( .A(round_reg[1332]), .B(round_reg[1012]), .Z(n26041) );
  XOR U27308 ( .A(round_reg[372]), .B(n26042), .Z(n26040) );
  XOR U27309 ( .A(round_reg[692]), .B(round_reg[52]), .Z(n26042) );
  XNOR U27310 ( .A(n26043), .B(n22296), .Z(n20581) );
  XOR U27311 ( .A(round_reg[1591]), .B(n23789), .Z(n22296) );
  ANDN U27312 ( .B(n22896), .A(n24622), .Z(n26043) );
  XOR U27313 ( .A(round_reg[780]), .B(n24389), .Z(n24622) );
  XOR U27314 ( .A(round_reg[1163]), .B(n24767), .Z(n22896) );
  XOR U27315 ( .A(n22880), .B(n26044), .Z(n26026) );
  XOR U27316 ( .A(n19502), .B(n15638), .Z(n26044) );
  XNOR U27317 ( .A(n26045), .B(n22886), .Z(n15638) );
  XOR U27318 ( .A(round_reg[1308]), .B(n23121), .Z(n22886) );
  AND U27319 ( .A(n22887), .B(n24625), .Z(n26045) );
  XNOR U27320 ( .A(round_reg[877]), .B(n24309), .Z(n24625) );
  XOR U27321 ( .A(n26049), .B(n26050), .Z(n25899) );
  XNOR U27322 ( .A(round_reg[1452]), .B(round_reg[1132]), .Z(n26050) );
  XOR U27323 ( .A(round_reg[172]), .B(n26051), .Z(n26049) );
  XOR U27324 ( .A(round_reg[812]), .B(round_reg[492]), .Z(n26051) );
  XOR U27325 ( .A(round_reg[1235]), .B(n24202), .Z(n22887) );
  XOR U27326 ( .A(n24868), .B(n25854), .Z(n24202) );
  XNOR U27327 ( .A(n26052), .B(n26053), .Z(n25854) );
  XNOR U27328 ( .A(round_reg[1490]), .B(round_reg[1170]), .Z(n26053) );
  XOR U27329 ( .A(round_reg[210]), .B(n26054), .Z(n26052) );
  XOR U27330 ( .A(round_reg[850]), .B(round_reg[530]), .Z(n26054) );
  XOR U27331 ( .A(n26055), .B(n26056), .Z(n24868) );
  XNOR U27332 ( .A(round_reg[19]), .B(round_reg[1299]), .Z(n26056) );
  XOR U27333 ( .A(round_reg[339]), .B(n26057), .Z(n26055) );
  XOR U27334 ( .A(round_reg[979]), .B(round_reg[659]), .Z(n26057) );
  XNOR U27335 ( .A(n26058), .B(n22290), .Z(n19502) );
  XOR U27336 ( .A(round_reg[1465]), .B(n24296), .Z(n22290) );
  AND U27337 ( .A(n24617), .B(n22894), .Z(n26058) );
  XOR U27338 ( .A(round_reg[1024]), .B(n24381), .Z(n22894) );
  XNOR U27339 ( .A(round_reg[656]), .B(n23915), .Z(n24617) );
  XNOR U27340 ( .A(n26059), .B(n22299), .Z(n22880) );
  XOR U27341 ( .A(round_reg[1526]), .B(n24274), .Z(n22299) );
  ANDN U27342 ( .B(n22889), .A(n24619), .Z(n26059) );
  XOR U27343 ( .A(round_reg[734]), .B(n23327), .Z(n24619) );
  XOR U27344 ( .A(n25529), .B(n25499), .Z(n23327) );
  XNOR U27345 ( .A(n26060), .B(n26061), .Z(n25499) );
  XNOR U27346 ( .A(round_reg[29]), .B(round_reg[1309]), .Z(n26061) );
  XOR U27347 ( .A(round_reg[349]), .B(n26062), .Z(n26060) );
  XOR U27348 ( .A(round_reg[989]), .B(round_reg[669]), .Z(n26062) );
  XOR U27349 ( .A(n26063), .B(n26064), .Z(n25529) );
  XNOR U27350 ( .A(round_reg[1438]), .B(round_reg[1118]), .Z(n26064) );
  XOR U27351 ( .A(round_reg[158]), .B(n26065), .Z(n26063) );
  XOR U27352 ( .A(round_reg[798]), .B(round_reg[478]), .Z(n26065) );
  XNOR U27353 ( .A(round_reg[1137]), .B(n24368), .Z(n22889) );
  IV U27354 ( .A(n24285), .Z(n24368) );
  XOR U27355 ( .A(n26067), .B(n26068), .Z(n25391) );
  XNOR U27356 ( .A(round_reg[1521]), .B(round_reg[1201]), .Z(n26068) );
  XOR U27357 ( .A(round_reg[241]), .B(n26069), .Z(n26067) );
  XOR U27358 ( .A(round_reg[881]), .B(round_reg[561]), .Z(n26069) );
  XOR U27359 ( .A(n26070), .B(n26071), .Z(n22260) );
  XOR U27360 ( .A(n20164), .B(n20072), .Z(n26071) );
  XOR U27361 ( .A(n26072), .B(n22502), .Z(n20072) );
  XOR U27362 ( .A(round_reg[523]), .B(n24767), .Z(n22502) );
  XOR U27363 ( .A(n25492), .B(n25468), .Z(n24767) );
  XNOR U27364 ( .A(n26073), .B(n26074), .Z(n25468) );
  XNOR U27365 ( .A(round_reg[138]), .B(round_reg[1098]), .Z(n26074) );
  XOR U27366 ( .A(round_reg[1418]), .B(n26075), .Z(n26073) );
  XOR U27367 ( .A(round_reg[778]), .B(round_reg[458]), .Z(n26075) );
  XOR U27368 ( .A(n26076), .B(n26077), .Z(n25492) );
  XNOR U27369 ( .A(round_reg[1547]), .B(round_reg[1227]), .Z(n26077) );
  XOR U27370 ( .A(round_reg[267]), .B(n26078), .Z(n26076) );
  XOR U27371 ( .A(round_reg[907]), .B(round_reg[587]), .Z(n26078) );
  NOR U27372 ( .A(n24629), .B(n22501), .Z(n26072) );
  XNOR U27373 ( .A(round_reg[187]), .B(n23250), .Z(n22501) );
  XOR U27374 ( .A(n26008), .B(n25772), .Z(n23250) );
  XNOR U27375 ( .A(n26079), .B(n26080), .Z(n25772) );
  XNOR U27376 ( .A(round_reg[1531]), .B(round_reg[1211]), .Z(n26080) );
  XOR U27377 ( .A(round_reg[251]), .B(n26081), .Z(n26079) );
  XOR U27378 ( .A(round_reg[891]), .B(round_reg[571]), .Z(n26081) );
  XOR U27379 ( .A(n26082), .B(n26083), .Z(n26008) );
  XNOR U27380 ( .A(round_reg[122]), .B(round_reg[1082]), .Z(n26083) );
  XOR U27381 ( .A(round_reg[1402]), .B(n26084), .Z(n26082) );
  XOR U27382 ( .A(round_reg[762]), .B(round_reg[442]), .Z(n26084) );
  XOR U27383 ( .A(round_reg[1372]), .B(n22119), .Z(n24629) );
  XOR U27384 ( .A(n26085), .B(n26086), .Z(n22119) );
  XNOR U27385 ( .A(n26087), .B(n22484), .Z(n20164) );
  XOR U27386 ( .A(round_reg[591]), .B(n22802), .Z(n22484) );
  XOR U27387 ( .A(n25165), .B(n25119), .Z(n22802) );
  XNOR U27388 ( .A(n26088), .B(n26089), .Z(n25119) );
  XNOR U27389 ( .A(round_reg[1486]), .B(round_reg[1166]), .Z(n26089) );
  XOR U27390 ( .A(round_reg[206]), .B(n26090), .Z(n26088) );
  XOR U27391 ( .A(round_reg[846]), .B(round_reg[526]), .Z(n26090) );
  XOR U27392 ( .A(n26091), .B(n26092), .Z(n25165) );
  XNOR U27393 ( .A(round_reg[15]), .B(round_reg[1295]), .Z(n26092) );
  XOR U27394 ( .A(round_reg[335]), .B(n26093), .Z(n26091) );
  XOR U27395 ( .A(round_reg[975]), .B(round_reg[655]), .Z(n26093) );
  AND U27396 ( .A(n23231), .B(n22485), .Z(n26087) );
  XOR U27397 ( .A(round_reg[246]), .B(n24274), .Z(n22485) );
  IV U27398 ( .A(n25233), .Z(n24274) );
  XNOR U27399 ( .A(n26095), .B(n26096), .Z(n25045) );
  XNOR U27400 ( .A(round_reg[1461]), .B(round_reg[1141]), .Z(n26096) );
  XOR U27401 ( .A(round_reg[181]), .B(n26097), .Z(n26095) );
  XOR U27402 ( .A(round_reg[821]), .B(round_reg[501]), .Z(n26097) );
  XNOR U27403 ( .A(round_reg[1466]), .B(n24493), .Z(n23231) );
  IV U27404 ( .A(n24451), .Z(n24493) );
  XNOR U27405 ( .A(n25908), .B(n26098), .Z(n24451) );
  XOR U27406 ( .A(n26099), .B(n26100), .Z(n25908) );
  XNOR U27407 ( .A(round_reg[121]), .B(round_reg[1081]), .Z(n26100) );
  XOR U27408 ( .A(round_reg[1401]), .B(n26101), .Z(n26099) );
  XOR U27409 ( .A(round_reg[761]), .B(round_reg[441]), .Z(n26101) );
  XOR U27410 ( .A(n22479), .B(n26102), .Z(n26070) );
  XOR U27411 ( .A(n18680), .B(n16464), .Z(n26102) );
  XNOR U27412 ( .A(n26103), .B(n22497), .Z(n16464) );
  XOR U27413 ( .A(round_reg[489]), .B(n22372), .Z(n22497) );
  XNOR U27414 ( .A(n26104), .B(n26105), .Z(n25777) );
  XNOR U27415 ( .A(round_reg[1513]), .B(round_reg[1193]), .Z(n26105) );
  XOR U27416 ( .A(round_reg[233]), .B(n26106), .Z(n26104) );
  XOR U27417 ( .A(round_reg[873]), .B(round_reg[553]), .Z(n26106) );
  XNOR U27418 ( .A(n26107), .B(n26108), .Z(n25598) );
  XNOR U27419 ( .A(round_reg[1064]), .B(round_reg[104]), .Z(n26108) );
  XOR U27420 ( .A(round_reg[1384]), .B(n26109), .Z(n26107) );
  XOR U27421 ( .A(round_reg[744]), .B(round_reg[424]), .Z(n26109) );
  AND U27422 ( .A(n23228), .B(n22498), .Z(n26103) );
  XOR U27423 ( .A(round_reg[64]), .B(n24381), .Z(n22498) );
  IV U27424 ( .A(n24305), .Z(n24381) );
  XNOR U27425 ( .A(n26110), .B(n26111), .Z(n25998) );
  XNOR U27426 ( .A(round_reg[128]), .B(round_reg[1088]), .Z(n26111) );
  XOR U27427 ( .A(round_reg[1408]), .B(n26112), .Z(n26110) );
  XOR U27428 ( .A(round_reg[768]), .B(round_reg[448]), .Z(n26112) );
  XOR U27429 ( .A(n26113), .B(n26114), .Z(n25943) );
  XNOR U27430 ( .A(round_reg[1343]), .B(round_reg[1023]), .Z(n26114) );
  XOR U27431 ( .A(round_reg[383]), .B(n26115), .Z(n26113) );
  XOR U27432 ( .A(round_reg[703]), .B(round_reg[63]), .Z(n26115) );
  XNOR U27433 ( .A(round_reg[1309]), .B(n23910), .Z(n23228) );
  XOR U27434 ( .A(n26116), .B(n25161), .Z(n23910) );
  XNOR U27435 ( .A(n26117), .B(n26118), .Z(n25161) );
  XNOR U27436 ( .A(round_reg[1373]), .B(round_reg[1053]), .Z(n26118) );
  XOR U27437 ( .A(round_reg[413]), .B(n26119), .Z(n26117) );
  XOR U27438 ( .A(round_reg[93]), .B(round_reg[733]), .Z(n26119) );
  XOR U27439 ( .A(n26120), .B(n22494), .Z(n18680) );
  XNOR U27440 ( .A(round_reg[419]), .B(n21920), .Z(n22494) );
  XOR U27441 ( .A(n25273), .B(n25186), .Z(n21920) );
  XNOR U27442 ( .A(n26121), .B(n26122), .Z(n25186) );
  XNOR U27443 ( .A(round_reg[1443]), .B(round_reg[1123]), .Z(n26122) );
  XOR U27444 ( .A(round_reg[163]), .B(n26123), .Z(n26121) );
  XOR U27445 ( .A(round_reg[803]), .B(round_reg[483]), .Z(n26123) );
  XOR U27446 ( .A(n26124), .B(n26125), .Z(n25273) );
  XNOR U27447 ( .A(round_reg[34]), .B(round_reg[1314]), .Z(n26125) );
  XOR U27448 ( .A(round_reg[354]), .B(n26126), .Z(n26124) );
  XOR U27449 ( .A(round_reg[994]), .B(round_reg[674]), .Z(n26126) );
  NOR U27450 ( .A(n23224), .B(n22493), .Z(n26120) );
  XNOR U27451 ( .A(round_reg[42]), .B(n22649), .Z(n22493) );
  XOR U27452 ( .A(n26127), .B(n26128), .Z(n25696) );
  XNOR U27453 ( .A(round_reg[106]), .B(round_reg[1066]), .Z(n26128) );
  XOR U27454 ( .A(round_reg[1386]), .B(n26129), .Z(n26127) );
  XOR U27455 ( .A(round_reg[746]), .B(round_reg[426]), .Z(n26129) );
  XOR U27456 ( .A(n26130), .B(n26131), .Z(n25438) );
  XNOR U27457 ( .A(round_reg[1577]), .B(round_reg[1257]), .Z(n26131) );
  XOR U27458 ( .A(round_reg[297]), .B(n26132), .Z(n26130) );
  XOR U27459 ( .A(round_reg[937]), .B(round_reg[617]), .Z(n26132) );
  XOR U27460 ( .A(round_reg[1592]), .B(n21775), .Z(n23224) );
  XNOR U27461 ( .A(n25871), .B(n25146), .Z(n21775) );
  XNOR U27462 ( .A(n26133), .B(n26134), .Z(n25146) );
  XNOR U27463 ( .A(round_reg[1336]), .B(round_reg[1016]), .Z(n26134) );
  XOR U27464 ( .A(round_reg[376]), .B(n26135), .Z(n26133) );
  XOR U27465 ( .A(round_reg[696]), .B(round_reg[56]), .Z(n26135) );
  XNOR U27466 ( .A(n26136), .B(n26137), .Z(n25871) );
  XNOR U27467 ( .A(round_reg[1527]), .B(round_reg[1207]), .Z(n26137) );
  XOR U27468 ( .A(round_reg[247]), .B(n26138), .Z(n26136) );
  XOR U27469 ( .A(round_reg[887]), .B(round_reg[567]), .Z(n26138) );
  XNOR U27470 ( .A(n26139), .B(n22488), .Z(n22479) );
  XOR U27471 ( .A(round_reg[368]), .B(n23445), .Z(n22488) );
  XOR U27472 ( .A(n26140), .B(n26141), .Z(n24688) );
  XNOR U27473 ( .A(round_reg[1583]), .B(round_reg[1263]), .Z(n26141) );
  XOR U27474 ( .A(round_reg[303]), .B(n26142), .Z(n26140) );
  XOR U27475 ( .A(round_reg[943]), .B(round_reg[623]), .Z(n26142) );
  XNOR U27476 ( .A(n26143), .B(n26144), .Z(n26066) );
  XNOR U27477 ( .A(round_reg[112]), .B(round_reg[1072]), .Z(n26144) );
  XOR U27478 ( .A(round_reg[1392]), .B(n26145), .Z(n26143) );
  XOR U27479 ( .A(round_reg[752]), .B(round_reg[432]), .Z(n26145) );
  ANDN U27480 ( .B(n22489), .A(n23234), .Z(n26139) );
  XOR U27481 ( .A(round_reg[1527]), .B(n23127), .Z(n23234) );
  XOR U27482 ( .A(n25057), .B(n26146), .Z(n23127) );
  XOR U27483 ( .A(n26147), .B(n26148), .Z(n25057) );
  XNOR U27484 ( .A(round_reg[1462]), .B(round_reg[1142]), .Z(n26148) );
  XOR U27485 ( .A(round_reg[182]), .B(n26149), .Z(n26147) );
  XOR U27486 ( .A(round_reg[822]), .B(round_reg[502]), .Z(n26149) );
  XNOR U27487 ( .A(round_reg[294]), .B(n22432), .Z(n22489) );
  XNOR U27488 ( .A(n26150), .B(n26151), .Z(n25768) );
  XNOR U27489 ( .A(round_reg[358]), .B(round_reg[1318]), .Z(n26151) );
  XOR U27490 ( .A(round_reg[38]), .B(n26152), .Z(n26150) );
  XOR U27491 ( .A(round_reg[998]), .B(round_reg[678]), .Z(n26152) );
  XNOR U27492 ( .A(n26153), .B(n26154), .Z(n25209) );
  XNOR U27493 ( .A(round_reg[1509]), .B(round_reg[1189]), .Z(n26154) );
  XOR U27494 ( .A(round_reg[229]), .B(n26155), .Z(n26153) );
  XOR U27495 ( .A(round_reg[869]), .B(round_reg[549]), .Z(n26155) );
  NOR U27496 ( .A(n13293), .B(n13295), .Z(n26018) );
  XNOR U27497 ( .A(n19056), .B(n21489), .Z(n13295) );
  XNOR U27498 ( .A(n26156), .B(n19574), .Z(n21489) );
  NOR U27499 ( .A(n25471), .B(n25470), .Z(n26156) );
  IV U27500 ( .A(n21082), .Z(n25471) );
  XOR U27501 ( .A(round_reg[464]), .B(n24568), .Z(n21082) );
  IV U27502 ( .A(n23577), .Z(n24568) );
  XOR U27503 ( .A(n25215), .B(n25199), .Z(n23577) );
  XNOR U27504 ( .A(n26157), .B(n26158), .Z(n25199) );
  XNOR U27505 ( .A(round_reg[1488]), .B(round_reg[1168]), .Z(n26158) );
  XOR U27506 ( .A(round_reg[208]), .B(n26159), .Z(n26157) );
  XOR U27507 ( .A(round_reg[848]), .B(round_reg[528]), .Z(n26159) );
  XOR U27508 ( .A(n26160), .B(n26161), .Z(n25215) );
  XNOR U27509 ( .A(round_reg[1359]), .B(round_reg[1039]), .Z(n26161) );
  XOR U27510 ( .A(round_reg[399]), .B(n26162), .Z(n26160) );
  XOR U27511 ( .A(round_reg[79]), .B(round_reg[719]), .Z(n26162) );
  IV U27512 ( .A(n16898), .Z(n19056) );
  XNOR U27513 ( .A(n19774), .B(n21434), .Z(n16898) );
  XNOR U27514 ( .A(n26163), .B(n26164), .Z(n21434) );
  XNOR U27515 ( .A(n18317), .B(n18561), .Z(n26164) );
  XOR U27516 ( .A(n26165), .B(n19967), .Z(n18561) );
  XOR U27517 ( .A(round_reg[1347]), .B(n21747), .Z(n19967) );
  XOR U27518 ( .A(n25286), .B(n25948), .Z(n21747) );
  XOR U27519 ( .A(n26166), .B(n26167), .Z(n25948) );
  XNOR U27520 ( .A(round_reg[2]), .B(round_reg[1282]), .Z(n26167) );
  XOR U27521 ( .A(round_reg[322]), .B(n26168), .Z(n26166) );
  XOR U27522 ( .A(round_reg[962]), .B(round_reg[642]), .Z(n26168) );
  XOR U27523 ( .A(n26169), .B(n26170), .Z(n25286) );
  XNOR U27524 ( .A(round_reg[131]), .B(round_reg[1091]), .Z(n26170) );
  XOR U27525 ( .A(round_reg[1411]), .B(n26171), .Z(n26169) );
  XOR U27526 ( .A(round_reg[771]), .B(round_reg[451]), .Z(n26171) );
  NOR U27527 ( .A(n21491), .B(n19966), .Z(n26165) );
  XNOR U27528 ( .A(round_reg[971]), .B(n21754), .Z(n19966) );
  XNOR U27529 ( .A(n26172), .B(n26173), .Z(n25663) );
  XNOR U27530 ( .A(round_reg[1546]), .B(round_reg[1226]), .Z(n26173) );
  XOR U27531 ( .A(round_reg[266]), .B(n26174), .Z(n26172) );
  XOR U27532 ( .A(round_reg[906]), .B(round_reg[586]), .Z(n26174) );
  XOR U27533 ( .A(round_reg[924]), .B(n24446), .Z(n21491) );
  IV U27534 ( .A(n24372), .Z(n24446) );
  XOR U27535 ( .A(n25546), .B(n25136), .Z(n24372) );
  XOR U27536 ( .A(n26176), .B(n26177), .Z(n25136) );
  XNOR U27537 ( .A(round_reg[28]), .B(round_reg[1308]), .Z(n26177) );
  XOR U27538 ( .A(round_reg[348]), .B(n26178), .Z(n26176) );
  XOR U27539 ( .A(round_reg[988]), .B(round_reg[668]), .Z(n26178) );
  XOR U27540 ( .A(n26179), .B(n26180), .Z(n25546) );
  XNOR U27541 ( .A(round_reg[1499]), .B(round_reg[1179]), .Z(n26180) );
  XOR U27542 ( .A(round_reg[219]), .B(n26181), .Z(n26179) );
  XOR U27543 ( .A(round_reg[859]), .B(round_reg[539]), .Z(n26181) );
  XNOR U27544 ( .A(n26182), .B(n19567), .Z(n18317) );
  XOR U27545 ( .A(round_reg[1441]), .B(n24694), .Z(n19567) );
  ANDN U27546 ( .B(n21484), .A(n19566), .Z(n26182) );
  XNOR U27547 ( .A(round_reg[1064]), .B(n25364), .Z(n19566) );
  IV U27548 ( .A(n25512), .Z(n25364) );
  XOR U27549 ( .A(n25437), .B(n24954), .Z(n25512) );
  XOR U27550 ( .A(n26183), .B(n26184), .Z(n24954) );
  XNOR U27551 ( .A(round_reg[359]), .B(round_reg[1319]), .Z(n26184) );
  XOR U27552 ( .A(round_reg[39]), .B(n26185), .Z(n26183) );
  XOR U27553 ( .A(round_reg[999]), .B(round_reg[679]), .Z(n26185) );
  XOR U27554 ( .A(n26186), .B(n26187), .Z(n25437) );
  XNOR U27555 ( .A(round_reg[1448]), .B(round_reg[1128]), .Z(n26187) );
  XOR U27556 ( .A(round_reg[168]), .B(n26188), .Z(n26186) );
  XOR U27557 ( .A(round_reg[808]), .B(round_reg[488]), .Z(n26188) );
  IV U27558 ( .A(n25457), .Z(n21484) );
  XOR U27559 ( .A(round_reg[696]), .B(n24082), .Z(n25457) );
  IV U27560 ( .A(n24208), .Z(n24082) );
  XNOR U27561 ( .A(n26189), .B(n26146), .Z(n24208) );
  XNOR U27562 ( .A(n26190), .B(n26191), .Z(n26146) );
  XNOR U27563 ( .A(round_reg[1591]), .B(round_reg[1271]), .Z(n26191) );
  XOR U27564 ( .A(round_reg[311]), .B(n26192), .Z(n26190) );
  XOR U27565 ( .A(round_reg[951]), .B(round_reg[631]), .Z(n26192) );
  XOR U27566 ( .A(n16332), .B(n26193), .Z(n26163) );
  XOR U27567 ( .A(n15907), .B(n17065), .Z(n26193) );
  XNOR U27568 ( .A(n26194), .B(n21091), .Z(n17065) );
  XOR U27569 ( .A(round_reg[1502]), .B(n22751), .Z(n21091) );
  XOR U27570 ( .A(n25669), .B(n25137), .Z(n22751) );
  XNOR U27571 ( .A(n26195), .B(n26196), .Z(n25137) );
  XNOR U27572 ( .A(round_reg[1437]), .B(round_reg[1117]), .Z(n26196) );
  XOR U27573 ( .A(round_reg[157]), .B(n26197), .Z(n26195) );
  XOR U27574 ( .A(round_reg[797]), .B(round_reg[477]), .Z(n26197) );
  XOR U27575 ( .A(n26198), .B(n26199), .Z(n25669) );
  XNOR U27576 ( .A(round_reg[1566]), .B(round_reg[1246]), .Z(n26199) );
  XOR U27577 ( .A(round_reg[286]), .B(n26200), .Z(n26198) );
  XOR U27578 ( .A(round_reg[926]), .B(round_reg[606]), .Z(n26200) );
  ANDN U27579 ( .B(n21095), .A(n21486), .Z(n26194) );
  XOR U27580 ( .A(round_reg[710]), .B(n23883), .Z(n21486) );
  XOR U27581 ( .A(n26201), .B(n26202), .Z(n23883) );
  XOR U27582 ( .A(round_reg[1113]), .B(n21613), .Z(n21095) );
  IV U27583 ( .A(n23944), .Z(n21613) );
  XOR U27584 ( .A(n24994), .B(n25527), .Z(n23944) );
  XOR U27585 ( .A(n26203), .B(n26204), .Z(n25527) );
  XNOR U27586 ( .A(round_reg[1368]), .B(round_reg[1048]), .Z(n26204) );
  XOR U27587 ( .A(round_reg[408]), .B(n26205), .Z(n26203) );
  XOR U27588 ( .A(round_reg[88]), .B(round_reg[728]), .Z(n26205) );
  XOR U27589 ( .A(n26206), .B(n26207), .Z(n24994) );
  XNOR U27590 ( .A(round_reg[1497]), .B(round_reg[1177]), .Z(n26207) );
  XOR U27591 ( .A(round_reg[217]), .B(n26208), .Z(n26206) );
  XOR U27592 ( .A(round_reg[857]), .B(round_reg[537]), .Z(n26208) );
  XOR U27593 ( .A(n24341), .B(n26210), .Z(n26209) );
  NAND U27594 ( .A(n21525), .B(n19791), .Z(n26210) );
  XOR U27595 ( .A(round_reg[1203]), .B(n24518), .Z(n19791) );
  XNOR U27596 ( .A(n26211), .B(n23828), .Z(n24518) );
  XOR U27597 ( .A(n26212), .B(n26213), .Z(n23828) );
  XNOR U27598 ( .A(round_reg[1458]), .B(round_reg[1138]), .Z(n26213) );
  XOR U27599 ( .A(round_reg[178]), .B(n26214), .Z(n26212) );
  XOR U27600 ( .A(round_reg[818]), .B(round_reg[498]), .Z(n26214) );
  XNOR U27601 ( .A(round_reg[820]), .B(n22230), .Z(n21525) );
  XNOR U27602 ( .A(n26216), .B(n26217), .Z(n25895) );
  XNOR U27603 ( .A(round_reg[115]), .B(round_reg[1075]), .Z(n26217) );
  XOR U27604 ( .A(round_reg[1395]), .B(n26218), .Z(n26216) );
  XOR U27605 ( .A(round_reg[755]), .B(round_reg[435]), .Z(n26218) );
  AND U27606 ( .A(n15691), .B(n11365), .Z(n24341) );
  IV U27607 ( .A(rc_i[5]), .Z(n11365) );
  IV U27608 ( .A(rc_i[3]), .Z(n15691) );
  XOR U27609 ( .A(round_reg[1567]), .B(n25328), .Z(n19790) );
  XNOR U27610 ( .A(n26219), .B(n19573), .Z(n16332) );
  XOR U27611 ( .A(round_reg[1284]), .B(n23016), .Z(n19573) );
  XNOR U27612 ( .A(n26220), .B(n26221), .Z(n25330) );
  XNOR U27613 ( .A(round_reg[1348]), .B(round_reg[1028]), .Z(n26221) );
  XOR U27614 ( .A(round_reg[388]), .B(n26222), .Z(n26220) );
  XOR U27615 ( .A(round_reg[708]), .B(round_reg[68]), .Z(n26222) );
  XNOR U27616 ( .A(n26223), .B(n26224), .Z(n25358) );
  XNOR U27617 ( .A(round_reg[1539]), .B(round_reg[1219]), .Z(n26224) );
  XOR U27618 ( .A(round_reg[259]), .B(n26225), .Z(n26223) );
  XOR U27619 ( .A(round_reg[899]), .B(round_reg[579]), .Z(n26225) );
  AND U27620 ( .A(n25470), .B(n19574), .Z(n26219) );
  XOR U27621 ( .A(round_reg[1275]), .B(n22517), .Z(n19574) );
  XNOR U27622 ( .A(n25129), .B(n26098), .Z(n22517) );
  XNOR U27623 ( .A(n26226), .B(n26227), .Z(n26098) );
  XNOR U27624 ( .A(round_reg[1530]), .B(round_reg[1210]), .Z(n26227) );
  XOR U27625 ( .A(round_reg[250]), .B(n26228), .Z(n26226) );
  XOR U27626 ( .A(round_reg[890]), .B(round_reg[570]), .Z(n26228) );
  XNOR U27627 ( .A(n26229), .B(n26230), .Z(n25129) );
  XNOR U27628 ( .A(round_reg[1339]), .B(round_reg[1019]), .Z(n26230) );
  XOR U27629 ( .A(round_reg[379]), .B(n26231), .Z(n26229) );
  XOR U27630 ( .A(round_reg[699]), .B(round_reg[59]), .Z(n26231) );
  XNOR U27631 ( .A(round_reg[853]), .B(n22984), .Z(n25470) );
  IV U27632 ( .A(n23664), .Z(n22984) );
  XOR U27633 ( .A(n26232), .B(n24867), .Z(n23664) );
  XOR U27634 ( .A(n26233), .B(n26234), .Z(n24867) );
  XNOR U27635 ( .A(round_reg[1428]), .B(round_reg[1108]), .Z(n26234) );
  XOR U27636 ( .A(round_reg[148]), .B(n26235), .Z(n26233) );
  XOR U27637 ( .A(round_reg[788]), .B(round_reg[468]), .Z(n26235) );
  XOR U27638 ( .A(n26236), .B(n26237), .Z(n19774) );
  XNOR U27639 ( .A(n18354), .B(n24140), .Z(n26237) );
  XNOR U27640 ( .A(n26238), .B(n24470), .Z(n24140) );
  XNOR U27641 ( .A(round_reg[695]), .B(n24715), .Z(n24470) );
  XNOR U27642 ( .A(n26239), .B(n26240), .Z(n25609) );
  XNOR U27643 ( .A(round_reg[119]), .B(round_reg[1079]), .Z(n26240) );
  XOR U27644 ( .A(round_reg[1399]), .B(n26241), .Z(n26239) );
  XOR U27645 ( .A(round_reg[759]), .B(round_reg[439]), .Z(n26241) );
  XNOR U27646 ( .A(n26242), .B(n26243), .Z(n26094) );
  XNOR U27647 ( .A(round_reg[1590]), .B(round_reg[1270]), .Z(n26243) );
  XOR U27648 ( .A(round_reg[310]), .B(n26244), .Z(n26242) );
  XOR U27649 ( .A(round_reg[950]), .B(round_reg[630]), .Z(n26244) );
  NOR U27650 ( .A(n23835), .B(n21441), .Z(n26238) );
  XOR U27651 ( .A(round_reg[220]), .B(n23253), .Z(n21441) );
  XNOR U27652 ( .A(round_reg[629]), .B(n23467), .Z(n23835) );
  XOR U27653 ( .A(n26215), .B(n25058), .Z(n23467) );
  XNOR U27654 ( .A(n26245), .B(n26246), .Z(n25058) );
  XNOR U27655 ( .A(round_reg[1333]), .B(round_reg[1013]), .Z(n26246) );
  XOR U27656 ( .A(round_reg[373]), .B(n26247), .Z(n26245) );
  XOR U27657 ( .A(round_reg[693]), .B(round_reg[53]), .Z(n26247) );
  XOR U27658 ( .A(n26248), .B(n26249), .Z(n26215) );
  XNOR U27659 ( .A(round_reg[1524]), .B(round_reg[1204]), .Z(n26249) );
  XOR U27660 ( .A(round_reg[244]), .B(n26250), .Z(n26248) );
  XOR U27661 ( .A(round_reg[884]), .B(round_reg[564]), .Z(n26250) );
  XNOR U27662 ( .A(n26251), .B(n25010), .Z(n18354) );
  IV U27663 ( .A(n24472), .Z(n25010) );
  XOR U27664 ( .A(round_reg[709]), .B(n24559), .Z(n24472) );
  IV U27665 ( .A(n23762), .Z(n24559) );
  XOR U27666 ( .A(n25729), .B(n25448), .Z(n23762) );
  XOR U27667 ( .A(n26252), .B(n26253), .Z(n25448) );
  XNOR U27668 ( .A(round_reg[133]), .B(round_reg[1093]), .Z(n26253) );
  XOR U27669 ( .A(round_reg[1413]), .B(n26254), .Z(n26252) );
  XOR U27670 ( .A(round_reg[773]), .B(round_reg[453]), .Z(n26254) );
  XOR U27671 ( .A(n26255), .B(n26256), .Z(n25729) );
  XNOR U27672 ( .A(round_reg[324]), .B(round_reg[1284]), .Z(n26256) );
  XOR U27673 ( .A(round_reg[4]), .B(n26257), .Z(n26255) );
  XOR U27674 ( .A(round_reg[964]), .B(round_reg[644]), .Z(n26257) );
  NOR U27675 ( .A(n23837), .B(n23839), .Z(n26251) );
  XNOR U27676 ( .A(round_reg[268]), .B(n23479), .Z(n23839) );
  IV U27677 ( .A(n24523), .Z(n23479) );
  XOR U27678 ( .A(n26258), .B(n25279), .Z(n24523) );
  XNOR U27679 ( .A(n26259), .B(n26260), .Z(n25279) );
  XNOR U27680 ( .A(round_reg[12]), .B(round_reg[1292]), .Z(n26260) );
  XOR U27681 ( .A(round_reg[332]), .B(n26261), .Z(n26259) );
  XOR U27682 ( .A(round_reg[972]), .B(round_reg[652]), .Z(n26261) );
  XNOR U27683 ( .A(round_reg[342]), .B(n23596), .Z(n23837) );
  XOR U27684 ( .A(n26232), .B(n25952), .Z(n23596) );
  XNOR U27685 ( .A(n26262), .B(n26263), .Z(n25952) );
  XNOR U27686 ( .A(round_reg[1366]), .B(round_reg[1046]), .Z(n26263) );
  XOR U27687 ( .A(round_reg[406]), .B(n26264), .Z(n26262) );
  XOR U27688 ( .A(round_reg[86]), .B(round_reg[726]), .Z(n26264) );
  XOR U27689 ( .A(n26265), .B(n26266), .Z(n26232) );
  XNOR U27690 ( .A(round_reg[1557]), .B(round_reg[1237]), .Z(n26266) );
  XOR U27691 ( .A(round_reg[277]), .B(n26267), .Z(n26265) );
  XOR U27692 ( .A(round_reg[917]), .B(round_reg[597]), .Z(n26267) );
  XNOR U27693 ( .A(n19349), .B(n26268), .Z(n26236) );
  XOR U27694 ( .A(n19301), .B(n24454), .Z(n26268) );
  XNOR U27695 ( .A(n26269), .B(n24476), .Z(n24454) );
  XOR U27696 ( .A(round_reg[819]), .B(n23621), .Z(n24476) );
  XNOR U27697 ( .A(n26270), .B(n26271), .Z(n25251) );
  XNOR U27698 ( .A(round_reg[114]), .B(round_reg[1074]), .Z(n26271) );
  XOR U27699 ( .A(round_reg[1394]), .B(n26272), .Z(n26270) );
  XOR U27700 ( .A(round_reg[754]), .B(round_reg[434]), .Z(n26272) );
  XOR U27701 ( .A(n26273), .B(n26274), .Z(n26039) );
  XNOR U27702 ( .A(round_reg[1523]), .B(round_reg[1203]), .Z(n26274) );
  XOR U27703 ( .A(round_reg[243]), .B(n26275), .Z(n26273) );
  XOR U27704 ( .A(round_reg[883]), .B(round_reg[563]), .Z(n26275) );
  ANDN U27705 ( .B(n24477), .A(n23185), .Z(n26269) );
  XOR U27706 ( .A(round_reg[16]), .B(n23915), .Z(n23185) );
  XNOR U27707 ( .A(n25504), .B(n25811), .Z(n23915) );
  XOR U27708 ( .A(n26276), .B(n26277), .Z(n25811) );
  XNOR U27709 ( .A(round_reg[1551]), .B(round_reg[1231]), .Z(n26277) );
  XOR U27710 ( .A(round_reg[271]), .B(n26278), .Z(n26276) );
  XOR U27711 ( .A(round_reg[911]), .B(round_reg[591]), .Z(n26278) );
  XOR U27712 ( .A(n26279), .B(n26280), .Z(n25504) );
  XNOR U27713 ( .A(round_reg[1360]), .B(round_reg[1040]), .Z(n26280) );
  XOR U27714 ( .A(round_reg[400]), .B(n26281), .Z(n26279) );
  XOR U27715 ( .A(round_reg[80]), .B(round_reg[720]), .Z(n26281) );
  XNOR U27716 ( .A(round_reg[393]), .B(n24448), .Z(n24477) );
  XNOR U27717 ( .A(n26282), .B(n26283), .Z(n25662) );
  XNOR U27718 ( .A(round_reg[137]), .B(round_reg[1097]), .Z(n26283) );
  XOR U27719 ( .A(round_reg[1417]), .B(n26284), .Z(n26282) );
  XOR U27720 ( .A(round_reg[777]), .B(round_reg[457]), .Z(n26284) );
  XNOR U27721 ( .A(n26285), .B(n26286), .Z(n24549) );
  XNOR U27722 ( .A(round_reg[328]), .B(round_reg[1288]), .Z(n26286) );
  XOR U27723 ( .A(round_reg[648]), .B(n26287), .Z(n26285) );
  XOR U27724 ( .A(round_reg[968]), .B(round_reg[8]), .Z(n26287) );
  XNOR U27725 ( .A(n26288), .B(n24981), .Z(n19301) );
  XOR U27726 ( .A(round_reg[852]), .B(n22979), .Z(n24981) );
  XNOR U27727 ( .A(n25192), .B(n24939), .Z(n22979) );
  XOR U27728 ( .A(n26289), .B(n26290), .Z(n24939) );
  XNOR U27729 ( .A(round_reg[1427]), .B(round_reg[1107]), .Z(n26290) );
  XOR U27730 ( .A(round_reg[147]), .B(n26291), .Z(n26289) );
  XOR U27731 ( .A(round_reg[787]), .B(round_reg[467]), .Z(n26291) );
  XOR U27732 ( .A(n26292), .B(n26293), .Z(n25192) );
  XNOR U27733 ( .A(round_reg[1556]), .B(round_reg[1236]), .Z(n26293) );
  XOR U27734 ( .A(round_reg[276]), .B(n26294), .Z(n26292) );
  XOR U27735 ( .A(round_reg[916]), .B(round_reg[596]), .Z(n26294) );
  ANDN U27736 ( .B(n24982), .A(n21447), .Z(n26288) );
  XNOR U27737 ( .A(round_reg[102]), .B(n23856), .Z(n21447) );
  IV U27738 ( .A(n23865), .Z(n23856) );
  XNOR U27739 ( .A(n26295), .B(n26296), .Z(n25744) );
  XNOR U27740 ( .A(round_reg[1446]), .B(round_reg[1126]), .Z(n26296) );
  XOR U27741 ( .A(round_reg[166]), .B(n26297), .Z(n26295) );
  XOR U27742 ( .A(round_reg[806]), .B(round_reg[486]), .Z(n26297) );
  XOR U27743 ( .A(round_reg[463]), .B(n23784), .Z(n24982) );
  IV U27744 ( .A(n22969), .Z(n23784) );
  XNOR U27745 ( .A(n24751), .B(n25238), .Z(n22969) );
  XNOR U27746 ( .A(n26299), .B(n26300), .Z(n25238) );
  XNOR U27747 ( .A(round_reg[1358]), .B(round_reg[1038]), .Z(n26300) );
  XOR U27748 ( .A(round_reg[398]), .B(n26301), .Z(n26299) );
  XOR U27749 ( .A(round_reg[78]), .B(round_reg[718]), .Z(n26301) );
  XOR U27750 ( .A(n26302), .B(n26303), .Z(n24751) );
  XNOR U27751 ( .A(round_reg[1487]), .B(round_reg[1167]), .Z(n26303) );
  XOR U27752 ( .A(round_reg[207]), .B(n26304), .Z(n26302) );
  XOR U27753 ( .A(round_reg[847]), .B(round_reg[527]), .Z(n26304) );
  XNOR U27754 ( .A(n26305), .B(n25004), .Z(n19349) );
  IV U27755 ( .A(n24479), .Z(n25004) );
  XOR U27756 ( .A(round_reg[923]), .B(n24294), .Z(n24479) );
  IV U27757 ( .A(n24156), .Z(n24294) );
  XNOR U27758 ( .A(n25485), .B(n26086), .Z(n24156) );
  XNOR U27759 ( .A(n26306), .B(n26307), .Z(n26086) );
  XNOR U27760 ( .A(round_reg[27]), .B(round_reg[1307]), .Z(n26307) );
  XOR U27761 ( .A(round_reg[347]), .B(n26308), .Z(n26306) );
  XOR U27762 ( .A(round_reg[987]), .B(round_reg[667]), .Z(n26308) );
  XOR U27763 ( .A(n26309), .B(n26310), .Z(n25485) );
  XNOR U27764 ( .A(round_reg[1498]), .B(round_reg[1178]), .Z(n26310) );
  XOR U27765 ( .A(round_reg[218]), .B(n26311), .Z(n26309) );
  XOR U27766 ( .A(round_reg[858]), .B(round_reg[538]), .Z(n26311) );
  ANDN U27767 ( .B(n24480), .A(n21451), .Z(n26305) );
  XNOR U27768 ( .A(round_reg[161]), .B(n24255), .Z(n21451) );
  IV U27769 ( .A(n24694), .Z(n24255) );
  XNOR U27770 ( .A(n26312), .B(n26313), .Z(n25071) );
  XNOR U27771 ( .A(round_reg[1376]), .B(round_reg[1056]), .Z(n26313) );
  XOR U27772 ( .A(round_reg[416]), .B(n26314), .Z(n26312) );
  XOR U27773 ( .A(round_reg[96]), .B(round_reg[736]), .Z(n26314) );
  XNOR U27774 ( .A(n26315), .B(n26316), .Z(n25274) );
  XNOR U27775 ( .A(round_reg[1505]), .B(round_reg[1185]), .Z(n26316) );
  XOR U27776 ( .A(round_reg[225]), .B(n26317), .Z(n26315) );
  XOR U27777 ( .A(round_reg[865]), .B(round_reg[545]), .Z(n26317) );
  XOR U27778 ( .A(round_reg[561]), .B(n23801), .Z(n24480) );
  IV U27779 ( .A(n23851), .Z(n23801) );
  XOR U27780 ( .A(n26318), .B(n25250), .Z(n23851) );
  XOR U27781 ( .A(n26319), .B(n26320), .Z(n25250) );
  XNOR U27782 ( .A(round_reg[1585]), .B(round_reg[1265]), .Z(n26320) );
  XOR U27783 ( .A(round_reg[305]), .B(n26321), .Z(n26319) );
  XOR U27784 ( .A(round_reg[945]), .B(round_reg[625]), .Z(n26321) );
  XNOR U27785 ( .A(n24792), .B(n17792), .Z(n13293) );
  IV U27786 ( .A(n18306), .Z(n17792) );
  XOR U27787 ( .A(n23458), .B(n21784), .Z(n18306) );
  XNOR U27788 ( .A(n26322), .B(n26323), .Z(n21784) );
  XNOR U27789 ( .A(n17199), .B(n20090), .Z(n26323) );
  XOR U27790 ( .A(n26324), .B(n22672), .Z(n20090) );
  XNOR U27791 ( .A(round_reg[311]), .B(n23789), .Z(n22672) );
  XNOR U27792 ( .A(n25563), .B(n25114), .Z(n23789) );
  XNOR U27793 ( .A(n26325), .B(n26326), .Z(n25114) );
  XNOR U27794 ( .A(round_reg[1335]), .B(round_reg[1015]), .Z(n26326) );
  XOR U27795 ( .A(round_reg[375]), .B(n26327), .Z(n26325) );
  XOR U27796 ( .A(round_reg[695]), .B(round_reg[55]), .Z(n26327) );
  XNOR U27797 ( .A(n26328), .B(n26329), .Z(n25563) );
  XNOR U27798 ( .A(round_reg[1526]), .B(round_reg[1206]), .Z(n26329) );
  XOR U27799 ( .A(round_reg[246]), .B(n26330), .Z(n26328) );
  XOR U27800 ( .A(round_reg[886]), .B(round_reg[566]), .Z(n26330) );
  ANDN U27801 ( .B(n22671), .A(n23380), .Z(n26324) );
  XNOR U27802 ( .A(n26331), .B(n22662), .Z(n17199) );
  XOR U27803 ( .A(round_reg[199]), .B(n24028), .Z(n22662) );
  IV U27804 ( .A(n24006), .Z(n24028) );
  XNOR U27805 ( .A(n25244), .B(n26202), .Z(n24006) );
  XNOR U27806 ( .A(n26332), .B(n26333), .Z(n26202) );
  XNOR U27807 ( .A(round_reg[134]), .B(round_reg[1094]), .Z(n26333) );
  XOR U27808 ( .A(round_reg[1414]), .B(n26334), .Z(n26332) );
  XOR U27809 ( .A(round_reg[774]), .B(round_reg[454]), .Z(n26334) );
  XOR U27810 ( .A(n26335), .B(n26336), .Z(n25244) );
  XNOR U27811 ( .A(round_reg[1543]), .B(round_reg[1223]), .Z(n26336) );
  XOR U27812 ( .A(round_reg[263]), .B(n26337), .Z(n26335) );
  XOR U27813 ( .A(round_reg[903]), .B(round_reg[583]), .Z(n26337) );
  ANDN U27814 ( .B(n22663), .A(n24796), .Z(n26331) );
  XOR U27815 ( .A(round_reg[1042]), .B(n21786), .Z(n24796) );
  XOR U27816 ( .A(n25124), .B(n25200), .Z(n21786) );
  XNOR U27817 ( .A(n26338), .B(n26339), .Z(n25200) );
  XNOR U27818 ( .A(round_reg[17]), .B(round_reg[1297]), .Z(n26339) );
  XOR U27819 ( .A(round_reg[337]), .B(n26340), .Z(n26338) );
  XOR U27820 ( .A(round_reg[977]), .B(round_reg[657]), .Z(n26340) );
  XOR U27821 ( .A(n26341), .B(n26342), .Z(n25124) );
  XNOR U27822 ( .A(round_reg[1426]), .B(round_reg[1106]), .Z(n26342) );
  XOR U27823 ( .A(round_reg[146]), .B(n26343), .Z(n26341) );
  XOR U27824 ( .A(round_reg[786]), .B(round_reg[466]), .Z(n26343) );
  XOR U27825 ( .A(round_reg[1419]), .B(n24552), .Z(n22663) );
  IV U27826 ( .A(n24237), .Z(n24552) );
  XOR U27827 ( .A(n26258), .B(n25172), .Z(n24237) );
  XOR U27828 ( .A(n26344), .B(n26345), .Z(n25172) );
  XNOR U27829 ( .A(round_reg[1354]), .B(round_reg[1034]), .Z(n26345) );
  XOR U27830 ( .A(round_reg[394]), .B(n26346), .Z(n26344) );
  XOR U27831 ( .A(round_reg[74]), .B(round_reg[714]), .Z(n26346) );
  XOR U27832 ( .A(n26347), .B(n26348), .Z(n26258) );
  XNOR U27833 ( .A(round_reg[1483]), .B(round_reg[1163]), .Z(n26348) );
  XOR U27834 ( .A(round_reg[203]), .B(n26349), .Z(n26347) );
  XOR U27835 ( .A(round_reg[843]), .B(round_reg[523]), .Z(n26349) );
  XOR U27836 ( .A(n22521), .B(n26350), .Z(n26322) );
  XOR U27837 ( .A(n17998), .B(n19338), .Z(n26350) );
  XNOR U27838 ( .A(n26351), .B(n22667), .Z(n19338) );
  XOR U27839 ( .A(round_reg[59]), .B(n22986), .Z(n22667) );
  XOR U27840 ( .A(n25793), .B(n26007), .Z(n22986) );
  XNOR U27841 ( .A(n26352), .B(n26353), .Z(n26007) );
  XNOR U27842 ( .A(round_reg[123]), .B(round_reg[1083]), .Z(n26353) );
  XOR U27843 ( .A(round_reg[1403]), .B(n26354), .Z(n26352) );
  XOR U27844 ( .A(round_reg[763]), .B(round_reg[443]), .Z(n26354) );
  XOR U27845 ( .A(n26355), .B(n26356), .Z(n25793) );
  XNOR U27846 ( .A(round_reg[1594]), .B(round_reg[1274]), .Z(n26356) );
  XOR U27847 ( .A(round_reg[314]), .B(n26357), .Z(n26355) );
  XOR U27848 ( .A(round_reg[954]), .B(round_reg[634]), .Z(n26357) );
  ANDN U27849 ( .B(n22668), .A(n23372), .Z(n26351) );
  XOR U27850 ( .A(round_reg[1181]), .B(n24887), .Z(n23372) );
  XOR U27851 ( .A(n26085), .B(n25398), .Z(n24887) );
  XNOR U27852 ( .A(n26358), .B(n26359), .Z(n25398) );
  XNOR U27853 ( .A(round_reg[1565]), .B(round_reg[1245]), .Z(n26359) );
  XOR U27854 ( .A(round_reg[285]), .B(n26360), .Z(n26358) );
  XOR U27855 ( .A(round_reg[925]), .B(round_reg[605]), .Z(n26360) );
  XOR U27856 ( .A(n26361), .B(n26362), .Z(n26085) );
  XNOR U27857 ( .A(round_reg[1436]), .B(round_reg[1116]), .Z(n26362) );
  XOR U27858 ( .A(round_reg[156]), .B(n26363), .Z(n26361) );
  XOR U27859 ( .A(round_reg[796]), .B(round_reg[476]), .Z(n26363) );
  XOR U27860 ( .A(round_reg[1545]), .B(n21185), .Z(n22668) );
  XOR U27861 ( .A(n25426), .B(n25467), .Z(n21185) );
  XNOR U27862 ( .A(n26364), .B(n26365), .Z(n25467) );
  XNOR U27863 ( .A(round_reg[329]), .B(round_reg[1289]), .Z(n26365) );
  XOR U27864 ( .A(round_reg[649]), .B(n26366), .Z(n26364) );
  XOR U27865 ( .A(round_reg[9]), .B(round_reg[969]), .Z(n26366) );
  XOR U27866 ( .A(n26367), .B(n26368), .Z(n25426) );
  XNOR U27867 ( .A(round_reg[1480]), .B(round_reg[1160]), .Z(n26368) );
  XOR U27868 ( .A(round_reg[200]), .B(n26369), .Z(n26367) );
  XOR U27869 ( .A(round_reg[840]), .B(round_reg[520]), .Z(n26369) );
  XNOR U27870 ( .A(n26370), .B(n22675), .Z(n17998) );
  XOR U27871 ( .A(round_reg[140]), .B(n24389), .Z(n22675) );
  XOR U27872 ( .A(n25459), .B(n26175), .Z(n24389) );
  XNOR U27873 ( .A(n26371), .B(n26372), .Z(n26175) );
  XNOR U27874 ( .A(round_reg[1355]), .B(round_reg[1035]), .Z(n26372) );
  XOR U27875 ( .A(round_reg[395]), .B(n26373), .Z(n26371) );
  XOR U27876 ( .A(round_reg[75]), .B(round_reg[715]), .Z(n26373) );
  XOR U27877 ( .A(n26374), .B(n26375), .Z(n25459) );
  XNOR U27878 ( .A(round_reg[1484]), .B(round_reg[1164]), .Z(n26375) );
  XOR U27879 ( .A(round_reg[204]), .B(n26376), .Z(n26374) );
  XOR U27880 ( .A(round_reg[844]), .B(round_reg[524]), .Z(n26376) );
  ANDN U27881 ( .B(n22676), .A(n23369), .Z(n26370) );
  XNOR U27882 ( .A(round_reg[1013]), .B(n21313), .Z(n23369) );
  XNOR U27883 ( .A(n25562), .B(n25607), .Z(n21313) );
  XNOR U27884 ( .A(n26377), .B(n26378), .Z(n25607) );
  XNOR U27885 ( .A(round_reg[1588]), .B(round_reg[1268]), .Z(n26378) );
  XOR U27886 ( .A(round_reg[308]), .B(n26379), .Z(n26377) );
  XOR U27887 ( .A(round_reg[948]), .B(round_reg[628]), .Z(n26379) );
  XOR U27888 ( .A(n26380), .B(n26381), .Z(n25562) );
  XNOR U27889 ( .A(round_reg[117]), .B(round_reg[1077]), .Z(n26381) );
  XOR U27890 ( .A(round_reg[1397]), .B(n26382), .Z(n26380) );
  XOR U27891 ( .A(round_reg[757]), .B(round_reg[437]), .Z(n26382) );
  XOR U27892 ( .A(round_reg[1389]), .B(n24183), .Z(n22676) );
  XNOR U27893 ( .A(n26383), .B(n26384), .Z(n25126) );
  XNOR U27894 ( .A(round_reg[1324]), .B(round_reg[1004]), .Z(n26384) );
  XOR U27895 ( .A(round_reg[364]), .B(n26385), .Z(n26383) );
  XOR U27896 ( .A(round_reg[684]), .B(round_reg[44]), .Z(n26385) );
  XNOR U27897 ( .A(n26386), .B(n26387), .Z(n24977) );
  XNOR U27898 ( .A(round_reg[1453]), .B(round_reg[1133]), .Z(n26387) );
  XOR U27899 ( .A(round_reg[173]), .B(n26388), .Z(n26386) );
  XOR U27900 ( .A(round_reg[813]), .B(round_reg[493]), .Z(n26388) );
  XNOR U27901 ( .A(n26389), .B(n22658), .Z(n22521) );
  XOR U27902 ( .A(round_reg[81]), .B(n21199), .Z(n22658) );
  ANDN U27903 ( .B(n22659), .A(n23377), .Z(n26389) );
  XOR U27904 ( .A(round_reg[1253]), .B(n25042), .Z(n23377) );
  XOR U27905 ( .A(n25439), .B(n26298), .Z(n25042) );
  XNOR U27906 ( .A(n26390), .B(n26391), .Z(n26298) );
  XNOR U27907 ( .A(round_reg[357]), .B(round_reg[1317]), .Z(n26391) );
  XOR U27908 ( .A(round_reg[37]), .B(n26392), .Z(n26390) );
  XOR U27909 ( .A(round_reg[997]), .B(round_reg[677]), .Z(n26392) );
  XOR U27910 ( .A(n26393), .B(n26394), .Z(n25439) );
  XNOR U27911 ( .A(round_reg[1508]), .B(round_reg[1188]), .Z(n26394) );
  XOR U27912 ( .A(round_reg[228]), .B(n26395), .Z(n26393) );
  XOR U27913 ( .A(round_reg[868]), .B(round_reg[548]), .Z(n26395) );
  XOR U27914 ( .A(round_reg[1326]), .B(n24828), .Z(n22659) );
  XNOR U27915 ( .A(n26048), .B(n24813), .Z(n24828) );
  XNOR U27916 ( .A(n26396), .B(n26397), .Z(n24813) );
  XNOR U27917 ( .A(round_reg[110]), .B(round_reg[1070]), .Z(n26397) );
  XOR U27918 ( .A(round_reg[1390]), .B(n26398), .Z(n26396) );
  XOR U27919 ( .A(round_reg[750]), .B(round_reg[430]), .Z(n26398) );
  XNOR U27920 ( .A(n26399), .B(n26400), .Z(n26048) );
  XNOR U27921 ( .A(round_reg[1581]), .B(round_reg[1261]), .Z(n26400) );
  XOR U27922 ( .A(round_reg[301]), .B(n26401), .Z(n26399) );
  XOR U27923 ( .A(round_reg[941]), .B(round_reg[621]), .Z(n26401) );
  XNOR U27924 ( .A(n26402), .B(n26403), .Z(n23458) );
  XNOR U27925 ( .A(n19504), .B(n17425), .Z(n26403) );
  XOR U27926 ( .A(n26404), .B(n22530), .Z(n17425) );
  XNOR U27927 ( .A(round_reg[1012]), .B(n22796), .Z(n22530) );
  XOR U27928 ( .A(n26211), .B(n25488), .Z(n22796) );
  XNOR U27929 ( .A(n26405), .B(n26406), .Z(n25488) );
  XNOR U27930 ( .A(round_reg[116]), .B(round_reg[1076]), .Z(n26406) );
  XOR U27931 ( .A(round_reg[1396]), .B(n26407), .Z(n26405) );
  XOR U27932 ( .A(round_reg[756]), .B(round_reg[436]), .Z(n26407) );
  XOR U27933 ( .A(n26408), .B(n26409), .Z(n26211) );
  XNOR U27934 ( .A(round_reg[1587]), .B(round_reg[1267]), .Z(n26409) );
  XOR U27935 ( .A(round_reg[307]), .B(n26410), .Z(n26408) );
  XOR U27936 ( .A(round_reg[947]), .B(round_reg[627]), .Z(n26410) );
  XOR U27937 ( .A(round_reg[539]), .B(n24342), .Z(n24362) );
  XOR U27938 ( .A(n25621), .B(n26047), .Z(n24342) );
  XNOR U27939 ( .A(n26411), .B(n26412), .Z(n26047) );
  XNOR U27940 ( .A(round_reg[1563]), .B(round_reg[1243]), .Z(n26412) );
  XOR U27941 ( .A(round_reg[283]), .B(n26413), .Z(n26411) );
  XOR U27942 ( .A(round_reg[923]), .B(round_reg[603]), .Z(n26413) );
  XOR U27943 ( .A(n26414), .B(n26415), .Z(n25621) );
  XNOR U27944 ( .A(round_reg[1434]), .B(round_reg[1114]), .Z(n26415) );
  XOR U27945 ( .A(round_reg[154]), .B(n26416), .Z(n26414) );
  XOR U27946 ( .A(round_reg[794]), .B(round_reg[474]), .Z(n26416) );
  XOR U27947 ( .A(round_reg[901]), .B(n22206), .Z(n22529) );
  XOR U27948 ( .A(n26201), .B(n25981), .Z(n22206) );
  XOR U27949 ( .A(n26417), .B(n26418), .Z(n25981) );
  XNOR U27950 ( .A(round_reg[1476]), .B(round_reg[1156]), .Z(n26418) );
  XOR U27951 ( .A(round_reg[196]), .B(n26419), .Z(n26417) );
  XOR U27952 ( .A(round_reg[836]), .B(round_reg[516]), .Z(n26419) );
  XOR U27953 ( .A(n26420), .B(n26421), .Z(n26201) );
  XNOR U27954 ( .A(round_reg[325]), .B(round_reg[1285]), .Z(n26421) );
  XOR U27955 ( .A(round_reg[5]), .B(n26422), .Z(n26420) );
  XOR U27956 ( .A(round_reg[965]), .B(round_reg[645]), .Z(n26422) );
  XNOR U27957 ( .A(n26423), .B(n20408), .Z(n19504) );
  XOR U27958 ( .A(round_reg[1180]), .B(n23253), .Z(n20408) );
  XNOR U27959 ( .A(n26116), .B(n26029), .Z(n23253) );
  XOR U27960 ( .A(n26424), .B(n26425), .Z(n26029) );
  XNOR U27961 ( .A(round_reg[1435]), .B(round_reg[1115]), .Z(n26425) );
  XOR U27962 ( .A(round_reg[155]), .B(n26426), .Z(n26424) );
  XOR U27963 ( .A(round_reg[795]), .B(round_reg[475]), .Z(n26426) );
  XOR U27964 ( .A(n26427), .B(n26428), .Z(n26116) );
  XNOR U27965 ( .A(round_reg[1564]), .B(round_reg[1244]), .Z(n26428) );
  XOR U27966 ( .A(round_reg[284]), .B(n26429), .Z(n26427) );
  XOR U27967 ( .A(round_reg[924]), .B(round_reg[604]), .Z(n26429) );
  ANDN U27968 ( .B(n22526), .A(n24357), .Z(n26423) );
  XOR U27969 ( .A(round_reg[435]), .B(n23475), .Z(n24357) );
  XOR U27970 ( .A(n25390), .B(n25606), .Z(n23475) );
  XNOR U27971 ( .A(n26430), .B(n26431), .Z(n25606) );
  XNOR U27972 ( .A(round_reg[1459]), .B(round_reg[1139]), .Z(n26431) );
  XOR U27973 ( .A(round_reg[179]), .B(n26432), .Z(n26430) );
  XOR U27974 ( .A(round_reg[819]), .B(round_reg[499]), .Z(n26432) );
  XOR U27975 ( .A(n26433), .B(n26434), .Z(n25390) );
  XNOR U27976 ( .A(round_reg[1330]), .B(round_reg[1010]), .Z(n26434) );
  XOR U27977 ( .A(round_reg[370]), .B(n26435), .Z(n26433) );
  XOR U27978 ( .A(round_reg[690]), .B(round_reg[50]), .Z(n26435) );
  XOR U27979 ( .A(round_reg[797]), .B(n23902), .Z(n22526) );
  IV U27980 ( .A(n24540), .Z(n23902) );
  XNOR U27981 ( .A(n25976), .B(n26046), .Z(n24540) );
  XNOR U27982 ( .A(n26436), .B(n26437), .Z(n26046) );
  XNOR U27983 ( .A(round_reg[1372]), .B(round_reg[1052]), .Z(n26437) );
  XOR U27984 ( .A(round_reg[412]), .B(n26438), .Z(n26436) );
  XOR U27985 ( .A(round_reg[92]), .B(round_reg[732]), .Z(n26438) );
  XOR U27986 ( .A(n26439), .B(n26440), .Z(n25976) );
  XNOR U27987 ( .A(round_reg[1501]), .B(round_reg[1181]), .Z(n26440) );
  XOR U27988 ( .A(round_reg[221]), .B(n26441), .Z(n26439) );
  XOR U27989 ( .A(round_reg[861]), .B(round_reg[541]), .Z(n26441) );
  XOR U27990 ( .A(n17516), .B(n26442), .Z(n26402) );
  XOR U27991 ( .A(n19078), .B(n18957), .Z(n26442) );
  XOR U27992 ( .A(n26443), .B(n20411), .Z(n18957) );
  XNOR U27993 ( .A(round_reg[1252]), .B(n25023), .Z(n20411) );
  XOR U27994 ( .A(n26444), .B(n26445), .Z(n24991) );
  XNOR U27995 ( .A(round_reg[356]), .B(round_reg[1316]), .Z(n26445) );
  XOR U27996 ( .A(round_reg[36]), .B(n26446), .Z(n26444) );
  XOR U27997 ( .A(round_reg[996]), .B(round_reg[676]), .Z(n26446) );
  XNOR U27998 ( .A(n26447), .B(n26448), .Z(n25535) );
  XNOR U27999 ( .A(round_reg[1507]), .B(round_reg[1187]), .Z(n26448) );
  XOR U28000 ( .A(round_reg[227]), .B(n26449), .Z(n26447) );
  XOR U28001 ( .A(round_reg[867]), .B(round_reg[547]), .Z(n26449) );
  ANDN U28002 ( .B(n22533), .A(n24350), .Z(n26443) );
  XNOR U28003 ( .A(round_reg[505]), .B(n25151), .Z(n24350) );
  IV U28004 ( .A(n24296), .Z(n25151) );
  XOR U28005 ( .A(n26189), .B(n25843), .Z(n24296) );
  XNOR U28006 ( .A(n26450), .B(n26451), .Z(n25843) );
  XNOR U28007 ( .A(round_reg[1529]), .B(round_reg[1209]), .Z(n26451) );
  XOR U28008 ( .A(round_reg[249]), .B(n26452), .Z(n26450) );
  XOR U28009 ( .A(round_reg[889]), .B(round_reg[569]), .Z(n26452) );
  XOR U28010 ( .A(n26453), .B(n26454), .Z(n26189) );
  XNOR U28011 ( .A(round_reg[120]), .B(round_reg[1080]), .Z(n26454) );
  XOR U28012 ( .A(round_reg[1400]), .B(n26455), .Z(n26453) );
  XOR U28013 ( .A(round_reg[760]), .B(round_reg[440]), .Z(n26455) );
  XOR U28014 ( .A(round_reg[894]), .B(n23588), .Z(n22533) );
  XOR U28015 ( .A(n25026), .B(n24822), .Z(n23588) );
  XNOR U28016 ( .A(n26456), .B(n26457), .Z(n24822) );
  XNOR U28017 ( .A(round_reg[1469]), .B(round_reg[1149]), .Z(n26457) );
  XOR U28018 ( .A(round_reg[189]), .B(n26458), .Z(n26456) );
  XOR U28019 ( .A(round_reg[829]), .B(round_reg[509]), .Z(n26458) );
  XOR U28020 ( .A(n26459), .B(n26460), .Z(n25026) );
  XNOR U28021 ( .A(round_reg[1598]), .B(round_reg[1278]), .Z(n26460) );
  XOR U28022 ( .A(round_reg[318]), .B(n26461), .Z(n26459) );
  XOR U28023 ( .A(round_reg[958]), .B(round_reg[638]), .Z(n26461) );
  XNOR U28024 ( .A(n26462), .B(n20416), .Z(n19078) );
  XOR U28025 ( .A(round_reg[1041]), .B(n21199), .Z(n20416) );
  XOR U28026 ( .A(n24750), .B(n25109), .Z(n21199) );
  XNOR U28027 ( .A(n26463), .B(n26464), .Z(n25109) );
  XNOR U28028 ( .A(round_reg[1425]), .B(round_reg[1105]), .Z(n26464) );
  XOR U28029 ( .A(round_reg[145]), .B(n26465), .Z(n26463) );
  XOR U28030 ( .A(round_reg[785]), .B(round_reg[465]), .Z(n26465) );
  XOR U28031 ( .A(n26466), .B(n26467), .Z(n24750) );
  XNOR U28032 ( .A(round_reg[16]), .B(round_reg[1296]), .Z(n26467) );
  XOR U28033 ( .A(round_reg[336]), .B(n26468), .Z(n26466) );
  XOR U28034 ( .A(round_reg[976]), .B(round_reg[656]), .Z(n26468) );
  AND U28035 ( .A(n24352), .B(n22535), .Z(n26462) );
  XNOR U28036 ( .A(round_reg[673]), .B(n24815), .Z(n22535) );
  XOR U28037 ( .A(n25033), .B(n25748), .Z(n24815) );
  XNOR U28038 ( .A(n26469), .B(n26470), .Z(n25748) );
  XNOR U28039 ( .A(round_reg[1377]), .B(round_reg[1057]), .Z(n26470) );
  XOR U28040 ( .A(round_reg[417]), .B(n26471), .Z(n26469) );
  XOR U28041 ( .A(round_reg[97]), .B(round_reg[737]), .Z(n26471) );
  XNOR U28042 ( .A(n26472), .B(n26473), .Z(n25033) );
  XNOR U28043 ( .A(round_reg[1568]), .B(round_reg[1248]), .Z(n26473) );
  XOR U28044 ( .A(round_reg[288]), .B(n26474), .Z(n26472) );
  XOR U28045 ( .A(round_reg[928]), .B(round_reg[608]), .Z(n26474) );
  XOR U28046 ( .A(round_reg[607]), .B(n25328), .Z(n24352) );
  XOR U28047 ( .A(n25160), .B(n25818), .Z(n25328) );
  XNOR U28048 ( .A(n26475), .B(n26476), .Z(n25818) );
  XNOR U28049 ( .A(round_reg[31]), .B(round_reg[1311]), .Z(n26476) );
  XOR U28050 ( .A(round_reg[351]), .B(n26477), .Z(n26475) );
  XOR U28051 ( .A(round_reg[991]), .B(round_reg[671]), .Z(n26477) );
  XNOR U28052 ( .A(n26478), .B(n26479), .Z(n25160) );
  XNOR U28053 ( .A(round_reg[1502]), .B(round_reg[1182]), .Z(n26479) );
  XOR U28054 ( .A(round_reg[222]), .B(n26480), .Z(n26478) );
  XOR U28055 ( .A(round_reg[862]), .B(round_reg[542]), .Z(n26480) );
  XNOR U28056 ( .A(n26481), .B(n20403), .Z(n17516) );
  XOR U28057 ( .A(round_reg[1090]), .B(n24161), .Z(n20403) );
  XOR U28058 ( .A(n24910), .B(n25681), .Z(n24161) );
  XNOR U28059 ( .A(n26482), .B(n26483), .Z(n25681) );
  XNOR U28060 ( .A(round_reg[1474]), .B(round_reg[1154]), .Z(n26483) );
  XOR U28061 ( .A(round_reg[194]), .B(n26484), .Z(n26482) );
  XOR U28062 ( .A(round_reg[834]), .B(round_reg[514]), .Z(n26484) );
  XOR U28063 ( .A(n26485), .B(n26486), .Z(n24910) );
  XNOR U28064 ( .A(round_reg[1345]), .B(round_reg[1025]), .Z(n26486) );
  XOR U28065 ( .A(round_reg[385]), .B(n26487), .Z(n26485) );
  XOR U28066 ( .A(round_reg[705]), .B(round_reg[65]), .Z(n26487) );
  AND U28067 ( .A(n24359), .B(n22537), .Z(n26481) );
  XNOR U28068 ( .A(round_reg[751]), .B(n23241), .Z(n22537) );
  XNOR U28069 ( .A(n26488), .B(n26489), .Z(n25393) );
  XNOR U28070 ( .A(round_reg[1455]), .B(round_reg[1135]), .Z(n26489) );
  XOR U28071 ( .A(round_reg[175]), .B(n26490), .Z(n26488) );
  XOR U28072 ( .A(round_reg[815]), .B(round_reg[495]), .Z(n26490) );
  XOR U28073 ( .A(n26491), .B(n26492), .Z(n25073) );
  XNOR U28074 ( .A(round_reg[1326]), .B(round_reg[1006]), .Z(n26492) );
  XOR U28075 ( .A(round_reg[366]), .B(n26493), .Z(n26491) );
  XOR U28076 ( .A(round_reg[686]), .B(round_reg[46]), .Z(n26493) );
  XNOR U28077 ( .A(round_reg[320]), .B(n23811), .Z(n24359) );
  IV U28078 ( .A(n24538), .Z(n23811) );
  XOR U28079 ( .A(n25932), .B(n24337), .Z(n24538) );
  XOR U28080 ( .A(n26494), .B(n26495), .Z(n24337) );
  XNOR U28081 ( .A(round_reg[1344]), .B(round_reg[1024]), .Z(n26495) );
  XOR U28082 ( .A(round_reg[384]), .B(n26496), .Z(n26494) );
  XOR U28083 ( .A(round_reg[704]), .B(round_reg[64]), .Z(n26496) );
  XOR U28084 ( .A(n26497), .B(n26498), .Z(n25932) );
  XNOR U28085 ( .A(round_reg[1599]), .B(round_reg[1279]), .Z(n26498) );
  XOR U28086 ( .A(round_reg[319]), .B(n26499), .Z(n26497) );
  XOR U28087 ( .A(round_reg[959]), .B(round_reg[639]), .Z(n26499) );
  XNOR U28088 ( .A(n26500), .B(n22671), .Z(n24792) );
  XOR U28089 ( .A(round_reg[1480]), .B(n21783), .Z(n22671) );
  XOR U28090 ( .A(n25154), .B(n25481), .Z(n21783) );
  XNOR U28091 ( .A(n26501), .B(n26502), .Z(n25481) );
  XNOR U28092 ( .A(round_reg[135]), .B(round_reg[1095]), .Z(n26502) );
  XOR U28093 ( .A(round_reg[1415]), .B(n26503), .Z(n26501) );
  XOR U28094 ( .A(round_reg[775]), .B(round_reg[455]), .Z(n26503) );
  XOR U28095 ( .A(n26504), .B(n26505), .Z(n25154) );
  XNOR U28096 ( .A(round_reg[1544]), .B(round_reg[1224]), .Z(n26505) );
  XOR U28097 ( .A(round_reg[264]), .B(n26506), .Z(n26504) );
  XOR U28098 ( .A(round_reg[904]), .B(round_reg[584]), .Z(n26506) );
  ANDN U28099 ( .B(n23380), .A(n23381), .Z(n26500) );
  XOR U28100 ( .A(round_reg[752]), .B(n24770), .Z(n23381) );
  IV U28101 ( .A(n25294), .Z(n24770) );
  XNOR U28102 ( .A(n26318), .B(n25904), .Z(n25294) );
  XNOR U28103 ( .A(n26507), .B(n26508), .Z(n25904) );
  XNOR U28104 ( .A(round_reg[1327]), .B(round_reg[1007]), .Z(n26508) );
  XOR U28105 ( .A(round_reg[367]), .B(n26509), .Z(n26507) );
  XOR U28106 ( .A(round_reg[687]), .B(round_reg[47]), .Z(n26509) );
  XOR U28107 ( .A(n26510), .B(n26511), .Z(n26318) );
  XNOR U28108 ( .A(round_reg[1456]), .B(round_reg[1136]), .Z(n26511) );
  XOR U28109 ( .A(round_reg[176]), .B(n26512), .Z(n26510) );
  XOR U28110 ( .A(round_reg[816]), .B(round_reg[496]), .Z(n26512) );
  XOR U28111 ( .A(round_reg[1091]), .B(n22757), .Z(n23380) );
  XOR U28112 ( .A(n25730), .B(n24880), .Z(n22757) );
  XNOR U28113 ( .A(n26513), .B(n26514), .Z(n24880) );
  XNOR U28114 ( .A(round_reg[1346]), .B(round_reg[1026]), .Z(n26514) );
  XOR U28115 ( .A(round_reg[386]), .B(n26515), .Z(n26513) );
  XOR U28116 ( .A(round_reg[706]), .B(round_reg[66]), .Z(n26515) );
  XOR U28117 ( .A(n26516), .B(n26517), .Z(n25730) );
  XNOR U28118 ( .A(round_reg[1475]), .B(round_reg[1155]), .Z(n26517) );
  XOR U28119 ( .A(round_reg[195]), .B(n26518), .Z(n26516) );
  XOR U28120 ( .A(round_reg[835]), .B(round_reg[515]), .Z(n26518) );
  IV U28121 ( .A(init), .Z(n1032) );
endmodule

