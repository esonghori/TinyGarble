
module mult_N128_CC2 ( clk, rst, a, b, c );
  input [127:0] a;
  input [63:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593,
         n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
         n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
         n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
         n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
         n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
         n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
         n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665,
         n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
         n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
         n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
         n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
         n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713,
         n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737,
         n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
         n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
         n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
         n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
         n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857,
         n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
         n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
         n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
         n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
         n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
         n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929,
         n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
         n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
         n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
         n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
         n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
         n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
         n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
         n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
         n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
         n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
         n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
         n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
         n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097,
         n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
         n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
         n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
         n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
         n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
         n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
         n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
         n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169,
         n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
         n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
         n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
         n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201,
         n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
         n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217,
         n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
         n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
         n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
         n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
         n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
         n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
         n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273,
         n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
         n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
         n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
         n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
         n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313,
         n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
         n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
         n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337,
         n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345,
         n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
         n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361,
         n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
         n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377,
         n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385,
         n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393,
         n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
         n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409,
         n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417,
         n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
         n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433,
         n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
         n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449,
         n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
         n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
         n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
         n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
         n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489,
         n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
         n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505,
         n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
         n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521,
         n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529,
         n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537,
         n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
         n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553,
         n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
         n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
         n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577,
         n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
         n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593,
         n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601,
         n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609,
         n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
         n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625,
         n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633,
         n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641,
         n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649,
         n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
         n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
         n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673,
         n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681,
         n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
         n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697,
         n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705,
         n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
         n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721,
         n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
         n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737,
         n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745,
         n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753,
         n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
         n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769,
         n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777,
         n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785,
         n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793,
         n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
         n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809,
         n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817,
         n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825,
         n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
         n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841,
         n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849,
         n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857,
         n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865,
         n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
         n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881,
         n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889,
         n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897,
         n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
         n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913,
         n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921,
         n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
         n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937,
         n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
         n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953,
         n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961,
         n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
         n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
         n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985,
         n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993,
         n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
         n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009,
         n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017,
         n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025,
         n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033,
         n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
         n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049,
         n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057,
         n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065,
         n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
         n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081,
         n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089,
         n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097,
         n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105,
         n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113,
         n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121,
         n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129,
         n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137,
         n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
         n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153,
         n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
         n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169,
         n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177,
         n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185,
         n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
         n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201,
         n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209,
         n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217,
         n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225,
         n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233,
         n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241,
         n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249,
         n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257,
         n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265,
         n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273,
         n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281,
         n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289,
         n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297,
         n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305,
         n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313,
         n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321,
         n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
         n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
         n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345,
         n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353,
         n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361,
         n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369,
         n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377,
         n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385,
         n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393,
         n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
         n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409,
         n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417,
         n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425,
         n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433,
         n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441,
         n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449,
         n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457,
         n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465,
         n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
         n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481,
         n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489,
         n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497,
         n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
         n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513,
         n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521,
         n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529,
         n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537,
         n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545,
         n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553,
         n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561,
         n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569,
         n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577,
         n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585,
         n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593,
         n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601,
         n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609,
         n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617,
         n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625,
         n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633,
         n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641,
         n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
         n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657,
         n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665,
         n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
         n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681,
         n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
         n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697,
         n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705,
         n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713,
         n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
         n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729,
         n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
         n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745,
         n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
         n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761,
         n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
         n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777,
         n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785,
         n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
         n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801,
         n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
         n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
         n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825,
         n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
         n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841,
         n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849,
         n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857,
         n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865,
         n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873,
         n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
         n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889,
         n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897,
         n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905,
         n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913,
         n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921,
         n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929,
         n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
         n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945,
         n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
         n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961,
         n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969,
         n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977,
         n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985,
         n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993,
         n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001,
         n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009,
         n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017,
         n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025,
         n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
         n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041,
         n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
         n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
         n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065,
         n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073,
         n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081,
         n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089,
         n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097,
         n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105,
         n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113,
         n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121,
         n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129,
         n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137,
         n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145,
         n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153,
         n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161,
         n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169,
         n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177,
         n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185,
         n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193,
         n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201,
         n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209,
         n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217,
         n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225,
         n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233,
         n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241,
         n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249,
         n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257,
         n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265,
         n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273,
         n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281,
         n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289,
         n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
         n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305,
         n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313,
         n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321,
         n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329,
         n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337,
         n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345,
         n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353,
         n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361,
         n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369,
         n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377,
         n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385,
         n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
         n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401,
         n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409,
         n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417,
         n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425,
         n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433,
         n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441,
         n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449,
         n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457,
         n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
         n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473,
         n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481,
         n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
         n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497,
         n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505,
         n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513,
         n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521,
         n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529,
         n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537,
         n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545,
         n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553,
         n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561,
         n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569,
         n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577,
         n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
         n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593,
         n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
         n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609,
         n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617,
         n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625,
         n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633,
         n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641,
         n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649,
         n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657,
         n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665,
         n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
         n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681,
         n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689,
         n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697,
         n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705,
         n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713,
         n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721,
         n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
         n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737,
         n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
         n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753,
         n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761,
         n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769,
         n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777,
         n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785,
         n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793,
         n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801,
         n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809,
         n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
         n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825,
         n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833,
         n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841,
         n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849,
         n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857,
         n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865,
         n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873,
         n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881,
         n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
         n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897,
         n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905,
         n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913,
         n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921,
         n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929,
         n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937,
         n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945,
         n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
         n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
         n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969,
         n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977,
         n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985,
         n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993,
         n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001,
         n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009,
         n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
         n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
         n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
         n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041,
         n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049,
         n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057,
         n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065,
         n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073,
         n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081,
         n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
         n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097,
         n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105,
         n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113,
         n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121,
         n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129,
         n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137,
         n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145,
         n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153,
         n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
         n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
         n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177,
         n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185,
         n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193,
         n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201,
         n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209,
         n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217,
         n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225,
         n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
         n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241,
         n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249,
         n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257,
         n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265,
         n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273,
         n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281,
         n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289,
         n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297,
         n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
         n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313,
         n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
         n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329,
         n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337,
         n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345,
         n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353,
         n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361,
         n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369,
         n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
         n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385,
         n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393,
         n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401,
         n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409,
         n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417,
         n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425,
         n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433,
         n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441,
         n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
         n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457,
         n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465,
         n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473,
         n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481,
         n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489,
         n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497,
         n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505,
         n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513,
         n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
         n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529,
         n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537,
         n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545,
         n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553,
         n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561,
         n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569,
         n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577,
         n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585,
         n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593,
         n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601,
         n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609,
         n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617,
         n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625,
         n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633,
         n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641,
         n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649,
         n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657,
         n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665,
         n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673,
         n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681,
         n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689,
         n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697,
         n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705,
         n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713,
         n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721,
         n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729,
         n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737,
         n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745,
         n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753,
         n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761,
         n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769,
         n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777,
         n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785,
         n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793,
         n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801,
         n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809,
         n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817,
         n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825,
         n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833,
         n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841,
         n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849,
         n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857,
         n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865,
         n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873,
         n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881,
         n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889,
         n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897,
         n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905,
         n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913,
         n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921,
         n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929,
         n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937,
         n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945,
         n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953,
         n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961,
         n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969,
         n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977,
         n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985,
         n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993,
         n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001,
         n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009,
         n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017,
         n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025,
         n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033,
         n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041,
         n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049,
         n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057,
         n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065,
         n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073,
         n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081,
         n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089,
         n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097,
         n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105,
         n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113,
         n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121,
         n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129,
         n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137,
         n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145,
         n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153,
         n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161,
         n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169,
         n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177,
         n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185,
         n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193,
         n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201,
         n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209,
         n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217,
         n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225,
         n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233,
         n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241,
         n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249,
         n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257,
         n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265,
         n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273,
         n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281,
         n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289,
         n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297,
         n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305,
         n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313,
         n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321,
         n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329,
         n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337,
         n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345,
         n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353,
         n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361,
         n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369,
         n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377,
         n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385,
         n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393,
         n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401,
         n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409,
         n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417,
         n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425,
         n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433,
         n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441,
         n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449,
         n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457,
         n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465,
         n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473,
         n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481,
         n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489,
         n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497,
         n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505,
         n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513,
         n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521,
         n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529,
         n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537,
         n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545,
         n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553,
         n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561,
         n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569,
         n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577,
         n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585,
         n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593,
         n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601,
         n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609,
         n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617,
         n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625,
         n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633,
         n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641,
         n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649,
         n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657,
         n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665,
         n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673,
         n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681,
         n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689,
         n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697,
         n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705,
         n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713,
         n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721,
         n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729,
         n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737,
         n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745,
         n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753,
         n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761,
         n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769,
         n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777,
         n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785,
         n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793,
         n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801,
         n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809,
         n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817,
         n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825,
         n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833,
         n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841,
         n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849,
         n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857,
         n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865,
         n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873,
         n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881,
         n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889,
         n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897,
         n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905,
         n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913,
         n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921,
         n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929,
         n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937,
         n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945,
         n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953,
         n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961,
         n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969,
         n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977,
         n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985,
         n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993,
         n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001,
         n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009,
         n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017,
         n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025,
         n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033,
         n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041,
         n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049,
         n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057,
         n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065,
         n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073,
         n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081,
         n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089,
         n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097,
         n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105,
         n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113,
         n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121,
         n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129,
         n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137,
         n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145,
         n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153,
         n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161,
         n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169,
         n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177,
         n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185,
         n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193,
         n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201,
         n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209,
         n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217,
         n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225,
         n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233,
         n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241,
         n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249,
         n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257,
         n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265,
         n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273,
         n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281,
         n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289,
         n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297,
         n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305,
         n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313,
         n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321,
         n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329,
         n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337,
         n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345,
         n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353,
         n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361,
         n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369,
         n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377,
         n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385,
         n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393,
         n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401,
         n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409,
         n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417,
         n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425,
         n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433,
         n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441,
         n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449,
         n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457,
         n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465,
         n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473,
         n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481,
         n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489,
         n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497,
         n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505,
         n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513,
         n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521,
         n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529,
         n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537,
         n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545,
         n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553,
         n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561,
         n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569,
         n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577,
         n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585,
         n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593,
         n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601,
         n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609,
         n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617,
         n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625,
         n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633,
         n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641,
         n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649,
         n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657,
         n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665,
         n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673,
         n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681,
         n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689,
         n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697,
         n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705,
         n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713,
         n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721,
         n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729,
         n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737,
         n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745,
         n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753,
         n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761,
         n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769,
         n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777,
         n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785,
         n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793,
         n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801,
         n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809,
         n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817,
         n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825,
         n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833,
         n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841,
         n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849,
         n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857,
         n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865,
         n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873,
         n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881,
         n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889,
         n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897,
         n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905,
         n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913,
         n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921,
         n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929,
         n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937,
         n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945,
         n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953,
         n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961,
         n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969,
         n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977,
         n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985,
         n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993,
         n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001,
         n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009,
         n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017,
         n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025,
         n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033,
         n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041,
         n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049,
         n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057,
         n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065,
         n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073,
         n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081,
         n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089,
         n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097,
         n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105,
         n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113,
         n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121,
         n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129,
         n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137,
         n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145,
         n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153,
         n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161,
         n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169,
         n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177,
         n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185,
         n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193,
         n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201,
         n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209,
         n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217,
         n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225,
         n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233,
         n32234, n32235, n32236, n32237, n32238, n32239, n32240, n32241,
         n32242, n32243, n32244, n32245, n32246, n32247, n32248, n32249,
         n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257,
         n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265,
         n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273,
         n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281,
         n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289,
         n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297,
         n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305,
         n32306, n32307, n32308, n32309, n32310, n32311, n32312, n32313,
         n32314, n32315, n32316, n32317, n32318, n32319, n32320, n32321,
         n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329,
         n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337,
         n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345,
         n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353,
         n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361,
         n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369,
         n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377,
         n32378, n32379, n32380, n32381, n32382, n32383, n32384, n32385,
         n32386, n32387, n32388, n32389, n32390, n32391, n32392, n32393,
         n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401,
         n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409,
         n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417,
         n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425,
         n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433,
         n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441,
         n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449,
         n32450, n32451, n32452, n32453, n32454, n32455, n32456, n32457,
         n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465,
         n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473,
         n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481,
         n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489,
         n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497,
         n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505,
         n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513,
         n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521,
         n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529,
         n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537,
         n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545,
         n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553,
         n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561,
         n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569,
         n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577,
         n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585,
         n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593,
         n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601,
         n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609,
         n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617,
         n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625,
         n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633,
         n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641,
         n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649,
         n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657,
         n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665,
         n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673,
         n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681,
         n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689,
         n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697,
         n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705,
         n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713,
         n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721,
         n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729,
         n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737,
         n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745,
         n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753,
         n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761,
         n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769,
         n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777,
         n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785,
         n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793,
         n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801,
         n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809,
         n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817,
         n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825,
         n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833,
         n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841,
         n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849,
         n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857,
         n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865,
         n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873,
         n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881,
         n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889,
         n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897,
         n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905,
         n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913,
         n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921,
         n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929,
         n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937,
         n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945,
         n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953,
         n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961,
         n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969,
         n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977,
         n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985,
         n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993,
         n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001,
         n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009,
         n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017,
         n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025,
         n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033,
         n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041,
         n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049,
         n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057,
         n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065,
         n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073,
         n33074, n33075, n33076, n33077, n33078, n33079, n33080, n33081,
         n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089,
         n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097,
         n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105,
         n33106, n33107, n33108, n33109, n33110, n33111, n33112, n33113,
         n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121,
         n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129,
         n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137,
         n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145,
         n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153,
         n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161,
         n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169,
         n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177,
         n33178, n33179, n33180, n33181, n33182, n33183, n33184, n33185,
         n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193,
         n33194, n33195, n33196, n33197, n33198, n33199, n33200, n33201,
         n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209,
         n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217,
         n33218, n33219, n33220, n33221, n33222, n33223, n33224, n33225,
         n33226, n33227, n33228, n33229, n33230, n33231, n33232, n33233,
         n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241,
         n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249,
         n33250, n33251, n33252, n33253, n33254, n33255, n33256, n33257,
         n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265,
         n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273,
         n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281,
         n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289,
         n33290, n33291, n33292, n33293, n33294, n33295, n33296, n33297,
         n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305,
         n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313,
         n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321,
         n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329,
         n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337,
         n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345,
         n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33353,
         n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361,
         n33362, n33363, n33364, n33365, n33366, n33367, n33368, n33369,
         n33370, n33371, n33372, n33373, n33374, n33375, n33376, n33377,
         n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385,
         n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393,
         n33394, n33395, n33396, n33397, n33398, n33399, n33400, n33401,
         n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409,
         n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417,
         n33418, n33419, n33420, n33421, n33422, n33423, n33424, n33425,
         n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433,
         n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441,
         n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449,
         n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457,
         n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465,
         n33466, n33467, n33468, n33469, n33470, n33471, n33472, n33473,
         n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481,
         n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489,
         n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497,
         n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505,
         n33506, n33507, n33508, n33509, n33510, n33511, n33512, n33513,
         n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521,
         n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529,
         n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537,
         n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545,
         n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553,
         n33554, n33555, n33556, n33557, n33558, n33559, n33560, n33561,
         n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569,
         n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577,
         n33578, n33579, n33580, n33581, n33582, n33583, n33584, n33585,
         n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593,
         n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601,
         n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609,
         n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617,
         n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625,
         n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633,
         n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641,
         n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649,
         n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657,
         n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665,
         n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673,
         n33674, n33675, n33676, n33677, n33678, n33679, n33680, n33681,
         n33682, n33683, n33684, n33685, n33686, n33687, n33688, n33689,
         n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697,
         n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705,
         n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713,
         n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721,
         n33722, n33723, n33724, n33725, n33726, n33727, n33728, n33729,
         n33730, n33731, n33732, n33733, n33734, n33735, n33736, n33737,
         n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745,
         n33746, n33747, n33748, n33749, n33750, n33751, n33752, n33753,
         n33754, n33755, n33756, n33757, n33758, n33759, n33760, n33761,
         n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769,
         n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777,
         n33778, n33779, n33780, n33781, n33782, n33783, n33784, n33785,
         n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793,
         n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801,
         n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809,
         n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817,
         n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825,
         n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833,
         n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841,
         n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849,
         n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857,
         n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865,
         n33866, n33867, n33868, n33869, n33870, n33871, n33872, n33873,
         n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881,
         n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889,
         n33890, n33891, n33892, n33893, n33894, n33895, n33896, n33897,
         n33898, n33899, n33900, n33901, n33902, n33903, n33904, n33905,
         n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913,
         n33914, n33915, n33916, n33917, n33918, n33919, n33920, n33921,
         n33922, n33923, n33924, n33925, n33926, n33927, n33928, n33929,
         n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937,
         n33938, n33939, n33940, n33941, n33942, n33943, n33944, n33945,
         n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953,
         n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961,
         n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969,
         n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977,
         n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985,
         n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993,
         n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001,
         n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009,
         n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017,
         n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025,
         n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033,
         n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041,
         n34042, n34043, n34044, n34045, n34046, n34047, n34048, n34049,
         n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057,
         n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065,
         n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073,
         n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081,
         n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089,
         n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097,
         n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105,
         n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113,
         n34114, n34115, n34116, n34117, n34118, n34119, n34120, n34121,
         n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129,
         n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137,
         n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145,
         n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153,
         n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161,
         n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169,
         n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177,
         n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185,
         n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193,
         n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201,
         n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209,
         n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217,
         n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225,
         n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233,
         n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241,
         n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249,
         n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257,
         n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265,
         n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273,
         n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281,
         n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289,
         n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297,
         n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305,
         n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313,
         n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321,
         n34322, n34323, n34324, n34325, n34326, n34327, n34328, n34329,
         n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337,
         n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345,
         n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353,
         n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361,
         n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369,
         n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377,
         n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385,
         n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393,
         n34394, n34395, n34396, n34397, n34398, n34399, n34400, n34401,
         n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409,
         n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417,
         n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425,
         n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433,
         n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441,
         n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449,
         n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457,
         n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465,
         n34466, n34467, n34468, n34469, n34470, n34471, n34472, n34473,
         n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481,
         n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489,
         n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497,
         n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505,
         n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513,
         n34514, n34515, n34516, n34517, n34518, n34519, n34520, n34521,
         n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529,
         n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537,
         n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545,
         n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553,
         n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561,
         n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569,
         n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577,
         n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585,
         n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593,
         n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601,
         n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609,
         n34610, n34611, n34612, n34613, n34614, n34615, n34616, n34617,
         n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625,
         n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633,
         n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641,
         n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649,
         n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657,
         n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665,
         n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673,
         n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681,
         n34682, n34683, n34684, n34685, n34686, n34687, n34688, n34689,
         n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697,
         n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705,
         n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713,
         n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721,
         n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729,
         n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737,
         n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745,
         n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753,
         n34754, n34755, n34756, n34757, n34758, n34759, n34760, n34761,
         n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769,
         n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777,
         n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785,
         n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793,
         n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801,
         n34802, n34803, n34804, n34805, n34806, n34807, n34808, n34809,
         n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817,
         n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825,
         n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833,
         n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841,
         n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849,
         n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857,
         n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865,
         n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873,
         n34874, n34875, n34876, n34877, n34878, n34879, n34880, n34881,
         n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889,
         n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897,
         n34898, n34899, n34900, n34901, n34902, n34903, n34904, n34905,
         n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913,
         n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921,
         n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929,
         n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937,
         n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945,
         n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953,
         n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961,
         n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969,
         n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977,
         n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985,
         n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993,
         n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001,
         n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009,
         n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017,
         n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025,
         n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033,
         n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041,
         n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049,
         n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057,
         n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065,
         n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073,
         n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081,
         n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089,
         n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097,
         n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105,
         n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113,
         n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121,
         n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129,
         n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137,
         n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145,
         n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153,
         n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161,
         n35162, n35163, n35164, n35165, n35166, n35167, n35168, n35169,
         n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177,
         n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185,
         n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193,
         n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201,
         n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209,
         n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217,
         n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225,
         n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233,
         n35234, n35235, n35236, n35237, n35238, n35239, n35240, n35241,
         n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249,
         n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257,
         n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265,
         n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273,
         n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281,
         n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289,
         n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297,
         n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305,
         n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313,
         n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321,
         n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329,
         n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337,
         n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345,
         n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353,
         n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361,
         n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369,
         n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377,
         n35378, n35379, n35380, n35381, n35382, n35383, n35384, n35385,
         n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393,
         n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401,
         n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35409,
         n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417,
         n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425,
         n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433,
         n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441,
         n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449,
         n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457,
         n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465,
         n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473,
         n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481,
         n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489,
         n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497,
         n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505,
         n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513,
         n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521,
         n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529,
         n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537,
         n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545,
         n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553,
         n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561,
         n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569,
         n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577;
  wire   [127:64] swire;
  wire   [255:128] sreg;

  DFF \sreg_reg[128]  ( .D(swire[64]), .CLK(clk), .RST(rst), .Q(sreg[128]) );
  DFF \sreg_reg[129]  ( .D(swire[65]), .CLK(clk), .RST(rst), .Q(sreg[129]) );
  DFF \sreg_reg[130]  ( .D(swire[66]), .CLK(clk), .RST(rst), .Q(sreg[130]) );
  DFF \sreg_reg[131]  ( .D(swire[67]), .CLK(clk), .RST(rst), .Q(sreg[131]) );
  DFF \sreg_reg[132]  ( .D(swire[68]), .CLK(clk), .RST(rst), .Q(sreg[132]) );
  DFF \sreg_reg[133]  ( .D(swire[69]), .CLK(clk), .RST(rst), .Q(sreg[133]) );
  DFF \sreg_reg[134]  ( .D(swire[70]), .CLK(clk), .RST(rst), .Q(sreg[134]) );
  DFF \sreg_reg[135]  ( .D(swire[71]), .CLK(clk), .RST(rst), .Q(sreg[135]) );
  DFF \sreg_reg[136]  ( .D(swire[72]), .CLK(clk), .RST(rst), .Q(sreg[136]) );
  DFF \sreg_reg[137]  ( .D(swire[73]), .CLK(clk), .RST(rst), .Q(sreg[137]) );
  DFF \sreg_reg[138]  ( .D(swire[74]), .CLK(clk), .RST(rst), .Q(sreg[138]) );
  DFF \sreg_reg[139]  ( .D(swire[75]), .CLK(clk), .RST(rst), .Q(sreg[139]) );
  DFF \sreg_reg[140]  ( .D(swire[76]), .CLK(clk), .RST(rst), .Q(sreg[140]) );
  DFF \sreg_reg[141]  ( .D(swire[77]), .CLK(clk), .RST(rst), .Q(sreg[141]) );
  DFF \sreg_reg[142]  ( .D(swire[78]), .CLK(clk), .RST(rst), .Q(sreg[142]) );
  DFF \sreg_reg[143]  ( .D(swire[79]), .CLK(clk), .RST(rst), .Q(sreg[143]) );
  DFF \sreg_reg[144]  ( .D(swire[80]), .CLK(clk), .RST(rst), .Q(sreg[144]) );
  DFF \sreg_reg[145]  ( .D(swire[81]), .CLK(clk), .RST(rst), .Q(sreg[145]) );
  DFF \sreg_reg[146]  ( .D(swire[82]), .CLK(clk), .RST(rst), .Q(sreg[146]) );
  DFF \sreg_reg[147]  ( .D(swire[83]), .CLK(clk), .RST(rst), .Q(sreg[147]) );
  DFF \sreg_reg[148]  ( .D(swire[84]), .CLK(clk), .RST(rst), .Q(sreg[148]) );
  DFF \sreg_reg[149]  ( .D(swire[85]), .CLK(clk), .RST(rst), .Q(sreg[149]) );
  DFF \sreg_reg[150]  ( .D(swire[86]), .CLK(clk), .RST(rst), .Q(sreg[150]) );
  DFF \sreg_reg[151]  ( .D(swire[87]), .CLK(clk), .RST(rst), .Q(sreg[151]) );
  DFF \sreg_reg[152]  ( .D(swire[88]), .CLK(clk), .RST(rst), .Q(sreg[152]) );
  DFF \sreg_reg[153]  ( .D(swire[89]), .CLK(clk), .RST(rst), .Q(sreg[153]) );
  DFF \sreg_reg[154]  ( .D(swire[90]), .CLK(clk), .RST(rst), .Q(sreg[154]) );
  DFF \sreg_reg[155]  ( .D(swire[91]), .CLK(clk), .RST(rst), .Q(sreg[155]) );
  DFF \sreg_reg[156]  ( .D(swire[92]), .CLK(clk), .RST(rst), .Q(sreg[156]) );
  DFF \sreg_reg[157]  ( .D(swire[93]), .CLK(clk), .RST(rst), .Q(sreg[157]) );
  DFF \sreg_reg[158]  ( .D(swire[94]), .CLK(clk), .RST(rst), .Q(sreg[158]) );
  DFF \sreg_reg[159]  ( .D(swire[95]), .CLK(clk), .RST(rst), .Q(sreg[159]) );
  DFF \sreg_reg[160]  ( .D(swire[96]), .CLK(clk), .RST(rst), .Q(sreg[160]) );
  DFF \sreg_reg[161]  ( .D(swire[97]), .CLK(clk), .RST(rst), .Q(sreg[161]) );
  DFF \sreg_reg[162]  ( .D(swire[98]), .CLK(clk), .RST(rst), .Q(sreg[162]) );
  DFF \sreg_reg[163]  ( .D(swire[99]), .CLK(clk), .RST(rst), .Q(sreg[163]) );
  DFF \sreg_reg[164]  ( .D(swire[100]), .CLK(clk), .RST(rst), .Q(sreg[164]) );
  DFF \sreg_reg[165]  ( .D(swire[101]), .CLK(clk), .RST(rst), .Q(sreg[165]) );
  DFF \sreg_reg[166]  ( .D(swire[102]), .CLK(clk), .RST(rst), .Q(sreg[166]) );
  DFF \sreg_reg[167]  ( .D(swire[103]), .CLK(clk), .RST(rst), .Q(sreg[167]) );
  DFF \sreg_reg[168]  ( .D(swire[104]), .CLK(clk), .RST(rst), .Q(sreg[168]) );
  DFF \sreg_reg[169]  ( .D(swire[105]), .CLK(clk), .RST(rst), .Q(sreg[169]) );
  DFF \sreg_reg[170]  ( .D(swire[106]), .CLK(clk), .RST(rst), .Q(sreg[170]) );
  DFF \sreg_reg[171]  ( .D(swire[107]), .CLK(clk), .RST(rst), .Q(sreg[171]) );
  DFF \sreg_reg[172]  ( .D(swire[108]), .CLK(clk), .RST(rst), .Q(sreg[172]) );
  DFF \sreg_reg[173]  ( .D(swire[109]), .CLK(clk), .RST(rst), .Q(sreg[173]) );
  DFF \sreg_reg[174]  ( .D(swire[110]), .CLK(clk), .RST(rst), .Q(sreg[174]) );
  DFF \sreg_reg[175]  ( .D(swire[111]), .CLK(clk), .RST(rst), .Q(sreg[175]) );
  DFF \sreg_reg[176]  ( .D(swire[112]), .CLK(clk), .RST(rst), .Q(sreg[176]) );
  DFF \sreg_reg[177]  ( .D(swire[113]), .CLK(clk), .RST(rst), .Q(sreg[177]) );
  DFF \sreg_reg[178]  ( .D(swire[114]), .CLK(clk), .RST(rst), .Q(sreg[178]) );
  DFF \sreg_reg[179]  ( .D(swire[115]), .CLK(clk), .RST(rst), .Q(sreg[179]) );
  DFF \sreg_reg[180]  ( .D(swire[116]), .CLK(clk), .RST(rst), .Q(sreg[180]) );
  DFF \sreg_reg[181]  ( .D(swire[117]), .CLK(clk), .RST(rst), .Q(sreg[181]) );
  DFF \sreg_reg[182]  ( .D(swire[118]), .CLK(clk), .RST(rst), .Q(sreg[182]) );
  DFF \sreg_reg[183]  ( .D(swire[119]), .CLK(clk), .RST(rst), .Q(sreg[183]) );
  DFF \sreg_reg[184]  ( .D(swire[120]), .CLK(clk), .RST(rst), .Q(sreg[184]) );
  DFF \sreg_reg[185]  ( .D(swire[121]), .CLK(clk), .RST(rst), .Q(sreg[185]) );
  DFF \sreg_reg[186]  ( .D(swire[122]), .CLK(clk), .RST(rst), .Q(sreg[186]) );
  DFF \sreg_reg[187]  ( .D(swire[123]), .CLK(clk), .RST(rst), .Q(sreg[187]) );
  DFF \sreg_reg[188]  ( .D(swire[124]), .CLK(clk), .RST(rst), .Q(sreg[188]) );
  DFF \sreg_reg[189]  ( .D(swire[125]), .CLK(clk), .RST(rst), .Q(sreg[189]) );
  DFF \sreg_reg[190]  ( .D(swire[126]), .CLK(clk), .RST(rst), .Q(sreg[190]) );
  DFF \sreg_reg[191]  ( .D(swire[127]), .CLK(clk), .RST(rst), .Q(sreg[191]) );
  DFF \sreg_reg[127]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[126]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[125]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[124]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[123]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[122]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[121]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[120]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[119]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[118]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[117]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[116]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[115]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[114]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[113]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[112]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[111]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[110]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[109]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[108]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[107]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[106]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[105]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[104]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[103]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[102]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[101]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[100]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[99]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[98]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[97]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[96]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[95]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[94]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[93]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[92]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[91]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[90]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[89]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[88]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[87]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[86]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[85]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[84]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[83]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[82]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[81]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[80]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[79]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[78]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[77]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[76]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[75]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[74]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[73]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[72]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[71]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[70]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[69]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[68]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[67]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[66]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[65]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[64]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XNOR U67 ( .A(n11705), .B(n11929), .Z(n11709) );
  XNOR U68 ( .A(n12824), .B(n13030), .Z(n12828) );
  XNOR U69 ( .A(n13943), .B(n14131), .Z(n13947) );
  XNOR U70 ( .A(n15062), .B(n15232), .Z(n15066) );
  XNOR U71 ( .A(n12123), .B(n12287), .Z(n12127) );
  XNOR U72 ( .A(n13242), .B(n13388), .Z(n13246) );
  XNOR U73 ( .A(n17300), .B(n17434), .Z(n17304) );
  XNOR U74 ( .A(n14361), .B(n14489), .Z(n14365) );
  XNOR U75 ( .A(n15480), .B(n15590), .Z(n15484) );
  XNOR U76 ( .A(n3100), .B(n3205), .Z(n3101) );
  XNOR U77 ( .A(n18802), .B(n18900), .Z(n18806) );
  XNOR U78 ( .A(n16599), .B(n16691), .Z(n16603) );
  XNOR U79 ( .A(n20647), .B(n20739), .Z(n20651) );
  XNOR U80 ( .A(n20289), .B(n20369), .Z(n20293) );
  XNOR U81 ( .A(n2375), .B(n2453), .Z(n2379) );
  XNOR U82 ( .A(n17718), .B(n17792), .Z(n17722) );
  XNOR U83 ( .A(n21766), .B(n21840), .Z(n21770) );
  XNOR U84 ( .A(n18837), .B(n18893), .Z(n18841) );
  XNOR U85 ( .A(n21786), .B(n21836), .Z(n21790) );
  XNOR U86 ( .A(n19956), .B(n19994), .Z(n19960) );
  XNOR U87 ( .A(n13460), .B(n13785), .Z(n13469) );
  XNOR U88 ( .A(n15698), .B(n15987), .Z(n15707) );
  XNOR U89 ( .A(n8191), .B(n8443), .Z(n8195) );
  XNOR U90 ( .A(n17936), .B(n18189), .Z(n17945) );
  XNOR U91 ( .A(n10969), .B(n10598), .Z(n10600) );
  XNOR U92 ( .A(n8211), .B(n8439), .Z(n8215) );
  XNOR U93 ( .A(n11715), .B(n11927), .Z(n11719) );
  XNOR U94 ( .A(n20174), .B(n20391), .Z(n20183) );
  XNOR U95 ( .A(n7101), .B(n7320), .Z(n7105) );
  XNOR U96 ( .A(n6349), .B(n6580), .Z(n6350) );
  XNOR U97 ( .A(n6378), .B(n6573), .Z(n6379) );
  XNOR U98 ( .A(n12834), .B(n13028), .Z(n12838) );
  XNOR U99 ( .A(n11740), .B(n11922), .Z(n11744) );
  XNOR U100 ( .A(n4840), .B(n5096), .Z(n4841) );
  XNOR U101 ( .A(n13953), .B(n14129), .Z(n13957) );
  XNOR U102 ( .A(n12859), .B(n13023), .Z(n12863) );
  XNOR U103 ( .A(n15072), .B(n15230), .Z(n15076) );
  XNOR U104 ( .A(n12133), .B(n12285), .Z(n12137) );
  XNOR U105 ( .A(n16549), .B(n16701), .Z(n16553) );
  XNOR U106 ( .A(n13978), .B(n14124), .Z(n13982) );
  XNOR U107 ( .A(n16191), .B(n16331), .Z(n16195) );
  XNOR U108 ( .A(n12148), .B(n12282), .Z(n12152) );
  XNOR U109 ( .A(n13252), .B(n13386), .Z(n13256) );
  XNOR U110 ( .A(n15097), .B(n15225), .Z(n15101) );
  XNOR U111 ( .A(n17310), .B(n17432), .Z(n17314) );
  XNOR U112 ( .A(n12163), .B(n12279), .Z(n12167) );
  XNOR U113 ( .A(n13267), .B(n13383), .Z(n13271) );
  XNOR U114 ( .A(n14371), .B(n14487), .Z(n14375) );
  XNOR U115 ( .A(n18787), .B(n18903), .Z(n18791) );
  XNOR U116 ( .A(n16216), .B(n16326), .Z(n16220) );
  XNOR U117 ( .A(n18429), .B(n18533), .Z(n18433) );
  XNOR U118 ( .A(n12178), .B(n12276), .Z(n12182) );
  XNOR U119 ( .A(n13282), .B(n13380), .Z(n13286) );
  XNOR U120 ( .A(n14386), .B(n14484), .Z(n14390) );
  XNOR U121 ( .A(n15490), .B(n15588), .Z(n15494) );
  XNOR U122 ( .A(n20642), .B(n20740), .Z(n20646) );
  XNOR U123 ( .A(n3107), .B(n3203), .Z(n3111) );
  XNOR U124 ( .A(n17335), .B(n17427), .Z(n17339) );
  XNOR U125 ( .A(n19548), .B(n19634), .Z(n19552) );
  XNOR U126 ( .A(n12193), .B(n12273), .Z(n12197) );
  XNOR U127 ( .A(n13297), .B(n13377), .Z(n13301) );
  XNOR U128 ( .A(n14401), .B(n14481), .Z(n14405) );
  XNOR U129 ( .A(n15505), .B(n15585), .Z(n15509) );
  XNOR U130 ( .A(n16609), .B(n16689), .Z(n16613) );
  XNOR U131 ( .A(n20657), .B(n20737), .Z(n20661) );
  XNOR U132 ( .A(n21761), .B(n21841), .Z(n21765) );
  XNOR U133 ( .A(n18454), .B(n18528), .Z(n18458) );
  XNOR U134 ( .A(n1998), .B(n2082), .Z(n2002) );
  XNOR U135 ( .A(n20299), .B(n20367), .Z(n20303) );
  XNOR U136 ( .A(n12208), .B(n12270), .Z(n12212) );
  XNOR U137 ( .A(n13312), .B(n13374), .Z(n13316) );
  XNOR U138 ( .A(n14416), .B(n14478), .Z(n14420) );
  XNOR U139 ( .A(n15520), .B(n15582), .Z(n15524) );
  XNOR U140 ( .A(n16624), .B(n16686), .Z(n16628) );
  XNOR U141 ( .A(n17728), .B(n17790), .Z(n17732) );
  XNOR U142 ( .A(n22144), .B(n22206), .Z(n22148) );
  XNOR U143 ( .A(n19941), .B(n19997), .Z(n19945) );
  XNOR U144 ( .A(n21781), .B(n21837), .Z(n21785) );
  XNOR U145 ( .A(n12223), .B(n12267), .Z(n12227) );
  XNOR U146 ( .A(n13327), .B(n13371), .Z(n13331) );
  XNOR U147 ( .A(n14431), .B(n14475), .Z(n14435) );
  XNOR U148 ( .A(n15535), .B(n15579), .Z(n15539) );
  XNOR U149 ( .A(n16639), .B(n16683), .Z(n16643) );
  XNOR U150 ( .A(n17743), .B(n17787), .Z(n17747) );
  XNOR U151 ( .A(n18847), .B(n18891), .Z(n18851) );
  XNOR U152 ( .A(n22164), .B(n22202), .Z(n22168) );
  XNOR U153 ( .A(n12238), .B(n12264), .Z(n12242) );
  XNOR U154 ( .A(n13342), .B(n13368), .Z(n13346) );
  XNOR U155 ( .A(n14446), .B(n14472), .Z(n14450) );
  XNOR U156 ( .A(n15550), .B(n15576), .Z(n15554) );
  XNOR U157 ( .A(n16654), .B(n16680), .Z(n16658) );
  XNOR U158 ( .A(n17758), .B(n17784), .Z(n17762) );
  XNOR U159 ( .A(n18862), .B(n18888), .Z(n18866) );
  XNOR U160 ( .A(n19966), .B(n19992), .Z(n19970) );
  XNOR U161 ( .A(n11968), .B(n12317), .Z(n11977) );
  XNOR U162 ( .A(n14206), .B(n14519), .Z(n14215) );
  XNOR U163 ( .A(n7769), .B(n8081), .Z(n7773) );
  XNOR U164 ( .A(n7784), .B(n8078), .Z(n7788) );
  XNOR U165 ( .A(n16444), .B(n16721), .Z(n16453) );
  XNOR U166 ( .A(n7799), .B(n8075), .Z(n7803) );
  XNOR U167 ( .A(n7819), .B(n8071), .Z(n7823) );
  XNOR U168 ( .A(n11690), .B(n11932), .Z(n11694) );
  XNOR U169 ( .A(n18682), .B(n18923), .Z(n18691) );
  XNOR U170 ( .A(n10595), .B(n10824), .Z(n10599) );
  XNOR U171 ( .A(n12073), .B(n12297), .Z(n12077) );
  XNOR U172 ( .A(n12809), .B(n13033), .Z(n12813) );
  XNOR U173 ( .A(n7839), .B(n8067), .Z(n7843) );
  XNOR U174 ( .A(n7481), .B(n7691), .Z(n7485) );
  XNOR U175 ( .A(n12088), .B(n12294), .Z(n12092) );
  XNOR U176 ( .A(n13192), .B(n13398), .Z(n13196) );
  XNOR U177 ( .A(n13928), .B(n14134), .Z(n13932) );
  XNOR U178 ( .A(n11725), .B(n11925), .Z(n11729) );
  XNOR U179 ( .A(n20920), .B(n21125), .Z(n20929) );
  XNOR U180 ( .A(n5972), .B(n6209), .Z(n5973) );
  XNOR U181 ( .A(n6755), .B(n6940), .Z(n6756) );
  XNOR U182 ( .A(n13207), .B(n13395), .Z(n13211) );
  XNOR U183 ( .A(n14311), .B(n14499), .Z(n14315) );
  XNOR U184 ( .A(n15047), .B(n15235), .Z(n15051) );
  XNOR U185 ( .A(n12108), .B(n12290), .Z(n12112) );
  XNOR U186 ( .A(n12844), .B(n13026), .Z(n12848) );
  XNOR U187 ( .A(n22412), .B(n22593), .Z(n22421) );
  XNOR U188 ( .A(n14326), .B(n14496), .Z(n14330) );
  XNOR U189 ( .A(n15430), .B(n15600), .Z(n15434) );
  XNOR U190 ( .A(n16166), .B(n16336), .Z(n16170) );
  XNOR U191 ( .A(n5276), .B(n5453), .Z(n5277) );
  XNOR U192 ( .A(n4086), .B(n4353), .Z(n4087) );
  XNOR U193 ( .A(n13227), .B(n13391), .Z(n13231) );
  XNOR U194 ( .A(n13963), .B(n14127), .Z(n13967) );
  XNOR U195 ( .A(n12501), .B(n12653), .Z(n12505) );
  XNOR U196 ( .A(n15445), .B(n15597), .Z(n15449) );
  XNOR U197 ( .A(n16181), .B(n16333), .Z(n16185) );
  XNOR U198 ( .A(n16917), .B(n17069), .Z(n16921) );
  XNOR U199 ( .A(n17653), .B(n17805), .Z(n17657) );
  XNOR U200 ( .A(n2955), .B(n3240), .Z(n2956) );
  XNOR U201 ( .A(n4550), .B(n4703), .Z(n4551) );
  XNOR U202 ( .A(n14346), .B(n14492), .Z(n14350) );
  XNOR U203 ( .A(n15082), .B(n15228), .Z(n15086) );
  XNOR U204 ( .A(n5293), .B(n5449), .Z(n5301) );
  XNOR U205 ( .A(n12516), .B(n12650), .Z(n12520) );
  XNOR U206 ( .A(n13620), .B(n13754), .Z(n13624) );
  XNOR U207 ( .A(n16564), .B(n16698), .Z(n16568) );
  XNOR U208 ( .A(n17668), .B(n17802), .Z(n17672) );
  XNOR U209 ( .A(n18404), .B(n18538), .Z(n18408) );
  XNOR U210 ( .A(n15465), .B(n15593), .Z(n15469) );
  XNOR U211 ( .A(n16201), .B(n16329), .Z(n16205) );
  XNOR U212 ( .A(n3825), .B(n3954), .Z(n3826) );
  XNOR U213 ( .A(n4567), .B(n4699), .Z(n4575) );
  XNOR U214 ( .A(n12531), .B(n12647), .Z(n12535) );
  XNOR U215 ( .A(n13635), .B(n13751), .Z(n13639) );
  XNOR U216 ( .A(n14739), .B(n14855), .Z(n14743) );
  XNOR U217 ( .A(n17683), .B(n17799), .Z(n17687) );
  XNOR U218 ( .A(n18419), .B(n18535), .Z(n18423) );
  XNOR U219 ( .A(n19155), .B(n19271), .Z(n19159) );
  XNOR U220 ( .A(n19891), .B(n20007), .Z(n19895) );
  XNOR U221 ( .A(n16584), .B(n16694), .Z(n16588) );
  XNOR U222 ( .A(n17320), .B(n17430), .Z(n17324) );
  XNOR U223 ( .A(n3477), .B(n3576), .Z(n3478) );
  XNOR U224 ( .A(n12546), .B(n12644), .Z(n12550) );
  XNOR U225 ( .A(n13650), .B(n13748), .Z(n13654) );
  XNOR U226 ( .A(n14754), .B(n14852), .Z(n14758) );
  XNOR U227 ( .A(n15858), .B(n15956), .Z(n15862) );
  XNOR U228 ( .A(n19170), .B(n19268), .Z(n19174) );
  XNOR U229 ( .A(n19906), .B(n20004), .Z(n19910) );
  XNOR U230 ( .A(n21010), .B(n21108), .Z(n21014) );
  XNOR U231 ( .A(n17703), .B(n17795), .Z(n17707) );
  XNOR U232 ( .A(n18439), .B(n18531), .Z(n18443) );
  XNOR U233 ( .A(n3117), .B(n3201), .Z(n3125) );
  XNOR U234 ( .A(n12561), .B(n12641), .Z(n12565) );
  XNOR U235 ( .A(n13665), .B(n13745), .Z(n13669) );
  XNOR U236 ( .A(n14769), .B(n14849), .Z(n14773) );
  XNOR U237 ( .A(n15873), .B(n15953), .Z(n15877) );
  XNOR U238 ( .A(n16977), .B(n17057), .Z(n16981) );
  XNOR U239 ( .A(n21025), .B(n21105), .Z(n21029) );
  XNOR U240 ( .A(n18822), .B(n18896), .Z(n18826) );
  XNOR U241 ( .A(n19558), .B(n19632), .Z(n19562) );
  XNOR U242 ( .A(n20294), .B(n20368), .Z(n20298) );
  XNOR U243 ( .A(n22134), .B(n22208), .Z(n22138) );
  XNOR U244 ( .A(n2380), .B(n2452), .Z(n2384) );
  XNOR U245 ( .A(n1264), .B(n1336), .Z(n1268) );
  XNOR U246 ( .A(n12576), .B(n12638), .Z(n12580) );
  XNOR U247 ( .A(n13680), .B(n13742), .Z(n13684) );
  XNOR U248 ( .A(n14784), .B(n14846), .Z(n14788) );
  XNOR U249 ( .A(n15888), .B(n15950), .Z(n15892) );
  XNOR U250 ( .A(n16992), .B(n17054), .Z(n16996) );
  XNOR U251 ( .A(n18096), .B(n18158), .Z(n18100) );
  XNOR U252 ( .A(n21408), .B(n21470), .Z(n21412) );
  XNOR U253 ( .A(n19573), .B(n19629), .Z(n19577) );
  XNOR U254 ( .A(n20309), .B(n20365), .Z(n20313) );
  XNOR U255 ( .A(n21045), .B(n21101), .Z(n21049) );
  XNOR U256 ( .A(n22149), .B(n22205), .Z(n22153) );
  XNOR U257 ( .A(n12591), .B(n12635), .Z(n12595) );
  XNOR U258 ( .A(n13695), .B(n13739), .Z(n13699) );
  XNOR U259 ( .A(n14799), .B(n14843), .Z(n14803) );
  XNOR U260 ( .A(n15903), .B(n15947), .Z(n15907) );
  XNOR U261 ( .A(n17007), .B(n17051), .Z(n17011) );
  XNOR U262 ( .A(n18111), .B(n18155), .Z(n18115) );
  XNOR U263 ( .A(n19215), .B(n19259), .Z(n19219) );
  XNOR U264 ( .A(n917), .B(n959), .Z(n921) );
  XNOR U265 ( .A(n1661), .B(n1703), .Z(n1665) );
  XNOR U266 ( .A(n22532), .B(n22570), .Z(n22536) );
  XNOR U267 ( .A(n10235), .B(n10372), .Z(n10229) );
  XNOR U268 ( .A(n21433), .B(n21465), .Z(n21437) );
  XNOR U269 ( .A(n12606), .B(n12632), .Z(n12610) );
  XNOR U270 ( .A(n13710), .B(n13736), .Z(n13714) );
  XNOR U271 ( .A(n14814), .B(n14840), .Z(n14818) );
  XNOR U272 ( .A(n15918), .B(n15944), .Z(n15922) );
  XNOR U273 ( .A(n17022), .B(n17048), .Z(n17026) );
  XNOR U274 ( .A(n18126), .B(n18152), .Z(n18130) );
  XNOR U275 ( .A(n19230), .B(n19256), .Z(n19234) );
  XNOR U276 ( .A(n20334), .B(n20360), .Z(n20338) );
  XNOR U277 ( .A(n21070), .B(n21096), .Z(n21074) );
  XNOR U278 ( .A(n22174), .B(n22200), .Z(n22178) );
  AND U279 ( .A(n63), .B(n64), .Z(n61) );
  XNOR U280 ( .A(n15643), .B(n16000), .Z(n15648) );
  XNOR U281 ( .A(n20059), .B(n20416), .Z(n20064) );
  XNOR U282 ( .A(n10495), .B(n10844), .Z(n10499) );
  XNOR U283 ( .A(n11231), .B(n11582), .Z(n11236) );
  XNOR U284 ( .A(n12705), .B(n13055), .Z(n12709) );
  XNOR U285 ( .A(n17121), .B(n17471), .Z(n17125) );
  XNOR U286 ( .A(n21537), .B(n21887), .Z(n21541) );
  XNOR U287 ( .A(n8111), .B(n8459), .Z(n8115) );
  XNOR U288 ( .A(n14182), .B(n14526), .Z(n14186) );
  XNOR U289 ( .A(n18598), .B(n18942), .Z(n18602) );
  XNOR U290 ( .A(n15659), .B(n15997), .Z(n15663) );
  XNOR U291 ( .A(n20075), .B(n20413), .Z(n20079) );
  XNOR U292 ( .A(n10878), .B(n11210), .Z(n10882) );
  XNOR U293 ( .A(n11615), .B(n11947), .Z(n11619) );
  XNOR U294 ( .A(n12351), .B(n12683), .Z(n12355) );
  XNOR U295 ( .A(n17136), .B(n17468), .Z(n17140) );
  XNOR U296 ( .A(n21552), .B(n21884), .Z(n21556) );
  XNOR U297 ( .A(n8126), .B(n8456), .Z(n8130) );
  XNOR U298 ( .A(n14197), .B(n14523), .Z(n14201) );
  XNOR U299 ( .A(n18613), .B(n18939), .Z(n18617) );
  XNOR U300 ( .A(n15674), .B(n15994), .Z(n15678) );
  XNOR U301 ( .A(n20090), .B(n20410), .Z(n20094) );
  XNOR U302 ( .A(n7759), .B(n8083), .Z(n7763) );
  XNOR U303 ( .A(n6992), .B(n7343), .Z(n6996) );
  XNOR U304 ( .A(n10525), .B(n10838), .Z(n10529) );
  XNOR U305 ( .A(n11262), .B(n11576), .Z(n11266) );
  XNOR U306 ( .A(n11998), .B(n12312), .Z(n12002) );
  XNOR U307 ( .A(n12734), .B(n13048), .Z(n12738) );
  XNOR U308 ( .A(n13470), .B(n13784), .Z(n13474) );
  XNOR U309 ( .A(n17151), .B(n17465), .Z(n17155) );
  XNOR U310 ( .A(n21567), .B(n21881), .Z(n21571) );
  XNOR U311 ( .A(n18628), .B(n18936), .Z(n18632) );
  XNOR U312 ( .A(n15689), .B(n15991), .Z(n15693) );
  XNOR U313 ( .A(n20105), .B(n20407), .Z(n20109) );
  XNOR U314 ( .A(n8151), .B(n8451), .Z(n8155) );
  XNOR U315 ( .A(n10908), .B(n11204), .Z(n10912) );
  XNOR U316 ( .A(n11645), .B(n11941), .Z(n11649) );
  XNOR U317 ( .A(n12381), .B(n12677), .Z(n12385) );
  XNOR U318 ( .A(n13117), .B(n13413), .Z(n13121) );
  XNOR U319 ( .A(n13853), .B(n14149), .Z(n13857) );
  XNOR U320 ( .A(n14589), .B(n14885), .Z(n14593) );
  XNOR U321 ( .A(n17166), .B(n17462), .Z(n17170) );
  XNOR U322 ( .A(n21582), .B(n21878), .Z(n21586) );
  XNOR U323 ( .A(n18643), .B(n18933), .Z(n18647) );
  XNOR U324 ( .A(n7017), .B(n7338), .Z(n7021) );
  XNOR U325 ( .A(n10924), .B(n10553), .Z(n10555) );
  XNOR U326 ( .A(n20120), .B(n20404), .Z(n20124) );
  XNOR U327 ( .A(n7789), .B(n8077), .Z(n7793) );
  XNOR U328 ( .A(n11292), .B(n11570), .Z(n11296) );
  XNOR U329 ( .A(n12028), .B(n12306), .Z(n12032) );
  XNOR U330 ( .A(n12764), .B(n13042), .Z(n12768) );
  XNOR U331 ( .A(n13500), .B(n13778), .Z(n13504) );
  XNOR U332 ( .A(n14236), .B(n14514), .Z(n14240) );
  XNOR U333 ( .A(n14972), .B(n15250), .Z(n14976) );
  XNOR U334 ( .A(n15708), .B(n15986), .Z(n15712) );
  XNOR U335 ( .A(n17181), .B(n17459), .Z(n17185) );
  XNOR U336 ( .A(n21597), .B(n21875), .Z(n21601) );
  XNOR U337 ( .A(n18658), .B(n18930), .Z(n18662) );
  XNOR U338 ( .A(n8176), .B(n8446), .Z(n8180) );
  XNOR U339 ( .A(n10939), .B(n10568), .Z(n10570) );
  XNOR U340 ( .A(n11308), .B(n10936), .Z(n10938) );
  XNOR U341 ( .A(n20135), .B(n20401), .Z(n20139) );
  XNOR U342 ( .A(n11675), .B(n11935), .Z(n11679) );
  XNOR U343 ( .A(n12411), .B(n12671), .Z(n12415) );
  XNOR U344 ( .A(n13147), .B(n13407), .Z(n13151) );
  XNOR U345 ( .A(n13883), .B(n14143), .Z(n13887) );
  XNOR U346 ( .A(n14619), .B(n14879), .Z(n14623) );
  XNOR U347 ( .A(n15355), .B(n15615), .Z(n15359) );
  XNOR U348 ( .A(n16091), .B(n16351), .Z(n16095) );
  XNOR U349 ( .A(n16827), .B(n17087), .Z(n16831) );
  XNOR U350 ( .A(n21612), .B(n21872), .Z(n21616) );
  XNOR U351 ( .A(n6282), .B(n6594), .Z(n6286) );
  XNOR U352 ( .A(n18673), .B(n18927), .Z(n18677) );
  XNOR U353 ( .A(n10954), .B(n10583), .Z(n10585) );
  XNOR U354 ( .A(n20150), .B(n20398), .Z(n20154) );
  XNOR U355 ( .A(n7437), .B(n7701), .Z(n7441) );
  XNOR U356 ( .A(n11322), .B(n11564), .Z(n11326) );
  XNOR U357 ( .A(n12058), .B(n12300), .Z(n12062) );
  XNOR U358 ( .A(n12794), .B(n13036), .Z(n12798) );
  XNOR U359 ( .A(n13530), .B(n13772), .Z(n13534) );
  XNOR U360 ( .A(n14266), .B(n14508), .Z(n14270) );
  XNOR U361 ( .A(n15002), .B(n15244), .Z(n15006) );
  XNOR U362 ( .A(n15738), .B(n15980), .Z(n15742) );
  XNOR U363 ( .A(n16474), .B(n16716), .Z(n16478) );
  XNOR U364 ( .A(n17210), .B(n17452), .Z(n17214) );
  XNOR U365 ( .A(n17946), .B(n18188), .Z(n17950) );
  XNOR U366 ( .A(n21627), .B(n21869), .Z(n21631) );
  XNOR U367 ( .A(n20165), .B(n20395), .Z(n20169) );
  XNOR U368 ( .A(n7452), .B(n7698), .Z(n7456) );
  XNOR U369 ( .A(n6307), .B(n6589), .Z(n6311) );
  XNOR U370 ( .A(n12447), .B(n12076), .Z(n12078) );
  XNOR U371 ( .A(n12441), .B(n12665), .Z(n12445) );
  XNOR U372 ( .A(n13177), .B(n13401), .Z(n13181) );
  XNOR U373 ( .A(n13913), .B(n14137), .Z(n13917) );
  XNOR U374 ( .A(n14649), .B(n14873), .Z(n14653) );
  XNOR U375 ( .A(n15385), .B(n15609), .Z(n15389) );
  XNOR U376 ( .A(n16121), .B(n16345), .Z(n16125) );
  XNOR U377 ( .A(n16857), .B(n17081), .Z(n16861) );
  XNOR U378 ( .A(n17593), .B(n17817), .Z(n17597) );
  XNOR U379 ( .A(n18329), .B(n18553), .Z(n18333) );
  XNOR U380 ( .A(n19065), .B(n19289), .Z(n19069) );
  XNOR U381 ( .A(n21642), .B(n21866), .Z(n21646) );
  XNOR U382 ( .A(n10973), .B(n11191), .Z(n10977) );
  XNOR U383 ( .A(n7479), .B(n7692), .Z(n7480) );
  XNOR U384 ( .A(n8221), .B(n8437), .Z(n8229) );
  XNOR U385 ( .A(n12456), .B(n12662), .Z(n12460) );
  XNOR U386 ( .A(n13566), .B(n13195), .Z(n13197) );
  XNOR U387 ( .A(n13560), .B(n13766), .Z(n13564) );
  XNOR U388 ( .A(n14296), .B(n14502), .Z(n14300) );
  XNOR U389 ( .A(n15032), .B(n15238), .Z(n15036) );
  XNOR U390 ( .A(n15768), .B(n15974), .Z(n15772) );
  XNOR U391 ( .A(n16504), .B(n16710), .Z(n16508) );
  XNOR U392 ( .A(n17240), .B(n17446), .Z(n17244) );
  XNOR U393 ( .A(n17976), .B(n18182), .Z(n17980) );
  XNOR U394 ( .A(n18712), .B(n18918), .Z(n18716) );
  XNOR U395 ( .A(n19448), .B(n19654), .Z(n19452) );
  XNOR U396 ( .A(n20184), .B(n20390), .Z(n20188) );
  XNOR U397 ( .A(n21657), .B(n21863), .Z(n21661) );
  XNOR U398 ( .A(n7106), .B(n7319), .Z(n7110) );
  XNOR U399 ( .A(n10620), .B(n10819), .Z(n10624) );
  XNOR U400 ( .A(n12093), .B(n12293), .Z(n12097) );
  XNOR U401 ( .A(n10999), .B(n10628), .Z(n10630) );
  XNOR U402 ( .A(n5974), .B(n6208), .Z(n5978) );
  XNOR U403 ( .A(n3662), .B(n3992), .Z(n3666) );
  XNOR U404 ( .A(n7496), .B(n7688), .Z(n7504) );
  XNOR U405 ( .A(n13575), .B(n13763), .Z(n13579) );
  XNOR U406 ( .A(n14685), .B(n14314), .Z(n14316) );
  XNOR U407 ( .A(n14679), .B(n14867), .Z(n14683) );
  XNOR U408 ( .A(n15415), .B(n15603), .Z(n15419) );
  XNOR U409 ( .A(n16151), .B(n16339), .Z(n16155) );
  XNOR U410 ( .A(n16887), .B(n17075), .Z(n16891) );
  XNOR U411 ( .A(n17623), .B(n17811), .Z(n17627) );
  XNOR U412 ( .A(n18359), .B(n18547), .Z(n18363) );
  XNOR U413 ( .A(n19095), .B(n19283), .Z(n19099) );
  XNOR U414 ( .A(n19831), .B(n20019), .Z(n19835) );
  XNOR U415 ( .A(n20567), .B(n20755), .Z(n20571) );
  XNOR U416 ( .A(n21303), .B(n21491), .Z(n21307) );
  XNOR U417 ( .A(n6385), .B(n6571), .Z(n6389) );
  XNOR U418 ( .A(n7128), .B(n7314), .Z(n7129) );
  XNOR U419 ( .A(n11009), .B(n10638), .Z(n10640) );
  XNOR U420 ( .A(n12482), .B(n12111), .Z(n12113) );
  XNOR U421 ( .A(n12476), .B(n12658), .Z(n12480) );
  XNOR U422 ( .A(n13212), .B(n13394), .Z(n13216) );
  XNOR U423 ( .A(n5201), .B(n5471), .Z(n5205) );
  XNOR U424 ( .A(n11014), .B(n10643), .Z(n10645) );
  XNOR U425 ( .A(n4842), .B(n5095), .Z(n4846) );
  XNOR U426 ( .A(n4059), .B(n4359), .Z(n4063) );
  XNOR U427 ( .A(n4869), .B(n5089), .Z(n4870) );
  XNOR U428 ( .A(n9742), .B(n9920), .Z(n9746) );
  XNOR U429 ( .A(n14694), .B(n14864), .Z(n14698) );
  XNOR U430 ( .A(n15804), .B(n15433), .Z(n15435) );
  XNOR U431 ( .A(n15798), .B(n15968), .Z(n15802) );
  XNOR U432 ( .A(n16534), .B(n16704), .Z(n16538) );
  XNOR U433 ( .A(n17270), .B(n17440), .Z(n17274) );
  XNOR U434 ( .A(n18006), .B(n18176), .Z(n18010) );
  XNOR U435 ( .A(n18742), .B(n18912), .Z(n18746) );
  XNOR U436 ( .A(n19478), .B(n19648), .Z(n19482) );
  XNOR U437 ( .A(n20214), .B(n20384), .Z(n20218) );
  XNOR U438 ( .A(n20950), .B(n21120), .Z(n20954) );
  XNOR U439 ( .A(n21686), .B(n21856), .Z(n21690) );
  XNOR U440 ( .A(n22422), .B(n22592), .Z(n22426) );
  XNOR U441 ( .A(n5636), .B(n5828), .Z(n5640) );
  XNOR U442 ( .A(n6404), .B(n6568), .Z(n6399) );
  XNOR U443 ( .A(n11755), .B(n11919), .Z(n11759) );
  XNOR U444 ( .A(n12491), .B(n12655), .Z(n12495) );
  XNOR U445 ( .A(n13601), .B(n13230), .Z(n13232) );
  XNOR U446 ( .A(n13595), .B(n13759), .Z(n13599) );
  XNOR U447 ( .A(n14331), .B(n14495), .Z(n14335) );
  XNOR U448 ( .A(n4898), .B(n5082), .Z(n4899) );
  XNOR U449 ( .A(n3709), .B(n3982), .Z(n3710) );
  XNOR U450 ( .A(n6032), .B(n6194), .Z(n6036) );
  XNOR U451 ( .A(n11029), .B(n10658), .Z(n10660) );
  XNOR U452 ( .A(n5283), .B(n5451), .Z(n5287) );
  XNOR U453 ( .A(n3310), .B(n3616), .Z(n3314) );
  XNOR U454 ( .A(n3738), .B(n3975), .Z(n3739) );
  XNOR U455 ( .A(n11771), .B(n11400), .Z(n11402) );
  XNOR U456 ( .A(n15813), .B(n15965), .Z(n15817) );
  XNOR U457 ( .A(n16923), .B(n16552), .Z(n16554) );
  XNOR U458 ( .A(n17285), .B(n17437), .Z(n17289) );
  XNOR U459 ( .A(n18021), .B(n18173), .Z(n18025) );
  XNOR U460 ( .A(n18757), .B(n18909), .Z(n18761) );
  XNOR U461 ( .A(n19493), .B(n19645), .Z(n19497) );
  XNOR U462 ( .A(n20229), .B(n20381), .Z(n20233) );
  XNOR U463 ( .A(n20965), .B(n21117), .Z(n20969) );
  XNOR U464 ( .A(n21701), .B(n21853), .Z(n21705) );
  XNOR U465 ( .A(n22437), .B(n22589), .Z(n22441) );
  XNOR U466 ( .A(n4504), .B(n4714), .Z(n4508) );
  XNOR U467 ( .A(n5670), .B(n5820), .Z(n5678) );
  XNOR U468 ( .A(n11039), .B(n10668), .Z(n10670) );
  XNOR U469 ( .A(n12138), .B(n12284), .Z(n12142) );
  XNOR U470 ( .A(n12874), .B(n13020), .Z(n12878) );
  XNOR U471 ( .A(n13610), .B(n13756), .Z(n13614) );
  XNOR U472 ( .A(n14720), .B(n14349), .Z(n14351) );
  XNOR U473 ( .A(n14714), .B(n14860), .Z(n14718) );
  XNOR U474 ( .A(n15450), .B(n15596), .Z(n15454) );
  XNOR U475 ( .A(n3767), .B(n3968), .Z(n3768) );
  XNOR U476 ( .A(n2577), .B(n2869), .Z(n2578) );
  XNOR U477 ( .A(n5305), .B(n5446), .Z(n5306) );
  XNOR U478 ( .A(n6791), .B(n6931), .Z(n6795) );
  XNOR U479 ( .A(n11044), .B(n10673), .Z(n10675) );
  XNOR U480 ( .A(n4533), .B(n4707), .Z(n4537) );
  XNOR U481 ( .A(n3344), .B(n3608), .Z(n3348) );
  XNOR U482 ( .A(n2606), .B(n2862), .Z(n2607) );
  XNOR U483 ( .A(n3796), .B(n3961), .Z(n3797) );
  XNOR U484 ( .A(n9771), .B(n9912), .Z(n9775) );
  XNOR U485 ( .A(n16932), .B(n17066), .Z(n16936) );
  XNOR U486 ( .A(n18042), .B(n17671), .Z(n17673) );
  XNOR U487 ( .A(n18036), .B(n18170), .Z(n18040) );
  XNOR U488 ( .A(n18772), .B(n18906), .Z(n18776) );
  XNOR U489 ( .A(n19508), .B(n19642), .Z(n19512) );
  XNOR U490 ( .A(n20244), .B(n20378), .Z(n20248) );
  XNOR U491 ( .A(n20980), .B(n21114), .Z(n20984) );
  XNOR U492 ( .A(n21716), .B(n21850), .Z(n21720) );
  XNOR U493 ( .A(n22452), .B(n22586), .Z(n22456) );
  XNOR U494 ( .A(n3373), .B(n3601), .Z(n3377) );
  XNOR U495 ( .A(n11785), .B(n11913), .Z(n11789) );
  XNOR U496 ( .A(n12521), .B(n12649), .Z(n12525) );
  XNOR U497 ( .A(n13257), .B(n13385), .Z(n13261) );
  XNOR U498 ( .A(n13993), .B(n14121), .Z(n13997) );
  XNOR U499 ( .A(n14729), .B(n14857), .Z(n14733) );
  XNOR U500 ( .A(n15839), .B(n15468), .Z(n15470) );
  XNOR U501 ( .A(n15833), .B(n15961), .Z(n15837) );
  XNOR U502 ( .A(n16569), .B(n16697), .Z(n16573) );
  XNOR U503 ( .A(n2635), .B(n2855), .Z(n2636) );
  XNOR U504 ( .A(n1445), .B(n1754), .Z(n1446) );
  XNOR U505 ( .A(n4202), .B(n4325), .Z(n4203) );
  XNOR U506 ( .A(n6061), .B(n6187), .Z(n6065) );
  XNOR U507 ( .A(n7549), .B(n7675), .Z(n7553) );
  XNOR U508 ( .A(n11059), .B(n10688), .Z(n10690) );
  XNOR U509 ( .A(n3402), .B(n3594), .Z(n3406) );
  XNOR U510 ( .A(n2211), .B(n2494), .Z(n2215) );
  XNOR U511 ( .A(n1474), .B(n1747), .Z(n1475) );
  XNOR U512 ( .A(n2664), .B(n2848), .Z(n2665) );
  XNOR U513 ( .A(n4953), .B(n5070), .Z(n4948) );
  XNOR U514 ( .A(n11801), .B(n11430), .Z(n11432) );
  XNOR U515 ( .A(n18051), .B(n18167), .Z(n18055) );
  XNOR U516 ( .A(n19161), .B(n18790), .Z(n18792) );
  XNOR U517 ( .A(n19523), .B(n19639), .Z(n19527) );
  XNOR U518 ( .A(n20259), .B(n20375), .Z(n20263) );
  XNOR U519 ( .A(n20995), .B(n21111), .Z(n20999) );
  XNOR U520 ( .A(n21731), .B(n21847), .Z(n21735) );
  XNOR U521 ( .A(n22467), .B(n22583), .Z(n22471) );
  XNOR U522 ( .A(n2240), .B(n2487), .Z(n2244) );
  XNOR U523 ( .A(n3431), .B(n3587), .Z(n3435) );
  XNOR U524 ( .A(n11069), .B(n10698), .Z(n10700) );
  XNOR U525 ( .A(n12168), .B(n12278), .Z(n12172) );
  XNOR U526 ( .A(n12904), .B(n13014), .Z(n12908) );
  XNOR U527 ( .A(n13640), .B(n13750), .Z(n13644) );
  XNOR U528 ( .A(n14376), .B(n14486), .Z(n14380) );
  XNOR U529 ( .A(n15112), .B(n15222), .Z(n15116) );
  XNOR U530 ( .A(n15848), .B(n15958), .Z(n15852) );
  XNOR U531 ( .A(n16958), .B(n16587), .Z(n16589) );
  XNOR U532 ( .A(n16952), .B(n17062), .Z(n16956) );
  XNOR U533 ( .A(n17688), .B(n17798), .Z(n17692) );
  XNOR U534 ( .A(n2693), .B(n2841), .Z(n2694) );
  XNOR U535 ( .A(n1503), .B(n1740), .Z(n1504) );
  XNOR U536 ( .A(n6820), .B(n6924), .Z(n6824) );
  XNOR U537 ( .A(n8308), .B(n8416), .Z(n8316) );
  XNOR U538 ( .A(n11074), .B(n10703), .Z(n10705) );
  XNOR U539 ( .A(n3460), .B(n3580), .Z(n3464) );
  XNOR U540 ( .A(n2269), .B(n2480), .Z(n2273) );
  XNOR U541 ( .A(n1532), .B(n1733), .Z(n1533) );
  XNOR U542 ( .A(n2722), .B(n2834), .Z(n2723) );
  XNOR U543 ( .A(n9800), .B(n9904), .Z(n9804) );
  XNOR U544 ( .A(n19538), .B(n19636), .Z(n19542) );
  XNOR U545 ( .A(n20274), .B(n20372), .Z(n20278) );
  XNOR U546 ( .A(n21746), .B(n21844), .Z(n21750) );
  XNOR U547 ( .A(n22482), .B(n22580), .Z(n22486) );
  XNOR U548 ( .A(n2298), .B(n2473), .Z(n2302) );
  XNOR U549 ( .A(n3479), .B(n3575), .Z(n3483) );
  XNOR U550 ( .A(n4228), .B(n4320), .Z(n4223) );
  XNOR U551 ( .A(n11815), .B(n11907), .Z(n11819) );
  XNOR U552 ( .A(n12551), .B(n12643), .Z(n12555) );
  XNOR U553 ( .A(n13287), .B(n13379), .Z(n13291) );
  XNOR U554 ( .A(n14023), .B(n14115), .Z(n14027) );
  XNOR U555 ( .A(n14759), .B(n14851), .Z(n14763) );
  XNOR U556 ( .A(n15495), .B(n15587), .Z(n15499) );
  XNOR U557 ( .A(n16231), .B(n16323), .Z(n16235) );
  XNOR U558 ( .A(n16967), .B(n17059), .Z(n16971) );
  XNOR U559 ( .A(n18077), .B(n17706), .Z(n17708) );
  XNOR U560 ( .A(n18071), .B(n18163), .Z(n18075) );
  XNOR U561 ( .A(n18807), .B(n18899), .Z(n18811) );
  XNOR U562 ( .A(n21015), .B(n21107), .Z(n21019) );
  XNOR U563 ( .A(n1561), .B(n1726), .Z(n1562) );
  XNOR U564 ( .A(n7578), .B(n7668), .Z(n7582) );
  XNOR U565 ( .A(n9071), .B(n9153), .Z(n9066) );
  XNOR U566 ( .A(n11089), .B(n10718), .Z(n10720) );
  XNOR U567 ( .A(n2327), .B(n2466), .Z(n2331) );
  XNOR U568 ( .A(n1590), .B(n1719), .Z(n1591) );
  XNOR U569 ( .A(n11831), .B(n11460), .Z(n11462) );
  XNOR U570 ( .A(n22497), .B(n22577), .Z(n22501) );
  XNOR U571 ( .A(n2356), .B(n2459), .Z(n2360) );
  XNOR U572 ( .A(n3126), .B(n3200), .Z(n3121) );
  XNOR U573 ( .A(n11099), .B(n10728), .Z(n10730) );
  XNOR U574 ( .A(n12198), .B(n12272), .Z(n12202) );
  XNOR U575 ( .A(n12934), .B(n13008), .Z(n12938) );
  XNOR U576 ( .A(n13670), .B(n13744), .Z(n13674) );
  XNOR U577 ( .A(n14406), .B(n14480), .Z(n14410) );
  XNOR U578 ( .A(n15142), .B(n15216), .Z(n15146) );
  XNOR U579 ( .A(n15878), .B(n15952), .Z(n15882) );
  XNOR U580 ( .A(n16614), .B(n16688), .Z(n16618) );
  XNOR U581 ( .A(n17350), .B(n17424), .Z(n17354) );
  XNOR U582 ( .A(n18086), .B(n18160), .Z(n18090) );
  XNOR U583 ( .A(n19196), .B(n18825), .Z(n18827) );
  XNOR U584 ( .A(n19190), .B(n19264), .Z(n19194) );
  XNOR U585 ( .A(n19926), .B(n20000), .Z(n19930) );
  XNOR U586 ( .A(n20662), .B(n20736), .Z(n20666) );
  XNOR U587 ( .A(n21398), .B(n21472), .Z(n21402) );
  XNOR U588 ( .A(n1619), .B(n1712), .Z(n1620) );
  XNOR U589 ( .A(n11104), .B(n10733), .Z(n10735) );
  XNOR U590 ( .A(n22139), .B(n22207), .Z(n22143) );
  XNOR U591 ( .A(n1641), .B(n1707), .Z(n1645) );
  XNOR U592 ( .A(n2385), .B(n2451), .Z(n2389) );
  XNOR U593 ( .A(n3883), .B(n3940), .Z(n3884) );
  XNOR U594 ( .A(n7602), .B(n7662), .Z(n7606) );
  XNOR U595 ( .A(n11845), .B(n11901), .Z(n11849) );
  XNOR U596 ( .A(n12581), .B(n12637), .Z(n12585) );
  XNOR U597 ( .A(n13317), .B(n13373), .Z(n13321) );
  XNOR U598 ( .A(n14053), .B(n14109), .Z(n14057) );
  XNOR U599 ( .A(n14789), .B(n14845), .Z(n14793) );
  XNOR U600 ( .A(n15525), .B(n15581), .Z(n15529) );
  XNOR U601 ( .A(n16261), .B(n16317), .Z(n16265) );
  XNOR U602 ( .A(n16997), .B(n17053), .Z(n17001) );
  XNOR U603 ( .A(n17733), .B(n17789), .Z(n17737) );
  XNOR U604 ( .A(n18469), .B(n18525), .Z(n18473) );
  XNOR U605 ( .A(n19205), .B(n19261), .Z(n19209) );
  XNOR U606 ( .A(n20315), .B(n19944), .Z(n19946) );
  XNOR U607 ( .A(n20677), .B(n20733), .Z(n20681) );
  XNOR U608 ( .A(n21413), .B(n21469), .Z(n21417) );
  XNOR U609 ( .A(n1274), .B(n1334), .Z(n1278) );
  XNOR U610 ( .A(n11119), .B(n10748), .Z(n10750) );
  XNOR U611 ( .A(n22890), .B(n22940), .Z(n22894) );
  XNOR U612 ( .A(n5380), .B(n5428), .Z(n5388) );
  XNOR U613 ( .A(n6124), .B(n6172), .Z(n6128) );
  XNOR U614 ( .A(n8728), .B(n8776), .Z(n8732) );
  XNOR U615 ( .A(n11124), .B(n10753), .Z(n10755) );
  XNOR U616 ( .A(n11861), .B(n11490), .Z(n11492) );
  XNOR U617 ( .A(n22527), .B(n22571), .Z(n22531) );
  XNOR U618 ( .A(n2033), .B(n2075), .Z(n2037) );
  XNOR U619 ( .A(n2778), .B(n2821), .Z(n2782) );
  XNOR U620 ( .A(n12228), .B(n12266), .Z(n12232) );
  XNOR U621 ( .A(n12964), .B(n13002), .Z(n12968) );
  XNOR U622 ( .A(n13700), .B(n13738), .Z(n13704) );
  XNOR U623 ( .A(n14436), .B(n14474), .Z(n14440) );
  XNOR U624 ( .A(n15172), .B(n15210), .Z(n15176) );
  XNOR U625 ( .A(n15908), .B(n15946), .Z(n15912) );
  XNOR U626 ( .A(n16644), .B(n16682), .Z(n16648) );
  XNOR U627 ( .A(n17380), .B(n17418), .Z(n17384) );
  XNOR U628 ( .A(n18116), .B(n18154), .Z(n18120) );
  XNOR U629 ( .A(n18852), .B(n18890), .Z(n18856) );
  XNOR U630 ( .A(n19588), .B(n19626), .Z(n19592) );
  XNOR U631 ( .A(n20324), .B(n20362), .Z(n20328) );
  XNOR U632 ( .A(n21060), .B(n21098), .Z(n21064) );
  XNOR U633 ( .A(n21796), .B(n21834), .Z(n21800) );
  XNOR U634 ( .A(n1294), .B(n1330), .Z(n1298) );
  XNOR U635 ( .A(n5021), .B(n5052), .Z(n5025) );
  XNOR U636 ( .A(n11508), .B(n11136), .Z(n11138) );
  XNOR U637 ( .A(n11876), .B(n11505), .Z(n11507) );
  XNOR U638 ( .A(n22910), .B(n22936), .Z(n22914) );
  XNOR U639 ( .A(n10770), .B(n10789), .Z(n10774) );
  XNOR U640 ( .A(n12243), .B(n12263), .Z(n12247) );
  XNOR U641 ( .A(n12979), .B(n12999), .Z(n12983) );
  XNOR U642 ( .A(n13715), .B(n13735), .Z(n13719) );
  XNOR U643 ( .A(n14451), .B(n14471), .Z(n14455) );
  XNOR U644 ( .A(n15187), .B(n15207), .Z(n15191) );
  XNOR U645 ( .A(n15923), .B(n15943), .Z(n15927) );
  XNOR U646 ( .A(n16659), .B(n16679), .Z(n16663) );
  XNOR U647 ( .A(n17395), .B(n17415), .Z(n17399) );
  XNOR U648 ( .A(n18131), .B(n18151), .Z(n18135) );
  XNOR U649 ( .A(n18867), .B(n18887), .Z(n18871) );
  XNOR U650 ( .A(n19603), .B(n19623), .Z(n19607) );
  XNOR U651 ( .A(n20339), .B(n20359), .Z(n20343) );
  XNOR U652 ( .A(n21075), .B(n21095), .Z(n21079) );
  XNOR U653 ( .A(n21811), .B(n21831), .Z(n21815) );
  XNOR U654 ( .A(n22547), .B(n22567), .Z(n22551) );
  AND U655 ( .A(n6158), .B(n6159), .Z(n5786) );
  ANDN U656 ( .B(n7646), .A(n7647), .Z(n7274) );
  ANDN U657 ( .B(n9134), .A(n9135), .Z(n8762) );
  AND U658 ( .A(n7), .B(n8), .Z(n5) );
  AND U659 ( .A(n15), .B(n16), .Z(n13) );
  AND U660 ( .A(n23), .B(n24), .Z(n21) );
  AND U661 ( .A(n31), .B(n32), .Z(n29) );
  AND U662 ( .A(n39), .B(n40), .Z(n37) );
  AND U663 ( .A(n47), .B(n48), .Z(n45) );
  AND U664 ( .A(n55), .B(n56), .Z(n53) );
  AND U665 ( .A(n65), .B(n66), .Z(n63) );
  XNOR U666 ( .A(n8100), .B(n8461), .Z(n8105) );
  XNOR U667 ( .A(n8844), .B(n9201), .Z(n8849) );
  XNOR U668 ( .A(n9587), .B(n9953), .Z(n9592) );
  XNOR U669 ( .A(n13435), .B(n13792), .Z(n13440) );
  XNOR U670 ( .A(n17851), .B(n18208), .Z(n17856) );
  XNOR U671 ( .A(n24197), .B(n24553), .Z(n24201) );
  XNOR U672 ( .A(n23377), .B(n23807), .Z(n23381) );
  XNOR U673 ( .A(n10863), .B(n11213), .Z(n10867) );
  XNOR U674 ( .A(n11595), .B(n11950), .Z(n11604) );
  XNOR U675 ( .A(n14913), .B(n15263), .Z(n14917) );
  XNOR U676 ( .A(n19329), .B(n19679), .Z(n19333) );
  XNOR U677 ( .A(n21905), .B(n22255), .Z(n21909) );
  XNOR U678 ( .A(n22641), .B(n22991), .Z(n22645) );
  XNOR U679 ( .A(n16390), .B(n16734), .Z(n16394) );
  XNOR U680 ( .A(n20806), .B(n21150), .Z(n20810) );
  XNOR U681 ( .A(n7739), .B(n8087), .Z(n7743) );
  XNOR U682 ( .A(n8860), .B(n9198), .Z(n8864) );
  XNOR U683 ( .A(n9603), .B(n9950), .Z(n9607) );
  XNOR U684 ( .A(n13451), .B(n13789), .Z(n13455) );
  XNOR U685 ( .A(n17867), .B(n18205), .Z(n17871) );
  XNOR U686 ( .A(n25628), .B(n25966), .Z(n25632) );
  XNOR U687 ( .A(n24932), .B(n25270), .Z(n24936) );
  XNOR U688 ( .A(n24212), .B(n24550), .Z(n24216) );
  XNOR U689 ( .A(n23392), .B(n23804), .Z(n23396) );
  XNOR U690 ( .A(n10510), .B(n10841), .Z(n10514) );
  XNOR U691 ( .A(n11247), .B(n11579), .Z(n11251) );
  XNOR U692 ( .A(n11983), .B(n12315), .Z(n11987) );
  XNOR U693 ( .A(n12714), .B(n13051), .Z(n12723) );
  XNOR U694 ( .A(n14928), .B(n15260), .Z(n14932) );
  XNOR U695 ( .A(n19344), .B(n19676), .Z(n19348) );
  XNOR U696 ( .A(n21920), .B(n22252), .Z(n21924) );
  XNOR U697 ( .A(n22656), .B(n22988), .Z(n22660) );
  XNOR U698 ( .A(n8498), .B(n8828), .Z(n8502) );
  XNOR U699 ( .A(n16405), .B(n16731), .Z(n16409) );
  XNOR U700 ( .A(n20821), .B(n21147), .Z(n20825) );
  XNOR U701 ( .A(n7372), .B(n7714), .Z(n7376) );
  XNOR U702 ( .A(n9618), .B(n9947), .Z(n9622) );
  XNOR U703 ( .A(n17882), .B(n18202), .Z(n17886) );
  XNOR U704 ( .A(n26315), .B(n26635), .Z(n26319) );
  XNOR U705 ( .A(n25643), .B(n25963), .Z(n25647) );
  XNOR U706 ( .A(n24947), .B(n25267), .Z(n24951) );
  XNOR U707 ( .A(n24227), .B(n24547), .Z(n24231) );
  XNOR U708 ( .A(n23407), .B(n23801), .Z(n23411) );
  XNOR U709 ( .A(n8136), .B(n8454), .Z(n8140) );
  XNOR U710 ( .A(n10893), .B(n11207), .Z(n10897) );
  XNOR U711 ( .A(n11630), .B(n11944), .Z(n11634) );
  XNOR U712 ( .A(n12366), .B(n12680), .Z(n12370) );
  XNOR U713 ( .A(n13102), .B(n13416), .Z(n13106) );
  XNOR U714 ( .A(n13833), .B(n14152), .Z(n13842) );
  XNOR U715 ( .A(n14943), .B(n15257), .Z(n14947) );
  XNOR U716 ( .A(n19359), .B(n19673), .Z(n19363) );
  XNOR U717 ( .A(n21935), .B(n22249), .Z(n21939) );
  XNOR U718 ( .A(n22671), .B(n22985), .Z(n22675) );
  XNOR U719 ( .A(n9253), .B(n9568), .Z(n9257) );
  XNOR U720 ( .A(n16420), .B(n16728), .Z(n16424) );
  XNOR U721 ( .A(n20836), .B(n21144), .Z(n20840) );
  XNOR U722 ( .A(n7002), .B(n7341), .Z(n7006) );
  XNOR U723 ( .A(n17897), .B(n18199), .Z(n17901) );
  XNOR U724 ( .A(n27602), .B(n27904), .Z(n27606) );
  XNOR U725 ( .A(n26978), .B(n27280), .Z(n26982) );
  XNOR U726 ( .A(n26330), .B(n26632), .Z(n26334) );
  XNOR U727 ( .A(n25658), .B(n25960), .Z(n25662) );
  XNOR U728 ( .A(n24962), .B(n25264), .Z(n24966) );
  XNOR U729 ( .A(n24242), .B(n24544), .Z(n24246) );
  XNOR U730 ( .A(n23422), .B(n23798), .Z(n23426) );
  XNOR U731 ( .A(n8895), .B(n9191), .Z(n8899) );
  XNOR U732 ( .A(n10540), .B(n10835), .Z(n10544) );
  XNOR U733 ( .A(n11277), .B(n11573), .Z(n11281) );
  XNOR U734 ( .A(n12013), .B(n12309), .Z(n12017) );
  XNOR U735 ( .A(n12749), .B(n13045), .Z(n12753) );
  XNOR U736 ( .A(n13485), .B(n13781), .Z(n13489) );
  XNOR U737 ( .A(n14221), .B(n14517), .Z(n14225) );
  XNOR U738 ( .A(n14952), .B(n15253), .Z(n14961) );
  XNOR U739 ( .A(n19374), .B(n19670), .Z(n19378) );
  XNOR U740 ( .A(n21950), .B(n22246), .Z(n21954) );
  XNOR U741 ( .A(n22686), .B(n22982), .Z(n22690) );
  XNOR U742 ( .A(n7779), .B(n8079), .Z(n7783) );
  XNOR U743 ( .A(n9643), .B(n9942), .Z(n9647) );
  XNOR U744 ( .A(n16435), .B(n16725), .Z(n16439) );
  XNOR U745 ( .A(n20851), .B(n21141), .Z(n20855) );
  XNOR U746 ( .A(n6257), .B(n6599), .Z(n6261) );
  XNOR U747 ( .A(n17912), .B(n18196), .Z(n17916) );
  XNOR U748 ( .A(n28217), .B(n28501), .Z(n28221) );
  XNOR U749 ( .A(n27617), .B(n27901), .Z(n27621) );
  XNOR U750 ( .A(n26993), .B(n27277), .Z(n26997) );
  XNOR U751 ( .A(n26345), .B(n26629), .Z(n26349) );
  XNOR U752 ( .A(n25673), .B(n25957), .Z(n25677) );
  XNOR U753 ( .A(n24977), .B(n25261), .Z(n24981) );
  XNOR U754 ( .A(n24257), .B(n24541), .Z(n24261) );
  XNOR U755 ( .A(n23437), .B(n23795), .Z(n23441) );
  XNOR U756 ( .A(n8538), .B(n8820), .Z(n8542) );
  XNOR U757 ( .A(n9278), .B(n9563), .Z(n9282) );
  XNOR U758 ( .A(n10929), .B(n10558), .Z(n10560) );
  XNOR U759 ( .A(n10923), .B(n11201), .Z(n10927) );
  XNOR U760 ( .A(n11660), .B(n11938), .Z(n11664) );
  XNOR U761 ( .A(n12396), .B(n12674), .Z(n12400) );
  XNOR U762 ( .A(n13132), .B(n13410), .Z(n13136) );
  XNOR U763 ( .A(n13868), .B(n14146), .Z(n13872) );
  XNOR U764 ( .A(n14604), .B(n14882), .Z(n14608) );
  XNOR U765 ( .A(n15340), .B(n15618), .Z(n15344) );
  XNOR U766 ( .A(n16071), .B(n16354), .Z(n16080) );
  XNOR U767 ( .A(n19389), .B(n19667), .Z(n19393) );
  XNOR U768 ( .A(n21965), .B(n22243), .Z(n21969) );
  XNOR U769 ( .A(n22701), .B(n22979), .Z(n22705) );
  XNOR U770 ( .A(n7027), .B(n7336), .Z(n7031) );
  XNOR U771 ( .A(n20866), .B(n21138), .Z(n20870) );
  XNOR U772 ( .A(n7417), .B(n7705), .Z(n7421) );
  XNOR U773 ( .A(n6272), .B(n6596), .Z(n6276) );
  XNOR U774 ( .A(n5508), .B(n5856), .Z(n5512) );
  XNOR U775 ( .A(n17927), .B(n18193), .Z(n17931) );
  XNOR U776 ( .A(n29360), .B(n29626), .Z(n29364) );
  XNOR U777 ( .A(n28808), .B(n29074), .Z(n28812) );
  XNOR U778 ( .A(n28232), .B(n28498), .Z(n28236) );
  XNOR U779 ( .A(n27632), .B(n27898), .Z(n27636) );
  XNOR U780 ( .A(n27008), .B(n27274), .Z(n27012) );
  XNOR U781 ( .A(n26360), .B(n26626), .Z(n26364) );
  XNOR U782 ( .A(n25688), .B(n25954), .Z(n25692) );
  XNOR U783 ( .A(n24992), .B(n25258), .Z(n24996) );
  XNOR U784 ( .A(n24272), .B(n24538), .Z(n24276) );
  XNOR U785 ( .A(n23452), .B(n23792), .Z(n23456) );
  XNOR U786 ( .A(n7804), .B(n8074), .Z(n7808) );
  XNOR U787 ( .A(n9668), .B(n9937), .Z(n9672) );
  XNOR U788 ( .A(n10944), .B(n10573), .Z(n10575) );
  XNOR U789 ( .A(n11313), .B(n10941), .Z(n10943) );
  XNOR U790 ( .A(n11307), .B(n11567), .Z(n11311) );
  XNOR U791 ( .A(n12043), .B(n12303), .Z(n12047) );
  XNOR U792 ( .A(n12779), .B(n13039), .Z(n12783) );
  XNOR U793 ( .A(n13515), .B(n13775), .Z(n13519) );
  XNOR U794 ( .A(n14251), .B(n14511), .Z(n14255) );
  XNOR U795 ( .A(n14987), .B(n15247), .Z(n14991) );
  XNOR U796 ( .A(n15723), .B(n15983), .Z(n15727) );
  XNOR U797 ( .A(n16459), .B(n16719), .Z(n16463) );
  XNOR U798 ( .A(n17190), .B(n17455), .Z(n17199) );
  XNOR U799 ( .A(n19404), .B(n19664), .Z(n19408) );
  XNOR U800 ( .A(n21980), .B(n22240), .Z(n21984) );
  XNOR U801 ( .A(n22716), .B(n22976), .Z(n22720) );
  XNOR U802 ( .A(n8930), .B(n9184), .Z(n8934) );
  XNOR U803 ( .A(n20881), .B(n21135), .Z(n20885) );
  XNOR U804 ( .A(n6669), .B(n6959), .Z(n6673) );
  XNOR U805 ( .A(n5905), .B(n6223), .Z(n5909) );
  XNOR U806 ( .A(n29903), .B(n30151), .Z(n29907) );
  XNOR U807 ( .A(n29375), .B(n29623), .Z(n29379) );
  XNOR U808 ( .A(n28823), .B(n29071), .Z(n28827) );
  XNOR U809 ( .A(n28247), .B(n28495), .Z(n28251) );
  XNOR U810 ( .A(n27647), .B(n27895), .Z(n27651) );
  XNOR U811 ( .A(n27023), .B(n27271), .Z(n27027) );
  XNOR U812 ( .A(n26375), .B(n26623), .Z(n26379) );
  XNOR U813 ( .A(n25703), .B(n25951), .Z(n25707) );
  XNOR U814 ( .A(n25007), .B(n25255), .Z(n25011) );
  XNOR U815 ( .A(n24287), .B(n24535), .Z(n24291) );
  XNOR U816 ( .A(n23467), .B(n23789), .Z(n23471) );
  XNOR U817 ( .A(n11328), .B(n10956), .Z(n10958) );
  XNOR U818 ( .A(n11696), .B(n11325), .Z(n11327) );
  XNOR U819 ( .A(n12064), .B(n11693), .Z(n11695) );
  XNOR U820 ( .A(n12432), .B(n12061), .Z(n12063) );
  XNOR U821 ( .A(n12426), .B(n12668), .Z(n12430) );
  XNOR U822 ( .A(n13162), .B(n13404), .Z(n13166) );
  XNOR U823 ( .A(n13898), .B(n14140), .Z(n13902) );
  XNOR U824 ( .A(n14634), .B(n14876), .Z(n14638) );
  XNOR U825 ( .A(n15370), .B(n15612), .Z(n15374) );
  XNOR U826 ( .A(n16106), .B(n16348), .Z(n16110) );
  XNOR U827 ( .A(n16842), .B(n17084), .Z(n16846) );
  XNOR U828 ( .A(n17578), .B(n17820), .Z(n17582) );
  XNOR U829 ( .A(n18309), .B(n18556), .Z(n18318) );
  XNOR U830 ( .A(n19419), .B(n19661), .Z(n19423) );
  XNOR U831 ( .A(n21995), .B(n22237), .Z(n21999) );
  XNOR U832 ( .A(n22731), .B(n22973), .Z(n22735) );
  XNOR U833 ( .A(n8945), .B(n9181), .Z(n8949) );
  XNOR U834 ( .A(n9688), .B(n9933), .Z(n9692) );
  XNOR U835 ( .A(n11333), .B(n10961), .Z(n10963) );
  XNOR U836 ( .A(n20896), .B(n21132), .Z(n20900) );
  XNOR U837 ( .A(n7062), .B(n7329), .Z(n7066) );
  XNOR U838 ( .A(n5920), .B(n6220), .Z(n5924) );
  XNOR U839 ( .A(n5156), .B(n5480), .Z(n5160) );
  XNOR U840 ( .A(n8578), .B(n8812), .Z(n8582) );
  XNOR U841 ( .A(n11338), .B(n10966), .Z(n10968) );
  XNOR U842 ( .A(n30902), .B(n31132), .Z(n30906) );
  XNOR U843 ( .A(n30422), .B(n30652), .Z(n30426) );
  XNOR U844 ( .A(n29918), .B(n30148), .Z(n29922) );
  XNOR U845 ( .A(n29390), .B(n29620), .Z(n29394) );
  XNOR U846 ( .A(n28838), .B(n29068), .Z(n28842) );
  XNOR U847 ( .A(n28262), .B(n28492), .Z(n28266) );
  XNOR U848 ( .A(n27662), .B(n27892), .Z(n27666) );
  XNOR U849 ( .A(n27038), .B(n27268), .Z(n27042) );
  XNOR U850 ( .A(n26390), .B(n26620), .Z(n26394) );
  XNOR U851 ( .A(n25718), .B(n25948), .Z(n25722) );
  XNOR U852 ( .A(n25022), .B(n25252), .Z(n25026) );
  XNOR U853 ( .A(n24302), .B(n24532), .Z(n24306) );
  XNOR U854 ( .A(n23482), .B(n23786), .Z(n23486) );
  XNOR U855 ( .A(n7834), .B(n8068), .Z(n7838) );
  XNOR U856 ( .A(n4396), .B(n4738), .Z(n4400) );
  XNOR U857 ( .A(n12815), .B(n12444), .Z(n12446) );
  XNOR U858 ( .A(n13183), .B(n12812), .Z(n12814) );
  XNOR U859 ( .A(n13551), .B(n13180), .Z(n13182) );
  XNOR U860 ( .A(n13545), .B(n13769), .Z(n13549) );
  XNOR U861 ( .A(n14281), .B(n14505), .Z(n14285) );
  XNOR U862 ( .A(n15017), .B(n15241), .Z(n15021) );
  XNOR U863 ( .A(n15753), .B(n15977), .Z(n15757) );
  XNOR U864 ( .A(n16489), .B(n16713), .Z(n16493) );
  XNOR U865 ( .A(n17225), .B(n17449), .Z(n17229) );
  XNOR U866 ( .A(n17961), .B(n18185), .Z(n17965) );
  XNOR U867 ( .A(n18697), .B(n18921), .Z(n18701) );
  XNOR U868 ( .A(n19428), .B(n19657), .Z(n19437) );
  XNOR U869 ( .A(n22010), .B(n22234), .Z(n22014) );
  XNOR U870 ( .A(n22746), .B(n22970), .Z(n22750) );
  XNOR U871 ( .A(n9703), .B(n9930), .Z(n9707) );
  XNOR U872 ( .A(n10605), .B(n10822), .Z(n10609) );
  XNOR U873 ( .A(n20911), .B(n21129), .Z(n20915) );
  XNOR U874 ( .A(n7099), .B(n7321), .Z(n7100) );
  XNOR U875 ( .A(n6699), .B(n6953), .Z(n6703) );
  XNOR U876 ( .A(n5935), .B(n6217), .Z(n5939) );
  XNOR U877 ( .A(n5171), .B(n5477), .Z(n5175) );
  XNOR U878 ( .A(n8593), .B(n8809), .Z(n8597) );
  XNOR U879 ( .A(n9333), .B(n9552), .Z(n9337) );
  XNOR U880 ( .A(n11721), .B(n11350), .Z(n11352) );
  XNOR U881 ( .A(n12083), .B(n12295), .Z(n12087) );
  XNOR U882 ( .A(n31373), .B(n31585), .Z(n31377) );
  XNOR U883 ( .A(n30917), .B(n31129), .Z(n30921) );
  XNOR U884 ( .A(n30437), .B(n30649), .Z(n30441) );
  XNOR U885 ( .A(n29933), .B(n30145), .Z(n29937) );
  XNOR U886 ( .A(n29405), .B(n29617), .Z(n29409) );
  XNOR U887 ( .A(n28853), .B(n29065), .Z(n28857) );
  XNOR U888 ( .A(n28277), .B(n28489), .Z(n28281) );
  XNOR U889 ( .A(n27677), .B(n27889), .Z(n27681) );
  XNOR U890 ( .A(n27053), .B(n27265), .Z(n27057) );
  XNOR U891 ( .A(n26405), .B(n26617), .Z(n26409) );
  XNOR U892 ( .A(n25733), .B(n25945), .Z(n25737) );
  XNOR U893 ( .A(n25037), .B(n25249), .Z(n25041) );
  XNOR U894 ( .A(n24317), .B(n24529), .Z(n24321) );
  XNOR U895 ( .A(n23497), .B(n23783), .Z(n23501) );
  XNOR U896 ( .A(n7467), .B(n7695), .Z(n7475) );
  XNOR U897 ( .A(n4411), .B(n4735), .Z(n4415) );
  XNOR U898 ( .A(n3647), .B(n3995), .Z(n3651) );
  XNOR U899 ( .A(n11358), .B(n10986), .Z(n10988) );
  XNOR U900 ( .A(n13934), .B(n13563), .Z(n13565) );
  XNOR U901 ( .A(n14302), .B(n13931), .Z(n13933) );
  XNOR U902 ( .A(n14670), .B(n14299), .Z(n14301) );
  XNOR U903 ( .A(n14664), .B(n14870), .Z(n14668) );
  XNOR U904 ( .A(n15400), .B(n15606), .Z(n15404) );
  XNOR U905 ( .A(n16136), .B(n16342), .Z(n16140) );
  XNOR U906 ( .A(n16872), .B(n17078), .Z(n16876) );
  XNOR U907 ( .A(n17608), .B(n17814), .Z(n17612) );
  XNOR U908 ( .A(n18344), .B(n18550), .Z(n18348) );
  XNOR U909 ( .A(n19080), .B(n19286), .Z(n19084) );
  XNOR U910 ( .A(n19816), .B(n20022), .Z(n19820) );
  XNOR U911 ( .A(n20547), .B(n20758), .Z(n20556) );
  XNOR U912 ( .A(n22025), .B(n22231), .Z(n22029) );
  XNOR U913 ( .A(n22761), .B(n22967), .Z(n22765) );
  XNOR U914 ( .A(n7486), .B(n7690), .Z(n7490) );
  XNOR U915 ( .A(n11363), .B(n10991), .Z(n10993) );
  XNOR U916 ( .A(n6332), .B(n6584), .Z(n6336) );
  XNOR U917 ( .A(n5568), .B(n5844), .Z(n5572) );
  XNOR U918 ( .A(n8235), .B(n8433), .Z(n8239) );
  XNOR U919 ( .A(n8984), .B(n9174), .Z(n8979) );
  XNOR U920 ( .A(n9723), .B(n9926), .Z(n9727) );
  XNOR U921 ( .A(n12466), .B(n12660), .Z(n12470) );
  XNOR U922 ( .A(n13202), .B(n13396), .Z(n13206) );
  XNOR U923 ( .A(n32383), .B(n32572), .Z(n32387) );
  XNOR U924 ( .A(n31991), .B(n32177), .Z(n31995) );
  XNOR U925 ( .A(n31388), .B(n31582), .Z(n31392) );
  XNOR U926 ( .A(n30932), .B(n31126), .Z(n30936) );
  XNOR U927 ( .A(n30452), .B(n30646), .Z(n30456) );
  XNOR U928 ( .A(n29948), .B(n30142), .Z(n29952) );
  XNOR U929 ( .A(n29420), .B(n29614), .Z(n29424) );
  XNOR U930 ( .A(n28868), .B(n29062), .Z(n28872) );
  XNOR U931 ( .A(n28292), .B(n28486), .Z(n28296) );
  XNOR U932 ( .A(n27692), .B(n27886), .Z(n27696) );
  XNOR U933 ( .A(n27068), .B(n27262), .Z(n27072) );
  XNOR U934 ( .A(n26420), .B(n26614), .Z(n26424) );
  XNOR U935 ( .A(n25748), .B(n25942), .Z(n25752) );
  XNOR U936 ( .A(n25052), .B(n25246), .Z(n25056) );
  XNOR U937 ( .A(n24332), .B(n24526), .Z(n24336) );
  XNOR U938 ( .A(n23512), .B(n23780), .Z(n23516) );
  XNOR U939 ( .A(n5595), .B(n5838), .Z(n5596) );
  XNOR U940 ( .A(n11373), .B(n11001), .Z(n11003) );
  XNOR U941 ( .A(n12103), .B(n12291), .Z(n12107) );
  XNOR U942 ( .A(n15053), .B(n14682), .Z(n14684) );
  XNOR U943 ( .A(n15421), .B(n15050), .Z(n15052) );
  XNOR U944 ( .A(n15789), .B(n15418), .Z(n15420) );
  XNOR U945 ( .A(n15783), .B(n15971), .Z(n15787) );
  XNOR U946 ( .A(n16519), .B(n16707), .Z(n16523) );
  XNOR U947 ( .A(n17255), .B(n17443), .Z(n17259) );
  XNOR U948 ( .A(n17991), .B(n18179), .Z(n17995) );
  XNOR U949 ( .A(n18727), .B(n18915), .Z(n18731) );
  XNOR U950 ( .A(n19463), .B(n19651), .Z(n19467) );
  XNOR U951 ( .A(n20199), .B(n20387), .Z(n20203) );
  XNOR U952 ( .A(n20935), .B(n21123), .Z(n20939) );
  XNOR U953 ( .A(n21666), .B(n21859), .Z(n21675) );
  XNOR U954 ( .A(n22776), .B(n22964), .Z(n22780) );
  XNOR U955 ( .A(n6743), .B(n6943), .Z(n6751) );
  XNOR U956 ( .A(n6003), .B(n6201), .Z(n6007) );
  XNOR U957 ( .A(n11378), .B(n11006), .Z(n11008) );
  XNOR U958 ( .A(n4818), .B(n5101), .Z(n4822) );
  XNOR U959 ( .A(n3672), .B(n3990), .Z(n3676) );
  XNOR U960 ( .A(n6762), .B(n6938), .Z(n6766) );
  XNOR U961 ( .A(n7508), .B(n7685), .Z(n7509) );
  XNOR U962 ( .A(n8250), .B(n8430), .Z(n8258) );
  XNOR U963 ( .A(n8994), .B(n9170), .Z(n8998) );
  XNOR U964 ( .A(n13585), .B(n13761), .Z(n13589) );
  XNOR U965 ( .A(n14321), .B(n14497), .Z(n14325) );
  XNOR U966 ( .A(n32769), .B(n32937), .Z(n32773) );
  XNOR U967 ( .A(n32398), .B(n32569), .Z(n32402) );
  XNOR U968 ( .A(n32006), .B(n32174), .Z(n32010) );
  XNOR U969 ( .A(n31403), .B(n31579), .Z(n31407) );
  XNOR U970 ( .A(n30947), .B(n31123), .Z(n30951) );
  XNOR U971 ( .A(n30467), .B(n30643), .Z(n30471) );
  XNOR U972 ( .A(n29963), .B(n30139), .Z(n29967) );
  XNOR U973 ( .A(n29435), .B(n29611), .Z(n29439) );
  XNOR U974 ( .A(n28883), .B(n29059), .Z(n28887) );
  XNOR U975 ( .A(n28307), .B(n28483), .Z(n28311) );
  XNOR U976 ( .A(n27707), .B(n27883), .Z(n27711) );
  XNOR U977 ( .A(n27083), .B(n27259), .Z(n27087) );
  XNOR U978 ( .A(n26435), .B(n26611), .Z(n26439) );
  XNOR U979 ( .A(n25763), .B(n25939), .Z(n25767) );
  XNOR U980 ( .A(n25067), .B(n25243), .Z(n25071) );
  XNOR U981 ( .A(n24347), .B(n24523), .Z(n24351) );
  XNOR U982 ( .A(n23527), .B(n23777), .Z(n23535) );
  XNOR U983 ( .A(n4463), .B(n4724), .Z(n4464) );
  XNOR U984 ( .A(n5653), .B(n5824), .Z(n5654) );
  XNOR U985 ( .A(n11388), .B(n11016), .Z(n11018) );
  XNOR U986 ( .A(n11756), .B(n11385), .Z(n11387) );
  XNOR U987 ( .A(n12118), .B(n12288), .Z(n12122) );
  XNOR U988 ( .A(n13222), .B(n13392), .Z(n13226) );
  XNOR U989 ( .A(n16172), .B(n15801), .Z(n15803) );
  XNOR U990 ( .A(n16540), .B(n16169), .Z(n16171) );
  XNOR U991 ( .A(n16908), .B(n16537), .Z(n16539) );
  XNOR U992 ( .A(n16902), .B(n17072), .Z(n16906) );
  XNOR U993 ( .A(n17638), .B(n17808), .Z(n17642) );
  XNOR U994 ( .A(n18374), .B(n18544), .Z(n18378) );
  XNOR U995 ( .A(n19110), .B(n19280), .Z(n19114) );
  XNOR U996 ( .A(n19846), .B(n20016), .Z(n19850) );
  XNOR U997 ( .A(n20582), .B(n20752), .Z(n20586) );
  XNOR U998 ( .A(n21318), .B(n21488), .Z(n21322) );
  XNOR U999 ( .A(n22054), .B(n22224), .Z(n22058) );
  XNOR U1000 ( .A(n22785), .B(n22960), .Z(n22794) );
  XNOR U1001 ( .A(n2535), .B(n2878), .Z(n2539) );
  XNOR U1002 ( .A(n6018), .B(n6198), .Z(n6026) );
  XNOR U1003 ( .A(n5254), .B(n5458), .Z(n5258) );
  XNOR U1004 ( .A(n4492), .B(n4717), .Z(n4493) );
  XNOR U1005 ( .A(n11024), .B(n10653), .Z(n10655) );
  XNOR U1006 ( .A(n11393), .B(n11021), .Z(n11023) );
  XNOR U1007 ( .A(n12497), .B(n12126), .Z(n12128) );
  XNOR U1008 ( .A(n5235), .B(n5463), .Z(n5243) );
  XNOR U1009 ( .A(n4069), .B(n4357), .Z(n4073) );
  XNOR U1010 ( .A(n6781), .B(n6935), .Z(n6776) );
  XNOR U1011 ( .A(n7520), .B(n7682), .Z(n7524) );
  XNOR U1012 ( .A(n8264), .B(n8426), .Z(n8268) );
  XNOR U1013 ( .A(n9013), .B(n9167), .Z(n9008) );
  XNOR U1014 ( .A(n9752), .B(n9918), .Z(n9756) );
  XNOR U1015 ( .A(n14704), .B(n14862), .Z(n14708) );
  XNOR U1016 ( .A(n15440), .B(n15598), .Z(n15444) );
  XNOR U1017 ( .A(n33451), .B(n33604), .Z(n33455) );
  XNOR U1018 ( .A(n33131), .B(n33281), .Z(n33135) );
  XNOR U1019 ( .A(n32784), .B(n32934), .Z(n32788) );
  XNOR U1020 ( .A(n32413), .B(n32566), .Z(n32417) );
  XNOR U1021 ( .A(n32021), .B(n32171), .Z(n32025) );
  XNOR U1022 ( .A(n31418), .B(n31576), .Z(n31422) );
  XNOR U1023 ( .A(n30962), .B(n31120), .Z(n30966) );
  XNOR U1024 ( .A(n30482), .B(n30640), .Z(n30486) );
  XNOR U1025 ( .A(n29978), .B(n30136), .Z(n29982) );
  XNOR U1026 ( .A(n29450), .B(n29608), .Z(n29454) );
  XNOR U1027 ( .A(n28898), .B(n29056), .Z(n28902) );
  XNOR U1028 ( .A(n28322), .B(n28480), .Z(n28326) );
  XNOR U1029 ( .A(n27722), .B(n27880), .Z(n27726) );
  XNOR U1030 ( .A(n27098), .B(n27256), .Z(n27102) );
  XNOR U1031 ( .A(n26450), .B(n26608), .Z(n26454) );
  XNOR U1032 ( .A(n25778), .B(n25936), .Z(n25782) );
  XNOR U1033 ( .A(n25082), .B(n25240), .Z(n25086) );
  XNOR U1034 ( .A(n24362), .B(n24520), .Z(n24366) );
  XNOR U1035 ( .A(n23541), .B(n23774), .Z(n23545) );
  XNOR U1036 ( .A(n4521), .B(n4710), .Z(n4522) );
  XNOR U1037 ( .A(n4475), .B(n4721), .Z(n4479) );
  XNOR U1038 ( .A(n3711), .B(n3981), .Z(n3715) );
  XNOR U1039 ( .A(n6037), .B(n6193), .Z(n6041) );
  XNOR U1040 ( .A(n11403), .B(n11031), .Z(n11033) );
  XNOR U1041 ( .A(n13237), .B(n13389), .Z(n13241) );
  XNOR U1042 ( .A(n14341), .B(n14493), .Z(n14345) );
  XNOR U1043 ( .A(n17291), .B(n16920), .Z(n16922) );
  XNOR U1044 ( .A(n17659), .B(n17288), .Z(n17290) );
  XNOR U1045 ( .A(n18027), .B(n17656), .Z(n17658) );
  XNOR U1046 ( .A(n18389), .B(n18541), .Z(n18393) );
  XNOR U1047 ( .A(n19125), .B(n19277), .Z(n19129) );
  XNOR U1048 ( .A(n19861), .B(n20013), .Z(n19865) );
  XNOR U1049 ( .A(n20597), .B(n20749), .Z(n20601) );
  XNOR U1050 ( .A(n21333), .B(n21485), .Z(n21337) );
  XNOR U1051 ( .A(n22069), .B(n22221), .Z(n22073) );
  XNOR U1052 ( .A(n22805), .B(n22957), .Z(n22809) );
  XNOR U1053 ( .A(n2550), .B(n2875), .Z(n2554) );
  XNOR U1054 ( .A(n1785), .B(n2133), .Z(n1789) );
  XNOR U1055 ( .A(n4122), .B(n4344), .Z(n4126) );
  XNOR U1056 ( .A(n3361), .B(n3604), .Z(n3362) );
  XNOR U1057 ( .A(n4927), .B(n5075), .Z(n4928) );
  XNOR U1058 ( .A(n11408), .B(n11036), .Z(n11038) );
  XNOR U1059 ( .A(n11770), .B(n11916), .Z(n11774) );
  XNOR U1060 ( .A(n12506), .B(n12652), .Z(n12510) );
  XNOR U1061 ( .A(n13616), .B(n13245), .Z(n13247) );
  XNOR U1062 ( .A(n3320), .B(n3614), .Z(n3328) );
  XNOR U1063 ( .A(n5679), .B(n5819), .Z(n5674) );
  XNOR U1064 ( .A(n7537), .B(n7678), .Z(n7538) );
  XNOR U1065 ( .A(n8279), .B(n8423), .Z(n8287) );
  XNOR U1066 ( .A(n9023), .B(n9163), .Z(n9027) );
  XNOR U1067 ( .A(n15823), .B(n15963), .Z(n15827) );
  XNOR U1068 ( .A(n16559), .B(n16699), .Z(n16563) );
  XNOR U1069 ( .A(n33765), .B(n33897), .Z(n33769) );
  XNOR U1070 ( .A(n33466), .B(n33601), .Z(n33470) );
  XNOR U1071 ( .A(n33146), .B(n33278), .Z(n33150) );
  XNOR U1072 ( .A(n32799), .B(n32931), .Z(n32803) );
  XNOR U1073 ( .A(n32428), .B(n32563), .Z(n32432) );
  XNOR U1074 ( .A(n32036), .B(n32168), .Z(n32040) );
  XNOR U1075 ( .A(n31433), .B(n31573), .Z(n31437) );
  XNOR U1076 ( .A(n30977), .B(n31117), .Z(n30981) );
  XNOR U1077 ( .A(n30497), .B(n30637), .Z(n30501) );
  XNOR U1078 ( .A(n29993), .B(n30133), .Z(n29997) );
  XNOR U1079 ( .A(n29465), .B(n29605), .Z(n29469) );
  XNOR U1080 ( .A(n28913), .B(n29053), .Z(n28917) );
  XNOR U1081 ( .A(n28337), .B(n28477), .Z(n28341) );
  XNOR U1082 ( .A(n27737), .B(n27877), .Z(n27741) );
  XNOR U1083 ( .A(n27113), .B(n27253), .Z(n27117) );
  XNOR U1084 ( .A(n26465), .B(n26605), .Z(n26469) );
  XNOR U1085 ( .A(n25793), .B(n25933), .Z(n25797) );
  XNOR U1086 ( .A(n25097), .B(n25237), .Z(n25101) );
  XNOR U1087 ( .A(n24377), .B(n24517), .Z(n24381) );
  XNOR U1088 ( .A(n23556), .B(n23771), .Z(n23560) );
  XNOR U1089 ( .A(n4151), .B(n4337), .Z(n4155) );
  XNOR U1090 ( .A(n3390), .B(n3597), .Z(n3391) );
  XNOR U1091 ( .A(n2962), .B(n3238), .Z(n2966) );
  XNOR U1092 ( .A(n2199), .B(n2497), .Z(n2200) );
  XNOR U1093 ( .A(n6796), .B(n6930), .Z(n6800) );
  XNOR U1094 ( .A(n11418), .B(n11046), .Z(n11048) );
  XNOR U1095 ( .A(n11786), .B(n11415), .Z(n11417) );
  XNOR U1096 ( .A(n14356), .B(n14490), .Z(n14360) );
  XNOR U1097 ( .A(n15460), .B(n15594), .Z(n15464) );
  XNOR U1098 ( .A(n18410), .B(n18039), .Z(n18041) );
  XNOR U1099 ( .A(n18778), .B(n18407), .Z(n18409) );
  XNOR U1100 ( .A(n19146), .B(n18775), .Z(n18777) );
  XNOR U1101 ( .A(n19140), .B(n19274), .Z(n19144) );
  XNOR U1102 ( .A(n19876), .B(n20010), .Z(n19880) );
  XNOR U1103 ( .A(n20612), .B(n20746), .Z(n20616) );
  XNOR U1104 ( .A(n21348), .B(n21482), .Z(n21352) );
  XNOR U1105 ( .A(n22084), .B(n22218), .Z(n22088) );
  XNOR U1106 ( .A(n22820), .B(n22954), .Z(n22824) );
  XNOR U1107 ( .A(n2182), .B(n2501), .Z(n2186) );
  XNOR U1108 ( .A(n1418), .B(n1760), .Z(n1422) );
  XNOR U1109 ( .A(n2991), .B(n3231), .Z(n2995) );
  XNOR U1110 ( .A(n2228), .B(n2490), .Z(n2229) );
  XNOR U1111 ( .A(n4180), .B(n4330), .Z(n4184) );
  XNOR U1112 ( .A(n3419), .B(n3590), .Z(n3420) );
  XNOR U1113 ( .A(n5312), .B(n5444), .Z(n5316) );
  XNOR U1114 ( .A(n11054), .B(n10683), .Z(n10685) );
  XNOR U1115 ( .A(n11423), .B(n11051), .Z(n11053) );
  XNOR U1116 ( .A(n12153), .B(n12281), .Z(n12157) );
  XNOR U1117 ( .A(n12889), .B(n13017), .Z(n12893) );
  XNOR U1118 ( .A(n13625), .B(n13753), .Z(n13629) );
  XNOR U1119 ( .A(n14735), .B(n14364), .Z(n14366) );
  XNOR U1120 ( .A(n8293), .B(n8419), .Z(n8297) );
  XNOR U1121 ( .A(n9042), .B(n9160), .Z(n9037) );
  XNOR U1122 ( .A(n9781), .B(n9910), .Z(n9785) );
  XNOR U1123 ( .A(n16942), .B(n17064), .Z(n16946) );
  XNOR U1124 ( .A(n17678), .B(n17800), .Z(n17682) );
  XNOR U1125 ( .A(n34303), .B(n34420), .Z(n34307) );
  XNOR U1126 ( .A(n34055), .B(n34169), .Z(n34059) );
  XNOR U1127 ( .A(n33780), .B(n33894), .Z(n33784) );
  XNOR U1128 ( .A(n33481), .B(n33598), .Z(n33485) );
  XNOR U1129 ( .A(n33161), .B(n33275), .Z(n33165) );
  XNOR U1130 ( .A(n32814), .B(n32928), .Z(n32818) );
  XNOR U1131 ( .A(n32443), .B(n32560), .Z(n32447) );
  XNOR U1132 ( .A(n32051), .B(n32165), .Z(n32055) );
  XNOR U1133 ( .A(n31448), .B(n31570), .Z(n31452) );
  XNOR U1134 ( .A(n30992), .B(n31114), .Z(n30996) );
  XNOR U1135 ( .A(n30512), .B(n30634), .Z(n30516) );
  XNOR U1136 ( .A(n30008), .B(n30130), .Z(n30012) );
  XNOR U1137 ( .A(n29480), .B(n29602), .Z(n29484) );
  XNOR U1138 ( .A(n28928), .B(n29050), .Z(n28932) );
  XNOR U1139 ( .A(n28352), .B(n28474), .Z(n28356) );
  XNOR U1140 ( .A(n27752), .B(n27874), .Z(n27756) );
  XNOR U1141 ( .A(n27128), .B(n27250), .Z(n27132) );
  XNOR U1142 ( .A(n26480), .B(n26602), .Z(n26484) );
  XNOR U1143 ( .A(n25808), .B(n25930), .Z(n25812) );
  XNOR U1144 ( .A(n25112), .B(n25234), .Z(n25116) );
  XNOR U1145 ( .A(n24392), .B(n24514), .Z(n24396) );
  XNOR U1146 ( .A(n23571), .B(n23768), .Z(n23575) );
  XNOR U1147 ( .A(n3448), .B(n3583), .Z(n3449) );
  XNOR U1148 ( .A(n3020), .B(n3224), .Z(n3024) );
  XNOR U1149 ( .A(n2257), .B(n2483), .Z(n2258) );
  XNOR U1150 ( .A(n1829), .B(n2123), .Z(n1833) );
  XNOR U1151 ( .A(n1068), .B(n1383), .Z(n1069) );
  XNOR U1152 ( .A(n4576), .B(n4698), .Z(n4571) );
  XNOR U1153 ( .A(n7554), .B(n7674), .Z(n7562) );
  XNOR U1154 ( .A(n11433), .B(n11061), .Z(n11063) );
  XNOR U1155 ( .A(n15475), .B(n15591), .Z(n15479) );
  XNOR U1156 ( .A(n16579), .B(n16695), .Z(n16583) );
  XNOR U1157 ( .A(n19529), .B(n19158), .Z(n19160) );
  XNOR U1158 ( .A(n19897), .B(n19526), .Z(n19528) );
  XNOR U1159 ( .A(n20265), .B(n19894), .Z(n19896) );
  XNOR U1160 ( .A(n20627), .B(n20743), .Z(n20631) );
  XNOR U1161 ( .A(n21363), .B(n21479), .Z(n21367) );
  XNOR U1162 ( .A(n22099), .B(n22215), .Z(n22103) );
  XNOR U1163 ( .A(n22835), .B(n22951), .Z(n22839) );
  XNOR U1164 ( .A(n1051), .B(n1387), .Z(n1055) );
  XNOR U1165 ( .A(n1858), .B(n2116), .Z(n1862) );
  XNOR U1166 ( .A(n1097), .B(n1376), .Z(n1098) );
  XNOR U1167 ( .A(n3049), .B(n3217), .Z(n3053) );
  XNOR U1168 ( .A(n2286), .B(n2476), .Z(n2287) );
  XNOR U1169 ( .A(n6071), .B(n6185), .Z(n6075) );
  XNOR U1170 ( .A(n11438), .B(n11066), .Z(n11068) );
  XNOR U1171 ( .A(n11800), .B(n11910), .Z(n11804) );
  XNOR U1172 ( .A(n12536), .B(n12646), .Z(n12540) );
  XNOR U1173 ( .A(n13272), .B(n13382), .Z(n13276) );
  XNOR U1174 ( .A(n14008), .B(n14118), .Z(n14012) );
  XNOR U1175 ( .A(n14744), .B(n14854), .Z(n14748) );
  XNOR U1176 ( .A(n15854), .B(n15483), .Z(n15485) );
  XNOR U1177 ( .A(n4214), .B(n4322), .Z(n4218) );
  XNOR U1178 ( .A(n5334), .B(n5439), .Z(n5335) );
  XNOR U1179 ( .A(n9052), .B(n9156), .Z(n9056) );
  XNOR U1180 ( .A(n18061), .B(n18165), .Z(n18065) );
  XNOR U1181 ( .A(n18797), .B(n18901), .Z(n18801) );
  XNOR U1182 ( .A(n34545), .B(n34641), .Z(n34549) );
  XNOR U1183 ( .A(n34318), .B(n34417), .Z(n34322) );
  XNOR U1184 ( .A(n34070), .B(n34166), .Z(n34074) );
  XNOR U1185 ( .A(n33795), .B(n33891), .Z(n33799) );
  XNOR U1186 ( .A(n33496), .B(n33595), .Z(n33500) );
  XNOR U1187 ( .A(n33176), .B(n33272), .Z(n33180) );
  XNOR U1188 ( .A(n32829), .B(n32925), .Z(n32833) );
  XNOR U1189 ( .A(n32458), .B(n32557), .Z(n32462) );
  XNOR U1190 ( .A(n32066), .B(n32162), .Z(n32070) );
  XNOR U1191 ( .A(n31463), .B(n31567), .Z(n31467) );
  XNOR U1192 ( .A(n31007), .B(n31111), .Z(n31011) );
  XNOR U1193 ( .A(n30527), .B(n30631), .Z(n30531) );
  XNOR U1194 ( .A(n30023), .B(n30127), .Z(n30027) );
  XNOR U1195 ( .A(n29495), .B(n29599), .Z(n29499) );
  XNOR U1196 ( .A(n28943), .B(n29047), .Z(n28947) );
  XNOR U1197 ( .A(n28367), .B(n28471), .Z(n28371) );
  XNOR U1198 ( .A(n27767), .B(n27871), .Z(n27771) );
  XNOR U1199 ( .A(n27143), .B(n27247), .Z(n27147) );
  XNOR U1200 ( .A(n26495), .B(n26599), .Z(n26499) );
  XNOR U1201 ( .A(n25823), .B(n25927), .Z(n25827) );
  XNOR U1202 ( .A(n25127), .B(n25231), .Z(n25131) );
  XNOR U1203 ( .A(n24407), .B(n24511), .Z(n24411) );
  XNOR U1204 ( .A(n23586), .B(n23765), .Z(n23590) );
  XNOR U1205 ( .A(n3078), .B(n3210), .Z(n3082) );
  XNOR U1206 ( .A(n2315), .B(n2469), .Z(n2316) );
  XNOR U1207 ( .A(n1887), .B(n2109), .Z(n1891) );
  XNOR U1208 ( .A(n1126), .B(n1369), .Z(n1127) );
  XNOR U1209 ( .A(n1080), .B(n1380), .Z(n1084) );
  XNOR U1210 ( .A(n4963), .B(n5066), .Z(n4967) );
  XNOR U1211 ( .A(n8317), .B(n8415), .Z(n8312) );
  XNOR U1212 ( .A(n11448), .B(n11076), .Z(n11078) );
  XNOR U1213 ( .A(n11816), .B(n11445), .Z(n11447) );
  XNOR U1214 ( .A(n16594), .B(n16692), .Z(n16598) );
  XNOR U1215 ( .A(n17698), .B(n17796), .Z(n17702) );
  XNOR U1216 ( .A(n19912), .B(n19541), .Z(n19543) );
  XNOR U1217 ( .A(n20280), .B(n19909), .Z(n19911) );
  XNOR U1218 ( .A(n20648), .B(n20277), .Z(n20279) );
  XNOR U1219 ( .A(n21384), .B(n21013), .Z(n21015) );
  XNOR U1220 ( .A(n21378), .B(n21476), .Z(n21382) );
  XNOR U1221 ( .A(n22114), .B(n22212), .Z(n22118) );
  XNOR U1222 ( .A(n22850), .B(n22948), .Z(n22854) );
  XNOR U1223 ( .A(n3851), .B(n3949), .Z(n3846) );
  XNOR U1224 ( .A(n1109), .B(n1373), .Z(n1113) );
  XNOR U1225 ( .A(n1916), .B(n2102), .Z(n1920) );
  XNOR U1226 ( .A(n1155), .B(n1362), .Z(n1156) );
  XNOR U1227 ( .A(n2344), .B(n2462), .Z(n2345) );
  XNOR U1228 ( .A(n6830), .B(n6922), .Z(n6838) );
  XNOR U1229 ( .A(n11084), .B(n10713), .Z(n10715) );
  XNOR U1230 ( .A(n11453), .B(n11081), .Z(n11083) );
  XNOR U1231 ( .A(n12183), .B(n12275), .Z(n12187) );
  XNOR U1232 ( .A(n12919), .B(n13011), .Z(n12923) );
  XNOR U1233 ( .A(n13655), .B(n13747), .Z(n13659) );
  XNOR U1234 ( .A(n14391), .B(n14483), .Z(n14395) );
  XNOR U1235 ( .A(n15127), .B(n15219), .Z(n15131) );
  XNOR U1236 ( .A(n15863), .B(n15955), .Z(n15867) );
  XNOR U1237 ( .A(n16973), .B(n16602), .Z(n16604) );
  XNOR U1238 ( .A(n6090), .B(n6180), .Z(n6094) );
  XNOR U1239 ( .A(n9810), .B(n9902), .Z(n9814) );
  XNOR U1240 ( .A(n19180), .B(n19266), .Z(n19184) );
  XNOR U1241 ( .A(n34939), .B(n35020), .Z(n34943) );
  XNOR U1242 ( .A(n34763), .B(n34841), .Z(n34767) );
  XNOR U1243 ( .A(n34560), .B(n34638), .Z(n34564) );
  XNOR U1244 ( .A(n34333), .B(n34414), .Z(n34337) );
  XNOR U1245 ( .A(n34085), .B(n34163), .Z(n34089) );
  XNOR U1246 ( .A(n33810), .B(n33888), .Z(n33814) );
  XNOR U1247 ( .A(n33511), .B(n33592), .Z(n33515) );
  XNOR U1248 ( .A(n33191), .B(n33269), .Z(n33195) );
  XNOR U1249 ( .A(n32844), .B(n32922), .Z(n32848) );
  XNOR U1250 ( .A(n32473), .B(n32554), .Z(n32477) );
  XNOR U1251 ( .A(n32081), .B(n32159), .Z(n32085) );
  XNOR U1252 ( .A(n31478), .B(n31564), .Z(n31482) );
  XNOR U1253 ( .A(n31022), .B(n31108), .Z(n31026) );
  XNOR U1254 ( .A(n30542), .B(n30628), .Z(n30546) );
  XNOR U1255 ( .A(n30038), .B(n30124), .Z(n30042) );
  XNOR U1256 ( .A(n29510), .B(n29596), .Z(n29514) );
  XNOR U1257 ( .A(n28958), .B(n29044), .Z(n28962) );
  XNOR U1258 ( .A(n28382), .B(n28468), .Z(n28386) );
  XNOR U1259 ( .A(n27782), .B(n27868), .Z(n27786) );
  XNOR U1260 ( .A(n27158), .B(n27244), .Z(n27162) );
  XNOR U1261 ( .A(n26510), .B(n26596), .Z(n26514) );
  XNOR U1262 ( .A(n25838), .B(n25924), .Z(n25842) );
  XNOR U1263 ( .A(n25142), .B(n25228), .Z(n25146) );
  XNOR U1264 ( .A(n24422), .B(n24508), .Z(n24426) );
  XNOR U1265 ( .A(n23601), .B(n23762), .Z(n23605) );
  XNOR U1266 ( .A(n1945), .B(n2095), .Z(n1949) );
  XNOR U1267 ( .A(n1184), .B(n1355), .Z(n1185) );
  XNOR U1268 ( .A(n1138), .B(n1366), .Z(n1142) );
  XNOR U1269 ( .A(n3489), .B(n3573), .Z(n3493) );
  XNOR U1270 ( .A(n4233), .B(n4317), .Z(n4237) );
  XNOR U1271 ( .A(n4982), .B(n5063), .Z(n4977) );
  XNOR U1272 ( .A(n5723), .B(n5807), .Z(n5727) );
  XNOR U1273 ( .A(n9074), .B(n9151), .Z(n9075) );
  XNOR U1274 ( .A(n11463), .B(n11091), .Z(n11093) );
  XNOR U1275 ( .A(n17713), .B(n17793), .Z(n17717) );
  XNOR U1276 ( .A(n18817), .B(n18897), .Z(n18821) );
  XNOR U1277 ( .A(n19921), .B(n20001), .Z(n19925) );
  XNOR U1278 ( .A(n21031), .B(n20660), .Z(n20662) );
  XNOR U1279 ( .A(n21399), .B(n21028), .Z(n21030) );
  XNOR U1280 ( .A(n21393), .B(n21473), .Z(n21397) );
  XNOR U1281 ( .A(n22129), .B(n22209), .Z(n22133) );
  XNOR U1282 ( .A(n22865), .B(n22945), .Z(n22869) );
  XNOR U1283 ( .A(n1167), .B(n1359), .Z(n1171) );
  XNOR U1284 ( .A(n1974), .B(n2088), .Z(n1978) );
  XNOR U1285 ( .A(n1213), .B(n1348), .Z(n1214) );
  XNOR U1286 ( .A(n7592), .B(n7666), .Z(n7587) );
  XNOR U1287 ( .A(n11468), .B(n11096), .Z(n11098) );
  XNOR U1288 ( .A(n11830), .B(n11904), .Z(n11834) );
  XNOR U1289 ( .A(n12566), .B(n12640), .Z(n12570) );
  XNOR U1290 ( .A(n13302), .B(n13376), .Z(n13306) );
  XNOR U1291 ( .A(n14038), .B(n14112), .Z(n14042) );
  XNOR U1292 ( .A(n14774), .B(n14848), .Z(n14778) );
  XNOR U1293 ( .A(n15510), .B(n15584), .Z(n15514) );
  XNOR U1294 ( .A(n16246), .B(n16320), .Z(n16250) );
  XNOR U1295 ( .A(n16982), .B(n17056), .Z(n16986) );
  XNOR U1296 ( .A(n18092), .B(n17721), .Z(n17723) );
  XNOR U1297 ( .A(n3129), .B(n3198), .Z(n3130) );
  XNOR U1298 ( .A(n6849), .B(n6917), .Z(n6853) );
  XNOR U1299 ( .A(n8337), .B(n8409), .Z(n8345) );
  XNOR U1300 ( .A(n35109), .B(n35169), .Z(n35113) );
  XNOR U1301 ( .A(n34954), .B(n35017), .Z(n34958) );
  XNOR U1302 ( .A(n34778), .B(n34838), .Z(n34782) );
  XNOR U1303 ( .A(n34575), .B(n34635), .Z(n34579) );
  XNOR U1304 ( .A(n34348), .B(n34411), .Z(n34352) );
  XNOR U1305 ( .A(n34100), .B(n34160), .Z(n34104) );
  XNOR U1306 ( .A(n33825), .B(n33885), .Z(n33829) );
  XNOR U1307 ( .A(n33526), .B(n33589), .Z(n33530) );
  XNOR U1308 ( .A(n33206), .B(n33266), .Z(n33210) );
  XNOR U1309 ( .A(n32859), .B(n32919), .Z(n32863) );
  XNOR U1310 ( .A(n32488), .B(n32551), .Z(n32492) );
  XNOR U1311 ( .A(n32096), .B(n32156), .Z(n32100) );
  XNOR U1312 ( .A(n31493), .B(n31561), .Z(n31497) );
  XNOR U1313 ( .A(n31037), .B(n31105), .Z(n31041) );
  XNOR U1314 ( .A(n30557), .B(n30625), .Z(n30561) );
  XNOR U1315 ( .A(n30053), .B(n30121), .Z(n30057) );
  XNOR U1316 ( .A(n29525), .B(n29593), .Z(n29529) );
  XNOR U1317 ( .A(n28973), .B(n29041), .Z(n28977) );
  XNOR U1318 ( .A(n28397), .B(n28465), .Z(n28401) );
  XNOR U1319 ( .A(n27797), .B(n27865), .Z(n27801) );
  XNOR U1320 ( .A(n27173), .B(n27241), .Z(n27177) );
  XNOR U1321 ( .A(n26525), .B(n26593), .Z(n26529) );
  XNOR U1322 ( .A(n25853), .B(n25921), .Z(n25857) );
  XNOR U1323 ( .A(n25157), .B(n25225), .Z(n25161) );
  XNOR U1324 ( .A(n24437), .B(n24505), .Z(n24441) );
  XNOR U1325 ( .A(n23616), .B(n23759), .Z(n23620) );
  XNOR U1326 ( .A(n1196), .B(n1352), .Z(n1200) );
  XNOR U1327 ( .A(n2758), .B(n2825), .Z(n2762) );
  XNOR U1328 ( .A(n4248), .B(n4314), .Z(n4256) );
  XNOR U1329 ( .A(n4992), .B(n5059), .Z(n4996) );
  XNOR U1330 ( .A(n5740), .B(n5803), .Z(n5741) );
  XNOR U1331 ( .A(n6482), .B(n6548), .Z(n6490) );
  XNOR U1332 ( .A(n9829), .B(n9896), .Z(n9833) );
  XNOR U1333 ( .A(n11478), .B(n11106), .Z(n11108) );
  XNOR U1334 ( .A(n11846), .B(n11475), .Z(n11477) );
  XNOR U1335 ( .A(n18832), .B(n18894), .Z(n18836) );
  XNOR U1336 ( .A(n19936), .B(n19998), .Z(n19940) );
  XNOR U1337 ( .A(n21040), .B(n21102), .Z(n21044) );
  XNOR U1338 ( .A(n21776), .B(n21838), .Z(n21780) );
  XNOR U1339 ( .A(n22880), .B(n22942), .Z(n22884) );
  XNOR U1340 ( .A(n1626), .B(n1710), .Z(n1630) );
  XNOR U1341 ( .A(n1225), .B(n1345), .Z(n1229) );
  XNOR U1342 ( .A(n1646), .B(n1706), .Z(n1650) );
  XNOR U1343 ( .A(n2390), .B(n2450), .Z(n2394) );
  XNOR U1344 ( .A(n11114), .B(n10743), .Z(n10745) );
  XNOR U1345 ( .A(n11483), .B(n11111), .Z(n11113) );
  XNOR U1346 ( .A(n12213), .B(n12269), .Z(n12217) );
  XNOR U1347 ( .A(n12949), .B(n13005), .Z(n12953) );
  XNOR U1348 ( .A(n13685), .B(n13741), .Z(n13689) );
  XNOR U1349 ( .A(n14421), .B(n14477), .Z(n14425) );
  XNOR U1350 ( .A(n15157), .B(n15213), .Z(n15161) );
  XNOR U1351 ( .A(n15893), .B(n15949), .Z(n15897) );
  XNOR U1352 ( .A(n16629), .B(n16685), .Z(n16633) );
  XNOR U1353 ( .A(n17365), .B(n17421), .Z(n17369) );
  XNOR U1354 ( .A(n18101), .B(n18157), .Z(n18105) );
  XNOR U1355 ( .A(n19211), .B(n18840), .Z(n18842) );
  XNOR U1356 ( .A(n21051), .B(n20680), .Z(n20682) );
  XNOR U1357 ( .A(n21419), .B(n21048), .Z(n21050) );
  XNOR U1358 ( .A(n22517), .B(n22573), .Z(n22521) );
  XNOR U1359 ( .A(n7607), .B(n7661), .Z(n7611) );
  XNOR U1360 ( .A(n9100), .B(n9146), .Z(n9095) );
  XNOR U1361 ( .A(n35310), .B(n35352), .Z(n35314) );
  XNOR U1362 ( .A(n35191), .B(n35236), .Z(n35195) );
  XNOR U1363 ( .A(n35051), .B(n35093), .Z(n35055) );
  XNOR U1364 ( .A(n34884), .B(n34926), .Z(n34888) );
  XNOR U1365 ( .A(n34693), .B(n34738), .Z(n34697) );
  XNOR U1366 ( .A(n34481), .B(n34523), .Z(n34485) );
  XNOR U1367 ( .A(n34242), .B(n34284), .Z(n34246) );
  XNOR U1368 ( .A(n33979), .B(n34024), .Z(n33983) );
  XNOR U1369 ( .A(n33695), .B(n33737), .Z(n33699) );
  XNOR U1370 ( .A(n33384), .B(n33426), .Z(n33388) );
  XNOR U1371 ( .A(n33049), .B(n33094), .Z(n33053) );
  XNOR U1372 ( .A(n32693), .B(n32735), .Z(n32697) );
  XNOR U1373 ( .A(n32310), .B(n32352), .Z(n32314) );
  XNOR U1374 ( .A(n31727), .B(n31948), .Z(n31731) );
  XNOR U1375 ( .A(n31283), .B(n31333), .Z(n31287) );
  XNOR U1376 ( .A(n30815), .B(n30865), .Z(n30819) );
  XNOR U1377 ( .A(n30323), .B(n30373), .Z(n30327) );
  XNOR U1378 ( .A(n29807), .B(n29857), .Z(n29811) );
  XNOR U1379 ( .A(n29267), .B(n29317), .Z(n29271) );
  XNOR U1380 ( .A(n28703), .B(n28753), .Z(n28707) );
  XNOR U1381 ( .A(n28115), .B(n28165), .Z(n28119) );
  XNOR U1382 ( .A(n27503), .B(n27553), .Z(n27507) );
  XNOR U1383 ( .A(n26867), .B(n26917), .Z(n26871) );
  XNOR U1384 ( .A(n26207), .B(n26257), .Z(n26211) );
  XNOR U1385 ( .A(n25523), .B(n25573), .Z(n25527) );
  XNOR U1386 ( .A(n24815), .B(n24865), .Z(n24819) );
  XNOR U1387 ( .A(n24080), .B(n24130), .Z(n24084) );
  XNOR U1388 ( .A(n1279), .B(n1333), .Z(n1283) );
  XNOR U1389 ( .A(n3518), .B(n3566), .Z(n3522) );
  XNOR U1390 ( .A(n4637), .B(n4682), .Z(n4638) );
  XNOR U1391 ( .A(n6871), .B(n6912), .Z(n6872) );
  XNOR U1392 ( .A(n11493), .B(n11121), .Z(n11123) );
  XNOR U1393 ( .A(n19951), .B(n19995), .Z(n19955) );
  XNOR U1394 ( .A(n22159), .B(n22203), .Z(n22163) );
  XNOR U1395 ( .A(n4267), .B(n4309), .Z(n4271) );
  XNOR U1396 ( .A(n11498), .B(n11126), .Z(n11128) );
  XNOR U1397 ( .A(n11860), .B(n11898), .Z(n11864) );
  XNOR U1398 ( .A(n12596), .B(n12634), .Z(n12600) );
  XNOR U1399 ( .A(n13332), .B(n13370), .Z(n13336) );
  XNOR U1400 ( .A(n14068), .B(n14106), .Z(n14072) );
  XNOR U1401 ( .A(n14804), .B(n14842), .Z(n14808) );
  XNOR U1402 ( .A(n15540), .B(n15578), .Z(n15544) );
  XNOR U1403 ( .A(n16276), .B(n16314), .Z(n16280) );
  XNOR U1404 ( .A(n17012), .B(n17050), .Z(n17016) );
  XNOR U1405 ( .A(n17748), .B(n17786), .Z(n17752) );
  XNOR U1406 ( .A(n18484), .B(n18522), .Z(n18488) );
  XNOR U1407 ( .A(n19220), .B(n19258), .Z(n19224) );
  XNOR U1408 ( .A(n20330), .B(n19959), .Z(n19961) );
  XNOR U1409 ( .A(n20692), .B(n20730), .Z(n20696) );
  XNOR U1410 ( .A(n21428), .B(n21466), .Z(n21432) );
  XNOR U1411 ( .A(n22538), .B(n22167), .Z(n22169) );
  XNOR U1412 ( .A(n22900), .B(n22938), .Z(n22904) );
  XNOR U1413 ( .A(n23641), .B(n23754), .Z(n23645) );
  XNOR U1414 ( .A(n1666), .B(n1702), .Z(n1670) );
  XNOR U1415 ( .A(n6134), .B(n6170), .Z(n6142) );
  XNOR U1416 ( .A(n7998), .B(n8030), .Z(n7993) );
  XNOR U1417 ( .A(n9110), .B(n9142), .Z(n9114) );
  XNOR U1418 ( .A(n35457), .B(n35481), .Z(n35461) );
  XNOR U1419 ( .A(n35374), .B(n35401), .Z(n35378) );
  XNOR U1420 ( .A(n35270), .B(n35294), .Z(n35274) );
  XNOR U1421 ( .A(n35139), .B(n35163), .Z(n35143) );
  XNOR U1422 ( .A(n34984), .B(n35011), .Z(n34988) );
  XNOR U1423 ( .A(n34808), .B(n34832), .Z(n34812) );
  XNOR U1424 ( .A(n34605), .B(n34629), .Z(n34609) );
  XNOR U1425 ( .A(n34378), .B(n34405), .Z(n34382) );
  XNOR U1426 ( .A(n34130), .B(n34154), .Z(n34134) );
  XNOR U1427 ( .A(n33855), .B(n33879), .Z(n33859) );
  XNOR U1428 ( .A(n33556), .B(n33583), .Z(n33560) );
  XNOR U1429 ( .A(n33236), .B(n33260), .Z(n33240) );
  XNOR U1430 ( .A(n32889), .B(n32913), .Z(n32893) );
  XNOR U1431 ( .A(n32518), .B(n32545), .Z(n32522) );
  XNOR U1432 ( .A(n32126), .B(n32150), .Z(n32130) );
  XNOR U1433 ( .A(n31523), .B(n31555), .Z(n31527) );
  XNOR U1434 ( .A(n31067), .B(n31099), .Z(n31071) );
  XNOR U1435 ( .A(n30587), .B(n30619), .Z(n30591) );
  XNOR U1436 ( .A(n30083), .B(n30115), .Z(n30087) );
  XNOR U1437 ( .A(n29555), .B(n29587), .Z(n29559) );
  XNOR U1438 ( .A(n29003), .B(n29035), .Z(n29007) );
  XNOR U1439 ( .A(n28427), .B(n28459), .Z(n28431) );
  XNOR U1440 ( .A(n27827), .B(n27859), .Z(n27831) );
  XNOR U1441 ( .A(n27203), .B(n27235), .Z(n27207) );
  XNOR U1442 ( .A(n26555), .B(n26587), .Z(n26559) );
  XNOR U1443 ( .A(n25883), .B(n25915), .Z(n25887) );
  XNOR U1444 ( .A(n25187), .B(n25219), .Z(n25191) );
  XNOR U1445 ( .A(n24467), .B(n24499), .Z(n24471) );
  XNOR U1446 ( .A(n927), .B(n957), .Z(n931) );
  XNOR U1447 ( .A(n2415), .B(n2445), .Z(n2419) );
  XNOR U1448 ( .A(n3161), .B(n3191), .Z(n3165) );
  XNOR U1449 ( .A(n3905), .B(n3935), .Z(n3909) );
  XNOR U1450 ( .A(n5394), .B(n5424), .Z(n5398) );
  XNOR U1451 ( .A(n6883), .B(n6909), .Z(n6887) );
  XNOR U1452 ( .A(n7626), .B(n7656), .Z(n7630) );
  XNOR U1453 ( .A(n8743), .B(n8773), .Z(n8751) );
  XNOR U1454 ( .A(n9858), .B(n9888), .Z(n9862) );
  XNOR U1455 ( .A(n11144), .B(n10773), .Z(n10775) );
  XNOR U1456 ( .A(n11513), .B(n11141), .Z(n11143) );
  XNOR U1457 ( .A(n11881), .B(n11510), .Z(n11512) );
  XNOR U1458 ( .A(n11875), .B(n11895), .Z(n11879) );
  XNOR U1459 ( .A(n12611), .B(n12631), .Z(n12615) );
  XNOR U1460 ( .A(n13347), .B(n13367), .Z(n13351) );
  XNOR U1461 ( .A(n14083), .B(n14103), .Z(n14087) );
  XNOR U1462 ( .A(n14819), .B(n14839), .Z(n14823) );
  XNOR U1463 ( .A(n15555), .B(n15575), .Z(n15559) );
  XNOR U1464 ( .A(n16291), .B(n16311), .Z(n16295) );
  XNOR U1465 ( .A(n17027), .B(n17047), .Z(n17031) );
  XNOR U1466 ( .A(n17763), .B(n17783), .Z(n17767) );
  XNOR U1467 ( .A(n18499), .B(n18519), .Z(n18503) );
  XNOR U1468 ( .A(n19235), .B(n19255), .Z(n19239) );
  XNOR U1469 ( .A(n19971), .B(n19991), .Z(n19975) );
  XNOR U1470 ( .A(n20707), .B(n20727), .Z(n20711) );
  XNOR U1471 ( .A(n21443), .B(n21463), .Z(n21447) );
  XNOR U1472 ( .A(n22179), .B(n22199), .Z(n22183) );
  XNOR U1473 ( .A(n22915), .B(n22935), .Z(n22919) );
  AND U1474 ( .A(n5414), .B(n5415), .Z(n5041) );
  AND U1475 ( .A(n6902), .B(n6903), .Z(n6530) );
  ANDN U1476 ( .B(n8390), .A(n8391), .Z(n8018) );
  ANDN U1477 ( .B(n9878), .A(n9879), .Z(n9506) );
  AND U1478 ( .A(n9), .B(n10), .Z(n7) );
  AND U1479 ( .A(n17), .B(n18), .Z(n15) );
  AND U1480 ( .A(n25), .B(n26), .Z(n23) );
  AND U1481 ( .A(n33), .B(n34), .Z(n31) );
  AND U1482 ( .A(n41), .B(n42), .Z(n39) );
  AND U1483 ( .A(n49), .B(n50), .Z(n47) );
  AND U1484 ( .A(n57), .B(n58), .Z(n55) );
  AND U1485 ( .A(n67), .B(n68), .Z(n65) );
  XNOR U1486 ( .A(n22267), .B(n22624), .Z(n22272) );
  XNOR U1487 ( .A(n24560), .B(n24916), .Z(n24564) );
  XNOR U1488 ( .A(n23825), .B(n24181), .Z(n23829) );
  XNOR U1489 ( .A(n8478), .B(n8832), .Z(n8482) );
  XNOR U1490 ( .A(n9218), .B(n9575), .Z(n9222) );
  XNOR U1491 ( .A(n9970), .B(n10474), .Z(n9974) );
  XNOR U1492 ( .A(n10869), .B(n10498), .Z(n10500) );
  XNOR U1493 ( .A(n11238), .B(n10866), .Z(n10868) );
  XNOR U1494 ( .A(n11606), .B(n11235), .Z(n11237) );
  XNOR U1495 ( .A(n11974), .B(n11603), .Z(n11605) );
  XNOR U1496 ( .A(n12337), .B(n12687), .Z(n12345) );
  XNOR U1497 ( .A(n13073), .B(n13423), .Z(n13077) );
  XNOR U1498 ( .A(n13809), .B(n14159), .Z(n13813) );
  XNOR U1499 ( .A(n14545), .B(n14895), .Z(n14549) );
  XNOR U1500 ( .A(n15281), .B(n15631), .Z(n15285) );
  XNOR U1501 ( .A(n16017), .B(n16367), .Z(n16021) );
  XNOR U1502 ( .A(n16753), .B(n17103), .Z(n16757) );
  XNOR U1503 ( .A(n17489), .B(n17839), .Z(n17493) );
  XNOR U1504 ( .A(n18225), .B(n18575), .Z(n18229) );
  XNOR U1505 ( .A(n18961), .B(n19311), .Z(n18965) );
  XNOR U1506 ( .A(n19697), .B(n20047), .Z(n19701) );
  XNOR U1507 ( .A(n20433), .B(n20783), .Z(n20437) );
  XNOR U1508 ( .A(n21169), .B(n21519), .Z(n21173) );
  XNOR U1509 ( .A(n23009), .B(n23359), .Z(n23013) );
  XNOR U1510 ( .A(n22283), .B(n22621), .Z(n22287) );
  XNOR U1511 ( .A(n25283), .B(n25621), .Z(n25287) );
  XNOR U1512 ( .A(n24575), .B(n24913), .Z(n24579) );
  XNOR U1513 ( .A(n23840), .B(n24178), .Z(n23844) );
  XNOR U1514 ( .A(n7744), .B(n8086), .Z(n7748) );
  XNOR U1515 ( .A(n8493), .B(n8829), .Z(n8497) );
  XNOR U1516 ( .A(n9233), .B(n9572), .Z(n9237) );
  XNOR U1517 ( .A(n9985), .B(n10468), .Z(n9989) );
  XNOR U1518 ( .A(n10884), .B(n10513), .Z(n10515) );
  XNOR U1519 ( .A(n11253), .B(n10881), .Z(n10883) );
  XNOR U1520 ( .A(n11621), .B(n11250), .Z(n11252) );
  XNOR U1521 ( .A(n11989), .B(n11618), .Z(n11620) );
  XNOR U1522 ( .A(n12357), .B(n11986), .Z(n11988) );
  XNOR U1523 ( .A(n12725), .B(n12354), .Z(n12356) );
  XNOR U1524 ( .A(n13093), .B(n12722), .Z(n12724) );
  XNOR U1525 ( .A(n13092), .B(n13420), .Z(n13087) );
  XNOR U1526 ( .A(n13824), .B(n14156), .Z(n13828) );
  XNOR U1527 ( .A(n14560), .B(n14892), .Z(n14564) );
  XNOR U1528 ( .A(n15296), .B(n15628), .Z(n15300) );
  XNOR U1529 ( .A(n16032), .B(n16364), .Z(n16036) );
  XNOR U1530 ( .A(n16768), .B(n17100), .Z(n16772) );
  XNOR U1531 ( .A(n17504), .B(n17836), .Z(n17508) );
  XNOR U1532 ( .A(n18240), .B(n18572), .Z(n18244) );
  XNOR U1533 ( .A(n18976), .B(n19308), .Z(n18980) );
  XNOR U1534 ( .A(n19712), .B(n20044), .Z(n19716) );
  XNOR U1535 ( .A(n20448), .B(n20780), .Z(n20452) );
  XNOR U1536 ( .A(n21184), .B(n21516), .Z(n21188) );
  XNOR U1537 ( .A(n23024), .B(n23356), .Z(n23028) );
  XNOR U1538 ( .A(n22298), .B(n22618), .Z(n22302) );
  XNOR U1539 ( .A(n26642), .B(n26962), .Z(n26646) );
  XNOR U1540 ( .A(n25982), .B(n26302), .Z(n25986) );
  XNOR U1541 ( .A(n25298), .B(n25618), .Z(n25302) );
  XNOR U1542 ( .A(n24590), .B(n24910), .Z(n24594) );
  XNOR U1543 ( .A(n23855), .B(n24175), .Z(n23859) );
  XNOR U1544 ( .A(n8508), .B(n8826), .Z(n8512) );
  XNOR U1545 ( .A(n9248), .B(n9569), .Z(n9252) );
  XNOR U1546 ( .A(n10000), .B(n10462), .Z(n10004) );
  XNOR U1547 ( .A(n10899), .B(n10528), .Z(n10530) );
  XNOR U1548 ( .A(n11268), .B(n10896), .Z(n10898) );
  XNOR U1549 ( .A(n11636), .B(n11265), .Z(n11267) );
  XNOR U1550 ( .A(n12004), .B(n11633), .Z(n11635) );
  XNOR U1551 ( .A(n12372), .B(n12001), .Z(n12003) );
  XNOR U1552 ( .A(n12740), .B(n12369), .Z(n12371) );
  XNOR U1553 ( .A(n13108), .B(n12737), .Z(n12739) );
  XNOR U1554 ( .A(n13476), .B(n13105), .Z(n13107) );
  XNOR U1555 ( .A(n13844), .B(n13473), .Z(n13475) );
  XNOR U1556 ( .A(n14212), .B(n13841), .Z(n13843) );
  XNOR U1557 ( .A(n14575), .B(n14889), .Z(n14583) );
  XNOR U1558 ( .A(n15311), .B(n15625), .Z(n15315) );
  XNOR U1559 ( .A(n16047), .B(n16361), .Z(n16051) );
  XNOR U1560 ( .A(n16783), .B(n17097), .Z(n16787) );
  XNOR U1561 ( .A(n17519), .B(n17833), .Z(n17523) );
  XNOR U1562 ( .A(n18255), .B(n18569), .Z(n18259) );
  XNOR U1563 ( .A(n18991), .B(n19305), .Z(n18995) );
  XNOR U1564 ( .A(n19727), .B(n20041), .Z(n19731) );
  XNOR U1565 ( .A(n20463), .B(n20777), .Z(n20467) );
  XNOR U1566 ( .A(n21199), .B(n21513), .Z(n21203) );
  XNOR U1567 ( .A(n23039), .B(n23353), .Z(n23043) );
  XNOR U1568 ( .A(n7382), .B(n7712), .Z(n7386) );
  XNOR U1569 ( .A(n6624), .B(n6968), .Z(n6628) );
  XNOR U1570 ( .A(n22313), .B(n22615), .Z(n22317) );
  XNOR U1571 ( .A(n27293), .B(n27595), .Z(n27297) );
  XNOR U1572 ( .A(n26657), .B(n26959), .Z(n26661) );
  XNOR U1573 ( .A(n25997), .B(n26299), .Z(n26001) );
  XNOR U1574 ( .A(n25313), .B(n25615), .Z(n25317) );
  XNOR U1575 ( .A(n24605), .B(n24907), .Z(n24609) );
  XNOR U1576 ( .A(n23870), .B(n24172), .Z(n23874) );
  XNOR U1577 ( .A(n8523), .B(n8823), .Z(n8527) );
  XNOR U1578 ( .A(n9263), .B(n9566), .Z(n9267) );
  XNOR U1579 ( .A(n10015), .B(n10456), .Z(n10019) );
  XNOR U1580 ( .A(n10914), .B(n10543), .Z(n10545) );
  XNOR U1581 ( .A(n11283), .B(n10911), .Z(n10913) );
  XNOR U1582 ( .A(n11651), .B(n11280), .Z(n11282) );
  XNOR U1583 ( .A(n12019), .B(n11648), .Z(n11650) );
  XNOR U1584 ( .A(n12387), .B(n12016), .Z(n12018) );
  XNOR U1585 ( .A(n12755), .B(n12384), .Z(n12386) );
  XNOR U1586 ( .A(n13123), .B(n12752), .Z(n12754) );
  XNOR U1587 ( .A(n13491), .B(n13120), .Z(n13122) );
  XNOR U1588 ( .A(n13859), .B(n13488), .Z(n13490) );
  XNOR U1589 ( .A(n14227), .B(n13856), .Z(n13858) );
  XNOR U1590 ( .A(n14595), .B(n14224), .Z(n14226) );
  XNOR U1591 ( .A(n14963), .B(n14592), .Z(n14594) );
  XNOR U1592 ( .A(n15331), .B(n14960), .Z(n14962) );
  XNOR U1593 ( .A(n15330), .B(n15622), .Z(n15325) );
  XNOR U1594 ( .A(n16062), .B(n16358), .Z(n16066) );
  XNOR U1595 ( .A(n16798), .B(n17094), .Z(n16802) );
  XNOR U1596 ( .A(n17534), .B(n17830), .Z(n17538) );
  XNOR U1597 ( .A(n18270), .B(n18566), .Z(n18274) );
  XNOR U1598 ( .A(n19006), .B(n19302), .Z(n19010) );
  XNOR U1599 ( .A(n19742), .B(n20038), .Z(n19746) );
  XNOR U1600 ( .A(n20478), .B(n20774), .Z(n20482) );
  XNOR U1601 ( .A(n21214), .B(n21510), .Z(n21218) );
  XNOR U1602 ( .A(n23054), .B(n23350), .Z(n23058) );
  XNOR U1603 ( .A(n7397), .B(n7709), .Z(n7401) );
  XNOR U1604 ( .A(n6639), .B(n6965), .Z(n6643) );
  XNOR U1605 ( .A(n5875), .B(n6229), .Z(n5879) );
  XNOR U1606 ( .A(n8161), .B(n8449), .Z(n8165) );
  XNOR U1607 ( .A(n22328), .B(n22612), .Z(n22332) );
  XNOR U1608 ( .A(n28508), .B(n28792), .Z(n28512) );
  XNOR U1609 ( .A(n27920), .B(n28204), .Z(n27924) );
  XNOR U1610 ( .A(n27308), .B(n27592), .Z(n27312) );
  XNOR U1611 ( .A(n26672), .B(n26956), .Z(n26676) );
  XNOR U1612 ( .A(n26012), .B(n26296), .Z(n26016) );
  XNOR U1613 ( .A(n25328), .B(n25612), .Z(n25332) );
  XNOR U1614 ( .A(n24620), .B(n24904), .Z(n24624) );
  XNOR U1615 ( .A(n23885), .B(n24169), .Z(n23889) );
  XNOR U1616 ( .A(n8910), .B(n9188), .Z(n8914) );
  XNOR U1617 ( .A(n9653), .B(n9940), .Z(n9657) );
  XNOR U1618 ( .A(n10555), .B(n10832), .Z(n10559) );
  XNOR U1619 ( .A(n11298), .B(n10926), .Z(n10928) );
  XNOR U1620 ( .A(n11666), .B(n11295), .Z(n11297) );
  XNOR U1621 ( .A(n12034), .B(n11663), .Z(n11665) );
  XNOR U1622 ( .A(n12402), .B(n12031), .Z(n12033) );
  XNOR U1623 ( .A(n12770), .B(n12399), .Z(n12401) );
  XNOR U1624 ( .A(n13138), .B(n12767), .Z(n12769) );
  XNOR U1625 ( .A(n13506), .B(n13135), .Z(n13137) );
  XNOR U1626 ( .A(n13874), .B(n13503), .Z(n13505) );
  XNOR U1627 ( .A(n14242), .B(n13871), .Z(n13873) );
  XNOR U1628 ( .A(n14610), .B(n14239), .Z(n14241) );
  XNOR U1629 ( .A(n14978), .B(n14607), .Z(n14609) );
  XNOR U1630 ( .A(n15346), .B(n14975), .Z(n14977) );
  XNOR U1631 ( .A(n15714), .B(n15343), .Z(n15345) );
  XNOR U1632 ( .A(n16082), .B(n15711), .Z(n15713) );
  XNOR U1633 ( .A(n16450), .B(n16079), .Z(n16081) );
  XNOR U1634 ( .A(n16813), .B(n17091), .Z(n16821) );
  XNOR U1635 ( .A(n17549), .B(n17827), .Z(n17553) );
  XNOR U1636 ( .A(n18285), .B(n18563), .Z(n18289) );
  XNOR U1637 ( .A(n19021), .B(n19299), .Z(n19025) );
  XNOR U1638 ( .A(n19757), .B(n20035), .Z(n19761) );
  XNOR U1639 ( .A(n20493), .B(n20771), .Z(n20497) );
  XNOR U1640 ( .A(n21229), .B(n21507), .Z(n21233) );
  XNOR U1641 ( .A(n23069), .B(n23347), .Z(n23073) );
  XNOR U1642 ( .A(n7794), .B(n8076), .Z(n7798) );
  XNOR U1643 ( .A(n7032), .B(n7335), .Z(n7036) );
  XNOR U1644 ( .A(n5890), .B(n6226), .Z(n5894) );
  XNOR U1645 ( .A(n22343), .B(n22609), .Z(n22347) );
  XNOR U1646 ( .A(n29087), .B(n29353), .Z(n29091) );
  XNOR U1647 ( .A(n28523), .B(n28789), .Z(n28527) );
  XNOR U1648 ( .A(n27935), .B(n28201), .Z(n27939) );
  XNOR U1649 ( .A(n27323), .B(n27589), .Z(n27327) );
  XNOR U1650 ( .A(n26687), .B(n26953), .Z(n26691) );
  XNOR U1651 ( .A(n26027), .B(n26293), .Z(n26031) );
  XNOR U1652 ( .A(n25343), .B(n25609), .Z(n25347) );
  XNOR U1653 ( .A(n24635), .B(n24901), .Z(n24639) );
  XNOR U1654 ( .A(n23900), .B(n24166), .Z(n23904) );
  XNOR U1655 ( .A(n5131), .B(n5485), .Z(n5135) );
  XNOR U1656 ( .A(n8553), .B(n8817), .Z(n8557) );
  XNOR U1657 ( .A(n9293), .B(n9560), .Z(n9297) );
  XNOR U1658 ( .A(n10045), .B(n10444), .Z(n10049) );
  XNOR U1659 ( .A(n10570), .B(n10829), .Z(n10574) );
  XNOR U1660 ( .A(n10938), .B(n11198), .Z(n10942) );
  XNOR U1661 ( .A(n11681), .B(n11310), .Z(n11312) );
  XNOR U1662 ( .A(n12049), .B(n11678), .Z(n11680) );
  XNOR U1663 ( .A(n12417), .B(n12046), .Z(n12048) );
  XNOR U1664 ( .A(n12785), .B(n12414), .Z(n12416) );
  XNOR U1665 ( .A(n13153), .B(n12782), .Z(n12784) );
  XNOR U1666 ( .A(n13521), .B(n13150), .Z(n13152) );
  XNOR U1667 ( .A(n13889), .B(n13518), .Z(n13520) );
  XNOR U1668 ( .A(n14257), .B(n13886), .Z(n13888) );
  XNOR U1669 ( .A(n14625), .B(n14254), .Z(n14256) );
  XNOR U1670 ( .A(n14993), .B(n14622), .Z(n14624) );
  XNOR U1671 ( .A(n15361), .B(n14990), .Z(n14992) );
  XNOR U1672 ( .A(n15729), .B(n15358), .Z(n15360) );
  XNOR U1673 ( .A(n16097), .B(n15726), .Z(n15728) );
  XNOR U1674 ( .A(n16465), .B(n16094), .Z(n16096) );
  XNOR U1675 ( .A(n16833), .B(n16462), .Z(n16464) );
  XNOR U1676 ( .A(n17201), .B(n16830), .Z(n16832) );
  XNOR U1677 ( .A(n17569), .B(n17198), .Z(n17200) );
  XNOR U1678 ( .A(n17568), .B(n17824), .Z(n17563) );
  XNOR U1679 ( .A(n18300), .B(n18560), .Z(n18304) );
  XNOR U1680 ( .A(n19036), .B(n19296), .Z(n19040) );
  XNOR U1681 ( .A(n19772), .B(n20032), .Z(n19776) );
  XNOR U1682 ( .A(n20508), .B(n20768), .Z(n20512) );
  XNOR U1683 ( .A(n21244), .B(n21504), .Z(n21248) );
  XNOR U1684 ( .A(n23084), .B(n23344), .Z(n23088) );
  XNOR U1685 ( .A(n7809), .B(n8073), .Z(n7813) );
  XNOR U1686 ( .A(n7047), .B(n7332), .Z(n7051) );
  XNOR U1687 ( .A(n6287), .B(n6593), .Z(n6291) );
  XNOR U1688 ( .A(n5523), .B(n5853), .Z(n5527) );
  XNOR U1689 ( .A(n22358), .B(n22606), .Z(n22362) );
  XNOR U1690 ( .A(n30158), .B(n30406), .Z(n30162) );
  XNOR U1691 ( .A(n29642), .B(n29890), .Z(n29646) );
  XNOR U1692 ( .A(n29102), .B(n29350), .Z(n29106) );
  XNOR U1693 ( .A(n28538), .B(n28786), .Z(n28542) );
  XNOR U1694 ( .A(n27950), .B(n28198), .Z(n27954) );
  XNOR U1695 ( .A(n27338), .B(n27586), .Z(n27342) );
  XNOR U1696 ( .A(n26702), .B(n26950), .Z(n26706) );
  XNOR U1697 ( .A(n26042), .B(n26290), .Z(n26046) );
  XNOR U1698 ( .A(n25358), .B(n25606), .Z(n25362) );
  XNOR U1699 ( .A(n24650), .B(n24898), .Z(n24654) );
  XNOR U1700 ( .A(n23915), .B(n24163), .Z(n23919) );
  XNOR U1701 ( .A(n4763), .B(n5112), .Z(n4767) );
  XNOR U1702 ( .A(n8568), .B(n8814), .Z(n8572) );
  XNOR U1703 ( .A(n9308), .B(n9557), .Z(n9312) );
  XNOR U1704 ( .A(n10060), .B(n10438), .Z(n10064) );
  XNOR U1705 ( .A(n10959), .B(n10588), .Z(n10590) );
  XNOR U1706 ( .A(n10953), .B(n11195), .Z(n10957) );
  XNOR U1707 ( .A(n12800), .B(n12429), .Z(n12431) );
  XNOR U1708 ( .A(n13168), .B(n12797), .Z(n12799) );
  XNOR U1709 ( .A(n13536), .B(n13165), .Z(n13167) );
  XNOR U1710 ( .A(n13904), .B(n13533), .Z(n13535) );
  XNOR U1711 ( .A(n14272), .B(n13901), .Z(n13903) );
  XNOR U1712 ( .A(n14640), .B(n14269), .Z(n14271) );
  XNOR U1713 ( .A(n15008), .B(n14637), .Z(n14639) );
  XNOR U1714 ( .A(n15376), .B(n15005), .Z(n15007) );
  XNOR U1715 ( .A(n15744), .B(n15373), .Z(n15375) );
  XNOR U1716 ( .A(n16112), .B(n15741), .Z(n15743) );
  XNOR U1717 ( .A(n16480), .B(n16109), .Z(n16111) );
  XNOR U1718 ( .A(n16848), .B(n16477), .Z(n16479) );
  XNOR U1719 ( .A(n17216), .B(n16845), .Z(n16847) );
  XNOR U1720 ( .A(n17584), .B(n17213), .Z(n17215) );
  XNOR U1721 ( .A(n17952), .B(n17581), .Z(n17583) );
  XNOR U1722 ( .A(n18320), .B(n17949), .Z(n17951) );
  XNOR U1723 ( .A(n18688), .B(n18317), .Z(n18319) );
  XNOR U1724 ( .A(n19051), .B(n19293), .Z(n19059) );
  XNOR U1725 ( .A(n19787), .B(n20029), .Z(n19791) );
  XNOR U1726 ( .A(n20523), .B(n20765), .Z(n20527) );
  XNOR U1727 ( .A(n21259), .B(n21501), .Z(n21263) );
  XNOR U1728 ( .A(n23099), .B(n23341), .Z(n23103) );
  XNOR U1729 ( .A(n7824), .B(n8070), .Z(n7828) );
  XNOR U1730 ( .A(n11695), .B(n11931), .Z(n11699) );
  XNOR U1731 ( .A(n12063), .B(n12299), .Z(n12067) );
  XNOR U1732 ( .A(n6684), .B(n6956), .Z(n6688) );
  XNOR U1733 ( .A(n5538), .B(n5850), .Z(n5542) );
  XNOR U1734 ( .A(n22373), .B(n22603), .Z(n22377) );
  XNOR U1735 ( .A(n30665), .B(n30895), .Z(n30669) );
  XNOR U1736 ( .A(n30173), .B(n30403), .Z(n30177) );
  XNOR U1737 ( .A(n29657), .B(n29887), .Z(n29661) );
  XNOR U1738 ( .A(n29117), .B(n29347), .Z(n29121) );
  XNOR U1739 ( .A(n28553), .B(n28783), .Z(n28557) );
  XNOR U1740 ( .A(n27965), .B(n28195), .Z(n27969) );
  XNOR U1741 ( .A(n27353), .B(n27583), .Z(n27357) );
  XNOR U1742 ( .A(n26717), .B(n26947), .Z(n26721) );
  XNOR U1743 ( .A(n26057), .B(n26287), .Z(n26061) );
  XNOR U1744 ( .A(n25373), .B(n25603), .Z(n25377) );
  XNOR U1745 ( .A(n24665), .B(n24895), .Z(n24669) );
  XNOR U1746 ( .A(n23930), .B(n24160), .Z(n23934) );
  XNOR U1747 ( .A(n4778), .B(n5109), .Z(n4782) );
  XNOR U1748 ( .A(n8955), .B(n9179), .Z(n8959) );
  XNOR U1749 ( .A(n9698), .B(n9931), .Z(n9702) );
  XNOR U1750 ( .A(n11711), .B(n11340), .Z(n11342) );
  XNOR U1751 ( .A(n12079), .B(n11708), .Z(n11710) );
  XNOR U1752 ( .A(n13919), .B(n13548), .Z(n13550) );
  XNOR U1753 ( .A(n14287), .B(n13916), .Z(n13918) );
  XNOR U1754 ( .A(n14655), .B(n14284), .Z(n14286) );
  XNOR U1755 ( .A(n15023), .B(n14652), .Z(n14654) );
  XNOR U1756 ( .A(n15391), .B(n15020), .Z(n15022) );
  XNOR U1757 ( .A(n15759), .B(n15388), .Z(n15390) );
  XNOR U1758 ( .A(n16127), .B(n15756), .Z(n15758) );
  XNOR U1759 ( .A(n16495), .B(n16124), .Z(n16126) );
  XNOR U1760 ( .A(n16863), .B(n16492), .Z(n16494) );
  XNOR U1761 ( .A(n17231), .B(n16860), .Z(n16862) );
  XNOR U1762 ( .A(n17599), .B(n17228), .Z(n17230) );
  XNOR U1763 ( .A(n17967), .B(n17596), .Z(n17598) );
  XNOR U1764 ( .A(n18335), .B(n17964), .Z(n17966) );
  XNOR U1765 ( .A(n18703), .B(n18332), .Z(n18334) );
  XNOR U1766 ( .A(n19071), .B(n18700), .Z(n18702) );
  XNOR U1767 ( .A(n19439), .B(n19068), .Z(n19070) );
  XNOR U1768 ( .A(n19807), .B(n19436), .Z(n19438) );
  XNOR U1769 ( .A(n19806), .B(n20026), .Z(n19801) );
  XNOR U1770 ( .A(n20538), .B(n20762), .Z(n20542) );
  XNOR U1771 ( .A(n21274), .B(n21498), .Z(n21278) );
  XNOR U1772 ( .A(n23114), .B(n23338), .Z(n23118) );
  XNOR U1773 ( .A(n7457), .B(n7697), .Z(n7461) );
  XNOR U1774 ( .A(n4019), .B(n4367), .Z(n4023) );
  XNOR U1775 ( .A(n10979), .B(n10608), .Z(n10610) );
  XNOR U1776 ( .A(n11348), .B(n10976), .Z(n10978) );
  XNOR U1777 ( .A(n11716), .B(n11345), .Z(n11347) );
  XNOR U1778 ( .A(n12446), .B(n12664), .Z(n12450) );
  XNOR U1779 ( .A(n12814), .B(n13032), .Z(n12818) );
  XNOR U1780 ( .A(n13182), .B(n13400), .Z(n13186) );
  XNOR U1781 ( .A(n5553), .B(n5847), .Z(n5557) );
  XNOR U1782 ( .A(n22388), .B(n22600), .Z(n22392) );
  XNOR U1783 ( .A(n31592), .B(n31975), .Z(n31596) );
  XNOR U1784 ( .A(n31148), .B(n31360), .Z(n31152) );
  XNOR U1785 ( .A(n30680), .B(n30892), .Z(n30684) );
  XNOR U1786 ( .A(n30188), .B(n30400), .Z(n30192) );
  XNOR U1787 ( .A(n29672), .B(n29884), .Z(n29676) );
  XNOR U1788 ( .A(n29132), .B(n29344), .Z(n29136) );
  XNOR U1789 ( .A(n28568), .B(n28780), .Z(n28572) );
  XNOR U1790 ( .A(n27980), .B(n28192), .Z(n27984) );
  XNOR U1791 ( .A(n27368), .B(n27580), .Z(n27372) );
  XNOR U1792 ( .A(n26732), .B(n26944), .Z(n26736) );
  XNOR U1793 ( .A(n26072), .B(n26284), .Z(n26076) );
  XNOR U1794 ( .A(n25388), .B(n25600), .Z(n25392) );
  XNOR U1795 ( .A(n24680), .B(n24892), .Z(n24684) );
  XNOR U1796 ( .A(n23945), .B(n24157), .Z(n23949) );
  XNOR U1797 ( .A(n6726), .B(n6947), .Z(n6727) );
  XNOR U1798 ( .A(n6322), .B(n6586), .Z(n6326) );
  XNOR U1799 ( .A(n4793), .B(n5106), .Z(n4797) );
  XNOR U1800 ( .A(n8230), .B(n8436), .Z(n8225) );
  XNOR U1801 ( .A(n8970), .B(n9176), .Z(n8974) );
  XNOR U1802 ( .A(n9713), .B(n9928), .Z(n9717) );
  XNOR U1803 ( .A(n13198), .B(n12827), .Z(n12829) );
  XNOR U1804 ( .A(n15038), .B(n14667), .Z(n14669) );
  XNOR U1805 ( .A(n15406), .B(n15035), .Z(n15037) );
  XNOR U1806 ( .A(n15774), .B(n15403), .Z(n15405) );
  XNOR U1807 ( .A(n16142), .B(n15771), .Z(n15773) );
  XNOR U1808 ( .A(n16510), .B(n16139), .Z(n16141) );
  XNOR U1809 ( .A(n16878), .B(n16507), .Z(n16509) );
  XNOR U1810 ( .A(n17246), .B(n16875), .Z(n16877) );
  XNOR U1811 ( .A(n17614), .B(n17243), .Z(n17245) );
  XNOR U1812 ( .A(n17982), .B(n17611), .Z(n17613) );
  XNOR U1813 ( .A(n18350), .B(n17979), .Z(n17981) );
  XNOR U1814 ( .A(n18718), .B(n18347), .Z(n18349) );
  XNOR U1815 ( .A(n19086), .B(n18715), .Z(n18717) );
  XNOR U1816 ( .A(n19454), .B(n19083), .Z(n19085) );
  XNOR U1817 ( .A(n19822), .B(n19451), .Z(n19453) );
  XNOR U1818 ( .A(n20190), .B(n19819), .Z(n19821) );
  XNOR U1819 ( .A(n20558), .B(n20187), .Z(n20189) );
  XNOR U1820 ( .A(n20926), .B(n20555), .Z(n20557) );
  XNOR U1821 ( .A(n21289), .B(n21495), .Z(n21297) );
  XNOR U1822 ( .A(n23129), .B(n23335), .Z(n23133) );
  XNOR U1823 ( .A(n7087), .B(n7324), .Z(n7095) );
  XNOR U1824 ( .A(n4034), .B(n4364), .Z(n4038) );
  XNOR U1825 ( .A(n3270), .B(n3624), .Z(n3274) );
  XNOR U1826 ( .A(n10994), .B(n10623), .Z(n10625) );
  XNOR U1827 ( .A(n10988), .B(n11188), .Z(n10992) );
  XNOR U1828 ( .A(n11731), .B(n11360), .Z(n11362) );
  XNOR U1829 ( .A(n12099), .B(n11728), .Z(n11730) );
  XNOR U1830 ( .A(n12467), .B(n12096), .Z(n12098) );
  XNOR U1831 ( .A(n12461), .B(n12661), .Z(n12465) );
  XNOR U1832 ( .A(n13565), .B(n13765), .Z(n13569) );
  XNOR U1833 ( .A(n13933), .B(n14133), .Z(n13937) );
  XNOR U1834 ( .A(n14301), .B(n14501), .Z(n14305) );
  XNOR U1835 ( .A(n5186), .B(n5474), .Z(n5190) );
  XNOR U1836 ( .A(n7491), .B(n7689), .Z(n7495) );
  XNOR U1837 ( .A(n22403), .B(n22597), .Z(n22407) );
  XNOR U1838 ( .A(n32190), .B(n32376), .Z(n32194) );
  XNOR U1839 ( .A(n31607), .B(n31972), .Z(n31611) );
  XNOR U1840 ( .A(n31163), .B(n31357), .Z(n31167) );
  XNOR U1841 ( .A(n30695), .B(n30889), .Z(n30699) );
  XNOR U1842 ( .A(n30203), .B(n30397), .Z(n30207) );
  XNOR U1843 ( .A(n29687), .B(n29881), .Z(n29691) );
  XNOR U1844 ( .A(n29147), .B(n29341), .Z(n29151) );
  XNOR U1845 ( .A(n28583), .B(n28777), .Z(n28587) );
  XNOR U1846 ( .A(n27995), .B(n28189), .Z(n27999) );
  XNOR U1847 ( .A(n27383), .B(n27577), .Z(n27387) );
  XNOR U1848 ( .A(n26747), .B(n26941), .Z(n26751) );
  XNOR U1849 ( .A(n26087), .B(n26281), .Z(n26091) );
  XNOR U1850 ( .A(n25403), .B(n25597), .Z(n25407) );
  XNOR U1851 ( .A(n24695), .B(n24889), .Z(n24699) );
  XNOR U1852 ( .A(n23960), .B(n24154), .Z(n23964) );
  XNOR U1853 ( .A(n6356), .B(n6578), .Z(n6360) );
  XNOR U1854 ( .A(n5955), .B(n6213), .Z(n5959) );
  XNOR U1855 ( .A(n4426), .B(n4732), .Z(n4430) );
  XNOR U1856 ( .A(n6380), .B(n6572), .Z(n6384) );
  XNOR U1857 ( .A(n8240), .B(n8432), .Z(n8244) );
  XNOR U1858 ( .A(n8987), .B(n9172), .Z(n8988) );
  XNOR U1859 ( .A(n9728), .B(n9925), .Z(n9736) );
  XNOR U1860 ( .A(n14317), .B(n13946), .Z(n13948) );
  XNOR U1861 ( .A(n16157), .B(n15786), .Z(n15788) );
  XNOR U1862 ( .A(n16525), .B(n16154), .Z(n16156) );
  XNOR U1863 ( .A(n16893), .B(n16522), .Z(n16524) );
  XNOR U1864 ( .A(n17261), .B(n16890), .Z(n16892) );
  XNOR U1865 ( .A(n17629), .B(n17258), .Z(n17260) );
  XNOR U1866 ( .A(n17997), .B(n17626), .Z(n17628) );
  XNOR U1867 ( .A(n18365), .B(n17994), .Z(n17996) );
  XNOR U1868 ( .A(n18733), .B(n18362), .Z(n18364) );
  XNOR U1869 ( .A(n19101), .B(n18730), .Z(n18732) );
  XNOR U1870 ( .A(n19469), .B(n19098), .Z(n19100) );
  XNOR U1871 ( .A(n19837), .B(n19466), .Z(n19468) );
  XNOR U1872 ( .A(n20205), .B(n19834), .Z(n19836) );
  XNOR U1873 ( .A(n20573), .B(n20202), .Z(n20204) );
  XNOR U1874 ( .A(n20941), .B(n20570), .Z(n20572) );
  XNOR U1875 ( .A(n21309), .B(n20938), .Z(n20940) );
  XNOR U1876 ( .A(n21677), .B(n21306), .Z(n21308) );
  XNOR U1877 ( .A(n22045), .B(n21674), .Z(n21676) );
  XNOR U1878 ( .A(n22044), .B(n22228), .Z(n22039) );
  XNOR U1879 ( .A(n23144), .B(n23332), .Z(n23148) );
  XNOR U1880 ( .A(n7125), .B(n7316), .Z(n7120) );
  XNOR U1881 ( .A(n5597), .B(n5837), .Z(n5601) );
  XNOR U1882 ( .A(n3667), .B(n3991), .Z(n3671) );
  XNOR U1883 ( .A(n2903), .B(n3251), .Z(n2907) );
  XNOR U1884 ( .A(n5624), .B(n5831), .Z(n5625) );
  XNOR U1885 ( .A(n11003), .B(n11185), .Z(n11007) );
  XNOR U1886 ( .A(n11746), .B(n11375), .Z(n11377) );
  XNOR U1887 ( .A(n12114), .B(n11743), .Z(n11745) );
  XNOR U1888 ( .A(n13218), .B(n12847), .Z(n12849) );
  XNOR U1889 ( .A(n13586), .B(n13215), .Z(n13217) );
  XNOR U1890 ( .A(n13580), .B(n13762), .Z(n13584) );
  XNOR U1891 ( .A(n14684), .B(n14866), .Z(n14688) );
  XNOR U1892 ( .A(n15052), .B(n15234), .Z(n15056) );
  XNOR U1893 ( .A(n15420), .B(n15602), .Z(n15424) );
  XNOR U1894 ( .A(n10640), .B(n10815), .Z(n10644) );
  XNOR U1895 ( .A(n12481), .B(n12657), .Z(n12485) );
  XNOR U1896 ( .A(n32944), .B(n33115), .Z(n32948) );
  XNOR U1897 ( .A(n32588), .B(n32756), .Z(n32592) );
  XNOR U1898 ( .A(n32205), .B(n32373), .Z(n32209) );
  XNOR U1899 ( .A(n31622), .B(n31969), .Z(n31626) );
  XNOR U1900 ( .A(n31178), .B(n31354), .Z(n31182) );
  XNOR U1901 ( .A(n30710), .B(n30886), .Z(n30714) );
  XNOR U1902 ( .A(n30218), .B(n30394), .Z(n30222) );
  XNOR U1903 ( .A(n29702), .B(n29878), .Z(n29706) );
  XNOR U1904 ( .A(n29162), .B(n29338), .Z(n29166) );
  XNOR U1905 ( .A(n28598), .B(n28774), .Z(n28602) );
  XNOR U1906 ( .A(n28010), .B(n28186), .Z(n28014) );
  XNOR U1907 ( .A(n27398), .B(n27574), .Z(n27402) );
  XNOR U1908 ( .A(n26762), .B(n26938), .Z(n26766) );
  XNOR U1909 ( .A(n26102), .B(n26278), .Z(n26106) );
  XNOR U1910 ( .A(n25418), .B(n25594), .Z(n25422) );
  XNOR U1911 ( .A(n24710), .B(n24886), .Z(n24714) );
  XNOR U1912 ( .A(n23975), .B(n24151), .Z(n23979) );
  XNOR U1913 ( .A(n5989), .B(n6205), .Z(n5997) );
  XNOR U1914 ( .A(n5206), .B(n5470), .Z(n5214) );
  XNOR U1915 ( .A(n4441), .B(n4729), .Z(n4445) );
  XNOR U1916 ( .A(n6767), .B(n6937), .Z(n6771) );
  XNOR U1917 ( .A(n7510), .B(n7684), .Z(n7514) );
  XNOR U1918 ( .A(n8259), .B(n8429), .Z(n8254) );
  XNOR U1919 ( .A(n8999), .B(n9169), .Z(n9003) );
  XNOR U1920 ( .A(n10651), .B(n10122), .Z(n10124) );
  XNOR U1921 ( .A(n15436), .B(n15065), .Z(n15067) );
  XNOR U1922 ( .A(n17276), .B(n16905), .Z(n16907) );
  XNOR U1923 ( .A(n17644), .B(n17273), .Z(n17275) );
  XNOR U1924 ( .A(n18012), .B(n17641), .Z(n17643) );
  XNOR U1925 ( .A(n18380), .B(n18009), .Z(n18011) );
  XNOR U1926 ( .A(n18748), .B(n18377), .Z(n18379) );
  XNOR U1927 ( .A(n19116), .B(n18745), .Z(n18747) );
  XNOR U1928 ( .A(n19484), .B(n19113), .Z(n19115) );
  XNOR U1929 ( .A(n19852), .B(n19481), .Z(n19483) );
  XNOR U1930 ( .A(n20220), .B(n19849), .Z(n19851) );
  XNOR U1931 ( .A(n20588), .B(n20217), .Z(n20219) );
  XNOR U1932 ( .A(n20956), .B(n20585), .Z(n20587) );
  XNOR U1933 ( .A(n21324), .B(n20953), .Z(n20955) );
  XNOR U1934 ( .A(n21692), .B(n21321), .Z(n21323) );
  XNOR U1935 ( .A(n22060), .B(n21689), .Z(n21691) );
  XNOR U1936 ( .A(n22428), .B(n22057), .Z(n22059) );
  XNOR U1937 ( .A(n22796), .B(n22425), .Z(n22427) );
  XNOR U1938 ( .A(n23164), .B(n22793), .Z(n22795) );
  XNOR U1939 ( .A(n23163), .B(n23329), .Z(n23158) );
  XNOR U1940 ( .A(n5230), .B(n5464), .Z(n5234) );
  XNOR U1941 ( .A(n4465), .B(n4723), .Z(n4469) );
  XNOR U1942 ( .A(n2918), .B(n3248), .Z(n2922) );
  XNOR U1943 ( .A(n4871), .B(n5088), .Z(n4875) );
  XNOR U1944 ( .A(n11018), .B(n11182), .Z(n11022) );
  XNOR U1945 ( .A(n13233), .B(n12862), .Z(n12864) );
  XNOR U1946 ( .A(n14337), .B(n13966), .Z(n13968) );
  XNOR U1947 ( .A(n14705), .B(n14334), .Z(n14336) );
  XNOR U1948 ( .A(n14699), .B(n14863), .Z(n14703) );
  XNOR U1949 ( .A(n15803), .B(n15967), .Z(n15807) );
  XNOR U1950 ( .A(n16171), .B(n16335), .Z(n16175) );
  XNOR U1951 ( .A(n16539), .B(n16703), .Z(n16543) );
  XNOR U1952 ( .A(n3305), .B(n3617), .Z(n3309) );
  XNOR U1953 ( .A(n2157), .B(n2506), .Z(n2161) );
  XNOR U1954 ( .A(n5641), .B(n5827), .Z(n5649) );
  XNOR U1955 ( .A(n4115), .B(n4346), .Z(n4116) );
  XNOR U1956 ( .A(n10655), .B(n10812), .Z(n10659) );
  XNOR U1957 ( .A(n11760), .B(n11918), .Z(n11764) );
  XNOR U1958 ( .A(n12496), .B(n12654), .Z(n12500) );
  XNOR U1959 ( .A(n13600), .B(n13758), .Z(n13604) );
  XNOR U1960 ( .A(n33294), .B(n33444), .Z(n33298) );
  XNOR U1961 ( .A(n32959), .B(n33112), .Z(n32963) );
  XNOR U1962 ( .A(n32603), .B(n32753), .Z(n32607) );
  XNOR U1963 ( .A(n32220), .B(n32370), .Z(n32224) );
  XNOR U1964 ( .A(n31637), .B(n31966), .Z(n31641) );
  XNOR U1965 ( .A(n31193), .B(n31351), .Z(n31197) );
  XNOR U1966 ( .A(n30725), .B(n30883), .Z(n30729) );
  XNOR U1967 ( .A(n30233), .B(n30391), .Z(n30237) );
  XNOR U1968 ( .A(n29717), .B(n29875), .Z(n29721) );
  XNOR U1969 ( .A(n29177), .B(n29335), .Z(n29181) );
  XNOR U1970 ( .A(n28613), .B(n28771), .Z(n28617) );
  XNOR U1971 ( .A(n28025), .B(n28183), .Z(n28029) );
  XNOR U1972 ( .A(n27413), .B(n27571), .Z(n27417) );
  XNOR U1973 ( .A(n26777), .B(n26935), .Z(n26781) );
  XNOR U1974 ( .A(n26117), .B(n26275), .Z(n26121) );
  XNOR U1975 ( .A(n25433), .B(n25591), .Z(n25437) );
  XNOR U1976 ( .A(n24725), .B(n24883), .Z(n24729) );
  XNOR U1977 ( .A(n23990), .B(n24148), .Z(n23994) );
  XNOR U1978 ( .A(n4900), .B(n5081), .Z(n4904) );
  XNOR U1979 ( .A(n4074), .B(n4356), .Z(n4082) );
  XNOR U1980 ( .A(n6784), .B(n6933), .Z(n6785) );
  XNOR U1981 ( .A(n7525), .B(n7681), .Z(n7533) );
  XNOR U1982 ( .A(n8269), .B(n8425), .Z(n8273) );
  XNOR U1983 ( .A(n9016), .B(n9165), .Z(n9017) );
  XNOR U1984 ( .A(n9757), .B(n9917), .Z(n9765) );
  XNOR U1985 ( .A(n16555), .B(n16184), .Z(n16186) );
  XNOR U1986 ( .A(n18395), .B(n18024), .Z(n18026) );
  XNOR U1987 ( .A(n18763), .B(n18392), .Z(n18394) );
  XNOR U1988 ( .A(n19131), .B(n18760), .Z(n18762) );
  XNOR U1989 ( .A(n19499), .B(n19128), .Z(n19130) );
  XNOR U1990 ( .A(n19867), .B(n19496), .Z(n19498) );
  XNOR U1991 ( .A(n20235), .B(n19864), .Z(n19866) );
  XNOR U1992 ( .A(n20603), .B(n20232), .Z(n20234) );
  XNOR U1993 ( .A(n20971), .B(n20600), .Z(n20602) );
  XNOR U1994 ( .A(n21339), .B(n20968), .Z(n20970) );
  XNOR U1995 ( .A(n21707), .B(n21336), .Z(n21338) );
  XNOR U1996 ( .A(n22075), .B(n21704), .Z(n21706) );
  XNOR U1997 ( .A(n22443), .B(n22072), .Z(n22074) );
  XNOR U1998 ( .A(n22811), .B(n22440), .Z(n22442) );
  XNOR U1999 ( .A(n23179), .B(n22808), .Z(n22810) );
  XNOR U2000 ( .A(n23173), .B(n23325), .Z(n23177) );
  XNOR U2001 ( .A(n4144), .B(n4339), .Z(n4145) );
  XNOR U2002 ( .A(n4480), .B(n4720), .Z(n4488) );
  XNOR U2003 ( .A(n3716), .B(n3980), .Z(n3720) );
  XNOR U2004 ( .A(n6042), .B(n6192), .Z(n6046) );
  XNOR U2005 ( .A(n11033), .B(n11179), .Z(n11037) );
  XNOR U2006 ( .A(n12512), .B(n12141), .Z(n12143) );
  XNOR U2007 ( .A(n14352), .B(n13981), .Z(n13983) );
  XNOR U2008 ( .A(n15456), .B(n15085), .Z(n15087) );
  XNOR U2009 ( .A(n15824), .B(n15453), .Z(n15455) );
  XNOR U2010 ( .A(n15818), .B(n15964), .Z(n15822) );
  XNOR U2011 ( .A(n16922), .B(n17068), .Z(n16926) );
  XNOR U2012 ( .A(n17290), .B(n17436), .Z(n17294) );
  XNOR U2013 ( .A(n17658), .B(n17804), .Z(n17662) );
  XNOR U2014 ( .A(n2555), .B(n2874), .Z(n2559) );
  XNOR U2015 ( .A(n1790), .B(n2132), .Z(n1794) );
  XNOR U2016 ( .A(n4509), .B(n4713), .Z(n4517) );
  XNOR U2017 ( .A(n3745), .B(n3973), .Z(n3749) );
  XNOR U2018 ( .A(n2984), .B(n3233), .Z(n2985) );
  XNOR U2019 ( .A(n4173), .B(n4332), .Z(n4174) );
  XNOR U2020 ( .A(n10670), .B(n10809), .Z(n10674) );
  XNOR U2021 ( .A(n11775), .B(n11915), .Z(n11779) );
  XNOR U2022 ( .A(n12879), .B(n13019), .Z(n12883) );
  XNOR U2023 ( .A(n13615), .B(n13755), .Z(n13619) );
  XNOR U2024 ( .A(n14719), .B(n14859), .Z(n14723) );
  XNOR U2025 ( .A(n33904), .B(n34039), .Z(n33908) );
  XNOR U2026 ( .A(n33620), .B(n33752), .Z(n33624) );
  XNOR U2027 ( .A(n33309), .B(n33441), .Z(n33313) );
  XNOR U2028 ( .A(n32974), .B(n33109), .Z(n32978) );
  XNOR U2029 ( .A(n32618), .B(n32750), .Z(n32622) );
  XNOR U2030 ( .A(n32235), .B(n32367), .Z(n32239) );
  XNOR U2031 ( .A(n31652), .B(n31963), .Z(n31656) );
  XNOR U2032 ( .A(n31208), .B(n31348), .Z(n31212) );
  XNOR U2033 ( .A(n30740), .B(n30880), .Z(n30744) );
  XNOR U2034 ( .A(n30248), .B(n30388), .Z(n30252) );
  XNOR U2035 ( .A(n29732), .B(n29872), .Z(n29736) );
  XNOR U2036 ( .A(n29192), .B(n29332), .Z(n29196) );
  XNOR U2037 ( .A(n28628), .B(n28768), .Z(n28632) );
  XNOR U2038 ( .A(n28040), .B(n28180), .Z(n28044) );
  XNOR U2039 ( .A(n27428), .B(n27568), .Z(n27432) );
  XNOR U2040 ( .A(n26792), .B(n26932), .Z(n26796) );
  XNOR U2041 ( .A(n26132), .B(n26272), .Z(n26136) );
  XNOR U2042 ( .A(n25448), .B(n25588), .Z(n25452) );
  XNOR U2043 ( .A(n24740), .B(n24880), .Z(n24744) );
  XNOR U2044 ( .A(n24005), .B(n24145), .Z(n24009) );
  XNOR U2045 ( .A(n5302), .B(n5448), .Z(n5297) );
  XNOR U2046 ( .A(n2943), .B(n3243), .Z(n2951) );
  XNOR U2047 ( .A(n4934), .B(n5073), .Z(n4938) );
  XNOR U2048 ( .A(n7539), .B(n7677), .Z(n7543) );
  XNOR U2049 ( .A(n8288), .B(n8422), .Z(n8283) );
  XNOR U2050 ( .A(n9028), .B(n9162), .Z(n9032) );
  XNOR U2051 ( .A(n10681), .B(n10151), .Z(n10153) );
  XNOR U2052 ( .A(n17674), .B(n17303), .Z(n17305) );
  XNOR U2053 ( .A(n19514), .B(n19143), .Z(n19145) );
  XNOR U2054 ( .A(n19882), .B(n19511), .Z(n19513) );
  XNOR U2055 ( .A(n20250), .B(n19879), .Z(n19881) );
  XNOR U2056 ( .A(n20618), .B(n20247), .Z(n20249) );
  XNOR U2057 ( .A(n20986), .B(n20615), .Z(n20617) );
  XNOR U2058 ( .A(n21354), .B(n20983), .Z(n20985) );
  XNOR U2059 ( .A(n21722), .B(n21351), .Z(n21353) );
  XNOR U2060 ( .A(n22090), .B(n21719), .Z(n21721) );
  XNOR U2061 ( .A(n22458), .B(n22087), .Z(n22089) );
  XNOR U2062 ( .A(n22826), .B(n22455), .Z(n22457) );
  XNOR U2063 ( .A(n23194), .B(n22823), .Z(n22825) );
  XNOR U2064 ( .A(n23188), .B(n23322), .Z(n23192) );
  XNOR U2065 ( .A(n4538), .B(n4706), .Z(n4546) );
  XNOR U2066 ( .A(n3774), .B(n3966), .Z(n3778) );
  XNOR U2067 ( .A(n3013), .B(n3226), .Z(n3014) );
  XNOR U2068 ( .A(n3349), .B(n3607), .Z(n3357) );
  XNOR U2069 ( .A(n2584), .B(n2867), .Z(n2588) );
  XNOR U2070 ( .A(n1822), .B(n2125), .Z(n1823) );
  XNOR U2071 ( .A(n6801), .B(n6929), .Z(n6809) );
  XNOR U2072 ( .A(n11048), .B(n11176), .Z(n11052) );
  XNOR U2073 ( .A(n12527), .B(n12156), .Z(n12158) );
  XNOR U2074 ( .A(n13631), .B(n13260), .Z(n13262) );
  XNOR U2075 ( .A(n15471), .B(n15100), .Z(n15102) );
  XNOR U2076 ( .A(n16575), .B(n16204), .Z(n16206) );
  XNOR U2077 ( .A(n16943), .B(n16572), .Z(n16574) );
  XNOR U2078 ( .A(n16937), .B(n17065), .Z(n16941) );
  XNOR U2079 ( .A(n18041), .B(n18169), .Z(n18045) );
  XNOR U2080 ( .A(n18409), .B(n18537), .Z(n18413) );
  XNOR U2081 ( .A(n18777), .B(n18905), .Z(n18781) );
  XNOR U2082 ( .A(n1805), .B(n2129), .Z(n1809) );
  XNOR U2083 ( .A(n1041), .B(n1389), .Z(n1045) );
  XNOR U2084 ( .A(n3378), .B(n3600), .Z(n3386) );
  XNOR U2085 ( .A(n2613), .B(n2860), .Z(n2617) );
  XNOR U2086 ( .A(n1851), .B(n2118), .Z(n1852) );
  XNOR U2087 ( .A(n3803), .B(n3959), .Z(n3807) );
  XNOR U2088 ( .A(n3042), .B(n3219), .Z(n3043) );
  XNOR U2089 ( .A(n6436), .B(n6559), .Z(n6437) );
  XNOR U2090 ( .A(n10685), .B(n10806), .Z(n10689) );
  XNOR U2091 ( .A(n11790), .B(n11912), .Z(n11794) );
  XNOR U2092 ( .A(n12894), .B(n13016), .Z(n12898) );
  XNOR U2093 ( .A(n13998), .B(n14120), .Z(n14002) );
  XNOR U2094 ( .A(n14734), .B(n14856), .Z(n14738) );
  XNOR U2095 ( .A(n15838), .B(n15960), .Z(n15842) );
  XNOR U2096 ( .A(n34182), .B(n34296), .Z(n34186) );
  XNOR U2097 ( .A(n33919), .B(n34036), .Z(n33923) );
  XNOR U2098 ( .A(n33635), .B(n33749), .Z(n33639) );
  XNOR U2099 ( .A(n33324), .B(n33438), .Z(n33328) );
  XNOR U2100 ( .A(n32989), .B(n33106), .Z(n32993) );
  XNOR U2101 ( .A(n32633), .B(n32747), .Z(n32637) );
  XNOR U2102 ( .A(n32250), .B(n32364), .Z(n32254) );
  XNOR U2103 ( .A(n31667), .B(n31960), .Z(n31671) );
  XNOR U2104 ( .A(n31223), .B(n31345), .Z(n31227) );
  XNOR U2105 ( .A(n30755), .B(n30877), .Z(n30759) );
  XNOR U2106 ( .A(n30263), .B(n30385), .Z(n30267) );
  XNOR U2107 ( .A(n29747), .B(n29869), .Z(n29751) );
  XNOR U2108 ( .A(n29207), .B(n29329), .Z(n29211) );
  XNOR U2109 ( .A(n28643), .B(n28765), .Z(n28647) );
  XNOR U2110 ( .A(n28055), .B(n28177), .Z(n28059) );
  XNOR U2111 ( .A(n27443), .B(n27565), .Z(n27447) );
  XNOR U2112 ( .A(n26807), .B(n26929), .Z(n26811) );
  XNOR U2113 ( .A(n26147), .B(n26269), .Z(n26151) );
  XNOR U2114 ( .A(n25463), .B(n25585), .Z(n25467) );
  XNOR U2115 ( .A(n24755), .B(n24877), .Z(n24759) );
  XNOR U2116 ( .A(n24020), .B(n24142), .Z(n24024) );
  XNOR U2117 ( .A(n3827), .B(n3953), .Z(n3831) );
  XNOR U2118 ( .A(n4579), .B(n4696), .Z(n4580) );
  XNOR U2119 ( .A(n5322), .B(n5442), .Z(n5330) );
  XNOR U2120 ( .A(n8298), .B(n8418), .Z(n8302) );
  XNOR U2121 ( .A(n9045), .B(n9158), .Z(n9046) );
  XNOR U2122 ( .A(n9786), .B(n9909), .Z(n9794) );
  XNOR U2123 ( .A(n18793), .B(n18422), .Z(n18424) );
  XNOR U2124 ( .A(n20633), .B(n20262), .Z(n20264) );
  XNOR U2125 ( .A(n21001), .B(n20630), .Z(n20632) );
  XNOR U2126 ( .A(n21369), .B(n20998), .Z(n21000) );
  XNOR U2127 ( .A(n21737), .B(n21366), .Z(n21368) );
  XNOR U2128 ( .A(n22105), .B(n21734), .Z(n21736) );
  XNOR U2129 ( .A(n22473), .B(n22102), .Z(n22104) );
  XNOR U2130 ( .A(n22841), .B(n22470), .Z(n22472) );
  XNOR U2131 ( .A(n23209), .B(n22838), .Z(n22840) );
  XNOR U2132 ( .A(n23203), .B(n23319), .Z(n23207) );
  XNOR U2133 ( .A(n3071), .B(n3212), .Z(n3072) );
  XNOR U2134 ( .A(n3407), .B(n3593), .Z(n3415) );
  XNOR U2135 ( .A(n2642), .B(n2853), .Z(n2646) );
  XNOR U2136 ( .A(n1880), .B(n2111), .Z(n1881) );
  XNOR U2137 ( .A(n2216), .B(n2493), .Z(n2224) );
  XNOR U2138 ( .A(n1452), .B(n1752), .Z(n1456) );
  XNOR U2139 ( .A(n691), .B(n1012), .Z(n692) );
  XNOR U2140 ( .A(n7563), .B(n7673), .Z(n7558) );
  XNOR U2141 ( .A(n11063), .B(n11173), .Z(n11067) );
  XNOR U2142 ( .A(n12542), .B(n12171), .Z(n12173) );
  XNOR U2143 ( .A(n13646), .B(n13275), .Z(n13277) );
  XNOR U2144 ( .A(n14750), .B(n14379), .Z(n14381) );
  XNOR U2145 ( .A(n16590), .B(n16219), .Z(n16221) );
  XNOR U2146 ( .A(n17694), .B(n17323), .Z(n17325) );
  XNOR U2147 ( .A(n18062), .B(n17691), .Z(n17693) );
  XNOR U2148 ( .A(n18056), .B(n18166), .Z(n18060) );
  XNOR U2149 ( .A(n19160), .B(n19270), .Z(n19164) );
  XNOR U2150 ( .A(n19528), .B(n19638), .Z(n19532) );
  XNOR U2151 ( .A(n19896), .B(n20006), .Z(n19900) );
  XNOR U2152 ( .A(n1056), .B(n1386), .Z(n1064) );
  XNOR U2153 ( .A(n2245), .B(n2486), .Z(n2253) );
  XNOR U2154 ( .A(n1481), .B(n1745), .Z(n1485) );
  XNOR U2155 ( .A(n720), .B(n1005), .Z(n721) );
  XNOR U2156 ( .A(n3436), .B(n3586), .Z(n3444) );
  XNOR U2157 ( .A(n2671), .B(n2846), .Z(n2675) );
  XNOR U2158 ( .A(n1909), .B(n2104), .Z(n1910) );
  XNOR U2159 ( .A(n7188), .B(n7299), .Z(n7192) );
  XNOR U2160 ( .A(n10700), .B(n10803), .Z(n10704) );
  XNOR U2161 ( .A(n11805), .B(n11909), .Z(n11809) );
  XNOR U2162 ( .A(n12909), .B(n13013), .Z(n12913) );
  XNOR U2163 ( .A(n14013), .B(n14117), .Z(n14017) );
  XNOR U2164 ( .A(n15117), .B(n15221), .Z(n15121) );
  XNOR U2165 ( .A(n15853), .B(n15957), .Z(n15857) );
  XNOR U2166 ( .A(n16957), .B(n17061), .Z(n16961) );
  XNOR U2167 ( .A(n34648), .B(n34747), .Z(n34652) );
  XNOR U2168 ( .A(n34436), .B(n34532), .Z(n34440) );
  XNOR U2169 ( .A(n34197), .B(n34293), .Z(n34201) );
  XNOR U2170 ( .A(n33934), .B(n34033), .Z(n33938) );
  XNOR U2171 ( .A(n33650), .B(n33746), .Z(n33654) );
  XNOR U2172 ( .A(n33339), .B(n33435), .Z(n33343) );
  XNOR U2173 ( .A(n33004), .B(n33103), .Z(n33008) );
  XNOR U2174 ( .A(n32648), .B(n32744), .Z(n32652) );
  XNOR U2175 ( .A(n32265), .B(n32361), .Z(n32269) );
  XNOR U2176 ( .A(n31682), .B(n31957), .Z(n31686) );
  XNOR U2177 ( .A(n31238), .B(n31342), .Z(n31242) );
  XNOR U2178 ( .A(n30770), .B(n30874), .Z(n30774) );
  XNOR U2179 ( .A(n30278), .B(n30382), .Z(n30282) );
  XNOR U2180 ( .A(n29762), .B(n29866), .Z(n29766) );
  XNOR U2181 ( .A(n29222), .B(n29326), .Z(n29226) );
  XNOR U2182 ( .A(n28658), .B(n28762), .Z(n28662) );
  XNOR U2183 ( .A(n28070), .B(n28174), .Z(n28074) );
  XNOR U2184 ( .A(n27458), .B(n27562), .Z(n27462) );
  XNOR U2185 ( .A(n26822), .B(n26926), .Z(n26826) );
  XNOR U2186 ( .A(n26162), .B(n26266), .Z(n26166) );
  XNOR U2187 ( .A(n25478), .B(n25582), .Z(n25482) );
  XNOR U2188 ( .A(n24770), .B(n24874), .Z(n24774) );
  XNOR U2189 ( .A(n24035), .B(n24139), .Z(n24039) );
  XNOR U2190 ( .A(n4591), .B(n4693), .Z(n4595) );
  XNOR U2191 ( .A(n5336), .B(n5438), .Z(n5340) );
  XNOR U2192 ( .A(n6085), .B(n6183), .Z(n6080) );
  XNOR U2193 ( .A(n9057), .B(n9155), .Z(n9061) );
  XNOR U2194 ( .A(n10711), .B(n10180), .Z(n10182) );
  XNOR U2195 ( .A(n21752), .B(n21381), .Z(n21383) );
  XNOR U2196 ( .A(n22120), .B(n21749), .Z(n21751) );
  XNOR U2197 ( .A(n22488), .B(n22117), .Z(n22119) );
  XNOR U2198 ( .A(n22856), .B(n22485), .Z(n22487) );
  XNOR U2199 ( .A(n23224), .B(n22853), .Z(n22855) );
  XNOR U2200 ( .A(n23218), .B(n23316), .Z(n23222) );
  XNOR U2201 ( .A(n3465), .B(n3579), .Z(n3473) );
  XNOR U2202 ( .A(n2700), .B(n2839), .Z(n2704) );
  XNOR U2203 ( .A(n1938), .B(n2097), .Z(n1939) );
  XNOR U2204 ( .A(n2274), .B(n2479), .Z(n2282) );
  XNOR U2205 ( .A(n1510), .B(n1738), .Z(n1514) );
  XNOR U2206 ( .A(n749), .B(n998), .Z(n750) );
  XNOR U2207 ( .A(n1085), .B(n1379), .Z(n1093) );
  XNOR U2208 ( .A(n2724), .B(n2833), .Z(n2728) );
  XNOR U2209 ( .A(n8320), .B(n8413), .Z(n8321) );
  XNOR U2210 ( .A(n11078), .B(n11170), .Z(n11082) );
  XNOR U2211 ( .A(n12557), .B(n12186), .Z(n12188) );
  XNOR U2212 ( .A(n13661), .B(n13290), .Z(n13292) );
  XNOR U2213 ( .A(n14765), .B(n14394), .Z(n14396) );
  XNOR U2214 ( .A(n15869), .B(n15498), .Z(n15500) );
  XNOR U2215 ( .A(n17709), .B(n17338), .Z(n17340) );
  XNOR U2216 ( .A(n18813), .B(n18442), .Z(n18444) );
  XNOR U2217 ( .A(n19181), .B(n18810), .Z(n18812) );
  XNOR U2218 ( .A(n19175), .B(n19267), .Z(n19179) );
  XNOR U2219 ( .A(n20279), .B(n20371), .Z(n20283) );
  XNOR U2220 ( .A(n1114), .B(n1372), .Z(n1122) );
  XNOR U2221 ( .A(n2303), .B(n2472), .Z(n2311) );
  XNOR U2222 ( .A(n1539), .B(n1731), .Z(n1543) );
  XNOR U2223 ( .A(n778), .B(n991), .Z(n779) );
  XNOR U2224 ( .A(n1967), .B(n2090), .Z(n1968) );
  XNOR U2225 ( .A(n7950), .B(n8040), .Z(n7954) );
  XNOR U2226 ( .A(n10715), .B(n10800), .Z(n10719) );
  XNOR U2227 ( .A(n11820), .B(n11906), .Z(n11824) );
  XNOR U2228 ( .A(n12924), .B(n13010), .Z(n12928) );
  XNOR U2229 ( .A(n14028), .B(n14114), .Z(n14032) );
  XNOR U2230 ( .A(n15132), .B(n15218), .Z(n15136) );
  XNOR U2231 ( .A(n16236), .B(n16322), .Z(n16240) );
  XNOR U2232 ( .A(n16972), .B(n17058), .Z(n16976) );
  XNOR U2233 ( .A(n18076), .B(n18162), .Z(n18080) );
  XNOR U2234 ( .A(n19916), .B(n20002), .Z(n19920) );
  XNOR U2235 ( .A(n21020), .B(n21106), .Z(n21024) );
  XNOR U2236 ( .A(n34854), .B(n34932), .Z(n34858) );
  XNOR U2237 ( .A(n34663), .B(n34744), .Z(n34667) );
  XNOR U2238 ( .A(n34451), .B(n34529), .Z(n34455) );
  XNOR U2239 ( .A(n34212), .B(n34290), .Z(n34216) );
  XNOR U2240 ( .A(n33949), .B(n34030), .Z(n33953) );
  XNOR U2241 ( .A(n33665), .B(n33743), .Z(n33669) );
  XNOR U2242 ( .A(n33354), .B(n33432), .Z(n33358) );
  XNOR U2243 ( .A(n33019), .B(n33100), .Z(n33023) );
  XNOR U2244 ( .A(n32663), .B(n32741), .Z(n32667) );
  XNOR U2245 ( .A(n32280), .B(n32358), .Z(n32284) );
  XNOR U2246 ( .A(n31697), .B(n31954), .Z(n31701) );
  XNOR U2247 ( .A(n31253), .B(n31339), .Z(n31257) );
  XNOR U2248 ( .A(n30785), .B(n30871), .Z(n30789) );
  XNOR U2249 ( .A(n30293), .B(n30379), .Z(n30297) );
  XNOR U2250 ( .A(n29777), .B(n29863), .Z(n29781) );
  XNOR U2251 ( .A(n29237), .B(n29323), .Z(n29241) );
  XNOR U2252 ( .A(n28673), .B(n28759), .Z(n28677) );
  XNOR U2253 ( .A(n28085), .B(n28171), .Z(n28089) );
  XNOR U2254 ( .A(n27473), .B(n27559), .Z(n27477) );
  XNOR U2255 ( .A(n26837), .B(n26923), .Z(n26841) );
  XNOR U2256 ( .A(n26177), .B(n26263), .Z(n26181) );
  XNOR U2257 ( .A(n25493), .B(n25579), .Z(n25497) );
  XNOR U2258 ( .A(n24785), .B(n24871), .Z(n24789) );
  XNOR U2259 ( .A(n24050), .B(n24136), .Z(n24054) );
  XNOR U2260 ( .A(n3861), .B(n3945), .Z(n3865) );
  XNOR U2261 ( .A(n4608), .B(n4689), .Z(n4609) );
  XNOR U2262 ( .A(n5351), .B(n5435), .Z(n5359) );
  XNOR U2263 ( .A(n6095), .B(n6179), .Z(n6099) );
  XNOR U2264 ( .A(n6842), .B(n6919), .Z(n6843) );
  XNOR U2265 ( .A(n9815), .B(n9901), .Z(n9823) );
  XNOR U2266 ( .A(n22503), .B(n22132), .Z(n22134) );
  XNOR U2267 ( .A(n22871), .B(n22500), .Z(n22502) );
  XNOR U2268 ( .A(n23239), .B(n22868), .Z(n22870) );
  XNOR U2269 ( .A(n23233), .B(n23313), .Z(n23237) );
  XNOR U2270 ( .A(n1996), .B(n2083), .Z(n1997) );
  XNOR U2271 ( .A(n2332), .B(n2465), .Z(n2340) );
  XNOR U2272 ( .A(n1568), .B(n1724), .Z(n1572) );
  XNOR U2273 ( .A(n807), .B(n984), .Z(n808) );
  XNOR U2274 ( .A(n1143), .B(n1365), .Z(n1151) );
  XNOR U2275 ( .A(n9076), .B(n9150), .Z(n9080) );
  XNOR U2276 ( .A(n11093), .B(n11167), .Z(n11097) );
  XNOR U2277 ( .A(n12572), .B(n12201), .Z(n12203) );
  XNOR U2278 ( .A(n13676), .B(n13305), .Z(n13307) );
  XNOR U2279 ( .A(n14780), .B(n14409), .Z(n14411) );
  XNOR U2280 ( .A(n15884), .B(n15513), .Z(n15515) );
  XNOR U2281 ( .A(n16988), .B(n16617), .Z(n16619) );
  XNOR U2282 ( .A(n18828), .B(n18457), .Z(n18459) );
  XNOR U2283 ( .A(n19932), .B(n19561), .Z(n19563) );
  XNOR U2284 ( .A(n20300), .B(n19929), .Z(n19931) );
  XNOR U2285 ( .A(n1172), .B(n1358), .Z(n1180) );
  XNOR U2286 ( .A(n2361), .B(n2458), .Z(n2369) );
  XNOR U2287 ( .A(n1597), .B(n1717), .Z(n1601) );
  XNOR U2288 ( .A(n836), .B(n977), .Z(n837) );
  XNOR U2289 ( .A(n8709), .B(n8781), .Z(n8713) );
  XNOR U2290 ( .A(n10730), .B(n10797), .Z(n10734) );
  XNOR U2291 ( .A(n11835), .B(n11903), .Z(n11839) );
  XNOR U2292 ( .A(n12939), .B(n13007), .Z(n12943) );
  XNOR U2293 ( .A(n14043), .B(n14111), .Z(n14047) );
  XNOR U2294 ( .A(n15147), .B(n15215), .Z(n15151) );
  XNOR U2295 ( .A(n16251), .B(n16319), .Z(n16255) );
  XNOR U2296 ( .A(n17355), .B(n17423), .Z(n17359) );
  XNOR U2297 ( .A(n18091), .B(n18159), .Z(n18095) );
  XNOR U2298 ( .A(n19195), .B(n19263), .Z(n19199) );
  XNOR U2299 ( .A(n20667), .B(n20735), .Z(n20671) );
  XNOR U2300 ( .A(n21403), .B(n21471), .Z(n21407) );
  XNOR U2301 ( .A(n35176), .B(n35239), .Z(n35180) );
  XNOR U2302 ( .A(n35036), .B(n35096), .Z(n35040) );
  XNOR U2303 ( .A(n34869), .B(n34929), .Z(n34873) );
  XNOR U2304 ( .A(n34678), .B(n34741), .Z(n34682) );
  XNOR U2305 ( .A(n34466), .B(n34526), .Z(n34470) );
  XNOR U2306 ( .A(n34227), .B(n34287), .Z(n34231) );
  XNOR U2307 ( .A(n33964), .B(n34027), .Z(n33968) );
  XNOR U2308 ( .A(n33680), .B(n33740), .Z(n33684) );
  XNOR U2309 ( .A(n33369), .B(n33429), .Z(n33373) );
  XNOR U2310 ( .A(n33034), .B(n33097), .Z(n33038) );
  XNOR U2311 ( .A(n32678), .B(n32738), .Z(n32682) );
  XNOR U2312 ( .A(n32295), .B(n32355), .Z(n32299) );
  XNOR U2313 ( .A(n31712), .B(n31951), .Z(n31716) );
  XNOR U2314 ( .A(n31268), .B(n31336), .Z(n31272) );
  XNOR U2315 ( .A(n30800), .B(n30868), .Z(n30804) );
  XNOR U2316 ( .A(n30308), .B(n30376), .Z(n30312) );
  XNOR U2317 ( .A(n29792), .B(n29860), .Z(n29796) );
  XNOR U2318 ( .A(n29252), .B(n29320), .Z(n29256) );
  XNOR U2319 ( .A(n28688), .B(n28756), .Z(n28692) );
  XNOR U2320 ( .A(n28100), .B(n28168), .Z(n28104) );
  XNOR U2321 ( .A(n27488), .B(n27556), .Z(n27492) );
  XNOR U2322 ( .A(n26852), .B(n26920), .Z(n26856) );
  XNOR U2323 ( .A(n26192), .B(n26260), .Z(n26196) );
  XNOR U2324 ( .A(n25508), .B(n25576), .Z(n25512) );
  XNOR U2325 ( .A(n24800), .B(n24868), .Z(n24804) );
  XNOR U2326 ( .A(n24065), .B(n24133), .Z(n24069) );
  XNOR U2327 ( .A(n3131), .B(n3197), .Z(n3135) );
  XNOR U2328 ( .A(n3880), .B(n3942), .Z(n3875) );
  XNOR U2329 ( .A(n4620), .B(n4686), .Z(n4624) );
  XNOR U2330 ( .A(n5365), .B(n5431), .Z(n5369) );
  XNOR U2331 ( .A(n6114), .B(n6176), .Z(n6109) );
  XNOR U2332 ( .A(n6854), .B(n6916), .Z(n6858) );
  XNOR U2333 ( .A(n7597), .B(n7663), .Z(n7601) );
  XNOR U2334 ( .A(n10741), .B(n10209), .Z(n10211) );
  XNOR U2335 ( .A(n22512), .B(n22574), .Z(n22516) );
  XNOR U2336 ( .A(n23248), .B(n23310), .Z(n23252) );
  XNOR U2337 ( .A(n2008), .B(n2080), .Z(n2012) );
  XNOR U2338 ( .A(n865), .B(n970), .Z(n866) );
  XNOR U2339 ( .A(n1201), .B(n1351), .Z(n1209) );
  XNOR U2340 ( .A(n1269), .B(n1335), .Z(n1273) );
  XNOR U2341 ( .A(n8349), .B(n8406), .Z(n8350) );
  XNOR U2342 ( .A(n9834), .B(n9895), .Z(n9838) );
  XNOR U2343 ( .A(n11108), .B(n11164), .Z(n11112) );
  XNOR U2344 ( .A(n12587), .B(n12216), .Z(n12218) );
  XNOR U2345 ( .A(n13691), .B(n13320), .Z(n13322) );
  XNOR U2346 ( .A(n14795), .B(n14424), .Z(n14426) );
  XNOR U2347 ( .A(n15899), .B(n15528), .Z(n15530) );
  XNOR U2348 ( .A(n17003), .B(n16632), .Z(n16634) );
  XNOR U2349 ( .A(n18107), .B(n17736), .Z(n17738) );
  XNOR U2350 ( .A(n19947), .B(n19576), .Z(n19578) );
  XNOR U2351 ( .A(n1249), .B(n1339), .Z(n1253) );
  XNOR U2352 ( .A(n1230), .B(n1344), .Z(n1238) );
  XNOR U2353 ( .A(n9464), .B(n9521), .Z(n9472) );
  XNOR U2354 ( .A(n10745), .B(n10794), .Z(n10749) );
  XNOR U2355 ( .A(n11850), .B(n11900), .Z(n11854) );
  XNOR U2356 ( .A(n12954), .B(n13004), .Z(n12958) );
  XNOR U2357 ( .A(n14058), .B(n14108), .Z(n14062) );
  XNOR U2358 ( .A(n15162), .B(n15212), .Z(n15166) );
  XNOR U2359 ( .A(n16266), .B(n16316), .Z(n16270) );
  XNOR U2360 ( .A(n17370), .B(n17420), .Z(n17374) );
  XNOR U2361 ( .A(n18474), .B(n18524), .Z(n18478) );
  XNOR U2362 ( .A(n19210), .B(n19260), .Z(n19214) );
  XNOR U2363 ( .A(n20314), .B(n20364), .Z(n20318) );
  XNOR U2364 ( .A(n21418), .B(n21468), .Z(n21422) );
  XNOR U2365 ( .A(n22154), .B(n22204), .Z(n22158) );
  XNOR U2366 ( .A(n35359), .B(n35404), .Z(n35363) );
  XNOR U2367 ( .A(n35255), .B(n35297), .Z(n35259) );
  XNOR U2368 ( .A(n35124), .B(n35166), .Z(n35128) );
  XNOR U2369 ( .A(n34969), .B(n35014), .Z(n34973) );
  XNOR U2370 ( .A(n34793), .B(n34835), .Z(n34797) );
  XNOR U2371 ( .A(n34590), .B(n34632), .Z(n34594) );
  XNOR U2372 ( .A(n34363), .B(n34408), .Z(n34367) );
  XNOR U2373 ( .A(n34115), .B(n34157), .Z(n34119) );
  XNOR U2374 ( .A(n33840), .B(n33882), .Z(n33844) );
  XNOR U2375 ( .A(n33541), .B(n33586), .Z(n33545) );
  XNOR U2376 ( .A(n33221), .B(n33263), .Z(n33225) );
  XNOR U2377 ( .A(n32874), .B(n32916), .Z(n32878) );
  XNOR U2378 ( .A(n32503), .B(n32548), .Z(n32507) );
  XNOR U2379 ( .A(n32111), .B(n32153), .Z(n32115) );
  XNOR U2380 ( .A(n31508), .B(n31558), .Z(n31512) );
  XNOR U2381 ( .A(n31052), .B(n31102), .Z(n31056) );
  XNOR U2382 ( .A(n30572), .B(n30622), .Z(n30576) );
  XNOR U2383 ( .A(n30068), .B(n30118), .Z(n30072) );
  XNOR U2384 ( .A(n29540), .B(n29590), .Z(n29544) );
  XNOR U2385 ( .A(n28988), .B(n29038), .Z(n28992) );
  XNOR U2386 ( .A(n28412), .B(n28462), .Z(n28416) );
  XNOR U2387 ( .A(n27812), .B(n27862), .Z(n27816) );
  XNOR U2388 ( .A(n27188), .B(n27238), .Z(n27192) );
  XNOR U2389 ( .A(n26540), .B(n26590), .Z(n26544) );
  XNOR U2390 ( .A(n25868), .B(n25918), .Z(n25872) );
  XNOR U2391 ( .A(n25172), .B(n25222), .Z(n25176) );
  XNOR U2392 ( .A(n24452), .B(n24502), .Z(n24456) );
  XNOR U2393 ( .A(n23631), .B(n23756), .Z(n23635) );
  XNOR U2394 ( .A(n1656), .B(n1704), .Z(n1660) );
  XNOR U2395 ( .A(n2400), .B(n2448), .Z(n2404) );
  XNOR U2396 ( .A(n3146), .B(n3194), .Z(n3150) );
  XNOR U2397 ( .A(n3890), .B(n3938), .Z(n3894) );
  XNOR U2398 ( .A(n5011), .B(n5056), .Z(n5006) );
  XNOR U2399 ( .A(n5752), .B(n5800), .Z(n5756) );
  XNOR U2400 ( .A(n6496), .B(n6544), .Z(n6500) );
  XNOR U2401 ( .A(n7241), .B(n7288), .Z(n7236) );
  XNOR U2402 ( .A(n7984), .B(n8032), .Z(n7988) );
  XNOR U2403 ( .A(n21055), .B(n21099), .Z(n21059) );
  XNOR U2404 ( .A(n22895), .B(n22939), .Z(n22899) );
  XNOR U2405 ( .A(n8733), .B(n8775), .Z(n8737) );
  XNOR U2406 ( .A(n11123), .B(n11161), .Z(n11127) );
  XNOR U2407 ( .A(n12602), .B(n12231), .Z(n12233) );
  XNOR U2408 ( .A(n13706), .B(n13335), .Z(n13337) );
  XNOR U2409 ( .A(n14810), .B(n14439), .Z(n14441) );
  XNOR U2410 ( .A(n15914), .B(n15543), .Z(n15545) );
  XNOR U2411 ( .A(n17018), .B(n16647), .Z(n16649) );
  XNOR U2412 ( .A(n18122), .B(n17751), .Z(n17753) );
  XNOR U2413 ( .A(n19226), .B(n18855), .Z(n18857) );
  XNOR U2414 ( .A(n21066), .B(n20695), .Z(n20697) );
  XNOR U2415 ( .A(n22170), .B(n21799), .Z(n21801) );
  XNOR U2416 ( .A(n11503), .B(n11131), .Z(n11133) );
  XNOR U2417 ( .A(n11865), .B(n11897), .Z(n11869) );
  XNOR U2418 ( .A(n12969), .B(n13001), .Z(n12973) );
  XNOR U2419 ( .A(n14073), .B(n14105), .Z(n14077) );
  XNOR U2420 ( .A(n15177), .B(n15209), .Z(n15181) );
  XNOR U2421 ( .A(n16281), .B(n16313), .Z(n16285) );
  XNOR U2422 ( .A(n17385), .B(n17417), .Z(n17389) );
  XNOR U2423 ( .A(n18489), .B(n18521), .Z(n18493) );
  XNOR U2424 ( .A(n19593), .B(n19625), .Z(n19597) );
  XNOR U2425 ( .A(n20329), .B(n20361), .Z(n20333) );
  XNOR U2426 ( .A(n21807), .B(n21436), .Z(n21438) );
  XNOR U2427 ( .A(n22537), .B(n22569), .Z(n22541) );
  XNOR U2428 ( .A(n35488), .B(n35515), .Z(n35492) );
  XNOR U2429 ( .A(n35420), .B(n35444), .Z(n35424) );
  XNOR U2430 ( .A(n35325), .B(n35349), .Z(n35329) );
  XNOR U2431 ( .A(n35206), .B(n35233), .Z(n35210) );
  XNOR U2432 ( .A(n35066), .B(n35090), .Z(n35070) );
  XNOR U2433 ( .A(n34899), .B(n34923), .Z(n34903) );
  XNOR U2434 ( .A(n34708), .B(n34735), .Z(n34712) );
  XNOR U2435 ( .A(n34496), .B(n34520), .Z(n34500) );
  XNOR U2436 ( .A(n34257), .B(n34281), .Z(n34261) );
  XNOR U2437 ( .A(n33994), .B(n34021), .Z(n33998) );
  XNOR U2438 ( .A(n33710), .B(n33734), .Z(n33714) );
  XNOR U2439 ( .A(n33399), .B(n33423), .Z(n33403) );
  XNOR U2440 ( .A(n33064), .B(n33091), .Z(n33068) );
  XNOR U2441 ( .A(n32708), .B(n32732), .Z(n32712) );
  XNOR U2442 ( .A(n32325), .B(n32349), .Z(n32329) );
  XNOR U2443 ( .A(n31742), .B(n31945), .Z(n31746) );
  XNOR U2444 ( .A(n31298), .B(n31330), .Z(n31302) );
  XNOR U2445 ( .A(n30830), .B(n30862), .Z(n30834) );
  XNOR U2446 ( .A(n30338), .B(n30370), .Z(n30342) );
  XNOR U2447 ( .A(n29822), .B(n29854), .Z(n29826) );
  XNOR U2448 ( .A(n29282), .B(n29314), .Z(n29286) );
  XNOR U2449 ( .A(n28718), .B(n28750), .Z(n28722) );
  XNOR U2450 ( .A(n28130), .B(n28162), .Z(n28134) );
  XNOR U2451 ( .A(n27518), .B(n27550), .Z(n27522) );
  XNOR U2452 ( .A(n26882), .B(n26914), .Z(n26886) );
  XNOR U2453 ( .A(n26222), .B(n26254), .Z(n26226) );
  XNOR U2454 ( .A(n25538), .B(n25570), .Z(n25542) );
  XNOR U2455 ( .A(n24830), .B(n24862), .Z(n24834) );
  XNOR U2456 ( .A(n24095), .B(n24127), .Z(n24099) );
  XNOR U2457 ( .A(n1299), .B(n1329), .Z(n1303) );
  XNOR U2458 ( .A(n2043), .B(n2073), .Z(n2047) );
  XNOR U2459 ( .A(n3533), .B(n3563), .Z(n3537) );
  XNOR U2460 ( .A(n4277), .B(n4307), .Z(n4281) );
  XNOR U2461 ( .A(n5769), .B(n5796), .Z(n5770) );
  XNOR U2462 ( .A(n7251), .B(n7284), .Z(n7255) );
  XNOR U2463 ( .A(n8001), .B(n8028), .Z(n8002) );
  XNOR U2464 ( .A(n10771), .B(n10238), .Z(n10240) );
  XNOR U2465 ( .A(n11139), .B(n10768), .Z(n10770) );
  XNOR U2466 ( .A(n23278), .B(n23304), .Z(n23282) );
  XNOR U2467 ( .A(n2793), .B(n2818), .Z(n2797) );
  XNOR U2468 ( .A(n5026), .B(n5051), .Z(n5030) );
  XNOR U2469 ( .A(n6888), .B(n6908), .Z(n6896) );
  XNOR U2470 ( .A(n8752), .B(n8772), .Z(n8747) );
  XNOR U2471 ( .A(n9488), .B(n9515), .Z(n9492) );
  XNOR U2472 ( .A(n12617), .B(n12246), .Z(n12248) );
  XNOR U2473 ( .A(n13721), .B(n13350), .Z(n13352) );
  XNOR U2474 ( .A(n14825), .B(n14454), .Z(n14456) );
  XNOR U2475 ( .A(n15929), .B(n15558), .Z(n15560) );
  XNOR U2476 ( .A(n17033), .B(n16662), .Z(n16664) );
  XNOR U2477 ( .A(n18137), .B(n17766), .Z(n17768) );
  XNOR U2478 ( .A(n19241), .B(n18870), .Z(n18872) );
  XNOR U2479 ( .A(n20345), .B(n19974), .Z(n19976) );
  XNOR U2480 ( .A(n22185), .B(n21814), .Z(n21816) );
  XNOR U2481 ( .A(n23289), .B(n22918), .Z(n22920) );
  XNOR U2482 ( .A(n11880), .B(n11894), .Z(n11884) );
  XNOR U2483 ( .A(n12984), .B(n12998), .Z(n12988) );
  XNOR U2484 ( .A(n14088), .B(n14102), .Z(n14092) );
  XNOR U2485 ( .A(n15192), .B(n15206), .Z(n15196) );
  XNOR U2486 ( .A(n16296), .B(n16310), .Z(n16300) );
  XNOR U2487 ( .A(n17400), .B(n17414), .Z(n17404) );
  XNOR U2488 ( .A(n18504), .B(n18518), .Z(n18508) );
  XNOR U2489 ( .A(n19608), .B(n19622), .Z(n19612) );
  XNOR U2490 ( .A(n20712), .B(n20726), .Z(n20716) );
  XNOR U2491 ( .A(n21448), .B(n21462), .Z(n21452) );
  XNOR U2492 ( .A(n22552), .B(n22566), .Z(n22556) );
  XOR U2493 ( .A(n11148), .B(n11155), .Z(n11152) );
  AND U2494 ( .A(n5786), .B(n5787), .Z(n5414) );
  AND U2495 ( .A(n7274), .B(n7275), .Z(n6902) );
  ANDN U2496 ( .B(n8762), .A(n8763), .Z(n8390) );
  NOR U2497 ( .A(n2), .B(n1), .Z(n9878) );
  AND U2498 ( .A(n11), .B(n12), .Z(n9) );
  AND U2499 ( .A(n19), .B(n20), .Z(n17) );
  AND U2500 ( .A(n27), .B(n28), .Z(n25) );
  AND U2501 ( .A(n35), .B(n36), .Z(n33) );
  AND U2502 ( .A(n43), .B(n44), .Z(n41) );
  AND U2503 ( .A(n51), .B(n52), .Z(n49) );
  AND U2504 ( .A(n59), .B(n60), .Z(n57) );
  XOR U2505 ( .A(n10352), .B(n65), .Z(n10351) );
  XNOR U2506 ( .A(n8106), .B(n8460), .Z(n8110) );
  XNOR U2507 ( .A(n8850), .B(n9200), .Z(n8854) );
  XNOR U2508 ( .A(n9593), .B(n9952), .Z(n9597) );
  XNOR U2509 ( .A(n24922), .B(n25272), .Z(n24926) );
  XNOR U2510 ( .A(n24202), .B(n24552), .Z(n24206) );
  XNOR U2511 ( .A(n23382), .B(n23806), .Z(n23386) );
  XNOR U2512 ( .A(n10874), .B(n10503), .Z(n10505) );
  XNOR U2513 ( .A(n11243), .B(n10871), .Z(n10873) );
  XNOR U2514 ( .A(n11611), .B(n11240), .Z(n11242) );
  XNOR U2515 ( .A(n11605), .B(n11949), .Z(n11609) );
  XNOR U2516 ( .A(n12346), .B(n12686), .Z(n12341) );
  XNOR U2517 ( .A(n13078), .B(n13422), .Z(n13082) );
  XNOR U2518 ( .A(n13814), .B(n14158), .Z(n13818) );
  XNOR U2519 ( .A(n14550), .B(n14894), .Z(n14554) );
  XNOR U2520 ( .A(n15286), .B(n15630), .Z(n15290) );
  XNOR U2521 ( .A(n16022), .B(n16366), .Z(n16026) );
  XNOR U2522 ( .A(n16758), .B(n17102), .Z(n16762) );
  XNOR U2523 ( .A(n17494), .B(n17838), .Z(n17498) );
  XNOR U2524 ( .A(n18230), .B(n18574), .Z(n18234) );
  XNOR U2525 ( .A(n18966), .B(n19310), .Z(n18970) );
  XNOR U2526 ( .A(n19702), .B(n20046), .Z(n19706) );
  XNOR U2527 ( .A(n20438), .B(n20782), .Z(n20442) );
  XNOR U2528 ( .A(n21174), .B(n21518), .Z(n21178) );
  XNOR U2529 ( .A(n21910), .B(n22254), .Z(n21914) );
  XNOR U2530 ( .A(n22646), .B(n22990), .Z(n22650) );
  XNOR U2531 ( .A(n7356), .B(n7717), .Z(n7361) );
  XNOR U2532 ( .A(n8865), .B(n9197), .Z(n8869) );
  XNOR U2533 ( .A(n9608), .B(n9949), .Z(n9612) );
  XNOR U2534 ( .A(n25633), .B(n25965), .Z(n25637) );
  XNOR U2535 ( .A(n24937), .B(n25269), .Z(n24941) );
  XNOR U2536 ( .A(n24217), .B(n24549), .Z(n24221) );
  XNOR U2537 ( .A(n23397), .B(n23803), .Z(n23401) );
  XNOR U2538 ( .A(n7749), .B(n8085), .Z(n7753) );
  XNOR U2539 ( .A(n10889), .B(n10518), .Z(n10520) );
  XNOR U2540 ( .A(n11258), .B(n10886), .Z(n10888) );
  XNOR U2541 ( .A(n11626), .B(n11255), .Z(n11257) );
  XNOR U2542 ( .A(n11620), .B(n11946), .Z(n11624) );
  XNOR U2543 ( .A(n11988), .B(n12314), .Z(n11992) );
  XNOR U2544 ( .A(n12356), .B(n12682), .Z(n12360) );
  XNOR U2545 ( .A(n12724), .B(n13050), .Z(n12728) );
  XNOR U2546 ( .A(n13087), .B(n13418), .Z(n13096) );
  XNOR U2547 ( .A(n13829), .B(n14155), .Z(n13837) );
  XNOR U2548 ( .A(n14565), .B(n14891), .Z(n14569) );
  XNOR U2549 ( .A(n15301), .B(n15627), .Z(n15305) );
  XNOR U2550 ( .A(n16037), .B(n16363), .Z(n16041) );
  XNOR U2551 ( .A(n16773), .B(n17099), .Z(n16777) );
  XNOR U2552 ( .A(n17509), .B(n17835), .Z(n17513) );
  XNOR U2553 ( .A(n18245), .B(n18571), .Z(n18249) );
  XNOR U2554 ( .A(n18981), .B(n19307), .Z(n18985) );
  XNOR U2555 ( .A(n19717), .B(n20043), .Z(n19721) );
  XNOR U2556 ( .A(n20453), .B(n20779), .Z(n20457) );
  XNOR U2557 ( .A(n21189), .B(n21515), .Z(n21193) );
  XNOR U2558 ( .A(n21925), .B(n22251), .Z(n21929) );
  XNOR U2559 ( .A(n22661), .B(n22987), .Z(n22665) );
  XNOR U2560 ( .A(n6987), .B(n7344), .Z(n6991) );
  XNOR U2561 ( .A(n8880), .B(n9194), .Z(n8884) );
  XNOR U2562 ( .A(n9623), .B(n9946), .Z(n9627) );
  XNOR U2563 ( .A(n26968), .B(n27282), .Z(n26972) );
  XNOR U2564 ( .A(n26320), .B(n26634), .Z(n26324) );
  XNOR U2565 ( .A(n25648), .B(n25962), .Z(n25652) );
  XNOR U2566 ( .A(n24952), .B(n25266), .Z(n24956) );
  XNOR U2567 ( .A(n24232), .B(n24546), .Z(n24236) );
  XNOR U2568 ( .A(n23412), .B(n23800), .Z(n23416) );
  XNOR U2569 ( .A(n7764), .B(n8082), .Z(n7768) );
  XNOR U2570 ( .A(n8513), .B(n8825), .Z(n8517) );
  XNOR U2571 ( .A(n10904), .B(n10533), .Z(n10535) );
  XNOR U2572 ( .A(n11273), .B(n10901), .Z(n10903) );
  XNOR U2573 ( .A(n11641), .B(n11270), .Z(n11272) );
  XNOR U2574 ( .A(n11635), .B(n11943), .Z(n11639) );
  XNOR U2575 ( .A(n12003), .B(n12311), .Z(n12007) );
  XNOR U2576 ( .A(n12371), .B(n12679), .Z(n12375) );
  XNOR U2577 ( .A(n12739), .B(n13047), .Z(n12743) );
  XNOR U2578 ( .A(n13107), .B(n13415), .Z(n13111) );
  XNOR U2579 ( .A(n13475), .B(n13783), .Z(n13479) );
  XNOR U2580 ( .A(n13843), .B(n14151), .Z(n13847) );
  XNOR U2581 ( .A(n14584), .B(n14888), .Z(n14579) );
  XNOR U2582 ( .A(n15316), .B(n15624), .Z(n15320) );
  XNOR U2583 ( .A(n16052), .B(n16360), .Z(n16056) );
  XNOR U2584 ( .A(n16788), .B(n17096), .Z(n16792) );
  XNOR U2585 ( .A(n17524), .B(n17832), .Z(n17528) );
  XNOR U2586 ( .A(n18260), .B(n18568), .Z(n18264) );
  XNOR U2587 ( .A(n18996), .B(n19304), .Z(n19000) );
  XNOR U2588 ( .A(n19732), .B(n20040), .Z(n19736) );
  XNOR U2589 ( .A(n20468), .B(n20776), .Z(n20472) );
  XNOR U2590 ( .A(n21204), .B(n21512), .Z(n21208) );
  XNOR U2591 ( .A(n21940), .B(n22248), .Z(n21944) );
  XNOR U2592 ( .A(n22676), .B(n22984), .Z(n22680) );
  XNOR U2593 ( .A(n6241), .B(n6602), .Z(n6246) );
  XNOR U2594 ( .A(n6629), .B(n6967), .Z(n6633) );
  XNOR U2595 ( .A(n9638), .B(n9943), .Z(n9642) );
  XNOR U2596 ( .A(n27607), .B(n27903), .Z(n27611) );
  XNOR U2597 ( .A(n26983), .B(n27279), .Z(n26987) );
  XNOR U2598 ( .A(n26335), .B(n26631), .Z(n26339) );
  XNOR U2599 ( .A(n25663), .B(n25959), .Z(n25667) );
  XNOR U2600 ( .A(n24967), .B(n25263), .Z(n24971) );
  XNOR U2601 ( .A(n24247), .B(n24543), .Z(n24251) );
  XNOR U2602 ( .A(n23427), .B(n23797), .Z(n23431) );
  XNOR U2603 ( .A(n7012), .B(n7339), .Z(n7016) );
  XNOR U2604 ( .A(n8156), .B(n8450), .Z(n8160) );
  XNOR U2605 ( .A(n8900), .B(n9190), .Z(n8904) );
  XNOR U2606 ( .A(n10919), .B(n10548), .Z(n10550) );
  XNOR U2607 ( .A(n11288), .B(n10916), .Z(n10918) );
  XNOR U2608 ( .A(n11656), .B(n11285), .Z(n11287) );
  XNOR U2609 ( .A(n11650), .B(n11940), .Z(n11654) );
  XNOR U2610 ( .A(n12018), .B(n12308), .Z(n12022) );
  XNOR U2611 ( .A(n12386), .B(n12676), .Z(n12390) );
  XNOR U2612 ( .A(n12754), .B(n13044), .Z(n12758) );
  XNOR U2613 ( .A(n13122), .B(n13412), .Z(n13126) );
  XNOR U2614 ( .A(n13490), .B(n13780), .Z(n13494) );
  XNOR U2615 ( .A(n13858), .B(n14148), .Z(n13862) );
  XNOR U2616 ( .A(n14226), .B(n14516), .Z(n14230) );
  XNOR U2617 ( .A(n14594), .B(n14884), .Z(n14598) );
  XNOR U2618 ( .A(n14962), .B(n15252), .Z(n14966) );
  XNOR U2619 ( .A(n15325), .B(n15620), .Z(n15334) );
  XNOR U2620 ( .A(n16067), .B(n16357), .Z(n16075) );
  XNOR U2621 ( .A(n16803), .B(n17093), .Z(n16807) );
  XNOR U2622 ( .A(n17539), .B(n17829), .Z(n17543) );
  XNOR U2623 ( .A(n18275), .B(n18565), .Z(n18279) );
  XNOR U2624 ( .A(n19011), .B(n19301), .Z(n19015) );
  XNOR U2625 ( .A(n19747), .B(n20037), .Z(n19751) );
  XNOR U2626 ( .A(n20483), .B(n20773), .Z(n20487) );
  XNOR U2627 ( .A(n21219), .B(n21509), .Z(n21223) );
  XNOR U2628 ( .A(n21955), .B(n22245), .Z(n21959) );
  XNOR U2629 ( .A(n22691), .B(n22981), .Z(n22695) );
  XNOR U2630 ( .A(n5880), .B(n6228), .Z(n5884) );
  XNOR U2631 ( .A(n10030), .B(n10450), .Z(n10034) );
  XNOR U2632 ( .A(n28798), .B(n29076), .Z(n28802) );
  XNOR U2633 ( .A(n28222), .B(n28500), .Z(n28226) );
  XNOR U2634 ( .A(n27622), .B(n27900), .Z(n27626) );
  XNOR U2635 ( .A(n26998), .B(n27276), .Z(n27002) );
  XNOR U2636 ( .A(n26350), .B(n26628), .Z(n26354) );
  XNOR U2637 ( .A(n25678), .B(n25956), .Z(n25682) );
  XNOR U2638 ( .A(n24982), .B(n25260), .Z(n24986) );
  XNOR U2639 ( .A(n24262), .B(n24540), .Z(n24266) );
  XNOR U2640 ( .A(n23442), .B(n23794), .Z(n23446) );
  XNOR U2641 ( .A(n7412), .B(n7706), .Z(n7416) );
  XNOR U2642 ( .A(n6267), .B(n6597), .Z(n6271) );
  XNOR U2643 ( .A(n8915), .B(n9187), .Z(n8919) );
  XNOR U2644 ( .A(n9658), .B(n9939), .Z(n9662) );
  XNOR U2645 ( .A(n11303), .B(n10931), .Z(n10933) );
  XNOR U2646 ( .A(n11671), .B(n11300), .Z(n11302) );
  XNOR U2647 ( .A(n11665), .B(n11937), .Z(n11669) );
  XNOR U2648 ( .A(n12033), .B(n12305), .Z(n12037) );
  XNOR U2649 ( .A(n12401), .B(n12673), .Z(n12405) );
  XNOR U2650 ( .A(n12769), .B(n13041), .Z(n12773) );
  XNOR U2651 ( .A(n13137), .B(n13409), .Z(n13141) );
  XNOR U2652 ( .A(n13505), .B(n13777), .Z(n13509) );
  XNOR U2653 ( .A(n13873), .B(n14145), .Z(n13877) );
  XNOR U2654 ( .A(n14241), .B(n14513), .Z(n14245) );
  XNOR U2655 ( .A(n14609), .B(n14881), .Z(n14613) );
  XNOR U2656 ( .A(n14977), .B(n15249), .Z(n14981) );
  XNOR U2657 ( .A(n15345), .B(n15617), .Z(n15349) );
  XNOR U2658 ( .A(n15713), .B(n15985), .Z(n15717) );
  XNOR U2659 ( .A(n16081), .B(n16353), .Z(n16085) );
  XNOR U2660 ( .A(n16822), .B(n17090), .Z(n16817) );
  XNOR U2661 ( .A(n17554), .B(n17826), .Z(n17558) );
  XNOR U2662 ( .A(n18290), .B(n18562), .Z(n18294) );
  XNOR U2663 ( .A(n19026), .B(n19298), .Z(n19030) );
  XNOR U2664 ( .A(n19762), .B(n20034), .Z(n19766) );
  XNOR U2665 ( .A(n20498), .B(n20770), .Z(n20502) );
  XNOR U2666 ( .A(n21234), .B(n21506), .Z(n21238) );
  XNOR U2667 ( .A(n21970), .B(n22242), .Z(n21974) );
  XNOR U2668 ( .A(n22706), .B(n22978), .Z(n22710) );
  XNOR U2669 ( .A(n6654), .B(n6962), .Z(n6658) );
  XNOR U2670 ( .A(n8548), .B(n8818), .Z(n8552) );
  XNOR U2671 ( .A(n29365), .B(n29625), .Z(n29369) );
  XNOR U2672 ( .A(n28813), .B(n29073), .Z(n28817) );
  XNOR U2673 ( .A(n28237), .B(n28497), .Z(n28241) );
  XNOR U2674 ( .A(n27637), .B(n27897), .Z(n27641) );
  XNOR U2675 ( .A(n27013), .B(n27273), .Z(n27017) );
  XNOR U2676 ( .A(n26365), .B(n26625), .Z(n26369) );
  XNOR U2677 ( .A(n25693), .B(n25953), .Z(n25697) );
  XNOR U2678 ( .A(n24997), .B(n25257), .Z(n25001) );
  XNOR U2679 ( .A(n24277), .B(n24537), .Z(n24281) );
  XNOR U2680 ( .A(n23457), .B(n23791), .Z(n23461) );
  XNOR U2681 ( .A(n7427), .B(n7703), .Z(n7431) );
  XNOR U2682 ( .A(n5518), .B(n5854), .Z(n5522) );
  XNOR U2683 ( .A(n9673), .B(n9936), .Z(n9677) );
  XNOR U2684 ( .A(n10949), .B(n10578), .Z(n10580) );
  XNOR U2685 ( .A(n11686), .B(n11315), .Z(n11317) );
  XNOR U2686 ( .A(n11680), .B(n11934), .Z(n11684) );
  XNOR U2687 ( .A(n12048), .B(n12302), .Z(n12052) );
  XNOR U2688 ( .A(n12416), .B(n12670), .Z(n12420) );
  XNOR U2689 ( .A(n12784), .B(n13038), .Z(n12788) );
  XNOR U2690 ( .A(n13152), .B(n13406), .Z(n13156) );
  XNOR U2691 ( .A(n13520), .B(n13774), .Z(n13524) );
  XNOR U2692 ( .A(n13888), .B(n14142), .Z(n13892) );
  XNOR U2693 ( .A(n14256), .B(n14510), .Z(n14260) );
  XNOR U2694 ( .A(n14624), .B(n14878), .Z(n14628) );
  XNOR U2695 ( .A(n14992), .B(n15246), .Z(n14996) );
  XNOR U2696 ( .A(n15360), .B(n15614), .Z(n15364) );
  XNOR U2697 ( .A(n15728), .B(n15982), .Z(n15732) );
  XNOR U2698 ( .A(n16096), .B(n16350), .Z(n16100) );
  XNOR U2699 ( .A(n16464), .B(n16718), .Z(n16468) );
  XNOR U2700 ( .A(n16832), .B(n17086), .Z(n16836) );
  XNOR U2701 ( .A(n17200), .B(n17454), .Z(n17204) );
  XNOR U2702 ( .A(n17563), .B(n17822), .Z(n17572) );
  XNOR U2703 ( .A(n18305), .B(n18559), .Z(n18313) );
  XNOR U2704 ( .A(n19041), .B(n19295), .Z(n19045) );
  XNOR U2705 ( .A(n19777), .B(n20031), .Z(n19781) );
  XNOR U2706 ( .A(n20513), .B(n20767), .Z(n20517) );
  XNOR U2707 ( .A(n21249), .B(n21503), .Z(n21253) );
  XNOR U2708 ( .A(n21985), .B(n22239), .Z(n21989) );
  XNOR U2709 ( .A(n22721), .B(n22975), .Z(n22725) );
  XNOR U2710 ( .A(n4758), .B(n5113), .Z(n4762) );
  XNOR U2711 ( .A(n8563), .B(n8815), .Z(n8567) );
  XNOR U2712 ( .A(n9303), .B(n9558), .Z(n9307) );
  XNOR U2713 ( .A(n11691), .B(n11320), .Z(n11322) );
  XNOR U2714 ( .A(n6292), .B(n6592), .Z(n6296) );
  XNOR U2715 ( .A(n30412), .B(n30654), .Z(n30416) );
  XNOR U2716 ( .A(n29908), .B(n30150), .Z(n29912) );
  XNOR U2717 ( .A(n29380), .B(n29622), .Z(n29384) );
  XNOR U2718 ( .A(n28828), .B(n29070), .Z(n28832) );
  XNOR U2719 ( .A(n28252), .B(n28494), .Z(n28256) );
  XNOR U2720 ( .A(n27652), .B(n27894), .Z(n27656) );
  XNOR U2721 ( .A(n27028), .B(n27270), .Z(n27032) );
  XNOR U2722 ( .A(n26380), .B(n26622), .Z(n26384) );
  XNOR U2723 ( .A(n25708), .B(n25950), .Z(n25712) );
  XNOR U2724 ( .A(n25012), .B(n25254), .Z(n25016) );
  XNOR U2725 ( .A(n24292), .B(n24534), .Z(n24296) );
  XNOR U2726 ( .A(n23472), .B(n23788), .Z(n23476) );
  XNOR U2727 ( .A(n7442), .B(n7700), .Z(n7446) );
  XNOR U2728 ( .A(n6679), .B(n6957), .Z(n6683) );
  XNOR U2729 ( .A(n5151), .B(n5481), .Z(n5155) );
  XNOR U2730 ( .A(n10964), .B(n10593), .Z(n10595) );
  XNOR U2731 ( .A(n11701), .B(n11330), .Z(n11332) );
  XNOR U2732 ( .A(n12431), .B(n12667), .Z(n12435) );
  XNOR U2733 ( .A(n12799), .B(n13035), .Z(n12803) );
  XNOR U2734 ( .A(n13167), .B(n13403), .Z(n13171) );
  XNOR U2735 ( .A(n13535), .B(n13771), .Z(n13539) );
  XNOR U2736 ( .A(n13903), .B(n14139), .Z(n13907) );
  XNOR U2737 ( .A(n14271), .B(n14507), .Z(n14275) );
  XNOR U2738 ( .A(n14639), .B(n14875), .Z(n14643) );
  XNOR U2739 ( .A(n15007), .B(n15243), .Z(n15011) );
  XNOR U2740 ( .A(n15375), .B(n15611), .Z(n15379) );
  XNOR U2741 ( .A(n15743), .B(n15979), .Z(n15747) );
  XNOR U2742 ( .A(n16111), .B(n16347), .Z(n16115) );
  XNOR U2743 ( .A(n16479), .B(n16715), .Z(n16483) );
  XNOR U2744 ( .A(n16847), .B(n17083), .Z(n16851) );
  XNOR U2745 ( .A(n17215), .B(n17451), .Z(n17219) );
  XNOR U2746 ( .A(n17583), .B(n17819), .Z(n17587) );
  XNOR U2747 ( .A(n17951), .B(n18187), .Z(n17955) );
  XNOR U2748 ( .A(n18319), .B(n18555), .Z(n18323) );
  XNOR U2749 ( .A(n19060), .B(n19292), .Z(n19055) );
  XNOR U2750 ( .A(n19792), .B(n20028), .Z(n19796) );
  XNOR U2751 ( .A(n20528), .B(n20764), .Z(n20532) );
  XNOR U2752 ( .A(n21264), .B(n21500), .Z(n21268) );
  XNOR U2753 ( .A(n22000), .B(n22236), .Z(n22004) );
  XNOR U2754 ( .A(n22736), .B(n22972), .Z(n22740) );
  XNOR U2755 ( .A(n4391), .B(n4739), .Z(n4395) );
  XNOR U2756 ( .A(n8206), .B(n8440), .Z(n8210) );
  XNOR U2757 ( .A(n8950), .B(n9180), .Z(n8954) );
  XNOR U2758 ( .A(n9693), .B(n9932), .Z(n9697) );
  XNOR U2759 ( .A(n11706), .B(n11335), .Z(n11337) );
  XNOR U2760 ( .A(n12068), .B(n12298), .Z(n12072) );
  XNOR U2761 ( .A(n5543), .B(n5849), .Z(n5547) );
  XNOR U2762 ( .A(n11343), .B(n10971), .Z(n10973) );
  XNOR U2763 ( .A(n30907), .B(n31131), .Z(n30911) );
  XNOR U2764 ( .A(n30427), .B(n30651), .Z(n30431) );
  XNOR U2765 ( .A(n29923), .B(n30147), .Z(n29927) );
  XNOR U2766 ( .A(n29395), .B(n29619), .Z(n29399) );
  XNOR U2767 ( .A(n28843), .B(n29067), .Z(n28847) );
  XNOR U2768 ( .A(n28267), .B(n28491), .Z(n28271) );
  XNOR U2769 ( .A(n27667), .B(n27891), .Z(n27671) );
  XNOR U2770 ( .A(n27043), .B(n27267), .Z(n27047) );
  XNOR U2771 ( .A(n26395), .B(n26619), .Z(n26399) );
  XNOR U2772 ( .A(n25723), .B(n25947), .Z(n25727) );
  XNOR U2773 ( .A(n25027), .B(n25251), .Z(n25031) );
  XNOR U2774 ( .A(n24307), .B(n24531), .Z(n24311) );
  XNOR U2775 ( .A(n23487), .B(n23785), .Z(n23491) );
  XNOR U2776 ( .A(n6694), .B(n6954), .Z(n6698) );
  XNOR U2777 ( .A(n5930), .B(n6218), .Z(n5934) );
  XNOR U2778 ( .A(n4783), .B(n5108), .Z(n4787) );
  XNOR U2779 ( .A(n11710), .B(n11928), .Z(n11714) );
  XNOR U2780 ( .A(n13550), .B(n13768), .Z(n13554) );
  XNOR U2781 ( .A(n13918), .B(n14136), .Z(n13922) );
  XNOR U2782 ( .A(n14286), .B(n14504), .Z(n14290) );
  XNOR U2783 ( .A(n14654), .B(n14872), .Z(n14658) );
  XNOR U2784 ( .A(n15022), .B(n15240), .Z(n15026) );
  XNOR U2785 ( .A(n15390), .B(n15608), .Z(n15394) );
  XNOR U2786 ( .A(n15758), .B(n15976), .Z(n15762) );
  XNOR U2787 ( .A(n16126), .B(n16344), .Z(n16130) );
  XNOR U2788 ( .A(n16494), .B(n16712), .Z(n16498) );
  XNOR U2789 ( .A(n16862), .B(n17080), .Z(n16866) );
  XNOR U2790 ( .A(n17230), .B(n17448), .Z(n17234) );
  XNOR U2791 ( .A(n17598), .B(n17816), .Z(n17602) );
  XNOR U2792 ( .A(n17966), .B(n18184), .Z(n17970) );
  XNOR U2793 ( .A(n18334), .B(n18552), .Z(n18338) );
  XNOR U2794 ( .A(n18702), .B(n18920), .Z(n18706) );
  XNOR U2795 ( .A(n19070), .B(n19288), .Z(n19074) );
  XNOR U2796 ( .A(n19438), .B(n19656), .Z(n19442) );
  XNOR U2797 ( .A(n19801), .B(n20024), .Z(n19810) );
  XNOR U2798 ( .A(n20543), .B(n20761), .Z(n20551) );
  XNOR U2799 ( .A(n21279), .B(n21497), .Z(n21283) );
  XNOR U2800 ( .A(n22015), .B(n22233), .Z(n22019) );
  XNOR U2801 ( .A(n22751), .B(n22969), .Z(n22755) );
  XNOR U2802 ( .A(n7077), .B(n7326), .Z(n7081) );
  XNOR U2803 ( .A(n4024), .B(n4366), .Z(n4028) );
  XNOR U2804 ( .A(n8965), .B(n9177), .Z(n8969) );
  XNOR U2805 ( .A(n9708), .B(n9929), .Z(n9712) );
  XNOR U2806 ( .A(n10984), .B(n10613), .Z(n10615) );
  XNOR U2807 ( .A(n11347), .B(n11559), .Z(n11351) );
  XNOR U2808 ( .A(n12451), .B(n12663), .Z(n12455) );
  XNOR U2809 ( .A(n13187), .B(n13399), .Z(n13191) );
  XNOR U2810 ( .A(n7853), .B(n8065), .Z(n7848) );
  XNOR U2811 ( .A(n11726), .B(n11355), .Z(n11357) );
  XNOR U2812 ( .A(n12462), .B(n12091), .Z(n12093) );
  XNOR U2813 ( .A(n31981), .B(n32179), .Z(n31985) );
  XNOR U2814 ( .A(n31378), .B(n31584), .Z(n31382) );
  XNOR U2815 ( .A(n30922), .B(n31128), .Z(n30926) );
  XNOR U2816 ( .A(n30442), .B(n30648), .Z(n30446) );
  XNOR U2817 ( .A(n29938), .B(n30144), .Z(n29942) );
  XNOR U2818 ( .A(n29410), .B(n29616), .Z(n29414) );
  XNOR U2819 ( .A(n28858), .B(n29064), .Z(n28862) );
  XNOR U2820 ( .A(n28282), .B(n28488), .Z(n28286) );
  XNOR U2821 ( .A(n27682), .B(n27888), .Z(n27686) );
  XNOR U2822 ( .A(n27058), .B(n27264), .Z(n27062) );
  XNOR U2823 ( .A(n26410), .B(n26616), .Z(n26414) );
  XNOR U2824 ( .A(n25738), .B(n25944), .Z(n25742) );
  XNOR U2825 ( .A(n25042), .B(n25248), .Z(n25046) );
  XNOR U2826 ( .A(n24322), .B(n24528), .Z(n24326) );
  XNOR U2827 ( .A(n23502), .B(n23782), .Z(n23506) );
  XNOR U2828 ( .A(n6728), .B(n6946), .Z(n6732) );
  XNOR U2829 ( .A(n5945), .B(n6215), .Z(n5949) );
  XNOR U2830 ( .A(n5181), .B(n5475), .Z(n5185) );
  XNOR U2831 ( .A(n12829), .B(n13029), .Z(n12833) );
  XNOR U2832 ( .A(n14669), .B(n14869), .Z(n14673) );
  XNOR U2833 ( .A(n15037), .B(n15237), .Z(n15041) );
  XNOR U2834 ( .A(n15405), .B(n15605), .Z(n15409) );
  XNOR U2835 ( .A(n15773), .B(n15973), .Z(n15777) );
  XNOR U2836 ( .A(n16141), .B(n16341), .Z(n16145) );
  XNOR U2837 ( .A(n16509), .B(n16709), .Z(n16513) );
  XNOR U2838 ( .A(n16877), .B(n17077), .Z(n16881) );
  XNOR U2839 ( .A(n17245), .B(n17445), .Z(n17249) );
  XNOR U2840 ( .A(n17613), .B(n17813), .Z(n17617) );
  XNOR U2841 ( .A(n17981), .B(n18181), .Z(n17985) );
  XNOR U2842 ( .A(n18349), .B(n18549), .Z(n18353) );
  XNOR U2843 ( .A(n18717), .B(n18917), .Z(n18721) );
  XNOR U2844 ( .A(n19085), .B(n19285), .Z(n19089) );
  XNOR U2845 ( .A(n19453), .B(n19653), .Z(n19457) );
  XNOR U2846 ( .A(n19821), .B(n20021), .Z(n19825) );
  XNOR U2847 ( .A(n20189), .B(n20389), .Z(n20193) );
  XNOR U2848 ( .A(n20557), .B(n20757), .Z(n20561) );
  XNOR U2849 ( .A(n21298), .B(n21494), .Z(n21293) );
  XNOR U2850 ( .A(n22030), .B(n22230), .Z(n22034) );
  XNOR U2851 ( .A(n22766), .B(n22966), .Z(n22770) );
  XNOR U2852 ( .A(n6714), .B(n6950), .Z(n6722) );
  XNOR U2853 ( .A(n4421), .B(n4733), .Z(n4425) );
  XNOR U2854 ( .A(n3657), .B(n3993), .Z(n3661) );
  XNOR U2855 ( .A(n7863), .B(n8061), .Z(n7867) );
  XNOR U2856 ( .A(n8610), .B(n8805), .Z(n8611) );
  XNOR U2857 ( .A(n9348), .B(n9549), .Z(n9356) );
  XNOR U2858 ( .A(n10100), .B(n10422), .Z(n10104) );
  XNOR U2859 ( .A(n10625), .B(n10818), .Z(n10629) );
  XNOR U2860 ( .A(n11736), .B(n11365), .Z(n11367) );
  XNOR U2861 ( .A(n11730), .B(n11924), .Z(n11734) );
  XNOR U2862 ( .A(n13570), .B(n13764), .Z(n13574) );
  XNOR U2863 ( .A(n14306), .B(n14500), .Z(n14310) );
  XNOR U2864 ( .A(n7116), .B(n7317), .Z(n7124) );
  XNOR U2865 ( .A(n2898), .B(n3252), .Z(n2902) );
  XNOR U2866 ( .A(n11741), .B(n11370), .Z(n11372) );
  XNOR U2867 ( .A(n12471), .B(n12659), .Z(n12475) );
  XNOR U2868 ( .A(n13581), .B(n13210), .Z(n13212) );
  XNOR U2869 ( .A(n32388), .B(n32571), .Z(n32392) );
  XNOR U2870 ( .A(n31996), .B(n32176), .Z(n32000) );
  XNOR U2871 ( .A(n31393), .B(n31581), .Z(n31397) );
  XNOR U2872 ( .A(n30937), .B(n31125), .Z(n30941) );
  XNOR U2873 ( .A(n30457), .B(n30645), .Z(n30461) );
  XNOR U2874 ( .A(n29953), .B(n30141), .Z(n29957) );
  XNOR U2875 ( .A(n29425), .B(n29613), .Z(n29429) );
  XNOR U2876 ( .A(n28873), .B(n29061), .Z(n28877) );
  XNOR U2877 ( .A(n28297), .B(n28485), .Z(n28301) );
  XNOR U2878 ( .A(n27697), .B(n27885), .Z(n27701) );
  XNOR U2879 ( .A(n27073), .B(n27261), .Z(n27077) );
  XNOR U2880 ( .A(n26425), .B(n26613), .Z(n26429) );
  XNOR U2881 ( .A(n25753), .B(n25941), .Z(n25757) );
  XNOR U2882 ( .A(n25057), .B(n25245), .Z(n25061) );
  XNOR U2883 ( .A(n24337), .B(n24525), .Z(n24341) );
  XNOR U2884 ( .A(n23517), .B(n23779), .Z(n23521) );
  XNOR U2885 ( .A(n6361), .B(n6577), .Z(n6365) );
  XNOR U2886 ( .A(n5218), .B(n5467), .Z(n5219) );
  XNOR U2887 ( .A(n5578), .B(n5842), .Z(n5582) );
  XNOR U2888 ( .A(n4813), .B(n5102), .Z(n4817) );
  XNOR U2889 ( .A(n13948), .B(n14130), .Z(n13952) );
  XNOR U2890 ( .A(n15788), .B(n15970), .Z(n15792) );
  XNOR U2891 ( .A(n16156), .B(n16338), .Z(n16160) );
  XNOR U2892 ( .A(n16524), .B(n16706), .Z(n16528) );
  XNOR U2893 ( .A(n16892), .B(n17074), .Z(n16896) );
  XNOR U2894 ( .A(n17260), .B(n17442), .Z(n17264) );
  XNOR U2895 ( .A(n17628), .B(n17810), .Z(n17632) );
  XNOR U2896 ( .A(n17996), .B(n18178), .Z(n18000) );
  XNOR U2897 ( .A(n18364), .B(n18546), .Z(n18368) );
  XNOR U2898 ( .A(n18732), .B(n18914), .Z(n18736) );
  XNOR U2899 ( .A(n19100), .B(n19282), .Z(n19104) );
  XNOR U2900 ( .A(n19468), .B(n19650), .Z(n19472) );
  XNOR U2901 ( .A(n19836), .B(n20018), .Z(n19840) );
  XNOR U2902 ( .A(n20204), .B(n20386), .Z(n20208) );
  XNOR U2903 ( .A(n20572), .B(n20754), .Z(n20576) );
  XNOR U2904 ( .A(n20940), .B(n21122), .Z(n20944) );
  XNOR U2905 ( .A(n21308), .B(n21490), .Z(n21312) );
  XNOR U2906 ( .A(n21676), .B(n21858), .Z(n21680) );
  XNOR U2907 ( .A(n22039), .B(n22226), .Z(n22048) );
  XNOR U2908 ( .A(n22781), .B(n22963), .Z(n22789) );
  XNOR U2909 ( .A(n5602), .B(n5836), .Z(n5606) );
  XNOR U2910 ( .A(n5969), .B(n6211), .Z(n5964) );
  XNOR U2911 ( .A(n4054), .B(n4360), .Z(n4058) );
  XNOR U2912 ( .A(n3290), .B(n3620), .Z(n3294) );
  XNOR U2913 ( .A(n5247), .B(n5460), .Z(n5248) );
  XNOR U2914 ( .A(n7130), .B(n7313), .Z(n7134) );
  XNOR U2915 ( .A(n7882), .B(n8058), .Z(n7877) );
  XNOR U2916 ( .A(n8622), .B(n8802), .Z(n8626) );
  XNOR U2917 ( .A(n9362), .B(n9545), .Z(n9366) );
  XNOR U2918 ( .A(n10119), .B(n10416), .Z(n10113) );
  XNOR U2919 ( .A(n11383), .B(n11011), .Z(n11013) );
  XNOR U2920 ( .A(n11751), .B(n11380), .Z(n11382) );
  XNOR U2921 ( .A(n11745), .B(n11921), .Z(n11749) );
  XNOR U2922 ( .A(n12849), .B(n13025), .Z(n12853) );
  XNOR U2923 ( .A(n14689), .B(n14865), .Z(n14693) );
  XNOR U2924 ( .A(n15425), .B(n15601), .Z(n15429) );
  XNOR U2925 ( .A(n2530), .B(n2879), .Z(n2534) );
  XNOR U2926 ( .A(n6013), .B(n6199), .Z(n6017) );
  XNOR U2927 ( .A(n12486), .B(n12656), .Z(n12490) );
  XNOR U2928 ( .A(n13590), .B(n13760), .Z(n13594) );
  XNOR U2929 ( .A(n14700), .B(n14329), .Z(n14331) );
  XNOR U2930 ( .A(n33121), .B(n33283), .Z(n33125) );
  XNOR U2931 ( .A(n32774), .B(n32936), .Z(n32778) );
  XNOR U2932 ( .A(n32403), .B(n32568), .Z(n32407) );
  XNOR U2933 ( .A(n32011), .B(n32173), .Z(n32015) );
  XNOR U2934 ( .A(n31408), .B(n31578), .Z(n31412) );
  XNOR U2935 ( .A(n30952), .B(n31122), .Z(n30956) );
  XNOR U2936 ( .A(n30472), .B(n30642), .Z(n30476) );
  XNOR U2937 ( .A(n29968), .B(n30138), .Z(n29972) );
  XNOR U2938 ( .A(n29440), .B(n29610), .Z(n29444) );
  XNOR U2939 ( .A(n28888), .B(n29058), .Z(n28892) );
  XNOR U2940 ( .A(n28312), .B(n28482), .Z(n28316) );
  XNOR U2941 ( .A(n27712), .B(n27882), .Z(n27716) );
  XNOR U2942 ( .A(n27088), .B(n27258), .Z(n27092) );
  XNOR U2943 ( .A(n26440), .B(n26610), .Z(n26444) );
  XNOR U2944 ( .A(n25768), .B(n25938), .Z(n25772) );
  XNOR U2945 ( .A(n25072), .B(n25242), .Z(n25076) );
  XNOR U2946 ( .A(n24352), .B(n24522), .Z(n24356) );
  XNOR U2947 ( .A(n23536), .B(n23776), .Z(n23530) );
  XNOR U2948 ( .A(n5998), .B(n6204), .Z(n5993) );
  XNOR U2949 ( .A(n4828), .B(n5099), .Z(n4836) );
  XNOR U2950 ( .A(n5655), .B(n5823), .Z(n5659) );
  XNOR U2951 ( .A(n11761), .B(n11390), .Z(n11392) );
  XNOR U2952 ( .A(n15067), .B(n15231), .Z(n15071) );
  XNOR U2953 ( .A(n16907), .B(n17071), .Z(n16911) );
  XNOR U2954 ( .A(n17275), .B(n17439), .Z(n17279) );
  XNOR U2955 ( .A(n17643), .B(n17807), .Z(n17647) );
  XNOR U2956 ( .A(n18011), .B(n18175), .Z(n18015) );
  XNOR U2957 ( .A(n18379), .B(n18543), .Z(n18383) );
  XNOR U2958 ( .A(n18747), .B(n18911), .Z(n18751) );
  XNOR U2959 ( .A(n19115), .B(n19279), .Z(n19119) );
  XNOR U2960 ( .A(n19483), .B(n19647), .Z(n19487) );
  XNOR U2961 ( .A(n19851), .B(n20015), .Z(n19855) );
  XNOR U2962 ( .A(n20219), .B(n20383), .Z(n20223) );
  XNOR U2963 ( .A(n20587), .B(n20751), .Z(n20591) );
  XNOR U2964 ( .A(n20955), .B(n21119), .Z(n20959) );
  XNOR U2965 ( .A(n21323), .B(n21487), .Z(n21327) );
  XNOR U2966 ( .A(n21691), .B(n21855), .Z(n21695) );
  XNOR U2967 ( .A(n22059), .B(n22223), .Z(n22063) );
  XNOR U2968 ( .A(n22427), .B(n22591), .Z(n22431) );
  XNOR U2969 ( .A(n22795), .B(n22959), .Z(n22799) );
  XNOR U2970 ( .A(n4852), .B(n5093), .Z(n4856) );
  XNOR U2971 ( .A(n3687), .B(n3987), .Z(n3691) );
  XNOR U2972 ( .A(n2923), .B(n3247), .Z(n2927) );
  XNOR U2973 ( .A(n4876), .B(n5087), .Z(n4880) );
  XNOR U2974 ( .A(n6407), .B(n6566), .Z(n6408) );
  XNOR U2975 ( .A(n7145), .B(n7310), .Z(n7153) );
  XNOR U2976 ( .A(n7892), .B(n8054), .Z(n7896) );
  XNOR U2977 ( .A(n8639), .B(n8798), .Z(n8640) );
  XNOR U2978 ( .A(n9377), .B(n9542), .Z(n9385) );
  XNOR U2979 ( .A(n10129), .B(n10411), .Z(n10133) );
  XNOR U2980 ( .A(n11398), .B(n11026), .Z(n11028) );
  XNOR U2981 ( .A(n11766), .B(n11395), .Z(n11397) );
  XNOR U2982 ( .A(n12128), .B(n12286), .Z(n12132) );
  XNOR U2983 ( .A(n12864), .B(n13022), .Z(n12868) );
  XNOR U2984 ( .A(n13968), .B(n14126), .Z(n13972) );
  XNOR U2985 ( .A(n15808), .B(n15966), .Z(n15812) );
  XNOR U2986 ( .A(n16544), .B(n16702), .Z(n16548) );
  XNOR U2987 ( .A(n4093), .B(n4351), .Z(n4097) );
  XNOR U2988 ( .A(n3332), .B(n3611), .Z(n3333) );
  XNOR U2989 ( .A(n2162), .B(n2505), .Z(n2166) );
  XNOR U2990 ( .A(n5264), .B(n5456), .Z(n5272) );
  XNOR U2991 ( .A(n13605), .B(n13757), .Z(n13609) );
  XNOR U2992 ( .A(n14709), .B(n14861), .Z(n14713) );
  XNOR U2993 ( .A(n15819), .B(n15448), .Z(n15450) );
  XNOR U2994 ( .A(n33456), .B(n33603), .Z(n33460) );
  XNOR U2995 ( .A(n33136), .B(n33280), .Z(n33140) );
  XNOR U2996 ( .A(n32789), .B(n32933), .Z(n32793) );
  XNOR U2997 ( .A(n32418), .B(n32565), .Z(n32422) );
  XNOR U2998 ( .A(n32026), .B(n32170), .Z(n32030) );
  XNOR U2999 ( .A(n31423), .B(n31575), .Z(n31427) );
  XNOR U3000 ( .A(n30967), .B(n31119), .Z(n30971) );
  XNOR U3001 ( .A(n30487), .B(n30639), .Z(n30491) );
  XNOR U3002 ( .A(n29983), .B(n30135), .Z(n29987) );
  XNOR U3003 ( .A(n29455), .B(n29607), .Z(n29459) );
  XNOR U3004 ( .A(n28903), .B(n29055), .Z(n28907) );
  XNOR U3005 ( .A(n28327), .B(n28479), .Z(n28331) );
  XNOR U3006 ( .A(n27727), .B(n27879), .Z(n27731) );
  XNOR U3007 ( .A(n27103), .B(n27255), .Z(n27107) );
  XNOR U3008 ( .A(n26455), .B(n26607), .Z(n26459) );
  XNOR U3009 ( .A(n25783), .B(n25935), .Z(n25787) );
  XNOR U3010 ( .A(n25087), .B(n25239), .Z(n25091) );
  XNOR U3011 ( .A(n24367), .B(n24519), .Z(n24371) );
  XNOR U3012 ( .A(n23546), .B(n23773), .Z(n23550) );
  XNOR U3013 ( .A(n4905), .B(n5080), .Z(n4909) );
  XNOR U3014 ( .A(n4083), .B(n4355), .Z(n4078) );
  XNOR U3015 ( .A(n3740), .B(n3974), .Z(n3744) );
  XNOR U3016 ( .A(n11776), .B(n11405), .Z(n11407) );
  XNOR U3017 ( .A(n16186), .B(n16332), .Z(n16190) );
  XNOR U3018 ( .A(n18026), .B(n18172), .Z(n18030) );
  XNOR U3019 ( .A(n18394), .B(n18540), .Z(n18398) );
  XNOR U3020 ( .A(n18762), .B(n18908), .Z(n18766) );
  XNOR U3021 ( .A(n19130), .B(n19276), .Z(n19134) );
  XNOR U3022 ( .A(n19498), .B(n19644), .Z(n19502) );
  XNOR U3023 ( .A(n19866), .B(n20012), .Z(n19870) );
  XNOR U3024 ( .A(n20234), .B(n20380), .Z(n20238) );
  XNOR U3025 ( .A(n20602), .B(n20748), .Z(n20606) );
  XNOR U3026 ( .A(n20970), .B(n21116), .Z(n20974) );
  XNOR U3027 ( .A(n21338), .B(n21484), .Z(n21342) );
  XNOR U3028 ( .A(n21706), .B(n21852), .Z(n21710) );
  XNOR U3029 ( .A(n22074), .B(n22220), .Z(n22078) );
  XNOR U3030 ( .A(n22442), .B(n22588), .Z(n22446) );
  XNOR U3031 ( .A(n22810), .B(n22956), .Z(n22814) );
  XNOR U3032 ( .A(n4489), .B(n4719), .Z(n4484) );
  XNOR U3033 ( .A(n2938), .B(n3244), .Z(n2942) );
  XNOR U3034 ( .A(n4929), .B(n5074), .Z(n4933) );
  XNOR U3035 ( .A(n6047), .B(n6191), .Z(n6055) );
  XNOR U3036 ( .A(n7159), .B(n7306), .Z(n7163) );
  XNOR U3037 ( .A(n7911), .B(n8051), .Z(n7906) );
  XNOR U3038 ( .A(n8651), .B(n8795), .Z(n8655) );
  XNOR U3039 ( .A(n9391), .B(n9538), .Z(n9395) );
  XNOR U3040 ( .A(n10148), .B(n10405), .Z(n10142) );
  XNOR U3041 ( .A(n11413), .B(n11041), .Z(n11043) );
  XNOR U3042 ( .A(n11781), .B(n11410), .Z(n11412) );
  XNOR U3043 ( .A(n12143), .B(n12283), .Z(n12147) );
  XNOR U3044 ( .A(n12511), .B(n12651), .Z(n12515) );
  XNOR U3045 ( .A(n13247), .B(n13387), .Z(n13251) );
  XNOR U3046 ( .A(n13983), .B(n14123), .Z(n13987) );
  XNOR U3047 ( .A(n15087), .B(n15227), .Z(n15091) );
  XNOR U3048 ( .A(n16927), .B(n17067), .Z(n16931) );
  XNOR U3049 ( .A(n17663), .B(n17803), .Z(n17667) );
  XNOR U3050 ( .A(n3769), .B(n3967), .Z(n3773) );
  XNOR U3051 ( .A(n3726), .B(n3978), .Z(n3734) );
  XNOR U3052 ( .A(n2177), .B(n2502), .Z(n2181) );
  XNOR U3053 ( .A(n1413), .B(n1761), .Z(n1417) );
  XNOR U3054 ( .A(n4518), .B(n4712), .Z(n4513) );
  XNOR U3055 ( .A(n5682), .B(n5817), .Z(n5683) );
  XNOR U3056 ( .A(n14724), .B(n14858), .Z(n14728) );
  XNOR U3057 ( .A(n15828), .B(n15962), .Z(n15832) );
  XNOR U3058 ( .A(n16938), .B(n16567), .Z(n16569) );
  XNOR U3059 ( .A(n34045), .B(n34171), .Z(n34049) );
  XNOR U3060 ( .A(n33770), .B(n33896), .Z(n33774) );
  XNOR U3061 ( .A(n33471), .B(n33600), .Z(n33475) );
  XNOR U3062 ( .A(n33151), .B(n33277), .Z(n33155) );
  XNOR U3063 ( .A(n32804), .B(n32930), .Z(n32808) );
  XNOR U3064 ( .A(n32433), .B(n32562), .Z(n32437) );
  XNOR U3065 ( .A(n32041), .B(n32167), .Z(n32045) );
  XNOR U3066 ( .A(n31438), .B(n31572), .Z(n31442) );
  XNOR U3067 ( .A(n30982), .B(n31116), .Z(n30986) );
  XNOR U3068 ( .A(n30502), .B(n30636), .Z(n30506) );
  XNOR U3069 ( .A(n29998), .B(n30132), .Z(n30002) );
  XNOR U3070 ( .A(n29470), .B(n29604), .Z(n29474) );
  XNOR U3071 ( .A(n28918), .B(n29052), .Z(n28922) );
  XNOR U3072 ( .A(n28342), .B(n28476), .Z(n28346) );
  XNOR U3073 ( .A(n27742), .B(n27876), .Z(n27746) );
  XNOR U3074 ( .A(n27118), .B(n27252), .Z(n27122) );
  XNOR U3075 ( .A(n26470), .B(n26604), .Z(n26474) );
  XNOR U3076 ( .A(n25798), .B(n25932), .Z(n25802) );
  XNOR U3077 ( .A(n25102), .B(n25236), .Z(n25106) );
  XNOR U3078 ( .A(n24382), .B(n24516), .Z(n24386) );
  XNOR U3079 ( .A(n23561), .B(n23770), .Z(n23565) );
  XNOR U3080 ( .A(n3755), .B(n3971), .Z(n3763) );
  XNOR U3081 ( .A(n4562), .B(n4700), .Z(n4566) );
  XNOR U3082 ( .A(n3798), .B(n3960), .Z(n3802) );
  XNOR U3083 ( .A(n11791), .B(n11420), .Z(n11422) );
  XNOR U3084 ( .A(n17305), .B(n17433), .Z(n17309) );
  XNOR U3085 ( .A(n19145), .B(n19273), .Z(n19149) );
  XNOR U3086 ( .A(n19513), .B(n19641), .Z(n19517) );
  XNOR U3087 ( .A(n19881), .B(n20009), .Z(n19885) );
  XNOR U3088 ( .A(n20249), .B(n20377), .Z(n20253) );
  XNOR U3089 ( .A(n20617), .B(n20745), .Z(n20621) );
  XNOR U3090 ( .A(n20985), .B(n21113), .Z(n20989) );
  XNOR U3091 ( .A(n21353), .B(n21481), .Z(n21357) );
  XNOR U3092 ( .A(n21721), .B(n21849), .Z(n21725) );
  XNOR U3093 ( .A(n22089), .B(n22217), .Z(n22093) );
  XNOR U3094 ( .A(n22457), .B(n22585), .Z(n22461) );
  XNOR U3095 ( .A(n22825), .B(n22953), .Z(n22829) );
  XNOR U3096 ( .A(n4547), .B(n4705), .Z(n4542) );
  XNOR U3097 ( .A(n2589), .B(n2866), .Z(n2593) );
  XNOR U3098 ( .A(n1824), .B(n2124), .Z(n1828) );
  XNOR U3099 ( .A(n2574), .B(n2871), .Z(n2569) );
  XNOR U3100 ( .A(n6810), .B(n6928), .Z(n6805) );
  XNOR U3101 ( .A(n7921), .B(n8047), .Z(n7925) );
  XNOR U3102 ( .A(n8668), .B(n8791), .Z(n8669) );
  XNOR U3103 ( .A(n9406), .B(n9535), .Z(n9414) );
  XNOR U3104 ( .A(n10158), .B(n10400), .Z(n10162) );
  XNOR U3105 ( .A(n11428), .B(n11056), .Z(n11058) );
  XNOR U3106 ( .A(n11796), .B(n11425), .Z(n11427) );
  XNOR U3107 ( .A(n12158), .B(n12280), .Z(n12162) );
  XNOR U3108 ( .A(n12526), .B(n12648), .Z(n12530) );
  XNOR U3109 ( .A(n13262), .B(n13384), .Z(n13266) );
  XNOR U3110 ( .A(n13630), .B(n13752), .Z(n13634) );
  XNOR U3111 ( .A(n14366), .B(n14488), .Z(n14370) );
  XNOR U3112 ( .A(n15102), .B(n15224), .Z(n15106) );
  XNOR U3113 ( .A(n16206), .B(n16328), .Z(n16210) );
  XNOR U3114 ( .A(n18046), .B(n18168), .Z(n18050) );
  XNOR U3115 ( .A(n18782), .B(n18904), .Z(n18786) );
  XNOR U3116 ( .A(n3784), .B(n3964), .Z(n3792) );
  XNOR U3117 ( .A(n2981), .B(n3235), .Z(n2976) );
  XNOR U3118 ( .A(n1810), .B(n2128), .Z(n1818) );
  XNOR U3119 ( .A(n1046), .B(n1388), .Z(n1050) );
  XNOR U3120 ( .A(n2618), .B(n2859), .Z(n2622) );
  XNOR U3121 ( .A(n1853), .B(n2117), .Z(n1857) );
  XNOR U3122 ( .A(n5694), .B(n5814), .Z(n5698) );
  XNOR U3123 ( .A(n6438), .B(n6558), .Z(n6442) );
  XNOR U3124 ( .A(n15843), .B(n15959), .Z(n15847) );
  XNOR U3125 ( .A(n16947), .B(n17063), .Z(n16951) );
  XNOR U3126 ( .A(n18057), .B(n17686), .Z(n17688) );
  XNOR U3127 ( .A(n34308), .B(n34419), .Z(n34312) );
  XNOR U3128 ( .A(n34060), .B(n34168), .Z(n34064) );
  XNOR U3129 ( .A(n33785), .B(n33893), .Z(n33789) );
  XNOR U3130 ( .A(n33486), .B(n33597), .Z(n33490) );
  XNOR U3131 ( .A(n33166), .B(n33274), .Z(n33170) );
  XNOR U3132 ( .A(n32819), .B(n32927), .Z(n32823) );
  XNOR U3133 ( .A(n32448), .B(n32559), .Z(n32452) );
  XNOR U3134 ( .A(n32056), .B(n32164), .Z(n32060) );
  XNOR U3135 ( .A(n31453), .B(n31569), .Z(n31457) );
  XNOR U3136 ( .A(n30997), .B(n31113), .Z(n31001) );
  XNOR U3137 ( .A(n30517), .B(n30633), .Z(n30521) );
  XNOR U3138 ( .A(n30013), .B(n30129), .Z(n30017) );
  XNOR U3139 ( .A(n29485), .B(n29601), .Z(n29489) );
  XNOR U3140 ( .A(n28933), .B(n29049), .Z(n28937) );
  XNOR U3141 ( .A(n28357), .B(n28473), .Z(n28361) );
  XNOR U3142 ( .A(n27757), .B(n27873), .Z(n27761) );
  XNOR U3143 ( .A(n27133), .B(n27249), .Z(n27137) );
  XNOR U3144 ( .A(n26485), .B(n26601), .Z(n26489) );
  XNOR U3145 ( .A(n25813), .B(n25929), .Z(n25817) );
  XNOR U3146 ( .A(n25117), .B(n25233), .Z(n25121) );
  XNOR U3147 ( .A(n24397), .B(n24513), .Z(n24401) );
  XNOR U3148 ( .A(n23576), .B(n23767), .Z(n23580) );
  XNOR U3149 ( .A(n3832), .B(n3952), .Z(n3836) );
  XNOR U3150 ( .A(n3010), .B(n3228), .Z(n3005) );
  XNOR U3151 ( .A(n3813), .B(n3957), .Z(n3821) );
  XNOR U3152 ( .A(n4581), .B(n4695), .Z(n4585) );
  XNOR U3153 ( .A(n5331), .B(n5441), .Z(n5326) );
  XNOR U3154 ( .A(n11806), .B(n11435), .Z(n11437) );
  XNOR U3155 ( .A(n18424), .B(n18534), .Z(n18428) );
  XNOR U3156 ( .A(n20264), .B(n20374), .Z(n20268) );
  XNOR U3157 ( .A(n20632), .B(n20742), .Z(n20636) );
  XNOR U3158 ( .A(n21000), .B(n21110), .Z(n21004) );
  XNOR U3159 ( .A(n21368), .B(n21478), .Z(n21372) );
  XNOR U3160 ( .A(n21736), .B(n21846), .Z(n21740) );
  XNOR U3161 ( .A(n22104), .B(n22214), .Z(n22108) );
  XNOR U3162 ( .A(n22472), .B(n22582), .Z(n22476) );
  XNOR U3163 ( .A(n22840), .B(n22950), .Z(n22844) );
  XNOR U3164 ( .A(n2647), .B(n2852), .Z(n2651) );
  XNOR U3165 ( .A(n1882), .B(n2110), .Z(n1886) );
  XNOR U3166 ( .A(n1839), .B(n2121), .Z(n1847) );
  XNOR U3167 ( .A(n1075), .B(n1381), .Z(n1079) );
  XNOR U3168 ( .A(n7566), .B(n7671), .Z(n7567) );
  XNOR U3169 ( .A(n8680), .B(n8788), .Z(n8684) );
  XNOR U3170 ( .A(n9420), .B(n9531), .Z(n9424) );
  XNOR U3171 ( .A(n10177), .B(n10394), .Z(n10171) );
  XNOR U3172 ( .A(n11443), .B(n11071), .Z(n11073) );
  XNOR U3173 ( .A(n11811), .B(n11440), .Z(n11442) );
  XNOR U3174 ( .A(n12173), .B(n12277), .Z(n12177) );
  XNOR U3175 ( .A(n12541), .B(n12645), .Z(n12545) );
  XNOR U3176 ( .A(n13277), .B(n13381), .Z(n13281) );
  XNOR U3177 ( .A(n13645), .B(n13749), .Z(n13649) );
  XNOR U3178 ( .A(n14381), .B(n14485), .Z(n14385) );
  XNOR U3179 ( .A(n14749), .B(n14853), .Z(n14753) );
  XNOR U3180 ( .A(n15485), .B(n15589), .Z(n15489) );
  XNOR U3181 ( .A(n16221), .B(n16325), .Z(n16225) );
  XNOR U3182 ( .A(n17325), .B(n17429), .Z(n17329) );
  XNOR U3183 ( .A(n19165), .B(n19269), .Z(n19169) );
  XNOR U3184 ( .A(n19901), .B(n20005), .Z(n19905) );
  XNOR U3185 ( .A(n3039), .B(n3221), .Z(n3034) );
  XNOR U3186 ( .A(n1065), .B(n1385), .Z(n1060) );
  XNOR U3187 ( .A(n1868), .B(n2114), .Z(n1876) );
  XNOR U3188 ( .A(n1104), .B(n1374), .Z(n1108) );
  XNOR U3189 ( .A(n2676), .B(n2845), .Z(n2680) );
  XNOR U3190 ( .A(n1911), .B(n2103), .Z(n1915) );
  XNOR U3191 ( .A(n6453), .B(n6555), .Z(n6461) );
  XNOR U3192 ( .A(n7193), .B(n7298), .Z(n7197) );
  XNOR U3193 ( .A(n16962), .B(n17060), .Z(n16966) );
  XNOR U3194 ( .A(n18066), .B(n18164), .Z(n18070) );
  XNOR U3195 ( .A(n19176), .B(n18805), .Z(n18807) );
  XNOR U3196 ( .A(n21016), .B(n20645), .Z(n20647) );
  XNOR U3197 ( .A(n34753), .B(n34843), .Z(n34757) );
  XNOR U3198 ( .A(n34550), .B(n34640), .Z(n34554) );
  XNOR U3199 ( .A(n34323), .B(n34416), .Z(n34327) );
  XNOR U3200 ( .A(n34075), .B(n34165), .Z(n34079) );
  XNOR U3201 ( .A(n33800), .B(n33890), .Z(n33804) );
  XNOR U3202 ( .A(n33501), .B(n33594), .Z(n33505) );
  XNOR U3203 ( .A(n33181), .B(n33271), .Z(n33185) );
  XNOR U3204 ( .A(n32834), .B(n32924), .Z(n32838) );
  XNOR U3205 ( .A(n32463), .B(n32556), .Z(n32467) );
  XNOR U3206 ( .A(n32071), .B(n32161), .Z(n32075) );
  XNOR U3207 ( .A(n31468), .B(n31566), .Z(n31472) );
  XNOR U3208 ( .A(n31012), .B(n31110), .Z(n31016) );
  XNOR U3209 ( .A(n30532), .B(n30630), .Z(n30536) );
  XNOR U3210 ( .A(n30028), .B(n30126), .Z(n30032) );
  XNOR U3211 ( .A(n29500), .B(n29598), .Z(n29504) );
  XNOR U3212 ( .A(n28948), .B(n29046), .Z(n28952) );
  XNOR U3213 ( .A(n28372), .B(n28470), .Z(n28376) );
  XNOR U3214 ( .A(n27772), .B(n27870), .Z(n27776) );
  XNOR U3215 ( .A(n27148), .B(n27246), .Z(n27152) );
  XNOR U3216 ( .A(n26500), .B(n26598), .Z(n26504) );
  XNOR U3217 ( .A(n25828), .B(n25926), .Z(n25832) );
  XNOR U3218 ( .A(n25132), .B(n25230), .Z(n25136) );
  XNOR U3219 ( .A(n24412), .B(n24510), .Z(n24416) );
  XNOR U3220 ( .A(n23591), .B(n23764), .Z(n23595) );
  XNOR U3221 ( .A(n3068), .B(n3214), .Z(n3063) );
  XNOR U3222 ( .A(n3854), .B(n3947), .Z(n3855) );
  XNOR U3223 ( .A(n4596), .B(n4692), .Z(n4604) );
  XNOR U3224 ( .A(n5341), .B(n5437), .Z(n5345) );
  XNOR U3225 ( .A(n6088), .B(n6181), .Z(n6089) );
  XNOR U3226 ( .A(n11821), .B(n11450), .Z(n11452) );
  XNOR U3227 ( .A(n19543), .B(n19635), .Z(n19547) );
  XNOR U3228 ( .A(n21383), .B(n21475), .Z(n21387) );
  XNOR U3229 ( .A(n21751), .B(n21843), .Z(n21755) );
  XNOR U3230 ( .A(n22119), .B(n22211), .Z(n22123) );
  XNOR U3231 ( .A(n22487), .B(n22579), .Z(n22491) );
  XNOR U3232 ( .A(n22855), .B(n22947), .Z(n22859) );
  XNOR U3233 ( .A(n2705), .B(n2838), .Z(n2709) );
  XNOR U3234 ( .A(n1940), .B(n2096), .Z(n1944) );
  XNOR U3235 ( .A(n1897), .B(n2107), .Z(n1905) );
  XNOR U3236 ( .A(n1133), .B(n1367), .Z(n1137) );
  XNOR U3237 ( .A(n1094), .B(n1378), .Z(n1089) );
  XNOR U3238 ( .A(n2729), .B(n2832), .Z(n2733) );
  XNOR U3239 ( .A(n8322), .B(n8412), .Z(n8326) );
  XNOR U3240 ( .A(n9435), .B(n9528), .Z(n9443) );
  XNOR U3241 ( .A(n10187), .B(n10389), .Z(n10191) );
  XNOR U3242 ( .A(n11458), .B(n11086), .Z(n11088) );
  XNOR U3243 ( .A(n11826), .B(n11455), .Z(n11457) );
  XNOR U3244 ( .A(n12188), .B(n12274), .Z(n12192) );
  XNOR U3245 ( .A(n12556), .B(n12642), .Z(n12560) );
  XNOR U3246 ( .A(n13292), .B(n13378), .Z(n13296) );
  XNOR U3247 ( .A(n13660), .B(n13746), .Z(n13664) );
  XNOR U3248 ( .A(n14396), .B(n14482), .Z(n14400) );
  XNOR U3249 ( .A(n14764), .B(n14850), .Z(n14768) );
  XNOR U3250 ( .A(n15500), .B(n15586), .Z(n15504) );
  XNOR U3251 ( .A(n15868), .B(n15954), .Z(n15872) );
  XNOR U3252 ( .A(n16604), .B(n16690), .Z(n16608) );
  XNOR U3253 ( .A(n17340), .B(n17426), .Z(n17344) );
  XNOR U3254 ( .A(n18444), .B(n18530), .Z(n18448) );
  XNOR U3255 ( .A(n20284), .B(n20370), .Z(n20288) );
  XNOR U3256 ( .A(n3097), .B(n3207), .Z(n3092) );
  XNOR U3257 ( .A(n1123), .B(n1371), .Z(n1118) );
  XNOR U3258 ( .A(n1926), .B(n2100), .Z(n1934) );
  XNOR U3259 ( .A(n1162), .B(n1360), .Z(n1166) );
  XNOR U3260 ( .A(n1969), .B(n2089), .Z(n1973) );
  XNOR U3261 ( .A(n7212), .B(n7295), .Z(n7207) );
  XNOR U3262 ( .A(n7955), .B(n8039), .Z(n7959) );
  XNOR U3263 ( .A(n18081), .B(n18161), .Z(n18085) );
  XNOR U3264 ( .A(n19185), .B(n19265), .Z(n19189) );
  XNOR U3265 ( .A(n20295), .B(n19924), .Z(n19926) );
  XNOR U3266 ( .A(n21767), .B(n21396), .Z(n21398) );
  XNOR U3267 ( .A(n22135), .B(n21764), .Z(n21766) );
  XNOR U3268 ( .A(n34944), .B(n35019), .Z(n34948) );
  XNOR U3269 ( .A(n34768), .B(n34840), .Z(n34772) );
  XNOR U3270 ( .A(n34565), .B(n34637), .Z(n34569) );
  XNOR U3271 ( .A(n34338), .B(n34413), .Z(n34342) );
  XNOR U3272 ( .A(n34090), .B(n34162), .Z(n34094) );
  XNOR U3273 ( .A(n33815), .B(n33887), .Z(n33819) );
  XNOR U3274 ( .A(n33516), .B(n33591), .Z(n33520) );
  XNOR U3275 ( .A(n33196), .B(n33268), .Z(n33200) );
  XNOR U3276 ( .A(n32849), .B(n32921), .Z(n32853) );
  XNOR U3277 ( .A(n32478), .B(n32553), .Z(n32482) );
  XNOR U3278 ( .A(n32086), .B(n32158), .Z(n32090) );
  XNOR U3279 ( .A(n31483), .B(n31563), .Z(n31487) );
  XNOR U3280 ( .A(n31027), .B(n31107), .Z(n31031) );
  XNOR U3281 ( .A(n30547), .B(n30627), .Z(n30551) );
  XNOR U3282 ( .A(n30043), .B(n30123), .Z(n30047) );
  XNOR U3283 ( .A(n29515), .B(n29595), .Z(n29519) );
  XNOR U3284 ( .A(n28963), .B(n29043), .Z(n28967) );
  XNOR U3285 ( .A(n28387), .B(n28467), .Z(n28391) );
  XNOR U3286 ( .A(n27787), .B(n27867), .Z(n27791) );
  XNOR U3287 ( .A(n27163), .B(n27243), .Z(n27167) );
  XNOR U3288 ( .A(n26515), .B(n26595), .Z(n26519) );
  XNOR U3289 ( .A(n25843), .B(n25923), .Z(n25847) );
  XNOR U3290 ( .A(n25147), .B(n25227), .Z(n25151) );
  XNOR U3291 ( .A(n24427), .B(n24507), .Z(n24431) );
  XNOR U3292 ( .A(n23606), .B(n23761), .Z(n23610) );
  XNOR U3293 ( .A(n3866), .B(n3944), .Z(n3870) );
  XNOR U3294 ( .A(n4610), .B(n4688), .Z(n4614) );
  XNOR U3295 ( .A(n5360), .B(n5434), .Z(n5355) );
  XNOR U3296 ( .A(n6100), .B(n6178), .Z(n6104) );
  XNOR U3297 ( .A(n6844), .B(n6918), .Z(n6848) );
  XNOR U3298 ( .A(n11836), .B(n11465), .Z(n11467) );
  XNOR U3299 ( .A(n22502), .B(n22576), .Z(n22506) );
  XNOR U3300 ( .A(n22870), .B(n22944), .Z(n22874) );
  XNOR U3301 ( .A(n1955), .B(n2093), .Z(n1963) );
  XNOR U3302 ( .A(n1191), .B(n1353), .Z(n1195) );
  XNOR U3303 ( .A(n1152), .B(n1364), .Z(n1147) );
  XNOR U3304 ( .A(n2748), .B(n2829), .Z(n2743) );
  XNOR U3305 ( .A(n9081), .B(n9149), .Z(n9085) );
  XNOR U3306 ( .A(n10206), .B(n10383), .Z(n10200) );
  XNOR U3307 ( .A(n11473), .B(n11101), .Z(n11103) );
  XNOR U3308 ( .A(n11841), .B(n11470), .Z(n11472) );
  XNOR U3309 ( .A(n12203), .B(n12271), .Z(n12207) );
  XNOR U3310 ( .A(n12571), .B(n12639), .Z(n12575) );
  XNOR U3311 ( .A(n13307), .B(n13375), .Z(n13311) );
  XNOR U3312 ( .A(n13675), .B(n13743), .Z(n13679) );
  XNOR U3313 ( .A(n14411), .B(n14479), .Z(n14415) );
  XNOR U3314 ( .A(n14779), .B(n14847), .Z(n14783) );
  XNOR U3315 ( .A(n15515), .B(n15583), .Z(n15519) );
  XNOR U3316 ( .A(n15883), .B(n15951), .Z(n15887) );
  XNOR U3317 ( .A(n16619), .B(n16687), .Z(n16623) );
  XNOR U3318 ( .A(n16987), .B(n17055), .Z(n16991) );
  XNOR U3319 ( .A(n17723), .B(n17791), .Z(n17727) );
  XNOR U3320 ( .A(n18459), .B(n18527), .Z(n18463) );
  XNOR U3321 ( .A(n19563), .B(n19631), .Z(n19567) );
  XNOR U3322 ( .A(n21035), .B(n21103), .Z(n21039) );
  XNOR U3323 ( .A(n1621), .B(n1711), .Z(n1625) );
  XNOR U3324 ( .A(n1181), .B(n1357), .Z(n1176) );
  XNOR U3325 ( .A(n1984), .B(n2086), .Z(n1992) );
  XNOR U3326 ( .A(n1220), .B(n1346), .Z(n1224) );
  XNOR U3327 ( .A(n7972), .B(n8035), .Z(n7973) );
  XNOR U3328 ( .A(n8714), .B(n8780), .Z(n8722) );
  XNOR U3329 ( .A(n19200), .B(n19262), .Z(n19204) );
  XNOR U3330 ( .A(n20304), .B(n20366), .Z(n20308) );
  XNOR U3331 ( .A(n21414), .B(n21043), .Z(n21045) );
  XNOR U3332 ( .A(n22150), .B(n21779), .Z(n21781) );
  XNOR U3333 ( .A(n22518), .B(n22147), .Z(n22149) );
  XNOR U3334 ( .A(n22886), .B(n22515), .Z(n22517) );
  XNOR U3335 ( .A(n23254), .B(n22883), .Z(n22885) );
  XNOR U3336 ( .A(n35245), .B(n35299), .Z(n35249) );
  XNOR U3337 ( .A(n35114), .B(n35168), .Z(n35118) );
  XNOR U3338 ( .A(n34959), .B(n35016), .Z(n34963) );
  XNOR U3339 ( .A(n34783), .B(n34837), .Z(n34787) );
  XNOR U3340 ( .A(n34580), .B(n34634), .Z(n34584) );
  XNOR U3341 ( .A(n34353), .B(n34410), .Z(n34357) );
  XNOR U3342 ( .A(n34105), .B(n34159), .Z(n34109) );
  XNOR U3343 ( .A(n33830), .B(n33884), .Z(n33834) );
  XNOR U3344 ( .A(n33531), .B(n33588), .Z(n33535) );
  XNOR U3345 ( .A(n33211), .B(n33265), .Z(n33215) );
  XNOR U3346 ( .A(n32864), .B(n32918), .Z(n32868) );
  XNOR U3347 ( .A(n32493), .B(n32550), .Z(n32497) );
  XNOR U3348 ( .A(n32101), .B(n32155), .Z(n32105) );
  XNOR U3349 ( .A(n31498), .B(n31560), .Z(n31502) );
  XNOR U3350 ( .A(n31042), .B(n31104), .Z(n31046) );
  XNOR U3351 ( .A(n30562), .B(n30624), .Z(n30566) );
  XNOR U3352 ( .A(n30058), .B(n30120), .Z(n30062) );
  XNOR U3353 ( .A(n29530), .B(n29592), .Z(n29534) );
  XNOR U3354 ( .A(n28978), .B(n29040), .Z(n28982) );
  XNOR U3355 ( .A(n28402), .B(n28464), .Z(n28406) );
  XNOR U3356 ( .A(n27802), .B(n27864), .Z(n27806) );
  XNOR U3357 ( .A(n27178), .B(n27240), .Z(n27182) );
  XNOR U3358 ( .A(n26530), .B(n26592), .Z(n26534) );
  XNOR U3359 ( .A(n25858), .B(n25920), .Z(n25862) );
  XNOR U3360 ( .A(n25162), .B(n25224), .Z(n25166) );
  XNOR U3361 ( .A(n24442), .B(n24504), .Z(n24446) );
  XNOR U3362 ( .A(n23621), .B(n23758), .Z(n23625) );
  XNOR U3363 ( .A(n887), .B(n965), .Z(n891) );
  XNOR U3364 ( .A(n3136), .B(n3196), .Z(n3140) );
  XNOR U3365 ( .A(n4625), .B(n4685), .Z(n4633) );
  XNOR U3366 ( .A(n5370), .B(n5430), .Z(n5374) );
  XNOR U3367 ( .A(n6117), .B(n6174), .Z(n6118) );
  XNOR U3368 ( .A(n6859), .B(n6915), .Z(n6867) );
  XNOR U3369 ( .A(n11851), .B(n11480), .Z(n11482) );
  XNOR U3370 ( .A(n2013), .B(n2079), .Z(n2017) );
  XNOR U3371 ( .A(n1210), .B(n1350), .Z(n1205) );
  XNOR U3372 ( .A(n3885), .B(n3939), .Z(n3889) );
  XNOR U3373 ( .A(n9839), .B(n9894), .Z(n9843) );
  XNOR U3374 ( .A(n11488), .B(n11116), .Z(n11118) );
  XNOR U3375 ( .A(n11856), .B(n11485), .Z(n11487) );
  XNOR U3376 ( .A(n12218), .B(n12268), .Z(n12222) );
  XNOR U3377 ( .A(n12586), .B(n12636), .Z(n12590) );
  XNOR U3378 ( .A(n13322), .B(n13372), .Z(n13326) );
  XNOR U3379 ( .A(n13690), .B(n13740), .Z(n13694) );
  XNOR U3380 ( .A(n14426), .B(n14476), .Z(n14430) );
  XNOR U3381 ( .A(n14794), .B(n14844), .Z(n14798) );
  XNOR U3382 ( .A(n15530), .B(n15580), .Z(n15534) );
  XNOR U3383 ( .A(n15898), .B(n15948), .Z(n15902) );
  XNOR U3384 ( .A(n16634), .B(n16684), .Z(n16638) );
  XNOR U3385 ( .A(n17002), .B(n17052), .Z(n17006) );
  XNOR U3386 ( .A(n17738), .B(n17788), .Z(n17742) );
  XNOR U3387 ( .A(n18106), .B(n18156), .Z(n18110) );
  XNOR U3388 ( .A(n18842), .B(n18892), .Z(n18846) );
  XNOR U3389 ( .A(n19578), .B(n19628), .Z(n19582) );
  XNOR U3390 ( .A(n20682), .B(n20732), .Z(n20686) );
  XNOR U3391 ( .A(n1254), .B(n1338), .Z(n1258) );
  XNOR U3392 ( .A(n1239), .B(n1343), .Z(n1234) );
  XNOR U3393 ( .A(n2028), .B(n2076), .Z(n2032) );
  XNOR U3394 ( .A(n2773), .B(n2822), .Z(n2777) );
  XNOR U3395 ( .A(n8356), .B(n8404), .Z(n8360) );
  XNOR U3396 ( .A(n9473), .B(n9520), .Z(n9468) );
  XNOR U3397 ( .A(n20319), .B(n20363), .Z(n20323) );
  XNOR U3398 ( .A(n21423), .B(n21467), .Z(n21427) );
  XNOR U3399 ( .A(n22533), .B(n22162), .Z(n22164) );
  XNOR U3400 ( .A(n22901), .B(n22530), .Z(n22532) );
  XNOR U3401 ( .A(n23269), .B(n22898), .Z(n22900) );
  XNOR U3402 ( .A(n23263), .B(n23307), .Z(n23267) );
  XNOR U3403 ( .A(n35410), .B(n35446), .Z(n35414) );
  XNOR U3404 ( .A(n35315), .B(n35351), .Z(n35319) );
  XNOR U3405 ( .A(n35196), .B(n35235), .Z(n35200) );
  XNOR U3406 ( .A(n35056), .B(n35092), .Z(n35060) );
  XNOR U3407 ( .A(n34889), .B(n34925), .Z(n34893) );
  XNOR U3408 ( .A(n34698), .B(n34737), .Z(n34702) );
  XNOR U3409 ( .A(n34486), .B(n34522), .Z(n34490) );
  XNOR U3410 ( .A(n34247), .B(n34283), .Z(n34251) );
  XNOR U3411 ( .A(n33984), .B(n34023), .Z(n33988) );
  XNOR U3412 ( .A(n33700), .B(n33736), .Z(n33704) );
  XNOR U3413 ( .A(n33389), .B(n33425), .Z(n33393) );
  XNOR U3414 ( .A(n33054), .B(n33093), .Z(n33058) );
  XNOR U3415 ( .A(n32698), .B(n32734), .Z(n32702) );
  XNOR U3416 ( .A(n32315), .B(n32351), .Z(n32319) );
  XNOR U3417 ( .A(n31732), .B(n31947), .Z(n31736) );
  XNOR U3418 ( .A(n31288), .B(n31332), .Z(n31292) );
  XNOR U3419 ( .A(n30820), .B(n30864), .Z(n30824) );
  XNOR U3420 ( .A(n30328), .B(n30372), .Z(n30332) );
  XNOR U3421 ( .A(n29812), .B(n29856), .Z(n29816) );
  XNOR U3422 ( .A(n29272), .B(n29316), .Z(n29276) );
  XNOR U3423 ( .A(n28708), .B(n28752), .Z(n28712) );
  XNOR U3424 ( .A(n28120), .B(n28164), .Z(n28124) );
  XNOR U3425 ( .A(n27508), .B(n27552), .Z(n27512) );
  XNOR U3426 ( .A(n26872), .B(n26916), .Z(n26876) );
  XNOR U3427 ( .A(n26212), .B(n26256), .Z(n26216) );
  XNOR U3428 ( .A(n25528), .B(n25572), .Z(n25532) );
  XNOR U3429 ( .A(n24820), .B(n24864), .Z(n24824) );
  XNOR U3430 ( .A(n24085), .B(n24129), .Z(n24089) );
  XNOR U3431 ( .A(n1284), .B(n1332), .Z(n1288) );
  XNOR U3432 ( .A(n3523), .B(n3565), .Z(n3527) );
  XNOR U3433 ( .A(n5014), .B(n5054), .Z(n5015) );
  XNOR U3434 ( .A(n5757), .B(n5799), .Z(n5765) );
  XNOR U3435 ( .A(n6501), .B(n6543), .Z(n6505) );
  XNOR U3436 ( .A(n7244), .B(n7286), .Z(n7245) );
  XNOR U3437 ( .A(n7989), .B(n8031), .Z(n7997) );
  XNOR U3438 ( .A(n9105), .B(n9143), .Z(n9109) );
  XNOR U3439 ( .A(n11129), .B(n10758), .Z(n10760) );
  XNOR U3440 ( .A(n11866), .B(n11495), .Z(n11497) );
  XNOR U3441 ( .A(n21434), .B(n21063), .Z(n21065) );
  XNOR U3442 ( .A(n4644), .B(n4680), .Z(n4648) );
  XNOR U3443 ( .A(n11871), .B(n11500), .Z(n11502) );
  XNOR U3444 ( .A(n12233), .B(n12265), .Z(n12237) );
  XNOR U3445 ( .A(n12601), .B(n12633), .Z(n12605) );
  XNOR U3446 ( .A(n13337), .B(n13369), .Z(n13341) );
  XNOR U3447 ( .A(n13705), .B(n13737), .Z(n13709) );
  XNOR U3448 ( .A(n14441), .B(n14473), .Z(n14445) );
  XNOR U3449 ( .A(n14809), .B(n14841), .Z(n14813) );
  XNOR U3450 ( .A(n15545), .B(n15577), .Z(n15549) );
  XNOR U3451 ( .A(n15913), .B(n15945), .Z(n15917) );
  XNOR U3452 ( .A(n16649), .B(n16681), .Z(n16653) );
  XNOR U3453 ( .A(n17017), .B(n17049), .Z(n17021) );
  XNOR U3454 ( .A(n17753), .B(n17785), .Z(n17757) );
  XNOR U3455 ( .A(n18121), .B(n18153), .Z(n18125) );
  XNOR U3456 ( .A(n18857), .B(n18889), .Z(n18861) );
  XNOR U3457 ( .A(n19225), .B(n19257), .Z(n19229) );
  XNOR U3458 ( .A(n19961), .B(n19993), .Z(n19965) );
  XNOR U3459 ( .A(n20697), .B(n20729), .Z(n20701) );
  XNOR U3460 ( .A(n21801), .B(n21833), .Z(n21805) );
  XNOR U3461 ( .A(n23646), .B(n23753), .Z(n23650) );
  XNOR U3462 ( .A(n1671), .B(n1701), .Z(n1675) );
  XNOR U3463 ( .A(n2788), .B(n2819), .Z(n2792) );
  XNOR U3464 ( .A(n11133), .B(n11159), .Z(n11137) );
  XNOR U3465 ( .A(n21438), .B(n21464), .Z(n21442) );
  XNOR U3466 ( .A(n22542), .B(n22568), .Z(n22546) );
  XNOR U3467 ( .A(n35521), .B(n35539), .Z(n35525) );
  XNOR U3468 ( .A(n35462), .B(n35480), .Z(n35466) );
  XNOR U3469 ( .A(n35379), .B(n35400), .Z(n35383) );
  XNOR U3470 ( .A(n35275), .B(n35293), .Z(n35279) );
  XNOR U3471 ( .A(n35144), .B(n35162), .Z(n35148) );
  XNOR U3472 ( .A(n34989), .B(n35010), .Z(n34993) );
  XNOR U3473 ( .A(n34813), .B(n34831), .Z(n34817) );
  XNOR U3474 ( .A(n34610), .B(n34628), .Z(n34614) );
  XNOR U3475 ( .A(n34383), .B(n34404), .Z(n34387) );
  XNOR U3476 ( .A(n34135), .B(n34153), .Z(n34139) );
  XNOR U3477 ( .A(n33860), .B(n33878), .Z(n33864) );
  XNOR U3478 ( .A(n33561), .B(n33582), .Z(n33565) );
  XNOR U3479 ( .A(n33241), .B(n33259), .Z(n33245) );
  XNOR U3480 ( .A(n32894), .B(n32912), .Z(n32898) );
  XNOR U3481 ( .A(n32523), .B(n32544), .Z(n32527) );
  XNOR U3482 ( .A(n32131), .B(n32149), .Z(n32135) );
  XNOR U3483 ( .A(n31528), .B(n31554), .Z(n31532) );
  XNOR U3484 ( .A(n31072), .B(n31098), .Z(n31076) );
  XNOR U3485 ( .A(n30592), .B(n30618), .Z(n30596) );
  XNOR U3486 ( .A(n30088), .B(n30114), .Z(n30092) );
  XNOR U3487 ( .A(n29560), .B(n29586), .Z(n29564) );
  XNOR U3488 ( .A(n29008), .B(n29034), .Z(n29012) );
  XNOR U3489 ( .A(n28432), .B(n28458), .Z(n28436) );
  XNOR U3490 ( .A(n27832), .B(n27858), .Z(n27836) );
  XNOR U3491 ( .A(n27208), .B(n27234), .Z(n27212) );
  XNOR U3492 ( .A(n26560), .B(n26586), .Z(n26564) );
  XNOR U3493 ( .A(n25888), .B(n25914), .Z(n25892) );
  XNOR U3494 ( .A(n25192), .B(n25218), .Z(n25196) );
  XNOR U3495 ( .A(n24472), .B(n24498), .Z(n24476) );
  XNOR U3496 ( .A(n1304), .B(n1328), .Z(n1308) );
  XNOR U3497 ( .A(n2420), .B(n2444), .Z(n2424) );
  XNOR U3498 ( .A(n3538), .B(n3562), .Z(n3542) );
  XNOR U3499 ( .A(n4282), .B(n4306), .Z(n4286) );
  XNOR U3500 ( .A(n5771), .B(n5795), .Z(n5775) );
  XNOR U3501 ( .A(n6520), .B(n6540), .Z(n6515) );
  XNOR U3502 ( .A(n7256), .B(n7283), .Z(n7260) );
  XNOR U3503 ( .A(n8003), .B(n8027), .Z(n8007) );
  XNOR U3504 ( .A(n9120), .B(n9140), .Z(n9128) );
  XNOR U3505 ( .A(n10240), .B(n10369), .Z(n10244) );
  XNOR U3506 ( .A(n21449), .B(n21078), .Z(n21080) );
  XNOR U3507 ( .A(n23283), .B(n23303), .Z(n23287) );
  XNOR U3508 ( .A(n5031), .B(n5050), .Z(n5039) );
  XNOR U3509 ( .A(n9868), .B(n9886), .Z(n9877) );
  XNOR U3510 ( .A(n11518), .B(n11146), .Z(n11148) );
  XNOR U3511 ( .A(n11512), .B(n11526), .Z(n11516) );
  XNOR U3512 ( .A(n12622), .B(n12251), .Z(n12253) );
  XNOR U3513 ( .A(n12616), .B(n12630), .Z(n12620) );
  XNOR U3514 ( .A(n13726), .B(n13355), .Z(n13357) );
  XNOR U3515 ( .A(n13720), .B(n13734), .Z(n13724) );
  XNOR U3516 ( .A(n14830), .B(n14459), .Z(n14461) );
  XNOR U3517 ( .A(n14824), .B(n14838), .Z(n14828) );
  XNOR U3518 ( .A(n15934), .B(n15563), .Z(n15565) );
  XNOR U3519 ( .A(n15928), .B(n15942), .Z(n15932) );
  XNOR U3520 ( .A(n17038), .B(n16667), .Z(n16669) );
  XNOR U3521 ( .A(n17032), .B(n17046), .Z(n17036) );
  XNOR U3522 ( .A(n18142), .B(n17771), .Z(n17773) );
  XNOR U3523 ( .A(n18136), .B(n18150), .Z(n18140) );
  XNOR U3524 ( .A(n19246), .B(n18875), .Z(n18877) );
  XNOR U3525 ( .A(n19240), .B(n19254), .Z(n19244) );
  XNOR U3526 ( .A(n20350), .B(n19979), .Z(n19981) );
  XNOR U3527 ( .A(n20344), .B(n20358), .Z(n20348) );
  XNOR U3528 ( .A(n21454), .B(n21083), .Z(n21085) );
  XNOR U3529 ( .A(n21816), .B(n21830), .Z(n21820) );
  XNOR U3530 ( .A(n22926), .B(n22555), .Z(n22557) );
  XNOR U3531 ( .A(n22920), .B(n22934), .Z(n22924) );
  XOR U3532 ( .A(n2802), .B(n2801), .Z(n2442) );
  NANDN U3533 ( .A(n2063), .B(n2064), .Z(n1691) );
  NANDN U3534 ( .A(n3553), .B(n3554), .Z(n3181) );
  NAND U3535 ( .A(n5041), .B(n5042), .Z(n4669) );
  AND U3536 ( .A(n6530), .B(n6531), .Z(n6158) );
  ANDN U3537 ( .B(n8018), .A(n8019), .Z(n7646) );
  ANDN U3538 ( .B(n9506), .A(n9507), .Z(n9134) );
  AND U3539 ( .A(n5), .B(n6), .Z(n3) );
  AND U3540 ( .A(n13), .B(n14), .Z(n11) );
  AND U3541 ( .A(n21), .B(n22), .Z(n19) );
  AND U3542 ( .A(n29), .B(n30), .Z(n27) );
  AND U3543 ( .A(n37), .B(n38), .Z(n35) );
  AND U3544 ( .A(n45), .B(n46), .Z(n43) );
  AND U3545 ( .A(n53), .B(n54), .Z(n51) );
  AND U3546 ( .A(n61), .B(n62), .Z(n59) );
  AND U3547 ( .A(n69), .B(n70), .Z(n67) );
  XNOR U3548 ( .A(n11963), .B(n12320), .Z(n11972) );
  XNOR U3549 ( .A(n12699), .B(n13056), .Z(n12704) );
  XNOR U3550 ( .A(n16379), .B(n16736), .Z(n16384) );
  XNOR U3551 ( .A(n17115), .B(n17472), .Z(n17120) );
  XNOR U3552 ( .A(n20795), .B(n21152), .Z(n20800) );
  XNOR U3553 ( .A(n21531), .B(n21888), .Z(n21536) );
  XNOR U3554 ( .A(n13441), .B(n13791), .Z(n13445) );
  XNOR U3555 ( .A(n14177), .B(n14527), .Z(n14181) );
  XNOR U3556 ( .A(n17857), .B(n18207), .Z(n17861) );
  XNOR U3557 ( .A(n18593), .B(n18943), .Z(n18597) );
  XNOR U3558 ( .A(n22273), .B(n22623), .Z(n22277) );
  XNOR U3559 ( .A(n24565), .B(n24915), .Z(n24569) );
  XNOR U3560 ( .A(n23830), .B(n24180), .Z(n23834) );
  XNOR U3561 ( .A(n8483), .B(n8831), .Z(n8487) );
  XNOR U3562 ( .A(n9223), .B(n9574), .Z(n9227) );
  XNOR U3563 ( .A(n9975), .B(n10472), .Z(n9979) );
  XNOR U3564 ( .A(n10500), .B(n10843), .Z(n10504) );
  XNOR U3565 ( .A(n10868), .B(n11212), .Z(n10872) );
  XNOR U3566 ( .A(n11237), .B(n11581), .Z(n11241) );
  XNOR U3567 ( .A(n11979), .B(n11608), .Z(n11610) );
  XNOR U3568 ( .A(n12347), .B(n11976), .Z(n11978) );
  XNOR U3569 ( .A(n14918), .B(n15262), .Z(n14922) );
  XNOR U3570 ( .A(n15654), .B(n15998), .Z(n15658) );
  XNOR U3571 ( .A(n19334), .B(n19678), .Z(n19338) );
  XNOR U3572 ( .A(n20070), .B(n20414), .Z(n20074) );
  XNOR U3573 ( .A(n23014), .B(n23358), .Z(n23018) );
  XNOR U3574 ( .A(n8116), .B(n8458), .Z(n8120) );
  XNOR U3575 ( .A(n12719), .B(n13053), .Z(n12714) );
  XNOR U3576 ( .A(n16395), .B(n16733), .Z(n16399) );
  XNOR U3577 ( .A(n17131), .B(n17469), .Z(n17135) );
  XNOR U3578 ( .A(n20811), .B(n21149), .Z(n20815) );
  XNOR U3579 ( .A(n21547), .B(n21885), .Z(n21551) );
  XNOR U3580 ( .A(n13456), .B(n13788), .Z(n13464) );
  XNOR U3581 ( .A(n14192), .B(n14524), .Z(n14196) );
  XNOR U3582 ( .A(n17872), .B(n18204), .Z(n17876) );
  XNOR U3583 ( .A(n18608), .B(n18940), .Z(n18612) );
  XNOR U3584 ( .A(n22288), .B(n22620), .Z(n22292) );
  XNOR U3585 ( .A(n25972), .B(n26304), .Z(n25976) );
  XNOR U3586 ( .A(n25288), .B(n25620), .Z(n25292) );
  XNOR U3587 ( .A(n24580), .B(n24912), .Z(n24584) );
  XNOR U3588 ( .A(n23845), .B(n24177), .Z(n23849) );
  XNOR U3589 ( .A(n7367), .B(n7715), .Z(n7371) );
  XNOR U3590 ( .A(n9238), .B(n9571), .Z(n9242) );
  XNOR U3591 ( .A(n9990), .B(n10466), .Z(n9994) );
  XNOR U3592 ( .A(n10515), .B(n10840), .Z(n10519) );
  XNOR U3593 ( .A(n10883), .B(n11209), .Z(n10887) );
  XNOR U3594 ( .A(n11252), .B(n11578), .Z(n11256) );
  XNOR U3595 ( .A(n11994), .B(n11623), .Z(n11625) );
  XNOR U3596 ( .A(n12362), .B(n11991), .Z(n11993) );
  XNOR U3597 ( .A(n12730), .B(n12359), .Z(n12361) );
  XNOR U3598 ( .A(n13098), .B(n12727), .Z(n12729) );
  XNOR U3599 ( .A(n13466), .B(n13095), .Z(n13097) );
  XNOR U3600 ( .A(n14933), .B(n15259), .Z(n14937) );
  XNOR U3601 ( .A(n15669), .B(n15995), .Z(n15673) );
  XNOR U3602 ( .A(n19349), .B(n19675), .Z(n19353) );
  XNOR U3603 ( .A(n20085), .B(n20411), .Z(n20089) );
  XNOR U3604 ( .A(n23029), .B(n23355), .Z(n23033) );
  XNOR U3605 ( .A(n8131), .B(n8455), .Z(n8135) );
  XNOR U3606 ( .A(n8875), .B(n9195), .Z(n8879) );
  XNOR U3607 ( .A(n16410), .B(n16730), .Z(n16414) );
  XNOR U3608 ( .A(n17146), .B(n17466), .Z(n17150) );
  XNOR U3609 ( .A(n20826), .B(n21146), .Z(n20830) );
  XNOR U3610 ( .A(n21562), .B(n21882), .Z(n21566) );
  XNOR U3611 ( .A(n14211), .B(n14521), .Z(n14206) );
  XNOR U3612 ( .A(n17887), .B(n18201), .Z(n17891) );
  XNOR U3613 ( .A(n18623), .B(n18937), .Z(n18627) );
  XNOR U3614 ( .A(n22303), .B(n22617), .Z(n22307) );
  XNOR U3615 ( .A(n26647), .B(n26961), .Z(n26651) );
  XNOR U3616 ( .A(n25987), .B(n26301), .Z(n25991) );
  XNOR U3617 ( .A(n25303), .B(n25617), .Z(n25307) );
  XNOR U3618 ( .A(n24595), .B(n24909), .Z(n24599) );
  XNOR U3619 ( .A(n23860), .B(n24174), .Z(n23864) );
  XNOR U3620 ( .A(n6997), .B(n7342), .Z(n7001) );
  XNOR U3621 ( .A(n10005), .B(n10460), .Z(n10009) );
  XNOR U3622 ( .A(n10530), .B(n10837), .Z(n10534) );
  XNOR U3623 ( .A(n10898), .B(n11206), .Z(n10902) );
  XNOR U3624 ( .A(n11267), .B(n11575), .Z(n11271) );
  XNOR U3625 ( .A(n12009), .B(n11638), .Z(n11640) );
  XNOR U3626 ( .A(n12377), .B(n12006), .Z(n12008) );
  XNOR U3627 ( .A(n12745), .B(n12374), .Z(n12376) );
  XNOR U3628 ( .A(n13113), .B(n12742), .Z(n12744) );
  XNOR U3629 ( .A(n13481), .B(n13110), .Z(n13112) );
  XNOR U3630 ( .A(n13849), .B(n13478), .Z(n13480) );
  XNOR U3631 ( .A(n14217), .B(n13846), .Z(n13848) );
  XNOR U3632 ( .A(n14585), .B(n14214), .Z(n14216) );
  XNOR U3633 ( .A(n14948), .B(n15256), .Z(n14956) );
  XNOR U3634 ( .A(n15684), .B(n15992), .Z(n15688) );
  XNOR U3635 ( .A(n19364), .B(n19672), .Z(n19368) );
  XNOR U3636 ( .A(n20100), .B(n20408), .Z(n20104) );
  XNOR U3637 ( .A(n23044), .B(n23352), .Z(n23048) );
  XNOR U3638 ( .A(n7387), .B(n7711), .Z(n7391) );
  XNOR U3639 ( .A(n8146), .B(n8452), .Z(n8150) );
  XNOR U3640 ( .A(n8890), .B(n9192), .Z(n8894) );
  XNOR U3641 ( .A(n9633), .B(n9944), .Z(n9637) );
  XNOR U3642 ( .A(n16425), .B(n16727), .Z(n16429) );
  XNOR U3643 ( .A(n17161), .B(n17463), .Z(n17165) );
  XNOR U3644 ( .A(n20841), .B(n21143), .Z(n20845) );
  XNOR U3645 ( .A(n21577), .B(n21879), .Z(n21581) );
  XNOR U3646 ( .A(n17902), .B(n18198), .Z(n17906) );
  XNOR U3647 ( .A(n18638), .B(n18934), .Z(n18642) );
  XNOR U3648 ( .A(n22318), .B(n22614), .Z(n22322) );
  XNOR U3649 ( .A(n27910), .B(n28206), .Z(n27914) );
  XNOR U3650 ( .A(n27298), .B(n27594), .Z(n27302) );
  XNOR U3651 ( .A(n26662), .B(n26958), .Z(n26666) );
  XNOR U3652 ( .A(n26002), .B(n26298), .Z(n26006) );
  XNOR U3653 ( .A(n25318), .B(n25614), .Z(n25322) );
  XNOR U3654 ( .A(n24610), .B(n24906), .Z(n24614) );
  XNOR U3655 ( .A(n23875), .B(n24171), .Z(n23879) );
  XNOR U3656 ( .A(n6252), .B(n6600), .Z(n6256) );
  XNOR U3657 ( .A(n10545), .B(n10834), .Z(n10549) );
  XNOR U3658 ( .A(n10913), .B(n11203), .Z(n10917) );
  XNOR U3659 ( .A(n11282), .B(n11572), .Z(n11286) );
  XNOR U3660 ( .A(n12024), .B(n11653), .Z(n11655) );
  XNOR U3661 ( .A(n12392), .B(n12021), .Z(n12023) );
  XNOR U3662 ( .A(n12760), .B(n12389), .Z(n12391) );
  XNOR U3663 ( .A(n13128), .B(n12757), .Z(n12759) );
  XNOR U3664 ( .A(n13496), .B(n13125), .Z(n13127) );
  XNOR U3665 ( .A(n13864), .B(n13493), .Z(n13495) );
  XNOR U3666 ( .A(n14232), .B(n13861), .Z(n13863) );
  XNOR U3667 ( .A(n14600), .B(n14229), .Z(n14231) );
  XNOR U3668 ( .A(n14968), .B(n14597), .Z(n14599) );
  XNOR U3669 ( .A(n15336), .B(n14965), .Z(n14967) );
  XNOR U3670 ( .A(n15704), .B(n15333), .Z(n15335) );
  XNOR U3671 ( .A(n15703), .B(n15989), .Z(n15698) );
  XNOR U3672 ( .A(n19379), .B(n19669), .Z(n19383) );
  XNOR U3673 ( .A(n20115), .B(n20405), .Z(n20119) );
  XNOR U3674 ( .A(n23059), .B(n23349), .Z(n23063) );
  XNOR U3675 ( .A(n7402), .B(n7708), .Z(n7406) );
  XNOR U3676 ( .A(n8905), .B(n9189), .Z(n8909) );
  XNOR U3677 ( .A(n9648), .B(n9941), .Z(n9652) );
  XNOR U3678 ( .A(n16440), .B(n16724), .Z(n16448) );
  XNOR U3679 ( .A(n17176), .B(n17460), .Z(n17180) );
  XNOR U3680 ( .A(n20856), .B(n21140), .Z(n20860) );
  XNOR U3681 ( .A(n21592), .B(n21876), .Z(n21596) );
  XNOR U3682 ( .A(n6644), .B(n6964), .Z(n6648) );
  XNOR U3683 ( .A(n17917), .B(n18195), .Z(n17921) );
  XNOR U3684 ( .A(n18653), .B(n18931), .Z(n18657) );
  XNOR U3685 ( .A(n22333), .B(n22611), .Z(n22337) );
  XNOR U3686 ( .A(n28513), .B(n28791), .Z(n28517) );
  XNOR U3687 ( .A(n27925), .B(n28203), .Z(n27929) );
  XNOR U3688 ( .A(n27313), .B(n27591), .Z(n27317) );
  XNOR U3689 ( .A(n26677), .B(n26955), .Z(n26681) );
  XNOR U3690 ( .A(n26017), .B(n26295), .Z(n26021) );
  XNOR U3691 ( .A(n25333), .B(n25611), .Z(n25337) );
  XNOR U3692 ( .A(n24625), .B(n24903), .Z(n24629) );
  XNOR U3693 ( .A(n23890), .B(n24168), .Z(n23894) );
  XNOR U3694 ( .A(n5503), .B(n5857), .Z(n5507) );
  XNOR U3695 ( .A(n8171), .B(n8447), .Z(n8175) );
  XNOR U3696 ( .A(n10934), .B(n10563), .Z(n10565) );
  XNOR U3697 ( .A(n10928), .B(n11200), .Z(n10932) );
  XNOR U3698 ( .A(n11297), .B(n11569), .Z(n11301) );
  XNOR U3699 ( .A(n12039), .B(n11668), .Z(n11670) );
  XNOR U3700 ( .A(n12407), .B(n12036), .Z(n12038) );
  XNOR U3701 ( .A(n12775), .B(n12404), .Z(n12406) );
  XNOR U3702 ( .A(n13143), .B(n12772), .Z(n12774) );
  XNOR U3703 ( .A(n13511), .B(n13140), .Z(n13142) );
  XNOR U3704 ( .A(n13879), .B(n13508), .Z(n13510) );
  XNOR U3705 ( .A(n14247), .B(n13876), .Z(n13878) );
  XNOR U3706 ( .A(n14615), .B(n14244), .Z(n14246) );
  XNOR U3707 ( .A(n14983), .B(n14612), .Z(n14614) );
  XNOR U3708 ( .A(n15351), .B(n14980), .Z(n14982) );
  XNOR U3709 ( .A(n15719), .B(n15348), .Z(n15350) );
  XNOR U3710 ( .A(n16087), .B(n15716), .Z(n15718) );
  XNOR U3711 ( .A(n16455), .B(n16084), .Z(n16086) );
  XNOR U3712 ( .A(n16823), .B(n16452), .Z(n16454) );
  XNOR U3713 ( .A(n19394), .B(n19666), .Z(n19398) );
  XNOR U3714 ( .A(n20130), .B(n20402), .Z(n20134) );
  XNOR U3715 ( .A(n23074), .B(n23346), .Z(n23078) );
  XNOR U3716 ( .A(n8920), .B(n9186), .Z(n8924) );
  XNOR U3717 ( .A(n9663), .B(n9938), .Z(n9667) );
  XNOR U3718 ( .A(n17195), .B(n17457), .Z(n17190) );
  XNOR U3719 ( .A(n20871), .B(n21137), .Z(n20875) );
  XNOR U3720 ( .A(n21607), .B(n21873), .Z(n21611) );
  XNOR U3721 ( .A(n6659), .B(n6961), .Z(n6663) );
  XNOR U3722 ( .A(n5895), .B(n6225), .Z(n5899) );
  XNOR U3723 ( .A(n17932), .B(n18192), .Z(n17940) );
  XNOR U3724 ( .A(n18668), .B(n18928), .Z(n18672) );
  XNOR U3725 ( .A(n22348), .B(n22608), .Z(n22352) );
  XNOR U3726 ( .A(n29632), .B(n29892), .Z(n29636) );
  XNOR U3727 ( .A(n29092), .B(n29352), .Z(n29096) );
  XNOR U3728 ( .A(n28528), .B(n28788), .Z(n28532) );
  XNOR U3729 ( .A(n27940), .B(n28200), .Z(n27944) );
  XNOR U3730 ( .A(n27328), .B(n27588), .Z(n27332) );
  XNOR U3731 ( .A(n26692), .B(n26952), .Z(n26696) );
  XNOR U3732 ( .A(n26032), .B(n26292), .Z(n26036) );
  XNOR U3733 ( .A(n25348), .B(n25608), .Z(n25352) );
  XNOR U3734 ( .A(n24640), .B(n24900), .Z(n24644) );
  XNOR U3735 ( .A(n23905), .B(n24165), .Z(n23909) );
  XNOR U3736 ( .A(n7042), .B(n7333), .Z(n7046) );
  XNOR U3737 ( .A(n5136), .B(n5484), .Z(n5140) );
  XNOR U3738 ( .A(n8186), .B(n8444), .Z(n8190) );
  XNOR U3739 ( .A(n11318), .B(n10946), .Z(n10948) );
  XNOR U3740 ( .A(n11312), .B(n11566), .Z(n11316) );
  XNOR U3741 ( .A(n12054), .B(n11683), .Z(n11685) );
  XNOR U3742 ( .A(n12422), .B(n12051), .Z(n12053) );
  XNOR U3743 ( .A(n12790), .B(n12419), .Z(n12421) );
  XNOR U3744 ( .A(n13158), .B(n12787), .Z(n12789) );
  XNOR U3745 ( .A(n13526), .B(n13155), .Z(n13157) );
  XNOR U3746 ( .A(n13894), .B(n13523), .Z(n13525) );
  XNOR U3747 ( .A(n14262), .B(n13891), .Z(n13893) );
  XNOR U3748 ( .A(n14630), .B(n14259), .Z(n14261) );
  XNOR U3749 ( .A(n14998), .B(n14627), .Z(n14629) );
  XNOR U3750 ( .A(n15366), .B(n14995), .Z(n14997) );
  XNOR U3751 ( .A(n15734), .B(n15363), .Z(n15365) );
  XNOR U3752 ( .A(n16102), .B(n15731), .Z(n15733) );
  XNOR U3753 ( .A(n16470), .B(n16099), .Z(n16101) );
  XNOR U3754 ( .A(n16838), .B(n16467), .Z(n16469) );
  XNOR U3755 ( .A(n17206), .B(n16835), .Z(n16837) );
  XNOR U3756 ( .A(n17574), .B(n17203), .Z(n17205) );
  XNOR U3757 ( .A(n17942), .B(n17571), .Z(n17573) );
  XNOR U3758 ( .A(n19409), .B(n19663), .Z(n19413) );
  XNOR U3759 ( .A(n20145), .B(n20399), .Z(n20149) );
  XNOR U3760 ( .A(n23089), .B(n23343), .Z(n23093) );
  XNOR U3761 ( .A(n8935), .B(n9183), .Z(n8939) );
  XNOR U3762 ( .A(n9678), .B(n9935), .Z(n9682) );
  XNOR U3763 ( .A(n11323), .B(n10951), .Z(n10953) );
  XNOR U3764 ( .A(n20886), .B(n21134), .Z(n20890) );
  XNOR U3765 ( .A(n21622), .B(n21870), .Z(n21626) );
  XNOR U3766 ( .A(n5528), .B(n5852), .Z(n5532) );
  XNOR U3767 ( .A(n10585), .B(n10826), .Z(n10589) );
  XNOR U3768 ( .A(n18687), .B(n18925), .Z(n18682) );
  XNOR U3769 ( .A(n22363), .B(n22605), .Z(n22367) );
  XNOR U3770 ( .A(n30163), .B(n30405), .Z(n30167) );
  XNOR U3771 ( .A(n29647), .B(n29889), .Z(n29651) );
  XNOR U3772 ( .A(n29107), .B(n29349), .Z(n29111) );
  XNOR U3773 ( .A(n28543), .B(n28785), .Z(n28547) );
  XNOR U3774 ( .A(n27955), .B(n28197), .Z(n27959) );
  XNOR U3775 ( .A(n27343), .B(n27585), .Z(n27347) );
  XNOR U3776 ( .A(n26707), .B(n26949), .Z(n26711) );
  XNOR U3777 ( .A(n26047), .B(n26289), .Z(n26051) );
  XNOR U3778 ( .A(n25363), .B(n25605), .Z(n25367) );
  XNOR U3779 ( .A(n24655), .B(n24897), .Z(n24659) );
  XNOR U3780 ( .A(n23920), .B(n24162), .Z(n23924) );
  XNOR U3781 ( .A(n7057), .B(n7330), .Z(n7061) );
  XNOR U3782 ( .A(n5915), .B(n6221), .Z(n5919) );
  XNOR U3783 ( .A(n4768), .B(n5111), .Z(n4772) );
  XNOR U3784 ( .A(n8201), .B(n8441), .Z(n8205) );
  XNOR U3785 ( .A(n12437), .B(n12066), .Z(n12068) );
  XNOR U3786 ( .A(n12805), .B(n12434), .Z(n12436) );
  XNOR U3787 ( .A(n13173), .B(n12802), .Z(n12804) );
  XNOR U3788 ( .A(n13541), .B(n13170), .Z(n13172) );
  XNOR U3789 ( .A(n13909), .B(n13538), .Z(n13540) );
  XNOR U3790 ( .A(n14277), .B(n13906), .Z(n13908) );
  XNOR U3791 ( .A(n14645), .B(n14274), .Z(n14276) );
  XNOR U3792 ( .A(n15013), .B(n14642), .Z(n14644) );
  XNOR U3793 ( .A(n15381), .B(n15010), .Z(n15012) );
  XNOR U3794 ( .A(n15749), .B(n15378), .Z(n15380) );
  XNOR U3795 ( .A(n16117), .B(n15746), .Z(n15748) );
  XNOR U3796 ( .A(n16485), .B(n16114), .Z(n16116) );
  XNOR U3797 ( .A(n16853), .B(n16482), .Z(n16484) );
  XNOR U3798 ( .A(n17221), .B(n16850), .Z(n16852) );
  XNOR U3799 ( .A(n17589), .B(n17218), .Z(n17220) );
  XNOR U3800 ( .A(n17957), .B(n17586), .Z(n17588) );
  XNOR U3801 ( .A(n18325), .B(n17954), .Z(n17956) );
  XNOR U3802 ( .A(n18693), .B(n18322), .Z(n18324) );
  XNOR U3803 ( .A(n19061), .B(n18690), .Z(n18692) );
  XNOR U3804 ( .A(n19424), .B(n19660), .Z(n19432) );
  XNOR U3805 ( .A(n20160), .B(n20396), .Z(n20164) );
  XNOR U3806 ( .A(n23104), .B(n23340), .Z(n23108) );
  XNOR U3807 ( .A(n6302), .B(n6590), .Z(n6306) );
  XNOR U3808 ( .A(n4008), .B(n4369), .Z(n4013) );
  XNOR U3809 ( .A(n9318), .B(n9555), .Z(n9322) );
  XNOR U3810 ( .A(n10070), .B(n10434), .Z(n10074) );
  XNOR U3811 ( .A(n11700), .B(n11930), .Z(n11704) );
  XNOR U3812 ( .A(n20901), .B(n21131), .Z(n20905) );
  XNOR U3813 ( .A(n21637), .B(n21867), .Z(n21641) );
  XNOR U3814 ( .A(n10968), .B(n11192), .Z(n10972) );
  XNOR U3815 ( .A(n11337), .B(n11561), .Z(n11341) );
  XNOR U3816 ( .A(n22378), .B(n22602), .Z(n22382) );
  XNOR U3817 ( .A(n31138), .B(n31362), .Z(n31142) );
  XNOR U3818 ( .A(n30670), .B(n30894), .Z(n30674) );
  XNOR U3819 ( .A(n30178), .B(n30402), .Z(n30182) );
  XNOR U3820 ( .A(n29662), .B(n29886), .Z(n29666) );
  XNOR U3821 ( .A(n29122), .B(n29346), .Z(n29126) );
  XNOR U3822 ( .A(n28558), .B(n28782), .Z(n28562) );
  XNOR U3823 ( .A(n27970), .B(n28194), .Z(n27974) );
  XNOR U3824 ( .A(n27358), .B(n27582), .Z(n27362) );
  XNOR U3825 ( .A(n26722), .B(n26946), .Z(n26726) );
  XNOR U3826 ( .A(n26062), .B(n26286), .Z(n26066) );
  XNOR U3827 ( .A(n25378), .B(n25602), .Z(n25382) );
  XNOR U3828 ( .A(n24670), .B(n24894), .Z(n24674) );
  XNOR U3829 ( .A(n23935), .B(n24159), .Z(n23939) );
  XNOR U3830 ( .A(n7072), .B(n7327), .Z(n7076) );
  XNOR U3831 ( .A(n5166), .B(n5478), .Z(n5170) );
  XNOR U3832 ( .A(n8216), .B(n8438), .Z(n8220) );
  XNOR U3833 ( .A(n8960), .B(n9178), .Z(n8964) );
  XNOR U3834 ( .A(n12078), .B(n12296), .Z(n12082) );
  XNOR U3835 ( .A(n13556), .B(n13185), .Z(n13187) );
  XNOR U3836 ( .A(n13924), .B(n13553), .Z(n13555) );
  XNOR U3837 ( .A(n14292), .B(n13921), .Z(n13923) );
  XNOR U3838 ( .A(n14660), .B(n14289), .Z(n14291) );
  XNOR U3839 ( .A(n15028), .B(n14657), .Z(n14659) );
  XNOR U3840 ( .A(n15396), .B(n15025), .Z(n15027) );
  XNOR U3841 ( .A(n15764), .B(n15393), .Z(n15395) );
  XNOR U3842 ( .A(n16132), .B(n15761), .Z(n15763) );
  XNOR U3843 ( .A(n16500), .B(n16129), .Z(n16131) );
  XNOR U3844 ( .A(n16868), .B(n16497), .Z(n16499) );
  XNOR U3845 ( .A(n17236), .B(n16865), .Z(n16867) );
  XNOR U3846 ( .A(n17604), .B(n17233), .Z(n17235) );
  XNOR U3847 ( .A(n17972), .B(n17601), .Z(n17603) );
  XNOR U3848 ( .A(n18340), .B(n17969), .Z(n17971) );
  XNOR U3849 ( .A(n18708), .B(n18337), .Z(n18339) );
  XNOR U3850 ( .A(n19076), .B(n18705), .Z(n18707) );
  XNOR U3851 ( .A(n19444), .B(n19073), .Z(n19075) );
  XNOR U3852 ( .A(n19812), .B(n19441), .Z(n19443) );
  XNOR U3853 ( .A(n20180), .B(n19809), .Z(n19811) );
  XNOR U3854 ( .A(n20179), .B(n20393), .Z(n20174) );
  XNOR U3855 ( .A(n23119), .B(n23337), .Z(n23123) );
  XNOR U3856 ( .A(n6317), .B(n6587), .Z(n6321) );
  XNOR U3857 ( .A(n4406), .B(n4736), .Z(n4410) );
  XNOR U3858 ( .A(n3642), .B(n3996), .Z(n3646) );
  XNOR U3859 ( .A(n10085), .B(n10428), .Z(n10089) );
  XNOR U3860 ( .A(n10610), .B(n10821), .Z(n10614) );
  XNOR U3861 ( .A(n11353), .B(n10981), .Z(n10983) );
  XNOR U3862 ( .A(n12819), .B(n13031), .Z(n12823) );
  XNOR U3863 ( .A(n20916), .B(n21128), .Z(n20924) );
  XNOR U3864 ( .A(n21652), .B(n21864), .Z(n21656) );
  XNOR U3865 ( .A(n5558), .B(n5846), .Z(n5562) );
  XNOR U3866 ( .A(n11720), .B(n11926), .Z(n11724) );
  XNOR U3867 ( .A(n12830), .B(n12459), .Z(n12461) );
  XNOR U3868 ( .A(n22393), .B(n22599), .Z(n22397) );
  XNOR U3869 ( .A(n31597), .B(n31974), .Z(n31601) );
  XNOR U3870 ( .A(n31153), .B(n31359), .Z(n31157) );
  XNOR U3871 ( .A(n30685), .B(n30891), .Z(n30689) );
  XNOR U3872 ( .A(n30193), .B(n30399), .Z(n30197) );
  XNOR U3873 ( .A(n29677), .B(n29883), .Z(n29681) );
  XNOR U3874 ( .A(n29137), .B(n29343), .Z(n29141) );
  XNOR U3875 ( .A(n28573), .B(n28779), .Z(n28577) );
  XNOR U3876 ( .A(n27985), .B(n28191), .Z(n27989) );
  XNOR U3877 ( .A(n27373), .B(n27579), .Z(n27377) );
  XNOR U3878 ( .A(n26737), .B(n26943), .Z(n26741) );
  XNOR U3879 ( .A(n26077), .B(n26283), .Z(n26081) );
  XNOR U3880 ( .A(n25393), .B(n25599), .Z(n25397) );
  XNOR U3881 ( .A(n24685), .B(n24891), .Z(n24689) );
  XNOR U3882 ( .A(n23950), .B(n24156), .Z(n23954) );
  XNOR U3883 ( .A(n7476), .B(n7694), .Z(n7471) );
  XNOR U3884 ( .A(n6709), .B(n6951), .Z(n6713) );
  XNOR U3885 ( .A(n4798), .B(n5105), .Z(n4802) );
  XNOR U3886 ( .A(n8233), .B(n8434), .Z(n8234) );
  XNOR U3887 ( .A(n8975), .B(n9175), .Z(n8983) );
  XNOR U3888 ( .A(n9718), .B(n9927), .Z(n9722) );
  XNOR U3889 ( .A(n13197), .B(n13397), .Z(n13201) );
  XNOR U3890 ( .A(n14675), .B(n14304), .Z(n14306) );
  XNOR U3891 ( .A(n15043), .B(n14672), .Z(n14674) );
  XNOR U3892 ( .A(n15411), .B(n15040), .Z(n15042) );
  XNOR U3893 ( .A(n15779), .B(n15408), .Z(n15410) );
  XNOR U3894 ( .A(n16147), .B(n15776), .Z(n15778) );
  XNOR U3895 ( .A(n16515), .B(n16144), .Z(n16146) );
  XNOR U3896 ( .A(n16883), .B(n16512), .Z(n16514) );
  XNOR U3897 ( .A(n17251), .B(n16880), .Z(n16882) );
  XNOR U3898 ( .A(n17619), .B(n17248), .Z(n17250) );
  XNOR U3899 ( .A(n17987), .B(n17616), .Z(n17618) );
  XNOR U3900 ( .A(n18355), .B(n17984), .Z(n17986) );
  XNOR U3901 ( .A(n18723), .B(n18352), .Z(n18354) );
  XNOR U3902 ( .A(n19091), .B(n18720), .Z(n18722) );
  XNOR U3903 ( .A(n19459), .B(n19088), .Z(n19090) );
  XNOR U3904 ( .A(n19827), .B(n19456), .Z(n19458) );
  XNOR U3905 ( .A(n20195), .B(n19824), .Z(n19826) );
  XNOR U3906 ( .A(n20563), .B(n20192), .Z(n20194) );
  XNOR U3907 ( .A(n20931), .B(n20560), .Z(n20562) );
  XNOR U3908 ( .A(n21299), .B(n20928), .Z(n20930) );
  XNOR U3909 ( .A(n23134), .B(n23334), .Z(n23138) );
  XNOR U3910 ( .A(n6733), .B(n6945), .Z(n6737) );
  XNOR U3911 ( .A(n5950), .B(n6214), .Z(n5954) );
  XNOR U3912 ( .A(n4039), .B(n4363), .Z(n4043) );
  XNOR U3913 ( .A(n3275), .B(n3623), .Z(n3279) );
  XNOR U3914 ( .A(n11368), .B(n10996), .Z(n10998) );
  XNOR U3915 ( .A(n11362), .B(n11556), .Z(n11366) );
  XNOR U3916 ( .A(n12104), .B(n11733), .Z(n11735) );
  XNOR U3917 ( .A(n12098), .B(n12292), .Z(n12102) );
  XNOR U3918 ( .A(n13938), .B(n14132), .Z(n13942) );
  XNOR U3919 ( .A(n21671), .B(n21861), .Z(n21666) );
  XNOR U3920 ( .A(n5191), .B(n5473), .Z(n5195) );
  XNOR U3921 ( .A(n6001), .B(n6202), .Z(n6002) );
  XNOR U3922 ( .A(n12839), .B(n13027), .Z(n12843) );
  XNOR U3923 ( .A(n13949), .B(n13578), .Z(n13580) );
  XNOR U3924 ( .A(n22408), .B(n22596), .Z(n22416) );
  XNOR U3925 ( .A(n32578), .B(n32758), .Z(n32582) );
  XNOR U3926 ( .A(n32195), .B(n32375), .Z(n32199) );
  XNOR U3927 ( .A(n31612), .B(n31971), .Z(n31616) );
  XNOR U3928 ( .A(n31168), .B(n31356), .Z(n31172) );
  XNOR U3929 ( .A(n30700), .B(n30888), .Z(n30704) );
  XNOR U3930 ( .A(n30208), .B(n30396), .Z(n30212) );
  XNOR U3931 ( .A(n29692), .B(n29880), .Z(n29696) );
  XNOR U3932 ( .A(n29152), .B(n29340), .Z(n29156) );
  XNOR U3933 ( .A(n28588), .B(n28776), .Z(n28592) );
  XNOR U3934 ( .A(n28000), .B(n28188), .Z(n28004) );
  XNOR U3935 ( .A(n27388), .B(n27576), .Z(n27392) );
  XNOR U3936 ( .A(n26752), .B(n26940), .Z(n26756) );
  XNOR U3937 ( .A(n26092), .B(n26280), .Z(n26096) );
  XNOR U3938 ( .A(n25408), .B(n25596), .Z(n25412) );
  XNOR U3939 ( .A(n24700), .B(n24888), .Z(n24704) );
  XNOR U3940 ( .A(n23965), .B(n24153), .Z(n23969) );
  XNOR U3941 ( .A(n6346), .B(n6582), .Z(n6341) );
  XNOR U3942 ( .A(n4431), .B(n4731), .Z(n4435) );
  XNOR U3943 ( .A(n6757), .B(n6939), .Z(n6761) );
  XNOR U3944 ( .A(n7505), .B(n7687), .Z(n7500) );
  XNOR U3945 ( .A(n8245), .B(n8431), .Z(n8249) );
  XNOR U3946 ( .A(n8989), .B(n9171), .Z(n8993) );
  XNOR U3947 ( .A(n9737), .B(n9924), .Z(n9731) );
  XNOR U3948 ( .A(n10635), .B(n10816), .Z(n10639) );
  XNOR U3949 ( .A(n14316), .B(n14498), .Z(n14320) );
  XNOR U3950 ( .A(n15794), .B(n15423), .Z(n15425) );
  XNOR U3951 ( .A(n16162), .B(n15791), .Z(n15793) );
  XNOR U3952 ( .A(n16530), .B(n16159), .Z(n16161) );
  XNOR U3953 ( .A(n16898), .B(n16527), .Z(n16529) );
  XNOR U3954 ( .A(n17266), .B(n16895), .Z(n16897) );
  XNOR U3955 ( .A(n17634), .B(n17263), .Z(n17265) );
  XNOR U3956 ( .A(n18002), .B(n17631), .Z(n17633) );
  XNOR U3957 ( .A(n18370), .B(n17999), .Z(n18001) );
  XNOR U3958 ( .A(n18738), .B(n18367), .Z(n18369) );
  XNOR U3959 ( .A(n19106), .B(n18735), .Z(n18737) );
  XNOR U3960 ( .A(n19474), .B(n19103), .Z(n19105) );
  XNOR U3961 ( .A(n19842), .B(n19471), .Z(n19473) );
  XNOR U3962 ( .A(n20210), .B(n19839), .Z(n19841) );
  XNOR U3963 ( .A(n20578), .B(n20207), .Z(n20209) );
  XNOR U3964 ( .A(n20946), .B(n20575), .Z(n20577) );
  XNOR U3965 ( .A(n21314), .B(n20943), .Z(n20945) );
  XNOR U3966 ( .A(n21682), .B(n21311), .Z(n21313) );
  XNOR U3967 ( .A(n22050), .B(n21679), .Z(n21681) );
  XNOR U3968 ( .A(n22418), .B(n22047), .Z(n22049) );
  XNOR U3969 ( .A(n23149), .B(n23331), .Z(n23153) );
  XNOR U3970 ( .A(n6366), .B(n6576), .Z(n6374) );
  XNOR U3971 ( .A(n5220), .B(n5466), .Z(n5224) );
  XNOR U3972 ( .A(n5583), .B(n5841), .Z(n5591) );
  XNOR U3973 ( .A(n2908), .B(n3250), .Z(n2912) );
  XNOR U3974 ( .A(n11377), .B(n11553), .Z(n11381) );
  XNOR U3975 ( .A(n12119), .B(n11748), .Z(n11750) );
  XNOR U3976 ( .A(n12113), .B(n12289), .Z(n12117) );
  XNOR U3977 ( .A(n12855), .B(n12484), .Z(n12486) );
  XNOR U3978 ( .A(n13223), .B(n12852), .Z(n12854) );
  XNOR U3979 ( .A(n13217), .B(n13393), .Z(n13221) );
  XNOR U3980 ( .A(n15057), .B(n15233), .Z(n15061) );
  XNOR U3981 ( .A(n5607), .B(n5835), .Z(n5611) );
  XNOR U3982 ( .A(n3295), .B(n3619), .Z(n3299) );
  XNOR U3983 ( .A(n2146), .B(n2508), .Z(n2151) );
  XNOR U3984 ( .A(n5631), .B(n5829), .Z(n5635) );
  XNOR U3985 ( .A(n13958), .B(n14128), .Z(n13962) );
  XNOR U3986 ( .A(n15068), .B(n14697), .Z(n14699) );
  XNOR U3987 ( .A(n32949), .B(n33114), .Z(n32953) );
  XNOR U3988 ( .A(n32593), .B(n32755), .Z(n32597) );
  XNOR U3989 ( .A(n32210), .B(n32372), .Z(n32214) );
  XNOR U3990 ( .A(n31627), .B(n31968), .Z(n31631) );
  XNOR U3991 ( .A(n31183), .B(n31353), .Z(n31187) );
  XNOR U3992 ( .A(n30715), .B(n30885), .Z(n30719) );
  XNOR U3993 ( .A(n30223), .B(n30393), .Z(n30227) );
  XNOR U3994 ( .A(n29707), .B(n29877), .Z(n29711) );
  XNOR U3995 ( .A(n29167), .B(n29337), .Z(n29171) );
  XNOR U3996 ( .A(n28603), .B(n28773), .Z(n28607) );
  XNOR U3997 ( .A(n28015), .B(n28185), .Z(n28019) );
  XNOR U3998 ( .A(n27403), .B(n27573), .Z(n27407) );
  XNOR U3999 ( .A(n26767), .B(n26937), .Z(n26771) );
  XNOR U4000 ( .A(n26107), .B(n26277), .Z(n26111) );
  XNOR U4001 ( .A(n25423), .B(n25593), .Z(n25427) );
  XNOR U4002 ( .A(n24715), .B(n24885), .Z(n24719) );
  XNOR U4003 ( .A(n23980), .B(n24150), .Z(n23984) );
  XNOR U4004 ( .A(n4446), .B(n4728), .Z(n4450) );
  XNOR U4005 ( .A(n3682), .B(n3988), .Z(n3686) );
  XNOR U4006 ( .A(n6030), .B(n6195), .Z(n6031) );
  XNOR U4007 ( .A(n6772), .B(n6936), .Z(n6780) );
  XNOR U4008 ( .A(n7515), .B(n7683), .Z(n7519) );
  XNOR U4009 ( .A(n8262), .B(n8427), .Z(n8263) );
  XNOR U4010 ( .A(n9004), .B(n9168), .Z(n9012) );
  XNOR U4011 ( .A(n9747), .B(n9919), .Z(n9751) );
  XNOR U4012 ( .A(n10650), .B(n10813), .Z(n10654) );
  XNOR U4013 ( .A(n12129), .B(n11758), .Z(n11760) );
  XNOR U4014 ( .A(n15435), .B(n15599), .Z(n15439) );
  XNOR U4015 ( .A(n16913), .B(n16542), .Z(n16544) );
  XNOR U4016 ( .A(n17281), .B(n16910), .Z(n16912) );
  XNOR U4017 ( .A(n17649), .B(n17278), .Z(n17280) );
  XNOR U4018 ( .A(n18017), .B(n17646), .Z(n17648) );
  XNOR U4019 ( .A(n18385), .B(n18014), .Z(n18016) );
  XNOR U4020 ( .A(n18753), .B(n18382), .Z(n18384) );
  XNOR U4021 ( .A(n19121), .B(n18750), .Z(n18752) );
  XNOR U4022 ( .A(n19489), .B(n19118), .Z(n19120) );
  XNOR U4023 ( .A(n19857), .B(n19486), .Z(n19488) );
  XNOR U4024 ( .A(n20225), .B(n19854), .Z(n19856) );
  XNOR U4025 ( .A(n20593), .B(n20222), .Z(n20224) );
  XNOR U4026 ( .A(n20961), .B(n20590), .Z(n20592) );
  XNOR U4027 ( .A(n21329), .B(n20958), .Z(n20960) );
  XNOR U4028 ( .A(n21697), .B(n21326), .Z(n21328) );
  XNOR U4029 ( .A(n22065), .B(n21694), .Z(n21696) );
  XNOR U4030 ( .A(n22433), .B(n22062), .Z(n22064) );
  XNOR U4031 ( .A(n22801), .B(n22430), .Z(n22432) );
  XNOR U4032 ( .A(n23169), .B(n22798), .Z(n22800) );
  XNOR U4033 ( .A(n23158), .B(n23327), .Z(n23167) );
  XNOR U4034 ( .A(n4470), .B(n4722), .Z(n4474) );
  XNOR U4035 ( .A(n4837), .B(n5098), .Z(n4832) );
  XNOR U4036 ( .A(n5660), .B(n5822), .Z(n5664) );
  XNOR U4037 ( .A(n11392), .B(n11550), .Z(n11396) );
  XNOR U4038 ( .A(n12134), .B(n11763), .Z(n11765) );
  XNOR U4039 ( .A(n12870), .B(n12499), .Z(n12501) );
  XNOR U4040 ( .A(n13238), .B(n12867), .Z(n12869) );
  XNOR U4041 ( .A(n13232), .B(n13390), .Z(n13236) );
  XNOR U4042 ( .A(n13974), .B(n13603), .Z(n13605) );
  XNOR U4043 ( .A(n14342), .B(n13971), .Z(n13973) );
  XNOR U4044 ( .A(n14336), .B(n14494), .Z(n14340) );
  XNOR U4045 ( .A(n16176), .B(n16334), .Z(n16180) );
  XNOR U4046 ( .A(n5244), .B(n5462), .Z(n5239) );
  XNOR U4047 ( .A(n2545), .B(n2876), .Z(n2549) );
  XNOR U4048 ( .A(n1780), .B(n2134), .Z(n1784) );
  XNOR U4049 ( .A(n4881), .B(n5086), .Z(n4885) );
  XNOR U4050 ( .A(n4117), .B(n4345), .Z(n4121) );
  XNOR U4051 ( .A(n15077), .B(n15229), .Z(n15081) );
  XNOR U4052 ( .A(n16187), .B(n15816), .Z(n15818) );
  XNOR U4053 ( .A(n33610), .B(n33754), .Z(n33614) );
  XNOR U4054 ( .A(n33299), .B(n33443), .Z(n33303) );
  XNOR U4055 ( .A(n32964), .B(n33111), .Z(n32968) );
  XNOR U4056 ( .A(n32608), .B(n32752), .Z(n32612) );
  XNOR U4057 ( .A(n32225), .B(n32369), .Z(n32229) );
  XNOR U4058 ( .A(n31642), .B(n31965), .Z(n31646) );
  XNOR U4059 ( .A(n31198), .B(n31350), .Z(n31202) );
  XNOR U4060 ( .A(n30730), .B(n30882), .Z(n30734) );
  XNOR U4061 ( .A(n30238), .B(n30390), .Z(n30242) );
  XNOR U4062 ( .A(n29722), .B(n29874), .Z(n29726) );
  XNOR U4063 ( .A(n29182), .B(n29334), .Z(n29186) );
  XNOR U4064 ( .A(n28618), .B(n28770), .Z(n28622) );
  XNOR U4065 ( .A(n28030), .B(n28182), .Z(n28034) );
  XNOR U4066 ( .A(n27418), .B(n27570), .Z(n27422) );
  XNOR U4067 ( .A(n26782), .B(n26934), .Z(n26786) );
  XNOR U4068 ( .A(n26122), .B(n26274), .Z(n26126) );
  XNOR U4069 ( .A(n25438), .B(n25590), .Z(n25442) );
  XNOR U4070 ( .A(n24730), .B(n24882), .Z(n24734) );
  XNOR U4071 ( .A(n23995), .B(n24147), .Z(n23999) );
  XNOR U4072 ( .A(n3315), .B(n3615), .Z(n3319) );
  XNOR U4073 ( .A(n5273), .B(n5455), .Z(n5268) );
  XNOR U4074 ( .A(n6786), .B(n6932), .Z(n6790) );
  XNOR U4075 ( .A(n7534), .B(n7680), .Z(n7529) );
  XNOR U4076 ( .A(n8274), .B(n8424), .Z(n8278) );
  XNOR U4077 ( .A(n9018), .B(n9164), .Z(n9022) );
  XNOR U4078 ( .A(n9766), .B(n9916), .Z(n9760) );
  XNOR U4079 ( .A(n10665), .B(n10810), .Z(n10669) );
  XNOR U4080 ( .A(n12144), .B(n11773), .Z(n11775) );
  XNOR U4081 ( .A(n13248), .B(n12877), .Z(n12879) );
  XNOR U4082 ( .A(n16554), .B(n16700), .Z(n16558) );
  XNOR U4083 ( .A(n18032), .B(n17661), .Z(n17663) );
  XNOR U4084 ( .A(n18400), .B(n18029), .Z(n18031) );
  XNOR U4085 ( .A(n18768), .B(n18397), .Z(n18399) );
  XNOR U4086 ( .A(n19136), .B(n18765), .Z(n18767) );
  XNOR U4087 ( .A(n19504), .B(n19133), .Z(n19135) );
  XNOR U4088 ( .A(n19872), .B(n19501), .Z(n19503) );
  XNOR U4089 ( .A(n20240), .B(n19869), .Z(n19871) );
  XNOR U4090 ( .A(n20608), .B(n20237), .Z(n20239) );
  XNOR U4091 ( .A(n20976), .B(n20605), .Z(n20607) );
  XNOR U4092 ( .A(n21344), .B(n20973), .Z(n20975) );
  XNOR U4093 ( .A(n21712), .B(n21341), .Z(n21343) );
  XNOR U4094 ( .A(n22080), .B(n21709), .Z(n21711) );
  XNOR U4095 ( .A(n22448), .B(n22077), .Z(n22079) );
  XNOR U4096 ( .A(n22816), .B(n22445), .Z(n22447) );
  XNOR U4097 ( .A(n23184), .B(n22813), .Z(n22815) );
  XNOR U4098 ( .A(n23178), .B(n23324), .Z(n23182) );
  XNOR U4099 ( .A(n4910), .B(n5079), .Z(n4914) );
  XNOR U4100 ( .A(n4146), .B(n4338), .Z(n4150) );
  XNOR U4101 ( .A(n4103), .B(n4349), .Z(n4111) );
  XNOR U4102 ( .A(n3339), .B(n3609), .Z(n3343) );
  XNOR U4103 ( .A(n3706), .B(n3984), .Z(n3701) );
  XNOR U4104 ( .A(n6419), .B(n6563), .Z(n6423) );
  XNOR U4105 ( .A(n11407), .B(n11547), .Z(n11411) );
  XNOR U4106 ( .A(n12149), .B(n11778), .Z(n11780) );
  XNOR U4107 ( .A(n12885), .B(n12514), .Z(n12516) );
  XNOR U4108 ( .A(n13253), .B(n12882), .Z(n12884) );
  XNOR U4109 ( .A(n13989), .B(n13618), .Z(n13620) );
  XNOR U4110 ( .A(n14357), .B(n13986), .Z(n13988) );
  XNOR U4111 ( .A(n14351), .B(n14491), .Z(n14355) );
  XNOR U4112 ( .A(n15093), .B(n14722), .Z(n14724) );
  XNOR U4113 ( .A(n15461), .B(n15090), .Z(n15092) );
  XNOR U4114 ( .A(n15455), .B(n15595), .Z(n15459) );
  XNOR U4115 ( .A(n17295), .B(n17435), .Z(n17299) );
  XNOR U4116 ( .A(n2579), .B(n2868), .Z(n2583) );
  XNOR U4117 ( .A(n1795), .B(n2131), .Z(n1799) );
  XNOR U4118 ( .A(n1030), .B(n1391), .Z(n1035) );
  XNOR U4119 ( .A(n4132), .B(n4342), .Z(n4140) );
  XNOR U4120 ( .A(n3368), .B(n3602), .Z(n3372) );
  XNOR U4121 ( .A(n4175), .B(n4331), .Z(n4179) );
  XNOR U4122 ( .A(n5307), .B(n5445), .Z(n5311) );
  XNOR U4123 ( .A(n6056), .B(n6190), .Z(n6051) );
  XNOR U4124 ( .A(n16196), .B(n16330), .Z(n16200) );
  XNOR U4125 ( .A(n17306), .B(n16935), .Z(n16937) );
  XNOR U4126 ( .A(n33909), .B(n34038), .Z(n33913) );
  XNOR U4127 ( .A(n33625), .B(n33751), .Z(n33629) );
  XNOR U4128 ( .A(n33314), .B(n33440), .Z(n33318) );
  XNOR U4129 ( .A(n32979), .B(n33108), .Z(n32983) );
  XNOR U4130 ( .A(n32623), .B(n32749), .Z(n32627) );
  XNOR U4131 ( .A(n32240), .B(n32366), .Z(n32244) );
  XNOR U4132 ( .A(n31657), .B(n31962), .Z(n31661) );
  XNOR U4133 ( .A(n31213), .B(n31347), .Z(n31217) );
  XNOR U4134 ( .A(n30745), .B(n30879), .Z(n30749) );
  XNOR U4135 ( .A(n30253), .B(n30387), .Z(n30257) );
  XNOR U4136 ( .A(n29737), .B(n29871), .Z(n29741) );
  XNOR U4137 ( .A(n29197), .B(n29331), .Z(n29201) );
  XNOR U4138 ( .A(n28633), .B(n28767), .Z(n28637) );
  XNOR U4139 ( .A(n28045), .B(n28179), .Z(n28049) );
  XNOR U4140 ( .A(n27433), .B(n27567), .Z(n27437) );
  XNOR U4141 ( .A(n26797), .B(n26931), .Z(n26801) );
  XNOR U4142 ( .A(n26137), .B(n26271), .Z(n26141) );
  XNOR U4143 ( .A(n25453), .B(n25587), .Z(n25457) );
  XNOR U4144 ( .A(n24745), .B(n24879), .Z(n24749) );
  XNOR U4145 ( .A(n24010), .B(n24144), .Z(n24014) );
  XNOR U4146 ( .A(n2565), .B(n2872), .Z(n2573) );
  XNOR U4147 ( .A(n2608), .B(n2861), .Z(n2612) );
  XNOR U4148 ( .A(n4939), .B(n5072), .Z(n4943) );
  XNOR U4149 ( .A(n7544), .B(n7676), .Z(n7548) );
  XNOR U4150 ( .A(n8291), .B(n8420), .Z(n8292) );
  XNOR U4151 ( .A(n9033), .B(n9161), .Z(n9041) );
  XNOR U4152 ( .A(n9776), .B(n9911), .Z(n9780) );
  XNOR U4153 ( .A(n10680), .B(n10807), .Z(n10684) );
  XNOR U4154 ( .A(n12159), .B(n11788), .Z(n11790) );
  XNOR U4155 ( .A(n13263), .B(n12892), .Z(n12894) );
  XNOR U4156 ( .A(n14367), .B(n13996), .Z(n13998) );
  XNOR U4157 ( .A(n17673), .B(n17801), .Z(n17677) );
  XNOR U4158 ( .A(n19151), .B(n18780), .Z(n18782) );
  XNOR U4159 ( .A(n19519), .B(n19148), .Z(n19150) );
  XNOR U4160 ( .A(n19887), .B(n19516), .Z(n19518) );
  XNOR U4161 ( .A(n20255), .B(n19884), .Z(n19886) );
  XNOR U4162 ( .A(n20623), .B(n20252), .Z(n20254) );
  XNOR U4163 ( .A(n20991), .B(n20620), .Z(n20622) );
  XNOR U4164 ( .A(n21359), .B(n20988), .Z(n20990) );
  XNOR U4165 ( .A(n21727), .B(n21356), .Z(n21358) );
  XNOR U4166 ( .A(n22095), .B(n21724), .Z(n21726) );
  XNOR U4167 ( .A(n22463), .B(n22092), .Z(n22094) );
  XNOR U4168 ( .A(n22831), .B(n22460), .Z(n22462) );
  XNOR U4169 ( .A(n23199), .B(n22828), .Z(n22830) );
  XNOR U4170 ( .A(n23193), .B(n23321), .Z(n23197) );
  XNOR U4171 ( .A(n4161), .B(n4335), .Z(n4169) );
  XNOR U4172 ( .A(n3397), .B(n3595), .Z(n3401) );
  XNOR U4173 ( .A(n3358), .B(n3606), .Z(n3353) );
  XNOR U4174 ( .A(n7174), .B(n7303), .Z(n7182) );
  XNOR U4175 ( .A(n11422), .B(n11544), .Z(n11426) );
  XNOR U4176 ( .A(n12164), .B(n11793), .Z(n11795) );
  XNOR U4177 ( .A(n12900), .B(n12529), .Z(n12531) );
  XNOR U4178 ( .A(n13268), .B(n12897), .Z(n12899) );
  XNOR U4179 ( .A(n14004), .B(n13633), .Z(n13635) );
  XNOR U4180 ( .A(n14372), .B(n14001), .Z(n14003) );
  XNOR U4181 ( .A(n15108), .B(n14737), .Z(n14739) );
  XNOR U4182 ( .A(n15476), .B(n15105), .Z(n15107) );
  XNOR U4183 ( .A(n15470), .B(n15592), .Z(n15474) );
  XNOR U4184 ( .A(n16212), .B(n15841), .Z(n15843) );
  XNOR U4185 ( .A(n16580), .B(n16209), .Z(n16211) );
  XNOR U4186 ( .A(n16574), .B(n16696), .Z(n16578) );
  XNOR U4187 ( .A(n18414), .B(n18536), .Z(n18418) );
  XNOR U4188 ( .A(n2637), .B(n2854), .Z(n2641) );
  XNOR U4189 ( .A(n2594), .B(n2865), .Z(n2602) );
  XNOR U4190 ( .A(n1428), .B(n1758), .Z(n1432) );
  XNOR U4191 ( .A(n664), .B(n1018), .Z(n668) );
  XNOR U4192 ( .A(n3387), .B(n3599), .Z(n3382) );
  XNOR U4193 ( .A(n4190), .B(n4328), .Z(n4198) );
  XNOR U4194 ( .A(n3426), .B(n3588), .Z(n3430) );
  XNOR U4195 ( .A(n4204), .B(n4324), .Z(n4208) );
  XNOR U4196 ( .A(n6066), .B(n6186), .Z(n6070) );
  XNOR U4197 ( .A(n6813), .B(n6926), .Z(n6814) );
  XNOR U4198 ( .A(n17315), .B(n17431), .Z(n17319) );
  XNOR U4199 ( .A(n18425), .B(n18054), .Z(n18056) );
  XNOR U4200 ( .A(n34426), .B(n34534), .Z(n34430) );
  XNOR U4201 ( .A(n34187), .B(n34295), .Z(n34191) );
  XNOR U4202 ( .A(n33924), .B(n34035), .Z(n33928) );
  XNOR U4203 ( .A(n33640), .B(n33748), .Z(n33644) );
  XNOR U4204 ( .A(n33329), .B(n33437), .Z(n33333) );
  XNOR U4205 ( .A(n32994), .B(n33105), .Z(n32998) );
  XNOR U4206 ( .A(n32638), .B(n32746), .Z(n32642) );
  XNOR U4207 ( .A(n32255), .B(n32363), .Z(n32259) );
  XNOR U4208 ( .A(n31672), .B(n31959), .Z(n31676) );
  XNOR U4209 ( .A(n31228), .B(n31344), .Z(n31232) );
  XNOR U4210 ( .A(n30760), .B(n30876), .Z(n30764) );
  XNOR U4211 ( .A(n30268), .B(n30384), .Z(n30272) );
  XNOR U4212 ( .A(n29752), .B(n29868), .Z(n29756) );
  XNOR U4213 ( .A(n29212), .B(n29328), .Z(n29216) );
  XNOR U4214 ( .A(n28648), .B(n28764), .Z(n28652) );
  XNOR U4215 ( .A(n28060), .B(n28176), .Z(n28064) );
  XNOR U4216 ( .A(n27448), .B(n27564), .Z(n27452) );
  XNOR U4217 ( .A(n26812), .B(n26928), .Z(n26816) );
  XNOR U4218 ( .A(n26152), .B(n26268), .Z(n26156) );
  XNOR U4219 ( .A(n25468), .B(n25584), .Z(n25472) );
  XNOR U4220 ( .A(n24760), .B(n24876), .Z(n24764) );
  XNOR U4221 ( .A(n24025), .B(n24141), .Z(n24029) );
  XNOR U4222 ( .A(n1819), .B(n2127), .Z(n1814) );
  XNOR U4223 ( .A(n2623), .B(n2858), .Z(n2631) );
  XNOR U4224 ( .A(n2666), .B(n2847), .Z(n2670) );
  XNOR U4225 ( .A(n4956), .B(n5068), .Z(n4957) );
  XNOR U4226 ( .A(n5699), .B(n5813), .Z(n5707) );
  XNOR U4227 ( .A(n8303), .B(n8417), .Z(n8307) );
  XNOR U4228 ( .A(n9047), .B(n9157), .Z(n9051) );
  XNOR U4229 ( .A(n9795), .B(n9908), .Z(n9789) );
  XNOR U4230 ( .A(n10695), .B(n10804), .Z(n10699) );
  XNOR U4231 ( .A(n12174), .B(n11803), .Z(n11805) );
  XNOR U4232 ( .A(n13278), .B(n12907), .Z(n12909) );
  XNOR U4233 ( .A(n14382), .B(n14011), .Z(n14013) );
  XNOR U4234 ( .A(n15486), .B(n15115), .Z(n15117) );
  XNOR U4235 ( .A(n18792), .B(n18902), .Z(n18796) );
  XNOR U4236 ( .A(n20270), .B(n19899), .Z(n19901) );
  XNOR U4237 ( .A(n20638), .B(n20267), .Z(n20269) );
  XNOR U4238 ( .A(n21006), .B(n20635), .Z(n20637) );
  XNOR U4239 ( .A(n21374), .B(n21003), .Z(n21005) );
  XNOR U4240 ( .A(n21742), .B(n21371), .Z(n21373) );
  XNOR U4241 ( .A(n22110), .B(n21739), .Z(n21741) );
  XNOR U4242 ( .A(n22478), .B(n22107), .Z(n22109) );
  XNOR U4243 ( .A(n22846), .B(n22475), .Z(n22477) );
  XNOR U4244 ( .A(n23214), .B(n22843), .Z(n22845) );
  XNOR U4245 ( .A(n23208), .B(n23318), .Z(n23212) );
  XNOR U4246 ( .A(n3455), .B(n3581), .Z(n3459) );
  XNOR U4247 ( .A(n3416), .B(n3592), .Z(n3411) );
  XNOR U4248 ( .A(n1457), .B(n1751), .Z(n1461) );
  XNOR U4249 ( .A(n693), .B(n1011), .Z(n697) );
  XNOR U4250 ( .A(n7940), .B(n8044), .Z(n7935) );
  XNOR U4251 ( .A(n11437), .B(n11541), .Z(n11441) );
  XNOR U4252 ( .A(n12179), .B(n11808), .Z(n11810) );
  XNOR U4253 ( .A(n12915), .B(n12544), .Z(n12546) );
  XNOR U4254 ( .A(n13283), .B(n12912), .Z(n12914) );
  XNOR U4255 ( .A(n14019), .B(n13648), .Z(n13650) );
  XNOR U4256 ( .A(n14387), .B(n14016), .Z(n14018) );
  XNOR U4257 ( .A(n15123), .B(n14752), .Z(n14754) );
  XNOR U4258 ( .A(n15491), .B(n15120), .Z(n15122) );
  XNOR U4259 ( .A(n16227), .B(n15856), .Z(n15858) );
  XNOR U4260 ( .A(n16595), .B(n16224), .Z(n16226) );
  XNOR U4261 ( .A(n16589), .B(n16693), .Z(n16593) );
  XNOR U4262 ( .A(n17331), .B(n16960), .Z(n16962) );
  XNOR U4263 ( .A(n17699), .B(n17328), .Z(n17330) );
  XNOR U4264 ( .A(n17693), .B(n17797), .Z(n17697) );
  XNOR U4265 ( .A(n19533), .B(n19637), .Z(n19537) );
  XNOR U4266 ( .A(n2695), .B(n2840), .Z(n2699) );
  XNOR U4267 ( .A(n2652), .B(n2851), .Z(n2660) );
  XNOR U4268 ( .A(n1848), .B(n2120), .Z(n1843) );
  XNOR U4269 ( .A(n679), .B(n1015), .Z(n687) );
  XNOR U4270 ( .A(n1486), .B(n1744), .Z(n1490) );
  XNOR U4271 ( .A(n722), .B(n1004), .Z(n726) );
  XNOR U4272 ( .A(n3445), .B(n3585), .Z(n3440) );
  XNOR U4273 ( .A(n3102), .B(n3204), .Z(n3106) );
  XNOR U4274 ( .A(n4219), .B(n4321), .Z(n4227) );
  XNOR U4275 ( .A(n6825), .B(n6923), .Z(n6829) );
  XNOR U4276 ( .A(n7568), .B(n7670), .Z(n7572) );
  XNOR U4277 ( .A(n18434), .B(n18532), .Z(n18438) );
  XNOR U4278 ( .A(n19544), .B(n19173), .Z(n19175) );
  XNOR U4279 ( .A(n34653), .B(n34746), .Z(n34657) );
  XNOR U4280 ( .A(n34441), .B(n34531), .Z(n34445) );
  XNOR U4281 ( .A(n34202), .B(n34292), .Z(n34206) );
  XNOR U4282 ( .A(n33939), .B(n34032), .Z(n33943) );
  XNOR U4283 ( .A(n33655), .B(n33745), .Z(n33659) );
  XNOR U4284 ( .A(n33344), .B(n33434), .Z(n33348) );
  XNOR U4285 ( .A(n33009), .B(n33102), .Z(n33013) );
  XNOR U4286 ( .A(n32653), .B(n32743), .Z(n32657) );
  XNOR U4287 ( .A(n32270), .B(n32360), .Z(n32274) );
  XNOR U4288 ( .A(n31687), .B(n31956), .Z(n31691) );
  XNOR U4289 ( .A(n31243), .B(n31341), .Z(n31247) );
  XNOR U4290 ( .A(n30775), .B(n30873), .Z(n30779) );
  XNOR U4291 ( .A(n30283), .B(n30381), .Z(n30287) );
  XNOR U4292 ( .A(n29767), .B(n29865), .Z(n29771) );
  XNOR U4293 ( .A(n29227), .B(n29325), .Z(n29231) );
  XNOR U4294 ( .A(n28663), .B(n28761), .Z(n28667) );
  XNOR U4295 ( .A(n28075), .B(n28173), .Z(n28079) );
  XNOR U4296 ( .A(n27463), .B(n27561), .Z(n27467) );
  XNOR U4297 ( .A(n26827), .B(n26925), .Z(n26831) );
  XNOR U4298 ( .A(n26167), .B(n26265), .Z(n26171) );
  XNOR U4299 ( .A(n25483), .B(n25581), .Z(n25487) );
  XNOR U4300 ( .A(n24775), .B(n24873), .Z(n24779) );
  XNOR U4301 ( .A(n24040), .B(n24138), .Z(n24044) );
  XNOR U4302 ( .A(n1877), .B(n2113), .Z(n1872) );
  XNOR U4303 ( .A(n2681), .B(n2844), .Z(n2689) );
  XNOR U4304 ( .A(n4968), .B(n5065), .Z(n4972) );
  XNOR U4305 ( .A(n5713), .B(n5809), .Z(n5717) );
  XNOR U4306 ( .A(n6462), .B(n6554), .Z(n6457) );
  XNOR U4307 ( .A(n9062), .B(n9154), .Z(n9070) );
  XNOR U4308 ( .A(n9805), .B(n9903), .Z(n9809) );
  XNOR U4309 ( .A(n10710), .B(n10801), .Z(n10714) );
  XNOR U4310 ( .A(n12189), .B(n11818), .Z(n11820) );
  XNOR U4311 ( .A(n13293), .B(n12922), .Z(n12924) );
  XNOR U4312 ( .A(n14397), .B(n14026), .Z(n14028) );
  XNOR U4313 ( .A(n15501), .B(n15130), .Z(n15132) );
  XNOR U4314 ( .A(n16605), .B(n16234), .Z(n16236) );
  XNOR U4315 ( .A(n19911), .B(n20003), .Z(n19915) );
  XNOR U4316 ( .A(n21389), .B(n21018), .Z(n21020) );
  XNOR U4317 ( .A(n21757), .B(n21386), .Z(n21388) );
  XNOR U4318 ( .A(n22125), .B(n21754), .Z(n21756) );
  XNOR U4319 ( .A(n22493), .B(n22122), .Z(n22124) );
  XNOR U4320 ( .A(n22861), .B(n22490), .Z(n22492) );
  XNOR U4321 ( .A(n23229), .B(n22858), .Z(n22860) );
  XNOR U4322 ( .A(n23223), .B(n23315), .Z(n23227) );
  XNOR U4323 ( .A(n3474), .B(n3578), .Z(n3469) );
  XNOR U4324 ( .A(n1515), .B(n1737), .Z(n1519) );
  XNOR U4325 ( .A(n751), .B(n997), .Z(n755) );
  XNOR U4326 ( .A(n708), .B(n1008), .Z(n716) );
  XNOR U4327 ( .A(n8697), .B(n8784), .Z(n8698) );
  XNOR U4328 ( .A(n11452), .B(n11538), .Z(n11456) );
  XNOR U4329 ( .A(n12194), .B(n11823), .Z(n11825) );
  XNOR U4330 ( .A(n12930), .B(n12559), .Z(n12561) );
  XNOR U4331 ( .A(n13298), .B(n12927), .Z(n12929) );
  XNOR U4332 ( .A(n14034), .B(n13663), .Z(n13665) );
  XNOR U4333 ( .A(n14402), .B(n14031), .Z(n14033) );
  XNOR U4334 ( .A(n15138), .B(n14767), .Z(n14769) );
  XNOR U4335 ( .A(n15506), .B(n15135), .Z(n15137) );
  XNOR U4336 ( .A(n16242), .B(n15871), .Z(n15873) );
  XNOR U4337 ( .A(n16610), .B(n16239), .Z(n16241) );
  XNOR U4338 ( .A(n17346), .B(n16975), .Z(n16977) );
  XNOR U4339 ( .A(n17714), .B(n17343), .Z(n17345) );
  XNOR U4340 ( .A(n17708), .B(n17794), .Z(n17712) );
  XNOR U4341 ( .A(n18450), .B(n18079), .Z(n18081) );
  XNOR U4342 ( .A(n18818), .B(n18447), .Z(n18449) );
  XNOR U4343 ( .A(n18812), .B(n18898), .Z(n18816) );
  XNOR U4344 ( .A(n20652), .B(n20738), .Z(n20656) );
  XNOR U4345 ( .A(n2710), .B(n2837), .Z(n2718) );
  XNOR U4346 ( .A(n1906), .B(n2106), .Z(n1901) );
  XNOR U4347 ( .A(n737), .B(n1001), .Z(n745) );
  XNOR U4348 ( .A(n1544), .B(n1730), .Z(n1548) );
  XNOR U4349 ( .A(n780), .B(n990), .Z(n784) );
  XNOR U4350 ( .A(n2734), .B(n2831), .Z(n2738) );
  XNOR U4351 ( .A(n7583), .B(n7667), .Z(n7591) );
  XNOR U4352 ( .A(n8327), .B(n8411), .Z(n8331) );
  XNOR U4353 ( .A(n19553), .B(n19633), .Z(n19557) );
  XNOR U4354 ( .A(n20663), .B(n20292), .Z(n20294) );
  XNOR U4355 ( .A(n35026), .B(n35098), .Z(n35030) );
  XNOR U4356 ( .A(n34859), .B(n34931), .Z(n34863) );
  XNOR U4357 ( .A(n34668), .B(n34743), .Z(n34672) );
  XNOR U4358 ( .A(n34456), .B(n34528), .Z(n34460) );
  XNOR U4359 ( .A(n34217), .B(n34289), .Z(n34221) );
  XNOR U4360 ( .A(n33954), .B(n34029), .Z(n33958) );
  XNOR U4361 ( .A(n33670), .B(n33742), .Z(n33674) );
  XNOR U4362 ( .A(n33359), .B(n33431), .Z(n33363) );
  XNOR U4363 ( .A(n33024), .B(n33099), .Z(n33028) );
  XNOR U4364 ( .A(n32668), .B(n32740), .Z(n32672) );
  XNOR U4365 ( .A(n32285), .B(n32357), .Z(n32289) );
  XNOR U4366 ( .A(n31702), .B(n31953), .Z(n31706) );
  XNOR U4367 ( .A(n31258), .B(n31338), .Z(n31262) );
  XNOR U4368 ( .A(n30790), .B(n30870), .Z(n30794) );
  XNOR U4369 ( .A(n30298), .B(n30378), .Z(n30302) );
  XNOR U4370 ( .A(n29782), .B(n29862), .Z(n29786) );
  XNOR U4371 ( .A(n29242), .B(n29322), .Z(n29246) );
  XNOR U4372 ( .A(n28678), .B(n28758), .Z(n28682) );
  XNOR U4373 ( .A(n28090), .B(n28170), .Z(n28094) );
  XNOR U4374 ( .A(n27478), .B(n27558), .Z(n27482) );
  XNOR U4375 ( .A(n26842), .B(n26922), .Z(n26846) );
  XNOR U4376 ( .A(n26182), .B(n26262), .Z(n26186) );
  XNOR U4377 ( .A(n25498), .B(n25578), .Z(n25502) );
  XNOR U4378 ( .A(n24790), .B(n24870), .Z(n24794) );
  XNOR U4379 ( .A(n24055), .B(n24135), .Z(n24059) );
  XNOR U4380 ( .A(n1935), .B(n2099), .Z(n1930) );
  XNOR U4381 ( .A(n2751), .B(n2827), .Z(n2752) );
  XNOR U4382 ( .A(n3494), .B(n3572), .Z(n3502) );
  XNOR U4383 ( .A(n4238), .B(n4316), .Z(n4242) );
  XNOR U4384 ( .A(n4985), .B(n5061), .Z(n4986) );
  XNOR U4385 ( .A(n5728), .B(n5806), .Z(n5736) );
  XNOR U4386 ( .A(n6472), .B(n6550), .Z(n6476) );
  XNOR U4387 ( .A(n7215), .B(n7293), .Z(n7216) );
  XNOR U4388 ( .A(n9824), .B(n9900), .Z(n9818) );
  XNOR U4389 ( .A(n10725), .B(n10798), .Z(n10729) );
  XNOR U4390 ( .A(n12204), .B(n11833), .Z(n11835) );
  XNOR U4391 ( .A(n13308), .B(n12937), .Z(n12939) );
  XNOR U4392 ( .A(n14412), .B(n14041), .Z(n14043) );
  XNOR U4393 ( .A(n15516), .B(n15145), .Z(n15147) );
  XNOR U4394 ( .A(n16620), .B(n16249), .Z(n16251) );
  XNOR U4395 ( .A(n17724), .B(n17353), .Z(n17355) );
  XNOR U4396 ( .A(n21030), .B(n21104), .Z(n21034) );
  XNOR U4397 ( .A(n22508), .B(n22137), .Z(n22139) );
  XNOR U4398 ( .A(n22876), .B(n22505), .Z(n22507) );
  XNOR U4399 ( .A(n23244), .B(n22873), .Z(n22875) );
  XNOR U4400 ( .A(n23238), .B(n23312), .Z(n23242) );
  XNOR U4401 ( .A(n1573), .B(n1723), .Z(n1577) );
  XNOR U4402 ( .A(n809), .B(n983), .Z(n813) );
  XNOR U4403 ( .A(n766), .B(n994), .Z(n774) );
  XNOR U4404 ( .A(n9449), .B(n9524), .Z(n9453) );
  XNOR U4405 ( .A(n11467), .B(n11535), .Z(n11471) );
  XNOR U4406 ( .A(n12209), .B(n11838), .Z(n11840) );
  XNOR U4407 ( .A(n12945), .B(n12574), .Z(n12576) );
  XNOR U4408 ( .A(n13313), .B(n12942), .Z(n12944) );
  XNOR U4409 ( .A(n14049), .B(n13678), .Z(n13680) );
  XNOR U4410 ( .A(n14417), .B(n14046), .Z(n14048) );
  XNOR U4411 ( .A(n15153), .B(n14782), .Z(n14784) );
  XNOR U4412 ( .A(n15521), .B(n15150), .Z(n15152) );
  XNOR U4413 ( .A(n16257), .B(n15886), .Z(n15888) );
  XNOR U4414 ( .A(n16625), .B(n16254), .Z(n16256) );
  XNOR U4415 ( .A(n17361), .B(n16990), .Z(n16992) );
  XNOR U4416 ( .A(n17729), .B(n17358), .Z(n17360) );
  XNOR U4417 ( .A(n18465), .B(n18094), .Z(n18096) );
  XNOR U4418 ( .A(n18833), .B(n18462), .Z(n18464) );
  XNOR U4419 ( .A(n18827), .B(n18895), .Z(n18831) );
  XNOR U4420 ( .A(n19569), .B(n19198), .Z(n19200) );
  XNOR U4421 ( .A(n19937), .B(n19566), .Z(n19568) );
  XNOR U4422 ( .A(n19931), .B(n19999), .Z(n19935) );
  XNOR U4423 ( .A(n21771), .B(n21839), .Z(n21775) );
  XNOR U4424 ( .A(n1242), .B(n1341), .Z(n1243) );
  XNOR U4425 ( .A(n1964), .B(n2092), .Z(n1959) );
  XNOR U4426 ( .A(n795), .B(n987), .Z(n803) );
  XNOR U4427 ( .A(n1602), .B(n1716), .Z(n1606) );
  XNOR U4428 ( .A(n838), .B(n976), .Z(n842) );
  XNOR U4429 ( .A(n8346), .B(n8408), .Z(n8341) );
  XNOR U4430 ( .A(n9086), .B(n9148), .Z(n9090) );
  XNOR U4431 ( .A(n20672), .B(n20734), .Z(n20676) );
  XNOR U4432 ( .A(n21782), .B(n21411), .Z(n21413) );
  XNOR U4433 ( .A(n35181), .B(n35238), .Z(n35185) );
  XNOR U4434 ( .A(n35041), .B(n35095), .Z(n35045) );
  XNOR U4435 ( .A(n34874), .B(n34928), .Z(n34878) );
  XNOR U4436 ( .A(n34683), .B(n34740), .Z(n34687) );
  XNOR U4437 ( .A(n34471), .B(n34525), .Z(n34475) );
  XNOR U4438 ( .A(n34232), .B(n34286), .Z(n34236) );
  XNOR U4439 ( .A(n33969), .B(n34026), .Z(n33973) );
  XNOR U4440 ( .A(n33685), .B(n33739), .Z(n33689) );
  XNOR U4441 ( .A(n33374), .B(n33428), .Z(n33378) );
  XNOR U4442 ( .A(n33039), .B(n33096), .Z(n33043) );
  XNOR U4443 ( .A(n32683), .B(n32737), .Z(n32687) );
  XNOR U4444 ( .A(n32300), .B(n32354), .Z(n32304) );
  XNOR U4445 ( .A(n31717), .B(n31950), .Z(n31721) );
  XNOR U4446 ( .A(n31273), .B(n31335), .Z(n31277) );
  XNOR U4447 ( .A(n30805), .B(n30867), .Z(n30809) );
  XNOR U4448 ( .A(n30313), .B(n30375), .Z(n30317) );
  XNOR U4449 ( .A(n29797), .B(n29859), .Z(n29801) );
  XNOR U4450 ( .A(n29257), .B(n29319), .Z(n29261) );
  XNOR U4451 ( .A(n28693), .B(n28755), .Z(n28697) );
  XNOR U4452 ( .A(n28105), .B(n28167), .Z(n28109) );
  XNOR U4453 ( .A(n27493), .B(n27555), .Z(n27497) );
  XNOR U4454 ( .A(n26857), .B(n26919), .Z(n26861) );
  XNOR U4455 ( .A(n26197), .B(n26259), .Z(n26201) );
  XNOR U4456 ( .A(n25513), .B(n25575), .Z(n25517) );
  XNOR U4457 ( .A(n24805), .B(n24867), .Z(n24809) );
  XNOR U4458 ( .A(n24070), .B(n24132), .Z(n24074) );
  XNOR U4459 ( .A(n1993), .B(n2085), .Z(n1988) );
  XNOR U4460 ( .A(n2018), .B(n2078), .Z(n2022) );
  XNOR U4461 ( .A(n2763), .B(n2824), .Z(n2767) );
  XNOR U4462 ( .A(n3508), .B(n3568), .Z(n3512) );
  XNOR U4463 ( .A(n4257), .B(n4313), .Z(n4252) );
  XNOR U4464 ( .A(n4997), .B(n5058), .Z(n5001) );
  XNOR U4465 ( .A(n5742), .B(n5802), .Z(n5746) );
  XNOR U4466 ( .A(n6491), .B(n6547), .Z(n6486) );
  XNOR U4467 ( .A(n7227), .B(n7290), .Z(n7231) );
  XNOR U4468 ( .A(n7974), .B(n8034), .Z(n7978) );
  XNOR U4469 ( .A(n10740), .B(n10795), .Z(n10744) );
  XNOR U4470 ( .A(n12219), .B(n11848), .Z(n11850) );
  XNOR U4471 ( .A(n13323), .B(n12952), .Z(n12954) );
  XNOR U4472 ( .A(n14427), .B(n14056), .Z(n14058) );
  XNOR U4473 ( .A(n15531), .B(n15160), .Z(n15162) );
  XNOR U4474 ( .A(n16635), .B(n16264), .Z(n16266) );
  XNOR U4475 ( .A(n17739), .B(n17368), .Z(n17370) );
  XNOR U4476 ( .A(n18843), .B(n18472), .Z(n18474) );
  XNOR U4477 ( .A(n22885), .B(n22941), .Z(n22889) );
  XNOR U4478 ( .A(n23253), .B(n23309), .Z(n23257) );
  XNOR U4479 ( .A(n824), .B(n980), .Z(n832) );
  XNOR U4480 ( .A(n10216), .B(n10378), .Z(n10220) );
  XNOR U4481 ( .A(n11482), .B(n11532), .Z(n11486) );
  XNOR U4482 ( .A(n12224), .B(n11853), .Z(n11855) );
  XNOR U4483 ( .A(n12960), .B(n12589), .Z(n12591) );
  XNOR U4484 ( .A(n13328), .B(n12957), .Z(n12959) );
  XNOR U4485 ( .A(n14064), .B(n13693), .Z(n13695) );
  XNOR U4486 ( .A(n14432), .B(n14061), .Z(n14063) );
  XNOR U4487 ( .A(n15168), .B(n14797), .Z(n14799) );
  XNOR U4488 ( .A(n15536), .B(n15165), .Z(n15167) );
  XNOR U4489 ( .A(n16272), .B(n15901), .Z(n15903) );
  XNOR U4490 ( .A(n16640), .B(n16269), .Z(n16271) );
  XNOR U4491 ( .A(n17376), .B(n17005), .Z(n17007) );
  XNOR U4492 ( .A(n17744), .B(n17373), .Z(n17375) );
  XNOR U4493 ( .A(n18480), .B(n18109), .Z(n18111) );
  XNOR U4494 ( .A(n18848), .B(n18477), .Z(n18479) );
  XNOR U4495 ( .A(n19584), .B(n19213), .Z(n19215) );
  XNOR U4496 ( .A(n19952), .B(n19581), .Z(n19583) );
  XNOR U4497 ( .A(n19946), .B(n19996), .Z(n19950) );
  XNOR U4498 ( .A(n20688), .B(n20317), .Z(n20319) );
  XNOR U4499 ( .A(n21056), .B(n20685), .Z(n20687) );
  XNOR U4500 ( .A(n21050), .B(n21100), .Z(n21054) );
  XNOR U4501 ( .A(n22522), .B(n22572), .Z(n22526) );
  XNOR U4502 ( .A(n872), .B(n968), .Z(n876) );
  XNOR U4503 ( .A(n853), .B(n973), .Z(n861) );
  XNOR U4504 ( .A(n9103), .B(n9144), .Z(n9104) );
  XNOR U4505 ( .A(n9844), .B(n9893), .Z(n9852) );
  XNOR U4506 ( .A(n21791), .B(n21835), .Z(n21795) );
  XNOR U4507 ( .A(n35364), .B(n35403), .Z(n35368) );
  XNOR U4508 ( .A(n35260), .B(n35296), .Z(n35264) );
  XNOR U4509 ( .A(n35129), .B(n35165), .Z(n35133) );
  XNOR U4510 ( .A(n34974), .B(n35013), .Z(n34978) );
  XNOR U4511 ( .A(n34798), .B(n34834), .Z(n34802) );
  XNOR U4512 ( .A(n34595), .B(n34631), .Z(n34599) );
  XNOR U4513 ( .A(n34368), .B(n34407), .Z(n34372) );
  XNOR U4514 ( .A(n34120), .B(n34156), .Z(n34124) );
  XNOR U4515 ( .A(n33845), .B(n33881), .Z(n33849) );
  XNOR U4516 ( .A(n33546), .B(n33585), .Z(n33550) );
  XNOR U4517 ( .A(n33226), .B(n33262), .Z(n33230) );
  XNOR U4518 ( .A(n32879), .B(n32915), .Z(n32883) );
  XNOR U4519 ( .A(n32508), .B(n32547), .Z(n32512) );
  XNOR U4520 ( .A(n32116), .B(n32152), .Z(n32120) );
  XNOR U4521 ( .A(n31513), .B(n31557), .Z(n31517) );
  XNOR U4522 ( .A(n31057), .B(n31101), .Z(n31061) );
  XNOR U4523 ( .A(n30577), .B(n30621), .Z(n30581) );
  XNOR U4524 ( .A(n30073), .B(n30117), .Z(n30077) );
  XNOR U4525 ( .A(n29545), .B(n29589), .Z(n29549) );
  XNOR U4526 ( .A(n28993), .B(n29037), .Z(n28997) );
  XNOR U4527 ( .A(n28417), .B(n28461), .Z(n28421) );
  XNOR U4528 ( .A(n27817), .B(n27861), .Z(n27821) );
  XNOR U4529 ( .A(n27193), .B(n27237), .Z(n27197) );
  XNOR U4530 ( .A(n26545), .B(n26589), .Z(n26549) );
  XNOR U4531 ( .A(n25873), .B(n25917), .Z(n25877) );
  XNOR U4532 ( .A(n25177), .B(n25221), .Z(n25181) );
  XNOR U4533 ( .A(n24457), .B(n24501), .Z(n24461) );
  XNOR U4534 ( .A(n23636), .B(n23755), .Z(n23640) );
  XNOR U4535 ( .A(n1259), .B(n1337), .Z(n1263) );
  XNOR U4536 ( .A(n902), .B(n962), .Z(n906) );
  XNOR U4537 ( .A(n2405), .B(n2447), .Z(n2409) );
  XNOR U4538 ( .A(n3151), .B(n3193), .Z(n3155) );
  XNOR U4539 ( .A(n3895), .B(n3937), .Z(n3899) );
  XNOR U4540 ( .A(n4639), .B(n4681), .Z(n4643) );
  XNOR U4541 ( .A(n5389), .B(n5427), .Z(n5384) );
  XNOR U4542 ( .A(n6129), .B(n6171), .Z(n6133) );
  XNOR U4543 ( .A(n6873), .B(n6911), .Z(n6877) );
  XNOR U4544 ( .A(n7621), .B(n7659), .Z(n7616) );
  XNOR U4545 ( .A(n8361), .B(n8403), .Z(n8365) );
  XNOR U4546 ( .A(n10755), .B(n10792), .Z(n10759) );
  XNOR U4547 ( .A(n12234), .B(n11863), .Z(n11865) );
  XNOR U4548 ( .A(n13338), .B(n12967), .Z(n12969) );
  XNOR U4549 ( .A(n14442), .B(n14071), .Z(n14073) );
  XNOR U4550 ( .A(n15546), .B(n15175), .Z(n15177) );
  XNOR U4551 ( .A(n16650), .B(n16279), .Z(n16281) );
  XNOR U4552 ( .A(n17754), .B(n17383), .Z(n17385) );
  XNOR U4553 ( .A(n18858), .B(n18487), .Z(n18489) );
  XNOR U4554 ( .A(n19962), .B(n19591), .Z(n19593) );
  XNOR U4555 ( .A(n1289), .B(n1331), .Z(n1293) );
  XNOR U4556 ( .A(n11134), .B(n10763), .Z(n10765) );
  XNOR U4557 ( .A(n11497), .B(n11529), .Z(n11501) );
  XNOR U4558 ( .A(n12239), .B(n11868), .Z(n11870) );
  XNOR U4559 ( .A(n12975), .B(n12604), .Z(n12606) );
  XNOR U4560 ( .A(n13343), .B(n12972), .Z(n12974) );
  XNOR U4561 ( .A(n14079), .B(n13708), .Z(n13710) );
  XNOR U4562 ( .A(n14447), .B(n14076), .Z(n14078) );
  XNOR U4563 ( .A(n15183), .B(n14812), .Z(n14814) );
  XNOR U4564 ( .A(n15551), .B(n15180), .Z(n15182) );
  XNOR U4565 ( .A(n16287), .B(n15916), .Z(n15918) );
  XNOR U4566 ( .A(n16655), .B(n16284), .Z(n16286) );
  XNOR U4567 ( .A(n17391), .B(n17020), .Z(n17022) );
  XNOR U4568 ( .A(n17759), .B(n17388), .Z(n17390) );
  XNOR U4569 ( .A(n18495), .B(n18124), .Z(n18126) );
  XNOR U4570 ( .A(n18863), .B(n18492), .Z(n18494) );
  XNOR U4571 ( .A(n19599), .B(n19228), .Z(n19230) );
  XNOR U4572 ( .A(n19967), .B(n19596), .Z(n19598) );
  XNOR U4573 ( .A(n20703), .B(n20332), .Z(n20334) );
  XNOR U4574 ( .A(n21071), .B(n20700), .Z(n20702) );
  XNOR U4575 ( .A(n21065), .B(n21097), .Z(n21069) );
  XNOR U4576 ( .A(n22175), .B(n21804), .Z(n21806) );
  XNOR U4577 ( .A(n22169), .B(n22201), .Z(n22173) );
  XNOR U4578 ( .A(n22905), .B(n22937), .Z(n22909) );
  XNOR U4579 ( .A(n9483), .B(n9516), .Z(n9487) );
  XNOR U4580 ( .A(n10230), .B(n10371), .Z(n10239) );
  XNOR U4581 ( .A(n35493), .B(n35514), .Z(n35497) );
  XNOR U4582 ( .A(n35425), .B(n35443), .Z(n35429) );
  XNOR U4583 ( .A(n35330), .B(n35348), .Z(n35334) );
  XNOR U4584 ( .A(n35211), .B(n35232), .Z(n35215) );
  XNOR U4585 ( .A(n35071), .B(n35089), .Z(n35075) );
  XNOR U4586 ( .A(n34904), .B(n34922), .Z(n34908) );
  XNOR U4587 ( .A(n34713), .B(n34734), .Z(n34717) );
  XNOR U4588 ( .A(n34501), .B(n34519), .Z(n34505) );
  XNOR U4589 ( .A(n34262), .B(n34280), .Z(n34266) );
  XNOR U4590 ( .A(n33999), .B(n34020), .Z(n34003) );
  XNOR U4591 ( .A(n33715), .B(n33733), .Z(n33719) );
  XNOR U4592 ( .A(n33404), .B(n33422), .Z(n33408) );
  XNOR U4593 ( .A(n33069), .B(n33090), .Z(n33073) );
  XNOR U4594 ( .A(n32713), .B(n32731), .Z(n32717) );
  XNOR U4595 ( .A(n32330), .B(n32348), .Z(n32334) );
  XNOR U4596 ( .A(n31747), .B(n31944), .Z(n31751) );
  XNOR U4597 ( .A(n31303), .B(n31329), .Z(n31307) );
  XNOR U4598 ( .A(n30835), .B(n30861), .Z(n30839) );
  XNOR U4599 ( .A(n30343), .B(n30369), .Z(n30347) );
  XNOR U4600 ( .A(n29827), .B(n29853), .Z(n29831) );
  XNOR U4601 ( .A(n29287), .B(n29313), .Z(n29291) );
  XNOR U4602 ( .A(n28723), .B(n28749), .Z(n28727) );
  XNOR U4603 ( .A(n28135), .B(n28161), .Z(n28139) );
  XNOR U4604 ( .A(n27523), .B(n27549), .Z(n27527) );
  XNOR U4605 ( .A(n26887), .B(n26913), .Z(n26891) );
  XNOR U4606 ( .A(n26227), .B(n26253), .Z(n26231) );
  XNOR U4607 ( .A(n25543), .B(n25569), .Z(n25547) );
  XNOR U4608 ( .A(n24835), .B(n24861), .Z(n24839) );
  XNOR U4609 ( .A(n24100), .B(n24126), .Z(n24104) );
  XNOR U4610 ( .A(n932), .B(n956), .Z(n936) );
  XNOR U4611 ( .A(n1676), .B(n1700), .Z(n1680) );
  XNOR U4612 ( .A(n3166), .B(n3190), .Z(n3170) );
  XNOR U4613 ( .A(n3910), .B(n3934), .Z(n3914) );
  XNOR U4614 ( .A(n4654), .B(n4678), .Z(n4658) );
  XNOR U4615 ( .A(n5399), .B(n5423), .Z(n5403) );
  XNOR U4616 ( .A(n6146), .B(n6167), .Z(n6147) );
  XNOR U4617 ( .A(n7631), .B(n7655), .Z(n7635) );
  XNOR U4618 ( .A(n8378), .B(n8399), .Z(n8379) );
  XNOR U4619 ( .A(n12249), .B(n11878), .Z(n11880) );
  XNOR U4620 ( .A(n13353), .B(n12982), .Z(n12984) );
  XNOR U4621 ( .A(n14457), .B(n14086), .Z(n14088) );
  XNOR U4622 ( .A(n15561), .B(n15190), .Z(n15192) );
  XNOR U4623 ( .A(n16665), .B(n16294), .Z(n16296) );
  XNOR U4624 ( .A(n17769), .B(n17398), .Z(n17400) );
  XNOR U4625 ( .A(n18873), .B(n18502), .Z(n18504) );
  XNOR U4626 ( .A(n19977), .B(n19606), .Z(n19608) );
  XNOR U4627 ( .A(n21081), .B(n20710), .Z(n20712) );
  XNOR U4628 ( .A(n22553), .B(n22182), .Z(n22184) );
  XNOR U4629 ( .A(n23656), .B(n23751), .Z(n23660) );
  XNOR U4630 ( .A(n2425), .B(n2443), .Z(n2433) );
  XNOR U4631 ( .A(n6897), .B(n6907), .Z(n6891) );
  XNOR U4632 ( .A(n9129), .B(n9139), .Z(n9123) );
  XNOR U4633 ( .A(n10775), .B(n10788), .Z(n10779) );
  XNOR U4634 ( .A(n11886), .B(n11515), .Z(n11517) );
  XNOR U4635 ( .A(n12254), .B(n11883), .Z(n11885) );
  XNOR U4636 ( .A(n12990), .B(n12619), .Z(n12621) );
  XNOR U4637 ( .A(n13358), .B(n12987), .Z(n12989) );
  XNOR U4638 ( .A(n14094), .B(n13723), .Z(n13725) );
  XNOR U4639 ( .A(n14462), .B(n14091), .Z(n14093) );
  XNOR U4640 ( .A(n15198), .B(n14827), .Z(n14829) );
  XNOR U4641 ( .A(n15566), .B(n15195), .Z(n15197) );
  XNOR U4642 ( .A(n16302), .B(n15931), .Z(n15933) );
  XNOR U4643 ( .A(n16670), .B(n16299), .Z(n16301) );
  XNOR U4644 ( .A(n17406), .B(n17035), .Z(n17037) );
  XNOR U4645 ( .A(n17774), .B(n17403), .Z(n17405) );
  XNOR U4646 ( .A(n18510), .B(n18139), .Z(n18141) );
  XNOR U4647 ( .A(n18878), .B(n18507), .Z(n18509) );
  XNOR U4648 ( .A(n19614), .B(n19243), .Z(n19245) );
  XNOR U4649 ( .A(n19982), .B(n19611), .Z(n19613) );
  XNOR U4650 ( .A(n20718), .B(n20347), .Z(n20349) );
  XNOR U4651 ( .A(n21086), .B(n20715), .Z(n20717) );
  XNOR U4652 ( .A(n21822), .B(n21451), .Z(n21453) );
  XNOR U4653 ( .A(n22190), .B(n21819), .Z(n21821) );
  XNOR U4654 ( .A(n22558), .B(n22187), .Z(n22189) );
  XNOR U4655 ( .A(n23294), .B(n22923), .Z(n22925) );
  XNOR U4656 ( .A(n23662), .B(n23291), .Z(n23293) );
  XOR U4657 ( .A(n10254), .B(n10366), .Z(n10248) );
  NANDN U4658 ( .A(n948), .B(n947), .Z(n444) );
  NANDN U4659 ( .A(n2435), .B(n2436), .Z(n2063) );
  NANDN U4660 ( .A(n3925), .B(n3926), .Z(n3553) );
  XOR U4661 ( .A(n4675), .B(n5041), .Z(n5043) );
  XOR U4662 ( .A(n5792), .B(n6158), .Z(n6160) );
  XOR U4663 ( .A(n7267), .B(n7274), .Z(n7276) );
  XNOR U4664 ( .A(n8390), .B(n8392), .Z(n8391) );
  XNOR U4665 ( .A(n9506), .B(n9508), .Z(n9507) );
  XOR U4666 ( .A(n10262), .B(n5), .Z(n10261) );
  XOR U4667 ( .A(n10271), .B(n11), .Z(n10270) );
  XOR U4668 ( .A(n10280), .B(n17), .Z(n10279) );
  XOR U4669 ( .A(n10289), .B(n23), .Z(n10288) );
  XOR U4670 ( .A(n10298), .B(n29), .Z(n10297) );
  XOR U4671 ( .A(n10307), .B(n35), .Z(n10306) );
  XOR U4672 ( .A(n10316), .B(n41), .Z(n10315) );
  XOR U4673 ( .A(n10325), .B(n47), .Z(n10324) );
  XOR U4674 ( .A(n10334), .B(n53), .Z(n10333) );
  XOR U4675 ( .A(n10343), .B(n59), .Z(n10342) );
  XOR U4676 ( .A(n10355), .B(n67), .Z(n10354) );
  XNOR U4677 ( .A(n24192), .B(n24554), .Z(n24196) );
  XNOR U4678 ( .A(n23371), .B(n23808), .Z(n23376) );
  XNOR U4679 ( .A(n10864), .B(n10493), .Z(n10495) );
  XNOR U4680 ( .A(n11233), .B(n10861), .Z(n10863) );
  XNOR U4681 ( .A(n11599), .B(n11952), .Z(n11595) );
  XNOR U4682 ( .A(n12331), .B(n12688), .Z(n12336) );
  XNOR U4683 ( .A(n13067), .B(n13424), .Z(n13072) );
  XNOR U4684 ( .A(n13803), .B(n14160), .Z(n13808) );
  XNOR U4685 ( .A(n14539), .B(n14896), .Z(n14544) );
  XNOR U4686 ( .A(n15275), .B(n15632), .Z(n15280) );
  XNOR U4687 ( .A(n16011), .B(n16368), .Z(n16016) );
  XNOR U4688 ( .A(n16747), .B(n17104), .Z(n16752) );
  XNOR U4689 ( .A(n17483), .B(n17840), .Z(n17488) );
  XNOR U4690 ( .A(n18219), .B(n18576), .Z(n18224) );
  XNOR U4691 ( .A(n18955), .B(n19312), .Z(n18960) );
  XNOR U4692 ( .A(n19691), .B(n20048), .Z(n19696) );
  XNOR U4693 ( .A(n20427), .B(n20784), .Z(n20432) );
  XNOR U4694 ( .A(n21163), .B(n21520), .Z(n21168) );
  XNOR U4695 ( .A(n21899), .B(n22256), .Z(n21904) );
  XNOR U4696 ( .A(n22635), .B(n22992), .Z(n22640) );
  XNOR U4697 ( .A(n7734), .B(n8088), .Z(n7738) );
  XNOR U4698 ( .A(n8855), .B(n9199), .Z(n8859) );
  XNOR U4699 ( .A(n9598), .B(n9951), .Z(n9602) );
  XNOR U4700 ( .A(n24927), .B(n25271), .Z(n24931) );
  XNOR U4701 ( .A(n24207), .B(n24551), .Z(n24211) );
  XNOR U4702 ( .A(n23387), .B(n23805), .Z(n23391) );
  XNOR U4703 ( .A(n10879), .B(n10508), .Z(n10510) );
  XNOR U4704 ( .A(n11248), .B(n10876), .Z(n10878) );
  XNOR U4705 ( .A(n11616), .B(n11245), .Z(n11247) );
  XNOR U4706 ( .A(n11610), .B(n11948), .Z(n11614) );
  XNOR U4707 ( .A(n11978), .B(n12316), .Z(n11982) );
  XNOR U4708 ( .A(n12341), .B(n12684), .Z(n12350) );
  XNOR U4709 ( .A(n13083), .B(n13421), .Z(n13091) );
  XNOR U4710 ( .A(n13819), .B(n14157), .Z(n13823) );
  XNOR U4711 ( .A(n14555), .B(n14893), .Z(n14559) );
  XNOR U4712 ( .A(n15291), .B(n15629), .Z(n15295) );
  XNOR U4713 ( .A(n16027), .B(n16365), .Z(n16031) );
  XNOR U4714 ( .A(n16763), .B(n17101), .Z(n16767) );
  XNOR U4715 ( .A(n17499), .B(n17837), .Z(n17503) );
  XNOR U4716 ( .A(n18235), .B(n18573), .Z(n18239) );
  XNOR U4717 ( .A(n18971), .B(n19309), .Z(n18975) );
  XNOR U4718 ( .A(n19707), .B(n20045), .Z(n19711) );
  XNOR U4719 ( .A(n20443), .B(n20781), .Z(n20447) );
  XNOR U4720 ( .A(n21179), .B(n21517), .Z(n21183) );
  XNOR U4721 ( .A(n21915), .B(n22253), .Z(n21919) );
  XNOR U4722 ( .A(n22651), .B(n22989), .Z(n22655) );
  XNOR U4723 ( .A(n8121), .B(n8457), .Z(n8125) );
  XNOR U4724 ( .A(n6981), .B(n7345), .Z(n6986) );
  XNOR U4725 ( .A(n8870), .B(n9196), .Z(n8874) );
  XNOR U4726 ( .A(n9613), .B(n9948), .Z(n9617) );
  XNOR U4727 ( .A(n26310), .B(n26636), .Z(n26314) );
  XNOR U4728 ( .A(n25638), .B(n25964), .Z(n25642) );
  XNOR U4729 ( .A(n24942), .B(n25268), .Z(n24946) );
  XNOR U4730 ( .A(n24222), .B(n24548), .Z(n24226) );
  XNOR U4731 ( .A(n23402), .B(n23802), .Z(n23406) );
  XNOR U4732 ( .A(n7754), .B(n8084), .Z(n7758) );
  XNOR U4733 ( .A(n10894), .B(n10523), .Z(n10525) );
  XNOR U4734 ( .A(n11263), .B(n10891), .Z(n10893) );
  XNOR U4735 ( .A(n11631), .B(n11260), .Z(n11262) );
  XNOR U4736 ( .A(n11625), .B(n11945), .Z(n11629) );
  XNOR U4737 ( .A(n11993), .B(n12313), .Z(n11997) );
  XNOR U4738 ( .A(n12361), .B(n12681), .Z(n12365) );
  XNOR U4739 ( .A(n12729), .B(n13049), .Z(n12733) );
  XNOR U4740 ( .A(n13097), .B(n13417), .Z(n13101) );
  XNOR U4741 ( .A(n13838), .B(n14154), .Z(n13833) );
  XNOR U4742 ( .A(n14570), .B(n14890), .Z(n14574) );
  XNOR U4743 ( .A(n15306), .B(n15626), .Z(n15310) );
  XNOR U4744 ( .A(n16042), .B(n16362), .Z(n16046) );
  XNOR U4745 ( .A(n16778), .B(n17098), .Z(n16782) );
  XNOR U4746 ( .A(n17514), .B(n17834), .Z(n17518) );
  XNOR U4747 ( .A(n18250), .B(n18570), .Z(n18254) );
  XNOR U4748 ( .A(n18986), .B(n19306), .Z(n18990) );
  XNOR U4749 ( .A(n19722), .B(n20042), .Z(n19726) );
  XNOR U4750 ( .A(n20458), .B(n20778), .Z(n20462) );
  XNOR U4751 ( .A(n21194), .B(n21514), .Z(n21198) );
  XNOR U4752 ( .A(n21930), .B(n22250), .Z(n21934) );
  XNOR U4753 ( .A(n22666), .B(n22986), .Z(n22670) );
  XNOR U4754 ( .A(n6619), .B(n6969), .Z(n6623) );
  XNOR U4755 ( .A(n8141), .B(n8453), .Z(n8145) );
  XNOR U4756 ( .A(n8885), .B(n9193), .Z(n8889) );
  XNOR U4757 ( .A(n9628), .B(n9945), .Z(n9632) );
  XNOR U4758 ( .A(n26973), .B(n27281), .Z(n26977) );
  XNOR U4759 ( .A(n26325), .B(n26633), .Z(n26329) );
  XNOR U4760 ( .A(n25653), .B(n25961), .Z(n25657) );
  XNOR U4761 ( .A(n24957), .B(n25265), .Z(n24961) );
  XNOR U4762 ( .A(n24237), .B(n24545), .Z(n24241) );
  XNOR U4763 ( .A(n23417), .B(n23799), .Z(n23421) );
  XNOR U4764 ( .A(n10909), .B(n10538), .Z(n10540) );
  XNOR U4765 ( .A(n11278), .B(n10906), .Z(n10908) );
  XNOR U4766 ( .A(n11646), .B(n11275), .Z(n11277) );
  XNOR U4767 ( .A(n11640), .B(n11942), .Z(n11644) );
  XNOR U4768 ( .A(n12008), .B(n12310), .Z(n12012) );
  XNOR U4769 ( .A(n12376), .B(n12678), .Z(n12380) );
  XNOR U4770 ( .A(n12744), .B(n13046), .Z(n12748) );
  XNOR U4771 ( .A(n13112), .B(n13414), .Z(n13116) );
  XNOR U4772 ( .A(n13480), .B(n13782), .Z(n13484) );
  XNOR U4773 ( .A(n13848), .B(n14150), .Z(n13852) );
  XNOR U4774 ( .A(n14216), .B(n14518), .Z(n14220) );
  XNOR U4775 ( .A(n14579), .B(n14886), .Z(n14588) );
  XNOR U4776 ( .A(n15321), .B(n15623), .Z(n15329) );
  XNOR U4777 ( .A(n16057), .B(n16359), .Z(n16061) );
  XNOR U4778 ( .A(n16793), .B(n17095), .Z(n16797) );
  XNOR U4779 ( .A(n17529), .B(n17831), .Z(n17533) );
  XNOR U4780 ( .A(n18265), .B(n18567), .Z(n18269) );
  XNOR U4781 ( .A(n19001), .B(n19303), .Z(n19005) );
  XNOR U4782 ( .A(n19737), .B(n20039), .Z(n19741) );
  XNOR U4783 ( .A(n20473), .B(n20775), .Z(n20477) );
  XNOR U4784 ( .A(n21209), .B(n21511), .Z(n21213) );
  XNOR U4785 ( .A(n21945), .B(n22247), .Z(n21949) );
  XNOR U4786 ( .A(n22681), .B(n22983), .Z(n22685) );
  XNOR U4787 ( .A(n7392), .B(n7710), .Z(n7396) );
  XNOR U4788 ( .A(n6634), .B(n6966), .Z(n6638) );
  XNOR U4789 ( .A(n5869), .B(n6230), .Z(n5874) );
  XNOR U4790 ( .A(n8528), .B(n8822), .Z(n8532) );
  XNOR U4791 ( .A(n9268), .B(n9565), .Z(n9272) );
  XNOR U4792 ( .A(n10020), .B(n10454), .Z(n10024) );
  XNOR U4793 ( .A(n28212), .B(n28502), .Z(n28216) );
  XNOR U4794 ( .A(n27612), .B(n27902), .Z(n27616) );
  XNOR U4795 ( .A(n26988), .B(n27278), .Z(n26992) );
  XNOR U4796 ( .A(n26340), .B(n26630), .Z(n26344) );
  XNOR U4797 ( .A(n25668), .B(n25958), .Z(n25672) );
  XNOR U4798 ( .A(n24972), .B(n25262), .Z(n24976) );
  XNOR U4799 ( .A(n24252), .B(n24542), .Z(n24256) );
  XNOR U4800 ( .A(n23432), .B(n23796), .Z(n23436) );
  XNOR U4801 ( .A(n11293), .B(n10921), .Z(n10923) );
  XNOR U4802 ( .A(n11661), .B(n11290), .Z(n11292) );
  XNOR U4803 ( .A(n11655), .B(n11939), .Z(n11659) );
  XNOR U4804 ( .A(n12023), .B(n12307), .Z(n12027) );
  XNOR U4805 ( .A(n12391), .B(n12675), .Z(n12395) );
  XNOR U4806 ( .A(n12759), .B(n13043), .Z(n12763) );
  XNOR U4807 ( .A(n13127), .B(n13411), .Z(n13131) );
  XNOR U4808 ( .A(n13495), .B(n13779), .Z(n13499) );
  XNOR U4809 ( .A(n13863), .B(n14147), .Z(n13867) );
  XNOR U4810 ( .A(n14231), .B(n14515), .Z(n14235) );
  XNOR U4811 ( .A(n14599), .B(n14883), .Z(n14603) );
  XNOR U4812 ( .A(n14967), .B(n15251), .Z(n14971) );
  XNOR U4813 ( .A(n15335), .B(n15619), .Z(n15339) );
  XNOR U4814 ( .A(n16076), .B(n16356), .Z(n16071) );
  XNOR U4815 ( .A(n16808), .B(n17092), .Z(n16812) );
  XNOR U4816 ( .A(n17544), .B(n17828), .Z(n17548) );
  XNOR U4817 ( .A(n18280), .B(n18564), .Z(n18284) );
  XNOR U4818 ( .A(n19016), .B(n19300), .Z(n19020) );
  XNOR U4819 ( .A(n19752), .B(n20036), .Z(n19756) );
  XNOR U4820 ( .A(n20488), .B(n20772), .Z(n20492) );
  XNOR U4821 ( .A(n21224), .B(n21508), .Z(n21228) );
  XNOR U4822 ( .A(n21960), .B(n22244), .Z(n21964) );
  XNOR U4823 ( .A(n22696), .B(n22980), .Z(n22700) );
  XNOR U4824 ( .A(n7407), .B(n7707), .Z(n7411) );
  XNOR U4825 ( .A(n6649), .B(n6963), .Z(n6653) );
  XNOR U4826 ( .A(n5885), .B(n6227), .Z(n5889) );
  XNOR U4827 ( .A(n8543), .B(n8819), .Z(n8547) );
  XNOR U4828 ( .A(n9283), .B(n9562), .Z(n9287) );
  XNOR U4829 ( .A(n10035), .B(n10448), .Z(n10039) );
  XNOR U4830 ( .A(n10560), .B(n10831), .Z(n10564) );
  XNOR U4831 ( .A(n28803), .B(n29075), .Z(n28807) );
  XNOR U4832 ( .A(n28227), .B(n28499), .Z(n28231) );
  XNOR U4833 ( .A(n27627), .B(n27899), .Z(n27631) );
  XNOR U4834 ( .A(n27003), .B(n27275), .Z(n27007) );
  XNOR U4835 ( .A(n26355), .B(n26627), .Z(n26359) );
  XNOR U4836 ( .A(n25683), .B(n25955), .Z(n25687) );
  XNOR U4837 ( .A(n24987), .B(n25259), .Z(n24991) );
  XNOR U4838 ( .A(n24267), .B(n24539), .Z(n24271) );
  XNOR U4839 ( .A(n23447), .B(n23793), .Z(n23451) );
  XNOR U4840 ( .A(n5125), .B(n5486), .Z(n5130) );
  XNOR U4841 ( .A(n11676), .B(n11305), .Z(n11307) );
  XNOR U4842 ( .A(n11670), .B(n11936), .Z(n11674) );
  XNOR U4843 ( .A(n12038), .B(n12304), .Z(n12042) );
  XNOR U4844 ( .A(n12406), .B(n12672), .Z(n12410) );
  XNOR U4845 ( .A(n12774), .B(n13040), .Z(n12778) );
  XNOR U4846 ( .A(n13142), .B(n13408), .Z(n13146) );
  XNOR U4847 ( .A(n13510), .B(n13776), .Z(n13514) );
  XNOR U4848 ( .A(n13878), .B(n14144), .Z(n13882) );
  XNOR U4849 ( .A(n14246), .B(n14512), .Z(n14250) );
  XNOR U4850 ( .A(n14614), .B(n14880), .Z(n14618) );
  XNOR U4851 ( .A(n14982), .B(n15248), .Z(n14986) );
  XNOR U4852 ( .A(n15350), .B(n15616), .Z(n15354) );
  XNOR U4853 ( .A(n15718), .B(n15984), .Z(n15722) );
  XNOR U4854 ( .A(n16086), .B(n16352), .Z(n16090) );
  XNOR U4855 ( .A(n16454), .B(n16720), .Z(n16458) );
  XNOR U4856 ( .A(n16817), .B(n17088), .Z(n16826) );
  XNOR U4857 ( .A(n17559), .B(n17825), .Z(n17567) );
  XNOR U4858 ( .A(n18295), .B(n18561), .Z(n18299) );
  XNOR U4859 ( .A(n19031), .B(n19297), .Z(n19035) );
  XNOR U4860 ( .A(n19767), .B(n20033), .Z(n19771) );
  XNOR U4861 ( .A(n20503), .B(n20769), .Z(n20507) );
  XNOR U4862 ( .A(n21239), .B(n21505), .Z(n21243) );
  XNOR U4863 ( .A(n21975), .B(n22241), .Z(n21979) );
  XNOR U4864 ( .A(n22711), .B(n22977), .Z(n22715) );
  XNOR U4865 ( .A(n7422), .B(n7704), .Z(n7426) );
  XNOR U4866 ( .A(n6664), .B(n6960), .Z(n6668) );
  XNOR U4867 ( .A(n5900), .B(n6224), .Z(n5904) );
  XNOR U4868 ( .A(n8558), .B(n8816), .Z(n8562) );
  XNOR U4869 ( .A(n9298), .B(n9559), .Z(n9302) );
  XNOR U4870 ( .A(n10050), .B(n10442), .Z(n10054) );
  XNOR U4871 ( .A(n10575), .B(n10828), .Z(n10579) );
  XNOR U4872 ( .A(n10943), .B(n11197), .Z(n10947) );
  XNOR U4873 ( .A(n29898), .B(n30152), .Z(n29902) );
  XNOR U4874 ( .A(n29370), .B(n29624), .Z(n29374) );
  XNOR U4875 ( .A(n28818), .B(n29072), .Z(n28822) );
  XNOR U4876 ( .A(n28242), .B(n28496), .Z(n28246) );
  XNOR U4877 ( .A(n27642), .B(n27896), .Z(n27646) );
  XNOR U4878 ( .A(n27018), .B(n27272), .Z(n27022) );
  XNOR U4879 ( .A(n26370), .B(n26624), .Z(n26374) );
  XNOR U4880 ( .A(n25698), .B(n25952), .Z(n25702) );
  XNOR U4881 ( .A(n25002), .B(n25256), .Z(n25006) );
  XNOR U4882 ( .A(n24282), .B(n24536), .Z(n24286) );
  XNOR U4883 ( .A(n23462), .B(n23790), .Z(n23466) );
  XNOR U4884 ( .A(n7814), .B(n8072), .Z(n7818) );
  XNOR U4885 ( .A(n5141), .B(n5483), .Z(n5145) );
  XNOR U4886 ( .A(n11685), .B(n11933), .Z(n11689) );
  XNOR U4887 ( .A(n12053), .B(n12301), .Z(n12057) );
  XNOR U4888 ( .A(n12421), .B(n12669), .Z(n12425) );
  XNOR U4889 ( .A(n12789), .B(n13037), .Z(n12793) );
  XNOR U4890 ( .A(n13157), .B(n13405), .Z(n13161) );
  XNOR U4891 ( .A(n13525), .B(n13773), .Z(n13529) );
  XNOR U4892 ( .A(n13893), .B(n14141), .Z(n13897) );
  XNOR U4893 ( .A(n14261), .B(n14509), .Z(n14265) );
  XNOR U4894 ( .A(n14629), .B(n14877), .Z(n14633) );
  XNOR U4895 ( .A(n14997), .B(n15245), .Z(n15001) );
  XNOR U4896 ( .A(n15365), .B(n15613), .Z(n15369) );
  XNOR U4897 ( .A(n15733), .B(n15981), .Z(n15737) );
  XNOR U4898 ( .A(n16101), .B(n16349), .Z(n16105) );
  XNOR U4899 ( .A(n16469), .B(n16717), .Z(n16473) );
  XNOR U4900 ( .A(n16837), .B(n17085), .Z(n16841) );
  XNOR U4901 ( .A(n17205), .B(n17453), .Z(n17209) );
  XNOR U4902 ( .A(n17573), .B(n17821), .Z(n17577) );
  XNOR U4903 ( .A(n18314), .B(n18558), .Z(n18309) );
  XNOR U4904 ( .A(n19046), .B(n19294), .Z(n19050) );
  XNOR U4905 ( .A(n19782), .B(n20030), .Z(n19786) );
  XNOR U4906 ( .A(n20518), .B(n20766), .Z(n20522) );
  XNOR U4907 ( .A(n21254), .B(n21502), .Z(n21258) );
  XNOR U4908 ( .A(n21990), .B(n22238), .Z(n21994) );
  XNOR U4909 ( .A(n22726), .B(n22974), .Z(n22730) );
  XNOR U4910 ( .A(n7052), .B(n7331), .Z(n7056) );
  XNOR U4911 ( .A(n4380), .B(n4741), .Z(n4385) );
  XNOR U4912 ( .A(n6297), .B(n6591), .Z(n6301) );
  XNOR U4913 ( .A(n5533), .B(n5851), .Z(n5537) );
  XNOR U4914 ( .A(n8573), .B(n8813), .Z(n8577) );
  XNOR U4915 ( .A(n9313), .B(n9556), .Z(n9317) );
  XNOR U4916 ( .A(n10065), .B(n10436), .Z(n10069) );
  XNOR U4917 ( .A(n10590), .B(n10825), .Z(n10594) );
  XNOR U4918 ( .A(n10958), .B(n11194), .Z(n10962) );
  XNOR U4919 ( .A(n11327), .B(n11563), .Z(n11331) );
  XNOR U4920 ( .A(n12069), .B(n11698), .Z(n11700) );
  XNOR U4921 ( .A(n30417), .B(n30653), .Z(n30421) );
  XNOR U4922 ( .A(n29913), .B(n30149), .Z(n29917) );
  XNOR U4923 ( .A(n29385), .B(n29621), .Z(n29389) );
  XNOR U4924 ( .A(n28833), .B(n29069), .Z(n28837) );
  XNOR U4925 ( .A(n28257), .B(n28493), .Z(n28261) );
  XNOR U4926 ( .A(n27657), .B(n27893), .Z(n27661) );
  XNOR U4927 ( .A(n27033), .B(n27269), .Z(n27037) );
  XNOR U4928 ( .A(n26385), .B(n26621), .Z(n26389) );
  XNOR U4929 ( .A(n25713), .B(n25949), .Z(n25717) );
  XNOR U4930 ( .A(n25017), .B(n25253), .Z(n25021) );
  XNOR U4931 ( .A(n24297), .B(n24533), .Z(n24301) );
  XNOR U4932 ( .A(n23477), .B(n23787), .Z(n23481) );
  XNOR U4933 ( .A(n7829), .B(n8069), .Z(n7833) );
  XNOR U4934 ( .A(n4773), .B(n5110), .Z(n4777) );
  XNOR U4935 ( .A(n12436), .B(n12666), .Z(n12440) );
  XNOR U4936 ( .A(n12804), .B(n13034), .Z(n12808) );
  XNOR U4937 ( .A(n13172), .B(n13402), .Z(n13176) );
  XNOR U4938 ( .A(n13540), .B(n13770), .Z(n13544) );
  XNOR U4939 ( .A(n13908), .B(n14138), .Z(n13912) );
  XNOR U4940 ( .A(n14276), .B(n14506), .Z(n14280) );
  XNOR U4941 ( .A(n14644), .B(n14874), .Z(n14648) );
  XNOR U4942 ( .A(n15012), .B(n15242), .Z(n15016) );
  XNOR U4943 ( .A(n15380), .B(n15610), .Z(n15384) );
  XNOR U4944 ( .A(n15748), .B(n15978), .Z(n15752) );
  XNOR U4945 ( .A(n16116), .B(n16346), .Z(n16120) );
  XNOR U4946 ( .A(n16484), .B(n16714), .Z(n16488) );
  XNOR U4947 ( .A(n16852), .B(n17082), .Z(n16856) );
  XNOR U4948 ( .A(n17220), .B(n17450), .Z(n17224) );
  XNOR U4949 ( .A(n17588), .B(n17818), .Z(n17592) );
  XNOR U4950 ( .A(n17956), .B(n18186), .Z(n17960) );
  XNOR U4951 ( .A(n18324), .B(n18554), .Z(n18328) );
  XNOR U4952 ( .A(n18692), .B(n18922), .Z(n18696) );
  XNOR U4953 ( .A(n19055), .B(n19290), .Z(n19064) );
  XNOR U4954 ( .A(n19797), .B(n20027), .Z(n19805) );
  XNOR U4955 ( .A(n20533), .B(n20763), .Z(n20537) );
  XNOR U4956 ( .A(n21269), .B(n21499), .Z(n21273) );
  XNOR U4957 ( .A(n22005), .B(n22235), .Z(n22009) );
  XNOR U4958 ( .A(n22741), .B(n22971), .Z(n22745) );
  XNOR U4959 ( .A(n7067), .B(n7328), .Z(n7071) );
  XNOR U4960 ( .A(n4014), .B(n4368), .Z(n4018) );
  XNOR U4961 ( .A(n10974), .B(n10603), .Z(n10605) );
  XNOR U4962 ( .A(n6312), .B(n6588), .Z(n6316) );
  XNOR U4963 ( .A(n5548), .B(n5848), .Z(n5552) );
  XNOR U4964 ( .A(n8588), .B(n8810), .Z(n8592) );
  XNOR U4965 ( .A(n9328), .B(n9553), .Z(n9332) );
  XNOR U4966 ( .A(n10080), .B(n10430), .Z(n10084) );
  XNOR U4967 ( .A(n11342), .B(n11560), .Z(n11346) );
  XNOR U4968 ( .A(n12084), .B(n11713), .Z(n11715) );
  XNOR U4969 ( .A(n12452), .B(n12081), .Z(n12083) );
  XNOR U4970 ( .A(n12820), .B(n12449), .Z(n12451) );
  XNOR U4971 ( .A(n13188), .B(n12817), .Z(n12819) );
  XNOR U4972 ( .A(n31368), .B(n31586), .Z(n31372) );
  XNOR U4973 ( .A(n30912), .B(n31130), .Z(n30916) );
  XNOR U4974 ( .A(n30432), .B(n30650), .Z(n30436) );
  XNOR U4975 ( .A(n29928), .B(n30146), .Z(n29932) );
  XNOR U4976 ( .A(n29400), .B(n29618), .Z(n29404) );
  XNOR U4977 ( .A(n28848), .B(n29066), .Z(n28852) );
  XNOR U4978 ( .A(n28272), .B(n28490), .Z(n28276) );
  XNOR U4979 ( .A(n27672), .B(n27890), .Z(n27676) );
  XNOR U4980 ( .A(n27048), .B(n27266), .Z(n27052) );
  XNOR U4981 ( .A(n26400), .B(n26618), .Z(n26404) );
  XNOR U4982 ( .A(n25728), .B(n25946), .Z(n25732) );
  XNOR U4983 ( .A(n25032), .B(n25250), .Z(n25036) );
  XNOR U4984 ( .A(n24312), .B(n24530), .Z(n24316) );
  XNOR U4985 ( .A(n23492), .B(n23784), .Z(n23496) );
  XNOR U4986 ( .A(n7844), .B(n8066), .Z(n7852) );
  XNOR U4987 ( .A(n4788), .B(n5107), .Z(n4792) );
  XNOR U4988 ( .A(n10978), .B(n11190), .Z(n10982) );
  XNOR U4989 ( .A(n13555), .B(n13767), .Z(n13559) );
  XNOR U4990 ( .A(n13923), .B(n14135), .Z(n13927) );
  XNOR U4991 ( .A(n14291), .B(n14503), .Z(n14295) );
  XNOR U4992 ( .A(n14659), .B(n14871), .Z(n14663) );
  XNOR U4993 ( .A(n15027), .B(n15239), .Z(n15031) );
  XNOR U4994 ( .A(n15395), .B(n15607), .Z(n15399) );
  XNOR U4995 ( .A(n15763), .B(n15975), .Z(n15767) );
  XNOR U4996 ( .A(n16131), .B(n16343), .Z(n16135) );
  XNOR U4997 ( .A(n16499), .B(n16711), .Z(n16503) );
  XNOR U4998 ( .A(n16867), .B(n17079), .Z(n16871) );
  XNOR U4999 ( .A(n17235), .B(n17447), .Z(n17239) );
  XNOR U5000 ( .A(n17603), .B(n17815), .Z(n17607) );
  XNOR U5001 ( .A(n17971), .B(n18183), .Z(n17975) );
  XNOR U5002 ( .A(n18339), .B(n18551), .Z(n18343) );
  XNOR U5003 ( .A(n18707), .B(n18919), .Z(n18711) );
  XNOR U5004 ( .A(n19075), .B(n19287), .Z(n19079) );
  XNOR U5005 ( .A(n19443), .B(n19655), .Z(n19447) );
  XNOR U5006 ( .A(n19811), .B(n20023), .Z(n19815) );
  XNOR U5007 ( .A(n20552), .B(n20760), .Z(n20547) );
  XNOR U5008 ( .A(n21284), .B(n21496), .Z(n21288) );
  XNOR U5009 ( .A(n22020), .B(n22232), .Z(n22024) );
  XNOR U5010 ( .A(n22756), .B(n22968), .Z(n22760) );
  XNOR U5011 ( .A(n7082), .B(n7325), .Z(n7086) );
  XNOR U5012 ( .A(n4029), .B(n4365), .Z(n4033) );
  XNOR U5013 ( .A(n3264), .B(n3625), .Z(n3269) );
  XNOR U5014 ( .A(n10989), .B(n10618), .Z(n10620) );
  XNOR U5015 ( .A(n6327), .B(n6585), .Z(n6331) );
  XNOR U5016 ( .A(n5563), .B(n5845), .Z(n5567) );
  XNOR U5017 ( .A(n7858), .B(n8062), .Z(n7862) );
  XNOR U5018 ( .A(n8607), .B(n8807), .Z(n8602) );
  XNOR U5019 ( .A(n9343), .B(n9550), .Z(n9347) );
  XNOR U5020 ( .A(n10095), .B(n10424), .Z(n10099) );
  XNOR U5021 ( .A(n11357), .B(n11557), .Z(n11361) );
  XNOR U5022 ( .A(n12835), .B(n12464), .Z(n12466) );
  XNOR U5023 ( .A(n13203), .B(n12832), .Z(n12834) );
  XNOR U5024 ( .A(n13571), .B(n13200), .Z(n13202) );
  XNOR U5025 ( .A(n13939), .B(n13568), .Z(n13570) );
  XNOR U5026 ( .A(n14307), .B(n13936), .Z(n13938) );
  XNOR U5027 ( .A(n31986), .B(n32178), .Z(n31990) );
  XNOR U5028 ( .A(n31383), .B(n31583), .Z(n31387) );
  XNOR U5029 ( .A(n30927), .B(n31127), .Z(n30931) );
  XNOR U5030 ( .A(n30447), .B(n30647), .Z(n30451) );
  XNOR U5031 ( .A(n29943), .B(n30143), .Z(n29947) );
  XNOR U5032 ( .A(n29415), .B(n29615), .Z(n29419) );
  XNOR U5033 ( .A(n28863), .B(n29063), .Z(n28867) );
  XNOR U5034 ( .A(n28287), .B(n28487), .Z(n28291) );
  XNOR U5035 ( .A(n27687), .B(n27887), .Z(n27691) );
  XNOR U5036 ( .A(n27063), .B(n27263), .Z(n27067) );
  XNOR U5037 ( .A(n26415), .B(n26615), .Z(n26419) );
  XNOR U5038 ( .A(n25743), .B(n25943), .Z(n25747) );
  XNOR U5039 ( .A(n25047), .B(n25247), .Z(n25051) );
  XNOR U5040 ( .A(n24327), .B(n24527), .Z(n24331) );
  XNOR U5041 ( .A(n23507), .B(n23781), .Z(n23511) );
  XNOR U5042 ( .A(n7111), .B(n7318), .Z(n7115) );
  XNOR U5043 ( .A(n6351), .B(n6579), .Z(n6355) );
  XNOR U5044 ( .A(n4803), .B(n5104), .Z(n4807) );
  XNOR U5045 ( .A(n10993), .B(n11187), .Z(n10997) );
  XNOR U5046 ( .A(n12472), .B(n12101), .Z(n12103) );
  XNOR U5047 ( .A(n12840), .B(n12469), .Z(n12471) );
  XNOR U5048 ( .A(n14674), .B(n14868), .Z(n14678) );
  XNOR U5049 ( .A(n15042), .B(n15236), .Z(n15046) );
  XNOR U5050 ( .A(n15410), .B(n15604), .Z(n15414) );
  XNOR U5051 ( .A(n15778), .B(n15972), .Z(n15782) );
  XNOR U5052 ( .A(n16146), .B(n16340), .Z(n16150) );
  XNOR U5053 ( .A(n16514), .B(n16708), .Z(n16518) );
  XNOR U5054 ( .A(n16882), .B(n17076), .Z(n16886) );
  XNOR U5055 ( .A(n17250), .B(n17444), .Z(n17254) );
  XNOR U5056 ( .A(n17618), .B(n17812), .Z(n17622) );
  XNOR U5057 ( .A(n17986), .B(n18180), .Z(n17990) );
  XNOR U5058 ( .A(n18354), .B(n18548), .Z(n18358) );
  XNOR U5059 ( .A(n18722), .B(n18916), .Z(n18726) );
  XNOR U5060 ( .A(n19090), .B(n19284), .Z(n19094) );
  XNOR U5061 ( .A(n19458), .B(n19652), .Z(n19462) );
  XNOR U5062 ( .A(n19826), .B(n20020), .Z(n19830) );
  XNOR U5063 ( .A(n20194), .B(n20388), .Z(n20198) );
  XNOR U5064 ( .A(n20562), .B(n20756), .Z(n20566) );
  XNOR U5065 ( .A(n20930), .B(n21124), .Z(n20934) );
  XNOR U5066 ( .A(n21293), .B(n21492), .Z(n21302) );
  XNOR U5067 ( .A(n22035), .B(n22229), .Z(n22043) );
  XNOR U5068 ( .A(n22771), .B(n22965), .Z(n22775) );
  XNOR U5069 ( .A(n6723), .B(n6949), .Z(n6718) );
  XNOR U5070 ( .A(n4044), .B(n4362), .Z(n4048) );
  XNOR U5071 ( .A(n3280), .B(n3622), .Z(n3284) );
  XNOR U5072 ( .A(n11004), .B(n10633), .Z(n10635) );
  XNOR U5073 ( .A(n11735), .B(n11923), .Z(n11739) );
  XNOR U5074 ( .A(n5960), .B(n6212), .Z(n5968) );
  XNOR U5075 ( .A(n5196), .B(n5472), .Z(n5200) );
  XNOR U5076 ( .A(n2519), .B(n2881), .Z(n2524) );
  XNOR U5077 ( .A(n7873), .B(n8059), .Z(n7881) );
  XNOR U5078 ( .A(n8617), .B(n8803), .Z(n8621) );
  XNOR U5079 ( .A(n9360), .B(n9546), .Z(n9361) );
  XNOR U5080 ( .A(n10110), .B(n10418), .Z(n10118) );
  XNOR U5081 ( .A(n11372), .B(n11554), .Z(n11376) );
  XNOR U5082 ( .A(n12850), .B(n12479), .Z(n12481) );
  XNOR U5083 ( .A(n13954), .B(n13583), .Z(n13585) );
  XNOR U5084 ( .A(n14322), .B(n13951), .Z(n13953) );
  XNOR U5085 ( .A(n14690), .B(n14319), .Z(n14321) );
  XNOR U5086 ( .A(n15058), .B(n14687), .Z(n14689) );
  XNOR U5087 ( .A(n15426), .B(n15055), .Z(n15057) );
  XNOR U5088 ( .A(n32764), .B(n32938), .Z(n32768) );
  XNOR U5089 ( .A(n32393), .B(n32570), .Z(n32397) );
  XNOR U5090 ( .A(n32001), .B(n32175), .Z(n32005) );
  XNOR U5091 ( .A(n31398), .B(n31580), .Z(n31402) );
  XNOR U5092 ( .A(n30942), .B(n31124), .Z(n30946) );
  XNOR U5093 ( .A(n30462), .B(n30644), .Z(n30466) );
  XNOR U5094 ( .A(n29958), .B(n30140), .Z(n29962) );
  XNOR U5095 ( .A(n29430), .B(n29612), .Z(n29434) );
  XNOR U5096 ( .A(n28878), .B(n29060), .Z(n28882) );
  XNOR U5097 ( .A(n28302), .B(n28484), .Z(n28306) );
  XNOR U5098 ( .A(n27702), .B(n27884), .Z(n27706) );
  XNOR U5099 ( .A(n27078), .B(n27260), .Z(n27082) );
  XNOR U5100 ( .A(n26430), .B(n26612), .Z(n26434) );
  XNOR U5101 ( .A(n25758), .B(n25940), .Z(n25762) );
  XNOR U5102 ( .A(n25062), .B(n25244), .Z(n25066) );
  XNOR U5103 ( .A(n24342), .B(n24524), .Z(n24346) );
  XNOR U5104 ( .A(n23522), .B(n23778), .Z(n23526) );
  XNOR U5105 ( .A(n6752), .B(n6942), .Z(n6747) );
  XNOR U5106 ( .A(n5984), .B(n6206), .Z(n5988) );
  XNOR U5107 ( .A(n4436), .B(n4730), .Z(n4440) );
  XNOR U5108 ( .A(n6008), .B(n6200), .Z(n6012) );
  XNOR U5109 ( .A(n11008), .B(n11184), .Z(n11012) );
  XNOR U5110 ( .A(n12487), .B(n12116), .Z(n12118) );
  XNOR U5111 ( .A(n13591), .B(n13220), .Z(n13222) );
  XNOR U5112 ( .A(n13959), .B(n13588), .Z(n13590) );
  XNOR U5113 ( .A(n15793), .B(n15969), .Z(n15797) );
  XNOR U5114 ( .A(n16161), .B(n16337), .Z(n16165) );
  XNOR U5115 ( .A(n16529), .B(n16705), .Z(n16533) );
  XNOR U5116 ( .A(n16897), .B(n17073), .Z(n16901) );
  XNOR U5117 ( .A(n17265), .B(n17441), .Z(n17269) );
  XNOR U5118 ( .A(n17633), .B(n17809), .Z(n17637) );
  XNOR U5119 ( .A(n18001), .B(n18177), .Z(n18005) );
  XNOR U5120 ( .A(n18369), .B(n18545), .Z(n18373) );
  XNOR U5121 ( .A(n18737), .B(n18913), .Z(n18741) );
  XNOR U5122 ( .A(n19105), .B(n19281), .Z(n19109) );
  XNOR U5123 ( .A(n19473), .B(n19649), .Z(n19477) );
  XNOR U5124 ( .A(n19841), .B(n20017), .Z(n19845) );
  XNOR U5125 ( .A(n20209), .B(n20385), .Z(n20213) );
  XNOR U5126 ( .A(n20577), .B(n20753), .Z(n20581) );
  XNOR U5127 ( .A(n20945), .B(n21121), .Z(n20949) );
  XNOR U5128 ( .A(n21313), .B(n21489), .Z(n21317) );
  XNOR U5129 ( .A(n21681), .B(n21857), .Z(n21685) );
  XNOR U5130 ( .A(n22049), .B(n22225), .Z(n22053) );
  XNOR U5131 ( .A(n22790), .B(n22962), .Z(n22785) );
  XNOR U5132 ( .A(n5225), .B(n5465), .Z(n5229) );
  XNOR U5133 ( .A(n3677), .B(n3989), .Z(n3681) );
  XNOR U5134 ( .A(n2913), .B(n3249), .Z(n2917) );
  XNOR U5135 ( .A(n5249), .B(n5459), .Z(n5253) );
  XNOR U5136 ( .A(n6395), .B(n6569), .Z(n6403) );
  XNOR U5137 ( .A(n11019), .B(n10648), .Z(n10650) );
  XNOR U5138 ( .A(n11750), .B(n11920), .Z(n11754) );
  XNOR U5139 ( .A(n12854), .B(n13024), .Z(n12858) );
  XNOR U5140 ( .A(n5215), .B(n5469), .Z(n5210) );
  XNOR U5141 ( .A(n2152), .B(n2507), .Z(n2156) );
  XNOR U5142 ( .A(n7140), .B(n7311), .Z(n7144) );
  XNOR U5143 ( .A(n7887), .B(n8055), .Z(n7891) );
  XNOR U5144 ( .A(n8636), .B(n8800), .Z(n8631) );
  XNOR U5145 ( .A(n9372), .B(n9543), .Z(n9376) );
  XNOR U5146 ( .A(n10124), .B(n10413), .Z(n10128) );
  XNOR U5147 ( .A(n11387), .B(n11551), .Z(n11391) );
  XNOR U5148 ( .A(n12865), .B(n12494), .Z(n12496) );
  XNOR U5149 ( .A(n13969), .B(n13598), .Z(n13600) );
  XNOR U5150 ( .A(n15073), .B(n14702), .Z(n14704) );
  XNOR U5151 ( .A(n15441), .B(n15070), .Z(n15072) );
  XNOR U5152 ( .A(n15809), .B(n15438), .Z(n15440) );
  XNOR U5153 ( .A(n16177), .B(n15806), .Z(n15808) );
  XNOR U5154 ( .A(n16545), .B(n16174), .Z(n16176) );
  XNOR U5155 ( .A(n33126), .B(n33282), .Z(n33130) );
  XNOR U5156 ( .A(n32779), .B(n32935), .Z(n32783) );
  XNOR U5157 ( .A(n32408), .B(n32567), .Z(n32412) );
  XNOR U5158 ( .A(n32016), .B(n32172), .Z(n32020) );
  XNOR U5159 ( .A(n31413), .B(n31577), .Z(n31417) );
  XNOR U5160 ( .A(n30957), .B(n31121), .Z(n30961) );
  XNOR U5161 ( .A(n30477), .B(n30641), .Z(n30481) );
  XNOR U5162 ( .A(n29973), .B(n30137), .Z(n29977) );
  XNOR U5163 ( .A(n29445), .B(n29609), .Z(n29449) );
  XNOR U5164 ( .A(n28893), .B(n29057), .Z(n28897) );
  XNOR U5165 ( .A(n28317), .B(n28481), .Z(n28321) );
  XNOR U5166 ( .A(n27717), .B(n27881), .Z(n27721) );
  XNOR U5167 ( .A(n27093), .B(n27257), .Z(n27097) );
  XNOR U5168 ( .A(n26445), .B(n26609), .Z(n26449) );
  XNOR U5169 ( .A(n25773), .B(n25937), .Z(n25777) );
  XNOR U5170 ( .A(n25077), .B(n25241), .Z(n25081) );
  XNOR U5171 ( .A(n24357), .B(n24521), .Z(n24361) );
  XNOR U5172 ( .A(n23531), .B(n23775), .Z(n23540) );
  XNOR U5173 ( .A(n5278), .B(n5452), .Z(n5282) );
  XNOR U5174 ( .A(n5621), .B(n5833), .Z(n5616) );
  XNOR U5175 ( .A(n4088), .B(n4352), .Z(n4092) );
  XNOR U5176 ( .A(n4451), .B(n4727), .Z(n4459) );
  XNOR U5177 ( .A(n11023), .B(n11181), .Z(n11027) );
  XNOR U5178 ( .A(n12502), .B(n12131), .Z(n12133) );
  XNOR U5179 ( .A(n13606), .B(n13235), .Z(n13237) );
  XNOR U5180 ( .A(n14710), .B(n14339), .Z(n14341) );
  XNOR U5181 ( .A(n15078), .B(n14707), .Z(n14709) );
  XNOR U5182 ( .A(n16912), .B(n17070), .Z(n16916) );
  XNOR U5183 ( .A(n17280), .B(n17438), .Z(n17284) );
  XNOR U5184 ( .A(n17648), .B(n17806), .Z(n17652) );
  XNOR U5185 ( .A(n18016), .B(n18174), .Z(n18020) );
  XNOR U5186 ( .A(n18384), .B(n18542), .Z(n18388) );
  XNOR U5187 ( .A(n18752), .B(n18910), .Z(n18756) );
  XNOR U5188 ( .A(n19120), .B(n19278), .Z(n19124) );
  XNOR U5189 ( .A(n19488), .B(n19646), .Z(n19492) );
  XNOR U5190 ( .A(n19856), .B(n20014), .Z(n19860) );
  XNOR U5191 ( .A(n20224), .B(n20382), .Z(n20228) );
  XNOR U5192 ( .A(n20592), .B(n20750), .Z(n20596) );
  XNOR U5193 ( .A(n20960), .B(n21118), .Z(n20964) );
  XNOR U5194 ( .A(n21328), .B(n21486), .Z(n21332) );
  XNOR U5195 ( .A(n21696), .B(n21854), .Z(n21700) );
  XNOR U5196 ( .A(n22064), .B(n22222), .Z(n22068) );
  XNOR U5197 ( .A(n22432), .B(n22590), .Z(n22436) );
  XNOR U5198 ( .A(n22800), .B(n22958), .Z(n22804) );
  XNOR U5199 ( .A(n4857), .B(n5092), .Z(n4865) );
  XNOR U5200 ( .A(n3692), .B(n3986), .Z(n3696) );
  XNOR U5201 ( .A(n2928), .B(n3246), .Z(n2932) );
  XNOR U5202 ( .A(n5650), .B(n5826), .Z(n5645) );
  XNOR U5203 ( .A(n4499), .B(n4715), .Z(n4503) );
  XNOR U5204 ( .A(n5665), .B(n5821), .Z(n5669) );
  XNOR U5205 ( .A(n11034), .B(n10663), .Z(n10665) );
  XNOR U5206 ( .A(n11765), .B(n11917), .Z(n11769) );
  XNOR U5207 ( .A(n12869), .B(n13021), .Z(n12873) );
  XNOR U5208 ( .A(n13973), .B(n14125), .Z(n13977) );
  XNOR U5209 ( .A(n2167), .B(n2504), .Z(n2171) );
  XNOR U5210 ( .A(n1402), .B(n1763), .Z(n1407) );
  XNOR U5211 ( .A(n4886), .B(n5085), .Z(n4894) );
  XNOR U5212 ( .A(n6414), .B(n6564), .Z(n6418) );
  XNOR U5213 ( .A(n7157), .B(n7307), .Z(n7158) );
  XNOR U5214 ( .A(n7902), .B(n8052), .Z(n7910) );
  XNOR U5215 ( .A(n8646), .B(n8796), .Z(n8650) );
  XNOR U5216 ( .A(n9389), .B(n9539), .Z(n9390) );
  XNOR U5217 ( .A(n10139), .B(n10407), .Z(n10147) );
  XNOR U5218 ( .A(n11402), .B(n11548), .Z(n11406) );
  XNOR U5219 ( .A(n12880), .B(n12509), .Z(n12511) );
  XNOR U5220 ( .A(n13984), .B(n13613), .Z(n13615) );
  XNOR U5221 ( .A(n15088), .B(n14717), .Z(n14719) );
  XNOR U5222 ( .A(n16192), .B(n15821), .Z(n15823) );
  XNOR U5223 ( .A(n16560), .B(n16189), .Z(n16191) );
  XNOR U5224 ( .A(n16928), .B(n16557), .Z(n16559) );
  XNOR U5225 ( .A(n17296), .B(n16925), .Z(n16927) );
  XNOR U5226 ( .A(n17664), .B(n17293), .Z(n17295) );
  XNOR U5227 ( .A(n33760), .B(n33898), .Z(n33764) );
  XNOR U5228 ( .A(n33461), .B(n33602), .Z(n33465) );
  XNOR U5229 ( .A(n33141), .B(n33279), .Z(n33145) );
  XNOR U5230 ( .A(n32794), .B(n32932), .Z(n32798) );
  XNOR U5231 ( .A(n32423), .B(n32564), .Z(n32427) );
  XNOR U5232 ( .A(n32031), .B(n32169), .Z(n32035) );
  XNOR U5233 ( .A(n31428), .B(n31574), .Z(n31432) );
  XNOR U5234 ( .A(n30972), .B(n31118), .Z(n30976) );
  XNOR U5235 ( .A(n30492), .B(n30638), .Z(n30496) );
  XNOR U5236 ( .A(n29988), .B(n30134), .Z(n29992) );
  XNOR U5237 ( .A(n29460), .B(n29606), .Z(n29464) );
  XNOR U5238 ( .A(n28908), .B(n29054), .Z(n28912) );
  XNOR U5239 ( .A(n28332), .B(n28478), .Z(n28336) );
  XNOR U5240 ( .A(n27732), .B(n27878), .Z(n27736) );
  XNOR U5241 ( .A(n27108), .B(n27254), .Z(n27112) );
  XNOR U5242 ( .A(n26460), .B(n26606), .Z(n26464) );
  XNOR U5243 ( .A(n25788), .B(n25934), .Z(n25792) );
  XNOR U5244 ( .A(n25092), .B(n25238), .Z(n25096) );
  XNOR U5245 ( .A(n24372), .B(n24518), .Z(n24376) );
  XNOR U5246 ( .A(n23551), .B(n23772), .Z(n23555) );
  XNOR U5247 ( .A(n4528), .B(n4708), .Z(n4532) );
  XNOR U5248 ( .A(n3721), .B(n3979), .Z(n3725) );
  XNOR U5249 ( .A(n2957), .B(n3239), .Z(n2961) );
  XNOR U5250 ( .A(n11038), .B(n11178), .Z(n11042) );
  XNOR U5251 ( .A(n12517), .B(n12146), .Z(n12148) );
  XNOR U5252 ( .A(n13621), .B(n13250), .Z(n13252) );
  XNOR U5253 ( .A(n14725), .B(n14354), .Z(n14356) );
  XNOR U5254 ( .A(n15829), .B(n15458), .Z(n15460) );
  XNOR U5255 ( .A(n16197), .B(n15826), .Z(n15828) );
  XNOR U5256 ( .A(n18031), .B(n18171), .Z(n18035) );
  XNOR U5257 ( .A(n18399), .B(n18539), .Z(n18403) );
  XNOR U5258 ( .A(n18767), .B(n18907), .Z(n18771) );
  XNOR U5259 ( .A(n19135), .B(n19275), .Z(n19139) );
  XNOR U5260 ( .A(n19503), .B(n19643), .Z(n19507) );
  XNOR U5261 ( .A(n19871), .B(n20011), .Z(n19875) );
  XNOR U5262 ( .A(n20239), .B(n20379), .Z(n20243) );
  XNOR U5263 ( .A(n20607), .B(n20747), .Z(n20611) );
  XNOR U5264 ( .A(n20975), .B(n21115), .Z(n20979) );
  XNOR U5265 ( .A(n21343), .B(n21483), .Z(n21347) );
  XNOR U5266 ( .A(n21711), .B(n21851), .Z(n21715) );
  XNOR U5267 ( .A(n22079), .B(n22219), .Z(n22083) );
  XNOR U5268 ( .A(n22447), .B(n22587), .Z(n22451) );
  XNOR U5269 ( .A(n22815), .B(n22955), .Z(n22819) );
  XNOR U5270 ( .A(n4915), .B(n5078), .Z(n4923) );
  XNOR U5271 ( .A(n4112), .B(n4348), .Z(n4107) );
  XNOR U5272 ( .A(n3329), .B(n3613), .Z(n3324) );
  XNOR U5273 ( .A(n2560), .B(n2873), .Z(n2564) );
  XNOR U5274 ( .A(n3750), .B(n3972), .Z(n3754) );
  XNOR U5275 ( .A(n2986), .B(n3232), .Z(n2990) );
  XNOR U5276 ( .A(n4557), .B(n4701), .Z(n4561) );
  XNOR U5277 ( .A(n11049), .B(n10678), .Z(n10680) );
  XNOR U5278 ( .A(n11780), .B(n11914), .Z(n11784) );
  XNOR U5279 ( .A(n12884), .B(n13018), .Z(n12888) );
  XNOR U5280 ( .A(n13988), .B(n14122), .Z(n13992) );
  XNOR U5281 ( .A(n15092), .B(n15226), .Z(n15096) );
  XNOR U5282 ( .A(n1800), .B(n2130), .Z(n1804) );
  XNOR U5283 ( .A(n1036), .B(n1390), .Z(n1040) );
  XNOR U5284 ( .A(n4141), .B(n4341), .Z(n4136) );
  XNOR U5285 ( .A(n5684), .B(n5816), .Z(n5688) );
  XNOR U5286 ( .A(n6433), .B(n6561), .Z(n6428) );
  XNOR U5287 ( .A(n7169), .B(n7304), .Z(n7173) );
  XNOR U5288 ( .A(n7916), .B(n8048), .Z(n7920) );
  XNOR U5289 ( .A(n8665), .B(n8793), .Z(n8660) );
  XNOR U5290 ( .A(n9401), .B(n9536), .Z(n9405) );
  XNOR U5291 ( .A(n10153), .B(n10402), .Z(n10157) );
  XNOR U5292 ( .A(n11417), .B(n11545), .Z(n11421) );
  XNOR U5293 ( .A(n12895), .B(n12524), .Z(n12526) );
  XNOR U5294 ( .A(n13999), .B(n13628), .Z(n13630) );
  XNOR U5295 ( .A(n15103), .B(n14732), .Z(n14734) );
  XNOR U5296 ( .A(n16207), .B(n15836), .Z(n15838) );
  XNOR U5297 ( .A(n17311), .B(n16940), .Z(n16942) );
  XNOR U5298 ( .A(n17679), .B(n17308), .Z(n17310) );
  XNOR U5299 ( .A(n18047), .B(n17676), .Z(n17678) );
  XNOR U5300 ( .A(n18415), .B(n18044), .Z(n18046) );
  XNOR U5301 ( .A(n18783), .B(n18412), .Z(n18414) );
  XNOR U5302 ( .A(n34050), .B(n34170), .Z(n34054) );
  XNOR U5303 ( .A(n33775), .B(n33895), .Z(n33779) );
  XNOR U5304 ( .A(n33476), .B(n33599), .Z(n33480) );
  XNOR U5305 ( .A(n33156), .B(n33276), .Z(n33160) );
  XNOR U5306 ( .A(n32809), .B(n32929), .Z(n32813) );
  XNOR U5307 ( .A(n32438), .B(n32561), .Z(n32442) );
  XNOR U5308 ( .A(n32046), .B(n32166), .Z(n32050) );
  XNOR U5309 ( .A(n31443), .B(n31571), .Z(n31447) );
  XNOR U5310 ( .A(n30987), .B(n31115), .Z(n30991) );
  XNOR U5311 ( .A(n30507), .B(n30635), .Z(n30511) );
  XNOR U5312 ( .A(n30003), .B(n30131), .Z(n30007) );
  XNOR U5313 ( .A(n29475), .B(n29603), .Z(n29479) );
  XNOR U5314 ( .A(n28923), .B(n29051), .Z(n28927) );
  XNOR U5315 ( .A(n28347), .B(n28475), .Z(n28351) );
  XNOR U5316 ( .A(n27747), .B(n27875), .Z(n27751) );
  XNOR U5317 ( .A(n27123), .B(n27251), .Z(n27127) );
  XNOR U5318 ( .A(n26475), .B(n26603), .Z(n26479) );
  XNOR U5319 ( .A(n25803), .B(n25931), .Z(n25807) );
  XNOR U5320 ( .A(n25107), .B(n25235), .Z(n25111) );
  XNOR U5321 ( .A(n24387), .B(n24515), .Z(n24391) );
  XNOR U5322 ( .A(n23566), .B(n23769), .Z(n23570) );
  XNOR U5323 ( .A(n3779), .B(n3965), .Z(n3783) );
  XNOR U5324 ( .A(n3015), .B(n3225), .Z(n3019) );
  XNOR U5325 ( .A(n2972), .B(n3236), .Z(n2980) );
  XNOR U5326 ( .A(n2206), .B(n2495), .Z(n2210) );
  XNOR U5327 ( .A(n5317), .B(n5443), .Z(n5321) );
  XNOR U5328 ( .A(n11053), .B(n11175), .Z(n11057) );
  XNOR U5329 ( .A(n12532), .B(n12161), .Z(n12163) );
  XNOR U5330 ( .A(n13636), .B(n13265), .Z(n13267) );
  XNOR U5331 ( .A(n14740), .B(n14369), .Z(n14371) );
  XNOR U5332 ( .A(n15844), .B(n15473), .Z(n15475) );
  XNOR U5333 ( .A(n16948), .B(n16577), .Z(n16579) );
  XNOR U5334 ( .A(n17316), .B(n16945), .Z(n16947) );
  XNOR U5335 ( .A(n19150), .B(n19272), .Z(n19154) );
  XNOR U5336 ( .A(n19518), .B(n19640), .Z(n19522) );
  XNOR U5337 ( .A(n19886), .B(n20008), .Z(n19890) );
  XNOR U5338 ( .A(n20254), .B(n20376), .Z(n20258) );
  XNOR U5339 ( .A(n20622), .B(n20744), .Z(n20626) );
  XNOR U5340 ( .A(n20990), .B(n21112), .Z(n20994) );
  XNOR U5341 ( .A(n21358), .B(n21480), .Z(n21362) );
  XNOR U5342 ( .A(n21726), .B(n21848), .Z(n21730) );
  XNOR U5343 ( .A(n22094), .B(n22216), .Z(n22098) );
  XNOR U5344 ( .A(n22462), .B(n22584), .Z(n22466) );
  XNOR U5345 ( .A(n22830), .B(n22952), .Z(n22834) );
  XNOR U5346 ( .A(n4170), .B(n4334), .Z(n4165) );
  XNOR U5347 ( .A(n1447), .B(n1753), .Z(n1451) );
  XNOR U5348 ( .A(n2196), .B(n2499), .Z(n2191) );
  XNOR U5349 ( .A(n3001), .B(n3229), .Z(n3009) );
  XNOR U5350 ( .A(n2235), .B(n2488), .Z(n2239) );
  XNOR U5351 ( .A(n3808), .B(n3958), .Z(n3812) );
  XNOR U5352 ( .A(n3044), .B(n3218), .Z(n3048) );
  XNOR U5353 ( .A(n11064), .B(n10693), .Z(n10695) );
  XNOR U5354 ( .A(n11795), .B(n11911), .Z(n11799) );
  XNOR U5355 ( .A(n12899), .B(n13015), .Z(n12903) );
  XNOR U5356 ( .A(n14003), .B(n14119), .Z(n14007) );
  XNOR U5357 ( .A(n15107), .B(n15223), .Z(n15111) );
  XNOR U5358 ( .A(n16211), .B(n16327), .Z(n16215) );
  XNOR U5359 ( .A(n1433), .B(n1757), .Z(n1441) );
  XNOR U5360 ( .A(n669), .B(n1017), .Z(n673) );
  XNOR U5361 ( .A(n1476), .B(n1746), .Z(n1480) );
  XNOR U5362 ( .A(n4199), .B(n4327), .Z(n4194) );
  XNOR U5363 ( .A(n6443), .B(n6557), .Z(n6447) );
  XNOR U5364 ( .A(n7186), .B(n7300), .Z(n7187) );
  XNOR U5365 ( .A(n7931), .B(n8045), .Z(n7939) );
  XNOR U5366 ( .A(n8675), .B(n8789), .Z(n8679) );
  XNOR U5367 ( .A(n9418), .B(n9532), .Z(n9419) );
  XNOR U5368 ( .A(n10168), .B(n10396), .Z(n10176) );
  XNOR U5369 ( .A(n11432), .B(n11542), .Z(n11436) );
  XNOR U5370 ( .A(n12910), .B(n12539), .Z(n12541) );
  XNOR U5371 ( .A(n14014), .B(n13643), .Z(n13645) );
  XNOR U5372 ( .A(n15118), .B(n14747), .Z(n14749) );
  XNOR U5373 ( .A(n16222), .B(n15851), .Z(n15853) );
  XNOR U5374 ( .A(n17326), .B(n16955), .Z(n16957) );
  XNOR U5375 ( .A(n18430), .B(n18059), .Z(n18061) );
  XNOR U5376 ( .A(n18798), .B(n18427), .Z(n18429) );
  XNOR U5377 ( .A(n19166), .B(n18795), .Z(n18797) );
  XNOR U5378 ( .A(n19534), .B(n19163), .Z(n19165) );
  XNOR U5379 ( .A(n19902), .B(n19531), .Z(n19533) );
  XNOR U5380 ( .A(n34540), .B(n34642), .Z(n34544) );
  XNOR U5381 ( .A(n34313), .B(n34418), .Z(n34317) );
  XNOR U5382 ( .A(n34065), .B(n34167), .Z(n34069) );
  XNOR U5383 ( .A(n33790), .B(n33892), .Z(n33794) );
  XNOR U5384 ( .A(n33491), .B(n33596), .Z(n33495) );
  XNOR U5385 ( .A(n33171), .B(n33273), .Z(n33175) );
  XNOR U5386 ( .A(n32824), .B(n32926), .Z(n32828) );
  XNOR U5387 ( .A(n32453), .B(n32558), .Z(n32457) );
  XNOR U5388 ( .A(n32061), .B(n32163), .Z(n32065) );
  XNOR U5389 ( .A(n31458), .B(n31568), .Z(n31462) );
  XNOR U5390 ( .A(n31002), .B(n31112), .Z(n31006) );
  XNOR U5391 ( .A(n30522), .B(n30632), .Z(n30526) );
  XNOR U5392 ( .A(n30018), .B(n30128), .Z(n30022) );
  XNOR U5393 ( .A(n29490), .B(n29600), .Z(n29494) );
  XNOR U5394 ( .A(n28938), .B(n29048), .Z(n28942) );
  XNOR U5395 ( .A(n28362), .B(n28472), .Z(n28366) );
  XNOR U5396 ( .A(n27762), .B(n27872), .Z(n27766) );
  XNOR U5397 ( .A(n27138), .B(n27248), .Z(n27142) );
  XNOR U5398 ( .A(n26490), .B(n26600), .Z(n26494) );
  XNOR U5399 ( .A(n25818), .B(n25928), .Z(n25822) );
  XNOR U5400 ( .A(n25122), .B(n25232), .Z(n25126) );
  XNOR U5401 ( .A(n24402), .B(n24512), .Z(n24406) );
  XNOR U5402 ( .A(n23581), .B(n23766), .Z(n23585) );
  XNOR U5403 ( .A(n3837), .B(n3951), .Z(n3841) );
  XNOR U5404 ( .A(n3073), .B(n3211), .Z(n3077) );
  XNOR U5405 ( .A(n3030), .B(n3222), .Z(n3038) );
  XNOR U5406 ( .A(n2264), .B(n2481), .Z(n2268) );
  XNOR U5407 ( .A(n2225), .B(n2492), .Z(n2220) );
  XNOR U5408 ( .A(n4586), .B(n4694), .Z(n4590) );
  XNOR U5409 ( .A(n6076), .B(n6184), .Z(n6084) );
  XNOR U5410 ( .A(n11068), .B(n11172), .Z(n11072) );
  XNOR U5411 ( .A(n12547), .B(n12176), .Z(n12178) );
  XNOR U5412 ( .A(n13651), .B(n13280), .Z(n13282) );
  XNOR U5413 ( .A(n14755), .B(n14384), .Z(n14386) );
  XNOR U5414 ( .A(n15859), .B(n15488), .Z(n15490) );
  XNOR U5415 ( .A(n16963), .B(n16592), .Z(n16594) );
  XNOR U5416 ( .A(n18067), .B(n17696), .Z(n17698) );
  XNOR U5417 ( .A(n18435), .B(n18064), .Z(n18066) );
  XNOR U5418 ( .A(n20269), .B(n20373), .Z(n20273) );
  XNOR U5419 ( .A(n20637), .B(n20741), .Z(n20641) );
  XNOR U5420 ( .A(n21005), .B(n21109), .Z(n21009) );
  XNOR U5421 ( .A(n21373), .B(n21477), .Z(n21377) );
  XNOR U5422 ( .A(n21741), .B(n21845), .Z(n21745) );
  XNOR U5423 ( .A(n22109), .B(n22213), .Z(n22113) );
  XNOR U5424 ( .A(n22477), .B(n22581), .Z(n22481) );
  XNOR U5425 ( .A(n22845), .B(n22949), .Z(n22849) );
  XNOR U5426 ( .A(n1505), .B(n1739), .Z(n1509) );
  XNOR U5427 ( .A(n1462), .B(n1750), .Z(n1470) );
  XNOR U5428 ( .A(n698), .B(n1010), .Z(n702) );
  XNOR U5429 ( .A(n2254), .B(n2485), .Z(n2249) );
  XNOR U5430 ( .A(n3059), .B(n3215), .Z(n3067) );
  XNOR U5431 ( .A(n2293), .B(n2474), .Z(n2297) );
  XNOR U5432 ( .A(n5711), .B(n5810), .Z(n5712) );
  XNOR U5433 ( .A(n11079), .B(n10708), .Z(n10710) );
  XNOR U5434 ( .A(n11810), .B(n11908), .Z(n11814) );
  XNOR U5435 ( .A(n12914), .B(n13012), .Z(n12918) );
  XNOR U5436 ( .A(n14018), .B(n14116), .Z(n14022) );
  XNOR U5437 ( .A(n15122), .B(n15220), .Z(n15126) );
  XNOR U5438 ( .A(n16226), .B(n16324), .Z(n16230) );
  XNOR U5439 ( .A(n17330), .B(n17428), .Z(n17334) );
  XNOR U5440 ( .A(n688), .B(n1014), .Z(n683) );
  XNOR U5441 ( .A(n1491), .B(n1743), .Z(n1499) );
  XNOR U5442 ( .A(n727), .B(n1003), .Z(n731) );
  XNOR U5443 ( .A(n1534), .B(n1732), .Z(n1538) );
  XNOR U5444 ( .A(n7198), .B(n7297), .Z(n7202) );
  XNOR U5445 ( .A(n7945), .B(n8041), .Z(n7949) );
  XNOR U5446 ( .A(n8694), .B(n8786), .Z(n8689) );
  XNOR U5447 ( .A(n9430), .B(n9529), .Z(n9434) );
  XNOR U5448 ( .A(n10182), .B(n10391), .Z(n10186) );
  XNOR U5449 ( .A(n11447), .B(n11539), .Z(n11451) );
  XNOR U5450 ( .A(n12925), .B(n12554), .Z(n12556) );
  XNOR U5451 ( .A(n14029), .B(n13658), .Z(n13660) );
  XNOR U5452 ( .A(n15133), .B(n14762), .Z(n14764) );
  XNOR U5453 ( .A(n16237), .B(n15866), .Z(n15868) );
  XNOR U5454 ( .A(n17341), .B(n16970), .Z(n16972) );
  XNOR U5455 ( .A(n18445), .B(n18074), .Z(n18076) );
  XNOR U5456 ( .A(n19549), .B(n19178), .Z(n19180) );
  XNOR U5457 ( .A(n19917), .B(n19546), .Z(n19548) );
  XNOR U5458 ( .A(n20285), .B(n19914), .Z(n19916) );
  XNOR U5459 ( .A(n20653), .B(n20282), .Z(n20284) );
  XNOR U5460 ( .A(n21021), .B(n20650), .Z(n20652) );
  XNOR U5461 ( .A(n34758), .B(n34842), .Z(n34762) );
  XNOR U5462 ( .A(n34555), .B(n34639), .Z(n34559) );
  XNOR U5463 ( .A(n34328), .B(n34415), .Z(n34332) );
  XNOR U5464 ( .A(n34080), .B(n34164), .Z(n34084) );
  XNOR U5465 ( .A(n33805), .B(n33889), .Z(n33809) );
  XNOR U5466 ( .A(n33506), .B(n33593), .Z(n33510) );
  XNOR U5467 ( .A(n33186), .B(n33270), .Z(n33190) );
  XNOR U5468 ( .A(n32839), .B(n32923), .Z(n32843) );
  XNOR U5469 ( .A(n32468), .B(n32555), .Z(n32472) );
  XNOR U5470 ( .A(n32076), .B(n32160), .Z(n32080) );
  XNOR U5471 ( .A(n31473), .B(n31565), .Z(n31477) );
  XNOR U5472 ( .A(n31017), .B(n31109), .Z(n31021) );
  XNOR U5473 ( .A(n30537), .B(n30629), .Z(n30541) );
  XNOR U5474 ( .A(n30033), .B(n30125), .Z(n30037) );
  XNOR U5475 ( .A(n29505), .B(n29597), .Z(n29509) );
  XNOR U5476 ( .A(n28953), .B(n29045), .Z(n28957) );
  XNOR U5477 ( .A(n28377), .B(n28469), .Z(n28381) );
  XNOR U5478 ( .A(n27777), .B(n27869), .Z(n27781) );
  XNOR U5479 ( .A(n27153), .B(n27245), .Z(n27157) );
  XNOR U5480 ( .A(n26505), .B(n26597), .Z(n26509) );
  XNOR U5481 ( .A(n25833), .B(n25925), .Z(n25837) );
  XNOR U5482 ( .A(n25137), .B(n25229), .Z(n25141) );
  XNOR U5483 ( .A(n24417), .B(n24509), .Z(n24421) );
  XNOR U5484 ( .A(n23596), .B(n23763), .Z(n23600) );
  XNOR U5485 ( .A(n3088), .B(n3208), .Z(n3096) );
  XNOR U5486 ( .A(n2322), .B(n2467), .Z(n2326) );
  XNOR U5487 ( .A(n2283), .B(n2478), .Z(n2278) );
  XNOR U5488 ( .A(n3112), .B(n3202), .Z(n3116) );
  XNOR U5489 ( .A(n3856), .B(n3946), .Z(n3860) );
  XNOR U5490 ( .A(n4605), .B(n4691), .Z(n4600) );
  XNOR U5491 ( .A(n5346), .B(n5436), .Z(n5350) );
  XNOR U5492 ( .A(n6839), .B(n6921), .Z(n6834) );
  XNOR U5493 ( .A(n11083), .B(n11169), .Z(n11087) );
  XNOR U5494 ( .A(n12562), .B(n12191), .Z(n12193) );
  XNOR U5495 ( .A(n13666), .B(n13295), .Z(n13297) );
  XNOR U5496 ( .A(n14770), .B(n14399), .Z(n14401) );
  XNOR U5497 ( .A(n15874), .B(n15503), .Z(n15505) );
  XNOR U5498 ( .A(n16978), .B(n16607), .Z(n16609) );
  XNOR U5499 ( .A(n18082), .B(n17711), .Z(n17713) );
  XNOR U5500 ( .A(n19186), .B(n18815), .Z(n18817) );
  XNOR U5501 ( .A(n19554), .B(n19183), .Z(n19185) );
  XNOR U5502 ( .A(n21388), .B(n21474), .Z(n21392) );
  XNOR U5503 ( .A(n21756), .B(n21842), .Z(n21760) );
  XNOR U5504 ( .A(n22124), .B(n22210), .Z(n22128) );
  XNOR U5505 ( .A(n22492), .B(n22578), .Z(n22496) );
  XNOR U5506 ( .A(n22860), .B(n22946), .Z(n22864) );
  XNOR U5507 ( .A(n1563), .B(n1725), .Z(n1567) );
  XNOR U5508 ( .A(n1520), .B(n1736), .Z(n1528) );
  XNOR U5509 ( .A(n756), .B(n996), .Z(n760) );
  XNOR U5510 ( .A(n717), .B(n1007), .Z(n712) );
  XNOR U5511 ( .A(n2312), .B(n2471), .Z(n2307) );
  XNOR U5512 ( .A(n2351), .B(n2460), .Z(n2355) );
  XNOR U5513 ( .A(n6467), .B(n6551), .Z(n6471) );
  XNOR U5514 ( .A(n11094), .B(n10723), .Z(n10725) );
  XNOR U5515 ( .A(n11825), .B(n11905), .Z(n11829) );
  XNOR U5516 ( .A(n12929), .B(n13009), .Z(n12933) );
  XNOR U5517 ( .A(n14033), .B(n14113), .Z(n14037) );
  XNOR U5518 ( .A(n15137), .B(n15217), .Z(n15141) );
  XNOR U5519 ( .A(n16241), .B(n16321), .Z(n16245) );
  XNOR U5520 ( .A(n17345), .B(n17425), .Z(n17349) );
  XNOR U5521 ( .A(n18449), .B(n18529), .Z(n18453) );
  XNOR U5522 ( .A(n746), .B(n1000), .Z(n741) );
  XNOR U5523 ( .A(n1549), .B(n1729), .Z(n1557) );
  XNOR U5524 ( .A(n785), .B(n989), .Z(n789) );
  XNOR U5525 ( .A(n1592), .B(n1718), .Z(n1596) );
  XNOR U5526 ( .A(n7960), .B(n8038), .Z(n7968) );
  XNOR U5527 ( .A(n8704), .B(n8782), .Z(n8708) );
  XNOR U5528 ( .A(n9447), .B(n9525), .Z(n9448) );
  XNOR U5529 ( .A(n10197), .B(n10385), .Z(n10205) );
  XNOR U5530 ( .A(n11462), .B(n11536), .Z(n11466) );
  XNOR U5531 ( .A(n12940), .B(n12569), .Z(n12571) );
  XNOR U5532 ( .A(n14044), .B(n13673), .Z(n13675) );
  XNOR U5533 ( .A(n15148), .B(n14777), .Z(n14779) );
  XNOR U5534 ( .A(n16252), .B(n15881), .Z(n15883) );
  XNOR U5535 ( .A(n17356), .B(n16985), .Z(n16987) );
  XNOR U5536 ( .A(n18460), .B(n18089), .Z(n18091) );
  XNOR U5537 ( .A(n19564), .B(n19193), .Z(n19195) );
  XNOR U5538 ( .A(n20668), .B(n20297), .Z(n20299) );
  XNOR U5539 ( .A(n21036), .B(n20665), .Z(n20667) );
  XNOR U5540 ( .A(n21404), .B(n21033), .Z(n21035) );
  XNOR U5541 ( .A(n21772), .B(n21401), .Z(n21403) );
  XNOR U5542 ( .A(n22140), .B(n21769), .Z(n21771) );
  XNOR U5543 ( .A(n35104), .B(n35170), .Z(n35108) );
  XNOR U5544 ( .A(n34949), .B(n35018), .Z(n34953) );
  XNOR U5545 ( .A(n34773), .B(n34839), .Z(n34777) );
  XNOR U5546 ( .A(n34570), .B(n34636), .Z(n34574) );
  XNOR U5547 ( .A(n34343), .B(n34412), .Z(n34347) );
  XNOR U5548 ( .A(n34095), .B(n34161), .Z(n34099) );
  XNOR U5549 ( .A(n33820), .B(n33886), .Z(n33824) );
  XNOR U5550 ( .A(n33521), .B(n33590), .Z(n33525) );
  XNOR U5551 ( .A(n33201), .B(n33267), .Z(n33205) );
  XNOR U5552 ( .A(n32854), .B(n32920), .Z(n32858) );
  XNOR U5553 ( .A(n32483), .B(n32552), .Z(n32487) );
  XNOR U5554 ( .A(n32091), .B(n32157), .Z(n32095) );
  XNOR U5555 ( .A(n31488), .B(n31562), .Z(n31492) );
  XNOR U5556 ( .A(n31032), .B(n31106), .Z(n31036) );
  XNOR U5557 ( .A(n30552), .B(n30626), .Z(n30556) );
  XNOR U5558 ( .A(n30048), .B(n30122), .Z(n30052) );
  XNOR U5559 ( .A(n29520), .B(n29594), .Z(n29524) );
  XNOR U5560 ( .A(n28968), .B(n29042), .Z(n28972) );
  XNOR U5561 ( .A(n28392), .B(n28466), .Z(n28396) );
  XNOR U5562 ( .A(n27792), .B(n27866), .Z(n27796) );
  XNOR U5563 ( .A(n27168), .B(n27242), .Z(n27172) );
  XNOR U5564 ( .A(n26520), .B(n26594), .Z(n26524) );
  XNOR U5565 ( .A(n25848), .B(n25922), .Z(n25852) );
  XNOR U5566 ( .A(n25152), .B(n25226), .Z(n25156) );
  XNOR U5567 ( .A(n24432), .B(n24506), .Z(n24436) );
  XNOR U5568 ( .A(n23611), .B(n23760), .Z(n23615) );
  XNOR U5569 ( .A(n2341), .B(n2464), .Z(n2336) );
  XNOR U5570 ( .A(n3871), .B(n3943), .Z(n3879) );
  XNOR U5571 ( .A(n4615), .B(n4687), .Z(n4619) );
  XNOR U5572 ( .A(n5363), .B(n5432), .Z(n5364) );
  XNOR U5573 ( .A(n6105), .B(n6177), .Z(n6113) );
  XNOR U5574 ( .A(n7595), .B(n7664), .Z(n7596) );
  XNOR U5575 ( .A(n11098), .B(n11166), .Z(n11102) );
  XNOR U5576 ( .A(n12577), .B(n12206), .Z(n12208) );
  XNOR U5577 ( .A(n13681), .B(n13310), .Z(n13312) );
  XNOR U5578 ( .A(n14785), .B(n14414), .Z(n14416) );
  XNOR U5579 ( .A(n15889), .B(n15518), .Z(n15520) );
  XNOR U5580 ( .A(n16993), .B(n16622), .Z(n16624) );
  XNOR U5581 ( .A(n18097), .B(n17726), .Z(n17728) );
  XNOR U5582 ( .A(n19201), .B(n18830), .Z(n18832) );
  XNOR U5583 ( .A(n20305), .B(n19934), .Z(n19936) );
  XNOR U5584 ( .A(n20673), .B(n20302), .Z(n20304) );
  XNOR U5585 ( .A(n22507), .B(n22575), .Z(n22511) );
  XNOR U5586 ( .A(n22875), .B(n22943), .Z(n22879) );
  XNOR U5587 ( .A(n2003), .B(n2081), .Z(n2007) );
  XNOR U5588 ( .A(n1578), .B(n1722), .Z(n1586) );
  XNOR U5589 ( .A(n814), .B(n982), .Z(n818) );
  XNOR U5590 ( .A(n775), .B(n993), .Z(n770) );
  XNOR U5591 ( .A(n2370), .B(n2457), .Z(n2365) );
  XNOR U5592 ( .A(n3506), .B(n3569), .Z(n3507) );
  XNOR U5593 ( .A(n7222), .B(n7291), .Z(n7226) );
  XNOR U5594 ( .A(n11109), .B(n10738), .Z(n10740) );
  XNOR U5595 ( .A(n11840), .B(n11902), .Z(n11844) );
  XNOR U5596 ( .A(n12944), .B(n13006), .Z(n12948) );
  XNOR U5597 ( .A(n14048), .B(n14110), .Z(n14052) );
  XNOR U5598 ( .A(n15152), .B(n15214), .Z(n15156) );
  XNOR U5599 ( .A(n16256), .B(n16318), .Z(n16260) );
  XNOR U5600 ( .A(n17360), .B(n17422), .Z(n17364) );
  XNOR U5601 ( .A(n18464), .B(n18526), .Z(n18468) );
  XNOR U5602 ( .A(n19568), .B(n19630), .Z(n19572) );
  XNOR U5603 ( .A(n1244), .B(n1340), .Z(n1248) );
  XNOR U5604 ( .A(n804), .B(n986), .Z(n799) );
  XNOR U5605 ( .A(n1607), .B(n1715), .Z(n1615) );
  XNOR U5606 ( .A(n843), .B(n975), .Z(n847) );
  XNOR U5607 ( .A(n8723), .B(n8779), .Z(n8718) );
  XNOR U5608 ( .A(n9459), .B(n9522), .Z(n9463) );
  XNOR U5609 ( .A(n10211), .B(n10380), .Z(n10215) );
  XNOR U5610 ( .A(n11477), .B(n11533), .Z(n11481) );
  XNOR U5611 ( .A(n12955), .B(n12584), .Z(n12586) );
  XNOR U5612 ( .A(n14059), .B(n13688), .Z(n13690) );
  XNOR U5613 ( .A(n15163), .B(n14792), .Z(n14794) );
  XNOR U5614 ( .A(n16267), .B(n15896), .Z(n15898) );
  XNOR U5615 ( .A(n17371), .B(n17000), .Z(n17002) );
  XNOR U5616 ( .A(n18475), .B(n18104), .Z(n18106) );
  XNOR U5617 ( .A(n19579), .B(n19208), .Z(n19210) );
  XNOR U5618 ( .A(n20683), .B(n20312), .Z(n20314) );
  XNOR U5619 ( .A(n21787), .B(n21416), .Z(n21418) );
  XNOR U5620 ( .A(n22155), .B(n21784), .Z(n21786) );
  XNOR U5621 ( .A(n22523), .B(n22152), .Z(n22154) );
  XNOR U5622 ( .A(n22891), .B(n22520), .Z(n22522) );
  XNOR U5623 ( .A(n23259), .B(n22888), .Z(n22890) );
  XNOR U5624 ( .A(n35250), .B(n35298), .Z(n35254) );
  XNOR U5625 ( .A(n35119), .B(n35167), .Z(n35123) );
  XNOR U5626 ( .A(n34964), .B(n35015), .Z(n34968) );
  XNOR U5627 ( .A(n34788), .B(n34836), .Z(n34792) );
  XNOR U5628 ( .A(n34585), .B(n34633), .Z(n34589) );
  XNOR U5629 ( .A(n34358), .B(n34409), .Z(n34362) );
  XNOR U5630 ( .A(n34110), .B(n34158), .Z(n34114) );
  XNOR U5631 ( .A(n33835), .B(n33883), .Z(n33839) );
  XNOR U5632 ( .A(n33536), .B(n33587), .Z(n33540) );
  XNOR U5633 ( .A(n33216), .B(n33264), .Z(n33220) );
  XNOR U5634 ( .A(n32869), .B(n32917), .Z(n32873) );
  XNOR U5635 ( .A(n32498), .B(n32549), .Z(n32502) );
  XNOR U5636 ( .A(n32106), .B(n32154), .Z(n32110) );
  XNOR U5637 ( .A(n31503), .B(n31559), .Z(n31507) );
  XNOR U5638 ( .A(n31047), .B(n31103), .Z(n31051) );
  XNOR U5639 ( .A(n30567), .B(n30623), .Z(n30571) );
  XNOR U5640 ( .A(n30063), .B(n30119), .Z(n30067) );
  XNOR U5641 ( .A(n29535), .B(n29591), .Z(n29539) );
  XNOR U5642 ( .A(n28983), .B(n29039), .Z(n28987) );
  XNOR U5643 ( .A(n28407), .B(n28463), .Z(n28411) );
  XNOR U5644 ( .A(n27807), .B(n27863), .Z(n27811) );
  XNOR U5645 ( .A(n27183), .B(n27239), .Z(n27187) );
  XNOR U5646 ( .A(n26535), .B(n26591), .Z(n26539) );
  XNOR U5647 ( .A(n25863), .B(n25919), .Z(n25867) );
  XNOR U5648 ( .A(n25167), .B(n25223), .Z(n25171) );
  XNOR U5649 ( .A(n24447), .B(n24503), .Z(n24451) );
  XNOR U5650 ( .A(n23626), .B(n23757), .Z(n23630) );
  XNOR U5651 ( .A(n892), .B(n964), .Z(n896) );
  XNOR U5652 ( .A(n1651), .B(n1705), .Z(n1655) );
  XNOR U5653 ( .A(n2395), .B(n2449), .Z(n2399) );
  XNOR U5654 ( .A(n3141), .B(n3195), .Z(n3145) );
  XNOR U5655 ( .A(n4634), .B(n4684), .Z(n4629) );
  XNOR U5656 ( .A(n5375), .B(n5429), .Z(n5379) );
  XNOR U5657 ( .A(n6119), .B(n6173), .Z(n6123) );
  XNOR U5658 ( .A(n6868), .B(n6914), .Z(n6863) );
  XNOR U5659 ( .A(n8351), .B(n8405), .Z(n8355) );
  XNOR U5660 ( .A(n11113), .B(n11163), .Z(n11117) );
  XNOR U5661 ( .A(n12592), .B(n12221), .Z(n12223) );
  XNOR U5662 ( .A(n13696), .B(n13325), .Z(n13327) );
  XNOR U5663 ( .A(n14800), .B(n14429), .Z(n14431) );
  XNOR U5664 ( .A(n15904), .B(n15533), .Z(n15535) );
  XNOR U5665 ( .A(n17008), .B(n16637), .Z(n16639) );
  XNOR U5666 ( .A(n18112), .B(n17741), .Z(n17743) );
  XNOR U5667 ( .A(n19216), .B(n18845), .Z(n18847) );
  XNOR U5668 ( .A(n20320), .B(n19949), .Z(n19951) );
  XNOR U5669 ( .A(n21424), .B(n21053), .Z(n21055) );
  XNOR U5670 ( .A(n21792), .B(n21421), .Z(n21423) );
  XNOR U5671 ( .A(n1636), .B(n1708), .Z(n1640) );
  XNOR U5672 ( .A(n833), .B(n979), .Z(n828) );
  XNOR U5673 ( .A(n4262), .B(n4310), .Z(n4266) );
  XNOR U5674 ( .A(n7612), .B(n7660), .Z(n7620) );
  XNOR U5675 ( .A(n10750), .B(n10793), .Z(n10754) );
  XNOR U5676 ( .A(n11855), .B(n11899), .Z(n11859) );
  XNOR U5677 ( .A(n12959), .B(n13003), .Z(n12963) );
  XNOR U5678 ( .A(n14063), .B(n14107), .Z(n14067) );
  XNOR U5679 ( .A(n15167), .B(n15211), .Z(n15171) );
  XNOR U5680 ( .A(n16271), .B(n16315), .Z(n16275) );
  XNOR U5681 ( .A(n17375), .B(n17419), .Z(n17379) );
  XNOR U5682 ( .A(n18479), .B(n18523), .Z(n18483) );
  XNOR U5683 ( .A(n19583), .B(n19627), .Z(n19587) );
  XNOR U5684 ( .A(n20687), .B(n20731), .Z(n20691) );
  XNOR U5685 ( .A(n877), .B(n967), .Z(n881) );
  XNOR U5686 ( .A(n862), .B(n972), .Z(n857) );
  XNOR U5687 ( .A(n9476), .B(n9518), .Z(n9477) );
  XNOR U5688 ( .A(n10226), .B(n10374), .Z(n10234) );
  XNOR U5689 ( .A(n11492), .B(n11530), .Z(n11496) );
  XNOR U5690 ( .A(n12970), .B(n12599), .Z(n12601) );
  XNOR U5691 ( .A(n14074), .B(n13703), .Z(n13705) );
  XNOR U5692 ( .A(n15178), .B(n14807), .Z(n14809) );
  XNOR U5693 ( .A(n16282), .B(n15911), .Z(n15913) );
  XNOR U5694 ( .A(n17386), .B(n17015), .Z(n17017) );
  XNOR U5695 ( .A(n18490), .B(n18119), .Z(n18121) );
  XNOR U5696 ( .A(n19594), .B(n19223), .Z(n19225) );
  XNOR U5697 ( .A(n20698), .B(n20327), .Z(n20329) );
  XNOR U5698 ( .A(n21802), .B(n21431), .Z(n21433) );
  XNOR U5699 ( .A(n22906), .B(n22535), .Z(n22537) );
  XNOR U5700 ( .A(n23274), .B(n22903), .Z(n22905) );
  XNOR U5701 ( .A(n23268), .B(n23306), .Z(n23272) );
  XNOR U5702 ( .A(n35452), .B(n35482), .Z(n35456) );
  XNOR U5703 ( .A(n35369), .B(n35402), .Z(n35373) );
  XNOR U5704 ( .A(n35265), .B(n35295), .Z(n35269) );
  XNOR U5705 ( .A(n35134), .B(n35164), .Z(n35138) );
  XNOR U5706 ( .A(n34979), .B(n35012), .Z(n34983) );
  XNOR U5707 ( .A(n34803), .B(n34833), .Z(n34807) );
  XNOR U5708 ( .A(n34600), .B(n34630), .Z(n34604) );
  XNOR U5709 ( .A(n34373), .B(n34406), .Z(n34377) );
  XNOR U5710 ( .A(n34125), .B(n34155), .Z(n34129) );
  XNOR U5711 ( .A(n33850), .B(n33880), .Z(n33854) );
  XNOR U5712 ( .A(n33551), .B(n33584), .Z(n33555) );
  XNOR U5713 ( .A(n33231), .B(n33261), .Z(n33235) );
  XNOR U5714 ( .A(n32884), .B(n32914), .Z(n32888) );
  XNOR U5715 ( .A(n32513), .B(n32546), .Z(n32517) );
  XNOR U5716 ( .A(n32121), .B(n32151), .Z(n32125) );
  XNOR U5717 ( .A(n31518), .B(n31556), .Z(n31522) );
  XNOR U5718 ( .A(n31062), .B(n31100), .Z(n31066) );
  XNOR U5719 ( .A(n30582), .B(n30620), .Z(n30586) );
  XNOR U5720 ( .A(n30078), .B(n30116), .Z(n30082) );
  XNOR U5721 ( .A(n29550), .B(n29588), .Z(n29554) );
  XNOR U5722 ( .A(n28998), .B(n29036), .Z(n29002) );
  XNOR U5723 ( .A(n28422), .B(n28460), .Z(n28426) );
  XNOR U5724 ( .A(n27822), .B(n27860), .Z(n27826) );
  XNOR U5725 ( .A(n27198), .B(n27236), .Z(n27202) );
  XNOR U5726 ( .A(n26550), .B(n26588), .Z(n26554) );
  XNOR U5727 ( .A(n25878), .B(n25916), .Z(n25882) );
  XNOR U5728 ( .A(n25182), .B(n25220), .Z(n25186) );
  XNOR U5729 ( .A(n24462), .B(n24500), .Z(n24466) );
  XNOR U5730 ( .A(n907), .B(n961), .Z(n911) );
  XNOR U5731 ( .A(n922), .B(n958), .Z(n926) );
  XNOR U5732 ( .A(n2410), .B(n2446), .Z(n2414) );
  XNOR U5733 ( .A(n3156), .B(n3192), .Z(n3160) );
  XNOR U5734 ( .A(n3900), .B(n3936), .Z(n3904) );
  XNOR U5735 ( .A(n5392), .B(n5425), .Z(n5393) );
  XNOR U5736 ( .A(n6506), .B(n6542), .Z(n6510) );
  XNOR U5737 ( .A(n7246), .B(n7285), .Z(n7250) );
  XNOR U5738 ( .A(n8738), .B(n8774), .Z(n8742) );
  XNOR U5739 ( .A(n11128), .B(n11160), .Z(n11132) );
  XNOR U5740 ( .A(n12607), .B(n12236), .Z(n12238) );
  XNOR U5741 ( .A(n13711), .B(n13340), .Z(n13342) );
  XNOR U5742 ( .A(n14815), .B(n14444), .Z(n14446) );
  XNOR U5743 ( .A(n15919), .B(n15548), .Z(n15550) );
  XNOR U5744 ( .A(n17023), .B(n16652), .Z(n16654) );
  XNOR U5745 ( .A(n18127), .B(n17756), .Z(n17758) );
  XNOR U5746 ( .A(n19231), .B(n18860), .Z(n18862) );
  XNOR U5747 ( .A(n20335), .B(n19964), .Z(n19966) );
  XNOR U5748 ( .A(n21439), .B(n21068), .Z(n21070) );
  XNOR U5749 ( .A(n22543), .B(n22172), .Z(n22174) );
  XNOR U5750 ( .A(n22911), .B(n22540), .Z(n22542) );
  XNOR U5751 ( .A(n4649), .B(n4679), .Z(n4653) );
  XNOR U5752 ( .A(n6143), .B(n6169), .Z(n6138) );
  XNOR U5753 ( .A(n8375), .B(n8401), .Z(n8370) );
  XNOR U5754 ( .A(n10765), .B(n10790), .Z(n10769) );
  XNOR U5755 ( .A(n11870), .B(n11896), .Z(n11874) );
  XNOR U5756 ( .A(n12974), .B(n13000), .Z(n12978) );
  XNOR U5757 ( .A(n14078), .B(n14104), .Z(n14082) );
  XNOR U5758 ( .A(n15182), .B(n15208), .Z(n15186) );
  XNOR U5759 ( .A(n16286), .B(n16312), .Z(n16290) );
  XNOR U5760 ( .A(n17390), .B(n17416), .Z(n17394) );
  XNOR U5761 ( .A(n18494), .B(n18520), .Z(n18498) );
  XNOR U5762 ( .A(n19598), .B(n19624), .Z(n19602) );
  XNOR U5763 ( .A(n20702), .B(n20728), .Z(n20706) );
  XNOR U5764 ( .A(n21806), .B(n21832), .Z(n21810) );
  XNOR U5765 ( .A(n23651), .B(n23752), .Z(n23655) );
  XNOR U5766 ( .A(n2048), .B(n2072), .Z(n2052) );
  XNOR U5767 ( .A(n9863), .B(n9887), .Z(n9867) );
  XNOR U5768 ( .A(n11507), .B(n11527), .Z(n11511) );
  XNOR U5769 ( .A(n12985), .B(n12614), .Z(n12616) );
  XNOR U5770 ( .A(n14089), .B(n13718), .Z(n13720) );
  XNOR U5771 ( .A(n15193), .B(n14822), .Z(n14824) );
  XNOR U5772 ( .A(n16297), .B(n15926), .Z(n15928) );
  XNOR U5773 ( .A(n17401), .B(n17030), .Z(n17032) );
  XNOR U5774 ( .A(n18505), .B(n18134), .Z(n18136) );
  XNOR U5775 ( .A(n19609), .B(n19238), .Z(n19240) );
  XNOR U5776 ( .A(n20713), .B(n20342), .Z(n20344) );
  XNOR U5777 ( .A(n21817), .B(n21446), .Z(n21448) );
  XNOR U5778 ( .A(n22921), .B(n22550), .Z(n22552) );
  XNOR U5779 ( .A(n35526), .B(n35538), .Z(n35530) );
  XNOR U5780 ( .A(n35467), .B(n35479), .Z(n35472) );
  XNOR U5781 ( .A(n35384), .B(n35399), .Z(n35393) );
  XNOR U5782 ( .A(n35280), .B(n35292), .Z(n35284) );
  XNOR U5783 ( .A(n35149), .B(n35161), .Z(n35154) );
  XNOR U5784 ( .A(n34994), .B(n35009), .Z(n35003) );
  XNOR U5785 ( .A(n34818), .B(n34830), .Z(n34822) );
  XNOR U5786 ( .A(n34615), .B(n34627), .Z(n34620) );
  XNOR U5787 ( .A(n34388), .B(n34403), .Z(n34397) );
  XNOR U5788 ( .A(n34140), .B(n34152), .Z(n34144) );
  XNOR U5789 ( .A(n33865), .B(n33877), .Z(n33870) );
  XNOR U5790 ( .A(n33566), .B(n33581), .Z(n33575) );
  XNOR U5791 ( .A(n33246), .B(n33258), .Z(n33250) );
  XNOR U5792 ( .A(n32899), .B(n32911), .Z(n32904) );
  XNOR U5793 ( .A(n32528), .B(n32543), .Z(n32537) );
  XNOR U5794 ( .A(n32136), .B(n32148), .Z(n32140) );
  XNOR U5795 ( .A(n31533), .B(n31553), .Z(n31542) );
  XNOR U5796 ( .A(n31077), .B(n31097), .Z(n31086) );
  XNOR U5797 ( .A(n30597), .B(n30617), .Z(n30606) );
  XNOR U5798 ( .A(n30093), .B(n30113), .Z(n30102) );
  XNOR U5799 ( .A(n29565), .B(n29585), .Z(n29574) );
  XNOR U5800 ( .A(n29013), .B(n29033), .Z(n29022) );
  XNOR U5801 ( .A(n28437), .B(n28457), .Z(n28446) );
  XNOR U5802 ( .A(n27837), .B(n27857), .Z(n27846) );
  XNOR U5803 ( .A(n27213), .B(n27233), .Z(n27222) );
  XNOR U5804 ( .A(n26565), .B(n26585), .Z(n26574) );
  XNOR U5805 ( .A(n25893), .B(n25913), .Z(n25902) );
  XNOR U5806 ( .A(n25197), .B(n25217), .Z(n25206) );
  XNOR U5807 ( .A(n24477), .B(n24497), .Z(n24486) );
  XNOR U5808 ( .A(n937), .B(n955), .Z(n946) );
  XNOR U5809 ( .A(n1681), .B(n1699), .Z(n1690) );
  XNOR U5810 ( .A(n2798), .B(n2817), .Z(n2806) );
  XNOR U5811 ( .A(n3543), .B(n3561), .Z(n3552) );
  XNOR U5812 ( .A(n4287), .B(n4305), .Z(n4296) );
  XNOR U5813 ( .A(n5776), .B(n5794), .Z(n5785) );
  XNOR U5814 ( .A(n7261), .B(n7282), .Z(n7265) );
  XNOR U5815 ( .A(n8008), .B(n8026), .Z(n8017) );
  XNOR U5816 ( .A(n9493), .B(n9514), .Z(n9497) );
  XNOR U5817 ( .A(n11143), .B(n11157), .Z(n11147) );
  XNOR U5818 ( .A(n12248), .B(n12262), .Z(n12252) );
  XNOR U5819 ( .A(n13352), .B(n13366), .Z(n13356) );
  XNOR U5820 ( .A(n14456), .B(n14470), .Z(n14460) );
  XNOR U5821 ( .A(n15560), .B(n15574), .Z(n15564) );
  XNOR U5822 ( .A(n16664), .B(n16678), .Z(n16668) );
  XNOR U5823 ( .A(n17768), .B(n17782), .Z(n17772) );
  XNOR U5824 ( .A(n18872), .B(n18886), .Z(n18876) );
  XNOR U5825 ( .A(n19976), .B(n19990), .Z(n19980) );
  XNOR U5826 ( .A(n21080), .B(n21094), .Z(n21084) );
  XNOR U5827 ( .A(n22184), .B(n22198), .Z(n22188) );
  XNOR U5828 ( .A(n23288), .B(n23302), .Z(n23292) );
  XNOR U5829 ( .A(n5039), .B(n5046), .Z(n5035) );
  XNOR U5830 ( .A(n6892), .B(n6906), .Z(n6900) );
  XNOR U5831 ( .A(n9124), .B(n9138), .Z(n9132) );
  XOR U5832 ( .A(n10780), .B(n10787), .Z(n10784) );
  XOR U5833 ( .A(n11885), .B(n11892), .Z(n11890) );
  XOR U5834 ( .A(n12989), .B(n12996), .Z(n12994) );
  XOR U5835 ( .A(n14093), .B(n14100), .Z(n14098) );
  XOR U5836 ( .A(n15197), .B(n15204), .Z(n15202) );
  XOR U5837 ( .A(n16301), .B(n16308), .Z(n16306) );
  XOR U5838 ( .A(n17405), .B(n17412), .Z(n17410) );
  XOR U5839 ( .A(n18509), .B(n18516), .Z(n18514) );
  XOR U5840 ( .A(n19613), .B(n19620), .Z(n19618) );
  XOR U5841 ( .A(n20717), .B(n20724), .Z(n20722) );
  XOR U5842 ( .A(n21821), .B(n21828), .Z(n21826) );
  XOR U5843 ( .A(n22925), .B(n22932), .Z(n22930) );
  ANDN U5844 ( .B(n1320), .A(n1319), .Z(n947) );
  NANDN U5845 ( .A(n2808), .B(n2809), .Z(n2435) );
  NANDN U5846 ( .A(n4297), .B(n4298), .Z(n3925) );
  XOR U5847 ( .A(n5049), .B(n5414), .Z(n5416) );
  XOR U5848 ( .A(n6164), .B(n6530), .Z(n6532) );
  XNOR U5849 ( .A(n7646), .B(n7648), .Z(n7647) );
  XNOR U5850 ( .A(n8762), .B(n8764), .Z(n8763) );
  XNOR U5851 ( .A(n9878), .B(n9880), .Z(n9879) );
  XOR U5852 ( .A(n10265), .B(n7), .Z(n10264) );
  XOR U5853 ( .A(n10274), .B(n13), .Z(n10273) );
  XOR U5854 ( .A(n10283), .B(n19), .Z(n10282) );
  XOR U5855 ( .A(n10292), .B(n25), .Z(n10291) );
  XOR U5856 ( .A(n10301), .B(n31), .Z(n10300) );
  XOR U5857 ( .A(n10310), .B(n37), .Z(n10309) );
  XOR U5858 ( .A(n10319), .B(n43), .Z(n10318) );
  XOR U5859 ( .A(n10328), .B(n49), .Z(n10327) );
  XOR U5860 ( .A(n10337), .B(n55), .Z(n10336) );
  XOR U5861 ( .A(n10346), .B(n61), .Z(n10345) );
  AND U5862 ( .A(n71), .B(n72), .Z(n69) );
  XNOR U5863 ( .A(n23819), .B(n24182), .Z(n23824) );
  XNOR U5864 ( .A(n8472), .B(n8833), .Z(n8477) );
  XNOR U5865 ( .A(n9212), .B(n9576), .Z(n9217) );
  XNOR U5866 ( .A(n9964), .B(n10476), .Z(n9969) );
  XNOR U5867 ( .A(n10489), .B(n10845), .Z(n10494) );
  XNOR U5868 ( .A(n10857), .B(n11214), .Z(n10862) );
  XNOR U5869 ( .A(n11601), .B(n11230), .Z(n11231) );
  XNOR U5870 ( .A(n14171), .B(n14528), .Z(n14176) );
  XNOR U5871 ( .A(n14907), .B(n15264), .Z(n14912) );
  XNOR U5872 ( .A(n18587), .B(n18944), .Z(n18592) );
  XNOR U5873 ( .A(n19323), .B(n19680), .Z(n19328) );
  XNOR U5874 ( .A(n23003), .B(n23360), .Z(n23008) );
  XNOR U5875 ( .A(n7728), .B(n8089), .Z(n7733) );
  XNOR U5876 ( .A(n11973), .B(n12319), .Z(n11968) );
  XNOR U5877 ( .A(n15649), .B(n15999), .Z(n15653) );
  XNOR U5878 ( .A(n16385), .B(n16735), .Z(n16389) );
  XNOR U5879 ( .A(n20065), .B(n20415), .Z(n20069) );
  XNOR U5880 ( .A(n20801), .B(n21151), .Z(n20805) );
  XNOR U5881 ( .A(n12710), .B(n13054), .Z(n12718) );
  XNOR U5882 ( .A(n13446), .B(n13790), .Z(n13450) );
  XNOR U5883 ( .A(n17126), .B(n17470), .Z(n17130) );
  XNOR U5884 ( .A(n17862), .B(n18206), .Z(n17866) );
  XNOR U5885 ( .A(n21542), .B(n21886), .Z(n21546) );
  XNOR U5886 ( .A(n22278), .B(n22622), .Z(n22282) );
  XNOR U5887 ( .A(n25278), .B(n25622), .Z(n25282) );
  XNOR U5888 ( .A(n24570), .B(n24914), .Z(n24574) );
  XNOR U5889 ( .A(n23835), .B(n24179), .Z(n23839) );
  XNOR U5890 ( .A(n8488), .B(n8830), .Z(n8492) );
  XNOR U5891 ( .A(n9228), .B(n9573), .Z(n9232) );
  XNOR U5892 ( .A(n9980), .B(n10470), .Z(n9984) );
  XNOR U5893 ( .A(n10505), .B(n10842), .Z(n10509) );
  XNOR U5894 ( .A(n10873), .B(n11211), .Z(n10877) );
  XNOR U5895 ( .A(n11242), .B(n11580), .Z(n11246) );
  XNOR U5896 ( .A(n11984), .B(n11613), .Z(n11615) );
  XNOR U5897 ( .A(n12352), .B(n11981), .Z(n11983) );
  XNOR U5898 ( .A(n12720), .B(n12349), .Z(n12351) );
  XNOR U5899 ( .A(n14187), .B(n14525), .Z(n14191) );
  XNOR U5900 ( .A(n14923), .B(n15261), .Z(n14927) );
  XNOR U5901 ( .A(n18603), .B(n18941), .Z(n18607) );
  XNOR U5902 ( .A(n19339), .B(n19677), .Z(n19343) );
  XNOR U5903 ( .A(n23019), .B(n23357), .Z(n23023) );
  XNOR U5904 ( .A(n7362), .B(n7716), .Z(n7366) );
  XNOR U5905 ( .A(n15664), .B(n15996), .Z(n15668) );
  XNOR U5906 ( .A(n16400), .B(n16732), .Z(n16404) );
  XNOR U5907 ( .A(n20080), .B(n20412), .Z(n20084) );
  XNOR U5908 ( .A(n20816), .B(n21148), .Z(n20820) );
  XNOR U5909 ( .A(n13465), .B(n13787), .Z(n13460) );
  XNOR U5910 ( .A(n17141), .B(n17467), .Z(n17145) );
  XNOR U5911 ( .A(n17877), .B(n18203), .Z(n17881) );
  XNOR U5912 ( .A(n21557), .B(n21883), .Z(n21561) );
  XNOR U5913 ( .A(n22293), .B(n22619), .Z(n22297) );
  XNOR U5914 ( .A(n25977), .B(n26303), .Z(n25981) );
  XNOR U5915 ( .A(n25293), .B(n25619), .Z(n25297) );
  XNOR U5916 ( .A(n24585), .B(n24911), .Z(n24589) );
  XNOR U5917 ( .A(n23850), .B(n24176), .Z(n23854) );
  XNOR U5918 ( .A(n8503), .B(n8827), .Z(n8507) );
  XNOR U5919 ( .A(n9243), .B(n9570), .Z(n9247) );
  XNOR U5920 ( .A(n9995), .B(n10464), .Z(n9999) );
  XNOR U5921 ( .A(n10520), .B(n10839), .Z(n10524) );
  XNOR U5922 ( .A(n10888), .B(n11208), .Z(n10892) );
  XNOR U5923 ( .A(n11257), .B(n11577), .Z(n11261) );
  XNOR U5924 ( .A(n11999), .B(n11628), .Z(n11630) );
  XNOR U5925 ( .A(n12367), .B(n11996), .Z(n11998) );
  XNOR U5926 ( .A(n12735), .B(n12364), .Z(n12366) );
  XNOR U5927 ( .A(n13103), .B(n12732), .Z(n12734) );
  XNOR U5928 ( .A(n13471), .B(n13100), .Z(n13102) );
  XNOR U5929 ( .A(n13839), .B(n13468), .Z(n13470) );
  XNOR U5930 ( .A(n14202), .B(n14522), .Z(n14210) );
  XNOR U5931 ( .A(n14938), .B(n15258), .Z(n14942) );
  XNOR U5932 ( .A(n18618), .B(n18938), .Z(n18622) );
  XNOR U5933 ( .A(n19354), .B(n19674), .Z(n19358) );
  XNOR U5934 ( .A(n23034), .B(n23354), .Z(n23038) );
  XNOR U5935 ( .A(n7377), .B(n7713), .Z(n7381) );
  XNOR U5936 ( .A(n6613), .B(n6970), .Z(n6618) );
  XNOR U5937 ( .A(n15679), .B(n15993), .Z(n15683) );
  XNOR U5938 ( .A(n16415), .B(n16729), .Z(n16419) );
  XNOR U5939 ( .A(n20095), .B(n20409), .Z(n20099) );
  XNOR U5940 ( .A(n20831), .B(n21145), .Z(n20835) );
  XNOR U5941 ( .A(n17156), .B(n17464), .Z(n17160) );
  XNOR U5942 ( .A(n17892), .B(n18200), .Z(n17896) );
  XNOR U5943 ( .A(n21572), .B(n21880), .Z(n21576) );
  XNOR U5944 ( .A(n22308), .B(n22616), .Z(n22312) );
  XNOR U5945 ( .A(n27288), .B(n27596), .Z(n27292) );
  XNOR U5946 ( .A(n26652), .B(n26960), .Z(n26656) );
  XNOR U5947 ( .A(n25992), .B(n26300), .Z(n25996) );
  XNOR U5948 ( .A(n25308), .B(n25616), .Z(n25312) );
  XNOR U5949 ( .A(n24600), .B(n24908), .Z(n24604) );
  XNOR U5950 ( .A(n23865), .B(n24173), .Z(n23869) );
  XNOR U5951 ( .A(n8518), .B(n8824), .Z(n8522) );
  XNOR U5952 ( .A(n9258), .B(n9567), .Z(n9262) );
  XNOR U5953 ( .A(n10010), .B(n10458), .Z(n10014) );
  XNOR U5954 ( .A(n10535), .B(n10836), .Z(n10539) );
  XNOR U5955 ( .A(n10903), .B(n11205), .Z(n10907) );
  XNOR U5956 ( .A(n11272), .B(n11574), .Z(n11276) );
  XNOR U5957 ( .A(n12014), .B(n11643), .Z(n11645) );
  XNOR U5958 ( .A(n12382), .B(n12011), .Z(n12013) );
  XNOR U5959 ( .A(n12750), .B(n12379), .Z(n12381) );
  XNOR U5960 ( .A(n13118), .B(n12747), .Z(n12749) );
  XNOR U5961 ( .A(n13486), .B(n13115), .Z(n13117) );
  XNOR U5962 ( .A(n13854), .B(n13483), .Z(n13485) );
  XNOR U5963 ( .A(n14222), .B(n13851), .Z(n13853) );
  XNOR U5964 ( .A(n14590), .B(n14219), .Z(n14221) );
  XNOR U5965 ( .A(n14958), .B(n14587), .Z(n14589) );
  XNOR U5966 ( .A(n14957), .B(n15255), .Z(n14952) );
  XNOR U5967 ( .A(n18633), .B(n18935), .Z(n18637) );
  XNOR U5968 ( .A(n19369), .B(n19671), .Z(n19373) );
  XNOR U5969 ( .A(n23049), .B(n23351), .Z(n23053) );
  XNOR U5970 ( .A(n7774), .B(n8080), .Z(n7778) );
  XNOR U5971 ( .A(n7007), .B(n7340), .Z(n7011) );
  XNOR U5972 ( .A(n6247), .B(n6601), .Z(n6251) );
  XNOR U5973 ( .A(n15694), .B(n15990), .Z(n15702) );
  XNOR U5974 ( .A(n16430), .B(n16726), .Z(n16434) );
  XNOR U5975 ( .A(n20110), .B(n20406), .Z(n20114) );
  XNOR U5976 ( .A(n20846), .B(n21142), .Z(n20850) );
  XNOR U5977 ( .A(n17171), .B(n17461), .Z(n17175) );
  XNOR U5978 ( .A(n17907), .B(n18197), .Z(n17911) );
  XNOR U5979 ( .A(n21587), .B(n21877), .Z(n21591) );
  XNOR U5980 ( .A(n22323), .B(n22613), .Z(n22327) );
  XNOR U5981 ( .A(n27915), .B(n28205), .Z(n27919) );
  XNOR U5982 ( .A(n27303), .B(n27593), .Z(n27307) );
  XNOR U5983 ( .A(n26667), .B(n26957), .Z(n26671) );
  XNOR U5984 ( .A(n26007), .B(n26297), .Z(n26011) );
  XNOR U5985 ( .A(n25323), .B(n25613), .Z(n25327) );
  XNOR U5986 ( .A(n24615), .B(n24905), .Z(n24619) );
  XNOR U5987 ( .A(n23880), .B(n24170), .Z(n23884) );
  XNOR U5988 ( .A(n8533), .B(n8821), .Z(n8537) );
  XNOR U5989 ( .A(n9273), .B(n9564), .Z(n9277) );
  XNOR U5990 ( .A(n10025), .B(n10452), .Z(n10029) );
  XNOR U5991 ( .A(n10550), .B(n10833), .Z(n10554) );
  XNOR U5992 ( .A(n10918), .B(n11202), .Z(n10922) );
  XNOR U5993 ( .A(n11287), .B(n11571), .Z(n11291) );
  XNOR U5994 ( .A(n12029), .B(n11658), .Z(n11660) );
  XNOR U5995 ( .A(n12397), .B(n12026), .Z(n12028) );
  XNOR U5996 ( .A(n12765), .B(n12394), .Z(n12396) );
  XNOR U5997 ( .A(n13133), .B(n12762), .Z(n12764) );
  XNOR U5998 ( .A(n13501), .B(n13130), .Z(n13132) );
  XNOR U5999 ( .A(n13869), .B(n13498), .Z(n13500) );
  XNOR U6000 ( .A(n14237), .B(n13866), .Z(n13868) );
  XNOR U6001 ( .A(n14605), .B(n14234), .Z(n14236) );
  XNOR U6002 ( .A(n14973), .B(n14602), .Z(n14604) );
  XNOR U6003 ( .A(n15341), .B(n14970), .Z(n14972) );
  XNOR U6004 ( .A(n15709), .B(n15338), .Z(n15340) );
  XNOR U6005 ( .A(n16077), .B(n15706), .Z(n15708) );
  XNOR U6006 ( .A(n18648), .B(n18932), .Z(n18652) );
  XNOR U6007 ( .A(n19384), .B(n19668), .Z(n19388) );
  XNOR U6008 ( .A(n23064), .B(n23348), .Z(n23068) );
  XNOR U6009 ( .A(n7022), .B(n7337), .Z(n7026) );
  XNOR U6010 ( .A(n6262), .B(n6598), .Z(n6266) );
  XNOR U6011 ( .A(n5497), .B(n5858), .Z(n5502) );
  XNOR U6012 ( .A(n8166), .B(n8448), .Z(n8170) );
  XNOR U6013 ( .A(n16449), .B(n16723), .Z(n16444) );
  XNOR U6014 ( .A(n20125), .B(n20403), .Z(n20129) );
  XNOR U6015 ( .A(n20861), .B(n21139), .Z(n20865) );
  XNOR U6016 ( .A(n17186), .B(n17458), .Z(n17194) );
  XNOR U6017 ( .A(n17922), .B(n18194), .Z(n17926) );
  XNOR U6018 ( .A(n21602), .B(n21874), .Z(n21606) );
  XNOR U6019 ( .A(n22338), .B(n22610), .Z(n22342) );
  XNOR U6020 ( .A(n29082), .B(n29354), .Z(n29086) );
  XNOR U6021 ( .A(n28518), .B(n28790), .Z(n28522) );
  XNOR U6022 ( .A(n27930), .B(n28202), .Z(n27934) );
  XNOR U6023 ( .A(n27318), .B(n27590), .Z(n27322) );
  XNOR U6024 ( .A(n26682), .B(n26954), .Z(n26686) );
  XNOR U6025 ( .A(n26022), .B(n26294), .Z(n26026) );
  XNOR U6026 ( .A(n25338), .B(n25610), .Z(n25342) );
  XNOR U6027 ( .A(n24630), .B(n24902), .Z(n24634) );
  XNOR U6028 ( .A(n23895), .B(n24167), .Z(n23899) );
  XNOR U6029 ( .A(n9288), .B(n9561), .Z(n9292) );
  XNOR U6030 ( .A(n10040), .B(n10446), .Z(n10044) );
  XNOR U6031 ( .A(n10565), .B(n10830), .Z(n10569) );
  XNOR U6032 ( .A(n10933), .B(n11199), .Z(n10937) );
  XNOR U6033 ( .A(n11302), .B(n11568), .Z(n11306) );
  XNOR U6034 ( .A(n12044), .B(n11673), .Z(n11675) );
  XNOR U6035 ( .A(n12412), .B(n12041), .Z(n12043) );
  XNOR U6036 ( .A(n12780), .B(n12409), .Z(n12411) );
  XNOR U6037 ( .A(n13148), .B(n12777), .Z(n12779) );
  XNOR U6038 ( .A(n13516), .B(n13145), .Z(n13147) );
  XNOR U6039 ( .A(n13884), .B(n13513), .Z(n13515) );
  XNOR U6040 ( .A(n14252), .B(n13881), .Z(n13883) );
  XNOR U6041 ( .A(n14620), .B(n14249), .Z(n14251) );
  XNOR U6042 ( .A(n14988), .B(n14617), .Z(n14619) );
  XNOR U6043 ( .A(n15356), .B(n14985), .Z(n14987) );
  XNOR U6044 ( .A(n15724), .B(n15353), .Z(n15355) );
  XNOR U6045 ( .A(n16092), .B(n15721), .Z(n15723) );
  XNOR U6046 ( .A(n16460), .B(n16089), .Z(n16091) );
  XNOR U6047 ( .A(n16828), .B(n16457), .Z(n16459) );
  XNOR U6048 ( .A(n17196), .B(n16825), .Z(n16827) );
  XNOR U6049 ( .A(n18663), .B(n18929), .Z(n18667) );
  XNOR U6050 ( .A(n19399), .B(n19665), .Z(n19403) );
  XNOR U6051 ( .A(n23079), .B(n23345), .Z(n23083) );
  XNOR U6052 ( .A(n7037), .B(n7334), .Z(n7041) );
  XNOR U6053 ( .A(n6277), .B(n6595), .Z(n6281) );
  XNOR U6054 ( .A(n5513), .B(n5855), .Z(n5517) );
  XNOR U6055 ( .A(n8181), .B(n8445), .Z(n8185) );
  XNOR U6056 ( .A(n8925), .B(n9185), .Z(n8929) );
  XNOR U6057 ( .A(n20140), .B(n20400), .Z(n20144) );
  XNOR U6058 ( .A(n20876), .B(n21136), .Z(n20880) );
  XNOR U6059 ( .A(n4752), .B(n5114), .Z(n4757) );
  XNOR U6060 ( .A(n17941), .B(n18191), .Z(n17936) );
  XNOR U6061 ( .A(n21617), .B(n21871), .Z(n21621) );
  XNOR U6062 ( .A(n22353), .B(n22607), .Z(n22357) );
  XNOR U6063 ( .A(n29637), .B(n29891), .Z(n29641) );
  XNOR U6064 ( .A(n29097), .B(n29351), .Z(n29101) );
  XNOR U6065 ( .A(n28533), .B(n28787), .Z(n28537) );
  XNOR U6066 ( .A(n27945), .B(n28199), .Z(n27949) );
  XNOR U6067 ( .A(n27333), .B(n27587), .Z(n27337) );
  XNOR U6068 ( .A(n26697), .B(n26951), .Z(n26701) );
  XNOR U6069 ( .A(n26037), .B(n26291), .Z(n26041) );
  XNOR U6070 ( .A(n25353), .B(n25607), .Z(n25357) );
  XNOR U6071 ( .A(n24645), .B(n24899), .Z(n24649) );
  XNOR U6072 ( .A(n23910), .B(n24164), .Z(n23914) );
  XNOR U6073 ( .A(n7432), .B(n7702), .Z(n7436) );
  XNOR U6074 ( .A(n10055), .B(n10440), .Z(n10059) );
  XNOR U6075 ( .A(n10580), .B(n10827), .Z(n10584) );
  XNOR U6076 ( .A(n10948), .B(n11196), .Z(n10952) );
  XNOR U6077 ( .A(n11317), .B(n11565), .Z(n11321) );
  XNOR U6078 ( .A(n12059), .B(n11688), .Z(n11690) );
  XNOR U6079 ( .A(n12427), .B(n12056), .Z(n12058) );
  XNOR U6080 ( .A(n12795), .B(n12424), .Z(n12426) );
  XNOR U6081 ( .A(n13163), .B(n12792), .Z(n12794) );
  XNOR U6082 ( .A(n13531), .B(n13160), .Z(n13162) );
  XNOR U6083 ( .A(n13899), .B(n13528), .Z(n13530) );
  XNOR U6084 ( .A(n14267), .B(n13896), .Z(n13898) );
  XNOR U6085 ( .A(n14635), .B(n14264), .Z(n14266) );
  XNOR U6086 ( .A(n15003), .B(n14632), .Z(n14634) );
  XNOR U6087 ( .A(n15371), .B(n15000), .Z(n15002) );
  XNOR U6088 ( .A(n15739), .B(n15368), .Z(n15370) );
  XNOR U6089 ( .A(n16107), .B(n15736), .Z(n15738) );
  XNOR U6090 ( .A(n16475), .B(n16104), .Z(n16106) );
  XNOR U6091 ( .A(n16843), .B(n16472), .Z(n16474) );
  XNOR U6092 ( .A(n17211), .B(n16840), .Z(n16842) );
  XNOR U6093 ( .A(n17579), .B(n17208), .Z(n17210) );
  XNOR U6094 ( .A(n17947), .B(n17576), .Z(n17578) );
  XNOR U6095 ( .A(n18315), .B(n17944), .Z(n17946) );
  XNOR U6096 ( .A(n18678), .B(n18926), .Z(n18686) );
  XNOR U6097 ( .A(n19414), .B(n19662), .Z(n19418) );
  XNOR U6098 ( .A(n23094), .B(n23342), .Z(n23098) );
  XNOR U6099 ( .A(n6674), .B(n6958), .Z(n6678) );
  XNOR U6100 ( .A(n5910), .B(n6222), .Z(n5914) );
  XNOR U6101 ( .A(n5146), .B(n5482), .Z(n5150) );
  XNOR U6102 ( .A(n8196), .B(n8442), .Z(n8200) );
  XNOR U6103 ( .A(n8940), .B(n9182), .Z(n8944) );
  XNOR U6104 ( .A(n9683), .B(n9934), .Z(n9687) );
  XNOR U6105 ( .A(n20155), .B(n20397), .Z(n20159) );
  XNOR U6106 ( .A(n20891), .B(n21133), .Z(n20895) );
  XNOR U6107 ( .A(n4386), .B(n4740), .Z(n4390) );
  XNOR U6108 ( .A(n21632), .B(n21868), .Z(n21636) );
  XNOR U6109 ( .A(n22368), .B(n22604), .Z(n22372) );
  XNOR U6110 ( .A(n30660), .B(n30896), .Z(n30664) );
  XNOR U6111 ( .A(n30168), .B(n30404), .Z(n30172) );
  XNOR U6112 ( .A(n29652), .B(n29888), .Z(n29656) );
  XNOR U6113 ( .A(n29112), .B(n29348), .Z(n29116) );
  XNOR U6114 ( .A(n28548), .B(n28784), .Z(n28552) );
  XNOR U6115 ( .A(n27960), .B(n28196), .Z(n27964) );
  XNOR U6116 ( .A(n27348), .B(n27584), .Z(n27352) );
  XNOR U6117 ( .A(n26712), .B(n26948), .Z(n26716) );
  XNOR U6118 ( .A(n26052), .B(n26288), .Z(n26056) );
  XNOR U6119 ( .A(n25368), .B(n25604), .Z(n25372) );
  XNOR U6120 ( .A(n24660), .B(n24896), .Z(n24664) );
  XNOR U6121 ( .A(n23925), .B(n24161), .Z(n23929) );
  XNOR U6122 ( .A(n7447), .B(n7699), .Z(n7451) );
  XNOR U6123 ( .A(n10963), .B(n11193), .Z(n10967) );
  XNOR U6124 ( .A(n11332), .B(n11562), .Z(n11336) );
  XNOR U6125 ( .A(n12074), .B(n11703), .Z(n11705) );
  XNOR U6126 ( .A(n12442), .B(n12071), .Z(n12073) );
  XNOR U6127 ( .A(n12810), .B(n12439), .Z(n12441) );
  XNOR U6128 ( .A(n13178), .B(n12807), .Z(n12809) );
  XNOR U6129 ( .A(n13546), .B(n13175), .Z(n13177) );
  XNOR U6130 ( .A(n13914), .B(n13543), .Z(n13545) );
  XNOR U6131 ( .A(n14282), .B(n13911), .Z(n13913) );
  XNOR U6132 ( .A(n14650), .B(n14279), .Z(n14281) );
  XNOR U6133 ( .A(n15018), .B(n14647), .Z(n14649) );
  XNOR U6134 ( .A(n15386), .B(n15015), .Z(n15017) );
  XNOR U6135 ( .A(n15754), .B(n15383), .Z(n15385) );
  XNOR U6136 ( .A(n16122), .B(n15751), .Z(n15753) );
  XNOR U6137 ( .A(n16490), .B(n16119), .Z(n16121) );
  XNOR U6138 ( .A(n16858), .B(n16487), .Z(n16489) );
  XNOR U6139 ( .A(n17226), .B(n16855), .Z(n16857) );
  XNOR U6140 ( .A(n17594), .B(n17223), .Z(n17225) );
  XNOR U6141 ( .A(n17962), .B(n17591), .Z(n17593) );
  XNOR U6142 ( .A(n18330), .B(n17959), .Z(n17961) );
  XNOR U6143 ( .A(n18698), .B(n18327), .Z(n18329) );
  XNOR U6144 ( .A(n19066), .B(n18695), .Z(n18697) );
  XNOR U6145 ( .A(n19434), .B(n19063), .Z(n19065) );
  XNOR U6146 ( .A(n19433), .B(n19659), .Z(n19428) );
  XNOR U6147 ( .A(n23109), .B(n23339), .Z(n23113) );
  XNOR U6148 ( .A(n6689), .B(n6955), .Z(n6693) );
  XNOR U6149 ( .A(n5925), .B(n6219), .Z(n5929) );
  XNOR U6150 ( .A(n5161), .B(n5479), .Z(n5165) );
  XNOR U6151 ( .A(n8583), .B(n8811), .Z(n8587) );
  XNOR U6152 ( .A(n9323), .B(n9554), .Z(n9327) );
  XNOR U6153 ( .A(n10075), .B(n10432), .Z(n10079) );
  XNOR U6154 ( .A(n10600), .B(n10823), .Z(n10604) );
  XNOR U6155 ( .A(n20170), .B(n20394), .Z(n20178) );
  XNOR U6156 ( .A(n20906), .B(n21130), .Z(n20910) );
  XNOR U6157 ( .A(n4401), .B(n4737), .Z(n4405) );
  XNOR U6158 ( .A(n3636), .B(n3997), .Z(n3641) );
  XNOR U6159 ( .A(n21647), .B(n21865), .Z(n21651) );
  XNOR U6160 ( .A(n22383), .B(n22601), .Z(n22387) );
  XNOR U6161 ( .A(n31143), .B(n31361), .Z(n31147) );
  XNOR U6162 ( .A(n30675), .B(n30893), .Z(n30679) );
  XNOR U6163 ( .A(n30183), .B(n30401), .Z(n30187) );
  XNOR U6164 ( .A(n29667), .B(n29885), .Z(n29671) );
  XNOR U6165 ( .A(n29127), .B(n29345), .Z(n29131) );
  XNOR U6166 ( .A(n28563), .B(n28781), .Z(n28567) );
  XNOR U6167 ( .A(n27975), .B(n28193), .Z(n27979) );
  XNOR U6168 ( .A(n27363), .B(n27581), .Z(n27367) );
  XNOR U6169 ( .A(n26727), .B(n26945), .Z(n26731) );
  XNOR U6170 ( .A(n26067), .B(n26285), .Z(n26071) );
  XNOR U6171 ( .A(n25383), .B(n25601), .Z(n25387) );
  XNOR U6172 ( .A(n24675), .B(n24893), .Z(n24679) );
  XNOR U6173 ( .A(n23940), .B(n24158), .Z(n23944) );
  XNOR U6174 ( .A(n7462), .B(n7696), .Z(n7466) );
  XNOR U6175 ( .A(n12089), .B(n11718), .Z(n11720) );
  XNOR U6176 ( .A(n12457), .B(n12086), .Z(n12088) );
  XNOR U6177 ( .A(n12825), .B(n12454), .Z(n12456) );
  XNOR U6178 ( .A(n13193), .B(n12822), .Z(n12824) );
  XNOR U6179 ( .A(n13561), .B(n13190), .Z(n13192) );
  XNOR U6180 ( .A(n13929), .B(n13558), .Z(n13560) );
  XNOR U6181 ( .A(n14297), .B(n13926), .Z(n13928) );
  XNOR U6182 ( .A(n14665), .B(n14294), .Z(n14296) );
  XNOR U6183 ( .A(n15033), .B(n14662), .Z(n14664) );
  XNOR U6184 ( .A(n15401), .B(n15030), .Z(n15032) );
  XNOR U6185 ( .A(n15769), .B(n15398), .Z(n15400) );
  XNOR U6186 ( .A(n16137), .B(n15766), .Z(n15768) );
  XNOR U6187 ( .A(n16505), .B(n16134), .Z(n16136) );
  XNOR U6188 ( .A(n16873), .B(n16502), .Z(n16504) );
  XNOR U6189 ( .A(n17241), .B(n16870), .Z(n16872) );
  XNOR U6190 ( .A(n17609), .B(n17238), .Z(n17240) );
  XNOR U6191 ( .A(n17977), .B(n17606), .Z(n17608) );
  XNOR U6192 ( .A(n18345), .B(n17974), .Z(n17976) );
  XNOR U6193 ( .A(n18713), .B(n18342), .Z(n18344) );
  XNOR U6194 ( .A(n19081), .B(n18710), .Z(n18712) );
  XNOR U6195 ( .A(n19449), .B(n19078), .Z(n19080) );
  XNOR U6196 ( .A(n19817), .B(n19446), .Z(n19448) );
  XNOR U6197 ( .A(n20185), .B(n19814), .Z(n19816) );
  XNOR U6198 ( .A(n20553), .B(n20182), .Z(n20184) );
  XNOR U6199 ( .A(n23124), .B(n23336), .Z(n23128) );
  XNOR U6200 ( .A(n6704), .B(n6952), .Z(n6708) );
  XNOR U6201 ( .A(n5940), .B(n6216), .Z(n5944) );
  XNOR U6202 ( .A(n5176), .B(n5476), .Z(n5180) );
  XNOR U6203 ( .A(n7856), .B(n8063), .Z(n7857) );
  XNOR U6204 ( .A(n8598), .B(n8808), .Z(n8606) );
  XNOR U6205 ( .A(n9338), .B(n9551), .Z(n9342) );
  XNOR U6206 ( .A(n10090), .B(n10426), .Z(n10094) );
  XNOR U6207 ( .A(n10615), .B(n10820), .Z(n10619) );
  XNOR U6208 ( .A(n10983), .B(n11189), .Z(n10987) );
  XNOR U6209 ( .A(n11352), .B(n11558), .Z(n11356) );
  XNOR U6210 ( .A(n12094), .B(n11723), .Z(n11725) );
  XNOR U6211 ( .A(n20925), .B(n21127), .Z(n20920) );
  XNOR U6212 ( .A(n4416), .B(n4734), .Z(n4420) );
  XNOR U6213 ( .A(n3652), .B(n3994), .Z(n3656) );
  XNOR U6214 ( .A(n21662), .B(n21862), .Z(n21670) );
  XNOR U6215 ( .A(n22398), .B(n22598), .Z(n22402) );
  XNOR U6216 ( .A(n32185), .B(n32377), .Z(n32189) );
  XNOR U6217 ( .A(n31602), .B(n31973), .Z(n31606) );
  XNOR U6218 ( .A(n31158), .B(n31358), .Z(n31162) );
  XNOR U6219 ( .A(n30690), .B(n30890), .Z(n30694) );
  XNOR U6220 ( .A(n30198), .B(n30398), .Z(n30202) );
  XNOR U6221 ( .A(n29682), .B(n29882), .Z(n29686) );
  XNOR U6222 ( .A(n29142), .B(n29342), .Z(n29146) );
  XNOR U6223 ( .A(n28578), .B(n28778), .Z(n28582) );
  XNOR U6224 ( .A(n27990), .B(n28190), .Z(n27994) );
  XNOR U6225 ( .A(n27378), .B(n27578), .Z(n27382) );
  XNOR U6226 ( .A(n26742), .B(n26942), .Z(n26746) );
  XNOR U6227 ( .A(n26082), .B(n26282), .Z(n26086) );
  XNOR U6228 ( .A(n25398), .B(n25598), .Z(n25402) );
  XNOR U6229 ( .A(n24690), .B(n24890), .Z(n24694) );
  XNOR U6230 ( .A(n23955), .B(n24155), .Z(n23959) );
  XNOR U6231 ( .A(n7096), .B(n7323), .Z(n7091) );
  XNOR U6232 ( .A(n2892), .B(n3253), .Z(n2897) );
  XNOR U6233 ( .A(n13208), .B(n12837), .Z(n12839) );
  XNOR U6234 ( .A(n13576), .B(n13205), .Z(n13207) );
  XNOR U6235 ( .A(n13944), .B(n13573), .Z(n13575) );
  XNOR U6236 ( .A(n14312), .B(n13941), .Z(n13943) );
  XNOR U6237 ( .A(n14680), .B(n14309), .Z(n14311) );
  XNOR U6238 ( .A(n15048), .B(n14677), .Z(n14679) );
  XNOR U6239 ( .A(n15416), .B(n15045), .Z(n15047) );
  XNOR U6240 ( .A(n15784), .B(n15413), .Z(n15415) );
  XNOR U6241 ( .A(n16152), .B(n15781), .Z(n15783) );
  XNOR U6242 ( .A(n16520), .B(n16149), .Z(n16151) );
  XNOR U6243 ( .A(n16888), .B(n16517), .Z(n16519) );
  XNOR U6244 ( .A(n17256), .B(n16885), .Z(n16887) );
  XNOR U6245 ( .A(n17624), .B(n17253), .Z(n17255) );
  XNOR U6246 ( .A(n17992), .B(n17621), .Z(n17623) );
  XNOR U6247 ( .A(n18360), .B(n17989), .Z(n17991) );
  XNOR U6248 ( .A(n18728), .B(n18357), .Z(n18359) );
  XNOR U6249 ( .A(n19096), .B(n18725), .Z(n18727) );
  XNOR U6250 ( .A(n19464), .B(n19093), .Z(n19095) );
  XNOR U6251 ( .A(n19832), .B(n19461), .Z(n19463) );
  XNOR U6252 ( .A(n20200), .B(n19829), .Z(n19831) );
  XNOR U6253 ( .A(n20568), .B(n20197), .Z(n20199) );
  XNOR U6254 ( .A(n20936), .B(n20565), .Z(n20567) );
  XNOR U6255 ( .A(n21304), .B(n20933), .Z(n20935) );
  XNOR U6256 ( .A(n21672), .B(n21301), .Z(n21303) );
  XNOR U6257 ( .A(n23139), .B(n23333), .Z(n23143) );
  XNOR U6258 ( .A(n6738), .B(n6944), .Z(n6742) );
  XNOR U6259 ( .A(n6337), .B(n6583), .Z(n6345) );
  XNOR U6260 ( .A(n5573), .B(n5843), .Z(n5577) );
  XNOR U6261 ( .A(n4808), .B(n5103), .Z(n4812) );
  XNOR U6262 ( .A(n7868), .B(n8060), .Z(n7872) );
  XNOR U6263 ( .A(n8612), .B(n8804), .Z(n8616) );
  XNOR U6264 ( .A(n9357), .B(n9548), .Z(n9352) );
  XNOR U6265 ( .A(n10105), .B(n10420), .Z(n10109) );
  XNOR U6266 ( .A(n10630), .B(n10817), .Z(n10634) );
  XNOR U6267 ( .A(n10998), .B(n11186), .Z(n11002) );
  XNOR U6268 ( .A(n11367), .B(n11555), .Z(n11371) );
  XNOR U6269 ( .A(n12109), .B(n11738), .Z(n11740) );
  XNOR U6270 ( .A(n12477), .B(n12106), .Z(n12108) );
  XNOR U6271 ( .A(n12845), .B(n12474), .Z(n12476) );
  XNOR U6272 ( .A(n13213), .B(n12842), .Z(n12844) );
  XNOR U6273 ( .A(n5979), .B(n6207), .Z(n5983) );
  XNOR U6274 ( .A(n4049), .B(n4361), .Z(n4053) );
  XNOR U6275 ( .A(n3285), .B(n3621), .Z(n3289) );
  XNOR U6276 ( .A(n22417), .B(n22595), .Z(n22412) );
  XNOR U6277 ( .A(n32583), .B(n32757), .Z(n32587) );
  XNOR U6278 ( .A(n32200), .B(n32374), .Z(n32204) );
  XNOR U6279 ( .A(n31617), .B(n31970), .Z(n31621) );
  XNOR U6280 ( .A(n31173), .B(n31355), .Z(n31177) );
  XNOR U6281 ( .A(n30705), .B(n30887), .Z(n30709) );
  XNOR U6282 ( .A(n30213), .B(n30395), .Z(n30217) );
  XNOR U6283 ( .A(n29697), .B(n29879), .Z(n29701) );
  XNOR U6284 ( .A(n29157), .B(n29339), .Z(n29161) );
  XNOR U6285 ( .A(n28593), .B(n28775), .Z(n28597) );
  XNOR U6286 ( .A(n28005), .B(n28187), .Z(n28009) );
  XNOR U6287 ( .A(n27393), .B(n27575), .Z(n27397) );
  XNOR U6288 ( .A(n26757), .B(n26939), .Z(n26761) );
  XNOR U6289 ( .A(n26097), .B(n26279), .Z(n26101) );
  XNOR U6290 ( .A(n25413), .B(n25595), .Z(n25417) );
  XNOR U6291 ( .A(n24705), .B(n24887), .Z(n24709) );
  XNOR U6292 ( .A(n23970), .B(n24152), .Z(n23974) );
  XNOR U6293 ( .A(n2525), .B(n2880), .Z(n2529) );
  XNOR U6294 ( .A(n5626), .B(n5830), .Z(n5630) );
  XNOR U6295 ( .A(n6390), .B(n6570), .Z(n6394) );
  XNOR U6296 ( .A(n14327), .B(n13956), .Z(n13958) );
  XNOR U6297 ( .A(n14695), .B(n14324), .Z(n14326) );
  XNOR U6298 ( .A(n15063), .B(n14692), .Z(n14694) );
  XNOR U6299 ( .A(n15431), .B(n15060), .Z(n15062) );
  XNOR U6300 ( .A(n15799), .B(n15428), .Z(n15430) );
  XNOR U6301 ( .A(n16167), .B(n15796), .Z(n15798) );
  XNOR U6302 ( .A(n16535), .B(n16164), .Z(n16166) );
  XNOR U6303 ( .A(n16903), .B(n16532), .Z(n16534) );
  XNOR U6304 ( .A(n17271), .B(n16900), .Z(n16902) );
  XNOR U6305 ( .A(n17639), .B(n17268), .Z(n17270) );
  XNOR U6306 ( .A(n18007), .B(n17636), .Z(n17638) );
  XNOR U6307 ( .A(n18375), .B(n18004), .Z(n18006) );
  XNOR U6308 ( .A(n18743), .B(n18372), .Z(n18374) );
  XNOR U6309 ( .A(n19111), .B(n18740), .Z(n18742) );
  XNOR U6310 ( .A(n19479), .B(n19108), .Z(n19110) );
  XNOR U6311 ( .A(n19847), .B(n19476), .Z(n19478) );
  XNOR U6312 ( .A(n20215), .B(n19844), .Z(n19846) );
  XNOR U6313 ( .A(n20583), .B(n20212), .Z(n20214) );
  XNOR U6314 ( .A(n20951), .B(n20580), .Z(n20582) );
  XNOR U6315 ( .A(n21319), .B(n20948), .Z(n20950) );
  XNOR U6316 ( .A(n21687), .B(n21316), .Z(n21318) );
  XNOR U6317 ( .A(n22055), .B(n21684), .Z(n21686) );
  XNOR U6318 ( .A(n22423), .B(n22052), .Z(n22054) );
  XNOR U6319 ( .A(n22791), .B(n22420), .Z(n22422) );
  XNOR U6320 ( .A(n23154), .B(n23330), .Z(n23162) );
  XNOR U6321 ( .A(n6375), .B(n6575), .Z(n6370) );
  XNOR U6322 ( .A(n5592), .B(n5840), .Z(n5587) );
  XNOR U6323 ( .A(n4823), .B(n5100), .Z(n4827) );
  XNOR U6324 ( .A(n7135), .B(n7312), .Z(n7139) );
  XNOR U6325 ( .A(n7885), .B(n8056), .Z(n7886) );
  XNOR U6326 ( .A(n8627), .B(n8801), .Z(n8635) );
  XNOR U6327 ( .A(n9367), .B(n9544), .Z(n9371) );
  XNOR U6328 ( .A(n10114), .B(n10415), .Z(n10123) );
  XNOR U6329 ( .A(n10645), .B(n10814), .Z(n10649) );
  XNOR U6330 ( .A(n11013), .B(n11183), .Z(n11017) );
  XNOR U6331 ( .A(n11382), .B(n11552), .Z(n11386) );
  XNOR U6332 ( .A(n12124), .B(n11753), .Z(n11755) );
  XNOR U6333 ( .A(n12492), .B(n12121), .Z(n12123) );
  XNOR U6334 ( .A(n12860), .B(n12489), .Z(n12491) );
  XNOR U6335 ( .A(n13228), .B(n12857), .Z(n12859) );
  XNOR U6336 ( .A(n13596), .B(n13225), .Z(n13227) );
  XNOR U6337 ( .A(n13964), .B(n13593), .Z(n13595) );
  XNOR U6338 ( .A(n14332), .B(n13961), .Z(n13963) );
  XNOR U6339 ( .A(n5612), .B(n5834), .Z(n5620) );
  XNOR U6340 ( .A(n4847), .B(n5094), .Z(n4851) );
  XNOR U6341 ( .A(n4064), .B(n4358), .Z(n4068) );
  XNOR U6342 ( .A(n3300), .B(n3618), .Z(n3304) );
  XNOR U6343 ( .A(n33289), .B(n33445), .Z(n33293) );
  XNOR U6344 ( .A(n32954), .B(n33113), .Z(n32958) );
  XNOR U6345 ( .A(n32598), .B(n32754), .Z(n32602) );
  XNOR U6346 ( .A(n32215), .B(n32371), .Z(n32219) );
  XNOR U6347 ( .A(n31632), .B(n31967), .Z(n31636) );
  XNOR U6348 ( .A(n31188), .B(n31352), .Z(n31192) );
  XNOR U6349 ( .A(n30720), .B(n30884), .Z(n30724) );
  XNOR U6350 ( .A(n30228), .B(n30392), .Z(n30232) );
  XNOR U6351 ( .A(n29712), .B(n29876), .Z(n29716) );
  XNOR U6352 ( .A(n29172), .B(n29336), .Z(n29176) );
  XNOR U6353 ( .A(n28608), .B(n28772), .Z(n28612) );
  XNOR U6354 ( .A(n28020), .B(n28184), .Z(n28024) );
  XNOR U6355 ( .A(n27408), .B(n27572), .Z(n27412) );
  XNOR U6356 ( .A(n26772), .B(n26936), .Z(n26776) );
  XNOR U6357 ( .A(n26112), .B(n26276), .Z(n26116) );
  XNOR U6358 ( .A(n25428), .B(n25592), .Z(n25432) );
  XNOR U6359 ( .A(n24720), .B(n24884), .Z(n24724) );
  XNOR U6360 ( .A(n23985), .B(n24149), .Z(n23989) );
  XNOR U6361 ( .A(n2540), .B(n2877), .Z(n2544) );
  XNOR U6362 ( .A(n1774), .B(n2135), .Z(n1779) );
  XNOR U6363 ( .A(n6027), .B(n6197), .Z(n6022) );
  XNOR U6364 ( .A(n5259), .B(n5457), .Z(n5263) );
  XNOR U6365 ( .A(n4494), .B(n4716), .Z(n4498) );
  XNOR U6366 ( .A(n15446), .B(n15075), .Z(n15077) );
  XNOR U6367 ( .A(n15814), .B(n15443), .Z(n15445) );
  XNOR U6368 ( .A(n16182), .B(n15811), .Z(n15813) );
  XNOR U6369 ( .A(n16550), .B(n16179), .Z(n16181) );
  XNOR U6370 ( .A(n16918), .B(n16547), .Z(n16549) );
  XNOR U6371 ( .A(n17286), .B(n16915), .Z(n16917) );
  XNOR U6372 ( .A(n17654), .B(n17283), .Z(n17285) );
  XNOR U6373 ( .A(n18022), .B(n17651), .Z(n17653) );
  XNOR U6374 ( .A(n18390), .B(n18019), .Z(n18021) );
  XNOR U6375 ( .A(n18758), .B(n18387), .Z(n18389) );
  XNOR U6376 ( .A(n19126), .B(n18755), .Z(n18757) );
  XNOR U6377 ( .A(n19494), .B(n19123), .Z(n19125) );
  XNOR U6378 ( .A(n19862), .B(n19491), .Z(n19493) );
  XNOR U6379 ( .A(n20230), .B(n19859), .Z(n19861) );
  XNOR U6380 ( .A(n20598), .B(n20227), .Z(n20229) );
  XNOR U6381 ( .A(n20966), .B(n20595), .Z(n20597) );
  XNOR U6382 ( .A(n21334), .B(n20963), .Z(n20965) );
  XNOR U6383 ( .A(n21702), .B(n21331), .Z(n21333) );
  XNOR U6384 ( .A(n22070), .B(n21699), .Z(n21701) );
  XNOR U6385 ( .A(n22438), .B(n22067), .Z(n22069) );
  XNOR U6386 ( .A(n22806), .B(n22435), .Z(n22437) );
  XNOR U6387 ( .A(n23174), .B(n22803), .Z(n22805) );
  XNOR U6388 ( .A(n23168), .B(n23326), .Z(n23172) );
  XNOR U6389 ( .A(n4460), .B(n4726), .Z(n4455) );
  XNOR U6390 ( .A(n6409), .B(n6565), .Z(n6413) );
  XNOR U6391 ( .A(n7154), .B(n7309), .Z(n7149) );
  XNOR U6392 ( .A(n7897), .B(n8053), .Z(n7901) );
  XNOR U6393 ( .A(n8641), .B(n8797), .Z(n8645) );
  XNOR U6394 ( .A(n9386), .B(n9541), .Z(n9381) );
  XNOR U6395 ( .A(n10134), .B(n10409), .Z(n10138) );
  XNOR U6396 ( .A(n10660), .B(n10811), .Z(n10664) );
  XNOR U6397 ( .A(n11028), .B(n11180), .Z(n11032) );
  XNOR U6398 ( .A(n11397), .B(n11549), .Z(n11401) );
  XNOR U6399 ( .A(n12139), .B(n11768), .Z(n11770) );
  XNOR U6400 ( .A(n12507), .B(n12136), .Z(n12138) );
  XNOR U6401 ( .A(n12875), .B(n12504), .Z(n12506) );
  XNOR U6402 ( .A(n13243), .B(n12872), .Z(n12874) );
  XNOR U6403 ( .A(n13611), .B(n13240), .Z(n13242) );
  XNOR U6404 ( .A(n13979), .B(n13608), .Z(n13610) );
  XNOR U6405 ( .A(n14347), .B(n13976), .Z(n13978) );
  XNOR U6406 ( .A(n14715), .B(n14344), .Z(n14346) );
  XNOR U6407 ( .A(n15083), .B(n14712), .Z(n14714) );
  XNOR U6408 ( .A(n15451), .B(n15080), .Z(n15082) );
  XNOR U6409 ( .A(n5288), .B(n5450), .Z(n5292) );
  XNOR U6410 ( .A(n4523), .B(n4709), .Z(n4527) );
  XNOR U6411 ( .A(n4866), .B(n5091), .Z(n4861) );
  XNOR U6412 ( .A(n4098), .B(n4350), .Z(n4102) );
  XNOR U6413 ( .A(n3334), .B(n3610), .Z(n3338) );
  XNOR U6414 ( .A(n3697), .B(n3985), .Z(n3705) );
  XNOR U6415 ( .A(n2933), .B(n3245), .Z(n2937) );
  XNOR U6416 ( .A(n33615), .B(n33753), .Z(n33619) );
  XNOR U6417 ( .A(n33304), .B(n33442), .Z(n33308) );
  XNOR U6418 ( .A(n32969), .B(n33110), .Z(n32973) );
  XNOR U6419 ( .A(n32613), .B(n32751), .Z(n32617) );
  XNOR U6420 ( .A(n32230), .B(n32368), .Z(n32234) );
  XNOR U6421 ( .A(n31647), .B(n31964), .Z(n31651) );
  XNOR U6422 ( .A(n31203), .B(n31349), .Z(n31207) );
  XNOR U6423 ( .A(n30735), .B(n30881), .Z(n30739) );
  XNOR U6424 ( .A(n30243), .B(n30389), .Z(n30247) );
  XNOR U6425 ( .A(n29727), .B(n29873), .Z(n29731) );
  XNOR U6426 ( .A(n29187), .B(n29333), .Z(n29191) );
  XNOR U6427 ( .A(n28623), .B(n28769), .Z(n28627) );
  XNOR U6428 ( .A(n28035), .B(n28181), .Z(n28039) );
  XNOR U6429 ( .A(n27423), .B(n27569), .Z(n27427) );
  XNOR U6430 ( .A(n26787), .B(n26933), .Z(n26791) );
  XNOR U6431 ( .A(n26127), .B(n26273), .Z(n26131) );
  XNOR U6432 ( .A(n25443), .B(n25589), .Z(n25447) );
  XNOR U6433 ( .A(n24735), .B(n24881), .Z(n24739) );
  XNOR U6434 ( .A(n24000), .B(n24146), .Z(n24004) );
  XNOR U6435 ( .A(n2172), .B(n2503), .Z(n2176) );
  XNOR U6436 ( .A(n1408), .B(n1762), .Z(n1412) );
  XNOR U6437 ( .A(n4895), .B(n5084), .Z(n4890) );
  XNOR U6438 ( .A(n4127), .B(n4343), .Z(n4131) );
  XNOR U6439 ( .A(n3363), .B(n3603), .Z(n3367) );
  XNOR U6440 ( .A(n4552), .B(n4702), .Z(n4556) );
  XNOR U6441 ( .A(n16565), .B(n16194), .Z(n16196) );
  XNOR U6442 ( .A(n16933), .B(n16562), .Z(n16564) );
  XNOR U6443 ( .A(n17301), .B(n16930), .Z(n16932) );
  XNOR U6444 ( .A(n17669), .B(n17298), .Z(n17300) );
  XNOR U6445 ( .A(n18037), .B(n17666), .Z(n17668) );
  XNOR U6446 ( .A(n18405), .B(n18034), .Z(n18036) );
  XNOR U6447 ( .A(n18773), .B(n18402), .Z(n18404) );
  XNOR U6448 ( .A(n19141), .B(n18770), .Z(n18772) );
  XNOR U6449 ( .A(n19509), .B(n19138), .Z(n19140) );
  XNOR U6450 ( .A(n19877), .B(n19506), .Z(n19508) );
  XNOR U6451 ( .A(n20245), .B(n19874), .Z(n19876) );
  XNOR U6452 ( .A(n20613), .B(n20242), .Z(n20244) );
  XNOR U6453 ( .A(n20981), .B(n20610), .Z(n20612) );
  XNOR U6454 ( .A(n21349), .B(n20978), .Z(n20980) );
  XNOR U6455 ( .A(n21717), .B(n21346), .Z(n21348) );
  XNOR U6456 ( .A(n22085), .B(n21714), .Z(n21716) );
  XNOR U6457 ( .A(n22453), .B(n22082), .Z(n22084) );
  XNOR U6458 ( .A(n22821), .B(n22450), .Z(n22452) );
  XNOR U6459 ( .A(n23189), .B(n22818), .Z(n22820) );
  XNOR U6460 ( .A(n23183), .B(n23323), .Z(n23187) );
  XNOR U6461 ( .A(n6424), .B(n6562), .Z(n6432) );
  XNOR U6462 ( .A(n7164), .B(n7305), .Z(n7168) );
  XNOR U6463 ( .A(n7914), .B(n8049), .Z(n7915) );
  XNOR U6464 ( .A(n8656), .B(n8794), .Z(n8664) );
  XNOR U6465 ( .A(n9396), .B(n9537), .Z(n9400) );
  XNOR U6466 ( .A(n10143), .B(n10404), .Z(n10152) );
  XNOR U6467 ( .A(n10675), .B(n10808), .Z(n10679) );
  XNOR U6468 ( .A(n11043), .B(n11177), .Z(n11047) );
  XNOR U6469 ( .A(n11412), .B(n11546), .Z(n11416) );
  XNOR U6470 ( .A(n12154), .B(n11783), .Z(n11785) );
  XNOR U6471 ( .A(n12522), .B(n12151), .Z(n12153) );
  XNOR U6472 ( .A(n12890), .B(n12519), .Z(n12521) );
  XNOR U6473 ( .A(n13258), .B(n12887), .Z(n12889) );
  XNOR U6474 ( .A(n13626), .B(n13255), .Z(n13257) );
  XNOR U6475 ( .A(n13994), .B(n13623), .Z(n13625) );
  XNOR U6476 ( .A(n14362), .B(n13991), .Z(n13993) );
  XNOR U6477 ( .A(n14730), .B(n14359), .Z(n14361) );
  XNOR U6478 ( .A(n15098), .B(n14727), .Z(n14729) );
  XNOR U6479 ( .A(n15466), .B(n15095), .Z(n15097) );
  XNOR U6480 ( .A(n15834), .B(n15463), .Z(n15465) );
  XNOR U6481 ( .A(n16202), .B(n15831), .Z(n15833) );
  XNOR U6482 ( .A(n16570), .B(n16199), .Z(n16201) );
  XNOR U6483 ( .A(n4924), .B(n5077), .Z(n4919) );
  XNOR U6484 ( .A(n4156), .B(n4336), .Z(n4160) );
  XNOR U6485 ( .A(n3392), .B(n3596), .Z(n3396) );
  XNOR U6486 ( .A(n3735), .B(n3977), .Z(n3730) );
  XNOR U6487 ( .A(n2967), .B(n3237), .Z(n2971) );
  XNOR U6488 ( .A(n2201), .B(n2496), .Z(n2205) );
  XNOR U6489 ( .A(n2952), .B(n3242), .Z(n2947) );
  XNOR U6490 ( .A(n6059), .B(n6188), .Z(n6060) );
  XNOR U6491 ( .A(n34177), .B(n34297), .Z(n34181) );
  XNOR U6492 ( .A(n33914), .B(n34037), .Z(n33918) );
  XNOR U6493 ( .A(n33630), .B(n33750), .Z(n33634) );
  XNOR U6494 ( .A(n33319), .B(n33439), .Z(n33323) );
  XNOR U6495 ( .A(n32984), .B(n33107), .Z(n32988) );
  XNOR U6496 ( .A(n32628), .B(n32748), .Z(n32632) );
  XNOR U6497 ( .A(n32245), .B(n32365), .Z(n32249) );
  XNOR U6498 ( .A(n31662), .B(n31961), .Z(n31666) );
  XNOR U6499 ( .A(n31218), .B(n31346), .Z(n31222) );
  XNOR U6500 ( .A(n30750), .B(n30878), .Z(n30754) );
  XNOR U6501 ( .A(n30258), .B(n30386), .Z(n30262) );
  XNOR U6502 ( .A(n29742), .B(n29870), .Z(n29746) );
  XNOR U6503 ( .A(n29202), .B(n29330), .Z(n29206) );
  XNOR U6504 ( .A(n28638), .B(n28766), .Z(n28642) );
  XNOR U6505 ( .A(n28050), .B(n28178), .Z(n28054) );
  XNOR U6506 ( .A(n27438), .B(n27566), .Z(n27442) );
  XNOR U6507 ( .A(n26802), .B(n26930), .Z(n26806) );
  XNOR U6508 ( .A(n26142), .B(n26270), .Z(n26146) );
  XNOR U6509 ( .A(n25458), .B(n25586), .Z(n25462) );
  XNOR U6510 ( .A(n24750), .B(n24878), .Z(n24754) );
  XNOR U6511 ( .A(n24015), .B(n24143), .Z(n24019) );
  XNOR U6512 ( .A(n2187), .B(n2500), .Z(n2195) );
  XNOR U6513 ( .A(n1423), .B(n1759), .Z(n1427) );
  XNOR U6514 ( .A(n658), .B(n1019), .Z(n663) );
  XNOR U6515 ( .A(n3764), .B(n3970), .Z(n3759) );
  XNOR U6516 ( .A(n2996), .B(n3230), .Z(n3000) );
  XNOR U6517 ( .A(n2230), .B(n2489), .Z(n2234) );
  XNOR U6518 ( .A(n4185), .B(n4329), .Z(n4189) );
  XNOR U6519 ( .A(n3421), .B(n3589), .Z(n3425) );
  XNOR U6520 ( .A(n4944), .B(n5071), .Z(n4952) );
  XNOR U6521 ( .A(n5689), .B(n5815), .Z(n5693) );
  XNOR U6522 ( .A(n17684), .B(n17313), .Z(n17315) );
  XNOR U6523 ( .A(n18052), .B(n17681), .Z(n17683) );
  XNOR U6524 ( .A(n18420), .B(n18049), .Z(n18051) );
  XNOR U6525 ( .A(n18788), .B(n18417), .Z(n18419) );
  XNOR U6526 ( .A(n19156), .B(n18785), .Z(n18787) );
  XNOR U6527 ( .A(n19524), .B(n19153), .Z(n19155) );
  XNOR U6528 ( .A(n19892), .B(n19521), .Z(n19523) );
  XNOR U6529 ( .A(n20260), .B(n19889), .Z(n19891) );
  XNOR U6530 ( .A(n20628), .B(n20257), .Z(n20259) );
  XNOR U6531 ( .A(n20996), .B(n20625), .Z(n20627) );
  XNOR U6532 ( .A(n21364), .B(n20993), .Z(n20995) );
  XNOR U6533 ( .A(n21732), .B(n21361), .Z(n21363) );
  XNOR U6534 ( .A(n22100), .B(n21729), .Z(n21731) );
  XNOR U6535 ( .A(n22468), .B(n22097), .Z(n22099) );
  XNOR U6536 ( .A(n22836), .B(n22465), .Z(n22467) );
  XNOR U6537 ( .A(n23204), .B(n22833), .Z(n22835) );
  XNOR U6538 ( .A(n23198), .B(n23320), .Z(n23202) );
  XNOR U6539 ( .A(n7183), .B(n7302), .Z(n7178) );
  XNOR U6540 ( .A(n7926), .B(n8046), .Z(n7930) );
  XNOR U6541 ( .A(n8670), .B(n8790), .Z(n8674) );
  XNOR U6542 ( .A(n9415), .B(n9534), .Z(n9410) );
  XNOR U6543 ( .A(n10163), .B(n10398), .Z(n10167) );
  XNOR U6544 ( .A(n10690), .B(n10805), .Z(n10694) );
  XNOR U6545 ( .A(n11058), .B(n11174), .Z(n11062) );
  XNOR U6546 ( .A(n11427), .B(n11543), .Z(n11431) );
  XNOR U6547 ( .A(n12169), .B(n11798), .Z(n11800) );
  XNOR U6548 ( .A(n12537), .B(n12166), .Z(n12168) );
  XNOR U6549 ( .A(n12905), .B(n12534), .Z(n12536) );
  XNOR U6550 ( .A(n13273), .B(n12902), .Z(n12904) );
  XNOR U6551 ( .A(n13641), .B(n13270), .Z(n13272) );
  XNOR U6552 ( .A(n14009), .B(n13638), .Z(n13640) );
  XNOR U6553 ( .A(n14377), .B(n14006), .Z(n14008) );
  XNOR U6554 ( .A(n14745), .B(n14374), .Z(n14376) );
  XNOR U6555 ( .A(n15113), .B(n14742), .Z(n14744) );
  XNOR U6556 ( .A(n15481), .B(n15110), .Z(n15112) );
  XNOR U6557 ( .A(n15849), .B(n15478), .Z(n15480) );
  XNOR U6558 ( .A(n16217), .B(n15846), .Z(n15848) );
  XNOR U6559 ( .A(n16585), .B(n16214), .Z(n16216) );
  XNOR U6560 ( .A(n16953), .B(n16582), .Z(n16584) );
  XNOR U6561 ( .A(n17321), .B(n16950), .Z(n16952) );
  XNOR U6562 ( .A(n17689), .B(n17318), .Z(n17320) );
  XNOR U6563 ( .A(n3450), .B(n3582), .Z(n3454) );
  XNOR U6564 ( .A(n3793), .B(n3963), .Z(n3788) );
  XNOR U6565 ( .A(n3025), .B(n3223), .Z(n3029) );
  XNOR U6566 ( .A(n2259), .B(n2482), .Z(n2263) );
  XNOR U6567 ( .A(n2603), .B(n2864), .Z(n2598) );
  XNOR U6568 ( .A(n1834), .B(n2122), .Z(n1838) );
  XNOR U6569 ( .A(n1070), .B(n1382), .Z(n1074) );
  XNOR U6570 ( .A(n4209), .B(n4323), .Z(n4213) );
  XNOR U6571 ( .A(n6815), .B(n6925), .Z(n6819) );
  XNOR U6572 ( .A(n34431), .B(n34533), .Z(n34435) );
  XNOR U6573 ( .A(n34192), .B(n34294), .Z(n34196) );
  XNOR U6574 ( .A(n33929), .B(n34034), .Z(n33933) );
  XNOR U6575 ( .A(n33645), .B(n33747), .Z(n33649) );
  XNOR U6576 ( .A(n33334), .B(n33436), .Z(n33338) );
  XNOR U6577 ( .A(n32999), .B(n33104), .Z(n33003) );
  XNOR U6578 ( .A(n32643), .B(n32745), .Z(n32647) );
  XNOR U6579 ( .A(n32260), .B(n32362), .Z(n32264) );
  XNOR U6580 ( .A(n31677), .B(n31958), .Z(n31681) );
  XNOR U6581 ( .A(n31233), .B(n31343), .Z(n31237) );
  XNOR U6582 ( .A(n30765), .B(n30875), .Z(n30769) );
  XNOR U6583 ( .A(n30273), .B(n30383), .Z(n30277) );
  XNOR U6584 ( .A(n29757), .B(n29867), .Z(n29761) );
  XNOR U6585 ( .A(n29217), .B(n29327), .Z(n29221) );
  XNOR U6586 ( .A(n28653), .B(n28763), .Z(n28657) );
  XNOR U6587 ( .A(n28065), .B(n28175), .Z(n28069) );
  XNOR U6588 ( .A(n27453), .B(n27563), .Z(n27457) );
  XNOR U6589 ( .A(n26817), .B(n26927), .Z(n26821) );
  XNOR U6590 ( .A(n26157), .B(n26267), .Z(n26161) );
  XNOR U6591 ( .A(n25473), .B(n25583), .Z(n25477) );
  XNOR U6592 ( .A(n24765), .B(n24875), .Z(n24769) );
  XNOR U6593 ( .A(n24030), .B(n24140), .Z(n24034) );
  XNOR U6594 ( .A(n1442), .B(n1756), .Z(n1437) );
  XNOR U6595 ( .A(n674), .B(n1016), .Z(n678) );
  XNOR U6596 ( .A(n2632), .B(n2857), .Z(n2627) );
  XNOR U6597 ( .A(n1863), .B(n2115), .Z(n1867) );
  XNOR U6598 ( .A(n1099), .B(n1375), .Z(n1103) );
  XNOR U6599 ( .A(n3822), .B(n3956), .Z(n3817) );
  XNOR U6600 ( .A(n3054), .B(n3216), .Z(n3058) );
  XNOR U6601 ( .A(n2288), .B(n2475), .Z(n2292) );
  XNOR U6602 ( .A(n4958), .B(n5067), .Z(n4962) );
  XNOR U6603 ( .A(n5708), .B(n5812), .Z(n5703) );
  XNOR U6604 ( .A(n6448), .B(n6556), .Z(n6452) );
  XNOR U6605 ( .A(n18803), .B(n18432), .Z(n18434) );
  XNOR U6606 ( .A(n19171), .B(n18800), .Z(n18802) );
  XNOR U6607 ( .A(n19539), .B(n19168), .Z(n19170) );
  XNOR U6608 ( .A(n19907), .B(n19536), .Z(n19538) );
  XNOR U6609 ( .A(n20275), .B(n19904), .Z(n19906) );
  XNOR U6610 ( .A(n20643), .B(n20272), .Z(n20274) );
  XNOR U6611 ( .A(n21011), .B(n20640), .Z(n20642) );
  XNOR U6612 ( .A(n21379), .B(n21008), .Z(n21010) );
  XNOR U6613 ( .A(n21747), .B(n21376), .Z(n21378) );
  XNOR U6614 ( .A(n22115), .B(n21744), .Z(n21746) );
  XNOR U6615 ( .A(n22483), .B(n22112), .Z(n22114) );
  XNOR U6616 ( .A(n22851), .B(n22480), .Z(n22482) );
  XNOR U6617 ( .A(n23219), .B(n22848), .Z(n22850) );
  XNOR U6618 ( .A(n23213), .B(n23317), .Z(n23217) );
  XNOR U6619 ( .A(n3842), .B(n3950), .Z(n3850) );
  XNOR U6620 ( .A(n7943), .B(n8042), .Z(n7944) );
  XNOR U6621 ( .A(n8685), .B(n8787), .Z(n8693) );
  XNOR U6622 ( .A(n9425), .B(n9530), .Z(n9429) );
  XNOR U6623 ( .A(n10172), .B(n10393), .Z(n10181) );
  XNOR U6624 ( .A(n10705), .B(n10802), .Z(n10709) );
  XNOR U6625 ( .A(n11073), .B(n11171), .Z(n11077) );
  XNOR U6626 ( .A(n11442), .B(n11540), .Z(n11446) );
  XNOR U6627 ( .A(n12184), .B(n11813), .Z(n11815) );
  XNOR U6628 ( .A(n12552), .B(n12181), .Z(n12183) );
  XNOR U6629 ( .A(n12920), .B(n12549), .Z(n12551) );
  XNOR U6630 ( .A(n13288), .B(n12917), .Z(n12919) );
  XNOR U6631 ( .A(n13656), .B(n13285), .Z(n13287) );
  XNOR U6632 ( .A(n14024), .B(n13653), .Z(n13655) );
  XNOR U6633 ( .A(n14392), .B(n14021), .Z(n14023) );
  XNOR U6634 ( .A(n14760), .B(n14389), .Z(n14391) );
  XNOR U6635 ( .A(n15128), .B(n14757), .Z(n14759) );
  XNOR U6636 ( .A(n15496), .B(n15125), .Z(n15127) );
  XNOR U6637 ( .A(n15864), .B(n15493), .Z(n15495) );
  XNOR U6638 ( .A(n16232), .B(n15861), .Z(n15863) );
  XNOR U6639 ( .A(n16600), .B(n16229), .Z(n16231) );
  XNOR U6640 ( .A(n16968), .B(n16597), .Z(n16599) );
  XNOR U6641 ( .A(n17336), .B(n16965), .Z(n16967) );
  XNOR U6642 ( .A(n17704), .B(n17333), .Z(n17335) );
  XNOR U6643 ( .A(n18072), .B(n17701), .Z(n17703) );
  XNOR U6644 ( .A(n18440), .B(n18069), .Z(n18071) );
  XNOR U6645 ( .A(n18808), .B(n18437), .Z(n18439) );
  XNOR U6646 ( .A(n3083), .B(n3209), .Z(n3087) );
  XNOR U6647 ( .A(n2317), .B(n2468), .Z(n2321) );
  XNOR U6648 ( .A(n2661), .B(n2850), .Z(n2656) );
  XNOR U6649 ( .A(n1892), .B(n2108), .Z(n1896) );
  XNOR U6650 ( .A(n1128), .B(n1368), .Z(n1132) );
  XNOR U6651 ( .A(n1471), .B(n1749), .Z(n1466) );
  XNOR U6652 ( .A(n703), .B(n1009), .Z(n707) );
  XNOR U6653 ( .A(n7573), .B(n7669), .Z(n7577) );
  XNOR U6654 ( .A(n34849), .B(n34933), .Z(n34853) );
  XNOR U6655 ( .A(n34658), .B(n34745), .Z(n34662) );
  XNOR U6656 ( .A(n34446), .B(n34530), .Z(n34450) );
  XNOR U6657 ( .A(n34207), .B(n34291), .Z(n34211) );
  XNOR U6658 ( .A(n33944), .B(n34031), .Z(n33948) );
  XNOR U6659 ( .A(n33660), .B(n33744), .Z(n33664) );
  XNOR U6660 ( .A(n33349), .B(n33433), .Z(n33353) );
  XNOR U6661 ( .A(n33014), .B(n33101), .Z(n33018) );
  XNOR U6662 ( .A(n32658), .B(n32742), .Z(n32662) );
  XNOR U6663 ( .A(n32275), .B(n32359), .Z(n32279) );
  XNOR U6664 ( .A(n31692), .B(n31955), .Z(n31696) );
  XNOR U6665 ( .A(n31248), .B(n31340), .Z(n31252) );
  XNOR U6666 ( .A(n30780), .B(n30872), .Z(n30784) );
  XNOR U6667 ( .A(n30288), .B(n30380), .Z(n30292) );
  XNOR U6668 ( .A(n29772), .B(n29864), .Z(n29776) );
  XNOR U6669 ( .A(n29232), .B(n29324), .Z(n29236) );
  XNOR U6670 ( .A(n28668), .B(n28760), .Z(n28672) );
  XNOR U6671 ( .A(n28080), .B(n28172), .Z(n28084) );
  XNOR U6672 ( .A(n27468), .B(n27560), .Z(n27472) );
  XNOR U6673 ( .A(n26832), .B(n26924), .Z(n26836) );
  XNOR U6674 ( .A(n26172), .B(n26264), .Z(n26176) );
  XNOR U6675 ( .A(n25488), .B(n25580), .Z(n25492) );
  XNOR U6676 ( .A(n24780), .B(n24872), .Z(n24784) );
  XNOR U6677 ( .A(n24045), .B(n24137), .Z(n24049) );
  XNOR U6678 ( .A(n340), .B(n631), .Z(n353) );
  XNOR U6679 ( .A(n1500), .B(n1742), .Z(n1495) );
  XNOR U6680 ( .A(n732), .B(n1002), .Z(n736) );
  XNOR U6681 ( .A(n2690), .B(n2843), .Z(n2685) );
  XNOR U6682 ( .A(n1921), .B(n2101), .Z(n1925) );
  XNOR U6683 ( .A(n1157), .B(n1361), .Z(n1161) );
  XNOR U6684 ( .A(n2346), .B(n2461), .Z(n2350) );
  XNOR U6685 ( .A(n3484), .B(n3574), .Z(n3488) );
  XNOR U6686 ( .A(n4231), .B(n4318), .Z(n4232) );
  XNOR U6687 ( .A(n4973), .B(n5064), .Z(n4981) );
  XNOR U6688 ( .A(n5718), .B(n5808), .Z(n5722) );
  XNOR U6689 ( .A(n6465), .B(n6552), .Z(n6466) );
  XNOR U6690 ( .A(n7203), .B(n7296), .Z(n7211) );
  XNOR U6691 ( .A(n19922), .B(n19551), .Z(n19553) );
  XNOR U6692 ( .A(n20290), .B(n19919), .Z(n19921) );
  XNOR U6693 ( .A(n20658), .B(n20287), .Z(n20289) );
  XNOR U6694 ( .A(n21026), .B(n20655), .Z(n20657) );
  XNOR U6695 ( .A(n21394), .B(n21023), .Z(n21025) );
  XNOR U6696 ( .A(n21762), .B(n21391), .Z(n21393) );
  XNOR U6697 ( .A(n22130), .B(n21759), .Z(n21761) );
  XNOR U6698 ( .A(n22498), .B(n22127), .Z(n22129) );
  XNOR U6699 ( .A(n22866), .B(n22495), .Z(n22497) );
  XNOR U6700 ( .A(n23234), .B(n22863), .Z(n22865) );
  XNOR U6701 ( .A(n23228), .B(n23314), .Z(n23232) );
  XNOR U6702 ( .A(n8699), .B(n8783), .Z(n8703) );
  XNOR U6703 ( .A(n9444), .B(n9527), .Z(n9439) );
  XNOR U6704 ( .A(n10192), .B(n10387), .Z(n10196) );
  XNOR U6705 ( .A(n10720), .B(n10799), .Z(n10724) );
  XNOR U6706 ( .A(n11088), .B(n11168), .Z(n11092) );
  XNOR U6707 ( .A(n11457), .B(n11537), .Z(n11461) );
  XNOR U6708 ( .A(n12199), .B(n11828), .Z(n11830) );
  XNOR U6709 ( .A(n12567), .B(n12196), .Z(n12198) );
  XNOR U6710 ( .A(n12935), .B(n12564), .Z(n12566) );
  XNOR U6711 ( .A(n13303), .B(n12932), .Z(n12934) );
  XNOR U6712 ( .A(n13671), .B(n13300), .Z(n13302) );
  XNOR U6713 ( .A(n14039), .B(n13668), .Z(n13670) );
  XNOR U6714 ( .A(n14407), .B(n14036), .Z(n14038) );
  XNOR U6715 ( .A(n14775), .B(n14404), .Z(n14406) );
  XNOR U6716 ( .A(n15143), .B(n14772), .Z(n14774) );
  XNOR U6717 ( .A(n15511), .B(n15140), .Z(n15142) );
  XNOR U6718 ( .A(n15879), .B(n15508), .Z(n15510) );
  XNOR U6719 ( .A(n16247), .B(n15876), .Z(n15878) );
  XNOR U6720 ( .A(n16615), .B(n16244), .Z(n16246) );
  XNOR U6721 ( .A(n16983), .B(n16612), .Z(n16614) );
  XNOR U6722 ( .A(n17351), .B(n16980), .Z(n16982) );
  XNOR U6723 ( .A(n17719), .B(n17348), .Z(n17350) );
  XNOR U6724 ( .A(n18087), .B(n17716), .Z(n17718) );
  XNOR U6725 ( .A(n18455), .B(n18084), .Z(n18086) );
  XNOR U6726 ( .A(n18823), .B(n18452), .Z(n18454) );
  XNOR U6727 ( .A(n19191), .B(n18820), .Z(n18822) );
  XNOR U6728 ( .A(n19559), .B(n19188), .Z(n19190) );
  XNOR U6729 ( .A(n19927), .B(n19556), .Z(n19558) );
  XNOR U6730 ( .A(n2719), .B(n2836), .Z(n2714) );
  XNOR U6731 ( .A(n1950), .B(n2094), .Z(n1954) );
  XNOR U6732 ( .A(n1186), .B(n1354), .Z(n1190) );
  XNOR U6733 ( .A(n1529), .B(n1735), .Z(n1524) );
  XNOR U6734 ( .A(n761), .B(n995), .Z(n765) );
  XNOR U6735 ( .A(n324), .B(n612), .Z(n363) );
  XNOR U6736 ( .A(n2739), .B(n2830), .Z(n2747) );
  XNOR U6737 ( .A(n8332), .B(n8410), .Z(n8336) );
  XNOR U6738 ( .A(n35031), .B(n35097), .Z(n35035) );
  XNOR U6739 ( .A(n34864), .B(n34930), .Z(n34868) );
  XNOR U6740 ( .A(n34673), .B(n34742), .Z(n34677) );
  XNOR U6741 ( .A(n34461), .B(n34527), .Z(n34465) );
  XNOR U6742 ( .A(n34222), .B(n34288), .Z(n34226) );
  XNOR U6743 ( .A(n33959), .B(n34028), .Z(n33963) );
  XNOR U6744 ( .A(n33675), .B(n33741), .Z(n33679) );
  XNOR U6745 ( .A(n33364), .B(n33430), .Z(n33368) );
  XNOR U6746 ( .A(n33029), .B(n33098), .Z(n33033) );
  XNOR U6747 ( .A(n32673), .B(n32739), .Z(n32677) );
  XNOR U6748 ( .A(n32290), .B(n32356), .Z(n32294) );
  XNOR U6749 ( .A(n31707), .B(n31952), .Z(n31711) );
  XNOR U6750 ( .A(n31263), .B(n31337), .Z(n31267) );
  XNOR U6751 ( .A(n30795), .B(n30869), .Z(n30799) );
  XNOR U6752 ( .A(n30303), .B(n30377), .Z(n30307) );
  XNOR U6753 ( .A(n29787), .B(n29861), .Z(n29791) );
  XNOR U6754 ( .A(n29247), .B(n29321), .Z(n29251) );
  XNOR U6755 ( .A(n28683), .B(n28757), .Z(n28687) );
  XNOR U6756 ( .A(n28095), .B(n28169), .Z(n28099) );
  XNOR U6757 ( .A(n27483), .B(n27557), .Z(n27487) );
  XNOR U6758 ( .A(n26847), .B(n26921), .Z(n26851) );
  XNOR U6759 ( .A(n26187), .B(n26261), .Z(n26191) );
  XNOR U6760 ( .A(n25503), .B(n25577), .Z(n25507) );
  XNOR U6761 ( .A(n24795), .B(n24869), .Z(n24799) );
  XNOR U6762 ( .A(n24060), .B(n24134), .Z(n24064) );
  XNOR U6763 ( .A(n308), .B(n593), .Z(n373) );
  XNOR U6764 ( .A(n1558), .B(n1728), .Z(n1553) );
  XNOR U6765 ( .A(n790), .B(n988), .Z(n794) );
  XNOR U6766 ( .A(n1979), .B(n2087), .Z(n1983) );
  XNOR U6767 ( .A(n1215), .B(n1347), .Z(n1219) );
  XNOR U6768 ( .A(n2753), .B(n2826), .Z(n2757) );
  XNOR U6769 ( .A(n3503), .B(n3571), .Z(n3498) );
  XNOR U6770 ( .A(n4243), .B(n4315), .Z(n4247) );
  XNOR U6771 ( .A(n4987), .B(n5060), .Z(n4991) );
  XNOR U6772 ( .A(n5737), .B(n5805), .Z(n5732) );
  XNOR U6773 ( .A(n6477), .B(n6549), .Z(n6481) );
  XNOR U6774 ( .A(n7217), .B(n7292), .Z(n7221) );
  XNOR U6775 ( .A(n7969), .B(n8037), .Z(n7964) );
  XNOR U6776 ( .A(n21041), .B(n20670), .Z(n20672) );
  XNOR U6777 ( .A(n21409), .B(n21038), .Z(n21040) );
  XNOR U6778 ( .A(n21777), .B(n21406), .Z(n21408) );
  XNOR U6779 ( .A(n22145), .B(n21774), .Z(n21776) );
  XNOR U6780 ( .A(n22513), .B(n22142), .Z(n22144) );
  XNOR U6781 ( .A(n22881), .B(n22510), .Z(n22512) );
  XNOR U6782 ( .A(n23249), .B(n22878), .Z(n22880) );
  XNOR U6783 ( .A(n23243), .B(n23311), .Z(n23247) );
  XNOR U6784 ( .A(n9454), .B(n9523), .Z(n9458) );
  XNOR U6785 ( .A(n10201), .B(n10382), .Z(n10210) );
  XNOR U6786 ( .A(n10735), .B(n10796), .Z(n10739) );
  XNOR U6787 ( .A(n11103), .B(n11165), .Z(n11107) );
  XNOR U6788 ( .A(n11472), .B(n11534), .Z(n11476) );
  XNOR U6789 ( .A(n12214), .B(n11843), .Z(n11845) );
  XNOR U6790 ( .A(n12582), .B(n12211), .Z(n12213) );
  XNOR U6791 ( .A(n12950), .B(n12579), .Z(n12581) );
  XNOR U6792 ( .A(n13318), .B(n12947), .Z(n12949) );
  XNOR U6793 ( .A(n13686), .B(n13315), .Z(n13317) );
  XNOR U6794 ( .A(n14054), .B(n13683), .Z(n13685) );
  XNOR U6795 ( .A(n14422), .B(n14051), .Z(n14053) );
  XNOR U6796 ( .A(n14790), .B(n14419), .Z(n14421) );
  XNOR U6797 ( .A(n15158), .B(n14787), .Z(n14789) );
  XNOR U6798 ( .A(n15526), .B(n15155), .Z(n15157) );
  XNOR U6799 ( .A(n15894), .B(n15523), .Z(n15525) );
  XNOR U6800 ( .A(n16262), .B(n15891), .Z(n15893) );
  XNOR U6801 ( .A(n16630), .B(n16259), .Z(n16261) );
  XNOR U6802 ( .A(n16998), .B(n16627), .Z(n16629) );
  XNOR U6803 ( .A(n17366), .B(n16995), .Z(n16997) );
  XNOR U6804 ( .A(n17734), .B(n17363), .Z(n17365) );
  XNOR U6805 ( .A(n18102), .B(n17731), .Z(n17733) );
  XNOR U6806 ( .A(n18470), .B(n18099), .Z(n18101) );
  XNOR U6807 ( .A(n18838), .B(n18467), .Z(n18469) );
  XNOR U6808 ( .A(n19206), .B(n18835), .Z(n18837) );
  XNOR U6809 ( .A(n19574), .B(n19203), .Z(n19205) );
  XNOR U6810 ( .A(n19942), .B(n19571), .Z(n19573) );
  XNOR U6811 ( .A(n20310), .B(n19939), .Z(n19941) );
  XNOR U6812 ( .A(n20678), .B(n20307), .Z(n20309) );
  XNOR U6813 ( .A(n21046), .B(n20675), .Z(n20677) );
  XNOR U6814 ( .A(n1587), .B(n1721), .Z(n1582) );
  XNOR U6815 ( .A(n819), .B(n981), .Z(n823) );
  XNOR U6816 ( .A(n292), .B(n574), .Z(n383) );
  XNOR U6817 ( .A(n9091), .B(n9147), .Z(n9099) );
  XNOR U6818 ( .A(n35305), .B(n35353), .Z(n35309) );
  XNOR U6819 ( .A(n35186), .B(n35237), .Z(n35190) );
  XNOR U6820 ( .A(n35046), .B(n35094), .Z(n35050) );
  XNOR U6821 ( .A(n34879), .B(n34927), .Z(n34883) );
  XNOR U6822 ( .A(n34688), .B(n34739), .Z(n34692) );
  XNOR U6823 ( .A(n34476), .B(n34524), .Z(n34480) );
  XNOR U6824 ( .A(n34237), .B(n34285), .Z(n34241) );
  XNOR U6825 ( .A(n33974), .B(n34025), .Z(n33978) );
  XNOR U6826 ( .A(n33690), .B(n33738), .Z(n33694) );
  XNOR U6827 ( .A(n33379), .B(n33427), .Z(n33383) );
  XNOR U6828 ( .A(n33044), .B(n33095), .Z(n33048) );
  XNOR U6829 ( .A(n32688), .B(n32736), .Z(n32692) );
  XNOR U6830 ( .A(n32305), .B(n32353), .Z(n32309) );
  XNOR U6831 ( .A(n31722), .B(n31949), .Z(n31726) );
  XNOR U6832 ( .A(n31278), .B(n31334), .Z(n31282) );
  XNOR U6833 ( .A(n30810), .B(n30866), .Z(n30814) );
  XNOR U6834 ( .A(n30318), .B(n30374), .Z(n30322) );
  XNOR U6835 ( .A(n29802), .B(n29858), .Z(n29806) );
  XNOR U6836 ( .A(n29262), .B(n29318), .Z(n29266) );
  XNOR U6837 ( .A(n28698), .B(n28754), .Z(n28702) );
  XNOR U6838 ( .A(n28110), .B(n28166), .Z(n28114) );
  XNOR U6839 ( .A(n27498), .B(n27554), .Z(n27502) );
  XNOR U6840 ( .A(n26862), .B(n26918), .Z(n26866) );
  XNOR U6841 ( .A(n26202), .B(n26258), .Z(n26206) );
  XNOR U6842 ( .A(n25518), .B(n25574), .Z(n25522) );
  XNOR U6843 ( .A(n24810), .B(n24866), .Z(n24814) );
  XNOR U6844 ( .A(n24075), .B(n24131), .Z(n24079) );
  XNOR U6845 ( .A(n1631), .B(n1709), .Z(n1635) );
  XNOR U6846 ( .A(n867), .B(n969), .Z(n871) );
  XNOR U6847 ( .A(n276), .B(n555), .Z(n393) );
  XNOR U6848 ( .A(n1616), .B(n1714), .Z(n1611) );
  XNOR U6849 ( .A(n848), .B(n974), .Z(n852) );
  XNOR U6850 ( .A(n2023), .B(n2077), .Z(n2027) );
  XNOR U6851 ( .A(n2768), .B(n2823), .Z(n2772) );
  XNOR U6852 ( .A(n3513), .B(n3567), .Z(n3517) );
  XNOR U6853 ( .A(n4260), .B(n4311), .Z(n4261) );
  XNOR U6854 ( .A(n5002), .B(n5057), .Z(n5010) );
  XNOR U6855 ( .A(n5747), .B(n5801), .Z(n5751) );
  XNOR U6856 ( .A(n6494), .B(n6545), .Z(n6495) );
  XNOR U6857 ( .A(n7232), .B(n7289), .Z(n7240) );
  XNOR U6858 ( .A(n7979), .B(n8033), .Z(n7983) );
  XNOR U6859 ( .A(n8726), .B(n8777), .Z(n8727) );
  XNOR U6860 ( .A(n22160), .B(n21789), .Z(n21791) );
  XNOR U6861 ( .A(n22528), .B(n22157), .Z(n22159) );
  XNOR U6862 ( .A(n22896), .B(n22525), .Z(n22527) );
  XNOR U6863 ( .A(n23264), .B(n22893), .Z(n22895) );
  XNOR U6864 ( .A(n23258), .B(n23308), .Z(n23262) );
  XNOR U6865 ( .A(n897), .B(n963), .Z(n901) );
  XNOR U6866 ( .A(n10221), .B(n10376), .Z(n10225) );
  XNOR U6867 ( .A(n11118), .B(n11162), .Z(n11122) );
  XNOR U6868 ( .A(n11487), .B(n11531), .Z(n11491) );
  XNOR U6869 ( .A(n12229), .B(n11858), .Z(n11860) );
  XNOR U6870 ( .A(n12597), .B(n12226), .Z(n12228) );
  XNOR U6871 ( .A(n12965), .B(n12594), .Z(n12596) );
  XNOR U6872 ( .A(n13333), .B(n12962), .Z(n12964) );
  XNOR U6873 ( .A(n13701), .B(n13330), .Z(n13332) );
  XNOR U6874 ( .A(n14069), .B(n13698), .Z(n13700) );
  XNOR U6875 ( .A(n14437), .B(n14066), .Z(n14068) );
  XNOR U6876 ( .A(n14805), .B(n14434), .Z(n14436) );
  XNOR U6877 ( .A(n15173), .B(n14802), .Z(n14804) );
  XNOR U6878 ( .A(n15541), .B(n15170), .Z(n15172) );
  XNOR U6879 ( .A(n15909), .B(n15538), .Z(n15540) );
  XNOR U6880 ( .A(n16277), .B(n15906), .Z(n15908) );
  XNOR U6881 ( .A(n16645), .B(n16274), .Z(n16276) );
  XNOR U6882 ( .A(n17013), .B(n16642), .Z(n16644) );
  XNOR U6883 ( .A(n17381), .B(n17010), .Z(n17012) );
  XNOR U6884 ( .A(n17749), .B(n17378), .Z(n17380) );
  XNOR U6885 ( .A(n18117), .B(n17746), .Z(n17748) );
  XNOR U6886 ( .A(n18485), .B(n18114), .Z(n18116) );
  XNOR U6887 ( .A(n18853), .B(n18482), .Z(n18484) );
  XNOR U6888 ( .A(n19221), .B(n18850), .Z(n18852) );
  XNOR U6889 ( .A(n19589), .B(n19218), .Z(n19220) );
  XNOR U6890 ( .A(n19957), .B(n19586), .Z(n19588) );
  XNOR U6891 ( .A(n20325), .B(n19954), .Z(n19956) );
  XNOR U6892 ( .A(n20693), .B(n20322), .Z(n20324) );
  XNOR U6893 ( .A(n21061), .B(n20690), .Z(n20692) );
  XNOR U6894 ( .A(n21429), .B(n21058), .Z(n21060) );
  XNOR U6895 ( .A(n21797), .B(n21426), .Z(n21428) );
  XNOR U6896 ( .A(n22165), .B(n21794), .Z(n21796) );
  XNOR U6897 ( .A(n260), .B(n536), .Z(n403) );
  XNOR U6898 ( .A(n9853), .B(n9892), .Z(n9847) );
  XNOR U6899 ( .A(n35415), .B(n35445), .Z(n35419) );
  XNOR U6900 ( .A(n35320), .B(n35350), .Z(n35324) );
  XNOR U6901 ( .A(n35201), .B(n35234), .Z(n35205) );
  XNOR U6902 ( .A(n35061), .B(n35091), .Z(n35065) );
  XNOR U6903 ( .A(n34894), .B(n34924), .Z(n34898) );
  XNOR U6904 ( .A(n34703), .B(n34736), .Z(n34707) );
  XNOR U6905 ( .A(n34491), .B(n34521), .Z(n34495) );
  XNOR U6906 ( .A(n34252), .B(n34282), .Z(n34256) );
  XNOR U6907 ( .A(n33989), .B(n34022), .Z(n33993) );
  XNOR U6908 ( .A(n33705), .B(n33735), .Z(n33709) );
  XNOR U6909 ( .A(n33394), .B(n33424), .Z(n33398) );
  XNOR U6910 ( .A(n33059), .B(n33092), .Z(n33063) );
  XNOR U6911 ( .A(n32703), .B(n32733), .Z(n32707) );
  XNOR U6912 ( .A(n32320), .B(n32350), .Z(n32324) );
  XNOR U6913 ( .A(n31737), .B(n31946), .Z(n31741) );
  XNOR U6914 ( .A(n31293), .B(n31331), .Z(n31297) );
  XNOR U6915 ( .A(n30825), .B(n30863), .Z(n30829) );
  XNOR U6916 ( .A(n30333), .B(n30371), .Z(n30337) );
  XNOR U6917 ( .A(n29817), .B(n29855), .Z(n29821) );
  XNOR U6918 ( .A(n29277), .B(n29315), .Z(n29281) );
  XNOR U6919 ( .A(n28713), .B(n28751), .Z(n28717) );
  XNOR U6920 ( .A(n28125), .B(n28163), .Z(n28129) );
  XNOR U6921 ( .A(n27513), .B(n27551), .Z(n27517) );
  XNOR U6922 ( .A(n26877), .B(n26915), .Z(n26881) );
  XNOR U6923 ( .A(n26217), .B(n26255), .Z(n26221) );
  XNOR U6924 ( .A(n25533), .B(n25571), .Z(n25537) );
  XNOR U6925 ( .A(n24825), .B(n24863), .Z(n24829) );
  XNOR U6926 ( .A(n24090), .B(n24128), .Z(n24094) );
  XNOR U6927 ( .A(n882), .B(n966), .Z(n886) );
  XNOR U6928 ( .A(n244), .B(n517), .Z(n413) );
  XNOR U6929 ( .A(n2038), .B(n2074), .Z(n2042) );
  XNOR U6930 ( .A(n2783), .B(n2820), .Z(n2787) );
  XNOR U6931 ( .A(n3528), .B(n3564), .Z(n3532) );
  XNOR U6932 ( .A(n4272), .B(n4308), .Z(n4276) );
  XNOR U6933 ( .A(n5016), .B(n5053), .Z(n5020) );
  XNOR U6934 ( .A(n5766), .B(n5798), .Z(n5761) );
  XNOR U6935 ( .A(n6878), .B(n6910), .Z(n6882) );
  XNOR U6936 ( .A(n7624), .B(n7657), .Z(n7625) );
  XNOR U6937 ( .A(n8366), .B(n8402), .Z(n8374) );
  XNOR U6938 ( .A(n9478), .B(n9517), .Z(n9482) );
  XNOR U6939 ( .A(n10760), .B(n10791), .Z(n10764) );
  XNOR U6940 ( .A(n23279), .B(n22908), .Z(n22910) );
  XNOR U6941 ( .A(n23273), .B(n23305), .Z(n23277) );
  XNOR U6942 ( .A(n912), .B(n960), .Z(n916) );
  XNOR U6943 ( .A(n6511), .B(n6541), .Z(n6519) );
  XNOR U6944 ( .A(n9115), .B(n9141), .Z(n9119) );
  XNOR U6945 ( .A(n11502), .B(n11528), .Z(n11506) );
  XNOR U6946 ( .A(n12244), .B(n11873), .Z(n11875) );
  XNOR U6947 ( .A(n12612), .B(n12241), .Z(n12243) );
  XNOR U6948 ( .A(n12980), .B(n12609), .Z(n12611) );
  XNOR U6949 ( .A(n13348), .B(n12977), .Z(n12979) );
  XNOR U6950 ( .A(n13716), .B(n13345), .Z(n13347) );
  XNOR U6951 ( .A(n14084), .B(n13713), .Z(n13715) );
  XNOR U6952 ( .A(n14452), .B(n14081), .Z(n14083) );
  XNOR U6953 ( .A(n14820), .B(n14449), .Z(n14451) );
  XNOR U6954 ( .A(n15188), .B(n14817), .Z(n14819) );
  XNOR U6955 ( .A(n15556), .B(n15185), .Z(n15187) );
  XNOR U6956 ( .A(n15924), .B(n15553), .Z(n15555) );
  XNOR U6957 ( .A(n16292), .B(n15921), .Z(n15923) );
  XNOR U6958 ( .A(n16660), .B(n16289), .Z(n16291) );
  XNOR U6959 ( .A(n17028), .B(n16657), .Z(n16659) );
  XNOR U6960 ( .A(n17396), .B(n17025), .Z(n17027) );
  XNOR U6961 ( .A(n17764), .B(n17393), .Z(n17395) );
  XNOR U6962 ( .A(n18132), .B(n17761), .Z(n17763) );
  XNOR U6963 ( .A(n18500), .B(n18129), .Z(n18131) );
  XNOR U6964 ( .A(n18868), .B(n18497), .Z(n18499) );
  XNOR U6965 ( .A(n19236), .B(n18865), .Z(n18867) );
  XNOR U6966 ( .A(n19604), .B(n19233), .Z(n19235) );
  XNOR U6967 ( .A(n19972), .B(n19601), .Z(n19603) );
  XNOR U6968 ( .A(n20340), .B(n19969), .Z(n19971) );
  XNOR U6969 ( .A(n20708), .B(n20337), .Z(n20339) );
  XNOR U6970 ( .A(n21076), .B(n20705), .Z(n20707) );
  XNOR U6971 ( .A(n21444), .B(n21073), .Z(n21075) );
  XNOR U6972 ( .A(n21812), .B(n21441), .Z(n21443) );
  XNOR U6973 ( .A(n22180), .B(n21809), .Z(n21811) );
  XNOR U6974 ( .A(n22548), .B(n22177), .Z(n22179) );
  XNOR U6975 ( .A(n22916), .B(n22545), .Z(n22547) );
  XNOR U6976 ( .A(n23284), .B(n22913), .Z(n22915) );
  XNOR U6977 ( .A(n11138), .B(n11158), .Z(n11142) );
  XNOR U6978 ( .A(n35545), .B(n35557), .Z(n35550) );
  XNOR U6979 ( .A(n35498), .B(n35513), .Z(n35507) );
  XNOR U6980 ( .A(n35430), .B(n35442), .Z(n35434) );
  XNOR U6981 ( .A(n35335), .B(n35347), .Z(n35340) );
  XNOR U6982 ( .A(n35216), .B(n35231), .Z(n35225) );
  XNOR U6983 ( .A(n35076), .B(n35088), .Z(n35080) );
  XNOR U6984 ( .A(n34909), .B(n34921), .Z(n34914) );
  XNOR U6985 ( .A(n34718), .B(n34733), .Z(n34727) );
  XNOR U6986 ( .A(n34506), .B(n34518), .Z(n34510) );
  XNOR U6987 ( .A(n34267), .B(n34279), .Z(n34272) );
  XNOR U6988 ( .A(n34004), .B(n34019), .Z(n34013) );
  XNOR U6989 ( .A(n33720), .B(n33732), .Z(n33724) );
  XNOR U6990 ( .A(n33409), .B(n33421), .Z(n33414) );
  XNOR U6991 ( .A(n33074), .B(n33089), .Z(n33083) );
  XNOR U6992 ( .A(n32718), .B(n32730), .Z(n32722) );
  XNOR U6993 ( .A(n32335), .B(n32347), .Z(n32340) );
  XNOR U6994 ( .A(n31752), .B(n31943), .Z(n31761) );
  XNOR U6995 ( .A(n31308), .B(n31328), .Z(n31317) );
  XNOR U6996 ( .A(n30840), .B(n30860), .Z(n30849) );
  XNOR U6997 ( .A(n30348), .B(n30368), .Z(n30357) );
  XNOR U6998 ( .A(n29832), .B(n29852), .Z(n29841) );
  XNOR U6999 ( .A(n29292), .B(n29312), .Z(n29301) );
  XNOR U7000 ( .A(n28728), .B(n28748), .Z(n28737) );
  XNOR U7001 ( .A(n28140), .B(n28160), .Z(n28149) );
  XNOR U7002 ( .A(n27528), .B(n27548), .Z(n27537) );
  XNOR U7003 ( .A(n26892), .B(n26912), .Z(n26901) );
  XNOR U7004 ( .A(n26232), .B(n26252), .Z(n26241) );
  XNOR U7005 ( .A(n25548), .B(n25568), .Z(n25557) );
  XNOR U7006 ( .A(n24840), .B(n24860), .Z(n24849) );
  XNOR U7007 ( .A(n24105), .B(n24125), .Z(n24114) );
  XNOR U7008 ( .A(n1309), .B(n1327), .Z(n1318) );
  XNOR U7009 ( .A(n2053), .B(n2071), .Z(n2062) );
  XNOR U7010 ( .A(n3171), .B(n3189), .Z(n3180) );
  XNOR U7011 ( .A(n3915), .B(n3933), .Z(n3924) );
  XNOR U7012 ( .A(n4659), .B(n4677), .Z(n4667) );
  XNOR U7013 ( .A(n5404), .B(n5422), .Z(n5413) );
  XNOR U7014 ( .A(n6148), .B(n6166), .Z(n6157) );
  XNOR U7015 ( .A(n7636), .B(n7654), .Z(n7645) );
  XNOR U7016 ( .A(n8380), .B(n8398), .Z(n8389) );
  XNOR U7017 ( .A(n10245), .B(n10367), .Z(n10253) );
  XNOR U7018 ( .A(n11149), .B(n10778), .Z(n10780) );
  XOR U7019 ( .A(n23660), .B(n23747), .Z(n23666) );
  XNOR U7020 ( .A(n2806), .B(n2813), .Z(n2802) );
  XOR U7021 ( .A(n7265), .B(n7278), .Z(n7273) );
  XOR U7022 ( .A(n9497), .B(n9510), .Z(n9505) );
  XOR U7023 ( .A(n11517), .B(n11524), .Z(n11522) );
  XOR U7024 ( .A(n12253), .B(n12260), .Z(n12258) );
  XOR U7025 ( .A(n12621), .B(n12628), .Z(n12626) );
  XOR U7026 ( .A(n13357), .B(n13364), .Z(n13362) );
  XOR U7027 ( .A(n13725), .B(n13732), .Z(n13730) );
  XOR U7028 ( .A(n14461), .B(n14468), .Z(n14466) );
  XOR U7029 ( .A(n14829), .B(n14836), .Z(n14834) );
  XOR U7030 ( .A(n15565), .B(n15572), .Z(n15570) );
  XOR U7031 ( .A(n15933), .B(n15940), .Z(n15938) );
  XOR U7032 ( .A(n16669), .B(n16676), .Z(n16674) );
  XOR U7033 ( .A(n17037), .B(n17044), .Z(n17042) );
  XOR U7034 ( .A(n17773), .B(n17780), .Z(n17778) );
  XOR U7035 ( .A(n18141), .B(n18148), .Z(n18146) );
  XOR U7036 ( .A(n18877), .B(n18884), .Z(n18882) );
  XOR U7037 ( .A(n19245), .B(n19252), .Z(n19250) );
  XOR U7038 ( .A(n19981), .B(n19988), .Z(n19986) );
  XOR U7039 ( .A(n20349), .B(n20356), .Z(n20354) );
  XOR U7040 ( .A(n21085), .B(n21092), .Z(n21090) );
  XOR U7041 ( .A(n21453), .B(n21460), .Z(n21458) );
  XOR U7042 ( .A(n22189), .B(n22196), .Z(n22194) );
  XOR U7043 ( .A(n22557), .B(n22564), .Z(n22562) );
  XOR U7044 ( .A(n23293), .B(n23300), .Z(n23298) );
  XOR U7045 ( .A(n5035), .B(n5034), .Z(n4676) );
  XNOR U7046 ( .A(n31932), .B(n31929), .Z(n31931) );
  NANDN U7047 ( .A(n1691), .B(n1692), .Z(n1319) );
  NANDN U7048 ( .A(n3181), .B(n3182), .Z(n2808) );
  NANDN U7049 ( .A(n4669), .B(n4670), .Z(n4297) );
  XOR U7050 ( .A(n5421), .B(n5786), .Z(n5788) );
  XOR U7051 ( .A(n6536), .B(n6902), .Z(n6904) );
  XNOR U7052 ( .A(n8018), .B(n8020), .Z(n8019) );
  XNOR U7053 ( .A(n9134), .B(n9136), .Z(n9135) );
  NANDN U7054 ( .A(n4), .B(n3), .Z(n1) );
  XOR U7055 ( .A(n10268), .B(n9), .Z(n10267) );
  XOR U7056 ( .A(n10277), .B(n15), .Z(n10276) );
  XOR U7057 ( .A(n10286), .B(n21), .Z(n10285) );
  XOR U7058 ( .A(n10295), .B(n27), .Z(n10294) );
  XOR U7059 ( .A(n10304), .B(n33), .Z(n10303) );
  XOR U7060 ( .A(n10313), .B(n39), .Z(n10312) );
  XOR U7061 ( .A(n10322), .B(n45), .Z(n10321) );
  XOR U7062 ( .A(n10331), .B(n51), .Z(n10330) );
  XOR U7063 ( .A(n10340), .B(n57), .Z(n10339) );
  XOR U7064 ( .A(n10349), .B(n63), .Z(n10348) );
  XOR U7065 ( .A(n10358), .B(n69), .Z(n10357) );
  XNOR U7066 ( .A(n1), .B(n2), .Z(swire[99]) );
  XOR U7067 ( .A(n3), .B(n4), .Z(swire[98]) );
  XNOR U7068 ( .A(n5), .B(n6), .Z(swire[97]) );
  XNOR U7069 ( .A(n7), .B(n8), .Z(swire[96]) );
  XNOR U7070 ( .A(n9), .B(n10), .Z(swire[95]) );
  XNOR U7071 ( .A(n11), .B(n12), .Z(swire[94]) );
  XNOR U7072 ( .A(n13), .B(n14), .Z(swire[93]) );
  XNOR U7073 ( .A(n15), .B(n16), .Z(swire[92]) );
  XNOR U7074 ( .A(n17), .B(n18), .Z(swire[91]) );
  XNOR U7075 ( .A(n19), .B(n20), .Z(swire[90]) );
  XNOR U7076 ( .A(n21), .B(n22), .Z(swire[89]) );
  XNOR U7077 ( .A(n23), .B(n24), .Z(swire[88]) );
  XNOR U7078 ( .A(n25), .B(n26), .Z(swire[87]) );
  XNOR U7079 ( .A(n27), .B(n28), .Z(swire[86]) );
  XNOR U7080 ( .A(n29), .B(n30), .Z(swire[85]) );
  XNOR U7081 ( .A(n31), .B(n32), .Z(swire[84]) );
  XNOR U7082 ( .A(n33), .B(n34), .Z(swire[83]) );
  XNOR U7083 ( .A(n35), .B(n36), .Z(swire[82]) );
  XNOR U7084 ( .A(n37), .B(n38), .Z(swire[81]) );
  XNOR U7085 ( .A(n39), .B(n40), .Z(swire[80]) );
  XNOR U7086 ( .A(n41), .B(n42), .Z(swire[79]) );
  XNOR U7087 ( .A(n43), .B(n44), .Z(swire[78]) );
  XNOR U7088 ( .A(n45), .B(n46), .Z(swire[77]) );
  XNOR U7089 ( .A(n47), .B(n48), .Z(swire[76]) );
  XNOR U7090 ( .A(n49), .B(n50), .Z(swire[75]) );
  XNOR U7091 ( .A(n51), .B(n52), .Z(swire[74]) );
  XNOR U7092 ( .A(n53), .B(n54), .Z(swire[73]) );
  XNOR U7093 ( .A(n55), .B(n56), .Z(swire[72]) );
  XNOR U7094 ( .A(n57), .B(n58), .Z(swire[71]) );
  XNOR U7095 ( .A(n59), .B(n60), .Z(swire[70]) );
  XNOR U7096 ( .A(n61), .B(n62), .Z(swire[69]) );
  XNOR U7097 ( .A(n63), .B(n64), .Z(swire[68]) );
  XNOR U7098 ( .A(n65), .B(n66), .Z(swire[67]) );
  XNOR U7099 ( .A(n67), .B(n68), .Z(swire[66]) );
  XNOR U7100 ( .A(n69), .B(n70), .Z(swire[65]) );
  XNOR U7101 ( .A(n71), .B(n72), .Z(swire[64]) );
  XOR U7102 ( .A(n73), .B(n74), .Z(swire[127]) );
  XOR U7103 ( .A(n75), .B(n76), .Z(n74) );
  XOR U7104 ( .A(n77), .B(n78), .Z(n76) );
  XOR U7105 ( .A(n79), .B(n80), .Z(n78) );
  XOR U7106 ( .A(n81), .B(n82), .Z(n80) );
  XOR U7107 ( .A(n83), .B(n84), .Z(n82) );
  AND U7108 ( .A(b[3]), .B(a[124]), .Z(n84) );
  AND U7109 ( .A(b[4]), .B(a[123]), .Z(n83) );
  XOR U7110 ( .A(n85), .B(n86), .Z(n81) );
  XOR U7111 ( .A(n87), .B(n88), .Z(n86) );
  XOR U7112 ( .A(n89), .B(n90), .Z(n88) );
  AND U7113 ( .A(b[9]), .B(a[118]), .Z(n90) );
  AND U7114 ( .A(b[10]), .B(a[117]), .Z(n89) );
  XOR U7115 ( .A(n91), .B(n92), .Z(n87) );
  XOR U7116 ( .A(n93), .B(n94), .Z(n92) );
  XOR U7117 ( .A(n95), .B(n96), .Z(n94) );
  AND U7118 ( .A(b[15]), .B(a[112]), .Z(n96) );
  AND U7119 ( .A(b[16]), .B(a[111]), .Z(n95) );
  XOR U7120 ( .A(n97), .B(n98), .Z(n93) );
  XOR U7121 ( .A(n99), .B(n100), .Z(n98) );
  XOR U7122 ( .A(n101), .B(n102), .Z(n100) );
  XOR U7123 ( .A(n103), .B(n104), .Z(n102) );
  XOR U7124 ( .A(n105), .B(n106), .Z(n104) );
  XOR U7125 ( .A(n107), .B(n108), .Z(n106) );
  XOR U7126 ( .A(n109), .B(n110), .Z(n108) );
  XOR U7127 ( .A(n111), .B(n112), .Z(n110) );
  XOR U7128 ( .A(n113), .B(n114), .Z(n112) );
  XOR U7129 ( .A(n115), .B(n116), .Z(n114) );
  XOR U7130 ( .A(n117), .B(n118), .Z(n116) );
  XOR U7131 ( .A(n119), .B(n120), .Z(n118) );
  XOR U7132 ( .A(n121), .B(n122), .Z(n120) );
  XOR U7133 ( .A(n123), .B(n124), .Z(n122) );
  XOR U7134 ( .A(n125), .B(n126), .Z(n124) );
  AND U7135 ( .A(b[45]), .B(a[82]), .Z(n126) );
  AND U7136 ( .A(b[51]), .B(a[76]), .Z(n125) );
  XOR U7137 ( .A(n127), .B(n128), .Z(n123) );
  XOR U7138 ( .A(n129), .B(n130), .Z(n128) );
  XOR U7139 ( .A(n131), .B(n132), .Z(n130) );
  XOR U7140 ( .A(n133), .B(n134), .Z(n132) );
  AND U7141 ( .A(b[52]), .B(a[75]), .Z(n134) );
  AND U7142 ( .A(b[57]), .B(a[70]), .Z(n133) );
  XOR U7143 ( .A(n135), .B(n136), .Z(n131) );
  AND U7144 ( .A(b[58]), .B(a[69]), .Z(n136) );
  AND U7145 ( .A(b[59]), .B(a[68]), .Z(n135) );
  XOR U7146 ( .A(n137), .B(n138), .Z(n129) );
  XOR U7147 ( .A(n139), .B(n140), .Z(n138) );
  AND U7148 ( .A(b[60]), .B(a[67]), .Z(n140) );
  AND U7149 ( .A(b[61]), .B(a[66]), .Z(n139) );
  XOR U7150 ( .A(n141), .B(n142), .Z(n137) );
  AND U7151 ( .A(b[62]), .B(a[65]), .Z(n142) );
  AND U7152 ( .A(b[63]), .B(a[64]), .Z(n141) );
  AND U7153 ( .A(b[46]), .B(a[81]), .Z(n127) );
  XOR U7154 ( .A(n143), .B(n144), .Z(n121) );
  XOR U7155 ( .A(n145), .B(n146), .Z(n144) );
  AND U7156 ( .A(b[53]), .B(a[74]), .Z(n146) );
  AND U7157 ( .A(b[54]), .B(a[73]), .Z(n145) );
  XOR U7158 ( .A(n147), .B(n148), .Z(n143) );
  AND U7159 ( .A(b[55]), .B(a[72]), .Z(n148) );
  AND U7160 ( .A(b[56]), .B(a[71]), .Z(n147) );
  AND U7161 ( .A(b[40]), .B(a[87]), .Z(n119) );
  AND U7162 ( .A(b[39]), .B(a[88]), .Z(n117) );
  XOR U7163 ( .A(n149), .B(n150), .Z(n115) );
  XOR U7164 ( .A(n151), .B(n152), .Z(n150) );
  AND U7165 ( .A(b[47]), .B(a[80]), .Z(n152) );
  AND U7166 ( .A(b[48]), .B(a[79]), .Z(n151) );
  XOR U7167 ( .A(n153), .B(n154), .Z(n149) );
  AND U7168 ( .A(b[49]), .B(a[78]), .Z(n154) );
  AND U7169 ( .A(b[50]), .B(a[77]), .Z(n153) );
  AND U7170 ( .A(b[34]), .B(a[93]), .Z(n113) );
  AND U7171 ( .A(b[33]), .B(a[94]), .Z(n111) );
  XOR U7172 ( .A(n155), .B(n156), .Z(n109) );
  XOR U7173 ( .A(n157), .B(n158), .Z(n156) );
  AND U7174 ( .A(b[41]), .B(a[86]), .Z(n158) );
  AND U7175 ( .A(b[42]), .B(a[85]), .Z(n157) );
  XOR U7176 ( .A(n159), .B(n160), .Z(n155) );
  AND U7177 ( .A(b[43]), .B(a[84]), .Z(n160) );
  AND U7178 ( .A(b[44]), .B(a[83]), .Z(n159) );
  AND U7179 ( .A(b[28]), .B(a[99]), .Z(n107) );
  AND U7180 ( .A(b[27]), .B(a[100]), .Z(n105) );
  XOR U7181 ( .A(n161), .B(n162), .Z(n103) );
  XOR U7182 ( .A(n163), .B(n164), .Z(n162) );
  AND U7183 ( .A(b[35]), .B(a[92]), .Z(n164) );
  AND U7184 ( .A(b[36]), .B(a[91]), .Z(n163) );
  XOR U7185 ( .A(n165), .B(n166), .Z(n161) );
  AND U7186 ( .A(b[37]), .B(a[90]), .Z(n166) );
  AND U7187 ( .A(b[38]), .B(a[89]), .Z(n165) );
  AND U7188 ( .A(b[22]), .B(a[105]), .Z(n101) );
  AND U7189 ( .A(b[21]), .B(a[106]), .Z(n99) );
  XOR U7190 ( .A(n167), .B(n168), .Z(n97) );
  XOR U7191 ( .A(n169), .B(n170), .Z(n168) );
  AND U7192 ( .A(b[29]), .B(a[98]), .Z(n170) );
  AND U7193 ( .A(b[30]), .B(a[97]), .Z(n169) );
  XOR U7194 ( .A(n171), .B(n172), .Z(n167) );
  AND U7195 ( .A(b[31]), .B(a[96]), .Z(n172) );
  AND U7196 ( .A(b[32]), .B(a[95]), .Z(n171) );
  XOR U7197 ( .A(n173), .B(n174), .Z(n91) );
  XOR U7198 ( .A(n175), .B(n176), .Z(n174) );
  AND U7199 ( .A(b[23]), .B(a[104]), .Z(n176) );
  AND U7200 ( .A(b[24]), .B(a[103]), .Z(n175) );
  XOR U7201 ( .A(n177), .B(n178), .Z(n173) );
  AND U7202 ( .A(b[25]), .B(a[102]), .Z(n178) );
  AND U7203 ( .A(b[26]), .B(a[101]), .Z(n177) );
  XOR U7204 ( .A(n179), .B(n180), .Z(n85) );
  XOR U7205 ( .A(n181), .B(n182), .Z(n180) );
  AND U7206 ( .A(b[17]), .B(a[110]), .Z(n182) );
  AND U7207 ( .A(b[18]), .B(a[109]), .Z(n181) );
  XOR U7208 ( .A(n183), .B(n184), .Z(n179) );
  AND U7209 ( .A(b[19]), .B(a[108]), .Z(n184) );
  AND U7210 ( .A(b[20]), .B(a[107]), .Z(n183) );
  XOR U7211 ( .A(n185), .B(n186), .Z(n79) );
  XOR U7212 ( .A(n187), .B(n188), .Z(n186) );
  AND U7213 ( .A(b[11]), .B(a[116]), .Z(n188) );
  AND U7214 ( .A(b[12]), .B(a[115]), .Z(n187) );
  XOR U7215 ( .A(n189), .B(n190), .Z(n185) );
  AND U7216 ( .A(b[13]), .B(a[114]), .Z(n190) );
  AND U7217 ( .A(b[14]), .B(a[113]), .Z(n189) );
  AND U7218 ( .A(a[127]), .B(b[0]), .Z(n77) );
  XOR U7219 ( .A(n191), .B(n192), .Z(n75) );
  AND U7220 ( .A(b[1]), .B(a[126]), .Z(n192) );
  AND U7221 ( .A(b[2]), .B(a[125]), .Z(n191) );
  XOR U7222 ( .A(n193), .B(n194), .Z(n73) );
  XOR U7223 ( .A(n195), .B(n196), .Z(n194) );
  AND U7224 ( .A(b[5]), .B(a[122]), .Z(n196) );
  AND U7225 ( .A(b[6]), .B(a[121]), .Z(n195) );
  XOR U7226 ( .A(n197), .B(n198), .Z(n193) );
  AND U7227 ( .A(b[7]), .B(a[120]), .Z(n198) );
  AND U7228 ( .A(b[8]), .B(a[119]), .Z(n197) );
  XOR U7229 ( .A(n199), .B(n200), .Z(swire[126]) );
  XOR U7230 ( .A(n201), .B(n202), .Z(n200) );
  XOR U7231 ( .A(n203), .B(n204), .Z(n202) );
  XOR U7232 ( .A(n205), .B(n206), .Z(n204) );
  XOR U7233 ( .A(n207), .B(n208), .Z(n206) );
  XOR U7234 ( .A(n209), .B(n210), .Z(n208) );
  AND U7235 ( .A(b[3]), .B(a[123]), .Z(n209) );
  XOR U7236 ( .A(n211), .B(n212), .Z(n207) );
  XOR U7237 ( .A(n213), .B(n214), .Z(n212) );
  XOR U7238 ( .A(n215), .B(n216), .Z(n214) );
  XOR U7239 ( .A(n217), .B(n218), .Z(n216) );
  AND U7240 ( .A(b[9]), .B(a[117]), .Z(n217) );
  XOR U7241 ( .A(n219), .B(n220), .Z(n215) );
  XOR U7242 ( .A(n221), .B(n222), .Z(n220) );
  XOR U7243 ( .A(n223), .B(n224), .Z(n222) );
  XOR U7244 ( .A(n225), .B(n223), .Z(n224) );
  AND U7245 ( .A(b[15]), .B(a[111]), .Z(n225) );
  XOR U7246 ( .A(n226), .B(n227), .Z(n223) );
  ANDN U7247 ( .B(n228), .A(n229), .Z(n226) );
  XOR U7248 ( .A(n230), .B(n231), .Z(n221) );
  XOR U7249 ( .A(n232), .B(n233), .Z(n231) );
  AND U7250 ( .A(b[20]), .B(a[106]), .Z(n232) );
  XOR U7251 ( .A(n233), .B(n234), .Z(n230) );
  XOR U7252 ( .A(n235), .B(n236), .Z(n234) );
  XOR U7253 ( .A(n237), .B(n238), .Z(n236) );
  XOR U7254 ( .A(n239), .B(n240), .Z(n238) );
  XOR U7255 ( .A(n241), .B(n239), .Z(n240) );
  AND U7256 ( .A(b[21]), .B(a[105]), .Z(n241) );
  XOR U7257 ( .A(n242), .B(n243), .Z(n239) );
  ANDN U7258 ( .B(n244), .A(n245), .Z(n242) );
  XOR U7259 ( .A(n246), .B(n247), .Z(n237) );
  XOR U7260 ( .A(n248), .B(n249), .Z(n247) );
  AND U7261 ( .A(b[26]), .B(a[100]), .Z(n248) );
  XOR U7262 ( .A(n249), .B(n250), .Z(n246) );
  XOR U7263 ( .A(n251), .B(n252), .Z(n250) );
  XOR U7264 ( .A(n253), .B(n254), .Z(n252) );
  XOR U7265 ( .A(n255), .B(n256), .Z(n254) );
  XOR U7266 ( .A(n257), .B(n255), .Z(n256) );
  AND U7267 ( .A(b[27]), .B(a[99]), .Z(n257) );
  XOR U7268 ( .A(n258), .B(n259), .Z(n255) );
  ANDN U7269 ( .B(n260), .A(n261), .Z(n258) );
  XOR U7270 ( .A(n262), .B(n263), .Z(n253) );
  XOR U7271 ( .A(n264), .B(n265), .Z(n263) );
  AND U7272 ( .A(b[32]), .B(a[94]), .Z(n264) );
  XOR U7273 ( .A(n265), .B(n266), .Z(n262) );
  XOR U7274 ( .A(n267), .B(n268), .Z(n266) );
  XOR U7275 ( .A(n269), .B(n270), .Z(n268) );
  XOR U7276 ( .A(n271), .B(n272), .Z(n270) );
  XOR U7277 ( .A(n273), .B(n271), .Z(n272) );
  AND U7278 ( .A(b[33]), .B(a[93]), .Z(n273) );
  XOR U7279 ( .A(n274), .B(n275), .Z(n271) );
  ANDN U7280 ( .B(n276), .A(n277), .Z(n274) );
  XOR U7281 ( .A(n278), .B(n279), .Z(n269) );
  XOR U7282 ( .A(n280), .B(n281), .Z(n279) );
  AND U7283 ( .A(b[38]), .B(a[88]), .Z(n280) );
  XOR U7284 ( .A(n281), .B(n282), .Z(n278) );
  XOR U7285 ( .A(n283), .B(n284), .Z(n282) );
  XOR U7286 ( .A(n285), .B(n286), .Z(n284) );
  XOR U7287 ( .A(n287), .B(n288), .Z(n286) );
  XOR U7288 ( .A(n289), .B(n287), .Z(n288) );
  AND U7289 ( .A(b[39]), .B(a[87]), .Z(n289) );
  XOR U7290 ( .A(n290), .B(n291), .Z(n287) );
  ANDN U7291 ( .B(n292), .A(n293), .Z(n290) );
  XOR U7292 ( .A(n294), .B(n295), .Z(n285) );
  XOR U7293 ( .A(n296), .B(n297), .Z(n295) );
  AND U7294 ( .A(b[44]), .B(a[82]), .Z(n296) );
  XOR U7295 ( .A(n297), .B(n298), .Z(n294) );
  XOR U7296 ( .A(n299), .B(n300), .Z(n298) );
  XOR U7297 ( .A(n301), .B(n302), .Z(n300) );
  XOR U7298 ( .A(n303), .B(n304), .Z(n302) );
  XOR U7299 ( .A(n305), .B(n303), .Z(n304) );
  AND U7300 ( .A(b[45]), .B(a[81]), .Z(n305) );
  XOR U7301 ( .A(n306), .B(n307), .Z(n303) );
  ANDN U7302 ( .B(n308), .A(n309), .Z(n306) );
  XOR U7303 ( .A(n310), .B(n311), .Z(n301) );
  XOR U7304 ( .A(n312), .B(n313), .Z(n311) );
  AND U7305 ( .A(b[50]), .B(a[76]), .Z(n312) );
  XOR U7306 ( .A(n313), .B(n314), .Z(n310) );
  XOR U7307 ( .A(n315), .B(n316), .Z(n314) );
  XOR U7308 ( .A(n317), .B(n318), .Z(n316) );
  XOR U7309 ( .A(n319), .B(n320), .Z(n318) );
  XOR U7310 ( .A(n321), .B(n319), .Z(n320) );
  AND U7311 ( .A(b[51]), .B(a[75]), .Z(n321) );
  XOR U7312 ( .A(n322), .B(n323), .Z(n319) );
  ANDN U7313 ( .B(n324), .A(n325), .Z(n322) );
  XOR U7314 ( .A(n326), .B(n327), .Z(n317) );
  XOR U7315 ( .A(n328), .B(n329), .Z(n327) );
  AND U7316 ( .A(b[56]), .B(a[70]), .Z(n328) );
  XOR U7317 ( .A(n329), .B(n330), .Z(n326) );
  XOR U7318 ( .A(n331), .B(n332), .Z(n330) );
  XOR U7319 ( .A(n333), .B(n334), .Z(n332) );
  XOR U7320 ( .A(n335), .B(n336), .Z(n334) );
  XOR U7321 ( .A(n337), .B(n335), .Z(n336) );
  AND U7322 ( .A(b[57]), .B(a[69]), .Z(n337) );
  XOR U7323 ( .A(n338), .B(n339), .Z(n335) );
  ANDN U7324 ( .B(n340), .A(n341), .Z(n338) );
  XOR U7325 ( .A(n342), .B(n343), .Z(n333) );
  AND U7326 ( .A(b[58]), .B(a[68]), .Z(n343) );
  AND U7327 ( .A(b[59]), .B(a[67]), .Z(n342) );
  XOR U7328 ( .A(n344), .B(n345), .Z(n331) );
  XOR U7329 ( .A(n346), .B(n347), .Z(n345) );
  AND U7330 ( .A(b[60]), .B(a[66]), .Z(n347) );
  AND U7331 ( .A(b[61]), .B(a[65]), .Z(n346) );
  XOR U7332 ( .A(n348), .B(n349), .Z(n344) );
  AND U7333 ( .A(b[62]), .B(a[64]), .Z(n349) );
  AND U7334 ( .A(a[63]), .B(b[63]), .Z(n348) );
  XOR U7335 ( .A(n350), .B(n351), .Z(n329) );
  AND U7336 ( .A(n352), .B(n353), .Z(n350) );
  XOR U7337 ( .A(n354), .B(n355), .Z(n315) );
  XOR U7338 ( .A(n356), .B(n357), .Z(n355) );
  AND U7339 ( .A(b[52]), .B(a[74]), .Z(n357) );
  AND U7340 ( .A(b[53]), .B(a[73]), .Z(n356) );
  XOR U7341 ( .A(n358), .B(n359), .Z(n354) );
  AND U7342 ( .A(b[54]), .B(a[72]), .Z(n359) );
  AND U7343 ( .A(b[55]), .B(a[71]), .Z(n358) );
  XOR U7344 ( .A(n360), .B(n361), .Z(n313) );
  AND U7345 ( .A(n362), .B(n363), .Z(n360) );
  XOR U7346 ( .A(n364), .B(n365), .Z(n299) );
  XOR U7347 ( .A(n366), .B(n367), .Z(n365) );
  AND U7348 ( .A(b[46]), .B(a[80]), .Z(n367) );
  AND U7349 ( .A(b[47]), .B(a[79]), .Z(n366) );
  XOR U7350 ( .A(n368), .B(n369), .Z(n364) );
  AND U7351 ( .A(b[48]), .B(a[78]), .Z(n369) );
  AND U7352 ( .A(b[49]), .B(a[77]), .Z(n368) );
  XOR U7353 ( .A(n370), .B(n371), .Z(n297) );
  AND U7354 ( .A(n372), .B(n373), .Z(n370) );
  XOR U7355 ( .A(n374), .B(n375), .Z(n283) );
  XOR U7356 ( .A(n376), .B(n377), .Z(n375) );
  AND U7357 ( .A(b[40]), .B(a[86]), .Z(n377) );
  AND U7358 ( .A(b[41]), .B(a[85]), .Z(n376) );
  XOR U7359 ( .A(n378), .B(n379), .Z(n374) );
  AND U7360 ( .A(b[42]), .B(a[84]), .Z(n379) );
  AND U7361 ( .A(b[43]), .B(a[83]), .Z(n378) );
  XOR U7362 ( .A(n380), .B(n381), .Z(n281) );
  AND U7363 ( .A(n382), .B(n383), .Z(n380) );
  XOR U7364 ( .A(n384), .B(n385), .Z(n267) );
  XOR U7365 ( .A(n386), .B(n387), .Z(n385) );
  AND U7366 ( .A(b[34]), .B(a[92]), .Z(n387) );
  AND U7367 ( .A(b[35]), .B(a[91]), .Z(n386) );
  XOR U7368 ( .A(n388), .B(n389), .Z(n384) );
  AND U7369 ( .A(b[36]), .B(a[90]), .Z(n389) );
  AND U7370 ( .A(b[37]), .B(a[89]), .Z(n388) );
  XOR U7371 ( .A(n390), .B(n391), .Z(n265) );
  AND U7372 ( .A(n392), .B(n393), .Z(n390) );
  XOR U7373 ( .A(n394), .B(n395), .Z(n251) );
  XOR U7374 ( .A(n396), .B(n397), .Z(n395) );
  AND U7375 ( .A(b[28]), .B(a[98]), .Z(n397) );
  AND U7376 ( .A(b[29]), .B(a[97]), .Z(n396) );
  XOR U7377 ( .A(n398), .B(n399), .Z(n394) );
  AND U7378 ( .A(b[30]), .B(a[96]), .Z(n399) );
  AND U7379 ( .A(b[31]), .B(a[95]), .Z(n398) );
  XOR U7380 ( .A(n400), .B(n401), .Z(n249) );
  AND U7381 ( .A(n402), .B(n403), .Z(n400) );
  XOR U7382 ( .A(n404), .B(n405), .Z(n235) );
  XOR U7383 ( .A(n406), .B(n407), .Z(n405) );
  AND U7384 ( .A(b[22]), .B(a[104]), .Z(n407) );
  AND U7385 ( .A(b[23]), .B(a[103]), .Z(n406) );
  XOR U7386 ( .A(n408), .B(n409), .Z(n404) );
  AND U7387 ( .A(b[24]), .B(a[102]), .Z(n409) );
  AND U7388 ( .A(b[25]), .B(a[101]), .Z(n408) );
  XOR U7389 ( .A(n410), .B(n411), .Z(n233) );
  AND U7390 ( .A(n412), .B(n413), .Z(n410) );
  XOR U7391 ( .A(n414), .B(n415), .Z(n219) );
  XOR U7392 ( .A(n416), .B(n417), .Z(n415) );
  AND U7393 ( .A(b[16]), .B(a[110]), .Z(n417) );
  AND U7394 ( .A(b[17]), .B(a[109]), .Z(n416) );
  XOR U7395 ( .A(n418), .B(n419), .Z(n414) );
  AND U7396 ( .A(b[18]), .B(a[108]), .Z(n419) );
  AND U7397 ( .A(b[19]), .B(a[107]), .Z(n418) );
  XOR U7398 ( .A(n420), .B(n218), .Z(n213) );
  XOR U7399 ( .A(n421), .B(n422), .Z(n218) );
  ANDN U7400 ( .B(n423), .A(n424), .Z(n421) );
  AND U7401 ( .A(b[10]), .B(a[116]), .Z(n420) );
  XOR U7402 ( .A(n425), .B(n426), .Z(n211) );
  XOR U7403 ( .A(n427), .B(n428), .Z(n426) );
  AND U7404 ( .A(b[11]), .B(a[115]), .Z(n428) );
  AND U7405 ( .A(b[12]), .B(a[114]), .Z(n427) );
  XOR U7406 ( .A(n429), .B(n430), .Z(n425) );
  AND U7407 ( .A(b[13]), .B(a[113]), .Z(n430) );
  AND U7408 ( .A(b[14]), .B(a[112]), .Z(n429) );
  XOR U7409 ( .A(n431), .B(n210), .Z(n205) );
  XNOR U7410 ( .A(n432), .B(n433), .Z(n210) );
  ANDN U7411 ( .B(n434), .A(n435), .Z(n432) );
  AND U7412 ( .A(b[4]), .B(a[122]), .Z(n431) );
  XOR U7413 ( .A(n436), .B(n437), .Z(n203) );
  XOR U7414 ( .A(n438), .B(n439), .Z(n437) );
  AND U7415 ( .A(b[5]), .B(a[121]), .Z(n439) );
  AND U7416 ( .A(b[6]), .B(a[120]), .Z(n438) );
  XOR U7417 ( .A(n440), .B(n441), .Z(n436) );
  AND U7418 ( .A(b[7]), .B(a[119]), .Z(n441) );
  AND U7419 ( .A(b[8]), .B(a[118]), .Z(n440) );
  AND U7420 ( .A(a[126]), .B(b[0]), .Z(n201) );
  XOR U7421 ( .A(n442), .B(n443), .Z(n199) );
  AND U7422 ( .A(b[1]), .B(a[125]), .Z(n443) );
  AND U7423 ( .A(b[2]), .B(a[124]), .Z(n442) );
  XNOR U7424 ( .A(n444), .B(n445), .Z(swire[125]) );
  XOR U7425 ( .A(n446), .B(n447), .Z(n445) );
  XNOR U7426 ( .A(n448), .B(n444), .Z(n447) );
  AND U7427 ( .A(a[125]), .B(b[0]), .Z(n448) );
  XOR U7428 ( .A(n449), .B(n450), .Z(n446) );
  XNOR U7429 ( .A(n451), .B(n452), .Z(n450) );
  AND U7430 ( .A(b[1]), .B(a[124]), .Z(n452) );
  XNOR U7431 ( .A(n435), .B(n453), .Z(n449) );
  XNOR U7432 ( .A(n451), .B(n434), .Z(n453) );
  XNOR U7433 ( .A(n454), .B(n433), .Z(n434) );
  AND U7434 ( .A(b[2]), .B(a[123]), .Z(n454) );
  OR U7435 ( .A(n455), .B(n456), .Z(n451) );
  XOR U7436 ( .A(n457), .B(n458), .Z(n435) );
  XNOR U7437 ( .A(n433), .B(n459), .Z(n458) );
  XOR U7438 ( .A(n460), .B(n461), .Z(n459) );
  XOR U7439 ( .A(n462), .B(n463), .Z(n461) );
  XOR U7440 ( .A(n464), .B(n465), .Z(n463) );
  XOR U7441 ( .A(n466), .B(n467), .Z(n465) );
  XOR U7442 ( .A(n468), .B(n469), .Z(n467) );
  XOR U7443 ( .A(n470), .B(n471), .Z(n469) );
  XOR U7444 ( .A(n472), .B(n473), .Z(n471) );
  XOR U7445 ( .A(n474), .B(n475), .Z(n473) );
  XOR U7446 ( .A(n423), .B(n476), .Z(n475) );
  XOR U7447 ( .A(n477), .B(n424), .Z(n476) );
  XOR U7448 ( .A(n478), .B(n479), .Z(n424) );
  XOR U7449 ( .A(n422), .B(n480), .Z(n479) );
  XOR U7450 ( .A(n481), .B(n482), .Z(n480) );
  XOR U7451 ( .A(n483), .B(n484), .Z(n482) );
  XOR U7452 ( .A(n485), .B(n486), .Z(n484) );
  XOR U7453 ( .A(n487), .B(n488), .Z(n486) );
  XOR U7454 ( .A(n489), .B(n490), .Z(n488) );
  XOR U7455 ( .A(n491), .B(n492), .Z(n490) );
  XOR U7456 ( .A(n493), .B(n494), .Z(n492) );
  XOR U7457 ( .A(n495), .B(n496), .Z(n494) );
  XOR U7458 ( .A(n228), .B(n497), .Z(n496) );
  XOR U7459 ( .A(n498), .B(n229), .Z(n497) );
  XOR U7460 ( .A(n499), .B(n500), .Z(n229) );
  XOR U7461 ( .A(n227), .B(n501), .Z(n500) );
  XOR U7462 ( .A(n502), .B(n503), .Z(n501) );
  XOR U7463 ( .A(n504), .B(n505), .Z(n503) );
  XOR U7464 ( .A(n506), .B(n507), .Z(n505) );
  XOR U7465 ( .A(n508), .B(n509), .Z(n507) );
  XOR U7466 ( .A(n510), .B(n511), .Z(n509) );
  XOR U7467 ( .A(n512), .B(n513), .Z(n511) );
  XOR U7468 ( .A(n514), .B(n515), .Z(n513) );
  XNOR U7469 ( .A(n413), .B(n412), .Z(n515) );
  XOR U7470 ( .A(n516), .B(n411), .Z(n412) );
  AND U7471 ( .A(b[19]), .B(a[106]), .Z(n516) );
  XOR U7472 ( .A(n411), .B(n245), .Z(n517) );
  XOR U7473 ( .A(n518), .B(n519), .Z(n245) );
  XOR U7474 ( .A(n243), .B(n520), .Z(n519) );
  XOR U7475 ( .A(n521), .B(n522), .Z(n520) );
  XOR U7476 ( .A(n523), .B(n524), .Z(n522) );
  XOR U7477 ( .A(n525), .B(n526), .Z(n524) );
  XOR U7478 ( .A(n527), .B(n528), .Z(n526) );
  XOR U7479 ( .A(n529), .B(n530), .Z(n528) );
  XOR U7480 ( .A(n531), .B(n532), .Z(n530) );
  XOR U7481 ( .A(n533), .B(n534), .Z(n532) );
  XNOR U7482 ( .A(n403), .B(n402), .Z(n534) );
  XOR U7483 ( .A(n535), .B(n401), .Z(n402) );
  AND U7484 ( .A(b[25]), .B(a[100]), .Z(n535) );
  XOR U7485 ( .A(n401), .B(n261), .Z(n536) );
  XOR U7486 ( .A(n537), .B(n538), .Z(n261) );
  XOR U7487 ( .A(n259), .B(n539), .Z(n538) );
  XOR U7488 ( .A(n540), .B(n541), .Z(n539) );
  XOR U7489 ( .A(n542), .B(n543), .Z(n541) );
  XOR U7490 ( .A(n544), .B(n545), .Z(n543) );
  XOR U7491 ( .A(n546), .B(n547), .Z(n545) );
  XOR U7492 ( .A(n548), .B(n549), .Z(n547) );
  XOR U7493 ( .A(n550), .B(n551), .Z(n549) );
  XOR U7494 ( .A(n552), .B(n553), .Z(n551) );
  XNOR U7495 ( .A(n393), .B(n392), .Z(n553) );
  XOR U7496 ( .A(n554), .B(n391), .Z(n392) );
  AND U7497 ( .A(b[31]), .B(a[94]), .Z(n554) );
  XOR U7498 ( .A(n391), .B(n277), .Z(n555) );
  XOR U7499 ( .A(n556), .B(n557), .Z(n277) );
  XOR U7500 ( .A(n275), .B(n558), .Z(n557) );
  XOR U7501 ( .A(n559), .B(n560), .Z(n558) );
  XOR U7502 ( .A(n561), .B(n562), .Z(n560) );
  XOR U7503 ( .A(n563), .B(n564), .Z(n562) );
  XOR U7504 ( .A(n565), .B(n566), .Z(n564) );
  XOR U7505 ( .A(n567), .B(n568), .Z(n566) );
  XOR U7506 ( .A(n569), .B(n570), .Z(n568) );
  XOR U7507 ( .A(n571), .B(n572), .Z(n570) );
  XNOR U7508 ( .A(n383), .B(n382), .Z(n572) );
  XOR U7509 ( .A(n573), .B(n381), .Z(n382) );
  AND U7510 ( .A(b[37]), .B(a[88]), .Z(n573) );
  XOR U7511 ( .A(n381), .B(n293), .Z(n574) );
  XOR U7512 ( .A(n575), .B(n576), .Z(n293) );
  XOR U7513 ( .A(n291), .B(n577), .Z(n576) );
  XOR U7514 ( .A(n578), .B(n579), .Z(n577) );
  XOR U7515 ( .A(n580), .B(n581), .Z(n579) );
  XOR U7516 ( .A(n582), .B(n583), .Z(n581) );
  XOR U7517 ( .A(n584), .B(n585), .Z(n583) );
  XOR U7518 ( .A(n586), .B(n587), .Z(n585) );
  XOR U7519 ( .A(n588), .B(n589), .Z(n587) );
  XOR U7520 ( .A(n590), .B(n591), .Z(n589) );
  XNOR U7521 ( .A(n373), .B(n372), .Z(n591) );
  XOR U7522 ( .A(n592), .B(n371), .Z(n372) );
  AND U7523 ( .A(b[43]), .B(a[82]), .Z(n592) );
  XOR U7524 ( .A(n371), .B(n309), .Z(n593) );
  XOR U7525 ( .A(n594), .B(n595), .Z(n309) );
  XOR U7526 ( .A(n307), .B(n596), .Z(n595) );
  XOR U7527 ( .A(n597), .B(n598), .Z(n596) );
  XOR U7528 ( .A(n599), .B(n600), .Z(n598) );
  XOR U7529 ( .A(n601), .B(n602), .Z(n600) );
  XOR U7530 ( .A(n603), .B(n604), .Z(n602) );
  XOR U7531 ( .A(n605), .B(n606), .Z(n604) );
  XOR U7532 ( .A(n607), .B(n608), .Z(n606) );
  XOR U7533 ( .A(n609), .B(n610), .Z(n608) );
  XNOR U7534 ( .A(n363), .B(n362), .Z(n610) );
  XOR U7535 ( .A(n611), .B(n361), .Z(n362) );
  AND U7536 ( .A(b[49]), .B(a[76]), .Z(n611) );
  XOR U7537 ( .A(n361), .B(n325), .Z(n612) );
  XOR U7538 ( .A(n613), .B(n614), .Z(n325) );
  XOR U7539 ( .A(n323), .B(n615), .Z(n614) );
  XOR U7540 ( .A(n616), .B(n617), .Z(n615) );
  XOR U7541 ( .A(n618), .B(n619), .Z(n617) );
  XOR U7542 ( .A(n620), .B(n621), .Z(n619) );
  XOR U7543 ( .A(n622), .B(n623), .Z(n621) );
  XOR U7544 ( .A(n624), .B(n625), .Z(n623) );
  XOR U7545 ( .A(n626), .B(n627), .Z(n625) );
  XOR U7546 ( .A(n628), .B(n629), .Z(n627) );
  XNOR U7547 ( .A(n353), .B(n352), .Z(n629) );
  XOR U7548 ( .A(n630), .B(n351), .Z(n352) );
  AND U7549 ( .A(b[55]), .B(a[70]), .Z(n630) );
  XOR U7550 ( .A(n351), .B(n341), .Z(n631) );
  XOR U7551 ( .A(n632), .B(n633), .Z(n341) );
  XOR U7552 ( .A(n339), .B(n634), .Z(n633) );
  XOR U7553 ( .A(n635), .B(n636), .Z(n634) );
  XOR U7554 ( .A(n637), .B(n638), .Z(n636) );
  XOR U7555 ( .A(n639), .B(n640), .Z(n638) );
  XOR U7556 ( .A(n641), .B(n642), .Z(n640) );
  XOR U7557 ( .A(n643), .B(n644), .Z(n642) );
  XOR U7558 ( .A(n645), .B(n646), .Z(n644) );
  XOR U7559 ( .A(n647), .B(n648), .Z(n646) );
  XOR U7560 ( .A(n649), .B(n650), .Z(n648) );
  XOR U7561 ( .A(n651), .B(n652), .Z(n650) );
  XOR U7562 ( .A(n653), .B(n654), .Z(n652) );
  NAND U7563 ( .A(b[62]), .B(a[63]), .Z(n654) );
  AND U7564 ( .A(a[62]), .B(b[63]), .Z(n653) );
  XOR U7565 ( .A(n655), .B(n651), .Z(n647) );
  XOR U7566 ( .A(n656), .B(n657), .Z(n651) );
  ANDN U7567 ( .B(n658), .A(n659), .Z(n656) );
  AND U7568 ( .A(b[61]), .B(a[64]), .Z(n655) );
  XOR U7569 ( .A(n660), .B(n649), .Z(n643) );
  XOR U7570 ( .A(n661), .B(n662), .Z(n649) );
  AND U7571 ( .A(n663), .B(n664), .Z(n661) );
  AND U7572 ( .A(b[60]), .B(a[65]), .Z(n660) );
  XOR U7573 ( .A(n665), .B(n645), .Z(n639) );
  XOR U7574 ( .A(n666), .B(n667), .Z(n645) );
  AND U7575 ( .A(n668), .B(n669), .Z(n666) );
  AND U7576 ( .A(b[59]), .B(a[66]), .Z(n665) );
  XOR U7577 ( .A(n670), .B(n641), .Z(n635) );
  XOR U7578 ( .A(n671), .B(n672), .Z(n641) );
  AND U7579 ( .A(n673), .B(n674), .Z(n671) );
  AND U7580 ( .A(b[58]), .B(a[67]), .Z(n670) );
  XOR U7581 ( .A(n675), .B(n637), .Z(n632) );
  XOR U7582 ( .A(n676), .B(n677), .Z(n637) );
  AND U7583 ( .A(n678), .B(n679), .Z(n676) );
  AND U7584 ( .A(b[57]), .B(a[68]), .Z(n675) );
  XOR U7585 ( .A(n680), .B(n681), .Z(n351) );
  AND U7586 ( .A(n682), .B(n683), .Z(n680) );
  XOR U7587 ( .A(n684), .B(n339), .Z(n340) );
  XOR U7588 ( .A(n685), .B(n686), .Z(n339) );
  AND U7589 ( .A(n687), .B(n688), .Z(n685) );
  AND U7590 ( .A(b[56]), .B(a[69]), .Z(n684) );
  XOR U7591 ( .A(n689), .B(n628), .Z(n624) );
  XOR U7592 ( .A(n690), .B(n691), .Z(n628) );
  AND U7593 ( .A(n692), .B(n693), .Z(n690) );
  AND U7594 ( .A(b[54]), .B(a[71]), .Z(n689) );
  XOR U7595 ( .A(n694), .B(n626), .Z(n620) );
  XOR U7596 ( .A(n695), .B(n696), .Z(n626) );
  AND U7597 ( .A(n697), .B(n698), .Z(n695) );
  AND U7598 ( .A(b[53]), .B(a[72]), .Z(n694) );
  XOR U7599 ( .A(n699), .B(n622), .Z(n616) );
  XOR U7600 ( .A(n700), .B(n701), .Z(n622) );
  AND U7601 ( .A(n702), .B(n703), .Z(n700) );
  AND U7602 ( .A(b[52]), .B(a[73]), .Z(n699) );
  XOR U7603 ( .A(n704), .B(n618), .Z(n613) );
  XOR U7604 ( .A(n705), .B(n706), .Z(n618) );
  AND U7605 ( .A(n707), .B(n708), .Z(n705) );
  AND U7606 ( .A(b[51]), .B(a[74]), .Z(n704) );
  XOR U7607 ( .A(n709), .B(n710), .Z(n361) );
  AND U7608 ( .A(n711), .B(n712), .Z(n709) );
  XOR U7609 ( .A(n713), .B(n323), .Z(n324) );
  XOR U7610 ( .A(n714), .B(n715), .Z(n323) );
  AND U7611 ( .A(n716), .B(n717), .Z(n714) );
  AND U7612 ( .A(b[50]), .B(a[75]), .Z(n713) );
  XOR U7613 ( .A(n718), .B(n609), .Z(n605) );
  XOR U7614 ( .A(n719), .B(n720), .Z(n609) );
  AND U7615 ( .A(n721), .B(n722), .Z(n719) );
  AND U7616 ( .A(b[48]), .B(a[77]), .Z(n718) );
  XOR U7617 ( .A(n723), .B(n607), .Z(n601) );
  XOR U7618 ( .A(n724), .B(n725), .Z(n607) );
  AND U7619 ( .A(n726), .B(n727), .Z(n724) );
  AND U7620 ( .A(b[47]), .B(a[78]), .Z(n723) );
  XOR U7621 ( .A(n728), .B(n603), .Z(n597) );
  XOR U7622 ( .A(n729), .B(n730), .Z(n603) );
  AND U7623 ( .A(n731), .B(n732), .Z(n729) );
  AND U7624 ( .A(b[46]), .B(a[79]), .Z(n728) );
  XOR U7625 ( .A(n733), .B(n599), .Z(n594) );
  XOR U7626 ( .A(n734), .B(n735), .Z(n599) );
  AND U7627 ( .A(n736), .B(n737), .Z(n734) );
  AND U7628 ( .A(b[45]), .B(a[80]), .Z(n733) );
  XOR U7629 ( .A(n738), .B(n739), .Z(n371) );
  AND U7630 ( .A(n740), .B(n741), .Z(n738) );
  XOR U7631 ( .A(n742), .B(n307), .Z(n308) );
  XOR U7632 ( .A(n743), .B(n744), .Z(n307) );
  AND U7633 ( .A(n745), .B(n746), .Z(n743) );
  AND U7634 ( .A(b[44]), .B(a[81]), .Z(n742) );
  XOR U7635 ( .A(n747), .B(n590), .Z(n586) );
  XOR U7636 ( .A(n748), .B(n749), .Z(n590) );
  AND U7637 ( .A(n750), .B(n751), .Z(n748) );
  AND U7638 ( .A(b[42]), .B(a[83]), .Z(n747) );
  XOR U7639 ( .A(n752), .B(n588), .Z(n582) );
  XOR U7640 ( .A(n753), .B(n754), .Z(n588) );
  AND U7641 ( .A(n755), .B(n756), .Z(n753) );
  AND U7642 ( .A(b[41]), .B(a[84]), .Z(n752) );
  XOR U7643 ( .A(n757), .B(n584), .Z(n578) );
  XOR U7644 ( .A(n758), .B(n759), .Z(n584) );
  AND U7645 ( .A(n760), .B(n761), .Z(n758) );
  AND U7646 ( .A(b[40]), .B(a[85]), .Z(n757) );
  XOR U7647 ( .A(n762), .B(n580), .Z(n575) );
  XOR U7648 ( .A(n763), .B(n764), .Z(n580) );
  AND U7649 ( .A(n765), .B(n766), .Z(n763) );
  AND U7650 ( .A(b[39]), .B(a[86]), .Z(n762) );
  XOR U7651 ( .A(n767), .B(n768), .Z(n381) );
  AND U7652 ( .A(n769), .B(n770), .Z(n767) );
  XOR U7653 ( .A(n771), .B(n291), .Z(n292) );
  XOR U7654 ( .A(n772), .B(n773), .Z(n291) );
  AND U7655 ( .A(n774), .B(n775), .Z(n772) );
  AND U7656 ( .A(b[38]), .B(a[87]), .Z(n771) );
  XOR U7657 ( .A(n776), .B(n571), .Z(n567) );
  XOR U7658 ( .A(n777), .B(n778), .Z(n571) );
  AND U7659 ( .A(n779), .B(n780), .Z(n777) );
  AND U7660 ( .A(b[36]), .B(a[89]), .Z(n776) );
  XOR U7661 ( .A(n781), .B(n569), .Z(n563) );
  XOR U7662 ( .A(n782), .B(n783), .Z(n569) );
  AND U7663 ( .A(n784), .B(n785), .Z(n782) );
  AND U7664 ( .A(b[35]), .B(a[90]), .Z(n781) );
  XOR U7665 ( .A(n786), .B(n565), .Z(n559) );
  XOR U7666 ( .A(n787), .B(n788), .Z(n565) );
  AND U7667 ( .A(n789), .B(n790), .Z(n787) );
  AND U7668 ( .A(b[34]), .B(a[91]), .Z(n786) );
  XOR U7669 ( .A(n791), .B(n561), .Z(n556) );
  XOR U7670 ( .A(n792), .B(n793), .Z(n561) );
  AND U7671 ( .A(n794), .B(n795), .Z(n792) );
  AND U7672 ( .A(b[33]), .B(a[92]), .Z(n791) );
  XOR U7673 ( .A(n796), .B(n797), .Z(n391) );
  AND U7674 ( .A(n798), .B(n799), .Z(n796) );
  XOR U7675 ( .A(n800), .B(n275), .Z(n276) );
  XOR U7676 ( .A(n801), .B(n802), .Z(n275) );
  AND U7677 ( .A(n803), .B(n804), .Z(n801) );
  AND U7678 ( .A(b[32]), .B(a[93]), .Z(n800) );
  XOR U7679 ( .A(n805), .B(n552), .Z(n548) );
  XOR U7680 ( .A(n806), .B(n807), .Z(n552) );
  AND U7681 ( .A(n808), .B(n809), .Z(n806) );
  AND U7682 ( .A(b[30]), .B(a[95]), .Z(n805) );
  XOR U7683 ( .A(n810), .B(n550), .Z(n544) );
  XOR U7684 ( .A(n811), .B(n812), .Z(n550) );
  AND U7685 ( .A(n813), .B(n814), .Z(n811) );
  AND U7686 ( .A(b[29]), .B(a[96]), .Z(n810) );
  XOR U7687 ( .A(n815), .B(n546), .Z(n540) );
  XOR U7688 ( .A(n816), .B(n817), .Z(n546) );
  AND U7689 ( .A(n818), .B(n819), .Z(n816) );
  AND U7690 ( .A(b[28]), .B(a[97]), .Z(n815) );
  XOR U7691 ( .A(n820), .B(n542), .Z(n537) );
  XOR U7692 ( .A(n821), .B(n822), .Z(n542) );
  AND U7693 ( .A(n823), .B(n824), .Z(n821) );
  AND U7694 ( .A(b[27]), .B(a[98]), .Z(n820) );
  XOR U7695 ( .A(n825), .B(n826), .Z(n401) );
  AND U7696 ( .A(n827), .B(n828), .Z(n825) );
  XOR U7697 ( .A(n829), .B(n259), .Z(n260) );
  XOR U7698 ( .A(n830), .B(n831), .Z(n259) );
  AND U7699 ( .A(n832), .B(n833), .Z(n830) );
  AND U7700 ( .A(b[26]), .B(a[99]), .Z(n829) );
  XOR U7701 ( .A(n834), .B(n533), .Z(n529) );
  XOR U7702 ( .A(n835), .B(n836), .Z(n533) );
  AND U7703 ( .A(n837), .B(n838), .Z(n835) );
  AND U7704 ( .A(b[24]), .B(a[101]), .Z(n834) );
  XOR U7705 ( .A(n839), .B(n531), .Z(n525) );
  XOR U7706 ( .A(n840), .B(n841), .Z(n531) );
  AND U7707 ( .A(n842), .B(n843), .Z(n840) );
  AND U7708 ( .A(b[23]), .B(a[102]), .Z(n839) );
  XOR U7709 ( .A(n844), .B(n527), .Z(n521) );
  XOR U7710 ( .A(n845), .B(n846), .Z(n527) );
  AND U7711 ( .A(n847), .B(n848), .Z(n845) );
  AND U7712 ( .A(b[22]), .B(a[103]), .Z(n844) );
  XOR U7713 ( .A(n849), .B(n523), .Z(n518) );
  XOR U7714 ( .A(n850), .B(n851), .Z(n523) );
  AND U7715 ( .A(n852), .B(n853), .Z(n850) );
  AND U7716 ( .A(b[21]), .B(a[104]), .Z(n849) );
  XOR U7717 ( .A(n854), .B(n855), .Z(n411) );
  AND U7718 ( .A(n856), .B(n857), .Z(n854) );
  XOR U7719 ( .A(n858), .B(n243), .Z(n244) );
  XOR U7720 ( .A(n859), .B(n860), .Z(n243) );
  AND U7721 ( .A(n861), .B(n862), .Z(n859) );
  AND U7722 ( .A(b[20]), .B(a[105]), .Z(n858) );
  XOR U7723 ( .A(n863), .B(n514), .Z(n510) );
  XOR U7724 ( .A(n864), .B(n865), .Z(n514) );
  AND U7725 ( .A(n866), .B(n867), .Z(n864) );
  AND U7726 ( .A(b[18]), .B(a[107]), .Z(n863) );
  XOR U7727 ( .A(n868), .B(n512), .Z(n506) );
  XOR U7728 ( .A(n869), .B(n870), .Z(n512) );
  AND U7729 ( .A(n871), .B(n872), .Z(n869) );
  AND U7730 ( .A(b[17]), .B(a[108]), .Z(n868) );
  XOR U7731 ( .A(n873), .B(n508), .Z(n502) );
  XOR U7732 ( .A(n874), .B(n875), .Z(n508) );
  AND U7733 ( .A(n876), .B(n877), .Z(n874) );
  AND U7734 ( .A(b[16]), .B(a[109]), .Z(n873) );
  XOR U7735 ( .A(n878), .B(n504), .Z(n499) );
  XOR U7736 ( .A(n879), .B(n880), .Z(n504) );
  AND U7737 ( .A(n881), .B(n882), .Z(n879) );
  AND U7738 ( .A(b[15]), .B(a[110]), .Z(n878) );
  XOR U7739 ( .A(n883), .B(n227), .Z(n228) );
  XOR U7740 ( .A(n884), .B(n885), .Z(n227) );
  AND U7741 ( .A(n886), .B(n887), .Z(n884) );
  AND U7742 ( .A(b[14]), .B(a[111]), .Z(n883) );
  XOR U7743 ( .A(n888), .B(n498), .Z(n493) );
  XOR U7744 ( .A(n889), .B(n890), .Z(n498) );
  AND U7745 ( .A(n891), .B(n892), .Z(n889) );
  AND U7746 ( .A(b[13]), .B(a[112]), .Z(n888) );
  XOR U7747 ( .A(n893), .B(n495), .Z(n489) );
  XOR U7748 ( .A(n894), .B(n895), .Z(n495) );
  AND U7749 ( .A(n896), .B(n897), .Z(n894) );
  AND U7750 ( .A(b[12]), .B(a[113]), .Z(n893) );
  XOR U7751 ( .A(n898), .B(n491), .Z(n485) );
  XOR U7752 ( .A(n899), .B(n900), .Z(n491) );
  AND U7753 ( .A(n901), .B(n902), .Z(n899) );
  AND U7754 ( .A(b[11]), .B(a[114]), .Z(n898) );
  XOR U7755 ( .A(n903), .B(n487), .Z(n481) );
  XOR U7756 ( .A(n904), .B(n905), .Z(n487) );
  AND U7757 ( .A(n906), .B(n907), .Z(n904) );
  AND U7758 ( .A(b[10]), .B(a[115]), .Z(n903) );
  XOR U7759 ( .A(n908), .B(n483), .Z(n478) );
  XOR U7760 ( .A(n909), .B(n910), .Z(n483) );
  AND U7761 ( .A(n911), .B(n912), .Z(n909) );
  AND U7762 ( .A(b[9]), .B(a[116]), .Z(n908) );
  XOR U7763 ( .A(n913), .B(n422), .Z(n423) );
  XOR U7764 ( .A(n914), .B(n915), .Z(n422) );
  AND U7765 ( .A(n916), .B(n917), .Z(n914) );
  AND U7766 ( .A(b[8]), .B(a[117]), .Z(n913) );
  XOR U7767 ( .A(n918), .B(n477), .Z(n472) );
  XOR U7768 ( .A(n919), .B(n920), .Z(n477) );
  AND U7769 ( .A(n921), .B(n922), .Z(n919) );
  AND U7770 ( .A(b[7]), .B(a[118]), .Z(n918) );
  XOR U7771 ( .A(n923), .B(n474), .Z(n468) );
  XOR U7772 ( .A(n924), .B(n925), .Z(n474) );
  AND U7773 ( .A(n926), .B(n927), .Z(n924) );
  AND U7774 ( .A(b[6]), .B(a[119]), .Z(n923) );
  XOR U7775 ( .A(n928), .B(n470), .Z(n464) );
  XOR U7776 ( .A(n929), .B(n930), .Z(n470) );
  AND U7777 ( .A(n931), .B(n932), .Z(n929) );
  AND U7778 ( .A(b[5]), .B(a[120]), .Z(n928) );
  XOR U7779 ( .A(n933), .B(n466), .Z(n460) );
  XOR U7780 ( .A(n934), .B(n935), .Z(n466) );
  AND U7781 ( .A(n936), .B(n937), .Z(n934) );
  AND U7782 ( .A(b[4]), .B(a[121]), .Z(n933) );
  XNOR U7783 ( .A(n938), .B(n939), .Z(n433) );
  NANDN U7784 ( .A(n940), .B(n941), .Z(n939) );
  XOR U7785 ( .A(n942), .B(n462), .Z(n457) );
  XNOR U7786 ( .A(n943), .B(n944), .Z(n462) );
  AND U7787 ( .A(n945), .B(n946), .Z(n943) );
  AND U7788 ( .A(b[3]), .B(a[122]), .Z(n942) );
  XOR U7789 ( .A(n947), .B(n948), .Z(swire[124]) );
  XOR U7790 ( .A(n456), .B(n949), .Z(n948) );
  XOR U7791 ( .A(n455), .B(n947), .Z(n949) );
  NAND U7792 ( .A(a[124]), .B(b[0]), .Z(n455) );
  XOR U7793 ( .A(n940), .B(n941), .Z(n456) );
  XOR U7794 ( .A(n938), .B(n950), .Z(n941) );
  NAND U7795 ( .A(b[1]), .B(a[123]), .Z(n950) );
  XOR U7796 ( .A(n946), .B(n951), .Z(n940) );
  XOR U7797 ( .A(n938), .B(n945), .Z(n951) );
  XNOR U7798 ( .A(n952), .B(n944), .Z(n945) );
  AND U7799 ( .A(b[2]), .B(a[122]), .Z(n952) );
  NANDN U7800 ( .A(n953), .B(n954), .Z(n938) );
  XOR U7801 ( .A(n944), .B(n936), .Z(n955) );
  XNOR U7802 ( .A(n935), .B(n931), .Z(n956) );
  XNOR U7803 ( .A(n930), .B(n926), .Z(n957) );
  XNOR U7804 ( .A(n925), .B(n921), .Z(n958) );
  XNOR U7805 ( .A(n920), .B(n916), .Z(n959) );
  XNOR U7806 ( .A(n915), .B(n911), .Z(n960) );
  XNOR U7807 ( .A(n910), .B(n906), .Z(n961) );
  XNOR U7808 ( .A(n905), .B(n901), .Z(n962) );
  XNOR U7809 ( .A(n900), .B(n896), .Z(n963) );
  XNOR U7810 ( .A(n895), .B(n891), .Z(n964) );
  XNOR U7811 ( .A(n890), .B(n886), .Z(n965) );
  XNOR U7812 ( .A(n885), .B(n881), .Z(n966) );
  XNOR U7813 ( .A(n880), .B(n876), .Z(n967) );
  XNOR U7814 ( .A(n875), .B(n871), .Z(n968) );
  XNOR U7815 ( .A(n870), .B(n866), .Z(n969) );
  XNOR U7816 ( .A(n857), .B(n856), .Z(n970) );
  XOR U7817 ( .A(n971), .B(n855), .Z(n856) );
  AND U7818 ( .A(b[18]), .B(a[106]), .Z(n971) );
  XNOR U7819 ( .A(n855), .B(n861), .Z(n972) );
  XNOR U7820 ( .A(n860), .B(n852), .Z(n973) );
  XNOR U7821 ( .A(n851), .B(n847), .Z(n974) );
  XNOR U7822 ( .A(n846), .B(n842), .Z(n975) );
  XNOR U7823 ( .A(n841), .B(n837), .Z(n976) );
  XNOR U7824 ( .A(n828), .B(n827), .Z(n977) );
  XOR U7825 ( .A(n978), .B(n826), .Z(n827) );
  AND U7826 ( .A(b[24]), .B(a[100]), .Z(n978) );
  XNOR U7827 ( .A(n826), .B(n832), .Z(n979) );
  XNOR U7828 ( .A(n831), .B(n823), .Z(n980) );
  XNOR U7829 ( .A(n822), .B(n818), .Z(n981) );
  XNOR U7830 ( .A(n817), .B(n813), .Z(n982) );
  XNOR U7831 ( .A(n812), .B(n808), .Z(n983) );
  XNOR U7832 ( .A(n799), .B(n798), .Z(n984) );
  XOR U7833 ( .A(n985), .B(n797), .Z(n798) );
  AND U7834 ( .A(b[30]), .B(a[94]), .Z(n985) );
  XNOR U7835 ( .A(n797), .B(n803), .Z(n986) );
  XNOR U7836 ( .A(n802), .B(n794), .Z(n987) );
  XNOR U7837 ( .A(n793), .B(n789), .Z(n988) );
  XNOR U7838 ( .A(n788), .B(n784), .Z(n989) );
  XNOR U7839 ( .A(n783), .B(n779), .Z(n990) );
  XNOR U7840 ( .A(n770), .B(n769), .Z(n991) );
  XOR U7841 ( .A(n992), .B(n768), .Z(n769) );
  AND U7842 ( .A(b[36]), .B(a[88]), .Z(n992) );
  XNOR U7843 ( .A(n768), .B(n774), .Z(n993) );
  XNOR U7844 ( .A(n773), .B(n765), .Z(n994) );
  XNOR U7845 ( .A(n764), .B(n760), .Z(n995) );
  XNOR U7846 ( .A(n759), .B(n755), .Z(n996) );
  XNOR U7847 ( .A(n754), .B(n750), .Z(n997) );
  XNOR U7848 ( .A(n741), .B(n740), .Z(n998) );
  XOR U7849 ( .A(n999), .B(n739), .Z(n740) );
  AND U7850 ( .A(b[42]), .B(a[82]), .Z(n999) );
  XNOR U7851 ( .A(n739), .B(n745), .Z(n1000) );
  XNOR U7852 ( .A(n744), .B(n736), .Z(n1001) );
  XNOR U7853 ( .A(n735), .B(n731), .Z(n1002) );
  XNOR U7854 ( .A(n730), .B(n726), .Z(n1003) );
  XNOR U7855 ( .A(n725), .B(n721), .Z(n1004) );
  XNOR U7856 ( .A(n712), .B(n711), .Z(n1005) );
  XOR U7857 ( .A(n1006), .B(n710), .Z(n711) );
  AND U7858 ( .A(b[48]), .B(a[76]), .Z(n1006) );
  XNOR U7859 ( .A(n710), .B(n716), .Z(n1007) );
  XNOR U7860 ( .A(n715), .B(n707), .Z(n1008) );
  XNOR U7861 ( .A(n706), .B(n702), .Z(n1009) );
  XNOR U7862 ( .A(n701), .B(n697), .Z(n1010) );
  XNOR U7863 ( .A(n696), .B(n692), .Z(n1011) );
  XNOR U7864 ( .A(n683), .B(n682), .Z(n1012) );
  XOR U7865 ( .A(n1013), .B(n681), .Z(n682) );
  AND U7866 ( .A(b[54]), .B(a[70]), .Z(n1013) );
  XNOR U7867 ( .A(n681), .B(n687), .Z(n1014) );
  XNOR U7868 ( .A(n686), .B(n678), .Z(n1015) );
  XNOR U7869 ( .A(n677), .B(n673), .Z(n1016) );
  XNOR U7870 ( .A(n672), .B(n668), .Z(n1017) );
  XNOR U7871 ( .A(n667), .B(n663), .Z(n1018) );
  XOR U7872 ( .A(n662), .B(n659), .Z(n1019) );
  XOR U7873 ( .A(n1020), .B(n1021), .Z(n659) );
  XOR U7874 ( .A(n657), .B(n1022), .Z(n1021) );
  XOR U7875 ( .A(n1023), .B(n1024), .Z(n1022) );
  XOR U7876 ( .A(n1025), .B(n1026), .Z(n1024) );
  NAND U7877 ( .A(a[62]), .B(b[62]), .Z(n1026) );
  AND U7878 ( .A(a[61]), .B(b[63]), .Z(n1025) );
  XOR U7879 ( .A(n1027), .B(n1023), .Z(n1020) );
  XOR U7880 ( .A(n1028), .B(n1029), .Z(n1023) );
  ANDN U7881 ( .B(n1030), .A(n1031), .Z(n1028) );
  AND U7882 ( .A(b[61]), .B(a[63]), .Z(n1027) );
  XOR U7883 ( .A(n1032), .B(n657), .Z(n658) );
  XOR U7884 ( .A(n1033), .B(n1034), .Z(n657) );
  AND U7885 ( .A(n1035), .B(n1036), .Z(n1033) );
  AND U7886 ( .A(b[60]), .B(a[64]), .Z(n1032) );
  XOR U7887 ( .A(n1037), .B(n662), .Z(n664) );
  XOR U7888 ( .A(n1038), .B(n1039), .Z(n662) );
  AND U7889 ( .A(n1040), .B(n1041), .Z(n1038) );
  AND U7890 ( .A(b[59]), .B(a[65]), .Z(n1037) );
  XOR U7891 ( .A(n1042), .B(n667), .Z(n669) );
  XOR U7892 ( .A(n1043), .B(n1044), .Z(n667) );
  AND U7893 ( .A(n1045), .B(n1046), .Z(n1043) );
  AND U7894 ( .A(b[58]), .B(a[66]), .Z(n1042) );
  XOR U7895 ( .A(n1047), .B(n672), .Z(n674) );
  XOR U7896 ( .A(n1048), .B(n1049), .Z(n672) );
  AND U7897 ( .A(n1050), .B(n1051), .Z(n1048) );
  AND U7898 ( .A(b[57]), .B(a[67]), .Z(n1047) );
  XOR U7899 ( .A(n1052), .B(n677), .Z(n679) );
  XOR U7900 ( .A(n1053), .B(n1054), .Z(n677) );
  AND U7901 ( .A(n1055), .B(n1056), .Z(n1053) );
  AND U7902 ( .A(b[56]), .B(a[68]), .Z(n1052) );
  XOR U7903 ( .A(n1057), .B(n1058), .Z(n681) );
  AND U7904 ( .A(n1059), .B(n1060), .Z(n1057) );
  XOR U7905 ( .A(n1061), .B(n686), .Z(n688) );
  XOR U7906 ( .A(n1062), .B(n1063), .Z(n686) );
  AND U7907 ( .A(n1064), .B(n1065), .Z(n1062) );
  AND U7908 ( .A(b[55]), .B(a[69]), .Z(n1061) );
  XOR U7909 ( .A(n1066), .B(n691), .Z(n693) );
  XOR U7910 ( .A(n1067), .B(n1068), .Z(n691) );
  AND U7911 ( .A(n1069), .B(n1070), .Z(n1067) );
  AND U7912 ( .A(b[53]), .B(a[71]), .Z(n1066) );
  XOR U7913 ( .A(n1071), .B(n696), .Z(n698) );
  XOR U7914 ( .A(n1072), .B(n1073), .Z(n696) );
  AND U7915 ( .A(n1074), .B(n1075), .Z(n1072) );
  AND U7916 ( .A(b[52]), .B(a[72]), .Z(n1071) );
  XOR U7917 ( .A(n1076), .B(n701), .Z(n703) );
  XOR U7918 ( .A(n1077), .B(n1078), .Z(n701) );
  AND U7919 ( .A(n1079), .B(n1080), .Z(n1077) );
  AND U7920 ( .A(b[51]), .B(a[73]), .Z(n1076) );
  XOR U7921 ( .A(n1081), .B(n706), .Z(n708) );
  XOR U7922 ( .A(n1082), .B(n1083), .Z(n706) );
  AND U7923 ( .A(n1084), .B(n1085), .Z(n1082) );
  AND U7924 ( .A(b[50]), .B(a[74]), .Z(n1081) );
  XOR U7925 ( .A(n1086), .B(n1087), .Z(n710) );
  AND U7926 ( .A(n1088), .B(n1089), .Z(n1086) );
  XOR U7927 ( .A(n1090), .B(n715), .Z(n717) );
  XOR U7928 ( .A(n1091), .B(n1092), .Z(n715) );
  AND U7929 ( .A(n1093), .B(n1094), .Z(n1091) );
  AND U7930 ( .A(b[49]), .B(a[75]), .Z(n1090) );
  XOR U7931 ( .A(n1095), .B(n720), .Z(n722) );
  XOR U7932 ( .A(n1096), .B(n1097), .Z(n720) );
  AND U7933 ( .A(n1098), .B(n1099), .Z(n1096) );
  AND U7934 ( .A(b[47]), .B(a[77]), .Z(n1095) );
  XOR U7935 ( .A(n1100), .B(n725), .Z(n727) );
  XOR U7936 ( .A(n1101), .B(n1102), .Z(n725) );
  AND U7937 ( .A(n1103), .B(n1104), .Z(n1101) );
  AND U7938 ( .A(b[46]), .B(a[78]), .Z(n1100) );
  XOR U7939 ( .A(n1105), .B(n730), .Z(n732) );
  XOR U7940 ( .A(n1106), .B(n1107), .Z(n730) );
  AND U7941 ( .A(n1108), .B(n1109), .Z(n1106) );
  AND U7942 ( .A(b[45]), .B(a[79]), .Z(n1105) );
  XOR U7943 ( .A(n1110), .B(n735), .Z(n737) );
  XOR U7944 ( .A(n1111), .B(n1112), .Z(n735) );
  AND U7945 ( .A(n1113), .B(n1114), .Z(n1111) );
  AND U7946 ( .A(b[44]), .B(a[80]), .Z(n1110) );
  XOR U7947 ( .A(n1115), .B(n1116), .Z(n739) );
  AND U7948 ( .A(n1117), .B(n1118), .Z(n1115) );
  XOR U7949 ( .A(n1119), .B(n744), .Z(n746) );
  XOR U7950 ( .A(n1120), .B(n1121), .Z(n744) );
  AND U7951 ( .A(n1122), .B(n1123), .Z(n1120) );
  AND U7952 ( .A(b[43]), .B(a[81]), .Z(n1119) );
  XOR U7953 ( .A(n1124), .B(n749), .Z(n751) );
  XOR U7954 ( .A(n1125), .B(n1126), .Z(n749) );
  AND U7955 ( .A(n1127), .B(n1128), .Z(n1125) );
  AND U7956 ( .A(b[41]), .B(a[83]), .Z(n1124) );
  XOR U7957 ( .A(n1129), .B(n754), .Z(n756) );
  XOR U7958 ( .A(n1130), .B(n1131), .Z(n754) );
  AND U7959 ( .A(n1132), .B(n1133), .Z(n1130) );
  AND U7960 ( .A(b[40]), .B(a[84]), .Z(n1129) );
  XOR U7961 ( .A(n1134), .B(n759), .Z(n761) );
  XOR U7962 ( .A(n1135), .B(n1136), .Z(n759) );
  AND U7963 ( .A(n1137), .B(n1138), .Z(n1135) );
  AND U7964 ( .A(b[39]), .B(a[85]), .Z(n1134) );
  XOR U7965 ( .A(n1139), .B(n764), .Z(n766) );
  XOR U7966 ( .A(n1140), .B(n1141), .Z(n764) );
  AND U7967 ( .A(n1142), .B(n1143), .Z(n1140) );
  AND U7968 ( .A(b[38]), .B(a[86]), .Z(n1139) );
  XOR U7969 ( .A(n1144), .B(n1145), .Z(n768) );
  AND U7970 ( .A(n1146), .B(n1147), .Z(n1144) );
  XOR U7971 ( .A(n1148), .B(n773), .Z(n775) );
  XOR U7972 ( .A(n1149), .B(n1150), .Z(n773) );
  AND U7973 ( .A(n1151), .B(n1152), .Z(n1149) );
  AND U7974 ( .A(b[37]), .B(a[87]), .Z(n1148) );
  XOR U7975 ( .A(n1153), .B(n778), .Z(n780) );
  XOR U7976 ( .A(n1154), .B(n1155), .Z(n778) );
  AND U7977 ( .A(n1156), .B(n1157), .Z(n1154) );
  AND U7978 ( .A(b[35]), .B(a[89]), .Z(n1153) );
  XOR U7979 ( .A(n1158), .B(n783), .Z(n785) );
  XOR U7980 ( .A(n1159), .B(n1160), .Z(n783) );
  AND U7981 ( .A(n1161), .B(n1162), .Z(n1159) );
  AND U7982 ( .A(b[34]), .B(a[90]), .Z(n1158) );
  XOR U7983 ( .A(n1163), .B(n788), .Z(n790) );
  XOR U7984 ( .A(n1164), .B(n1165), .Z(n788) );
  AND U7985 ( .A(n1166), .B(n1167), .Z(n1164) );
  AND U7986 ( .A(b[33]), .B(a[91]), .Z(n1163) );
  XOR U7987 ( .A(n1168), .B(n793), .Z(n795) );
  XOR U7988 ( .A(n1169), .B(n1170), .Z(n793) );
  AND U7989 ( .A(n1171), .B(n1172), .Z(n1169) );
  AND U7990 ( .A(b[32]), .B(a[92]), .Z(n1168) );
  XOR U7991 ( .A(n1173), .B(n1174), .Z(n797) );
  AND U7992 ( .A(n1175), .B(n1176), .Z(n1173) );
  XOR U7993 ( .A(n1177), .B(n802), .Z(n804) );
  XOR U7994 ( .A(n1178), .B(n1179), .Z(n802) );
  AND U7995 ( .A(n1180), .B(n1181), .Z(n1178) );
  AND U7996 ( .A(b[31]), .B(a[93]), .Z(n1177) );
  XOR U7997 ( .A(n1182), .B(n807), .Z(n809) );
  XOR U7998 ( .A(n1183), .B(n1184), .Z(n807) );
  AND U7999 ( .A(n1185), .B(n1186), .Z(n1183) );
  AND U8000 ( .A(b[29]), .B(a[95]), .Z(n1182) );
  XOR U8001 ( .A(n1187), .B(n812), .Z(n814) );
  XOR U8002 ( .A(n1188), .B(n1189), .Z(n812) );
  AND U8003 ( .A(n1190), .B(n1191), .Z(n1188) );
  AND U8004 ( .A(b[28]), .B(a[96]), .Z(n1187) );
  XOR U8005 ( .A(n1192), .B(n817), .Z(n819) );
  XOR U8006 ( .A(n1193), .B(n1194), .Z(n817) );
  AND U8007 ( .A(n1195), .B(n1196), .Z(n1193) );
  AND U8008 ( .A(b[27]), .B(a[97]), .Z(n1192) );
  XOR U8009 ( .A(n1197), .B(n822), .Z(n824) );
  XOR U8010 ( .A(n1198), .B(n1199), .Z(n822) );
  AND U8011 ( .A(n1200), .B(n1201), .Z(n1198) );
  AND U8012 ( .A(b[26]), .B(a[98]), .Z(n1197) );
  XOR U8013 ( .A(n1202), .B(n1203), .Z(n826) );
  AND U8014 ( .A(n1204), .B(n1205), .Z(n1202) );
  XOR U8015 ( .A(n1206), .B(n831), .Z(n833) );
  XOR U8016 ( .A(n1207), .B(n1208), .Z(n831) );
  AND U8017 ( .A(n1209), .B(n1210), .Z(n1207) );
  AND U8018 ( .A(b[25]), .B(a[99]), .Z(n1206) );
  XOR U8019 ( .A(n1211), .B(n836), .Z(n838) );
  XOR U8020 ( .A(n1212), .B(n1213), .Z(n836) );
  AND U8021 ( .A(n1214), .B(n1215), .Z(n1212) );
  AND U8022 ( .A(b[23]), .B(a[101]), .Z(n1211) );
  XOR U8023 ( .A(n1216), .B(n841), .Z(n843) );
  XOR U8024 ( .A(n1217), .B(n1218), .Z(n841) );
  AND U8025 ( .A(n1219), .B(n1220), .Z(n1217) );
  AND U8026 ( .A(b[22]), .B(a[102]), .Z(n1216) );
  XOR U8027 ( .A(n1221), .B(n846), .Z(n848) );
  XOR U8028 ( .A(n1222), .B(n1223), .Z(n846) );
  AND U8029 ( .A(n1224), .B(n1225), .Z(n1222) );
  AND U8030 ( .A(b[21]), .B(a[103]), .Z(n1221) );
  XOR U8031 ( .A(n1226), .B(n851), .Z(n853) );
  XOR U8032 ( .A(n1227), .B(n1228), .Z(n851) );
  AND U8033 ( .A(n1229), .B(n1230), .Z(n1227) );
  AND U8034 ( .A(b[20]), .B(a[104]), .Z(n1226) );
  XOR U8035 ( .A(n1231), .B(n1232), .Z(n855) );
  AND U8036 ( .A(n1233), .B(n1234), .Z(n1231) );
  XOR U8037 ( .A(n1235), .B(n860), .Z(n862) );
  XOR U8038 ( .A(n1236), .B(n1237), .Z(n860) );
  AND U8039 ( .A(n1238), .B(n1239), .Z(n1236) );
  AND U8040 ( .A(b[19]), .B(a[105]), .Z(n1235) );
  XOR U8041 ( .A(n1240), .B(n865), .Z(n867) );
  XOR U8042 ( .A(n1241), .B(n1242), .Z(n865) );
  AND U8043 ( .A(n1243), .B(n1244), .Z(n1241) );
  AND U8044 ( .A(b[17]), .B(a[107]), .Z(n1240) );
  XOR U8045 ( .A(n1245), .B(n870), .Z(n872) );
  XOR U8046 ( .A(n1246), .B(n1247), .Z(n870) );
  AND U8047 ( .A(n1248), .B(n1249), .Z(n1246) );
  AND U8048 ( .A(b[16]), .B(a[108]), .Z(n1245) );
  XOR U8049 ( .A(n1250), .B(n875), .Z(n877) );
  XOR U8050 ( .A(n1251), .B(n1252), .Z(n875) );
  AND U8051 ( .A(n1253), .B(n1254), .Z(n1251) );
  AND U8052 ( .A(b[15]), .B(a[109]), .Z(n1250) );
  XOR U8053 ( .A(n1255), .B(n880), .Z(n882) );
  XOR U8054 ( .A(n1256), .B(n1257), .Z(n880) );
  AND U8055 ( .A(n1258), .B(n1259), .Z(n1256) );
  AND U8056 ( .A(b[14]), .B(a[110]), .Z(n1255) );
  XOR U8057 ( .A(n1260), .B(n885), .Z(n887) );
  XOR U8058 ( .A(n1261), .B(n1262), .Z(n885) );
  AND U8059 ( .A(n1263), .B(n1264), .Z(n1261) );
  AND U8060 ( .A(b[13]), .B(a[111]), .Z(n1260) );
  XOR U8061 ( .A(n1265), .B(n890), .Z(n892) );
  XOR U8062 ( .A(n1266), .B(n1267), .Z(n890) );
  AND U8063 ( .A(n1268), .B(n1269), .Z(n1266) );
  AND U8064 ( .A(b[12]), .B(a[112]), .Z(n1265) );
  XOR U8065 ( .A(n1270), .B(n895), .Z(n897) );
  XOR U8066 ( .A(n1271), .B(n1272), .Z(n895) );
  AND U8067 ( .A(n1273), .B(n1274), .Z(n1271) );
  AND U8068 ( .A(b[11]), .B(a[113]), .Z(n1270) );
  XOR U8069 ( .A(n1275), .B(n900), .Z(n902) );
  XOR U8070 ( .A(n1276), .B(n1277), .Z(n900) );
  AND U8071 ( .A(n1278), .B(n1279), .Z(n1276) );
  AND U8072 ( .A(b[10]), .B(a[114]), .Z(n1275) );
  XOR U8073 ( .A(n1280), .B(n905), .Z(n907) );
  XOR U8074 ( .A(n1281), .B(n1282), .Z(n905) );
  AND U8075 ( .A(n1283), .B(n1284), .Z(n1281) );
  AND U8076 ( .A(b[9]), .B(a[115]), .Z(n1280) );
  XOR U8077 ( .A(n1285), .B(n910), .Z(n912) );
  XOR U8078 ( .A(n1286), .B(n1287), .Z(n910) );
  AND U8079 ( .A(n1288), .B(n1289), .Z(n1286) );
  AND U8080 ( .A(b[8]), .B(a[116]), .Z(n1285) );
  XOR U8081 ( .A(n1290), .B(n915), .Z(n917) );
  XOR U8082 ( .A(n1291), .B(n1292), .Z(n915) );
  AND U8083 ( .A(n1293), .B(n1294), .Z(n1291) );
  AND U8084 ( .A(b[7]), .B(a[117]), .Z(n1290) );
  XOR U8085 ( .A(n1295), .B(n920), .Z(n922) );
  XOR U8086 ( .A(n1296), .B(n1297), .Z(n920) );
  AND U8087 ( .A(n1298), .B(n1299), .Z(n1296) );
  AND U8088 ( .A(b[6]), .B(a[118]), .Z(n1295) );
  XOR U8089 ( .A(n1300), .B(n925), .Z(n927) );
  XOR U8090 ( .A(n1301), .B(n1302), .Z(n925) );
  AND U8091 ( .A(n1303), .B(n1304), .Z(n1301) );
  AND U8092 ( .A(b[5]), .B(a[119]), .Z(n1300) );
  XOR U8093 ( .A(n1305), .B(n930), .Z(n932) );
  XOR U8094 ( .A(n1306), .B(n1307), .Z(n930) );
  AND U8095 ( .A(n1308), .B(n1309), .Z(n1306) );
  AND U8096 ( .A(b[4]), .B(a[120]), .Z(n1305) );
  XNOR U8097 ( .A(n1310), .B(n1311), .Z(n944) );
  NANDN U8098 ( .A(n1312), .B(n1313), .Z(n1311) );
  XOR U8099 ( .A(n1314), .B(n935), .Z(n937) );
  XNOR U8100 ( .A(n1315), .B(n1316), .Z(n935) );
  AND U8101 ( .A(n1317), .B(n1318), .Z(n1315) );
  AND U8102 ( .A(b[3]), .B(a[121]), .Z(n1314) );
  XOR U8103 ( .A(n1319), .B(n1320), .Z(swire[123]) );
  XOR U8104 ( .A(n954), .B(n1321), .Z(n1320) );
  XNOR U8105 ( .A(n953), .B(n1319), .Z(n1321) );
  NAND U8106 ( .A(a[123]), .B(b[0]), .Z(n953) );
  XNOR U8107 ( .A(n1312), .B(n1313), .Z(n954) );
  XOR U8108 ( .A(n1310), .B(n1322), .Z(n1313) );
  NAND U8109 ( .A(b[1]), .B(a[122]), .Z(n1322) );
  XOR U8110 ( .A(n1318), .B(n1323), .Z(n1312) );
  XOR U8111 ( .A(n1310), .B(n1317), .Z(n1323) );
  XNOR U8112 ( .A(n1324), .B(n1316), .Z(n1317) );
  AND U8113 ( .A(b[2]), .B(a[121]), .Z(n1324) );
  NANDN U8114 ( .A(n1325), .B(n1326), .Z(n1310) );
  XOR U8115 ( .A(n1316), .B(n1308), .Z(n1327) );
  XNOR U8116 ( .A(n1307), .B(n1303), .Z(n1328) );
  XNOR U8117 ( .A(n1302), .B(n1298), .Z(n1329) );
  XNOR U8118 ( .A(n1297), .B(n1293), .Z(n1330) );
  XNOR U8119 ( .A(n1292), .B(n1288), .Z(n1331) );
  XNOR U8120 ( .A(n1287), .B(n1283), .Z(n1332) );
  XNOR U8121 ( .A(n1282), .B(n1278), .Z(n1333) );
  XNOR U8122 ( .A(n1277), .B(n1273), .Z(n1334) );
  XNOR U8123 ( .A(n1272), .B(n1268), .Z(n1335) );
  XNOR U8124 ( .A(n1267), .B(n1263), .Z(n1336) );
  XNOR U8125 ( .A(n1262), .B(n1258), .Z(n1337) );
  XNOR U8126 ( .A(n1257), .B(n1253), .Z(n1338) );
  XNOR U8127 ( .A(n1252), .B(n1248), .Z(n1339) );
  XNOR U8128 ( .A(n1247), .B(n1243), .Z(n1340) );
  XNOR U8129 ( .A(n1234), .B(n1233), .Z(n1341) );
  XOR U8130 ( .A(n1342), .B(n1232), .Z(n1233) );
  AND U8131 ( .A(b[17]), .B(a[106]), .Z(n1342) );
  XNOR U8132 ( .A(n1232), .B(n1238), .Z(n1343) );
  XNOR U8133 ( .A(n1237), .B(n1229), .Z(n1344) );
  XNOR U8134 ( .A(n1228), .B(n1224), .Z(n1345) );
  XNOR U8135 ( .A(n1223), .B(n1219), .Z(n1346) );
  XNOR U8136 ( .A(n1218), .B(n1214), .Z(n1347) );
  XNOR U8137 ( .A(n1205), .B(n1204), .Z(n1348) );
  XOR U8138 ( .A(n1349), .B(n1203), .Z(n1204) );
  AND U8139 ( .A(b[23]), .B(a[100]), .Z(n1349) );
  XNOR U8140 ( .A(n1203), .B(n1209), .Z(n1350) );
  XNOR U8141 ( .A(n1208), .B(n1200), .Z(n1351) );
  XNOR U8142 ( .A(n1199), .B(n1195), .Z(n1352) );
  XNOR U8143 ( .A(n1194), .B(n1190), .Z(n1353) );
  XNOR U8144 ( .A(n1189), .B(n1185), .Z(n1354) );
  XNOR U8145 ( .A(n1176), .B(n1175), .Z(n1355) );
  XOR U8146 ( .A(n1356), .B(n1174), .Z(n1175) );
  AND U8147 ( .A(b[29]), .B(a[94]), .Z(n1356) );
  XNOR U8148 ( .A(n1174), .B(n1180), .Z(n1357) );
  XNOR U8149 ( .A(n1179), .B(n1171), .Z(n1358) );
  XNOR U8150 ( .A(n1170), .B(n1166), .Z(n1359) );
  XNOR U8151 ( .A(n1165), .B(n1161), .Z(n1360) );
  XNOR U8152 ( .A(n1160), .B(n1156), .Z(n1361) );
  XNOR U8153 ( .A(n1147), .B(n1146), .Z(n1362) );
  XOR U8154 ( .A(n1363), .B(n1145), .Z(n1146) );
  AND U8155 ( .A(b[35]), .B(a[88]), .Z(n1363) );
  XNOR U8156 ( .A(n1145), .B(n1151), .Z(n1364) );
  XNOR U8157 ( .A(n1150), .B(n1142), .Z(n1365) );
  XNOR U8158 ( .A(n1141), .B(n1137), .Z(n1366) );
  XNOR U8159 ( .A(n1136), .B(n1132), .Z(n1367) );
  XNOR U8160 ( .A(n1131), .B(n1127), .Z(n1368) );
  XNOR U8161 ( .A(n1118), .B(n1117), .Z(n1369) );
  XOR U8162 ( .A(n1370), .B(n1116), .Z(n1117) );
  AND U8163 ( .A(b[41]), .B(a[82]), .Z(n1370) );
  XNOR U8164 ( .A(n1116), .B(n1122), .Z(n1371) );
  XNOR U8165 ( .A(n1121), .B(n1113), .Z(n1372) );
  XNOR U8166 ( .A(n1112), .B(n1108), .Z(n1373) );
  XNOR U8167 ( .A(n1107), .B(n1103), .Z(n1374) );
  XNOR U8168 ( .A(n1102), .B(n1098), .Z(n1375) );
  XNOR U8169 ( .A(n1089), .B(n1088), .Z(n1376) );
  XOR U8170 ( .A(n1377), .B(n1087), .Z(n1088) );
  AND U8171 ( .A(b[47]), .B(a[76]), .Z(n1377) );
  XNOR U8172 ( .A(n1087), .B(n1093), .Z(n1378) );
  XNOR U8173 ( .A(n1092), .B(n1084), .Z(n1379) );
  XNOR U8174 ( .A(n1083), .B(n1079), .Z(n1380) );
  XNOR U8175 ( .A(n1078), .B(n1074), .Z(n1381) );
  XNOR U8176 ( .A(n1073), .B(n1069), .Z(n1382) );
  XNOR U8177 ( .A(n1060), .B(n1059), .Z(n1383) );
  XOR U8178 ( .A(n1384), .B(n1058), .Z(n1059) );
  AND U8179 ( .A(b[53]), .B(a[70]), .Z(n1384) );
  XNOR U8180 ( .A(n1058), .B(n1064), .Z(n1385) );
  XNOR U8181 ( .A(n1063), .B(n1055), .Z(n1386) );
  XNOR U8182 ( .A(n1054), .B(n1050), .Z(n1387) );
  XNOR U8183 ( .A(n1049), .B(n1045), .Z(n1388) );
  XNOR U8184 ( .A(n1044), .B(n1040), .Z(n1389) );
  XNOR U8185 ( .A(n1039), .B(n1035), .Z(n1390) );
  XOR U8186 ( .A(n1034), .B(n1031), .Z(n1391) );
  XOR U8187 ( .A(n1392), .B(n1393), .Z(n1031) );
  XOR U8188 ( .A(n1029), .B(n1394), .Z(n1393) );
  XOR U8189 ( .A(n1395), .B(n1396), .Z(n1394) );
  XOR U8190 ( .A(n1397), .B(n1398), .Z(n1396) );
  NAND U8191 ( .A(a[61]), .B(b[62]), .Z(n1398) );
  AND U8192 ( .A(a[60]), .B(b[63]), .Z(n1397) );
  XOR U8193 ( .A(n1399), .B(n1395), .Z(n1392) );
  XOR U8194 ( .A(n1400), .B(n1401), .Z(n1395) );
  ANDN U8195 ( .B(n1402), .A(n1403), .Z(n1400) );
  AND U8196 ( .A(b[61]), .B(a[62]), .Z(n1399) );
  XOR U8197 ( .A(n1404), .B(n1029), .Z(n1030) );
  XOR U8198 ( .A(n1405), .B(n1406), .Z(n1029) );
  AND U8199 ( .A(n1407), .B(n1408), .Z(n1405) );
  AND U8200 ( .A(b[60]), .B(a[63]), .Z(n1404) );
  XOR U8201 ( .A(n1409), .B(n1034), .Z(n1036) );
  XOR U8202 ( .A(n1410), .B(n1411), .Z(n1034) );
  AND U8203 ( .A(n1412), .B(n1413), .Z(n1410) );
  AND U8204 ( .A(b[59]), .B(a[64]), .Z(n1409) );
  XOR U8205 ( .A(n1414), .B(n1039), .Z(n1041) );
  XOR U8206 ( .A(n1415), .B(n1416), .Z(n1039) );
  AND U8207 ( .A(n1417), .B(n1418), .Z(n1415) );
  AND U8208 ( .A(b[58]), .B(a[65]), .Z(n1414) );
  XOR U8209 ( .A(n1419), .B(n1044), .Z(n1046) );
  XOR U8210 ( .A(n1420), .B(n1421), .Z(n1044) );
  AND U8211 ( .A(n1422), .B(n1423), .Z(n1420) );
  AND U8212 ( .A(b[57]), .B(a[66]), .Z(n1419) );
  XOR U8213 ( .A(n1424), .B(n1049), .Z(n1051) );
  XOR U8214 ( .A(n1425), .B(n1426), .Z(n1049) );
  AND U8215 ( .A(n1427), .B(n1428), .Z(n1425) );
  AND U8216 ( .A(b[56]), .B(a[67]), .Z(n1424) );
  XOR U8217 ( .A(n1429), .B(n1054), .Z(n1056) );
  XOR U8218 ( .A(n1430), .B(n1431), .Z(n1054) );
  AND U8219 ( .A(n1432), .B(n1433), .Z(n1430) );
  AND U8220 ( .A(b[55]), .B(a[68]), .Z(n1429) );
  XOR U8221 ( .A(n1434), .B(n1435), .Z(n1058) );
  AND U8222 ( .A(n1436), .B(n1437), .Z(n1434) );
  XOR U8223 ( .A(n1438), .B(n1063), .Z(n1065) );
  XOR U8224 ( .A(n1439), .B(n1440), .Z(n1063) );
  AND U8225 ( .A(n1441), .B(n1442), .Z(n1439) );
  AND U8226 ( .A(b[54]), .B(a[69]), .Z(n1438) );
  XOR U8227 ( .A(n1443), .B(n1068), .Z(n1070) );
  XOR U8228 ( .A(n1444), .B(n1445), .Z(n1068) );
  AND U8229 ( .A(n1446), .B(n1447), .Z(n1444) );
  AND U8230 ( .A(b[52]), .B(a[71]), .Z(n1443) );
  XOR U8231 ( .A(n1448), .B(n1073), .Z(n1075) );
  XOR U8232 ( .A(n1449), .B(n1450), .Z(n1073) );
  AND U8233 ( .A(n1451), .B(n1452), .Z(n1449) );
  AND U8234 ( .A(b[51]), .B(a[72]), .Z(n1448) );
  XOR U8235 ( .A(n1453), .B(n1078), .Z(n1080) );
  XOR U8236 ( .A(n1454), .B(n1455), .Z(n1078) );
  AND U8237 ( .A(n1456), .B(n1457), .Z(n1454) );
  AND U8238 ( .A(b[50]), .B(a[73]), .Z(n1453) );
  XOR U8239 ( .A(n1458), .B(n1083), .Z(n1085) );
  XOR U8240 ( .A(n1459), .B(n1460), .Z(n1083) );
  AND U8241 ( .A(n1461), .B(n1462), .Z(n1459) );
  AND U8242 ( .A(b[49]), .B(a[74]), .Z(n1458) );
  XOR U8243 ( .A(n1463), .B(n1464), .Z(n1087) );
  AND U8244 ( .A(n1465), .B(n1466), .Z(n1463) );
  XOR U8245 ( .A(n1467), .B(n1092), .Z(n1094) );
  XOR U8246 ( .A(n1468), .B(n1469), .Z(n1092) );
  AND U8247 ( .A(n1470), .B(n1471), .Z(n1468) );
  AND U8248 ( .A(b[48]), .B(a[75]), .Z(n1467) );
  XOR U8249 ( .A(n1472), .B(n1097), .Z(n1099) );
  XOR U8250 ( .A(n1473), .B(n1474), .Z(n1097) );
  AND U8251 ( .A(n1475), .B(n1476), .Z(n1473) );
  AND U8252 ( .A(b[46]), .B(a[77]), .Z(n1472) );
  XOR U8253 ( .A(n1477), .B(n1102), .Z(n1104) );
  XOR U8254 ( .A(n1478), .B(n1479), .Z(n1102) );
  AND U8255 ( .A(n1480), .B(n1481), .Z(n1478) );
  AND U8256 ( .A(b[45]), .B(a[78]), .Z(n1477) );
  XOR U8257 ( .A(n1482), .B(n1107), .Z(n1109) );
  XOR U8258 ( .A(n1483), .B(n1484), .Z(n1107) );
  AND U8259 ( .A(n1485), .B(n1486), .Z(n1483) );
  AND U8260 ( .A(b[44]), .B(a[79]), .Z(n1482) );
  XOR U8261 ( .A(n1487), .B(n1112), .Z(n1114) );
  XOR U8262 ( .A(n1488), .B(n1489), .Z(n1112) );
  AND U8263 ( .A(n1490), .B(n1491), .Z(n1488) );
  AND U8264 ( .A(b[43]), .B(a[80]), .Z(n1487) );
  XOR U8265 ( .A(n1492), .B(n1493), .Z(n1116) );
  AND U8266 ( .A(n1494), .B(n1495), .Z(n1492) );
  XOR U8267 ( .A(n1496), .B(n1121), .Z(n1123) );
  XOR U8268 ( .A(n1497), .B(n1498), .Z(n1121) );
  AND U8269 ( .A(n1499), .B(n1500), .Z(n1497) );
  AND U8270 ( .A(b[42]), .B(a[81]), .Z(n1496) );
  XOR U8271 ( .A(n1501), .B(n1126), .Z(n1128) );
  XOR U8272 ( .A(n1502), .B(n1503), .Z(n1126) );
  AND U8273 ( .A(n1504), .B(n1505), .Z(n1502) );
  AND U8274 ( .A(b[40]), .B(a[83]), .Z(n1501) );
  XOR U8275 ( .A(n1506), .B(n1131), .Z(n1133) );
  XOR U8276 ( .A(n1507), .B(n1508), .Z(n1131) );
  AND U8277 ( .A(n1509), .B(n1510), .Z(n1507) );
  AND U8278 ( .A(b[39]), .B(a[84]), .Z(n1506) );
  XOR U8279 ( .A(n1511), .B(n1136), .Z(n1138) );
  XOR U8280 ( .A(n1512), .B(n1513), .Z(n1136) );
  AND U8281 ( .A(n1514), .B(n1515), .Z(n1512) );
  AND U8282 ( .A(b[38]), .B(a[85]), .Z(n1511) );
  XOR U8283 ( .A(n1516), .B(n1141), .Z(n1143) );
  XOR U8284 ( .A(n1517), .B(n1518), .Z(n1141) );
  AND U8285 ( .A(n1519), .B(n1520), .Z(n1517) );
  AND U8286 ( .A(b[37]), .B(a[86]), .Z(n1516) );
  XOR U8287 ( .A(n1521), .B(n1522), .Z(n1145) );
  AND U8288 ( .A(n1523), .B(n1524), .Z(n1521) );
  XOR U8289 ( .A(n1525), .B(n1150), .Z(n1152) );
  XOR U8290 ( .A(n1526), .B(n1527), .Z(n1150) );
  AND U8291 ( .A(n1528), .B(n1529), .Z(n1526) );
  AND U8292 ( .A(b[36]), .B(a[87]), .Z(n1525) );
  XOR U8293 ( .A(n1530), .B(n1155), .Z(n1157) );
  XOR U8294 ( .A(n1531), .B(n1532), .Z(n1155) );
  AND U8295 ( .A(n1533), .B(n1534), .Z(n1531) );
  AND U8296 ( .A(b[34]), .B(a[89]), .Z(n1530) );
  XOR U8297 ( .A(n1535), .B(n1160), .Z(n1162) );
  XOR U8298 ( .A(n1536), .B(n1537), .Z(n1160) );
  AND U8299 ( .A(n1538), .B(n1539), .Z(n1536) );
  AND U8300 ( .A(b[33]), .B(a[90]), .Z(n1535) );
  XOR U8301 ( .A(n1540), .B(n1165), .Z(n1167) );
  XOR U8302 ( .A(n1541), .B(n1542), .Z(n1165) );
  AND U8303 ( .A(n1543), .B(n1544), .Z(n1541) );
  AND U8304 ( .A(b[32]), .B(a[91]), .Z(n1540) );
  XOR U8305 ( .A(n1545), .B(n1170), .Z(n1172) );
  XOR U8306 ( .A(n1546), .B(n1547), .Z(n1170) );
  AND U8307 ( .A(n1548), .B(n1549), .Z(n1546) );
  AND U8308 ( .A(b[31]), .B(a[92]), .Z(n1545) );
  XOR U8309 ( .A(n1550), .B(n1551), .Z(n1174) );
  AND U8310 ( .A(n1552), .B(n1553), .Z(n1550) );
  XOR U8311 ( .A(n1554), .B(n1179), .Z(n1181) );
  XOR U8312 ( .A(n1555), .B(n1556), .Z(n1179) );
  AND U8313 ( .A(n1557), .B(n1558), .Z(n1555) );
  AND U8314 ( .A(b[30]), .B(a[93]), .Z(n1554) );
  XOR U8315 ( .A(n1559), .B(n1184), .Z(n1186) );
  XOR U8316 ( .A(n1560), .B(n1561), .Z(n1184) );
  AND U8317 ( .A(n1562), .B(n1563), .Z(n1560) );
  AND U8318 ( .A(b[28]), .B(a[95]), .Z(n1559) );
  XOR U8319 ( .A(n1564), .B(n1189), .Z(n1191) );
  XOR U8320 ( .A(n1565), .B(n1566), .Z(n1189) );
  AND U8321 ( .A(n1567), .B(n1568), .Z(n1565) );
  AND U8322 ( .A(b[27]), .B(a[96]), .Z(n1564) );
  XOR U8323 ( .A(n1569), .B(n1194), .Z(n1196) );
  XOR U8324 ( .A(n1570), .B(n1571), .Z(n1194) );
  AND U8325 ( .A(n1572), .B(n1573), .Z(n1570) );
  AND U8326 ( .A(b[26]), .B(a[97]), .Z(n1569) );
  XOR U8327 ( .A(n1574), .B(n1199), .Z(n1201) );
  XOR U8328 ( .A(n1575), .B(n1576), .Z(n1199) );
  AND U8329 ( .A(n1577), .B(n1578), .Z(n1575) );
  AND U8330 ( .A(b[25]), .B(a[98]), .Z(n1574) );
  XOR U8331 ( .A(n1579), .B(n1580), .Z(n1203) );
  AND U8332 ( .A(n1581), .B(n1582), .Z(n1579) );
  XOR U8333 ( .A(n1583), .B(n1208), .Z(n1210) );
  XOR U8334 ( .A(n1584), .B(n1585), .Z(n1208) );
  AND U8335 ( .A(n1586), .B(n1587), .Z(n1584) );
  AND U8336 ( .A(b[24]), .B(a[99]), .Z(n1583) );
  XOR U8337 ( .A(n1588), .B(n1213), .Z(n1215) );
  XOR U8338 ( .A(n1589), .B(n1590), .Z(n1213) );
  AND U8339 ( .A(n1591), .B(n1592), .Z(n1589) );
  AND U8340 ( .A(b[22]), .B(a[101]), .Z(n1588) );
  XOR U8341 ( .A(n1593), .B(n1218), .Z(n1220) );
  XOR U8342 ( .A(n1594), .B(n1595), .Z(n1218) );
  AND U8343 ( .A(n1596), .B(n1597), .Z(n1594) );
  AND U8344 ( .A(b[21]), .B(a[102]), .Z(n1593) );
  XOR U8345 ( .A(n1598), .B(n1223), .Z(n1225) );
  XOR U8346 ( .A(n1599), .B(n1600), .Z(n1223) );
  AND U8347 ( .A(n1601), .B(n1602), .Z(n1599) );
  AND U8348 ( .A(b[20]), .B(a[103]), .Z(n1598) );
  XOR U8349 ( .A(n1603), .B(n1228), .Z(n1230) );
  XOR U8350 ( .A(n1604), .B(n1605), .Z(n1228) );
  AND U8351 ( .A(n1606), .B(n1607), .Z(n1604) );
  AND U8352 ( .A(b[19]), .B(a[104]), .Z(n1603) );
  XOR U8353 ( .A(n1608), .B(n1609), .Z(n1232) );
  AND U8354 ( .A(n1610), .B(n1611), .Z(n1608) );
  XOR U8355 ( .A(n1612), .B(n1237), .Z(n1239) );
  XOR U8356 ( .A(n1613), .B(n1614), .Z(n1237) );
  AND U8357 ( .A(n1615), .B(n1616), .Z(n1613) );
  AND U8358 ( .A(b[18]), .B(a[105]), .Z(n1612) );
  XOR U8359 ( .A(n1617), .B(n1242), .Z(n1244) );
  XOR U8360 ( .A(n1618), .B(n1619), .Z(n1242) );
  AND U8361 ( .A(n1620), .B(n1621), .Z(n1618) );
  AND U8362 ( .A(b[16]), .B(a[107]), .Z(n1617) );
  XOR U8363 ( .A(n1622), .B(n1247), .Z(n1249) );
  XOR U8364 ( .A(n1623), .B(n1624), .Z(n1247) );
  AND U8365 ( .A(n1625), .B(n1626), .Z(n1623) );
  AND U8366 ( .A(b[15]), .B(a[108]), .Z(n1622) );
  XOR U8367 ( .A(n1627), .B(n1252), .Z(n1254) );
  XOR U8368 ( .A(n1628), .B(n1629), .Z(n1252) );
  AND U8369 ( .A(n1630), .B(n1631), .Z(n1628) );
  AND U8370 ( .A(b[14]), .B(a[109]), .Z(n1627) );
  XOR U8371 ( .A(n1632), .B(n1257), .Z(n1259) );
  XOR U8372 ( .A(n1633), .B(n1634), .Z(n1257) );
  AND U8373 ( .A(n1635), .B(n1636), .Z(n1633) );
  AND U8374 ( .A(b[13]), .B(a[110]), .Z(n1632) );
  XOR U8375 ( .A(n1637), .B(n1262), .Z(n1264) );
  XOR U8376 ( .A(n1638), .B(n1639), .Z(n1262) );
  AND U8377 ( .A(n1640), .B(n1641), .Z(n1638) );
  AND U8378 ( .A(b[12]), .B(a[111]), .Z(n1637) );
  XOR U8379 ( .A(n1642), .B(n1267), .Z(n1269) );
  XOR U8380 ( .A(n1643), .B(n1644), .Z(n1267) );
  AND U8381 ( .A(n1645), .B(n1646), .Z(n1643) );
  AND U8382 ( .A(b[11]), .B(a[112]), .Z(n1642) );
  XOR U8383 ( .A(n1647), .B(n1272), .Z(n1274) );
  XOR U8384 ( .A(n1648), .B(n1649), .Z(n1272) );
  AND U8385 ( .A(n1650), .B(n1651), .Z(n1648) );
  AND U8386 ( .A(b[10]), .B(a[113]), .Z(n1647) );
  XOR U8387 ( .A(n1652), .B(n1277), .Z(n1279) );
  XOR U8388 ( .A(n1653), .B(n1654), .Z(n1277) );
  AND U8389 ( .A(n1655), .B(n1656), .Z(n1653) );
  AND U8390 ( .A(b[9]), .B(a[114]), .Z(n1652) );
  XOR U8391 ( .A(n1657), .B(n1282), .Z(n1284) );
  XOR U8392 ( .A(n1658), .B(n1659), .Z(n1282) );
  AND U8393 ( .A(n1660), .B(n1661), .Z(n1658) );
  AND U8394 ( .A(b[8]), .B(a[115]), .Z(n1657) );
  XOR U8395 ( .A(n1662), .B(n1287), .Z(n1289) );
  XOR U8396 ( .A(n1663), .B(n1664), .Z(n1287) );
  AND U8397 ( .A(n1665), .B(n1666), .Z(n1663) );
  AND U8398 ( .A(b[7]), .B(a[116]), .Z(n1662) );
  XOR U8399 ( .A(n1667), .B(n1292), .Z(n1294) );
  XOR U8400 ( .A(n1668), .B(n1669), .Z(n1292) );
  AND U8401 ( .A(n1670), .B(n1671), .Z(n1668) );
  AND U8402 ( .A(b[6]), .B(a[117]), .Z(n1667) );
  XOR U8403 ( .A(n1672), .B(n1297), .Z(n1299) );
  XOR U8404 ( .A(n1673), .B(n1674), .Z(n1297) );
  AND U8405 ( .A(n1675), .B(n1676), .Z(n1673) );
  AND U8406 ( .A(b[5]), .B(a[118]), .Z(n1672) );
  XOR U8407 ( .A(n1677), .B(n1302), .Z(n1304) );
  XOR U8408 ( .A(n1678), .B(n1679), .Z(n1302) );
  AND U8409 ( .A(n1680), .B(n1681), .Z(n1678) );
  AND U8410 ( .A(b[4]), .B(a[119]), .Z(n1677) );
  XNOR U8411 ( .A(n1682), .B(n1683), .Z(n1316) );
  NANDN U8412 ( .A(n1684), .B(n1685), .Z(n1683) );
  XOR U8413 ( .A(n1686), .B(n1307), .Z(n1309) );
  XNOR U8414 ( .A(n1687), .B(n1688), .Z(n1307) );
  AND U8415 ( .A(n1689), .B(n1690), .Z(n1687) );
  AND U8416 ( .A(b[3]), .B(a[120]), .Z(n1686) );
  XOR U8417 ( .A(n1691), .B(n1692), .Z(swire[122]) );
  XOR U8418 ( .A(n1326), .B(n1693), .Z(n1692) );
  XNOR U8419 ( .A(n1325), .B(n1691), .Z(n1693) );
  NAND U8420 ( .A(a[122]), .B(b[0]), .Z(n1325) );
  XNOR U8421 ( .A(n1684), .B(n1685), .Z(n1326) );
  XOR U8422 ( .A(n1682), .B(n1694), .Z(n1685) );
  NAND U8423 ( .A(b[1]), .B(a[121]), .Z(n1694) );
  XOR U8424 ( .A(n1690), .B(n1695), .Z(n1684) );
  XOR U8425 ( .A(n1682), .B(n1689), .Z(n1695) );
  XNOR U8426 ( .A(n1696), .B(n1688), .Z(n1689) );
  AND U8427 ( .A(b[2]), .B(a[120]), .Z(n1696) );
  NANDN U8428 ( .A(n1697), .B(n1698), .Z(n1682) );
  XOR U8429 ( .A(n1688), .B(n1680), .Z(n1699) );
  XNOR U8430 ( .A(n1679), .B(n1675), .Z(n1700) );
  XNOR U8431 ( .A(n1674), .B(n1670), .Z(n1701) );
  XNOR U8432 ( .A(n1669), .B(n1665), .Z(n1702) );
  XNOR U8433 ( .A(n1664), .B(n1660), .Z(n1703) );
  XNOR U8434 ( .A(n1659), .B(n1655), .Z(n1704) );
  XNOR U8435 ( .A(n1654), .B(n1650), .Z(n1705) );
  XNOR U8436 ( .A(n1649), .B(n1645), .Z(n1706) );
  XNOR U8437 ( .A(n1644), .B(n1640), .Z(n1707) );
  XNOR U8438 ( .A(n1639), .B(n1635), .Z(n1708) );
  XNOR U8439 ( .A(n1634), .B(n1630), .Z(n1709) );
  XNOR U8440 ( .A(n1629), .B(n1625), .Z(n1710) );
  XNOR U8441 ( .A(n1624), .B(n1620), .Z(n1711) );
  XNOR U8442 ( .A(n1611), .B(n1610), .Z(n1712) );
  XOR U8443 ( .A(n1713), .B(n1609), .Z(n1610) );
  AND U8444 ( .A(b[16]), .B(a[106]), .Z(n1713) );
  XNOR U8445 ( .A(n1609), .B(n1615), .Z(n1714) );
  XNOR U8446 ( .A(n1614), .B(n1606), .Z(n1715) );
  XNOR U8447 ( .A(n1605), .B(n1601), .Z(n1716) );
  XNOR U8448 ( .A(n1600), .B(n1596), .Z(n1717) );
  XNOR U8449 ( .A(n1595), .B(n1591), .Z(n1718) );
  XNOR U8450 ( .A(n1582), .B(n1581), .Z(n1719) );
  XOR U8451 ( .A(n1720), .B(n1580), .Z(n1581) );
  AND U8452 ( .A(b[22]), .B(a[100]), .Z(n1720) );
  XNOR U8453 ( .A(n1580), .B(n1586), .Z(n1721) );
  XNOR U8454 ( .A(n1585), .B(n1577), .Z(n1722) );
  XNOR U8455 ( .A(n1576), .B(n1572), .Z(n1723) );
  XNOR U8456 ( .A(n1571), .B(n1567), .Z(n1724) );
  XNOR U8457 ( .A(n1566), .B(n1562), .Z(n1725) );
  XNOR U8458 ( .A(n1553), .B(n1552), .Z(n1726) );
  XOR U8459 ( .A(n1727), .B(n1551), .Z(n1552) );
  AND U8460 ( .A(b[28]), .B(a[94]), .Z(n1727) );
  XNOR U8461 ( .A(n1551), .B(n1557), .Z(n1728) );
  XNOR U8462 ( .A(n1556), .B(n1548), .Z(n1729) );
  XNOR U8463 ( .A(n1547), .B(n1543), .Z(n1730) );
  XNOR U8464 ( .A(n1542), .B(n1538), .Z(n1731) );
  XNOR U8465 ( .A(n1537), .B(n1533), .Z(n1732) );
  XNOR U8466 ( .A(n1524), .B(n1523), .Z(n1733) );
  XOR U8467 ( .A(n1734), .B(n1522), .Z(n1523) );
  AND U8468 ( .A(b[34]), .B(a[88]), .Z(n1734) );
  XNOR U8469 ( .A(n1522), .B(n1528), .Z(n1735) );
  XNOR U8470 ( .A(n1527), .B(n1519), .Z(n1736) );
  XNOR U8471 ( .A(n1518), .B(n1514), .Z(n1737) );
  XNOR U8472 ( .A(n1513), .B(n1509), .Z(n1738) );
  XNOR U8473 ( .A(n1508), .B(n1504), .Z(n1739) );
  XNOR U8474 ( .A(n1495), .B(n1494), .Z(n1740) );
  XOR U8475 ( .A(n1741), .B(n1493), .Z(n1494) );
  AND U8476 ( .A(b[40]), .B(a[82]), .Z(n1741) );
  XNOR U8477 ( .A(n1493), .B(n1499), .Z(n1742) );
  XNOR U8478 ( .A(n1498), .B(n1490), .Z(n1743) );
  XNOR U8479 ( .A(n1489), .B(n1485), .Z(n1744) );
  XNOR U8480 ( .A(n1484), .B(n1480), .Z(n1745) );
  XNOR U8481 ( .A(n1479), .B(n1475), .Z(n1746) );
  XNOR U8482 ( .A(n1466), .B(n1465), .Z(n1747) );
  XOR U8483 ( .A(n1748), .B(n1464), .Z(n1465) );
  AND U8484 ( .A(b[46]), .B(a[76]), .Z(n1748) );
  XNOR U8485 ( .A(n1464), .B(n1470), .Z(n1749) );
  XNOR U8486 ( .A(n1469), .B(n1461), .Z(n1750) );
  XNOR U8487 ( .A(n1460), .B(n1456), .Z(n1751) );
  XNOR U8488 ( .A(n1455), .B(n1451), .Z(n1752) );
  XNOR U8489 ( .A(n1450), .B(n1446), .Z(n1753) );
  XNOR U8490 ( .A(n1437), .B(n1436), .Z(n1754) );
  XOR U8491 ( .A(n1755), .B(n1435), .Z(n1436) );
  AND U8492 ( .A(b[52]), .B(a[70]), .Z(n1755) );
  XNOR U8493 ( .A(n1435), .B(n1441), .Z(n1756) );
  XNOR U8494 ( .A(n1440), .B(n1432), .Z(n1757) );
  XNOR U8495 ( .A(n1431), .B(n1427), .Z(n1758) );
  XNOR U8496 ( .A(n1426), .B(n1422), .Z(n1759) );
  XNOR U8497 ( .A(n1421), .B(n1417), .Z(n1760) );
  XNOR U8498 ( .A(n1416), .B(n1412), .Z(n1761) );
  XNOR U8499 ( .A(n1411), .B(n1407), .Z(n1762) );
  XOR U8500 ( .A(n1406), .B(n1403), .Z(n1763) );
  XOR U8501 ( .A(n1764), .B(n1765), .Z(n1403) );
  XOR U8502 ( .A(n1401), .B(n1766), .Z(n1765) );
  XOR U8503 ( .A(n1767), .B(n1768), .Z(n1766) );
  XOR U8504 ( .A(n1769), .B(n1770), .Z(n1768) );
  NAND U8505 ( .A(a[60]), .B(b[62]), .Z(n1770) );
  AND U8506 ( .A(a[59]), .B(b[63]), .Z(n1769) );
  XOR U8507 ( .A(n1771), .B(n1767), .Z(n1764) );
  XOR U8508 ( .A(n1772), .B(n1773), .Z(n1767) );
  ANDN U8509 ( .B(n1774), .A(n1775), .Z(n1772) );
  AND U8510 ( .A(a[61]), .B(b[61]), .Z(n1771) );
  XOR U8511 ( .A(n1776), .B(n1401), .Z(n1402) );
  XOR U8512 ( .A(n1777), .B(n1778), .Z(n1401) );
  AND U8513 ( .A(n1779), .B(n1780), .Z(n1777) );
  AND U8514 ( .A(b[60]), .B(a[62]), .Z(n1776) );
  XOR U8515 ( .A(n1781), .B(n1406), .Z(n1408) );
  XOR U8516 ( .A(n1782), .B(n1783), .Z(n1406) );
  AND U8517 ( .A(n1784), .B(n1785), .Z(n1782) );
  AND U8518 ( .A(b[59]), .B(a[63]), .Z(n1781) );
  XOR U8519 ( .A(n1786), .B(n1411), .Z(n1413) );
  XOR U8520 ( .A(n1787), .B(n1788), .Z(n1411) );
  AND U8521 ( .A(n1789), .B(n1790), .Z(n1787) );
  AND U8522 ( .A(b[58]), .B(a[64]), .Z(n1786) );
  XOR U8523 ( .A(n1791), .B(n1416), .Z(n1418) );
  XOR U8524 ( .A(n1792), .B(n1793), .Z(n1416) );
  AND U8525 ( .A(n1794), .B(n1795), .Z(n1792) );
  AND U8526 ( .A(b[57]), .B(a[65]), .Z(n1791) );
  XOR U8527 ( .A(n1796), .B(n1421), .Z(n1423) );
  XOR U8528 ( .A(n1797), .B(n1798), .Z(n1421) );
  AND U8529 ( .A(n1799), .B(n1800), .Z(n1797) );
  AND U8530 ( .A(b[56]), .B(a[66]), .Z(n1796) );
  XOR U8531 ( .A(n1801), .B(n1426), .Z(n1428) );
  XOR U8532 ( .A(n1802), .B(n1803), .Z(n1426) );
  AND U8533 ( .A(n1804), .B(n1805), .Z(n1802) );
  AND U8534 ( .A(b[55]), .B(a[67]), .Z(n1801) );
  XOR U8535 ( .A(n1806), .B(n1431), .Z(n1433) );
  XOR U8536 ( .A(n1807), .B(n1808), .Z(n1431) );
  AND U8537 ( .A(n1809), .B(n1810), .Z(n1807) );
  AND U8538 ( .A(b[54]), .B(a[68]), .Z(n1806) );
  XOR U8539 ( .A(n1811), .B(n1812), .Z(n1435) );
  AND U8540 ( .A(n1813), .B(n1814), .Z(n1811) );
  XOR U8541 ( .A(n1815), .B(n1440), .Z(n1442) );
  XOR U8542 ( .A(n1816), .B(n1817), .Z(n1440) );
  AND U8543 ( .A(n1818), .B(n1819), .Z(n1816) );
  AND U8544 ( .A(b[53]), .B(a[69]), .Z(n1815) );
  XOR U8545 ( .A(n1820), .B(n1445), .Z(n1447) );
  XOR U8546 ( .A(n1821), .B(n1822), .Z(n1445) );
  AND U8547 ( .A(n1823), .B(n1824), .Z(n1821) );
  AND U8548 ( .A(b[51]), .B(a[71]), .Z(n1820) );
  XOR U8549 ( .A(n1825), .B(n1450), .Z(n1452) );
  XOR U8550 ( .A(n1826), .B(n1827), .Z(n1450) );
  AND U8551 ( .A(n1828), .B(n1829), .Z(n1826) );
  AND U8552 ( .A(b[50]), .B(a[72]), .Z(n1825) );
  XOR U8553 ( .A(n1830), .B(n1455), .Z(n1457) );
  XOR U8554 ( .A(n1831), .B(n1832), .Z(n1455) );
  AND U8555 ( .A(n1833), .B(n1834), .Z(n1831) );
  AND U8556 ( .A(b[49]), .B(a[73]), .Z(n1830) );
  XOR U8557 ( .A(n1835), .B(n1460), .Z(n1462) );
  XOR U8558 ( .A(n1836), .B(n1837), .Z(n1460) );
  AND U8559 ( .A(n1838), .B(n1839), .Z(n1836) );
  AND U8560 ( .A(b[48]), .B(a[74]), .Z(n1835) );
  XOR U8561 ( .A(n1840), .B(n1841), .Z(n1464) );
  AND U8562 ( .A(n1842), .B(n1843), .Z(n1840) );
  XOR U8563 ( .A(n1844), .B(n1469), .Z(n1471) );
  XOR U8564 ( .A(n1845), .B(n1846), .Z(n1469) );
  AND U8565 ( .A(n1847), .B(n1848), .Z(n1845) );
  AND U8566 ( .A(b[47]), .B(a[75]), .Z(n1844) );
  XOR U8567 ( .A(n1849), .B(n1474), .Z(n1476) );
  XOR U8568 ( .A(n1850), .B(n1851), .Z(n1474) );
  AND U8569 ( .A(n1852), .B(n1853), .Z(n1850) );
  AND U8570 ( .A(b[45]), .B(a[77]), .Z(n1849) );
  XOR U8571 ( .A(n1854), .B(n1479), .Z(n1481) );
  XOR U8572 ( .A(n1855), .B(n1856), .Z(n1479) );
  AND U8573 ( .A(n1857), .B(n1858), .Z(n1855) );
  AND U8574 ( .A(b[44]), .B(a[78]), .Z(n1854) );
  XOR U8575 ( .A(n1859), .B(n1484), .Z(n1486) );
  XOR U8576 ( .A(n1860), .B(n1861), .Z(n1484) );
  AND U8577 ( .A(n1862), .B(n1863), .Z(n1860) );
  AND U8578 ( .A(b[43]), .B(a[79]), .Z(n1859) );
  XOR U8579 ( .A(n1864), .B(n1489), .Z(n1491) );
  XOR U8580 ( .A(n1865), .B(n1866), .Z(n1489) );
  AND U8581 ( .A(n1867), .B(n1868), .Z(n1865) );
  AND U8582 ( .A(b[42]), .B(a[80]), .Z(n1864) );
  XOR U8583 ( .A(n1869), .B(n1870), .Z(n1493) );
  AND U8584 ( .A(n1871), .B(n1872), .Z(n1869) );
  XOR U8585 ( .A(n1873), .B(n1498), .Z(n1500) );
  XOR U8586 ( .A(n1874), .B(n1875), .Z(n1498) );
  AND U8587 ( .A(n1876), .B(n1877), .Z(n1874) );
  AND U8588 ( .A(b[41]), .B(a[81]), .Z(n1873) );
  XOR U8589 ( .A(n1878), .B(n1503), .Z(n1505) );
  XOR U8590 ( .A(n1879), .B(n1880), .Z(n1503) );
  AND U8591 ( .A(n1881), .B(n1882), .Z(n1879) );
  AND U8592 ( .A(b[39]), .B(a[83]), .Z(n1878) );
  XOR U8593 ( .A(n1883), .B(n1508), .Z(n1510) );
  XOR U8594 ( .A(n1884), .B(n1885), .Z(n1508) );
  AND U8595 ( .A(n1886), .B(n1887), .Z(n1884) );
  AND U8596 ( .A(b[38]), .B(a[84]), .Z(n1883) );
  XOR U8597 ( .A(n1888), .B(n1513), .Z(n1515) );
  XOR U8598 ( .A(n1889), .B(n1890), .Z(n1513) );
  AND U8599 ( .A(n1891), .B(n1892), .Z(n1889) );
  AND U8600 ( .A(b[37]), .B(a[85]), .Z(n1888) );
  XOR U8601 ( .A(n1893), .B(n1518), .Z(n1520) );
  XOR U8602 ( .A(n1894), .B(n1895), .Z(n1518) );
  AND U8603 ( .A(n1896), .B(n1897), .Z(n1894) );
  AND U8604 ( .A(b[36]), .B(a[86]), .Z(n1893) );
  XOR U8605 ( .A(n1898), .B(n1899), .Z(n1522) );
  AND U8606 ( .A(n1900), .B(n1901), .Z(n1898) );
  XOR U8607 ( .A(n1902), .B(n1527), .Z(n1529) );
  XOR U8608 ( .A(n1903), .B(n1904), .Z(n1527) );
  AND U8609 ( .A(n1905), .B(n1906), .Z(n1903) );
  AND U8610 ( .A(b[35]), .B(a[87]), .Z(n1902) );
  XOR U8611 ( .A(n1907), .B(n1532), .Z(n1534) );
  XOR U8612 ( .A(n1908), .B(n1909), .Z(n1532) );
  AND U8613 ( .A(n1910), .B(n1911), .Z(n1908) );
  AND U8614 ( .A(b[33]), .B(a[89]), .Z(n1907) );
  XOR U8615 ( .A(n1912), .B(n1537), .Z(n1539) );
  XOR U8616 ( .A(n1913), .B(n1914), .Z(n1537) );
  AND U8617 ( .A(n1915), .B(n1916), .Z(n1913) );
  AND U8618 ( .A(b[32]), .B(a[90]), .Z(n1912) );
  XOR U8619 ( .A(n1917), .B(n1542), .Z(n1544) );
  XOR U8620 ( .A(n1918), .B(n1919), .Z(n1542) );
  AND U8621 ( .A(n1920), .B(n1921), .Z(n1918) );
  AND U8622 ( .A(b[31]), .B(a[91]), .Z(n1917) );
  XOR U8623 ( .A(n1922), .B(n1547), .Z(n1549) );
  XOR U8624 ( .A(n1923), .B(n1924), .Z(n1547) );
  AND U8625 ( .A(n1925), .B(n1926), .Z(n1923) );
  AND U8626 ( .A(b[30]), .B(a[92]), .Z(n1922) );
  XOR U8627 ( .A(n1927), .B(n1928), .Z(n1551) );
  AND U8628 ( .A(n1929), .B(n1930), .Z(n1927) );
  XOR U8629 ( .A(n1931), .B(n1556), .Z(n1558) );
  XOR U8630 ( .A(n1932), .B(n1933), .Z(n1556) );
  AND U8631 ( .A(n1934), .B(n1935), .Z(n1932) );
  AND U8632 ( .A(b[29]), .B(a[93]), .Z(n1931) );
  XOR U8633 ( .A(n1936), .B(n1561), .Z(n1563) );
  XOR U8634 ( .A(n1937), .B(n1938), .Z(n1561) );
  AND U8635 ( .A(n1939), .B(n1940), .Z(n1937) );
  AND U8636 ( .A(b[27]), .B(a[95]), .Z(n1936) );
  XOR U8637 ( .A(n1941), .B(n1566), .Z(n1568) );
  XOR U8638 ( .A(n1942), .B(n1943), .Z(n1566) );
  AND U8639 ( .A(n1944), .B(n1945), .Z(n1942) );
  AND U8640 ( .A(b[26]), .B(a[96]), .Z(n1941) );
  XOR U8641 ( .A(n1946), .B(n1571), .Z(n1573) );
  XOR U8642 ( .A(n1947), .B(n1948), .Z(n1571) );
  AND U8643 ( .A(n1949), .B(n1950), .Z(n1947) );
  AND U8644 ( .A(b[25]), .B(a[97]), .Z(n1946) );
  XOR U8645 ( .A(n1951), .B(n1576), .Z(n1578) );
  XOR U8646 ( .A(n1952), .B(n1953), .Z(n1576) );
  AND U8647 ( .A(n1954), .B(n1955), .Z(n1952) );
  AND U8648 ( .A(b[24]), .B(a[98]), .Z(n1951) );
  XOR U8649 ( .A(n1956), .B(n1957), .Z(n1580) );
  AND U8650 ( .A(n1958), .B(n1959), .Z(n1956) );
  XOR U8651 ( .A(n1960), .B(n1585), .Z(n1587) );
  XOR U8652 ( .A(n1961), .B(n1962), .Z(n1585) );
  AND U8653 ( .A(n1963), .B(n1964), .Z(n1961) );
  AND U8654 ( .A(b[23]), .B(a[99]), .Z(n1960) );
  XOR U8655 ( .A(n1965), .B(n1590), .Z(n1592) );
  XOR U8656 ( .A(n1966), .B(n1967), .Z(n1590) );
  AND U8657 ( .A(n1968), .B(n1969), .Z(n1966) );
  AND U8658 ( .A(b[21]), .B(a[101]), .Z(n1965) );
  XOR U8659 ( .A(n1970), .B(n1595), .Z(n1597) );
  XOR U8660 ( .A(n1971), .B(n1972), .Z(n1595) );
  AND U8661 ( .A(n1973), .B(n1974), .Z(n1971) );
  AND U8662 ( .A(b[20]), .B(a[102]), .Z(n1970) );
  XOR U8663 ( .A(n1975), .B(n1600), .Z(n1602) );
  XOR U8664 ( .A(n1976), .B(n1977), .Z(n1600) );
  AND U8665 ( .A(n1978), .B(n1979), .Z(n1976) );
  AND U8666 ( .A(b[19]), .B(a[103]), .Z(n1975) );
  XOR U8667 ( .A(n1980), .B(n1605), .Z(n1607) );
  XOR U8668 ( .A(n1981), .B(n1982), .Z(n1605) );
  AND U8669 ( .A(n1983), .B(n1984), .Z(n1981) );
  AND U8670 ( .A(b[18]), .B(a[104]), .Z(n1980) );
  XOR U8671 ( .A(n1985), .B(n1986), .Z(n1609) );
  AND U8672 ( .A(n1987), .B(n1988), .Z(n1985) );
  XOR U8673 ( .A(n1989), .B(n1614), .Z(n1616) );
  XOR U8674 ( .A(n1990), .B(n1991), .Z(n1614) );
  AND U8675 ( .A(n1992), .B(n1993), .Z(n1990) );
  AND U8676 ( .A(b[17]), .B(a[105]), .Z(n1989) );
  XOR U8677 ( .A(n1994), .B(n1619), .Z(n1621) );
  XOR U8678 ( .A(n1995), .B(n1996), .Z(n1619) );
  AND U8679 ( .A(n1997), .B(n1998), .Z(n1995) );
  AND U8680 ( .A(b[15]), .B(a[107]), .Z(n1994) );
  XOR U8681 ( .A(n1999), .B(n1624), .Z(n1626) );
  XOR U8682 ( .A(n2000), .B(n2001), .Z(n1624) );
  AND U8683 ( .A(n2002), .B(n2003), .Z(n2000) );
  AND U8684 ( .A(b[14]), .B(a[108]), .Z(n1999) );
  XOR U8685 ( .A(n2004), .B(n1629), .Z(n1631) );
  XOR U8686 ( .A(n2005), .B(n2006), .Z(n1629) );
  AND U8687 ( .A(n2007), .B(n2008), .Z(n2005) );
  AND U8688 ( .A(b[13]), .B(a[109]), .Z(n2004) );
  XOR U8689 ( .A(n2009), .B(n1634), .Z(n1636) );
  XOR U8690 ( .A(n2010), .B(n2011), .Z(n1634) );
  AND U8691 ( .A(n2012), .B(n2013), .Z(n2010) );
  AND U8692 ( .A(b[12]), .B(a[110]), .Z(n2009) );
  XOR U8693 ( .A(n2014), .B(n1639), .Z(n1641) );
  XOR U8694 ( .A(n2015), .B(n2016), .Z(n1639) );
  AND U8695 ( .A(n2017), .B(n2018), .Z(n2015) );
  AND U8696 ( .A(b[11]), .B(a[111]), .Z(n2014) );
  XOR U8697 ( .A(n2019), .B(n1644), .Z(n1646) );
  XOR U8698 ( .A(n2020), .B(n2021), .Z(n1644) );
  AND U8699 ( .A(n2022), .B(n2023), .Z(n2020) );
  AND U8700 ( .A(b[10]), .B(a[112]), .Z(n2019) );
  XOR U8701 ( .A(n2024), .B(n1649), .Z(n1651) );
  XOR U8702 ( .A(n2025), .B(n2026), .Z(n1649) );
  AND U8703 ( .A(n2027), .B(n2028), .Z(n2025) );
  AND U8704 ( .A(b[9]), .B(a[113]), .Z(n2024) );
  XOR U8705 ( .A(n2029), .B(n1654), .Z(n1656) );
  XOR U8706 ( .A(n2030), .B(n2031), .Z(n1654) );
  AND U8707 ( .A(n2032), .B(n2033), .Z(n2030) );
  AND U8708 ( .A(b[8]), .B(a[114]), .Z(n2029) );
  XOR U8709 ( .A(n2034), .B(n1659), .Z(n1661) );
  XOR U8710 ( .A(n2035), .B(n2036), .Z(n1659) );
  AND U8711 ( .A(n2037), .B(n2038), .Z(n2035) );
  AND U8712 ( .A(b[7]), .B(a[115]), .Z(n2034) );
  XOR U8713 ( .A(n2039), .B(n1664), .Z(n1666) );
  XOR U8714 ( .A(n2040), .B(n2041), .Z(n1664) );
  AND U8715 ( .A(n2042), .B(n2043), .Z(n2040) );
  AND U8716 ( .A(b[6]), .B(a[116]), .Z(n2039) );
  XOR U8717 ( .A(n2044), .B(n1669), .Z(n1671) );
  XOR U8718 ( .A(n2045), .B(n2046), .Z(n1669) );
  AND U8719 ( .A(n2047), .B(n2048), .Z(n2045) );
  AND U8720 ( .A(b[5]), .B(a[117]), .Z(n2044) );
  XOR U8721 ( .A(n2049), .B(n1674), .Z(n1676) );
  XOR U8722 ( .A(n2050), .B(n2051), .Z(n1674) );
  AND U8723 ( .A(n2052), .B(n2053), .Z(n2050) );
  AND U8724 ( .A(b[4]), .B(a[118]), .Z(n2049) );
  XNOR U8725 ( .A(n2054), .B(n2055), .Z(n1688) );
  NANDN U8726 ( .A(n2056), .B(n2057), .Z(n2055) );
  XOR U8727 ( .A(n2058), .B(n1679), .Z(n1681) );
  XNOR U8728 ( .A(n2059), .B(n2060), .Z(n1679) );
  AND U8729 ( .A(n2061), .B(n2062), .Z(n2059) );
  AND U8730 ( .A(b[3]), .B(a[119]), .Z(n2058) );
  XOR U8731 ( .A(n2063), .B(n2064), .Z(swire[121]) );
  XOR U8732 ( .A(n1698), .B(n2065), .Z(n2064) );
  XNOR U8733 ( .A(n1697), .B(n2063), .Z(n2065) );
  NAND U8734 ( .A(a[121]), .B(b[0]), .Z(n1697) );
  XNOR U8735 ( .A(n2056), .B(n2057), .Z(n1698) );
  XOR U8736 ( .A(n2054), .B(n2066), .Z(n2057) );
  NAND U8737 ( .A(b[1]), .B(a[120]), .Z(n2066) );
  XOR U8738 ( .A(n2062), .B(n2067), .Z(n2056) );
  XOR U8739 ( .A(n2054), .B(n2061), .Z(n2067) );
  XNOR U8740 ( .A(n2068), .B(n2060), .Z(n2061) );
  AND U8741 ( .A(b[2]), .B(a[119]), .Z(n2068) );
  NANDN U8742 ( .A(n2069), .B(n2070), .Z(n2054) );
  XOR U8743 ( .A(n2060), .B(n2052), .Z(n2071) );
  XNOR U8744 ( .A(n2051), .B(n2047), .Z(n2072) );
  XNOR U8745 ( .A(n2046), .B(n2042), .Z(n2073) );
  XNOR U8746 ( .A(n2041), .B(n2037), .Z(n2074) );
  XNOR U8747 ( .A(n2036), .B(n2032), .Z(n2075) );
  XNOR U8748 ( .A(n2031), .B(n2027), .Z(n2076) );
  XNOR U8749 ( .A(n2026), .B(n2022), .Z(n2077) );
  XNOR U8750 ( .A(n2021), .B(n2017), .Z(n2078) );
  XNOR U8751 ( .A(n2016), .B(n2012), .Z(n2079) );
  XNOR U8752 ( .A(n2011), .B(n2007), .Z(n2080) );
  XNOR U8753 ( .A(n2006), .B(n2002), .Z(n2081) );
  XNOR U8754 ( .A(n2001), .B(n1997), .Z(n2082) );
  XNOR U8755 ( .A(n1988), .B(n1987), .Z(n2083) );
  XOR U8756 ( .A(n2084), .B(n1986), .Z(n1987) );
  AND U8757 ( .A(b[15]), .B(a[106]), .Z(n2084) );
  XNOR U8758 ( .A(n1986), .B(n1992), .Z(n2085) );
  XNOR U8759 ( .A(n1991), .B(n1983), .Z(n2086) );
  XNOR U8760 ( .A(n1982), .B(n1978), .Z(n2087) );
  XNOR U8761 ( .A(n1977), .B(n1973), .Z(n2088) );
  XNOR U8762 ( .A(n1972), .B(n1968), .Z(n2089) );
  XNOR U8763 ( .A(n1959), .B(n1958), .Z(n2090) );
  XOR U8764 ( .A(n2091), .B(n1957), .Z(n1958) );
  AND U8765 ( .A(b[21]), .B(a[100]), .Z(n2091) );
  XNOR U8766 ( .A(n1957), .B(n1963), .Z(n2092) );
  XNOR U8767 ( .A(n1962), .B(n1954), .Z(n2093) );
  XNOR U8768 ( .A(n1953), .B(n1949), .Z(n2094) );
  XNOR U8769 ( .A(n1948), .B(n1944), .Z(n2095) );
  XNOR U8770 ( .A(n1943), .B(n1939), .Z(n2096) );
  XNOR U8771 ( .A(n1930), .B(n1929), .Z(n2097) );
  XOR U8772 ( .A(n2098), .B(n1928), .Z(n1929) );
  AND U8773 ( .A(b[27]), .B(a[94]), .Z(n2098) );
  XNOR U8774 ( .A(n1928), .B(n1934), .Z(n2099) );
  XNOR U8775 ( .A(n1933), .B(n1925), .Z(n2100) );
  XNOR U8776 ( .A(n1924), .B(n1920), .Z(n2101) );
  XNOR U8777 ( .A(n1919), .B(n1915), .Z(n2102) );
  XNOR U8778 ( .A(n1914), .B(n1910), .Z(n2103) );
  XNOR U8779 ( .A(n1901), .B(n1900), .Z(n2104) );
  XOR U8780 ( .A(n2105), .B(n1899), .Z(n1900) );
  AND U8781 ( .A(b[33]), .B(a[88]), .Z(n2105) );
  XNOR U8782 ( .A(n1899), .B(n1905), .Z(n2106) );
  XNOR U8783 ( .A(n1904), .B(n1896), .Z(n2107) );
  XNOR U8784 ( .A(n1895), .B(n1891), .Z(n2108) );
  XNOR U8785 ( .A(n1890), .B(n1886), .Z(n2109) );
  XNOR U8786 ( .A(n1885), .B(n1881), .Z(n2110) );
  XNOR U8787 ( .A(n1872), .B(n1871), .Z(n2111) );
  XOR U8788 ( .A(n2112), .B(n1870), .Z(n1871) );
  AND U8789 ( .A(b[39]), .B(a[82]), .Z(n2112) );
  XNOR U8790 ( .A(n1870), .B(n1876), .Z(n2113) );
  XNOR U8791 ( .A(n1875), .B(n1867), .Z(n2114) );
  XNOR U8792 ( .A(n1866), .B(n1862), .Z(n2115) );
  XNOR U8793 ( .A(n1861), .B(n1857), .Z(n2116) );
  XNOR U8794 ( .A(n1856), .B(n1852), .Z(n2117) );
  XNOR U8795 ( .A(n1843), .B(n1842), .Z(n2118) );
  XOR U8796 ( .A(n2119), .B(n1841), .Z(n1842) );
  AND U8797 ( .A(b[45]), .B(a[76]), .Z(n2119) );
  XNOR U8798 ( .A(n1841), .B(n1847), .Z(n2120) );
  XNOR U8799 ( .A(n1846), .B(n1838), .Z(n2121) );
  XNOR U8800 ( .A(n1837), .B(n1833), .Z(n2122) );
  XNOR U8801 ( .A(n1832), .B(n1828), .Z(n2123) );
  XNOR U8802 ( .A(n1827), .B(n1823), .Z(n2124) );
  XNOR U8803 ( .A(n1814), .B(n1813), .Z(n2125) );
  XOR U8804 ( .A(n2126), .B(n1812), .Z(n1813) );
  AND U8805 ( .A(b[51]), .B(a[70]), .Z(n2126) );
  XNOR U8806 ( .A(n1812), .B(n1818), .Z(n2127) );
  XNOR U8807 ( .A(n1817), .B(n1809), .Z(n2128) );
  XNOR U8808 ( .A(n1808), .B(n1804), .Z(n2129) );
  XNOR U8809 ( .A(n1803), .B(n1799), .Z(n2130) );
  XNOR U8810 ( .A(n1798), .B(n1794), .Z(n2131) );
  XNOR U8811 ( .A(n1793), .B(n1789), .Z(n2132) );
  XNOR U8812 ( .A(n1788), .B(n1784), .Z(n2133) );
  XNOR U8813 ( .A(n1783), .B(n1779), .Z(n2134) );
  XOR U8814 ( .A(n1778), .B(n1775), .Z(n2135) );
  XOR U8815 ( .A(n2136), .B(n2137), .Z(n1775) );
  XOR U8816 ( .A(n1773), .B(n2138), .Z(n2137) );
  XOR U8817 ( .A(n2139), .B(n2140), .Z(n2138) );
  XOR U8818 ( .A(n2141), .B(n2142), .Z(n2140) );
  NAND U8819 ( .A(a[59]), .B(b[62]), .Z(n2142) );
  AND U8820 ( .A(a[58]), .B(b[63]), .Z(n2141) );
  XOR U8821 ( .A(n2143), .B(n2139), .Z(n2136) );
  XOR U8822 ( .A(n2144), .B(n2145), .Z(n2139) );
  ANDN U8823 ( .B(n2146), .A(n2147), .Z(n2144) );
  AND U8824 ( .A(a[60]), .B(b[61]), .Z(n2143) );
  XOR U8825 ( .A(n2148), .B(n1773), .Z(n1774) );
  XOR U8826 ( .A(n2149), .B(n2150), .Z(n1773) );
  AND U8827 ( .A(n2151), .B(n2152), .Z(n2149) );
  AND U8828 ( .A(b[60]), .B(a[61]), .Z(n2148) );
  XOR U8829 ( .A(n2153), .B(n1778), .Z(n1780) );
  XOR U8830 ( .A(n2154), .B(n2155), .Z(n1778) );
  AND U8831 ( .A(n2156), .B(n2157), .Z(n2154) );
  AND U8832 ( .A(b[59]), .B(a[62]), .Z(n2153) );
  XOR U8833 ( .A(n2158), .B(n1783), .Z(n1785) );
  XOR U8834 ( .A(n2159), .B(n2160), .Z(n1783) );
  AND U8835 ( .A(n2161), .B(n2162), .Z(n2159) );
  AND U8836 ( .A(b[58]), .B(a[63]), .Z(n2158) );
  XOR U8837 ( .A(n2163), .B(n1788), .Z(n1790) );
  XOR U8838 ( .A(n2164), .B(n2165), .Z(n1788) );
  AND U8839 ( .A(n2166), .B(n2167), .Z(n2164) );
  AND U8840 ( .A(b[57]), .B(a[64]), .Z(n2163) );
  XOR U8841 ( .A(n2168), .B(n1793), .Z(n1795) );
  XOR U8842 ( .A(n2169), .B(n2170), .Z(n1793) );
  AND U8843 ( .A(n2171), .B(n2172), .Z(n2169) );
  AND U8844 ( .A(b[56]), .B(a[65]), .Z(n2168) );
  XOR U8845 ( .A(n2173), .B(n1798), .Z(n1800) );
  XOR U8846 ( .A(n2174), .B(n2175), .Z(n1798) );
  AND U8847 ( .A(n2176), .B(n2177), .Z(n2174) );
  AND U8848 ( .A(b[55]), .B(a[66]), .Z(n2173) );
  XOR U8849 ( .A(n2178), .B(n1803), .Z(n1805) );
  XOR U8850 ( .A(n2179), .B(n2180), .Z(n1803) );
  AND U8851 ( .A(n2181), .B(n2182), .Z(n2179) );
  AND U8852 ( .A(b[54]), .B(a[67]), .Z(n2178) );
  XOR U8853 ( .A(n2183), .B(n1808), .Z(n1810) );
  XOR U8854 ( .A(n2184), .B(n2185), .Z(n1808) );
  AND U8855 ( .A(n2186), .B(n2187), .Z(n2184) );
  AND U8856 ( .A(b[53]), .B(a[68]), .Z(n2183) );
  XOR U8857 ( .A(n2188), .B(n2189), .Z(n1812) );
  AND U8858 ( .A(n2190), .B(n2191), .Z(n2188) );
  XOR U8859 ( .A(n2192), .B(n1817), .Z(n1819) );
  XOR U8860 ( .A(n2193), .B(n2194), .Z(n1817) );
  AND U8861 ( .A(n2195), .B(n2196), .Z(n2193) );
  AND U8862 ( .A(b[52]), .B(a[69]), .Z(n2192) );
  XOR U8863 ( .A(n2197), .B(n1822), .Z(n1824) );
  XOR U8864 ( .A(n2198), .B(n2199), .Z(n1822) );
  AND U8865 ( .A(n2200), .B(n2201), .Z(n2198) );
  AND U8866 ( .A(b[50]), .B(a[71]), .Z(n2197) );
  XOR U8867 ( .A(n2202), .B(n1827), .Z(n1829) );
  XOR U8868 ( .A(n2203), .B(n2204), .Z(n1827) );
  AND U8869 ( .A(n2205), .B(n2206), .Z(n2203) );
  AND U8870 ( .A(b[49]), .B(a[72]), .Z(n2202) );
  XOR U8871 ( .A(n2207), .B(n1832), .Z(n1834) );
  XOR U8872 ( .A(n2208), .B(n2209), .Z(n1832) );
  AND U8873 ( .A(n2210), .B(n2211), .Z(n2208) );
  AND U8874 ( .A(b[48]), .B(a[73]), .Z(n2207) );
  XOR U8875 ( .A(n2212), .B(n1837), .Z(n1839) );
  XOR U8876 ( .A(n2213), .B(n2214), .Z(n1837) );
  AND U8877 ( .A(n2215), .B(n2216), .Z(n2213) );
  AND U8878 ( .A(b[47]), .B(a[74]), .Z(n2212) );
  XOR U8879 ( .A(n2217), .B(n2218), .Z(n1841) );
  AND U8880 ( .A(n2219), .B(n2220), .Z(n2217) );
  XOR U8881 ( .A(n2221), .B(n1846), .Z(n1848) );
  XOR U8882 ( .A(n2222), .B(n2223), .Z(n1846) );
  AND U8883 ( .A(n2224), .B(n2225), .Z(n2222) );
  AND U8884 ( .A(b[46]), .B(a[75]), .Z(n2221) );
  XOR U8885 ( .A(n2226), .B(n1851), .Z(n1853) );
  XOR U8886 ( .A(n2227), .B(n2228), .Z(n1851) );
  AND U8887 ( .A(n2229), .B(n2230), .Z(n2227) );
  AND U8888 ( .A(b[44]), .B(a[77]), .Z(n2226) );
  XOR U8889 ( .A(n2231), .B(n1856), .Z(n1858) );
  XOR U8890 ( .A(n2232), .B(n2233), .Z(n1856) );
  AND U8891 ( .A(n2234), .B(n2235), .Z(n2232) );
  AND U8892 ( .A(b[43]), .B(a[78]), .Z(n2231) );
  XOR U8893 ( .A(n2236), .B(n1861), .Z(n1863) );
  XOR U8894 ( .A(n2237), .B(n2238), .Z(n1861) );
  AND U8895 ( .A(n2239), .B(n2240), .Z(n2237) );
  AND U8896 ( .A(b[42]), .B(a[79]), .Z(n2236) );
  XOR U8897 ( .A(n2241), .B(n1866), .Z(n1868) );
  XOR U8898 ( .A(n2242), .B(n2243), .Z(n1866) );
  AND U8899 ( .A(n2244), .B(n2245), .Z(n2242) );
  AND U8900 ( .A(b[41]), .B(a[80]), .Z(n2241) );
  XOR U8901 ( .A(n2246), .B(n2247), .Z(n1870) );
  AND U8902 ( .A(n2248), .B(n2249), .Z(n2246) );
  XOR U8903 ( .A(n2250), .B(n1875), .Z(n1877) );
  XOR U8904 ( .A(n2251), .B(n2252), .Z(n1875) );
  AND U8905 ( .A(n2253), .B(n2254), .Z(n2251) );
  AND U8906 ( .A(b[40]), .B(a[81]), .Z(n2250) );
  XOR U8907 ( .A(n2255), .B(n1880), .Z(n1882) );
  XOR U8908 ( .A(n2256), .B(n2257), .Z(n1880) );
  AND U8909 ( .A(n2258), .B(n2259), .Z(n2256) );
  AND U8910 ( .A(b[38]), .B(a[83]), .Z(n2255) );
  XOR U8911 ( .A(n2260), .B(n1885), .Z(n1887) );
  XOR U8912 ( .A(n2261), .B(n2262), .Z(n1885) );
  AND U8913 ( .A(n2263), .B(n2264), .Z(n2261) );
  AND U8914 ( .A(b[37]), .B(a[84]), .Z(n2260) );
  XOR U8915 ( .A(n2265), .B(n1890), .Z(n1892) );
  XOR U8916 ( .A(n2266), .B(n2267), .Z(n1890) );
  AND U8917 ( .A(n2268), .B(n2269), .Z(n2266) );
  AND U8918 ( .A(b[36]), .B(a[85]), .Z(n2265) );
  XOR U8919 ( .A(n2270), .B(n1895), .Z(n1897) );
  XOR U8920 ( .A(n2271), .B(n2272), .Z(n1895) );
  AND U8921 ( .A(n2273), .B(n2274), .Z(n2271) );
  AND U8922 ( .A(b[35]), .B(a[86]), .Z(n2270) );
  XOR U8923 ( .A(n2275), .B(n2276), .Z(n1899) );
  AND U8924 ( .A(n2277), .B(n2278), .Z(n2275) );
  XOR U8925 ( .A(n2279), .B(n1904), .Z(n1906) );
  XOR U8926 ( .A(n2280), .B(n2281), .Z(n1904) );
  AND U8927 ( .A(n2282), .B(n2283), .Z(n2280) );
  AND U8928 ( .A(b[34]), .B(a[87]), .Z(n2279) );
  XOR U8929 ( .A(n2284), .B(n1909), .Z(n1911) );
  XOR U8930 ( .A(n2285), .B(n2286), .Z(n1909) );
  AND U8931 ( .A(n2287), .B(n2288), .Z(n2285) );
  AND U8932 ( .A(b[32]), .B(a[89]), .Z(n2284) );
  XOR U8933 ( .A(n2289), .B(n1914), .Z(n1916) );
  XOR U8934 ( .A(n2290), .B(n2291), .Z(n1914) );
  AND U8935 ( .A(n2292), .B(n2293), .Z(n2290) );
  AND U8936 ( .A(b[31]), .B(a[90]), .Z(n2289) );
  XOR U8937 ( .A(n2294), .B(n1919), .Z(n1921) );
  XOR U8938 ( .A(n2295), .B(n2296), .Z(n1919) );
  AND U8939 ( .A(n2297), .B(n2298), .Z(n2295) );
  AND U8940 ( .A(b[30]), .B(a[91]), .Z(n2294) );
  XOR U8941 ( .A(n2299), .B(n1924), .Z(n1926) );
  XOR U8942 ( .A(n2300), .B(n2301), .Z(n1924) );
  AND U8943 ( .A(n2302), .B(n2303), .Z(n2300) );
  AND U8944 ( .A(b[29]), .B(a[92]), .Z(n2299) );
  XOR U8945 ( .A(n2304), .B(n2305), .Z(n1928) );
  AND U8946 ( .A(n2306), .B(n2307), .Z(n2304) );
  XOR U8947 ( .A(n2308), .B(n1933), .Z(n1935) );
  XOR U8948 ( .A(n2309), .B(n2310), .Z(n1933) );
  AND U8949 ( .A(n2311), .B(n2312), .Z(n2309) );
  AND U8950 ( .A(b[28]), .B(a[93]), .Z(n2308) );
  XOR U8951 ( .A(n2313), .B(n1938), .Z(n1940) );
  XOR U8952 ( .A(n2314), .B(n2315), .Z(n1938) );
  AND U8953 ( .A(n2316), .B(n2317), .Z(n2314) );
  AND U8954 ( .A(b[26]), .B(a[95]), .Z(n2313) );
  XOR U8955 ( .A(n2318), .B(n1943), .Z(n1945) );
  XOR U8956 ( .A(n2319), .B(n2320), .Z(n1943) );
  AND U8957 ( .A(n2321), .B(n2322), .Z(n2319) );
  AND U8958 ( .A(b[25]), .B(a[96]), .Z(n2318) );
  XOR U8959 ( .A(n2323), .B(n1948), .Z(n1950) );
  XOR U8960 ( .A(n2324), .B(n2325), .Z(n1948) );
  AND U8961 ( .A(n2326), .B(n2327), .Z(n2324) );
  AND U8962 ( .A(b[24]), .B(a[97]), .Z(n2323) );
  XOR U8963 ( .A(n2328), .B(n1953), .Z(n1955) );
  XOR U8964 ( .A(n2329), .B(n2330), .Z(n1953) );
  AND U8965 ( .A(n2331), .B(n2332), .Z(n2329) );
  AND U8966 ( .A(b[23]), .B(a[98]), .Z(n2328) );
  XOR U8967 ( .A(n2333), .B(n2334), .Z(n1957) );
  AND U8968 ( .A(n2335), .B(n2336), .Z(n2333) );
  XOR U8969 ( .A(n2337), .B(n1962), .Z(n1964) );
  XOR U8970 ( .A(n2338), .B(n2339), .Z(n1962) );
  AND U8971 ( .A(n2340), .B(n2341), .Z(n2338) );
  AND U8972 ( .A(b[22]), .B(a[99]), .Z(n2337) );
  XOR U8973 ( .A(n2342), .B(n1967), .Z(n1969) );
  XOR U8974 ( .A(n2343), .B(n2344), .Z(n1967) );
  AND U8975 ( .A(n2345), .B(n2346), .Z(n2343) );
  AND U8976 ( .A(b[20]), .B(a[101]), .Z(n2342) );
  XOR U8977 ( .A(n2347), .B(n1972), .Z(n1974) );
  XOR U8978 ( .A(n2348), .B(n2349), .Z(n1972) );
  AND U8979 ( .A(n2350), .B(n2351), .Z(n2348) );
  AND U8980 ( .A(b[19]), .B(a[102]), .Z(n2347) );
  XOR U8981 ( .A(n2352), .B(n1977), .Z(n1979) );
  XOR U8982 ( .A(n2353), .B(n2354), .Z(n1977) );
  AND U8983 ( .A(n2355), .B(n2356), .Z(n2353) );
  AND U8984 ( .A(b[18]), .B(a[103]), .Z(n2352) );
  XOR U8985 ( .A(n2357), .B(n1982), .Z(n1984) );
  XOR U8986 ( .A(n2358), .B(n2359), .Z(n1982) );
  AND U8987 ( .A(n2360), .B(n2361), .Z(n2358) );
  AND U8988 ( .A(b[17]), .B(a[104]), .Z(n2357) );
  XOR U8989 ( .A(n2362), .B(n2363), .Z(n1986) );
  AND U8990 ( .A(n2364), .B(n2365), .Z(n2362) );
  XOR U8991 ( .A(n2366), .B(n1991), .Z(n1993) );
  XOR U8992 ( .A(n2367), .B(n2368), .Z(n1991) );
  AND U8993 ( .A(n2369), .B(n2370), .Z(n2367) );
  AND U8994 ( .A(b[16]), .B(a[105]), .Z(n2366) );
  XOR U8995 ( .A(n2371), .B(n1996), .Z(n1998) );
  XOR U8996 ( .A(n2372), .B(n2373), .Z(n1996) );
  AND U8997 ( .A(n2374), .B(n2375), .Z(n2372) );
  AND U8998 ( .A(b[14]), .B(a[107]), .Z(n2371) );
  XOR U8999 ( .A(n2376), .B(n2001), .Z(n2003) );
  XOR U9000 ( .A(n2377), .B(n2378), .Z(n2001) );
  AND U9001 ( .A(n2379), .B(n2380), .Z(n2377) );
  AND U9002 ( .A(b[13]), .B(a[108]), .Z(n2376) );
  XOR U9003 ( .A(n2381), .B(n2006), .Z(n2008) );
  XOR U9004 ( .A(n2382), .B(n2383), .Z(n2006) );
  AND U9005 ( .A(n2384), .B(n2385), .Z(n2382) );
  AND U9006 ( .A(b[12]), .B(a[109]), .Z(n2381) );
  XOR U9007 ( .A(n2386), .B(n2011), .Z(n2013) );
  XOR U9008 ( .A(n2387), .B(n2388), .Z(n2011) );
  AND U9009 ( .A(n2389), .B(n2390), .Z(n2387) );
  AND U9010 ( .A(b[11]), .B(a[110]), .Z(n2386) );
  XOR U9011 ( .A(n2391), .B(n2016), .Z(n2018) );
  XOR U9012 ( .A(n2392), .B(n2393), .Z(n2016) );
  AND U9013 ( .A(n2394), .B(n2395), .Z(n2392) );
  AND U9014 ( .A(b[10]), .B(a[111]), .Z(n2391) );
  XOR U9015 ( .A(n2396), .B(n2021), .Z(n2023) );
  XOR U9016 ( .A(n2397), .B(n2398), .Z(n2021) );
  AND U9017 ( .A(n2399), .B(n2400), .Z(n2397) );
  AND U9018 ( .A(b[9]), .B(a[112]), .Z(n2396) );
  XOR U9019 ( .A(n2401), .B(n2026), .Z(n2028) );
  XOR U9020 ( .A(n2402), .B(n2403), .Z(n2026) );
  AND U9021 ( .A(n2404), .B(n2405), .Z(n2402) );
  AND U9022 ( .A(b[8]), .B(a[113]), .Z(n2401) );
  XOR U9023 ( .A(n2406), .B(n2031), .Z(n2033) );
  XOR U9024 ( .A(n2407), .B(n2408), .Z(n2031) );
  AND U9025 ( .A(n2409), .B(n2410), .Z(n2407) );
  AND U9026 ( .A(b[7]), .B(a[114]), .Z(n2406) );
  XOR U9027 ( .A(n2411), .B(n2036), .Z(n2038) );
  XOR U9028 ( .A(n2412), .B(n2413), .Z(n2036) );
  AND U9029 ( .A(n2414), .B(n2415), .Z(n2412) );
  AND U9030 ( .A(b[6]), .B(a[115]), .Z(n2411) );
  XOR U9031 ( .A(n2416), .B(n2041), .Z(n2043) );
  XOR U9032 ( .A(n2417), .B(n2418), .Z(n2041) );
  AND U9033 ( .A(n2419), .B(n2420), .Z(n2417) );
  AND U9034 ( .A(b[5]), .B(a[116]), .Z(n2416) );
  XOR U9035 ( .A(n2421), .B(n2046), .Z(n2048) );
  XOR U9036 ( .A(n2422), .B(n2423), .Z(n2046) );
  AND U9037 ( .A(n2424), .B(n2425), .Z(n2422) );
  AND U9038 ( .A(b[4]), .B(a[117]), .Z(n2421) );
  XNOR U9039 ( .A(n2426), .B(n2427), .Z(n2060) );
  NANDN U9040 ( .A(n2428), .B(n2429), .Z(n2427) );
  XOR U9041 ( .A(n2430), .B(n2051), .Z(n2053) );
  XNOR U9042 ( .A(n2431), .B(n2432), .Z(n2051) );
  AND U9043 ( .A(n2433), .B(n2434), .Z(n2431) );
  AND U9044 ( .A(b[3]), .B(a[118]), .Z(n2430) );
  XOR U9045 ( .A(n2435), .B(n2436), .Z(swire[120]) );
  XOR U9046 ( .A(n2070), .B(n2437), .Z(n2436) );
  XNOR U9047 ( .A(n2069), .B(n2435), .Z(n2437) );
  NAND U9048 ( .A(a[120]), .B(b[0]), .Z(n2069) );
  XNOR U9049 ( .A(n2428), .B(n2429), .Z(n2070) );
  XOR U9050 ( .A(n2426), .B(n2438), .Z(n2429) );
  NAND U9051 ( .A(b[1]), .B(a[119]), .Z(n2438) );
  XOR U9052 ( .A(n2433), .B(n2439), .Z(n2428) );
  XOR U9053 ( .A(n2426), .B(n2434), .Z(n2439) );
  XNOR U9054 ( .A(n2440), .B(n2432), .Z(n2434) );
  AND U9055 ( .A(b[2]), .B(a[118]), .Z(n2440) );
  NANDN U9056 ( .A(n2441), .B(n2442), .Z(n2426) );
  XOR U9057 ( .A(n2432), .B(n2424), .Z(n2443) );
  XNOR U9058 ( .A(n2423), .B(n2419), .Z(n2444) );
  XNOR U9059 ( .A(n2418), .B(n2414), .Z(n2445) );
  XNOR U9060 ( .A(n2413), .B(n2409), .Z(n2446) );
  XNOR U9061 ( .A(n2408), .B(n2404), .Z(n2447) );
  XNOR U9062 ( .A(n2403), .B(n2399), .Z(n2448) );
  XNOR U9063 ( .A(n2398), .B(n2394), .Z(n2449) );
  XNOR U9064 ( .A(n2393), .B(n2389), .Z(n2450) );
  XNOR U9065 ( .A(n2388), .B(n2384), .Z(n2451) );
  XNOR U9066 ( .A(n2383), .B(n2379), .Z(n2452) );
  XNOR U9067 ( .A(n2378), .B(n2374), .Z(n2453) );
  XOR U9068 ( .A(n2454), .B(n2455), .Z(n2374) );
  XNOR U9069 ( .A(n2365), .B(n2364), .Z(n2455) );
  XOR U9070 ( .A(n2456), .B(n2363), .Z(n2364) );
  AND U9071 ( .A(b[14]), .B(a[106]), .Z(n2456) );
  XNOR U9072 ( .A(n2363), .B(n2369), .Z(n2457) );
  XNOR U9073 ( .A(n2368), .B(n2360), .Z(n2458) );
  XNOR U9074 ( .A(n2359), .B(n2355), .Z(n2459) );
  XNOR U9075 ( .A(n2354), .B(n2350), .Z(n2460) );
  XNOR U9076 ( .A(n2349), .B(n2345), .Z(n2461) );
  XNOR U9077 ( .A(n2336), .B(n2335), .Z(n2462) );
  XOR U9078 ( .A(n2463), .B(n2334), .Z(n2335) );
  AND U9079 ( .A(b[20]), .B(a[100]), .Z(n2463) );
  XNOR U9080 ( .A(n2334), .B(n2340), .Z(n2464) );
  XNOR U9081 ( .A(n2339), .B(n2331), .Z(n2465) );
  XNOR U9082 ( .A(n2330), .B(n2326), .Z(n2466) );
  XNOR U9083 ( .A(n2325), .B(n2321), .Z(n2467) );
  XNOR U9084 ( .A(n2320), .B(n2316), .Z(n2468) );
  XNOR U9085 ( .A(n2307), .B(n2306), .Z(n2469) );
  XOR U9086 ( .A(n2470), .B(n2305), .Z(n2306) );
  AND U9087 ( .A(b[26]), .B(a[94]), .Z(n2470) );
  XNOR U9088 ( .A(n2305), .B(n2311), .Z(n2471) );
  XNOR U9089 ( .A(n2310), .B(n2302), .Z(n2472) );
  XNOR U9090 ( .A(n2301), .B(n2297), .Z(n2473) );
  XNOR U9091 ( .A(n2296), .B(n2292), .Z(n2474) );
  XNOR U9092 ( .A(n2291), .B(n2287), .Z(n2475) );
  XNOR U9093 ( .A(n2278), .B(n2277), .Z(n2476) );
  XOR U9094 ( .A(n2477), .B(n2276), .Z(n2277) );
  AND U9095 ( .A(b[32]), .B(a[88]), .Z(n2477) );
  XNOR U9096 ( .A(n2276), .B(n2282), .Z(n2478) );
  XNOR U9097 ( .A(n2281), .B(n2273), .Z(n2479) );
  XNOR U9098 ( .A(n2272), .B(n2268), .Z(n2480) );
  XNOR U9099 ( .A(n2267), .B(n2263), .Z(n2481) );
  XNOR U9100 ( .A(n2262), .B(n2258), .Z(n2482) );
  XNOR U9101 ( .A(n2249), .B(n2248), .Z(n2483) );
  XOR U9102 ( .A(n2484), .B(n2247), .Z(n2248) );
  AND U9103 ( .A(b[38]), .B(a[82]), .Z(n2484) );
  XNOR U9104 ( .A(n2247), .B(n2253), .Z(n2485) );
  XNOR U9105 ( .A(n2252), .B(n2244), .Z(n2486) );
  XNOR U9106 ( .A(n2243), .B(n2239), .Z(n2487) );
  XNOR U9107 ( .A(n2238), .B(n2234), .Z(n2488) );
  XNOR U9108 ( .A(n2233), .B(n2229), .Z(n2489) );
  XNOR U9109 ( .A(n2220), .B(n2219), .Z(n2490) );
  XOR U9110 ( .A(n2491), .B(n2218), .Z(n2219) );
  AND U9111 ( .A(b[44]), .B(a[76]), .Z(n2491) );
  XNOR U9112 ( .A(n2218), .B(n2224), .Z(n2492) );
  XNOR U9113 ( .A(n2223), .B(n2215), .Z(n2493) );
  XNOR U9114 ( .A(n2214), .B(n2210), .Z(n2494) );
  XNOR U9115 ( .A(n2209), .B(n2205), .Z(n2495) );
  XNOR U9116 ( .A(n2204), .B(n2200), .Z(n2496) );
  XNOR U9117 ( .A(n2191), .B(n2190), .Z(n2497) );
  XOR U9118 ( .A(n2498), .B(n2189), .Z(n2190) );
  AND U9119 ( .A(b[50]), .B(a[70]), .Z(n2498) );
  XNOR U9120 ( .A(n2189), .B(n2195), .Z(n2499) );
  XNOR U9121 ( .A(n2194), .B(n2186), .Z(n2500) );
  XNOR U9122 ( .A(n2185), .B(n2181), .Z(n2501) );
  XNOR U9123 ( .A(n2180), .B(n2176), .Z(n2502) );
  XNOR U9124 ( .A(n2175), .B(n2171), .Z(n2503) );
  XNOR U9125 ( .A(n2170), .B(n2166), .Z(n2504) );
  XNOR U9126 ( .A(n2165), .B(n2161), .Z(n2505) );
  XNOR U9127 ( .A(n2160), .B(n2156), .Z(n2506) );
  XNOR U9128 ( .A(n2155), .B(n2151), .Z(n2507) );
  XOR U9129 ( .A(n2150), .B(n2147), .Z(n2508) );
  XOR U9130 ( .A(n2509), .B(n2510), .Z(n2147) );
  XOR U9131 ( .A(n2145), .B(n2511), .Z(n2510) );
  XOR U9132 ( .A(n2512), .B(n2513), .Z(n2511) );
  XOR U9133 ( .A(n2514), .B(n2515), .Z(n2513) );
  NAND U9134 ( .A(a[58]), .B(b[62]), .Z(n2515) );
  AND U9135 ( .A(a[57]), .B(b[63]), .Z(n2514) );
  XOR U9136 ( .A(n2516), .B(n2512), .Z(n2509) );
  XOR U9137 ( .A(n2517), .B(n2518), .Z(n2512) );
  ANDN U9138 ( .B(n2519), .A(n2520), .Z(n2517) );
  AND U9139 ( .A(a[59]), .B(b[61]), .Z(n2516) );
  XOR U9140 ( .A(n2521), .B(n2145), .Z(n2146) );
  XOR U9141 ( .A(n2522), .B(n2523), .Z(n2145) );
  AND U9142 ( .A(n2524), .B(n2525), .Z(n2522) );
  AND U9143 ( .A(a[60]), .B(b[60]), .Z(n2521) );
  XOR U9144 ( .A(n2526), .B(n2150), .Z(n2152) );
  XOR U9145 ( .A(n2527), .B(n2528), .Z(n2150) );
  AND U9146 ( .A(n2529), .B(n2530), .Z(n2527) );
  AND U9147 ( .A(b[59]), .B(a[61]), .Z(n2526) );
  XOR U9148 ( .A(n2531), .B(n2155), .Z(n2157) );
  XOR U9149 ( .A(n2532), .B(n2533), .Z(n2155) );
  AND U9150 ( .A(n2534), .B(n2535), .Z(n2532) );
  AND U9151 ( .A(b[58]), .B(a[62]), .Z(n2531) );
  XOR U9152 ( .A(n2536), .B(n2160), .Z(n2162) );
  XOR U9153 ( .A(n2537), .B(n2538), .Z(n2160) );
  AND U9154 ( .A(n2539), .B(n2540), .Z(n2537) );
  AND U9155 ( .A(b[57]), .B(a[63]), .Z(n2536) );
  XOR U9156 ( .A(n2541), .B(n2165), .Z(n2167) );
  XOR U9157 ( .A(n2542), .B(n2543), .Z(n2165) );
  AND U9158 ( .A(n2544), .B(n2545), .Z(n2542) );
  AND U9159 ( .A(b[56]), .B(a[64]), .Z(n2541) );
  XOR U9160 ( .A(n2546), .B(n2170), .Z(n2172) );
  XOR U9161 ( .A(n2547), .B(n2548), .Z(n2170) );
  AND U9162 ( .A(n2549), .B(n2550), .Z(n2547) );
  AND U9163 ( .A(b[55]), .B(a[65]), .Z(n2546) );
  XOR U9164 ( .A(n2551), .B(n2175), .Z(n2177) );
  XOR U9165 ( .A(n2552), .B(n2553), .Z(n2175) );
  AND U9166 ( .A(n2554), .B(n2555), .Z(n2552) );
  AND U9167 ( .A(b[54]), .B(a[66]), .Z(n2551) );
  XOR U9168 ( .A(n2556), .B(n2180), .Z(n2182) );
  XOR U9169 ( .A(n2557), .B(n2558), .Z(n2180) );
  AND U9170 ( .A(n2559), .B(n2560), .Z(n2557) );
  AND U9171 ( .A(b[53]), .B(a[67]), .Z(n2556) );
  XOR U9172 ( .A(n2561), .B(n2185), .Z(n2187) );
  XOR U9173 ( .A(n2562), .B(n2563), .Z(n2185) );
  AND U9174 ( .A(n2564), .B(n2565), .Z(n2562) );
  AND U9175 ( .A(b[52]), .B(a[68]), .Z(n2561) );
  XOR U9176 ( .A(n2566), .B(n2567), .Z(n2189) );
  AND U9177 ( .A(n2568), .B(n2569), .Z(n2566) );
  XOR U9178 ( .A(n2570), .B(n2194), .Z(n2196) );
  XOR U9179 ( .A(n2571), .B(n2572), .Z(n2194) );
  AND U9180 ( .A(n2573), .B(n2574), .Z(n2571) );
  AND U9181 ( .A(b[51]), .B(a[69]), .Z(n2570) );
  XOR U9182 ( .A(n2575), .B(n2199), .Z(n2201) );
  XOR U9183 ( .A(n2576), .B(n2577), .Z(n2199) );
  AND U9184 ( .A(n2578), .B(n2579), .Z(n2576) );
  AND U9185 ( .A(b[49]), .B(a[71]), .Z(n2575) );
  XOR U9186 ( .A(n2580), .B(n2204), .Z(n2206) );
  XOR U9187 ( .A(n2581), .B(n2582), .Z(n2204) );
  AND U9188 ( .A(n2583), .B(n2584), .Z(n2581) );
  AND U9189 ( .A(b[48]), .B(a[72]), .Z(n2580) );
  XOR U9190 ( .A(n2585), .B(n2209), .Z(n2211) );
  XOR U9191 ( .A(n2586), .B(n2587), .Z(n2209) );
  AND U9192 ( .A(n2588), .B(n2589), .Z(n2586) );
  AND U9193 ( .A(b[47]), .B(a[73]), .Z(n2585) );
  XOR U9194 ( .A(n2590), .B(n2214), .Z(n2216) );
  XOR U9195 ( .A(n2591), .B(n2592), .Z(n2214) );
  AND U9196 ( .A(n2593), .B(n2594), .Z(n2591) );
  AND U9197 ( .A(b[46]), .B(a[74]), .Z(n2590) );
  XOR U9198 ( .A(n2595), .B(n2596), .Z(n2218) );
  AND U9199 ( .A(n2597), .B(n2598), .Z(n2595) );
  XOR U9200 ( .A(n2599), .B(n2223), .Z(n2225) );
  XOR U9201 ( .A(n2600), .B(n2601), .Z(n2223) );
  AND U9202 ( .A(n2602), .B(n2603), .Z(n2600) );
  AND U9203 ( .A(b[45]), .B(a[75]), .Z(n2599) );
  XOR U9204 ( .A(n2604), .B(n2228), .Z(n2230) );
  XOR U9205 ( .A(n2605), .B(n2606), .Z(n2228) );
  AND U9206 ( .A(n2607), .B(n2608), .Z(n2605) );
  AND U9207 ( .A(b[43]), .B(a[77]), .Z(n2604) );
  XOR U9208 ( .A(n2609), .B(n2233), .Z(n2235) );
  XOR U9209 ( .A(n2610), .B(n2611), .Z(n2233) );
  AND U9210 ( .A(n2612), .B(n2613), .Z(n2610) );
  AND U9211 ( .A(b[42]), .B(a[78]), .Z(n2609) );
  XOR U9212 ( .A(n2614), .B(n2238), .Z(n2240) );
  XOR U9213 ( .A(n2615), .B(n2616), .Z(n2238) );
  AND U9214 ( .A(n2617), .B(n2618), .Z(n2615) );
  AND U9215 ( .A(b[41]), .B(a[79]), .Z(n2614) );
  XOR U9216 ( .A(n2619), .B(n2243), .Z(n2245) );
  XOR U9217 ( .A(n2620), .B(n2621), .Z(n2243) );
  AND U9218 ( .A(n2622), .B(n2623), .Z(n2620) );
  AND U9219 ( .A(b[40]), .B(a[80]), .Z(n2619) );
  XOR U9220 ( .A(n2624), .B(n2625), .Z(n2247) );
  AND U9221 ( .A(n2626), .B(n2627), .Z(n2624) );
  XOR U9222 ( .A(n2628), .B(n2252), .Z(n2254) );
  XOR U9223 ( .A(n2629), .B(n2630), .Z(n2252) );
  AND U9224 ( .A(n2631), .B(n2632), .Z(n2629) );
  AND U9225 ( .A(b[39]), .B(a[81]), .Z(n2628) );
  XOR U9226 ( .A(n2633), .B(n2257), .Z(n2259) );
  XOR U9227 ( .A(n2634), .B(n2635), .Z(n2257) );
  AND U9228 ( .A(n2636), .B(n2637), .Z(n2634) );
  AND U9229 ( .A(b[37]), .B(a[83]), .Z(n2633) );
  XOR U9230 ( .A(n2638), .B(n2262), .Z(n2264) );
  XOR U9231 ( .A(n2639), .B(n2640), .Z(n2262) );
  AND U9232 ( .A(n2641), .B(n2642), .Z(n2639) );
  AND U9233 ( .A(b[36]), .B(a[84]), .Z(n2638) );
  XOR U9234 ( .A(n2643), .B(n2267), .Z(n2269) );
  XOR U9235 ( .A(n2644), .B(n2645), .Z(n2267) );
  AND U9236 ( .A(n2646), .B(n2647), .Z(n2644) );
  AND U9237 ( .A(b[35]), .B(a[85]), .Z(n2643) );
  XOR U9238 ( .A(n2648), .B(n2272), .Z(n2274) );
  XOR U9239 ( .A(n2649), .B(n2650), .Z(n2272) );
  AND U9240 ( .A(n2651), .B(n2652), .Z(n2649) );
  AND U9241 ( .A(b[34]), .B(a[86]), .Z(n2648) );
  XOR U9242 ( .A(n2653), .B(n2654), .Z(n2276) );
  AND U9243 ( .A(n2655), .B(n2656), .Z(n2653) );
  XOR U9244 ( .A(n2657), .B(n2281), .Z(n2283) );
  XOR U9245 ( .A(n2658), .B(n2659), .Z(n2281) );
  AND U9246 ( .A(n2660), .B(n2661), .Z(n2658) );
  AND U9247 ( .A(b[33]), .B(a[87]), .Z(n2657) );
  XOR U9248 ( .A(n2662), .B(n2286), .Z(n2288) );
  XOR U9249 ( .A(n2663), .B(n2664), .Z(n2286) );
  AND U9250 ( .A(n2665), .B(n2666), .Z(n2663) );
  AND U9251 ( .A(b[31]), .B(a[89]), .Z(n2662) );
  XOR U9252 ( .A(n2667), .B(n2291), .Z(n2293) );
  XOR U9253 ( .A(n2668), .B(n2669), .Z(n2291) );
  AND U9254 ( .A(n2670), .B(n2671), .Z(n2668) );
  AND U9255 ( .A(b[30]), .B(a[90]), .Z(n2667) );
  XOR U9256 ( .A(n2672), .B(n2296), .Z(n2298) );
  XOR U9257 ( .A(n2673), .B(n2674), .Z(n2296) );
  AND U9258 ( .A(n2675), .B(n2676), .Z(n2673) );
  AND U9259 ( .A(b[29]), .B(a[91]), .Z(n2672) );
  XOR U9260 ( .A(n2677), .B(n2301), .Z(n2303) );
  XOR U9261 ( .A(n2678), .B(n2679), .Z(n2301) );
  AND U9262 ( .A(n2680), .B(n2681), .Z(n2678) );
  AND U9263 ( .A(b[28]), .B(a[92]), .Z(n2677) );
  XOR U9264 ( .A(n2682), .B(n2683), .Z(n2305) );
  AND U9265 ( .A(n2684), .B(n2685), .Z(n2682) );
  XOR U9266 ( .A(n2686), .B(n2310), .Z(n2312) );
  XOR U9267 ( .A(n2687), .B(n2688), .Z(n2310) );
  AND U9268 ( .A(n2689), .B(n2690), .Z(n2687) );
  AND U9269 ( .A(b[27]), .B(a[93]), .Z(n2686) );
  XOR U9270 ( .A(n2691), .B(n2315), .Z(n2317) );
  XOR U9271 ( .A(n2692), .B(n2693), .Z(n2315) );
  AND U9272 ( .A(n2694), .B(n2695), .Z(n2692) );
  AND U9273 ( .A(b[25]), .B(a[95]), .Z(n2691) );
  XOR U9274 ( .A(n2696), .B(n2320), .Z(n2322) );
  XOR U9275 ( .A(n2697), .B(n2698), .Z(n2320) );
  AND U9276 ( .A(n2699), .B(n2700), .Z(n2697) );
  AND U9277 ( .A(b[24]), .B(a[96]), .Z(n2696) );
  XOR U9278 ( .A(n2701), .B(n2325), .Z(n2327) );
  XOR U9279 ( .A(n2702), .B(n2703), .Z(n2325) );
  AND U9280 ( .A(n2704), .B(n2705), .Z(n2702) );
  AND U9281 ( .A(b[23]), .B(a[97]), .Z(n2701) );
  XOR U9282 ( .A(n2706), .B(n2330), .Z(n2332) );
  XOR U9283 ( .A(n2707), .B(n2708), .Z(n2330) );
  AND U9284 ( .A(n2709), .B(n2710), .Z(n2707) );
  AND U9285 ( .A(b[22]), .B(a[98]), .Z(n2706) );
  XOR U9286 ( .A(n2711), .B(n2712), .Z(n2334) );
  AND U9287 ( .A(n2713), .B(n2714), .Z(n2711) );
  XOR U9288 ( .A(n2715), .B(n2339), .Z(n2341) );
  XOR U9289 ( .A(n2716), .B(n2717), .Z(n2339) );
  AND U9290 ( .A(n2718), .B(n2719), .Z(n2716) );
  AND U9291 ( .A(b[21]), .B(a[99]), .Z(n2715) );
  XOR U9292 ( .A(n2720), .B(n2344), .Z(n2346) );
  XOR U9293 ( .A(n2721), .B(n2722), .Z(n2344) );
  AND U9294 ( .A(n2723), .B(n2724), .Z(n2721) );
  AND U9295 ( .A(b[19]), .B(a[101]), .Z(n2720) );
  XOR U9296 ( .A(n2725), .B(n2349), .Z(n2351) );
  XOR U9297 ( .A(n2726), .B(n2727), .Z(n2349) );
  AND U9298 ( .A(n2728), .B(n2729), .Z(n2726) );
  AND U9299 ( .A(b[18]), .B(a[102]), .Z(n2725) );
  XOR U9300 ( .A(n2730), .B(n2354), .Z(n2356) );
  XOR U9301 ( .A(n2731), .B(n2732), .Z(n2354) );
  AND U9302 ( .A(n2733), .B(n2734), .Z(n2731) );
  AND U9303 ( .A(b[17]), .B(a[103]), .Z(n2730) );
  XOR U9304 ( .A(n2735), .B(n2359), .Z(n2361) );
  XOR U9305 ( .A(n2736), .B(n2737), .Z(n2359) );
  AND U9306 ( .A(n2738), .B(n2739), .Z(n2736) );
  AND U9307 ( .A(b[16]), .B(a[104]), .Z(n2735) );
  XOR U9308 ( .A(n2740), .B(n2741), .Z(n2363) );
  AND U9309 ( .A(n2742), .B(n2743), .Z(n2740) );
  XOR U9310 ( .A(n2744), .B(n2368), .Z(n2370) );
  XOR U9311 ( .A(n2745), .B(n2746), .Z(n2368) );
  AND U9312 ( .A(n2747), .B(n2748), .Z(n2745) );
  AND U9313 ( .A(b[15]), .B(a[105]), .Z(n2744) );
  IV U9314 ( .A(n2373), .Z(n2454) );
  XOR U9315 ( .A(n2749), .B(n2373), .Z(n2375) );
  XOR U9316 ( .A(n2750), .B(n2751), .Z(n2373) );
  AND U9317 ( .A(n2752), .B(n2753), .Z(n2750) );
  AND U9318 ( .A(b[13]), .B(a[107]), .Z(n2749) );
  XOR U9319 ( .A(n2754), .B(n2378), .Z(n2380) );
  XOR U9320 ( .A(n2755), .B(n2756), .Z(n2378) );
  AND U9321 ( .A(n2757), .B(n2758), .Z(n2755) );
  AND U9322 ( .A(b[12]), .B(a[108]), .Z(n2754) );
  XOR U9323 ( .A(n2759), .B(n2383), .Z(n2385) );
  XOR U9324 ( .A(n2760), .B(n2761), .Z(n2383) );
  AND U9325 ( .A(n2762), .B(n2763), .Z(n2760) );
  AND U9326 ( .A(b[11]), .B(a[109]), .Z(n2759) );
  XOR U9327 ( .A(n2764), .B(n2388), .Z(n2390) );
  XOR U9328 ( .A(n2765), .B(n2766), .Z(n2388) );
  AND U9329 ( .A(n2767), .B(n2768), .Z(n2765) );
  AND U9330 ( .A(b[10]), .B(a[110]), .Z(n2764) );
  XOR U9331 ( .A(n2769), .B(n2393), .Z(n2395) );
  XOR U9332 ( .A(n2770), .B(n2771), .Z(n2393) );
  AND U9333 ( .A(n2772), .B(n2773), .Z(n2770) );
  AND U9334 ( .A(b[9]), .B(a[111]), .Z(n2769) );
  XOR U9335 ( .A(n2774), .B(n2398), .Z(n2400) );
  XOR U9336 ( .A(n2775), .B(n2776), .Z(n2398) );
  AND U9337 ( .A(n2777), .B(n2778), .Z(n2775) );
  AND U9338 ( .A(b[8]), .B(a[112]), .Z(n2774) );
  XOR U9339 ( .A(n2779), .B(n2403), .Z(n2405) );
  XOR U9340 ( .A(n2780), .B(n2781), .Z(n2403) );
  AND U9341 ( .A(n2782), .B(n2783), .Z(n2780) );
  AND U9342 ( .A(b[7]), .B(a[113]), .Z(n2779) );
  XOR U9343 ( .A(n2784), .B(n2408), .Z(n2410) );
  XOR U9344 ( .A(n2785), .B(n2786), .Z(n2408) );
  AND U9345 ( .A(n2787), .B(n2788), .Z(n2785) );
  AND U9346 ( .A(b[6]), .B(a[114]), .Z(n2784) );
  XOR U9347 ( .A(n2789), .B(n2413), .Z(n2415) );
  XOR U9348 ( .A(n2790), .B(n2791), .Z(n2413) );
  AND U9349 ( .A(n2792), .B(n2793), .Z(n2790) );
  AND U9350 ( .A(b[5]), .B(a[115]), .Z(n2789) );
  XOR U9351 ( .A(n2794), .B(n2418), .Z(n2420) );
  XOR U9352 ( .A(n2795), .B(n2796), .Z(n2418) );
  AND U9353 ( .A(n2797), .B(n2798), .Z(n2795) );
  AND U9354 ( .A(b[4]), .B(a[116]), .Z(n2794) );
  XOR U9355 ( .A(n2799), .B(n2800), .Z(n2432) );
  NAND U9356 ( .A(n2801), .B(n2802), .Z(n2800) );
  XOR U9357 ( .A(n2803), .B(n2423), .Z(n2425) );
  XNOR U9358 ( .A(n2804), .B(n2805), .Z(n2423) );
  ANDN U9359 ( .B(n2806), .A(n2807), .Z(n2804) );
  AND U9360 ( .A(b[3]), .B(a[117]), .Z(n2803) );
  XOR U9361 ( .A(n2808), .B(n2809), .Z(swire[119]) );
  XOR U9362 ( .A(n2442), .B(n2810), .Z(n2809) );
  XNOR U9363 ( .A(n2441), .B(n2808), .Z(n2810) );
  NAND U9364 ( .A(a[119]), .B(b[0]), .Z(n2441) );
  XOR U9365 ( .A(n2811), .B(n2812), .Z(n2801) );
  NAND U9366 ( .A(b[1]), .B(a[118]), .Z(n2812) );
  XNOR U9367 ( .A(n2811), .B(n2807), .Z(n2813) );
  XOR U9368 ( .A(n2814), .B(n2805), .Z(n2807) );
  AND U9369 ( .A(b[2]), .B(a[117]), .Z(n2814) );
  IV U9370 ( .A(n2799), .Z(n2811) );
  ANDN U9371 ( .B(n2815), .A(n2816), .Z(n2799) );
  XOR U9372 ( .A(n2805), .B(n2797), .Z(n2817) );
  XNOR U9373 ( .A(n2796), .B(n2792), .Z(n2818) );
  XNOR U9374 ( .A(n2791), .B(n2787), .Z(n2819) );
  XNOR U9375 ( .A(n2786), .B(n2782), .Z(n2820) );
  XNOR U9376 ( .A(n2781), .B(n2777), .Z(n2821) );
  XNOR U9377 ( .A(n2776), .B(n2772), .Z(n2822) );
  XNOR U9378 ( .A(n2771), .B(n2767), .Z(n2823) );
  XNOR U9379 ( .A(n2766), .B(n2762), .Z(n2824) );
  XNOR U9380 ( .A(n2761), .B(n2757), .Z(n2825) );
  XNOR U9381 ( .A(n2756), .B(n2752), .Z(n2826) );
  XNOR U9382 ( .A(n2743), .B(n2742), .Z(n2827) );
  XOR U9383 ( .A(n2828), .B(n2741), .Z(n2742) );
  AND U9384 ( .A(b[13]), .B(a[106]), .Z(n2828) );
  XNOR U9385 ( .A(n2741), .B(n2747), .Z(n2829) );
  XNOR U9386 ( .A(n2746), .B(n2738), .Z(n2830) );
  XNOR U9387 ( .A(n2737), .B(n2733), .Z(n2831) );
  XNOR U9388 ( .A(n2732), .B(n2728), .Z(n2832) );
  XNOR U9389 ( .A(n2727), .B(n2723), .Z(n2833) );
  XNOR U9390 ( .A(n2714), .B(n2713), .Z(n2834) );
  XOR U9391 ( .A(n2835), .B(n2712), .Z(n2713) );
  AND U9392 ( .A(b[19]), .B(a[100]), .Z(n2835) );
  XNOR U9393 ( .A(n2712), .B(n2718), .Z(n2836) );
  XNOR U9394 ( .A(n2717), .B(n2709), .Z(n2837) );
  XNOR U9395 ( .A(n2708), .B(n2704), .Z(n2838) );
  XNOR U9396 ( .A(n2703), .B(n2699), .Z(n2839) );
  XNOR U9397 ( .A(n2698), .B(n2694), .Z(n2840) );
  XNOR U9398 ( .A(n2685), .B(n2684), .Z(n2841) );
  XOR U9399 ( .A(n2842), .B(n2683), .Z(n2684) );
  AND U9400 ( .A(b[25]), .B(a[94]), .Z(n2842) );
  XNOR U9401 ( .A(n2683), .B(n2689), .Z(n2843) );
  XNOR U9402 ( .A(n2688), .B(n2680), .Z(n2844) );
  XNOR U9403 ( .A(n2679), .B(n2675), .Z(n2845) );
  XNOR U9404 ( .A(n2674), .B(n2670), .Z(n2846) );
  XNOR U9405 ( .A(n2669), .B(n2665), .Z(n2847) );
  XNOR U9406 ( .A(n2656), .B(n2655), .Z(n2848) );
  XOR U9407 ( .A(n2849), .B(n2654), .Z(n2655) );
  AND U9408 ( .A(b[31]), .B(a[88]), .Z(n2849) );
  XNOR U9409 ( .A(n2654), .B(n2660), .Z(n2850) );
  XNOR U9410 ( .A(n2659), .B(n2651), .Z(n2851) );
  XNOR U9411 ( .A(n2650), .B(n2646), .Z(n2852) );
  XNOR U9412 ( .A(n2645), .B(n2641), .Z(n2853) );
  XNOR U9413 ( .A(n2640), .B(n2636), .Z(n2854) );
  XNOR U9414 ( .A(n2627), .B(n2626), .Z(n2855) );
  XOR U9415 ( .A(n2856), .B(n2625), .Z(n2626) );
  AND U9416 ( .A(b[37]), .B(a[82]), .Z(n2856) );
  XNOR U9417 ( .A(n2625), .B(n2631), .Z(n2857) );
  XNOR U9418 ( .A(n2630), .B(n2622), .Z(n2858) );
  XNOR U9419 ( .A(n2621), .B(n2617), .Z(n2859) );
  XNOR U9420 ( .A(n2616), .B(n2612), .Z(n2860) );
  XNOR U9421 ( .A(n2611), .B(n2607), .Z(n2861) );
  XNOR U9422 ( .A(n2598), .B(n2597), .Z(n2862) );
  XOR U9423 ( .A(n2863), .B(n2596), .Z(n2597) );
  AND U9424 ( .A(b[43]), .B(a[76]), .Z(n2863) );
  XNOR U9425 ( .A(n2596), .B(n2602), .Z(n2864) );
  XNOR U9426 ( .A(n2601), .B(n2593), .Z(n2865) );
  XNOR U9427 ( .A(n2592), .B(n2588), .Z(n2866) );
  XNOR U9428 ( .A(n2587), .B(n2583), .Z(n2867) );
  XNOR U9429 ( .A(n2582), .B(n2578), .Z(n2868) );
  XNOR U9430 ( .A(n2569), .B(n2568), .Z(n2869) );
  XOR U9431 ( .A(n2870), .B(n2567), .Z(n2568) );
  AND U9432 ( .A(b[49]), .B(a[70]), .Z(n2870) );
  XNOR U9433 ( .A(n2567), .B(n2573), .Z(n2871) );
  XNOR U9434 ( .A(n2572), .B(n2564), .Z(n2872) );
  XNOR U9435 ( .A(n2563), .B(n2559), .Z(n2873) );
  XNOR U9436 ( .A(n2558), .B(n2554), .Z(n2874) );
  XNOR U9437 ( .A(n2553), .B(n2549), .Z(n2875) );
  XNOR U9438 ( .A(n2548), .B(n2544), .Z(n2876) );
  XNOR U9439 ( .A(n2543), .B(n2539), .Z(n2877) );
  XNOR U9440 ( .A(n2538), .B(n2534), .Z(n2878) );
  XNOR U9441 ( .A(n2533), .B(n2529), .Z(n2879) );
  XNOR U9442 ( .A(n2528), .B(n2524), .Z(n2880) );
  XOR U9443 ( .A(n2523), .B(n2520), .Z(n2881) );
  XOR U9444 ( .A(n2882), .B(n2883), .Z(n2520) );
  XOR U9445 ( .A(n2518), .B(n2884), .Z(n2883) );
  XOR U9446 ( .A(n2885), .B(n2886), .Z(n2884) );
  XOR U9447 ( .A(n2887), .B(n2888), .Z(n2886) );
  NAND U9448 ( .A(a[57]), .B(b[62]), .Z(n2888) );
  AND U9449 ( .A(a[56]), .B(b[63]), .Z(n2887) );
  XOR U9450 ( .A(n2889), .B(n2885), .Z(n2882) );
  XOR U9451 ( .A(n2890), .B(n2891), .Z(n2885) );
  ANDN U9452 ( .B(n2892), .A(n2893), .Z(n2890) );
  AND U9453 ( .A(a[58]), .B(b[61]), .Z(n2889) );
  XOR U9454 ( .A(n2894), .B(n2518), .Z(n2519) );
  XOR U9455 ( .A(n2895), .B(n2896), .Z(n2518) );
  AND U9456 ( .A(n2897), .B(n2898), .Z(n2895) );
  AND U9457 ( .A(a[59]), .B(b[60]), .Z(n2894) );
  XOR U9458 ( .A(n2899), .B(n2523), .Z(n2525) );
  XOR U9459 ( .A(n2900), .B(n2901), .Z(n2523) );
  AND U9460 ( .A(n2902), .B(n2903), .Z(n2900) );
  AND U9461 ( .A(b[59]), .B(a[60]), .Z(n2899) );
  XOR U9462 ( .A(n2904), .B(n2528), .Z(n2530) );
  XOR U9463 ( .A(n2905), .B(n2906), .Z(n2528) );
  AND U9464 ( .A(n2907), .B(n2908), .Z(n2905) );
  AND U9465 ( .A(b[58]), .B(a[61]), .Z(n2904) );
  XOR U9466 ( .A(n2909), .B(n2533), .Z(n2535) );
  XOR U9467 ( .A(n2910), .B(n2911), .Z(n2533) );
  AND U9468 ( .A(n2912), .B(n2913), .Z(n2910) );
  AND U9469 ( .A(b[57]), .B(a[62]), .Z(n2909) );
  XOR U9470 ( .A(n2914), .B(n2538), .Z(n2540) );
  XOR U9471 ( .A(n2915), .B(n2916), .Z(n2538) );
  AND U9472 ( .A(n2917), .B(n2918), .Z(n2915) );
  AND U9473 ( .A(b[56]), .B(a[63]), .Z(n2914) );
  XOR U9474 ( .A(n2919), .B(n2543), .Z(n2545) );
  XOR U9475 ( .A(n2920), .B(n2921), .Z(n2543) );
  AND U9476 ( .A(n2922), .B(n2923), .Z(n2920) );
  AND U9477 ( .A(b[55]), .B(a[64]), .Z(n2919) );
  XOR U9478 ( .A(n2924), .B(n2548), .Z(n2550) );
  XOR U9479 ( .A(n2925), .B(n2926), .Z(n2548) );
  AND U9480 ( .A(n2927), .B(n2928), .Z(n2925) );
  AND U9481 ( .A(b[54]), .B(a[65]), .Z(n2924) );
  XOR U9482 ( .A(n2929), .B(n2553), .Z(n2555) );
  XOR U9483 ( .A(n2930), .B(n2931), .Z(n2553) );
  AND U9484 ( .A(n2932), .B(n2933), .Z(n2930) );
  AND U9485 ( .A(b[53]), .B(a[66]), .Z(n2929) );
  XOR U9486 ( .A(n2934), .B(n2558), .Z(n2560) );
  XOR U9487 ( .A(n2935), .B(n2936), .Z(n2558) );
  AND U9488 ( .A(n2937), .B(n2938), .Z(n2935) );
  AND U9489 ( .A(b[52]), .B(a[67]), .Z(n2934) );
  XOR U9490 ( .A(n2939), .B(n2563), .Z(n2565) );
  XOR U9491 ( .A(n2940), .B(n2941), .Z(n2563) );
  AND U9492 ( .A(n2942), .B(n2943), .Z(n2940) );
  AND U9493 ( .A(b[51]), .B(a[68]), .Z(n2939) );
  XOR U9494 ( .A(n2944), .B(n2945), .Z(n2567) );
  AND U9495 ( .A(n2946), .B(n2947), .Z(n2944) );
  XOR U9496 ( .A(n2948), .B(n2572), .Z(n2574) );
  XOR U9497 ( .A(n2949), .B(n2950), .Z(n2572) );
  AND U9498 ( .A(n2951), .B(n2952), .Z(n2949) );
  AND U9499 ( .A(b[50]), .B(a[69]), .Z(n2948) );
  XOR U9500 ( .A(n2953), .B(n2577), .Z(n2579) );
  XOR U9501 ( .A(n2954), .B(n2955), .Z(n2577) );
  AND U9502 ( .A(n2956), .B(n2957), .Z(n2954) );
  AND U9503 ( .A(b[48]), .B(a[71]), .Z(n2953) );
  XOR U9504 ( .A(n2958), .B(n2582), .Z(n2584) );
  XOR U9505 ( .A(n2959), .B(n2960), .Z(n2582) );
  AND U9506 ( .A(n2961), .B(n2962), .Z(n2959) );
  AND U9507 ( .A(b[47]), .B(a[72]), .Z(n2958) );
  XOR U9508 ( .A(n2963), .B(n2587), .Z(n2589) );
  XOR U9509 ( .A(n2964), .B(n2965), .Z(n2587) );
  AND U9510 ( .A(n2966), .B(n2967), .Z(n2964) );
  AND U9511 ( .A(b[46]), .B(a[73]), .Z(n2963) );
  XOR U9512 ( .A(n2968), .B(n2592), .Z(n2594) );
  XOR U9513 ( .A(n2969), .B(n2970), .Z(n2592) );
  AND U9514 ( .A(n2971), .B(n2972), .Z(n2969) );
  AND U9515 ( .A(b[45]), .B(a[74]), .Z(n2968) );
  XOR U9516 ( .A(n2973), .B(n2974), .Z(n2596) );
  AND U9517 ( .A(n2975), .B(n2976), .Z(n2973) );
  XOR U9518 ( .A(n2977), .B(n2601), .Z(n2603) );
  XOR U9519 ( .A(n2978), .B(n2979), .Z(n2601) );
  AND U9520 ( .A(n2980), .B(n2981), .Z(n2978) );
  AND U9521 ( .A(b[44]), .B(a[75]), .Z(n2977) );
  XOR U9522 ( .A(n2982), .B(n2606), .Z(n2608) );
  XOR U9523 ( .A(n2983), .B(n2984), .Z(n2606) );
  AND U9524 ( .A(n2985), .B(n2986), .Z(n2983) );
  AND U9525 ( .A(b[42]), .B(a[77]), .Z(n2982) );
  XOR U9526 ( .A(n2987), .B(n2611), .Z(n2613) );
  XOR U9527 ( .A(n2988), .B(n2989), .Z(n2611) );
  AND U9528 ( .A(n2990), .B(n2991), .Z(n2988) );
  AND U9529 ( .A(b[41]), .B(a[78]), .Z(n2987) );
  XOR U9530 ( .A(n2992), .B(n2616), .Z(n2618) );
  XOR U9531 ( .A(n2993), .B(n2994), .Z(n2616) );
  AND U9532 ( .A(n2995), .B(n2996), .Z(n2993) );
  AND U9533 ( .A(b[40]), .B(a[79]), .Z(n2992) );
  XOR U9534 ( .A(n2997), .B(n2621), .Z(n2623) );
  XOR U9535 ( .A(n2998), .B(n2999), .Z(n2621) );
  AND U9536 ( .A(n3000), .B(n3001), .Z(n2998) );
  AND U9537 ( .A(b[39]), .B(a[80]), .Z(n2997) );
  XOR U9538 ( .A(n3002), .B(n3003), .Z(n2625) );
  AND U9539 ( .A(n3004), .B(n3005), .Z(n3002) );
  XOR U9540 ( .A(n3006), .B(n2630), .Z(n2632) );
  XOR U9541 ( .A(n3007), .B(n3008), .Z(n2630) );
  AND U9542 ( .A(n3009), .B(n3010), .Z(n3007) );
  AND U9543 ( .A(b[38]), .B(a[81]), .Z(n3006) );
  XOR U9544 ( .A(n3011), .B(n2635), .Z(n2637) );
  XOR U9545 ( .A(n3012), .B(n3013), .Z(n2635) );
  AND U9546 ( .A(n3014), .B(n3015), .Z(n3012) );
  AND U9547 ( .A(b[36]), .B(a[83]), .Z(n3011) );
  XOR U9548 ( .A(n3016), .B(n2640), .Z(n2642) );
  XOR U9549 ( .A(n3017), .B(n3018), .Z(n2640) );
  AND U9550 ( .A(n3019), .B(n3020), .Z(n3017) );
  AND U9551 ( .A(b[35]), .B(a[84]), .Z(n3016) );
  XOR U9552 ( .A(n3021), .B(n2645), .Z(n2647) );
  XOR U9553 ( .A(n3022), .B(n3023), .Z(n2645) );
  AND U9554 ( .A(n3024), .B(n3025), .Z(n3022) );
  AND U9555 ( .A(b[34]), .B(a[85]), .Z(n3021) );
  XOR U9556 ( .A(n3026), .B(n2650), .Z(n2652) );
  XOR U9557 ( .A(n3027), .B(n3028), .Z(n2650) );
  AND U9558 ( .A(n3029), .B(n3030), .Z(n3027) );
  AND U9559 ( .A(b[33]), .B(a[86]), .Z(n3026) );
  XOR U9560 ( .A(n3031), .B(n3032), .Z(n2654) );
  AND U9561 ( .A(n3033), .B(n3034), .Z(n3031) );
  XOR U9562 ( .A(n3035), .B(n2659), .Z(n2661) );
  XOR U9563 ( .A(n3036), .B(n3037), .Z(n2659) );
  AND U9564 ( .A(n3038), .B(n3039), .Z(n3036) );
  AND U9565 ( .A(b[32]), .B(a[87]), .Z(n3035) );
  XOR U9566 ( .A(n3040), .B(n2664), .Z(n2666) );
  XOR U9567 ( .A(n3041), .B(n3042), .Z(n2664) );
  AND U9568 ( .A(n3043), .B(n3044), .Z(n3041) );
  AND U9569 ( .A(b[30]), .B(a[89]), .Z(n3040) );
  XOR U9570 ( .A(n3045), .B(n2669), .Z(n2671) );
  XOR U9571 ( .A(n3046), .B(n3047), .Z(n2669) );
  AND U9572 ( .A(n3048), .B(n3049), .Z(n3046) );
  AND U9573 ( .A(b[29]), .B(a[90]), .Z(n3045) );
  XOR U9574 ( .A(n3050), .B(n2674), .Z(n2676) );
  XOR U9575 ( .A(n3051), .B(n3052), .Z(n2674) );
  AND U9576 ( .A(n3053), .B(n3054), .Z(n3051) );
  AND U9577 ( .A(b[28]), .B(a[91]), .Z(n3050) );
  XOR U9578 ( .A(n3055), .B(n2679), .Z(n2681) );
  XOR U9579 ( .A(n3056), .B(n3057), .Z(n2679) );
  AND U9580 ( .A(n3058), .B(n3059), .Z(n3056) );
  AND U9581 ( .A(b[27]), .B(a[92]), .Z(n3055) );
  XOR U9582 ( .A(n3060), .B(n3061), .Z(n2683) );
  AND U9583 ( .A(n3062), .B(n3063), .Z(n3060) );
  XOR U9584 ( .A(n3064), .B(n2688), .Z(n2690) );
  XOR U9585 ( .A(n3065), .B(n3066), .Z(n2688) );
  AND U9586 ( .A(n3067), .B(n3068), .Z(n3065) );
  AND U9587 ( .A(b[26]), .B(a[93]), .Z(n3064) );
  XOR U9588 ( .A(n3069), .B(n2693), .Z(n2695) );
  XOR U9589 ( .A(n3070), .B(n3071), .Z(n2693) );
  AND U9590 ( .A(n3072), .B(n3073), .Z(n3070) );
  AND U9591 ( .A(b[24]), .B(a[95]), .Z(n3069) );
  XOR U9592 ( .A(n3074), .B(n2698), .Z(n2700) );
  XOR U9593 ( .A(n3075), .B(n3076), .Z(n2698) );
  AND U9594 ( .A(n3077), .B(n3078), .Z(n3075) );
  AND U9595 ( .A(b[23]), .B(a[96]), .Z(n3074) );
  XOR U9596 ( .A(n3079), .B(n2703), .Z(n2705) );
  XOR U9597 ( .A(n3080), .B(n3081), .Z(n2703) );
  AND U9598 ( .A(n3082), .B(n3083), .Z(n3080) );
  AND U9599 ( .A(b[22]), .B(a[97]), .Z(n3079) );
  XOR U9600 ( .A(n3084), .B(n2708), .Z(n2710) );
  XOR U9601 ( .A(n3085), .B(n3086), .Z(n2708) );
  AND U9602 ( .A(n3087), .B(n3088), .Z(n3085) );
  AND U9603 ( .A(b[21]), .B(a[98]), .Z(n3084) );
  XOR U9604 ( .A(n3089), .B(n3090), .Z(n2712) );
  AND U9605 ( .A(n3091), .B(n3092), .Z(n3089) );
  XOR U9606 ( .A(n3093), .B(n2717), .Z(n2719) );
  XOR U9607 ( .A(n3094), .B(n3095), .Z(n2717) );
  AND U9608 ( .A(n3096), .B(n3097), .Z(n3094) );
  AND U9609 ( .A(b[20]), .B(a[99]), .Z(n3093) );
  XOR U9610 ( .A(n3098), .B(n2722), .Z(n2724) );
  XOR U9611 ( .A(n3099), .B(n3100), .Z(n2722) );
  AND U9612 ( .A(n3101), .B(n3102), .Z(n3099) );
  AND U9613 ( .A(b[18]), .B(a[101]), .Z(n3098) );
  XOR U9614 ( .A(n3103), .B(n2727), .Z(n2729) );
  XOR U9615 ( .A(n3104), .B(n3105), .Z(n2727) );
  AND U9616 ( .A(n3106), .B(n3107), .Z(n3104) );
  AND U9617 ( .A(b[17]), .B(a[102]), .Z(n3103) );
  XOR U9618 ( .A(n3108), .B(n2732), .Z(n2734) );
  XOR U9619 ( .A(n3109), .B(n3110), .Z(n2732) );
  AND U9620 ( .A(n3111), .B(n3112), .Z(n3109) );
  AND U9621 ( .A(b[16]), .B(a[103]), .Z(n3108) );
  XOR U9622 ( .A(n3113), .B(n2737), .Z(n2739) );
  XOR U9623 ( .A(n3114), .B(n3115), .Z(n2737) );
  AND U9624 ( .A(n3116), .B(n3117), .Z(n3114) );
  AND U9625 ( .A(b[15]), .B(a[104]), .Z(n3113) );
  XOR U9626 ( .A(n3118), .B(n3119), .Z(n2741) );
  AND U9627 ( .A(n3120), .B(n3121), .Z(n3118) );
  XOR U9628 ( .A(n3122), .B(n2746), .Z(n2748) );
  XOR U9629 ( .A(n3123), .B(n3124), .Z(n2746) );
  AND U9630 ( .A(n3125), .B(n3126), .Z(n3123) );
  AND U9631 ( .A(b[14]), .B(a[105]), .Z(n3122) );
  XOR U9632 ( .A(n3127), .B(n2751), .Z(n2753) );
  XOR U9633 ( .A(n3128), .B(n3129), .Z(n2751) );
  AND U9634 ( .A(n3130), .B(n3131), .Z(n3128) );
  AND U9635 ( .A(b[12]), .B(a[107]), .Z(n3127) );
  XOR U9636 ( .A(n3132), .B(n2756), .Z(n2758) );
  XOR U9637 ( .A(n3133), .B(n3134), .Z(n2756) );
  AND U9638 ( .A(n3135), .B(n3136), .Z(n3133) );
  AND U9639 ( .A(b[11]), .B(a[108]), .Z(n3132) );
  XOR U9640 ( .A(n3137), .B(n2761), .Z(n2763) );
  XOR U9641 ( .A(n3138), .B(n3139), .Z(n2761) );
  AND U9642 ( .A(n3140), .B(n3141), .Z(n3138) );
  AND U9643 ( .A(b[10]), .B(a[109]), .Z(n3137) );
  XOR U9644 ( .A(n3142), .B(n2766), .Z(n2768) );
  XOR U9645 ( .A(n3143), .B(n3144), .Z(n2766) );
  AND U9646 ( .A(n3145), .B(n3146), .Z(n3143) );
  AND U9647 ( .A(b[9]), .B(a[110]), .Z(n3142) );
  XOR U9648 ( .A(n3147), .B(n2771), .Z(n2773) );
  XOR U9649 ( .A(n3148), .B(n3149), .Z(n2771) );
  AND U9650 ( .A(n3150), .B(n3151), .Z(n3148) );
  AND U9651 ( .A(b[8]), .B(a[111]), .Z(n3147) );
  XOR U9652 ( .A(n3152), .B(n2776), .Z(n2778) );
  XOR U9653 ( .A(n3153), .B(n3154), .Z(n2776) );
  AND U9654 ( .A(n3155), .B(n3156), .Z(n3153) );
  AND U9655 ( .A(b[7]), .B(a[112]), .Z(n3152) );
  XOR U9656 ( .A(n3157), .B(n2781), .Z(n2783) );
  XOR U9657 ( .A(n3158), .B(n3159), .Z(n2781) );
  AND U9658 ( .A(n3160), .B(n3161), .Z(n3158) );
  AND U9659 ( .A(b[6]), .B(a[113]), .Z(n3157) );
  XOR U9660 ( .A(n3162), .B(n2786), .Z(n2788) );
  XOR U9661 ( .A(n3163), .B(n3164), .Z(n2786) );
  AND U9662 ( .A(n3165), .B(n3166), .Z(n3163) );
  AND U9663 ( .A(b[5]), .B(a[114]), .Z(n3162) );
  XOR U9664 ( .A(n3167), .B(n2791), .Z(n2793) );
  XOR U9665 ( .A(n3168), .B(n3169), .Z(n2791) );
  AND U9666 ( .A(n3170), .B(n3171), .Z(n3168) );
  AND U9667 ( .A(b[4]), .B(a[115]), .Z(n3167) );
  XOR U9668 ( .A(n3172), .B(n3173), .Z(n2805) );
  NANDN U9669 ( .A(n3174), .B(n3175), .Z(n3173) );
  XOR U9670 ( .A(n3176), .B(n2796), .Z(n2798) );
  XNOR U9671 ( .A(n3177), .B(n3178), .Z(n2796) );
  AND U9672 ( .A(n3179), .B(n3180), .Z(n3177) );
  AND U9673 ( .A(b[3]), .B(a[116]), .Z(n3176) );
  XOR U9674 ( .A(n3181), .B(n3182), .Z(swire[118]) );
  XOR U9675 ( .A(n2815), .B(n3183), .Z(n3182) );
  XNOR U9676 ( .A(n2816), .B(n3181), .Z(n3183) );
  NAND U9677 ( .A(a[118]), .B(b[0]), .Z(n2816) );
  XNOR U9678 ( .A(n3175), .B(n3174), .Z(n2815) );
  XOR U9679 ( .A(n3172), .B(n3184), .Z(n3174) );
  NAND U9680 ( .A(b[1]), .B(a[117]), .Z(n3184) );
  XNOR U9681 ( .A(n3180), .B(n3185), .Z(n3175) );
  XNOR U9682 ( .A(n3172), .B(n3179), .Z(n3185) );
  XNOR U9683 ( .A(n3186), .B(n3178), .Z(n3179) );
  AND U9684 ( .A(b[2]), .B(a[116]), .Z(n3186) );
  ANDN U9685 ( .B(n3187), .A(n3188), .Z(n3172) );
  XOR U9686 ( .A(n3178), .B(n3170), .Z(n3189) );
  XNOR U9687 ( .A(n3169), .B(n3165), .Z(n3190) );
  XNOR U9688 ( .A(n3164), .B(n3160), .Z(n3191) );
  XNOR U9689 ( .A(n3159), .B(n3155), .Z(n3192) );
  XNOR U9690 ( .A(n3154), .B(n3150), .Z(n3193) );
  XNOR U9691 ( .A(n3149), .B(n3145), .Z(n3194) );
  XNOR U9692 ( .A(n3144), .B(n3140), .Z(n3195) );
  XNOR U9693 ( .A(n3139), .B(n3135), .Z(n3196) );
  XNOR U9694 ( .A(n3134), .B(n3130), .Z(n3197) );
  XNOR U9695 ( .A(n3121), .B(n3120), .Z(n3198) );
  XOR U9696 ( .A(n3199), .B(n3119), .Z(n3120) );
  AND U9697 ( .A(b[12]), .B(a[106]), .Z(n3199) );
  XNOR U9698 ( .A(n3119), .B(n3125), .Z(n3200) );
  XNOR U9699 ( .A(n3124), .B(n3116), .Z(n3201) );
  XNOR U9700 ( .A(n3115), .B(n3111), .Z(n3202) );
  XNOR U9701 ( .A(n3110), .B(n3106), .Z(n3203) );
  XNOR U9702 ( .A(n3105), .B(n3101), .Z(n3204) );
  XNOR U9703 ( .A(n3092), .B(n3091), .Z(n3205) );
  XOR U9704 ( .A(n3206), .B(n3090), .Z(n3091) );
  AND U9705 ( .A(b[18]), .B(a[100]), .Z(n3206) );
  XNOR U9706 ( .A(n3090), .B(n3096), .Z(n3207) );
  XNOR U9707 ( .A(n3095), .B(n3087), .Z(n3208) );
  XNOR U9708 ( .A(n3086), .B(n3082), .Z(n3209) );
  XNOR U9709 ( .A(n3081), .B(n3077), .Z(n3210) );
  XNOR U9710 ( .A(n3076), .B(n3072), .Z(n3211) );
  XNOR U9711 ( .A(n3063), .B(n3062), .Z(n3212) );
  XOR U9712 ( .A(n3213), .B(n3061), .Z(n3062) );
  AND U9713 ( .A(b[24]), .B(a[94]), .Z(n3213) );
  XNOR U9714 ( .A(n3061), .B(n3067), .Z(n3214) );
  XNOR U9715 ( .A(n3066), .B(n3058), .Z(n3215) );
  XNOR U9716 ( .A(n3057), .B(n3053), .Z(n3216) );
  XNOR U9717 ( .A(n3052), .B(n3048), .Z(n3217) );
  XNOR U9718 ( .A(n3047), .B(n3043), .Z(n3218) );
  XNOR U9719 ( .A(n3034), .B(n3033), .Z(n3219) );
  XOR U9720 ( .A(n3220), .B(n3032), .Z(n3033) );
  AND U9721 ( .A(b[30]), .B(a[88]), .Z(n3220) );
  XNOR U9722 ( .A(n3032), .B(n3038), .Z(n3221) );
  XNOR U9723 ( .A(n3037), .B(n3029), .Z(n3222) );
  XNOR U9724 ( .A(n3028), .B(n3024), .Z(n3223) );
  XNOR U9725 ( .A(n3023), .B(n3019), .Z(n3224) );
  XNOR U9726 ( .A(n3018), .B(n3014), .Z(n3225) );
  XNOR U9727 ( .A(n3005), .B(n3004), .Z(n3226) );
  XOR U9728 ( .A(n3227), .B(n3003), .Z(n3004) );
  AND U9729 ( .A(b[36]), .B(a[82]), .Z(n3227) );
  XNOR U9730 ( .A(n3003), .B(n3009), .Z(n3228) );
  XNOR U9731 ( .A(n3008), .B(n3000), .Z(n3229) );
  XNOR U9732 ( .A(n2999), .B(n2995), .Z(n3230) );
  XNOR U9733 ( .A(n2994), .B(n2990), .Z(n3231) );
  XNOR U9734 ( .A(n2989), .B(n2985), .Z(n3232) );
  XNOR U9735 ( .A(n2976), .B(n2975), .Z(n3233) );
  XOR U9736 ( .A(n3234), .B(n2974), .Z(n2975) );
  AND U9737 ( .A(b[42]), .B(a[76]), .Z(n3234) );
  XNOR U9738 ( .A(n2974), .B(n2980), .Z(n3235) );
  XNOR U9739 ( .A(n2979), .B(n2971), .Z(n3236) );
  XNOR U9740 ( .A(n2970), .B(n2966), .Z(n3237) );
  XNOR U9741 ( .A(n2965), .B(n2961), .Z(n3238) );
  XNOR U9742 ( .A(n2960), .B(n2956), .Z(n3239) );
  XNOR U9743 ( .A(n2947), .B(n2946), .Z(n3240) );
  XOR U9744 ( .A(n3241), .B(n2945), .Z(n2946) );
  AND U9745 ( .A(b[48]), .B(a[70]), .Z(n3241) );
  XNOR U9746 ( .A(n2945), .B(n2951), .Z(n3242) );
  XNOR U9747 ( .A(n2950), .B(n2942), .Z(n3243) );
  XNOR U9748 ( .A(n2941), .B(n2937), .Z(n3244) );
  XNOR U9749 ( .A(n2936), .B(n2932), .Z(n3245) );
  XNOR U9750 ( .A(n2931), .B(n2927), .Z(n3246) );
  XNOR U9751 ( .A(n2926), .B(n2922), .Z(n3247) );
  XNOR U9752 ( .A(n2921), .B(n2917), .Z(n3248) );
  XNOR U9753 ( .A(n2916), .B(n2912), .Z(n3249) );
  XNOR U9754 ( .A(n2911), .B(n2907), .Z(n3250) );
  XNOR U9755 ( .A(n2906), .B(n2902), .Z(n3251) );
  XNOR U9756 ( .A(n2901), .B(n2897), .Z(n3252) );
  XOR U9757 ( .A(n2896), .B(n2893), .Z(n3253) );
  XOR U9758 ( .A(n3254), .B(n3255), .Z(n2893) );
  XOR U9759 ( .A(n2891), .B(n3256), .Z(n3255) );
  XOR U9760 ( .A(n3257), .B(n3258), .Z(n3256) );
  XOR U9761 ( .A(n3259), .B(n3260), .Z(n3258) );
  NAND U9762 ( .A(a[56]), .B(b[62]), .Z(n3260) );
  AND U9763 ( .A(a[55]), .B(b[63]), .Z(n3259) );
  XOR U9764 ( .A(n3261), .B(n3257), .Z(n3254) );
  XOR U9765 ( .A(n3262), .B(n3263), .Z(n3257) );
  ANDN U9766 ( .B(n3264), .A(n3265), .Z(n3262) );
  AND U9767 ( .A(a[57]), .B(b[61]), .Z(n3261) );
  XOR U9768 ( .A(n3266), .B(n2891), .Z(n2892) );
  XOR U9769 ( .A(n3267), .B(n3268), .Z(n2891) );
  AND U9770 ( .A(n3269), .B(n3270), .Z(n3267) );
  AND U9771 ( .A(a[58]), .B(b[60]), .Z(n3266) );
  XOR U9772 ( .A(n3271), .B(n2896), .Z(n2898) );
  XOR U9773 ( .A(n3272), .B(n3273), .Z(n2896) );
  AND U9774 ( .A(n3274), .B(n3275), .Z(n3272) );
  AND U9775 ( .A(a[59]), .B(b[59]), .Z(n3271) );
  XOR U9776 ( .A(n3276), .B(n2901), .Z(n2903) );
  XOR U9777 ( .A(n3277), .B(n3278), .Z(n2901) );
  AND U9778 ( .A(n3279), .B(n3280), .Z(n3277) );
  AND U9779 ( .A(b[58]), .B(a[60]), .Z(n3276) );
  XOR U9780 ( .A(n3281), .B(n2906), .Z(n2908) );
  XOR U9781 ( .A(n3282), .B(n3283), .Z(n2906) );
  AND U9782 ( .A(n3284), .B(n3285), .Z(n3282) );
  AND U9783 ( .A(b[57]), .B(a[61]), .Z(n3281) );
  XOR U9784 ( .A(n3286), .B(n2911), .Z(n2913) );
  XOR U9785 ( .A(n3287), .B(n3288), .Z(n2911) );
  AND U9786 ( .A(n3289), .B(n3290), .Z(n3287) );
  AND U9787 ( .A(b[56]), .B(a[62]), .Z(n3286) );
  XOR U9788 ( .A(n3291), .B(n2916), .Z(n2918) );
  XOR U9789 ( .A(n3292), .B(n3293), .Z(n2916) );
  AND U9790 ( .A(n3294), .B(n3295), .Z(n3292) );
  AND U9791 ( .A(b[55]), .B(a[63]), .Z(n3291) );
  XOR U9792 ( .A(n3296), .B(n2921), .Z(n2923) );
  XOR U9793 ( .A(n3297), .B(n3298), .Z(n2921) );
  AND U9794 ( .A(n3299), .B(n3300), .Z(n3297) );
  AND U9795 ( .A(b[54]), .B(a[64]), .Z(n3296) );
  XOR U9796 ( .A(n3301), .B(n2926), .Z(n2928) );
  XOR U9797 ( .A(n3302), .B(n3303), .Z(n2926) );
  AND U9798 ( .A(n3304), .B(n3305), .Z(n3302) );
  AND U9799 ( .A(b[53]), .B(a[65]), .Z(n3301) );
  XOR U9800 ( .A(n3306), .B(n2931), .Z(n2933) );
  XOR U9801 ( .A(n3307), .B(n3308), .Z(n2931) );
  AND U9802 ( .A(n3309), .B(n3310), .Z(n3307) );
  AND U9803 ( .A(b[52]), .B(a[66]), .Z(n3306) );
  XOR U9804 ( .A(n3311), .B(n2936), .Z(n2938) );
  XOR U9805 ( .A(n3312), .B(n3313), .Z(n2936) );
  AND U9806 ( .A(n3314), .B(n3315), .Z(n3312) );
  AND U9807 ( .A(b[51]), .B(a[67]), .Z(n3311) );
  XOR U9808 ( .A(n3316), .B(n2941), .Z(n2943) );
  XOR U9809 ( .A(n3317), .B(n3318), .Z(n2941) );
  AND U9810 ( .A(n3319), .B(n3320), .Z(n3317) );
  AND U9811 ( .A(b[50]), .B(a[68]), .Z(n3316) );
  XOR U9812 ( .A(n3321), .B(n3322), .Z(n2945) );
  AND U9813 ( .A(n3323), .B(n3324), .Z(n3321) );
  XOR U9814 ( .A(n3325), .B(n2950), .Z(n2952) );
  XOR U9815 ( .A(n3326), .B(n3327), .Z(n2950) );
  AND U9816 ( .A(n3328), .B(n3329), .Z(n3326) );
  AND U9817 ( .A(b[49]), .B(a[69]), .Z(n3325) );
  XOR U9818 ( .A(n3330), .B(n2955), .Z(n2957) );
  XOR U9819 ( .A(n3331), .B(n3332), .Z(n2955) );
  AND U9820 ( .A(n3333), .B(n3334), .Z(n3331) );
  AND U9821 ( .A(b[47]), .B(a[71]), .Z(n3330) );
  XOR U9822 ( .A(n3335), .B(n2960), .Z(n2962) );
  XOR U9823 ( .A(n3336), .B(n3337), .Z(n2960) );
  AND U9824 ( .A(n3338), .B(n3339), .Z(n3336) );
  AND U9825 ( .A(b[46]), .B(a[72]), .Z(n3335) );
  XOR U9826 ( .A(n3340), .B(n2965), .Z(n2967) );
  XOR U9827 ( .A(n3341), .B(n3342), .Z(n2965) );
  AND U9828 ( .A(n3343), .B(n3344), .Z(n3341) );
  AND U9829 ( .A(b[45]), .B(a[73]), .Z(n3340) );
  XOR U9830 ( .A(n3345), .B(n2970), .Z(n2972) );
  XOR U9831 ( .A(n3346), .B(n3347), .Z(n2970) );
  AND U9832 ( .A(n3348), .B(n3349), .Z(n3346) );
  AND U9833 ( .A(b[44]), .B(a[74]), .Z(n3345) );
  XOR U9834 ( .A(n3350), .B(n3351), .Z(n2974) );
  AND U9835 ( .A(n3352), .B(n3353), .Z(n3350) );
  XOR U9836 ( .A(n3354), .B(n2979), .Z(n2981) );
  XOR U9837 ( .A(n3355), .B(n3356), .Z(n2979) );
  AND U9838 ( .A(n3357), .B(n3358), .Z(n3355) );
  AND U9839 ( .A(b[43]), .B(a[75]), .Z(n3354) );
  XOR U9840 ( .A(n3359), .B(n2984), .Z(n2986) );
  XOR U9841 ( .A(n3360), .B(n3361), .Z(n2984) );
  AND U9842 ( .A(n3362), .B(n3363), .Z(n3360) );
  AND U9843 ( .A(b[41]), .B(a[77]), .Z(n3359) );
  XOR U9844 ( .A(n3364), .B(n2989), .Z(n2991) );
  XOR U9845 ( .A(n3365), .B(n3366), .Z(n2989) );
  AND U9846 ( .A(n3367), .B(n3368), .Z(n3365) );
  AND U9847 ( .A(b[40]), .B(a[78]), .Z(n3364) );
  XOR U9848 ( .A(n3369), .B(n2994), .Z(n2996) );
  XOR U9849 ( .A(n3370), .B(n3371), .Z(n2994) );
  AND U9850 ( .A(n3372), .B(n3373), .Z(n3370) );
  AND U9851 ( .A(b[39]), .B(a[79]), .Z(n3369) );
  XOR U9852 ( .A(n3374), .B(n2999), .Z(n3001) );
  XOR U9853 ( .A(n3375), .B(n3376), .Z(n2999) );
  AND U9854 ( .A(n3377), .B(n3378), .Z(n3375) );
  AND U9855 ( .A(b[38]), .B(a[80]), .Z(n3374) );
  XOR U9856 ( .A(n3379), .B(n3380), .Z(n3003) );
  AND U9857 ( .A(n3381), .B(n3382), .Z(n3379) );
  XOR U9858 ( .A(n3383), .B(n3008), .Z(n3010) );
  XOR U9859 ( .A(n3384), .B(n3385), .Z(n3008) );
  AND U9860 ( .A(n3386), .B(n3387), .Z(n3384) );
  AND U9861 ( .A(b[37]), .B(a[81]), .Z(n3383) );
  XOR U9862 ( .A(n3388), .B(n3013), .Z(n3015) );
  XOR U9863 ( .A(n3389), .B(n3390), .Z(n3013) );
  AND U9864 ( .A(n3391), .B(n3392), .Z(n3389) );
  AND U9865 ( .A(b[35]), .B(a[83]), .Z(n3388) );
  XOR U9866 ( .A(n3393), .B(n3018), .Z(n3020) );
  XOR U9867 ( .A(n3394), .B(n3395), .Z(n3018) );
  AND U9868 ( .A(n3396), .B(n3397), .Z(n3394) );
  AND U9869 ( .A(b[34]), .B(a[84]), .Z(n3393) );
  XOR U9870 ( .A(n3398), .B(n3023), .Z(n3025) );
  XOR U9871 ( .A(n3399), .B(n3400), .Z(n3023) );
  AND U9872 ( .A(n3401), .B(n3402), .Z(n3399) );
  AND U9873 ( .A(b[33]), .B(a[85]), .Z(n3398) );
  XOR U9874 ( .A(n3403), .B(n3028), .Z(n3030) );
  XOR U9875 ( .A(n3404), .B(n3405), .Z(n3028) );
  AND U9876 ( .A(n3406), .B(n3407), .Z(n3404) );
  AND U9877 ( .A(b[32]), .B(a[86]), .Z(n3403) );
  XOR U9878 ( .A(n3408), .B(n3409), .Z(n3032) );
  AND U9879 ( .A(n3410), .B(n3411), .Z(n3408) );
  XOR U9880 ( .A(n3412), .B(n3037), .Z(n3039) );
  XOR U9881 ( .A(n3413), .B(n3414), .Z(n3037) );
  AND U9882 ( .A(n3415), .B(n3416), .Z(n3413) );
  AND U9883 ( .A(b[31]), .B(a[87]), .Z(n3412) );
  XOR U9884 ( .A(n3417), .B(n3042), .Z(n3044) );
  XOR U9885 ( .A(n3418), .B(n3419), .Z(n3042) );
  AND U9886 ( .A(n3420), .B(n3421), .Z(n3418) );
  AND U9887 ( .A(b[29]), .B(a[89]), .Z(n3417) );
  XOR U9888 ( .A(n3422), .B(n3047), .Z(n3049) );
  XOR U9889 ( .A(n3423), .B(n3424), .Z(n3047) );
  AND U9890 ( .A(n3425), .B(n3426), .Z(n3423) );
  AND U9891 ( .A(b[28]), .B(a[90]), .Z(n3422) );
  XOR U9892 ( .A(n3427), .B(n3052), .Z(n3054) );
  XOR U9893 ( .A(n3428), .B(n3429), .Z(n3052) );
  AND U9894 ( .A(n3430), .B(n3431), .Z(n3428) );
  AND U9895 ( .A(b[27]), .B(a[91]), .Z(n3427) );
  XOR U9896 ( .A(n3432), .B(n3057), .Z(n3059) );
  XOR U9897 ( .A(n3433), .B(n3434), .Z(n3057) );
  AND U9898 ( .A(n3435), .B(n3436), .Z(n3433) );
  AND U9899 ( .A(b[26]), .B(a[92]), .Z(n3432) );
  XOR U9900 ( .A(n3437), .B(n3438), .Z(n3061) );
  AND U9901 ( .A(n3439), .B(n3440), .Z(n3437) );
  XOR U9902 ( .A(n3441), .B(n3066), .Z(n3068) );
  XOR U9903 ( .A(n3442), .B(n3443), .Z(n3066) );
  AND U9904 ( .A(n3444), .B(n3445), .Z(n3442) );
  AND U9905 ( .A(b[25]), .B(a[93]), .Z(n3441) );
  XOR U9906 ( .A(n3446), .B(n3071), .Z(n3073) );
  XOR U9907 ( .A(n3447), .B(n3448), .Z(n3071) );
  AND U9908 ( .A(n3449), .B(n3450), .Z(n3447) );
  AND U9909 ( .A(b[23]), .B(a[95]), .Z(n3446) );
  XOR U9910 ( .A(n3451), .B(n3076), .Z(n3078) );
  XOR U9911 ( .A(n3452), .B(n3453), .Z(n3076) );
  AND U9912 ( .A(n3454), .B(n3455), .Z(n3452) );
  AND U9913 ( .A(b[22]), .B(a[96]), .Z(n3451) );
  XOR U9914 ( .A(n3456), .B(n3081), .Z(n3083) );
  XOR U9915 ( .A(n3457), .B(n3458), .Z(n3081) );
  AND U9916 ( .A(n3459), .B(n3460), .Z(n3457) );
  AND U9917 ( .A(b[21]), .B(a[97]), .Z(n3456) );
  XOR U9918 ( .A(n3461), .B(n3086), .Z(n3088) );
  XOR U9919 ( .A(n3462), .B(n3463), .Z(n3086) );
  AND U9920 ( .A(n3464), .B(n3465), .Z(n3462) );
  AND U9921 ( .A(b[20]), .B(a[98]), .Z(n3461) );
  XOR U9922 ( .A(n3466), .B(n3467), .Z(n3090) );
  AND U9923 ( .A(n3468), .B(n3469), .Z(n3466) );
  XOR U9924 ( .A(n3470), .B(n3095), .Z(n3097) );
  XOR U9925 ( .A(n3471), .B(n3472), .Z(n3095) );
  AND U9926 ( .A(n3473), .B(n3474), .Z(n3471) );
  AND U9927 ( .A(b[19]), .B(a[99]), .Z(n3470) );
  XOR U9928 ( .A(n3475), .B(n3100), .Z(n3102) );
  XOR U9929 ( .A(n3476), .B(n3477), .Z(n3100) );
  AND U9930 ( .A(n3478), .B(n3479), .Z(n3476) );
  AND U9931 ( .A(b[17]), .B(a[101]), .Z(n3475) );
  XOR U9932 ( .A(n3480), .B(n3105), .Z(n3107) );
  XOR U9933 ( .A(n3481), .B(n3482), .Z(n3105) );
  AND U9934 ( .A(n3483), .B(n3484), .Z(n3481) );
  AND U9935 ( .A(b[16]), .B(a[102]), .Z(n3480) );
  XOR U9936 ( .A(n3485), .B(n3110), .Z(n3112) );
  XOR U9937 ( .A(n3486), .B(n3487), .Z(n3110) );
  AND U9938 ( .A(n3488), .B(n3489), .Z(n3486) );
  AND U9939 ( .A(b[15]), .B(a[103]), .Z(n3485) );
  XOR U9940 ( .A(n3490), .B(n3115), .Z(n3117) );
  XOR U9941 ( .A(n3491), .B(n3492), .Z(n3115) );
  AND U9942 ( .A(n3493), .B(n3494), .Z(n3491) );
  AND U9943 ( .A(b[14]), .B(a[104]), .Z(n3490) );
  XOR U9944 ( .A(n3495), .B(n3496), .Z(n3119) );
  AND U9945 ( .A(n3497), .B(n3498), .Z(n3495) );
  XOR U9946 ( .A(n3499), .B(n3124), .Z(n3126) );
  XOR U9947 ( .A(n3500), .B(n3501), .Z(n3124) );
  AND U9948 ( .A(n3502), .B(n3503), .Z(n3500) );
  AND U9949 ( .A(b[13]), .B(a[105]), .Z(n3499) );
  XOR U9950 ( .A(n3504), .B(n3129), .Z(n3131) );
  XOR U9951 ( .A(n3505), .B(n3506), .Z(n3129) );
  AND U9952 ( .A(n3507), .B(n3508), .Z(n3505) );
  AND U9953 ( .A(b[11]), .B(a[107]), .Z(n3504) );
  XOR U9954 ( .A(n3509), .B(n3134), .Z(n3136) );
  XOR U9955 ( .A(n3510), .B(n3511), .Z(n3134) );
  AND U9956 ( .A(n3512), .B(n3513), .Z(n3510) );
  AND U9957 ( .A(b[10]), .B(a[108]), .Z(n3509) );
  XOR U9958 ( .A(n3514), .B(n3139), .Z(n3141) );
  XOR U9959 ( .A(n3515), .B(n3516), .Z(n3139) );
  AND U9960 ( .A(n3517), .B(n3518), .Z(n3515) );
  AND U9961 ( .A(b[9]), .B(a[109]), .Z(n3514) );
  XOR U9962 ( .A(n3519), .B(n3144), .Z(n3146) );
  XOR U9963 ( .A(n3520), .B(n3521), .Z(n3144) );
  AND U9964 ( .A(n3522), .B(n3523), .Z(n3520) );
  AND U9965 ( .A(b[8]), .B(a[110]), .Z(n3519) );
  XOR U9966 ( .A(n3524), .B(n3149), .Z(n3151) );
  XOR U9967 ( .A(n3525), .B(n3526), .Z(n3149) );
  AND U9968 ( .A(n3527), .B(n3528), .Z(n3525) );
  AND U9969 ( .A(b[7]), .B(a[111]), .Z(n3524) );
  XOR U9970 ( .A(n3529), .B(n3154), .Z(n3156) );
  XOR U9971 ( .A(n3530), .B(n3531), .Z(n3154) );
  AND U9972 ( .A(n3532), .B(n3533), .Z(n3530) );
  AND U9973 ( .A(b[6]), .B(a[112]), .Z(n3529) );
  XOR U9974 ( .A(n3534), .B(n3159), .Z(n3161) );
  XOR U9975 ( .A(n3535), .B(n3536), .Z(n3159) );
  AND U9976 ( .A(n3537), .B(n3538), .Z(n3535) );
  AND U9977 ( .A(b[5]), .B(a[113]), .Z(n3534) );
  XOR U9978 ( .A(n3539), .B(n3164), .Z(n3166) );
  XOR U9979 ( .A(n3540), .B(n3541), .Z(n3164) );
  AND U9980 ( .A(n3542), .B(n3543), .Z(n3540) );
  AND U9981 ( .A(b[4]), .B(a[114]), .Z(n3539) );
  XNOR U9982 ( .A(n3544), .B(n3545), .Z(n3178) );
  NANDN U9983 ( .A(n3546), .B(n3547), .Z(n3545) );
  XOR U9984 ( .A(n3548), .B(n3169), .Z(n3171) );
  XNOR U9985 ( .A(n3549), .B(n3550), .Z(n3169) );
  AND U9986 ( .A(n3551), .B(n3552), .Z(n3549) );
  AND U9987 ( .A(b[3]), .B(a[115]), .Z(n3548) );
  XOR U9988 ( .A(n3553), .B(n3554), .Z(swire[117]) );
  XOR U9989 ( .A(n3187), .B(n3555), .Z(n3554) );
  XNOR U9990 ( .A(n3188), .B(n3553), .Z(n3555) );
  NAND U9991 ( .A(a[117]), .B(b[0]), .Z(n3188) );
  XNOR U9992 ( .A(n3546), .B(n3547), .Z(n3187) );
  XOR U9993 ( .A(n3544), .B(n3556), .Z(n3547) );
  NAND U9994 ( .A(b[1]), .B(a[116]), .Z(n3556) );
  XOR U9995 ( .A(n3552), .B(n3557), .Z(n3546) );
  XOR U9996 ( .A(n3544), .B(n3551), .Z(n3557) );
  XNOR U9997 ( .A(n3558), .B(n3550), .Z(n3551) );
  AND U9998 ( .A(b[2]), .B(a[115]), .Z(n3558) );
  NANDN U9999 ( .A(n3559), .B(n3560), .Z(n3544) );
  XOR U10000 ( .A(n3550), .B(n3542), .Z(n3561) );
  XNOR U10001 ( .A(n3541), .B(n3537), .Z(n3562) );
  XNOR U10002 ( .A(n3536), .B(n3532), .Z(n3563) );
  XNOR U10003 ( .A(n3531), .B(n3527), .Z(n3564) );
  XNOR U10004 ( .A(n3526), .B(n3522), .Z(n3565) );
  XNOR U10005 ( .A(n3521), .B(n3517), .Z(n3566) );
  XNOR U10006 ( .A(n3516), .B(n3512), .Z(n3567) );
  XNOR U10007 ( .A(n3511), .B(n3507), .Z(n3568) );
  XNOR U10008 ( .A(n3498), .B(n3497), .Z(n3569) );
  XOR U10009 ( .A(n3570), .B(n3496), .Z(n3497) );
  AND U10010 ( .A(b[11]), .B(a[106]), .Z(n3570) );
  XNOR U10011 ( .A(n3496), .B(n3502), .Z(n3571) );
  XNOR U10012 ( .A(n3501), .B(n3493), .Z(n3572) );
  XNOR U10013 ( .A(n3492), .B(n3488), .Z(n3573) );
  XNOR U10014 ( .A(n3487), .B(n3483), .Z(n3574) );
  XNOR U10015 ( .A(n3482), .B(n3478), .Z(n3575) );
  XNOR U10016 ( .A(n3469), .B(n3468), .Z(n3576) );
  XOR U10017 ( .A(n3577), .B(n3467), .Z(n3468) );
  AND U10018 ( .A(b[17]), .B(a[100]), .Z(n3577) );
  XNOR U10019 ( .A(n3467), .B(n3473), .Z(n3578) );
  XNOR U10020 ( .A(n3472), .B(n3464), .Z(n3579) );
  XNOR U10021 ( .A(n3463), .B(n3459), .Z(n3580) );
  XNOR U10022 ( .A(n3458), .B(n3454), .Z(n3581) );
  XNOR U10023 ( .A(n3453), .B(n3449), .Z(n3582) );
  XNOR U10024 ( .A(n3440), .B(n3439), .Z(n3583) );
  XOR U10025 ( .A(n3584), .B(n3438), .Z(n3439) );
  AND U10026 ( .A(b[23]), .B(a[94]), .Z(n3584) );
  XNOR U10027 ( .A(n3438), .B(n3444), .Z(n3585) );
  XNOR U10028 ( .A(n3443), .B(n3435), .Z(n3586) );
  XNOR U10029 ( .A(n3434), .B(n3430), .Z(n3587) );
  XNOR U10030 ( .A(n3429), .B(n3425), .Z(n3588) );
  XNOR U10031 ( .A(n3424), .B(n3420), .Z(n3589) );
  XNOR U10032 ( .A(n3411), .B(n3410), .Z(n3590) );
  XOR U10033 ( .A(n3591), .B(n3409), .Z(n3410) );
  AND U10034 ( .A(b[29]), .B(a[88]), .Z(n3591) );
  XNOR U10035 ( .A(n3409), .B(n3415), .Z(n3592) );
  XNOR U10036 ( .A(n3414), .B(n3406), .Z(n3593) );
  XNOR U10037 ( .A(n3405), .B(n3401), .Z(n3594) );
  XNOR U10038 ( .A(n3400), .B(n3396), .Z(n3595) );
  XNOR U10039 ( .A(n3395), .B(n3391), .Z(n3596) );
  XNOR U10040 ( .A(n3382), .B(n3381), .Z(n3597) );
  XOR U10041 ( .A(n3598), .B(n3380), .Z(n3381) );
  AND U10042 ( .A(b[35]), .B(a[82]), .Z(n3598) );
  XNOR U10043 ( .A(n3380), .B(n3386), .Z(n3599) );
  XNOR U10044 ( .A(n3385), .B(n3377), .Z(n3600) );
  XNOR U10045 ( .A(n3376), .B(n3372), .Z(n3601) );
  XNOR U10046 ( .A(n3371), .B(n3367), .Z(n3602) );
  XNOR U10047 ( .A(n3366), .B(n3362), .Z(n3603) );
  XNOR U10048 ( .A(n3353), .B(n3352), .Z(n3604) );
  XOR U10049 ( .A(n3605), .B(n3351), .Z(n3352) );
  AND U10050 ( .A(b[41]), .B(a[76]), .Z(n3605) );
  XNOR U10051 ( .A(n3351), .B(n3357), .Z(n3606) );
  XNOR U10052 ( .A(n3356), .B(n3348), .Z(n3607) );
  XNOR U10053 ( .A(n3347), .B(n3343), .Z(n3608) );
  XNOR U10054 ( .A(n3342), .B(n3338), .Z(n3609) );
  XNOR U10055 ( .A(n3337), .B(n3333), .Z(n3610) );
  XNOR U10056 ( .A(n3324), .B(n3323), .Z(n3611) );
  XOR U10057 ( .A(n3612), .B(n3322), .Z(n3323) );
  AND U10058 ( .A(b[47]), .B(a[70]), .Z(n3612) );
  XNOR U10059 ( .A(n3322), .B(n3328), .Z(n3613) );
  XNOR U10060 ( .A(n3327), .B(n3319), .Z(n3614) );
  XNOR U10061 ( .A(n3318), .B(n3314), .Z(n3615) );
  XNOR U10062 ( .A(n3313), .B(n3309), .Z(n3616) );
  XNOR U10063 ( .A(n3308), .B(n3304), .Z(n3617) );
  XNOR U10064 ( .A(n3303), .B(n3299), .Z(n3618) );
  XNOR U10065 ( .A(n3298), .B(n3294), .Z(n3619) );
  XNOR U10066 ( .A(n3293), .B(n3289), .Z(n3620) );
  XNOR U10067 ( .A(n3288), .B(n3284), .Z(n3621) );
  XNOR U10068 ( .A(n3283), .B(n3279), .Z(n3622) );
  XNOR U10069 ( .A(n3278), .B(n3274), .Z(n3623) );
  XNOR U10070 ( .A(n3273), .B(n3269), .Z(n3624) );
  XOR U10071 ( .A(n3268), .B(n3265), .Z(n3625) );
  XOR U10072 ( .A(n3626), .B(n3627), .Z(n3265) );
  XOR U10073 ( .A(n3263), .B(n3628), .Z(n3627) );
  XOR U10074 ( .A(n3629), .B(n3630), .Z(n3628) );
  XOR U10075 ( .A(n3631), .B(n3632), .Z(n3630) );
  NAND U10076 ( .A(a[55]), .B(b[62]), .Z(n3632) );
  AND U10077 ( .A(a[54]), .B(b[63]), .Z(n3631) );
  XOR U10078 ( .A(n3633), .B(n3629), .Z(n3626) );
  XOR U10079 ( .A(n3634), .B(n3635), .Z(n3629) );
  ANDN U10080 ( .B(n3636), .A(n3637), .Z(n3634) );
  AND U10081 ( .A(a[56]), .B(b[61]), .Z(n3633) );
  XOR U10082 ( .A(n3638), .B(n3263), .Z(n3264) );
  XOR U10083 ( .A(n3639), .B(n3640), .Z(n3263) );
  AND U10084 ( .A(n3641), .B(n3642), .Z(n3639) );
  AND U10085 ( .A(a[57]), .B(b[60]), .Z(n3638) );
  XOR U10086 ( .A(n3643), .B(n3268), .Z(n3270) );
  XOR U10087 ( .A(n3644), .B(n3645), .Z(n3268) );
  AND U10088 ( .A(n3646), .B(n3647), .Z(n3644) );
  AND U10089 ( .A(a[58]), .B(b[59]), .Z(n3643) );
  XOR U10090 ( .A(n3648), .B(n3273), .Z(n3275) );
  XOR U10091 ( .A(n3649), .B(n3650), .Z(n3273) );
  AND U10092 ( .A(n3651), .B(n3652), .Z(n3649) );
  AND U10093 ( .A(b[58]), .B(a[59]), .Z(n3648) );
  XOR U10094 ( .A(n3653), .B(n3278), .Z(n3280) );
  XOR U10095 ( .A(n3654), .B(n3655), .Z(n3278) );
  AND U10096 ( .A(n3656), .B(n3657), .Z(n3654) );
  AND U10097 ( .A(b[57]), .B(a[60]), .Z(n3653) );
  XOR U10098 ( .A(n3658), .B(n3283), .Z(n3285) );
  XOR U10099 ( .A(n3659), .B(n3660), .Z(n3283) );
  AND U10100 ( .A(n3661), .B(n3662), .Z(n3659) );
  AND U10101 ( .A(b[56]), .B(a[61]), .Z(n3658) );
  XOR U10102 ( .A(n3663), .B(n3288), .Z(n3290) );
  XOR U10103 ( .A(n3664), .B(n3665), .Z(n3288) );
  AND U10104 ( .A(n3666), .B(n3667), .Z(n3664) );
  AND U10105 ( .A(b[55]), .B(a[62]), .Z(n3663) );
  XOR U10106 ( .A(n3668), .B(n3293), .Z(n3295) );
  XOR U10107 ( .A(n3669), .B(n3670), .Z(n3293) );
  AND U10108 ( .A(n3671), .B(n3672), .Z(n3669) );
  AND U10109 ( .A(b[54]), .B(a[63]), .Z(n3668) );
  XOR U10110 ( .A(n3673), .B(n3298), .Z(n3300) );
  XOR U10111 ( .A(n3674), .B(n3675), .Z(n3298) );
  AND U10112 ( .A(n3676), .B(n3677), .Z(n3674) );
  AND U10113 ( .A(b[53]), .B(a[64]), .Z(n3673) );
  XOR U10114 ( .A(n3678), .B(n3303), .Z(n3305) );
  XOR U10115 ( .A(n3679), .B(n3680), .Z(n3303) );
  AND U10116 ( .A(n3681), .B(n3682), .Z(n3679) );
  AND U10117 ( .A(b[52]), .B(a[65]), .Z(n3678) );
  XOR U10118 ( .A(n3683), .B(n3308), .Z(n3310) );
  XOR U10119 ( .A(n3684), .B(n3685), .Z(n3308) );
  AND U10120 ( .A(n3686), .B(n3687), .Z(n3684) );
  AND U10121 ( .A(b[51]), .B(a[66]), .Z(n3683) );
  XOR U10122 ( .A(n3688), .B(n3313), .Z(n3315) );
  XOR U10123 ( .A(n3689), .B(n3690), .Z(n3313) );
  AND U10124 ( .A(n3691), .B(n3692), .Z(n3689) );
  AND U10125 ( .A(b[50]), .B(a[67]), .Z(n3688) );
  XOR U10126 ( .A(n3693), .B(n3318), .Z(n3320) );
  XOR U10127 ( .A(n3694), .B(n3695), .Z(n3318) );
  AND U10128 ( .A(n3696), .B(n3697), .Z(n3694) );
  AND U10129 ( .A(b[49]), .B(a[68]), .Z(n3693) );
  XOR U10130 ( .A(n3698), .B(n3699), .Z(n3322) );
  AND U10131 ( .A(n3700), .B(n3701), .Z(n3698) );
  XOR U10132 ( .A(n3702), .B(n3327), .Z(n3329) );
  XOR U10133 ( .A(n3703), .B(n3704), .Z(n3327) );
  AND U10134 ( .A(n3705), .B(n3706), .Z(n3703) );
  AND U10135 ( .A(b[48]), .B(a[69]), .Z(n3702) );
  XOR U10136 ( .A(n3707), .B(n3332), .Z(n3334) );
  XOR U10137 ( .A(n3708), .B(n3709), .Z(n3332) );
  AND U10138 ( .A(n3710), .B(n3711), .Z(n3708) );
  AND U10139 ( .A(b[46]), .B(a[71]), .Z(n3707) );
  XOR U10140 ( .A(n3712), .B(n3337), .Z(n3339) );
  XOR U10141 ( .A(n3713), .B(n3714), .Z(n3337) );
  AND U10142 ( .A(n3715), .B(n3716), .Z(n3713) );
  AND U10143 ( .A(b[45]), .B(a[72]), .Z(n3712) );
  XOR U10144 ( .A(n3717), .B(n3342), .Z(n3344) );
  XOR U10145 ( .A(n3718), .B(n3719), .Z(n3342) );
  AND U10146 ( .A(n3720), .B(n3721), .Z(n3718) );
  AND U10147 ( .A(b[44]), .B(a[73]), .Z(n3717) );
  XOR U10148 ( .A(n3722), .B(n3347), .Z(n3349) );
  XOR U10149 ( .A(n3723), .B(n3724), .Z(n3347) );
  AND U10150 ( .A(n3725), .B(n3726), .Z(n3723) );
  AND U10151 ( .A(b[43]), .B(a[74]), .Z(n3722) );
  XOR U10152 ( .A(n3727), .B(n3728), .Z(n3351) );
  AND U10153 ( .A(n3729), .B(n3730), .Z(n3727) );
  XOR U10154 ( .A(n3731), .B(n3356), .Z(n3358) );
  XOR U10155 ( .A(n3732), .B(n3733), .Z(n3356) );
  AND U10156 ( .A(n3734), .B(n3735), .Z(n3732) );
  AND U10157 ( .A(b[42]), .B(a[75]), .Z(n3731) );
  XOR U10158 ( .A(n3736), .B(n3361), .Z(n3363) );
  XOR U10159 ( .A(n3737), .B(n3738), .Z(n3361) );
  AND U10160 ( .A(n3739), .B(n3740), .Z(n3737) );
  AND U10161 ( .A(b[40]), .B(a[77]), .Z(n3736) );
  XOR U10162 ( .A(n3741), .B(n3366), .Z(n3368) );
  XOR U10163 ( .A(n3742), .B(n3743), .Z(n3366) );
  AND U10164 ( .A(n3744), .B(n3745), .Z(n3742) );
  AND U10165 ( .A(b[39]), .B(a[78]), .Z(n3741) );
  XOR U10166 ( .A(n3746), .B(n3371), .Z(n3373) );
  XOR U10167 ( .A(n3747), .B(n3748), .Z(n3371) );
  AND U10168 ( .A(n3749), .B(n3750), .Z(n3747) );
  AND U10169 ( .A(b[38]), .B(a[79]), .Z(n3746) );
  XOR U10170 ( .A(n3751), .B(n3376), .Z(n3378) );
  XOR U10171 ( .A(n3752), .B(n3753), .Z(n3376) );
  AND U10172 ( .A(n3754), .B(n3755), .Z(n3752) );
  AND U10173 ( .A(b[37]), .B(a[80]), .Z(n3751) );
  XOR U10174 ( .A(n3756), .B(n3757), .Z(n3380) );
  AND U10175 ( .A(n3758), .B(n3759), .Z(n3756) );
  XOR U10176 ( .A(n3760), .B(n3385), .Z(n3387) );
  XOR U10177 ( .A(n3761), .B(n3762), .Z(n3385) );
  AND U10178 ( .A(n3763), .B(n3764), .Z(n3761) );
  AND U10179 ( .A(b[36]), .B(a[81]), .Z(n3760) );
  XOR U10180 ( .A(n3765), .B(n3390), .Z(n3392) );
  XOR U10181 ( .A(n3766), .B(n3767), .Z(n3390) );
  AND U10182 ( .A(n3768), .B(n3769), .Z(n3766) );
  AND U10183 ( .A(b[34]), .B(a[83]), .Z(n3765) );
  XOR U10184 ( .A(n3770), .B(n3395), .Z(n3397) );
  XOR U10185 ( .A(n3771), .B(n3772), .Z(n3395) );
  AND U10186 ( .A(n3773), .B(n3774), .Z(n3771) );
  AND U10187 ( .A(b[33]), .B(a[84]), .Z(n3770) );
  XOR U10188 ( .A(n3775), .B(n3400), .Z(n3402) );
  XOR U10189 ( .A(n3776), .B(n3777), .Z(n3400) );
  AND U10190 ( .A(n3778), .B(n3779), .Z(n3776) );
  AND U10191 ( .A(b[32]), .B(a[85]), .Z(n3775) );
  XOR U10192 ( .A(n3780), .B(n3405), .Z(n3407) );
  XOR U10193 ( .A(n3781), .B(n3782), .Z(n3405) );
  AND U10194 ( .A(n3783), .B(n3784), .Z(n3781) );
  AND U10195 ( .A(b[31]), .B(a[86]), .Z(n3780) );
  XOR U10196 ( .A(n3785), .B(n3786), .Z(n3409) );
  AND U10197 ( .A(n3787), .B(n3788), .Z(n3785) );
  XOR U10198 ( .A(n3789), .B(n3414), .Z(n3416) );
  XOR U10199 ( .A(n3790), .B(n3791), .Z(n3414) );
  AND U10200 ( .A(n3792), .B(n3793), .Z(n3790) );
  AND U10201 ( .A(b[30]), .B(a[87]), .Z(n3789) );
  XOR U10202 ( .A(n3794), .B(n3419), .Z(n3421) );
  XOR U10203 ( .A(n3795), .B(n3796), .Z(n3419) );
  AND U10204 ( .A(n3797), .B(n3798), .Z(n3795) );
  AND U10205 ( .A(b[28]), .B(a[89]), .Z(n3794) );
  XOR U10206 ( .A(n3799), .B(n3424), .Z(n3426) );
  XOR U10207 ( .A(n3800), .B(n3801), .Z(n3424) );
  AND U10208 ( .A(n3802), .B(n3803), .Z(n3800) );
  AND U10209 ( .A(b[27]), .B(a[90]), .Z(n3799) );
  XOR U10210 ( .A(n3804), .B(n3429), .Z(n3431) );
  XOR U10211 ( .A(n3805), .B(n3806), .Z(n3429) );
  AND U10212 ( .A(n3807), .B(n3808), .Z(n3805) );
  AND U10213 ( .A(b[26]), .B(a[91]), .Z(n3804) );
  XOR U10214 ( .A(n3809), .B(n3434), .Z(n3436) );
  XOR U10215 ( .A(n3810), .B(n3811), .Z(n3434) );
  AND U10216 ( .A(n3812), .B(n3813), .Z(n3810) );
  AND U10217 ( .A(b[25]), .B(a[92]), .Z(n3809) );
  XOR U10218 ( .A(n3814), .B(n3815), .Z(n3438) );
  AND U10219 ( .A(n3816), .B(n3817), .Z(n3814) );
  XOR U10220 ( .A(n3818), .B(n3443), .Z(n3445) );
  XOR U10221 ( .A(n3819), .B(n3820), .Z(n3443) );
  AND U10222 ( .A(n3821), .B(n3822), .Z(n3819) );
  AND U10223 ( .A(b[24]), .B(a[93]), .Z(n3818) );
  XOR U10224 ( .A(n3823), .B(n3448), .Z(n3450) );
  XOR U10225 ( .A(n3824), .B(n3825), .Z(n3448) );
  AND U10226 ( .A(n3826), .B(n3827), .Z(n3824) );
  AND U10227 ( .A(b[22]), .B(a[95]), .Z(n3823) );
  XOR U10228 ( .A(n3828), .B(n3453), .Z(n3455) );
  XOR U10229 ( .A(n3829), .B(n3830), .Z(n3453) );
  AND U10230 ( .A(n3831), .B(n3832), .Z(n3829) );
  AND U10231 ( .A(b[21]), .B(a[96]), .Z(n3828) );
  XOR U10232 ( .A(n3833), .B(n3458), .Z(n3460) );
  XOR U10233 ( .A(n3834), .B(n3835), .Z(n3458) );
  AND U10234 ( .A(n3836), .B(n3837), .Z(n3834) );
  AND U10235 ( .A(b[20]), .B(a[97]), .Z(n3833) );
  XOR U10236 ( .A(n3838), .B(n3463), .Z(n3465) );
  XOR U10237 ( .A(n3839), .B(n3840), .Z(n3463) );
  AND U10238 ( .A(n3841), .B(n3842), .Z(n3839) );
  AND U10239 ( .A(b[19]), .B(a[98]), .Z(n3838) );
  XOR U10240 ( .A(n3843), .B(n3844), .Z(n3467) );
  AND U10241 ( .A(n3845), .B(n3846), .Z(n3843) );
  XOR U10242 ( .A(n3847), .B(n3472), .Z(n3474) );
  XOR U10243 ( .A(n3848), .B(n3849), .Z(n3472) );
  AND U10244 ( .A(n3850), .B(n3851), .Z(n3848) );
  AND U10245 ( .A(b[18]), .B(a[99]), .Z(n3847) );
  XOR U10246 ( .A(n3852), .B(n3477), .Z(n3479) );
  XOR U10247 ( .A(n3853), .B(n3854), .Z(n3477) );
  AND U10248 ( .A(n3855), .B(n3856), .Z(n3853) );
  AND U10249 ( .A(b[16]), .B(a[101]), .Z(n3852) );
  XOR U10250 ( .A(n3857), .B(n3482), .Z(n3484) );
  XOR U10251 ( .A(n3858), .B(n3859), .Z(n3482) );
  AND U10252 ( .A(n3860), .B(n3861), .Z(n3858) );
  AND U10253 ( .A(b[15]), .B(a[102]), .Z(n3857) );
  XOR U10254 ( .A(n3862), .B(n3487), .Z(n3489) );
  XOR U10255 ( .A(n3863), .B(n3864), .Z(n3487) );
  AND U10256 ( .A(n3865), .B(n3866), .Z(n3863) );
  AND U10257 ( .A(b[14]), .B(a[103]), .Z(n3862) );
  XOR U10258 ( .A(n3867), .B(n3492), .Z(n3494) );
  XOR U10259 ( .A(n3868), .B(n3869), .Z(n3492) );
  AND U10260 ( .A(n3870), .B(n3871), .Z(n3868) );
  AND U10261 ( .A(b[13]), .B(a[104]), .Z(n3867) );
  XOR U10262 ( .A(n3872), .B(n3873), .Z(n3496) );
  AND U10263 ( .A(n3874), .B(n3875), .Z(n3872) );
  XOR U10264 ( .A(n3876), .B(n3501), .Z(n3503) );
  XOR U10265 ( .A(n3877), .B(n3878), .Z(n3501) );
  AND U10266 ( .A(n3879), .B(n3880), .Z(n3877) );
  AND U10267 ( .A(b[12]), .B(a[105]), .Z(n3876) );
  XOR U10268 ( .A(n3881), .B(n3506), .Z(n3508) );
  XOR U10269 ( .A(n3882), .B(n3883), .Z(n3506) );
  AND U10270 ( .A(n3884), .B(n3885), .Z(n3882) );
  AND U10271 ( .A(b[10]), .B(a[107]), .Z(n3881) );
  XOR U10272 ( .A(n3886), .B(n3511), .Z(n3513) );
  XOR U10273 ( .A(n3887), .B(n3888), .Z(n3511) );
  AND U10274 ( .A(n3889), .B(n3890), .Z(n3887) );
  AND U10275 ( .A(b[9]), .B(a[108]), .Z(n3886) );
  XOR U10276 ( .A(n3891), .B(n3516), .Z(n3518) );
  XOR U10277 ( .A(n3892), .B(n3893), .Z(n3516) );
  AND U10278 ( .A(n3894), .B(n3895), .Z(n3892) );
  AND U10279 ( .A(b[8]), .B(a[109]), .Z(n3891) );
  XOR U10280 ( .A(n3896), .B(n3521), .Z(n3523) );
  XOR U10281 ( .A(n3897), .B(n3898), .Z(n3521) );
  AND U10282 ( .A(n3899), .B(n3900), .Z(n3897) );
  AND U10283 ( .A(b[7]), .B(a[110]), .Z(n3896) );
  XOR U10284 ( .A(n3901), .B(n3526), .Z(n3528) );
  XOR U10285 ( .A(n3902), .B(n3903), .Z(n3526) );
  AND U10286 ( .A(n3904), .B(n3905), .Z(n3902) );
  AND U10287 ( .A(b[6]), .B(a[111]), .Z(n3901) );
  XOR U10288 ( .A(n3906), .B(n3531), .Z(n3533) );
  XOR U10289 ( .A(n3907), .B(n3908), .Z(n3531) );
  AND U10290 ( .A(n3909), .B(n3910), .Z(n3907) );
  AND U10291 ( .A(b[5]), .B(a[112]), .Z(n3906) );
  XOR U10292 ( .A(n3911), .B(n3536), .Z(n3538) );
  XOR U10293 ( .A(n3912), .B(n3913), .Z(n3536) );
  AND U10294 ( .A(n3914), .B(n3915), .Z(n3912) );
  AND U10295 ( .A(b[4]), .B(a[113]), .Z(n3911) );
  XNOR U10296 ( .A(n3916), .B(n3917), .Z(n3550) );
  NANDN U10297 ( .A(n3918), .B(n3919), .Z(n3917) );
  XOR U10298 ( .A(n3920), .B(n3541), .Z(n3543) );
  XNOR U10299 ( .A(n3921), .B(n3922), .Z(n3541) );
  AND U10300 ( .A(n3923), .B(n3924), .Z(n3921) );
  AND U10301 ( .A(b[3]), .B(a[114]), .Z(n3920) );
  XOR U10302 ( .A(n3925), .B(n3926), .Z(swire[116]) );
  XOR U10303 ( .A(n3560), .B(n3927), .Z(n3926) );
  XNOR U10304 ( .A(n3559), .B(n3925), .Z(n3927) );
  NAND U10305 ( .A(a[116]), .B(b[0]), .Z(n3559) );
  XNOR U10306 ( .A(n3918), .B(n3919), .Z(n3560) );
  XOR U10307 ( .A(n3916), .B(n3928), .Z(n3919) );
  NAND U10308 ( .A(b[1]), .B(a[115]), .Z(n3928) );
  XOR U10309 ( .A(n3924), .B(n3929), .Z(n3918) );
  XOR U10310 ( .A(n3916), .B(n3923), .Z(n3929) );
  XNOR U10311 ( .A(n3930), .B(n3922), .Z(n3923) );
  AND U10312 ( .A(b[2]), .B(a[114]), .Z(n3930) );
  NANDN U10313 ( .A(n3931), .B(n3932), .Z(n3916) );
  XOR U10314 ( .A(n3922), .B(n3914), .Z(n3933) );
  XNOR U10315 ( .A(n3913), .B(n3909), .Z(n3934) );
  XNOR U10316 ( .A(n3908), .B(n3904), .Z(n3935) );
  XNOR U10317 ( .A(n3903), .B(n3899), .Z(n3936) );
  XNOR U10318 ( .A(n3898), .B(n3894), .Z(n3937) );
  XNOR U10319 ( .A(n3893), .B(n3889), .Z(n3938) );
  XNOR U10320 ( .A(n3888), .B(n3884), .Z(n3939) );
  XNOR U10321 ( .A(n3875), .B(n3874), .Z(n3940) );
  XOR U10322 ( .A(n3941), .B(n3873), .Z(n3874) );
  AND U10323 ( .A(b[10]), .B(a[106]), .Z(n3941) );
  XNOR U10324 ( .A(n3873), .B(n3879), .Z(n3942) );
  XNOR U10325 ( .A(n3878), .B(n3870), .Z(n3943) );
  XNOR U10326 ( .A(n3869), .B(n3865), .Z(n3944) );
  XNOR U10327 ( .A(n3864), .B(n3860), .Z(n3945) );
  XNOR U10328 ( .A(n3859), .B(n3855), .Z(n3946) );
  XNOR U10329 ( .A(n3846), .B(n3845), .Z(n3947) );
  XOR U10330 ( .A(n3948), .B(n3844), .Z(n3845) );
  AND U10331 ( .A(b[16]), .B(a[100]), .Z(n3948) );
  XNOR U10332 ( .A(n3844), .B(n3850), .Z(n3949) );
  XNOR U10333 ( .A(n3849), .B(n3841), .Z(n3950) );
  XNOR U10334 ( .A(n3840), .B(n3836), .Z(n3951) );
  XNOR U10335 ( .A(n3835), .B(n3831), .Z(n3952) );
  XNOR U10336 ( .A(n3830), .B(n3826), .Z(n3953) );
  XNOR U10337 ( .A(n3817), .B(n3816), .Z(n3954) );
  XOR U10338 ( .A(n3955), .B(n3815), .Z(n3816) );
  AND U10339 ( .A(b[22]), .B(a[94]), .Z(n3955) );
  XNOR U10340 ( .A(n3815), .B(n3821), .Z(n3956) );
  XNOR U10341 ( .A(n3820), .B(n3812), .Z(n3957) );
  XNOR U10342 ( .A(n3811), .B(n3807), .Z(n3958) );
  XNOR U10343 ( .A(n3806), .B(n3802), .Z(n3959) );
  XNOR U10344 ( .A(n3801), .B(n3797), .Z(n3960) );
  XNOR U10345 ( .A(n3788), .B(n3787), .Z(n3961) );
  XOR U10346 ( .A(n3962), .B(n3786), .Z(n3787) );
  AND U10347 ( .A(b[28]), .B(a[88]), .Z(n3962) );
  XNOR U10348 ( .A(n3786), .B(n3792), .Z(n3963) );
  XNOR U10349 ( .A(n3791), .B(n3783), .Z(n3964) );
  XNOR U10350 ( .A(n3782), .B(n3778), .Z(n3965) );
  XNOR U10351 ( .A(n3777), .B(n3773), .Z(n3966) );
  XNOR U10352 ( .A(n3772), .B(n3768), .Z(n3967) );
  XNOR U10353 ( .A(n3759), .B(n3758), .Z(n3968) );
  XOR U10354 ( .A(n3969), .B(n3757), .Z(n3758) );
  AND U10355 ( .A(b[34]), .B(a[82]), .Z(n3969) );
  XNOR U10356 ( .A(n3757), .B(n3763), .Z(n3970) );
  XNOR U10357 ( .A(n3762), .B(n3754), .Z(n3971) );
  XNOR U10358 ( .A(n3753), .B(n3749), .Z(n3972) );
  XNOR U10359 ( .A(n3748), .B(n3744), .Z(n3973) );
  XNOR U10360 ( .A(n3743), .B(n3739), .Z(n3974) );
  XNOR U10361 ( .A(n3730), .B(n3729), .Z(n3975) );
  XOR U10362 ( .A(n3976), .B(n3728), .Z(n3729) );
  AND U10363 ( .A(b[40]), .B(a[76]), .Z(n3976) );
  XNOR U10364 ( .A(n3728), .B(n3734), .Z(n3977) );
  XNOR U10365 ( .A(n3733), .B(n3725), .Z(n3978) );
  XNOR U10366 ( .A(n3724), .B(n3720), .Z(n3979) );
  XNOR U10367 ( .A(n3719), .B(n3715), .Z(n3980) );
  XNOR U10368 ( .A(n3714), .B(n3710), .Z(n3981) );
  XNOR U10369 ( .A(n3701), .B(n3700), .Z(n3982) );
  XOR U10370 ( .A(n3983), .B(n3699), .Z(n3700) );
  AND U10371 ( .A(b[46]), .B(a[70]), .Z(n3983) );
  XNOR U10372 ( .A(n3699), .B(n3705), .Z(n3984) );
  XNOR U10373 ( .A(n3704), .B(n3696), .Z(n3985) );
  XNOR U10374 ( .A(n3695), .B(n3691), .Z(n3986) );
  XNOR U10375 ( .A(n3690), .B(n3686), .Z(n3987) );
  XNOR U10376 ( .A(n3685), .B(n3681), .Z(n3988) );
  XNOR U10377 ( .A(n3680), .B(n3676), .Z(n3989) );
  XNOR U10378 ( .A(n3675), .B(n3671), .Z(n3990) );
  XNOR U10379 ( .A(n3670), .B(n3666), .Z(n3991) );
  XNOR U10380 ( .A(n3665), .B(n3661), .Z(n3992) );
  XNOR U10381 ( .A(n3660), .B(n3656), .Z(n3993) );
  XNOR U10382 ( .A(n3655), .B(n3651), .Z(n3994) );
  XNOR U10383 ( .A(n3650), .B(n3646), .Z(n3995) );
  XNOR U10384 ( .A(n3645), .B(n3641), .Z(n3996) );
  XOR U10385 ( .A(n3640), .B(n3637), .Z(n3997) );
  XOR U10386 ( .A(n3998), .B(n3999), .Z(n3637) );
  XOR U10387 ( .A(n3635), .B(n4000), .Z(n3999) );
  XOR U10388 ( .A(n4001), .B(n4002), .Z(n4000) );
  XOR U10389 ( .A(n4003), .B(n4004), .Z(n4002) );
  NAND U10390 ( .A(a[54]), .B(b[62]), .Z(n4004) );
  AND U10391 ( .A(a[53]), .B(b[63]), .Z(n4003) );
  XOR U10392 ( .A(n4005), .B(n4001), .Z(n3998) );
  XOR U10393 ( .A(n4006), .B(n4007), .Z(n4001) );
  ANDN U10394 ( .B(n4008), .A(n4009), .Z(n4006) );
  AND U10395 ( .A(a[55]), .B(b[61]), .Z(n4005) );
  XOR U10396 ( .A(n4010), .B(n3635), .Z(n3636) );
  XOR U10397 ( .A(n4011), .B(n4012), .Z(n3635) );
  AND U10398 ( .A(n4013), .B(n4014), .Z(n4011) );
  AND U10399 ( .A(a[56]), .B(b[60]), .Z(n4010) );
  XOR U10400 ( .A(n4015), .B(n3640), .Z(n3642) );
  XOR U10401 ( .A(n4016), .B(n4017), .Z(n3640) );
  AND U10402 ( .A(n4018), .B(n4019), .Z(n4016) );
  AND U10403 ( .A(a[57]), .B(b[59]), .Z(n4015) );
  XOR U10404 ( .A(n4020), .B(n3645), .Z(n3647) );
  XOR U10405 ( .A(n4021), .B(n4022), .Z(n3645) );
  AND U10406 ( .A(n4023), .B(n4024), .Z(n4021) );
  AND U10407 ( .A(a[58]), .B(b[58]), .Z(n4020) );
  XOR U10408 ( .A(n4025), .B(n3650), .Z(n3652) );
  XOR U10409 ( .A(n4026), .B(n4027), .Z(n3650) );
  AND U10410 ( .A(n4028), .B(n4029), .Z(n4026) );
  AND U10411 ( .A(b[57]), .B(a[59]), .Z(n4025) );
  XOR U10412 ( .A(n4030), .B(n3655), .Z(n3657) );
  XOR U10413 ( .A(n4031), .B(n4032), .Z(n3655) );
  AND U10414 ( .A(n4033), .B(n4034), .Z(n4031) );
  AND U10415 ( .A(b[56]), .B(a[60]), .Z(n4030) );
  XOR U10416 ( .A(n4035), .B(n3660), .Z(n3662) );
  XOR U10417 ( .A(n4036), .B(n4037), .Z(n3660) );
  AND U10418 ( .A(n4038), .B(n4039), .Z(n4036) );
  AND U10419 ( .A(b[55]), .B(a[61]), .Z(n4035) );
  XOR U10420 ( .A(n4040), .B(n3665), .Z(n3667) );
  XOR U10421 ( .A(n4041), .B(n4042), .Z(n3665) );
  AND U10422 ( .A(n4043), .B(n4044), .Z(n4041) );
  AND U10423 ( .A(b[54]), .B(a[62]), .Z(n4040) );
  XOR U10424 ( .A(n4045), .B(n3670), .Z(n3672) );
  XOR U10425 ( .A(n4046), .B(n4047), .Z(n3670) );
  AND U10426 ( .A(n4048), .B(n4049), .Z(n4046) );
  AND U10427 ( .A(b[53]), .B(a[63]), .Z(n4045) );
  XOR U10428 ( .A(n4050), .B(n3675), .Z(n3677) );
  XOR U10429 ( .A(n4051), .B(n4052), .Z(n3675) );
  AND U10430 ( .A(n4053), .B(n4054), .Z(n4051) );
  AND U10431 ( .A(b[52]), .B(a[64]), .Z(n4050) );
  XOR U10432 ( .A(n4055), .B(n3680), .Z(n3682) );
  XOR U10433 ( .A(n4056), .B(n4057), .Z(n3680) );
  AND U10434 ( .A(n4058), .B(n4059), .Z(n4056) );
  AND U10435 ( .A(b[51]), .B(a[65]), .Z(n4055) );
  XOR U10436 ( .A(n4060), .B(n3685), .Z(n3687) );
  XOR U10437 ( .A(n4061), .B(n4062), .Z(n3685) );
  AND U10438 ( .A(n4063), .B(n4064), .Z(n4061) );
  AND U10439 ( .A(b[50]), .B(a[66]), .Z(n4060) );
  XOR U10440 ( .A(n4065), .B(n3690), .Z(n3692) );
  XOR U10441 ( .A(n4066), .B(n4067), .Z(n3690) );
  AND U10442 ( .A(n4068), .B(n4069), .Z(n4066) );
  AND U10443 ( .A(b[49]), .B(a[67]), .Z(n4065) );
  XOR U10444 ( .A(n4070), .B(n3695), .Z(n3697) );
  XOR U10445 ( .A(n4071), .B(n4072), .Z(n3695) );
  AND U10446 ( .A(n4073), .B(n4074), .Z(n4071) );
  AND U10447 ( .A(b[48]), .B(a[68]), .Z(n4070) );
  XOR U10448 ( .A(n4075), .B(n4076), .Z(n3699) );
  AND U10449 ( .A(n4077), .B(n4078), .Z(n4075) );
  XOR U10450 ( .A(n4079), .B(n3704), .Z(n3706) );
  XOR U10451 ( .A(n4080), .B(n4081), .Z(n3704) );
  AND U10452 ( .A(n4082), .B(n4083), .Z(n4080) );
  AND U10453 ( .A(b[47]), .B(a[69]), .Z(n4079) );
  XOR U10454 ( .A(n4084), .B(n3709), .Z(n3711) );
  XOR U10455 ( .A(n4085), .B(n4086), .Z(n3709) );
  AND U10456 ( .A(n4087), .B(n4088), .Z(n4085) );
  AND U10457 ( .A(b[45]), .B(a[71]), .Z(n4084) );
  XOR U10458 ( .A(n4089), .B(n3714), .Z(n3716) );
  XOR U10459 ( .A(n4090), .B(n4091), .Z(n3714) );
  AND U10460 ( .A(n4092), .B(n4093), .Z(n4090) );
  AND U10461 ( .A(b[44]), .B(a[72]), .Z(n4089) );
  XOR U10462 ( .A(n4094), .B(n3719), .Z(n3721) );
  XOR U10463 ( .A(n4095), .B(n4096), .Z(n3719) );
  AND U10464 ( .A(n4097), .B(n4098), .Z(n4095) );
  AND U10465 ( .A(b[43]), .B(a[73]), .Z(n4094) );
  XOR U10466 ( .A(n4099), .B(n3724), .Z(n3726) );
  XOR U10467 ( .A(n4100), .B(n4101), .Z(n3724) );
  AND U10468 ( .A(n4102), .B(n4103), .Z(n4100) );
  AND U10469 ( .A(b[42]), .B(a[74]), .Z(n4099) );
  XOR U10470 ( .A(n4104), .B(n4105), .Z(n3728) );
  AND U10471 ( .A(n4106), .B(n4107), .Z(n4104) );
  XOR U10472 ( .A(n4108), .B(n3733), .Z(n3735) );
  XOR U10473 ( .A(n4109), .B(n4110), .Z(n3733) );
  AND U10474 ( .A(n4111), .B(n4112), .Z(n4109) );
  AND U10475 ( .A(b[41]), .B(a[75]), .Z(n4108) );
  XOR U10476 ( .A(n4113), .B(n3738), .Z(n3740) );
  XOR U10477 ( .A(n4114), .B(n4115), .Z(n3738) );
  AND U10478 ( .A(n4116), .B(n4117), .Z(n4114) );
  AND U10479 ( .A(b[39]), .B(a[77]), .Z(n4113) );
  XOR U10480 ( .A(n4118), .B(n3743), .Z(n3745) );
  XOR U10481 ( .A(n4119), .B(n4120), .Z(n3743) );
  AND U10482 ( .A(n4121), .B(n4122), .Z(n4119) );
  AND U10483 ( .A(b[38]), .B(a[78]), .Z(n4118) );
  XOR U10484 ( .A(n4123), .B(n3748), .Z(n3750) );
  XOR U10485 ( .A(n4124), .B(n4125), .Z(n3748) );
  AND U10486 ( .A(n4126), .B(n4127), .Z(n4124) );
  AND U10487 ( .A(b[37]), .B(a[79]), .Z(n4123) );
  XOR U10488 ( .A(n4128), .B(n3753), .Z(n3755) );
  XOR U10489 ( .A(n4129), .B(n4130), .Z(n3753) );
  AND U10490 ( .A(n4131), .B(n4132), .Z(n4129) );
  AND U10491 ( .A(b[36]), .B(a[80]), .Z(n4128) );
  XOR U10492 ( .A(n4133), .B(n4134), .Z(n3757) );
  AND U10493 ( .A(n4135), .B(n4136), .Z(n4133) );
  XOR U10494 ( .A(n4137), .B(n3762), .Z(n3764) );
  XOR U10495 ( .A(n4138), .B(n4139), .Z(n3762) );
  AND U10496 ( .A(n4140), .B(n4141), .Z(n4138) );
  AND U10497 ( .A(b[35]), .B(a[81]), .Z(n4137) );
  XOR U10498 ( .A(n4142), .B(n3767), .Z(n3769) );
  XOR U10499 ( .A(n4143), .B(n4144), .Z(n3767) );
  AND U10500 ( .A(n4145), .B(n4146), .Z(n4143) );
  AND U10501 ( .A(b[33]), .B(a[83]), .Z(n4142) );
  XOR U10502 ( .A(n4147), .B(n3772), .Z(n3774) );
  XOR U10503 ( .A(n4148), .B(n4149), .Z(n3772) );
  AND U10504 ( .A(n4150), .B(n4151), .Z(n4148) );
  AND U10505 ( .A(b[32]), .B(a[84]), .Z(n4147) );
  XOR U10506 ( .A(n4152), .B(n3777), .Z(n3779) );
  XOR U10507 ( .A(n4153), .B(n4154), .Z(n3777) );
  AND U10508 ( .A(n4155), .B(n4156), .Z(n4153) );
  AND U10509 ( .A(b[31]), .B(a[85]), .Z(n4152) );
  XOR U10510 ( .A(n4157), .B(n3782), .Z(n3784) );
  XOR U10511 ( .A(n4158), .B(n4159), .Z(n3782) );
  AND U10512 ( .A(n4160), .B(n4161), .Z(n4158) );
  AND U10513 ( .A(b[30]), .B(a[86]), .Z(n4157) );
  XOR U10514 ( .A(n4162), .B(n4163), .Z(n3786) );
  AND U10515 ( .A(n4164), .B(n4165), .Z(n4162) );
  XOR U10516 ( .A(n4166), .B(n3791), .Z(n3793) );
  XOR U10517 ( .A(n4167), .B(n4168), .Z(n3791) );
  AND U10518 ( .A(n4169), .B(n4170), .Z(n4167) );
  AND U10519 ( .A(b[29]), .B(a[87]), .Z(n4166) );
  XOR U10520 ( .A(n4171), .B(n3796), .Z(n3798) );
  XOR U10521 ( .A(n4172), .B(n4173), .Z(n3796) );
  AND U10522 ( .A(n4174), .B(n4175), .Z(n4172) );
  AND U10523 ( .A(b[27]), .B(a[89]), .Z(n4171) );
  XOR U10524 ( .A(n4176), .B(n3801), .Z(n3803) );
  XOR U10525 ( .A(n4177), .B(n4178), .Z(n3801) );
  AND U10526 ( .A(n4179), .B(n4180), .Z(n4177) );
  AND U10527 ( .A(b[26]), .B(a[90]), .Z(n4176) );
  XOR U10528 ( .A(n4181), .B(n3806), .Z(n3808) );
  XOR U10529 ( .A(n4182), .B(n4183), .Z(n3806) );
  AND U10530 ( .A(n4184), .B(n4185), .Z(n4182) );
  AND U10531 ( .A(b[25]), .B(a[91]), .Z(n4181) );
  XOR U10532 ( .A(n4186), .B(n3811), .Z(n3813) );
  XOR U10533 ( .A(n4187), .B(n4188), .Z(n3811) );
  AND U10534 ( .A(n4189), .B(n4190), .Z(n4187) );
  AND U10535 ( .A(b[24]), .B(a[92]), .Z(n4186) );
  XOR U10536 ( .A(n4191), .B(n4192), .Z(n3815) );
  AND U10537 ( .A(n4193), .B(n4194), .Z(n4191) );
  XOR U10538 ( .A(n4195), .B(n3820), .Z(n3822) );
  XOR U10539 ( .A(n4196), .B(n4197), .Z(n3820) );
  AND U10540 ( .A(n4198), .B(n4199), .Z(n4196) );
  AND U10541 ( .A(b[23]), .B(a[93]), .Z(n4195) );
  XOR U10542 ( .A(n4200), .B(n3825), .Z(n3827) );
  XOR U10543 ( .A(n4201), .B(n4202), .Z(n3825) );
  AND U10544 ( .A(n4203), .B(n4204), .Z(n4201) );
  AND U10545 ( .A(b[21]), .B(a[95]), .Z(n4200) );
  XOR U10546 ( .A(n4205), .B(n3830), .Z(n3832) );
  XOR U10547 ( .A(n4206), .B(n4207), .Z(n3830) );
  AND U10548 ( .A(n4208), .B(n4209), .Z(n4206) );
  AND U10549 ( .A(b[20]), .B(a[96]), .Z(n4205) );
  XOR U10550 ( .A(n4210), .B(n3835), .Z(n3837) );
  XOR U10551 ( .A(n4211), .B(n4212), .Z(n3835) );
  AND U10552 ( .A(n4213), .B(n4214), .Z(n4211) );
  AND U10553 ( .A(b[19]), .B(a[97]), .Z(n4210) );
  XOR U10554 ( .A(n4215), .B(n3840), .Z(n3842) );
  XOR U10555 ( .A(n4216), .B(n4217), .Z(n3840) );
  AND U10556 ( .A(n4218), .B(n4219), .Z(n4216) );
  AND U10557 ( .A(b[18]), .B(a[98]), .Z(n4215) );
  XOR U10558 ( .A(n4220), .B(n4221), .Z(n3844) );
  AND U10559 ( .A(n4222), .B(n4223), .Z(n4220) );
  XOR U10560 ( .A(n4224), .B(n3849), .Z(n3851) );
  XOR U10561 ( .A(n4225), .B(n4226), .Z(n3849) );
  AND U10562 ( .A(n4227), .B(n4228), .Z(n4225) );
  AND U10563 ( .A(b[17]), .B(a[99]), .Z(n4224) );
  XOR U10564 ( .A(n4229), .B(n3854), .Z(n3856) );
  XOR U10565 ( .A(n4230), .B(n4231), .Z(n3854) );
  AND U10566 ( .A(n4232), .B(n4233), .Z(n4230) );
  AND U10567 ( .A(b[15]), .B(a[101]), .Z(n4229) );
  XOR U10568 ( .A(n4234), .B(n3859), .Z(n3861) );
  XOR U10569 ( .A(n4235), .B(n4236), .Z(n3859) );
  AND U10570 ( .A(n4237), .B(n4238), .Z(n4235) );
  AND U10571 ( .A(b[14]), .B(a[102]), .Z(n4234) );
  XOR U10572 ( .A(n4239), .B(n3864), .Z(n3866) );
  XOR U10573 ( .A(n4240), .B(n4241), .Z(n3864) );
  AND U10574 ( .A(n4242), .B(n4243), .Z(n4240) );
  AND U10575 ( .A(b[13]), .B(a[103]), .Z(n4239) );
  XOR U10576 ( .A(n4244), .B(n3869), .Z(n3871) );
  XOR U10577 ( .A(n4245), .B(n4246), .Z(n3869) );
  AND U10578 ( .A(n4247), .B(n4248), .Z(n4245) );
  AND U10579 ( .A(b[12]), .B(a[104]), .Z(n4244) );
  XOR U10580 ( .A(n4249), .B(n4250), .Z(n3873) );
  AND U10581 ( .A(n4251), .B(n4252), .Z(n4249) );
  XOR U10582 ( .A(n4253), .B(n3878), .Z(n3880) );
  XOR U10583 ( .A(n4254), .B(n4255), .Z(n3878) );
  AND U10584 ( .A(n4256), .B(n4257), .Z(n4254) );
  AND U10585 ( .A(b[11]), .B(a[105]), .Z(n4253) );
  XOR U10586 ( .A(n4258), .B(n3883), .Z(n3885) );
  XOR U10587 ( .A(n4259), .B(n4260), .Z(n3883) );
  AND U10588 ( .A(n4261), .B(n4262), .Z(n4259) );
  AND U10589 ( .A(b[9]), .B(a[107]), .Z(n4258) );
  XOR U10590 ( .A(n4263), .B(n3888), .Z(n3890) );
  XOR U10591 ( .A(n4264), .B(n4265), .Z(n3888) );
  AND U10592 ( .A(n4266), .B(n4267), .Z(n4264) );
  AND U10593 ( .A(b[8]), .B(a[108]), .Z(n4263) );
  XOR U10594 ( .A(n4268), .B(n3893), .Z(n3895) );
  XOR U10595 ( .A(n4269), .B(n4270), .Z(n3893) );
  AND U10596 ( .A(n4271), .B(n4272), .Z(n4269) );
  AND U10597 ( .A(b[7]), .B(a[109]), .Z(n4268) );
  XOR U10598 ( .A(n4273), .B(n3898), .Z(n3900) );
  XOR U10599 ( .A(n4274), .B(n4275), .Z(n3898) );
  AND U10600 ( .A(n4276), .B(n4277), .Z(n4274) );
  AND U10601 ( .A(b[6]), .B(a[110]), .Z(n4273) );
  XOR U10602 ( .A(n4278), .B(n3903), .Z(n3905) );
  XOR U10603 ( .A(n4279), .B(n4280), .Z(n3903) );
  AND U10604 ( .A(n4281), .B(n4282), .Z(n4279) );
  AND U10605 ( .A(b[5]), .B(a[111]), .Z(n4278) );
  XOR U10606 ( .A(n4283), .B(n3908), .Z(n3910) );
  XOR U10607 ( .A(n4284), .B(n4285), .Z(n3908) );
  AND U10608 ( .A(n4286), .B(n4287), .Z(n4284) );
  AND U10609 ( .A(b[4]), .B(a[112]), .Z(n4283) );
  XNOR U10610 ( .A(n4288), .B(n4289), .Z(n3922) );
  NANDN U10611 ( .A(n4290), .B(n4291), .Z(n4289) );
  XOR U10612 ( .A(n4292), .B(n3913), .Z(n3915) );
  XNOR U10613 ( .A(n4293), .B(n4294), .Z(n3913) );
  AND U10614 ( .A(n4295), .B(n4296), .Z(n4293) );
  AND U10615 ( .A(b[3]), .B(a[113]), .Z(n4292) );
  XOR U10616 ( .A(n4297), .B(n4298), .Z(swire[115]) );
  XOR U10617 ( .A(n3932), .B(n4299), .Z(n4298) );
  XNOR U10618 ( .A(n3931), .B(n4297), .Z(n4299) );
  NAND U10619 ( .A(a[115]), .B(b[0]), .Z(n3931) );
  XNOR U10620 ( .A(n4290), .B(n4291), .Z(n3932) );
  XOR U10621 ( .A(n4288), .B(n4300), .Z(n4291) );
  NAND U10622 ( .A(b[1]), .B(a[114]), .Z(n4300) );
  XOR U10623 ( .A(n4296), .B(n4301), .Z(n4290) );
  XOR U10624 ( .A(n4288), .B(n4295), .Z(n4301) );
  XNOR U10625 ( .A(n4302), .B(n4294), .Z(n4295) );
  AND U10626 ( .A(b[2]), .B(a[113]), .Z(n4302) );
  NANDN U10627 ( .A(n4303), .B(n4304), .Z(n4288) );
  XOR U10628 ( .A(n4294), .B(n4286), .Z(n4305) );
  XNOR U10629 ( .A(n4285), .B(n4281), .Z(n4306) );
  XNOR U10630 ( .A(n4280), .B(n4276), .Z(n4307) );
  XNOR U10631 ( .A(n4275), .B(n4271), .Z(n4308) );
  XNOR U10632 ( .A(n4270), .B(n4266), .Z(n4309) );
  XNOR U10633 ( .A(n4265), .B(n4261), .Z(n4310) );
  XNOR U10634 ( .A(n4252), .B(n4251), .Z(n4311) );
  XOR U10635 ( .A(n4312), .B(n4250), .Z(n4251) );
  AND U10636 ( .A(b[9]), .B(a[106]), .Z(n4312) );
  XNOR U10637 ( .A(n4250), .B(n4256), .Z(n4313) );
  XNOR U10638 ( .A(n4255), .B(n4247), .Z(n4314) );
  XNOR U10639 ( .A(n4246), .B(n4242), .Z(n4315) );
  XNOR U10640 ( .A(n4241), .B(n4237), .Z(n4316) );
  XNOR U10641 ( .A(n4236), .B(n4232), .Z(n4317) );
  XNOR U10642 ( .A(n4223), .B(n4222), .Z(n4318) );
  XOR U10643 ( .A(n4319), .B(n4221), .Z(n4222) );
  AND U10644 ( .A(b[15]), .B(a[100]), .Z(n4319) );
  XNOR U10645 ( .A(n4221), .B(n4227), .Z(n4320) );
  XNOR U10646 ( .A(n4226), .B(n4218), .Z(n4321) );
  XNOR U10647 ( .A(n4217), .B(n4213), .Z(n4322) );
  XNOR U10648 ( .A(n4212), .B(n4208), .Z(n4323) );
  XNOR U10649 ( .A(n4207), .B(n4203), .Z(n4324) );
  XNOR U10650 ( .A(n4194), .B(n4193), .Z(n4325) );
  XOR U10651 ( .A(n4326), .B(n4192), .Z(n4193) );
  AND U10652 ( .A(b[21]), .B(a[94]), .Z(n4326) );
  XNOR U10653 ( .A(n4192), .B(n4198), .Z(n4327) );
  XNOR U10654 ( .A(n4197), .B(n4189), .Z(n4328) );
  XNOR U10655 ( .A(n4188), .B(n4184), .Z(n4329) );
  XNOR U10656 ( .A(n4183), .B(n4179), .Z(n4330) );
  XNOR U10657 ( .A(n4178), .B(n4174), .Z(n4331) );
  XNOR U10658 ( .A(n4165), .B(n4164), .Z(n4332) );
  XOR U10659 ( .A(n4333), .B(n4163), .Z(n4164) );
  AND U10660 ( .A(b[27]), .B(a[88]), .Z(n4333) );
  XNOR U10661 ( .A(n4163), .B(n4169), .Z(n4334) );
  XNOR U10662 ( .A(n4168), .B(n4160), .Z(n4335) );
  XNOR U10663 ( .A(n4159), .B(n4155), .Z(n4336) );
  XNOR U10664 ( .A(n4154), .B(n4150), .Z(n4337) );
  XNOR U10665 ( .A(n4149), .B(n4145), .Z(n4338) );
  XNOR U10666 ( .A(n4136), .B(n4135), .Z(n4339) );
  XOR U10667 ( .A(n4340), .B(n4134), .Z(n4135) );
  AND U10668 ( .A(b[33]), .B(a[82]), .Z(n4340) );
  XNOR U10669 ( .A(n4134), .B(n4140), .Z(n4341) );
  XNOR U10670 ( .A(n4139), .B(n4131), .Z(n4342) );
  XNOR U10671 ( .A(n4130), .B(n4126), .Z(n4343) );
  XNOR U10672 ( .A(n4125), .B(n4121), .Z(n4344) );
  XNOR U10673 ( .A(n4120), .B(n4116), .Z(n4345) );
  XNOR U10674 ( .A(n4107), .B(n4106), .Z(n4346) );
  XOR U10675 ( .A(n4347), .B(n4105), .Z(n4106) );
  AND U10676 ( .A(b[39]), .B(a[76]), .Z(n4347) );
  XNOR U10677 ( .A(n4105), .B(n4111), .Z(n4348) );
  XNOR U10678 ( .A(n4110), .B(n4102), .Z(n4349) );
  XNOR U10679 ( .A(n4101), .B(n4097), .Z(n4350) );
  XNOR U10680 ( .A(n4096), .B(n4092), .Z(n4351) );
  XNOR U10681 ( .A(n4091), .B(n4087), .Z(n4352) );
  XNOR U10682 ( .A(n4078), .B(n4077), .Z(n4353) );
  XOR U10683 ( .A(n4354), .B(n4076), .Z(n4077) );
  AND U10684 ( .A(b[45]), .B(a[70]), .Z(n4354) );
  XNOR U10685 ( .A(n4076), .B(n4082), .Z(n4355) );
  XNOR U10686 ( .A(n4081), .B(n4073), .Z(n4356) );
  XNOR U10687 ( .A(n4072), .B(n4068), .Z(n4357) );
  XNOR U10688 ( .A(n4067), .B(n4063), .Z(n4358) );
  XNOR U10689 ( .A(n4062), .B(n4058), .Z(n4359) );
  XNOR U10690 ( .A(n4057), .B(n4053), .Z(n4360) );
  XNOR U10691 ( .A(n4052), .B(n4048), .Z(n4361) );
  XNOR U10692 ( .A(n4047), .B(n4043), .Z(n4362) );
  XNOR U10693 ( .A(n4042), .B(n4038), .Z(n4363) );
  XNOR U10694 ( .A(n4037), .B(n4033), .Z(n4364) );
  XNOR U10695 ( .A(n4032), .B(n4028), .Z(n4365) );
  XNOR U10696 ( .A(n4027), .B(n4023), .Z(n4366) );
  XNOR U10697 ( .A(n4022), .B(n4018), .Z(n4367) );
  XNOR U10698 ( .A(n4017), .B(n4013), .Z(n4368) );
  XOR U10699 ( .A(n4012), .B(n4009), .Z(n4369) );
  XOR U10700 ( .A(n4370), .B(n4371), .Z(n4009) );
  XOR U10701 ( .A(n4007), .B(n4372), .Z(n4371) );
  XOR U10702 ( .A(n4373), .B(n4374), .Z(n4372) );
  XOR U10703 ( .A(n4375), .B(n4376), .Z(n4374) );
  NAND U10704 ( .A(a[53]), .B(b[62]), .Z(n4376) );
  AND U10705 ( .A(a[52]), .B(b[63]), .Z(n4375) );
  XOR U10706 ( .A(n4377), .B(n4373), .Z(n4370) );
  XOR U10707 ( .A(n4378), .B(n4379), .Z(n4373) );
  ANDN U10708 ( .B(n4380), .A(n4381), .Z(n4378) );
  AND U10709 ( .A(a[54]), .B(b[61]), .Z(n4377) );
  XOR U10710 ( .A(n4382), .B(n4007), .Z(n4008) );
  XOR U10711 ( .A(n4383), .B(n4384), .Z(n4007) );
  AND U10712 ( .A(n4385), .B(n4386), .Z(n4383) );
  AND U10713 ( .A(a[55]), .B(b[60]), .Z(n4382) );
  XOR U10714 ( .A(n4387), .B(n4012), .Z(n4014) );
  XOR U10715 ( .A(n4388), .B(n4389), .Z(n4012) );
  AND U10716 ( .A(n4390), .B(n4391), .Z(n4388) );
  AND U10717 ( .A(a[56]), .B(b[59]), .Z(n4387) );
  XOR U10718 ( .A(n4392), .B(n4017), .Z(n4019) );
  XOR U10719 ( .A(n4393), .B(n4394), .Z(n4017) );
  AND U10720 ( .A(n4395), .B(n4396), .Z(n4393) );
  AND U10721 ( .A(a[57]), .B(b[58]), .Z(n4392) );
  XOR U10722 ( .A(n4397), .B(n4022), .Z(n4024) );
  XOR U10723 ( .A(n4398), .B(n4399), .Z(n4022) );
  AND U10724 ( .A(n4400), .B(n4401), .Z(n4398) );
  AND U10725 ( .A(b[57]), .B(a[58]), .Z(n4397) );
  XOR U10726 ( .A(n4402), .B(n4027), .Z(n4029) );
  XOR U10727 ( .A(n4403), .B(n4404), .Z(n4027) );
  AND U10728 ( .A(n4405), .B(n4406), .Z(n4403) );
  AND U10729 ( .A(b[56]), .B(a[59]), .Z(n4402) );
  XOR U10730 ( .A(n4407), .B(n4032), .Z(n4034) );
  XOR U10731 ( .A(n4408), .B(n4409), .Z(n4032) );
  AND U10732 ( .A(n4410), .B(n4411), .Z(n4408) );
  AND U10733 ( .A(b[55]), .B(a[60]), .Z(n4407) );
  XOR U10734 ( .A(n4412), .B(n4037), .Z(n4039) );
  XOR U10735 ( .A(n4413), .B(n4414), .Z(n4037) );
  AND U10736 ( .A(n4415), .B(n4416), .Z(n4413) );
  AND U10737 ( .A(b[54]), .B(a[61]), .Z(n4412) );
  XOR U10738 ( .A(n4417), .B(n4042), .Z(n4044) );
  XOR U10739 ( .A(n4418), .B(n4419), .Z(n4042) );
  AND U10740 ( .A(n4420), .B(n4421), .Z(n4418) );
  AND U10741 ( .A(b[53]), .B(a[62]), .Z(n4417) );
  XOR U10742 ( .A(n4422), .B(n4047), .Z(n4049) );
  XOR U10743 ( .A(n4423), .B(n4424), .Z(n4047) );
  AND U10744 ( .A(n4425), .B(n4426), .Z(n4423) );
  AND U10745 ( .A(b[52]), .B(a[63]), .Z(n4422) );
  XOR U10746 ( .A(n4427), .B(n4052), .Z(n4054) );
  XOR U10747 ( .A(n4428), .B(n4429), .Z(n4052) );
  AND U10748 ( .A(n4430), .B(n4431), .Z(n4428) );
  AND U10749 ( .A(b[51]), .B(a[64]), .Z(n4427) );
  XOR U10750 ( .A(n4432), .B(n4057), .Z(n4059) );
  XOR U10751 ( .A(n4433), .B(n4434), .Z(n4057) );
  AND U10752 ( .A(n4435), .B(n4436), .Z(n4433) );
  AND U10753 ( .A(b[50]), .B(a[65]), .Z(n4432) );
  XOR U10754 ( .A(n4437), .B(n4062), .Z(n4064) );
  XOR U10755 ( .A(n4438), .B(n4439), .Z(n4062) );
  AND U10756 ( .A(n4440), .B(n4441), .Z(n4438) );
  AND U10757 ( .A(b[49]), .B(a[66]), .Z(n4437) );
  XOR U10758 ( .A(n4442), .B(n4067), .Z(n4069) );
  XOR U10759 ( .A(n4443), .B(n4444), .Z(n4067) );
  AND U10760 ( .A(n4445), .B(n4446), .Z(n4443) );
  AND U10761 ( .A(b[48]), .B(a[67]), .Z(n4442) );
  XOR U10762 ( .A(n4447), .B(n4072), .Z(n4074) );
  XOR U10763 ( .A(n4448), .B(n4449), .Z(n4072) );
  AND U10764 ( .A(n4450), .B(n4451), .Z(n4448) );
  AND U10765 ( .A(b[47]), .B(a[68]), .Z(n4447) );
  XOR U10766 ( .A(n4452), .B(n4453), .Z(n4076) );
  AND U10767 ( .A(n4454), .B(n4455), .Z(n4452) );
  XOR U10768 ( .A(n4456), .B(n4081), .Z(n4083) );
  XOR U10769 ( .A(n4457), .B(n4458), .Z(n4081) );
  AND U10770 ( .A(n4459), .B(n4460), .Z(n4457) );
  AND U10771 ( .A(b[46]), .B(a[69]), .Z(n4456) );
  XOR U10772 ( .A(n4461), .B(n4086), .Z(n4088) );
  XOR U10773 ( .A(n4462), .B(n4463), .Z(n4086) );
  AND U10774 ( .A(n4464), .B(n4465), .Z(n4462) );
  AND U10775 ( .A(b[44]), .B(a[71]), .Z(n4461) );
  XOR U10776 ( .A(n4466), .B(n4091), .Z(n4093) );
  XOR U10777 ( .A(n4467), .B(n4468), .Z(n4091) );
  AND U10778 ( .A(n4469), .B(n4470), .Z(n4467) );
  AND U10779 ( .A(b[43]), .B(a[72]), .Z(n4466) );
  XOR U10780 ( .A(n4471), .B(n4096), .Z(n4098) );
  XOR U10781 ( .A(n4472), .B(n4473), .Z(n4096) );
  AND U10782 ( .A(n4474), .B(n4475), .Z(n4472) );
  AND U10783 ( .A(b[42]), .B(a[73]), .Z(n4471) );
  XOR U10784 ( .A(n4476), .B(n4101), .Z(n4103) );
  XOR U10785 ( .A(n4477), .B(n4478), .Z(n4101) );
  AND U10786 ( .A(n4479), .B(n4480), .Z(n4477) );
  AND U10787 ( .A(b[41]), .B(a[74]), .Z(n4476) );
  XOR U10788 ( .A(n4481), .B(n4482), .Z(n4105) );
  AND U10789 ( .A(n4483), .B(n4484), .Z(n4481) );
  XOR U10790 ( .A(n4485), .B(n4110), .Z(n4112) );
  XOR U10791 ( .A(n4486), .B(n4487), .Z(n4110) );
  AND U10792 ( .A(n4488), .B(n4489), .Z(n4486) );
  AND U10793 ( .A(b[40]), .B(a[75]), .Z(n4485) );
  XOR U10794 ( .A(n4490), .B(n4115), .Z(n4117) );
  XOR U10795 ( .A(n4491), .B(n4492), .Z(n4115) );
  AND U10796 ( .A(n4493), .B(n4494), .Z(n4491) );
  AND U10797 ( .A(b[38]), .B(a[77]), .Z(n4490) );
  XOR U10798 ( .A(n4495), .B(n4120), .Z(n4122) );
  XOR U10799 ( .A(n4496), .B(n4497), .Z(n4120) );
  AND U10800 ( .A(n4498), .B(n4499), .Z(n4496) );
  AND U10801 ( .A(b[37]), .B(a[78]), .Z(n4495) );
  XOR U10802 ( .A(n4500), .B(n4125), .Z(n4127) );
  XOR U10803 ( .A(n4501), .B(n4502), .Z(n4125) );
  AND U10804 ( .A(n4503), .B(n4504), .Z(n4501) );
  AND U10805 ( .A(b[36]), .B(a[79]), .Z(n4500) );
  XOR U10806 ( .A(n4505), .B(n4130), .Z(n4132) );
  XOR U10807 ( .A(n4506), .B(n4507), .Z(n4130) );
  AND U10808 ( .A(n4508), .B(n4509), .Z(n4506) );
  AND U10809 ( .A(b[35]), .B(a[80]), .Z(n4505) );
  XOR U10810 ( .A(n4510), .B(n4511), .Z(n4134) );
  AND U10811 ( .A(n4512), .B(n4513), .Z(n4510) );
  XOR U10812 ( .A(n4514), .B(n4139), .Z(n4141) );
  XOR U10813 ( .A(n4515), .B(n4516), .Z(n4139) );
  AND U10814 ( .A(n4517), .B(n4518), .Z(n4515) );
  AND U10815 ( .A(b[34]), .B(a[81]), .Z(n4514) );
  XOR U10816 ( .A(n4519), .B(n4144), .Z(n4146) );
  XOR U10817 ( .A(n4520), .B(n4521), .Z(n4144) );
  AND U10818 ( .A(n4522), .B(n4523), .Z(n4520) );
  AND U10819 ( .A(b[32]), .B(a[83]), .Z(n4519) );
  XOR U10820 ( .A(n4524), .B(n4149), .Z(n4151) );
  XOR U10821 ( .A(n4525), .B(n4526), .Z(n4149) );
  AND U10822 ( .A(n4527), .B(n4528), .Z(n4525) );
  AND U10823 ( .A(b[31]), .B(a[84]), .Z(n4524) );
  XOR U10824 ( .A(n4529), .B(n4154), .Z(n4156) );
  XOR U10825 ( .A(n4530), .B(n4531), .Z(n4154) );
  AND U10826 ( .A(n4532), .B(n4533), .Z(n4530) );
  AND U10827 ( .A(b[30]), .B(a[85]), .Z(n4529) );
  XOR U10828 ( .A(n4534), .B(n4159), .Z(n4161) );
  XOR U10829 ( .A(n4535), .B(n4536), .Z(n4159) );
  AND U10830 ( .A(n4537), .B(n4538), .Z(n4535) );
  AND U10831 ( .A(b[29]), .B(a[86]), .Z(n4534) );
  XOR U10832 ( .A(n4539), .B(n4540), .Z(n4163) );
  AND U10833 ( .A(n4541), .B(n4542), .Z(n4539) );
  XOR U10834 ( .A(n4543), .B(n4168), .Z(n4170) );
  XOR U10835 ( .A(n4544), .B(n4545), .Z(n4168) );
  AND U10836 ( .A(n4546), .B(n4547), .Z(n4544) );
  AND U10837 ( .A(b[28]), .B(a[87]), .Z(n4543) );
  XOR U10838 ( .A(n4548), .B(n4173), .Z(n4175) );
  XOR U10839 ( .A(n4549), .B(n4550), .Z(n4173) );
  AND U10840 ( .A(n4551), .B(n4552), .Z(n4549) );
  AND U10841 ( .A(b[26]), .B(a[89]), .Z(n4548) );
  XOR U10842 ( .A(n4553), .B(n4178), .Z(n4180) );
  XOR U10843 ( .A(n4554), .B(n4555), .Z(n4178) );
  AND U10844 ( .A(n4556), .B(n4557), .Z(n4554) );
  AND U10845 ( .A(b[25]), .B(a[90]), .Z(n4553) );
  XOR U10846 ( .A(n4558), .B(n4183), .Z(n4185) );
  XOR U10847 ( .A(n4559), .B(n4560), .Z(n4183) );
  AND U10848 ( .A(n4561), .B(n4562), .Z(n4559) );
  AND U10849 ( .A(b[24]), .B(a[91]), .Z(n4558) );
  XOR U10850 ( .A(n4563), .B(n4188), .Z(n4190) );
  XOR U10851 ( .A(n4564), .B(n4565), .Z(n4188) );
  AND U10852 ( .A(n4566), .B(n4567), .Z(n4564) );
  AND U10853 ( .A(b[23]), .B(a[92]), .Z(n4563) );
  XOR U10854 ( .A(n4568), .B(n4569), .Z(n4192) );
  AND U10855 ( .A(n4570), .B(n4571), .Z(n4568) );
  XOR U10856 ( .A(n4572), .B(n4197), .Z(n4199) );
  XOR U10857 ( .A(n4573), .B(n4574), .Z(n4197) );
  AND U10858 ( .A(n4575), .B(n4576), .Z(n4573) );
  AND U10859 ( .A(b[22]), .B(a[93]), .Z(n4572) );
  XOR U10860 ( .A(n4577), .B(n4202), .Z(n4204) );
  XOR U10861 ( .A(n4578), .B(n4579), .Z(n4202) );
  AND U10862 ( .A(n4580), .B(n4581), .Z(n4578) );
  AND U10863 ( .A(b[20]), .B(a[95]), .Z(n4577) );
  XOR U10864 ( .A(n4582), .B(n4207), .Z(n4209) );
  XOR U10865 ( .A(n4583), .B(n4584), .Z(n4207) );
  AND U10866 ( .A(n4585), .B(n4586), .Z(n4583) );
  AND U10867 ( .A(b[19]), .B(a[96]), .Z(n4582) );
  XOR U10868 ( .A(n4587), .B(n4212), .Z(n4214) );
  XOR U10869 ( .A(n4588), .B(n4589), .Z(n4212) );
  AND U10870 ( .A(n4590), .B(n4591), .Z(n4588) );
  AND U10871 ( .A(b[18]), .B(a[97]), .Z(n4587) );
  XOR U10872 ( .A(n4592), .B(n4217), .Z(n4219) );
  XOR U10873 ( .A(n4593), .B(n4594), .Z(n4217) );
  AND U10874 ( .A(n4595), .B(n4596), .Z(n4593) );
  AND U10875 ( .A(b[17]), .B(a[98]), .Z(n4592) );
  XOR U10876 ( .A(n4597), .B(n4598), .Z(n4221) );
  AND U10877 ( .A(n4599), .B(n4600), .Z(n4597) );
  XOR U10878 ( .A(n4601), .B(n4226), .Z(n4228) );
  XOR U10879 ( .A(n4602), .B(n4603), .Z(n4226) );
  AND U10880 ( .A(n4604), .B(n4605), .Z(n4602) );
  AND U10881 ( .A(b[16]), .B(a[99]), .Z(n4601) );
  XOR U10882 ( .A(n4606), .B(n4231), .Z(n4233) );
  XOR U10883 ( .A(n4607), .B(n4608), .Z(n4231) );
  AND U10884 ( .A(n4609), .B(n4610), .Z(n4607) );
  AND U10885 ( .A(b[14]), .B(a[101]), .Z(n4606) );
  XOR U10886 ( .A(n4611), .B(n4236), .Z(n4238) );
  XOR U10887 ( .A(n4612), .B(n4613), .Z(n4236) );
  AND U10888 ( .A(n4614), .B(n4615), .Z(n4612) );
  AND U10889 ( .A(b[13]), .B(a[102]), .Z(n4611) );
  XOR U10890 ( .A(n4616), .B(n4241), .Z(n4243) );
  XOR U10891 ( .A(n4617), .B(n4618), .Z(n4241) );
  AND U10892 ( .A(n4619), .B(n4620), .Z(n4617) );
  AND U10893 ( .A(b[12]), .B(a[103]), .Z(n4616) );
  XOR U10894 ( .A(n4621), .B(n4246), .Z(n4248) );
  XOR U10895 ( .A(n4622), .B(n4623), .Z(n4246) );
  AND U10896 ( .A(n4624), .B(n4625), .Z(n4622) );
  AND U10897 ( .A(b[11]), .B(a[104]), .Z(n4621) );
  XOR U10898 ( .A(n4626), .B(n4627), .Z(n4250) );
  AND U10899 ( .A(n4628), .B(n4629), .Z(n4626) );
  XOR U10900 ( .A(n4630), .B(n4255), .Z(n4257) );
  XOR U10901 ( .A(n4631), .B(n4632), .Z(n4255) );
  AND U10902 ( .A(n4633), .B(n4634), .Z(n4631) );
  AND U10903 ( .A(b[10]), .B(a[105]), .Z(n4630) );
  XOR U10904 ( .A(n4635), .B(n4260), .Z(n4262) );
  XOR U10905 ( .A(n4636), .B(n4637), .Z(n4260) );
  AND U10906 ( .A(n4638), .B(n4639), .Z(n4636) );
  AND U10907 ( .A(b[8]), .B(a[107]), .Z(n4635) );
  XOR U10908 ( .A(n4640), .B(n4265), .Z(n4267) );
  XOR U10909 ( .A(n4641), .B(n4642), .Z(n4265) );
  AND U10910 ( .A(n4643), .B(n4644), .Z(n4641) );
  AND U10911 ( .A(b[7]), .B(a[108]), .Z(n4640) );
  XOR U10912 ( .A(n4645), .B(n4270), .Z(n4272) );
  XOR U10913 ( .A(n4646), .B(n4647), .Z(n4270) );
  AND U10914 ( .A(n4648), .B(n4649), .Z(n4646) );
  AND U10915 ( .A(b[6]), .B(a[109]), .Z(n4645) );
  XOR U10916 ( .A(n4650), .B(n4275), .Z(n4277) );
  XOR U10917 ( .A(n4651), .B(n4652), .Z(n4275) );
  AND U10918 ( .A(n4653), .B(n4654), .Z(n4651) );
  AND U10919 ( .A(b[5]), .B(a[110]), .Z(n4650) );
  XOR U10920 ( .A(n4655), .B(n4280), .Z(n4282) );
  XOR U10921 ( .A(n4656), .B(n4657), .Z(n4280) );
  AND U10922 ( .A(n4658), .B(n4659), .Z(n4656) );
  AND U10923 ( .A(b[4]), .B(a[111]), .Z(n4655) );
  XNOR U10924 ( .A(n4660), .B(n4661), .Z(n4294) );
  NANDN U10925 ( .A(n4662), .B(n4663), .Z(n4661) );
  XOR U10926 ( .A(n4664), .B(n4285), .Z(n4287) );
  XNOR U10927 ( .A(n4665), .B(n4666), .Z(n4285) );
  AND U10928 ( .A(n4667), .B(n4668), .Z(n4665) );
  AND U10929 ( .A(b[3]), .B(a[112]), .Z(n4664) );
  XOR U10930 ( .A(n4669), .B(n4670), .Z(swire[114]) );
  XOR U10931 ( .A(n4304), .B(n4671), .Z(n4670) );
  XNOR U10932 ( .A(n4303), .B(n4669), .Z(n4671) );
  NAND U10933 ( .A(a[114]), .B(b[0]), .Z(n4303) );
  XNOR U10934 ( .A(n4662), .B(n4663), .Z(n4304) );
  XOR U10935 ( .A(n4660), .B(n4672), .Z(n4663) );
  NAND U10936 ( .A(b[1]), .B(a[113]), .Z(n4672) );
  XOR U10937 ( .A(n4667), .B(n4673), .Z(n4662) );
  XOR U10938 ( .A(n4660), .B(n4668), .Z(n4673) );
  XNOR U10939 ( .A(n4674), .B(n4666), .Z(n4668) );
  AND U10940 ( .A(b[2]), .B(a[112]), .Z(n4674) );
  NANDN U10941 ( .A(n4675), .B(n4676), .Z(n4660) );
  XOR U10942 ( .A(n4666), .B(n4658), .Z(n4677) );
  XNOR U10943 ( .A(n4657), .B(n4653), .Z(n4678) );
  XNOR U10944 ( .A(n4652), .B(n4648), .Z(n4679) );
  XNOR U10945 ( .A(n4647), .B(n4643), .Z(n4680) );
  XNOR U10946 ( .A(n4642), .B(n4638), .Z(n4681) );
  XNOR U10947 ( .A(n4629), .B(n4628), .Z(n4682) );
  XOR U10948 ( .A(n4683), .B(n4627), .Z(n4628) );
  AND U10949 ( .A(b[8]), .B(a[106]), .Z(n4683) );
  XNOR U10950 ( .A(n4627), .B(n4633), .Z(n4684) );
  XNOR U10951 ( .A(n4632), .B(n4624), .Z(n4685) );
  XNOR U10952 ( .A(n4623), .B(n4619), .Z(n4686) );
  XNOR U10953 ( .A(n4618), .B(n4614), .Z(n4687) );
  XNOR U10954 ( .A(n4613), .B(n4609), .Z(n4688) );
  XNOR U10955 ( .A(n4600), .B(n4599), .Z(n4689) );
  XOR U10956 ( .A(n4690), .B(n4598), .Z(n4599) );
  AND U10957 ( .A(b[14]), .B(a[100]), .Z(n4690) );
  XNOR U10958 ( .A(n4598), .B(n4604), .Z(n4691) );
  XNOR U10959 ( .A(n4603), .B(n4595), .Z(n4692) );
  XNOR U10960 ( .A(n4594), .B(n4590), .Z(n4693) );
  XNOR U10961 ( .A(n4589), .B(n4585), .Z(n4694) );
  XNOR U10962 ( .A(n4584), .B(n4580), .Z(n4695) );
  XNOR U10963 ( .A(n4571), .B(n4570), .Z(n4696) );
  XOR U10964 ( .A(n4697), .B(n4569), .Z(n4570) );
  AND U10965 ( .A(b[20]), .B(a[94]), .Z(n4697) );
  XNOR U10966 ( .A(n4569), .B(n4575), .Z(n4698) );
  XNOR U10967 ( .A(n4574), .B(n4566), .Z(n4699) );
  XNOR U10968 ( .A(n4565), .B(n4561), .Z(n4700) );
  XNOR U10969 ( .A(n4560), .B(n4556), .Z(n4701) );
  XNOR U10970 ( .A(n4555), .B(n4551), .Z(n4702) );
  XNOR U10971 ( .A(n4542), .B(n4541), .Z(n4703) );
  XOR U10972 ( .A(n4704), .B(n4540), .Z(n4541) );
  AND U10973 ( .A(b[26]), .B(a[88]), .Z(n4704) );
  XNOR U10974 ( .A(n4540), .B(n4546), .Z(n4705) );
  XNOR U10975 ( .A(n4545), .B(n4537), .Z(n4706) );
  XNOR U10976 ( .A(n4536), .B(n4532), .Z(n4707) );
  XNOR U10977 ( .A(n4531), .B(n4527), .Z(n4708) );
  XNOR U10978 ( .A(n4526), .B(n4522), .Z(n4709) );
  XNOR U10979 ( .A(n4513), .B(n4512), .Z(n4710) );
  XOR U10980 ( .A(n4711), .B(n4511), .Z(n4512) );
  AND U10981 ( .A(b[32]), .B(a[82]), .Z(n4711) );
  XNOR U10982 ( .A(n4511), .B(n4517), .Z(n4712) );
  XNOR U10983 ( .A(n4516), .B(n4508), .Z(n4713) );
  XNOR U10984 ( .A(n4507), .B(n4503), .Z(n4714) );
  XNOR U10985 ( .A(n4502), .B(n4498), .Z(n4715) );
  XNOR U10986 ( .A(n4497), .B(n4493), .Z(n4716) );
  XNOR U10987 ( .A(n4484), .B(n4483), .Z(n4717) );
  XOR U10988 ( .A(n4718), .B(n4482), .Z(n4483) );
  AND U10989 ( .A(b[38]), .B(a[76]), .Z(n4718) );
  XNOR U10990 ( .A(n4482), .B(n4488), .Z(n4719) );
  XNOR U10991 ( .A(n4487), .B(n4479), .Z(n4720) );
  XNOR U10992 ( .A(n4478), .B(n4474), .Z(n4721) );
  XNOR U10993 ( .A(n4473), .B(n4469), .Z(n4722) );
  XNOR U10994 ( .A(n4468), .B(n4464), .Z(n4723) );
  XNOR U10995 ( .A(n4455), .B(n4454), .Z(n4724) );
  XOR U10996 ( .A(n4725), .B(n4453), .Z(n4454) );
  AND U10997 ( .A(b[44]), .B(a[70]), .Z(n4725) );
  XNOR U10998 ( .A(n4453), .B(n4459), .Z(n4726) );
  XNOR U10999 ( .A(n4458), .B(n4450), .Z(n4727) );
  XNOR U11000 ( .A(n4449), .B(n4445), .Z(n4728) );
  XNOR U11001 ( .A(n4444), .B(n4440), .Z(n4729) );
  XNOR U11002 ( .A(n4439), .B(n4435), .Z(n4730) );
  XNOR U11003 ( .A(n4434), .B(n4430), .Z(n4731) );
  XNOR U11004 ( .A(n4429), .B(n4425), .Z(n4732) );
  XNOR U11005 ( .A(n4424), .B(n4420), .Z(n4733) );
  XNOR U11006 ( .A(n4419), .B(n4415), .Z(n4734) );
  XNOR U11007 ( .A(n4414), .B(n4410), .Z(n4735) );
  XNOR U11008 ( .A(n4409), .B(n4405), .Z(n4736) );
  XNOR U11009 ( .A(n4404), .B(n4400), .Z(n4737) );
  XNOR U11010 ( .A(n4399), .B(n4395), .Z(n4738) );
  XNOR U11011 ( .A(n4394), .B(n4390), .Z(n4739) );
  XNOR U11012 ( .A(n4389), .B(n4385), .Z(n4740) );
  XOR U11013 ( .A(n4384), .B(n4381), .Z(n4741) );
  XOR U11014 ( .A(n4742), .B(n4743), .Z(n4381) );
  XOR U11015 ( .A(n4379), .B(n4744), .Z(n4743) );
  XOR U11016 ( .A(n4745), .B(n4746), .Z(n4744) );
  XOR U11017 ( .A(n4747), .B(n4748), .Z(n4746) );
  NAND U11018 ( .A(a[52]), .B(b[62]), .Z(n4748) );
  AND U11019 ( .A(a[51]), .B(b[63]), .Z(n4747) );
  XOR U11020 ( .A(n4749), .B(n4745), .Z(n4742) );
  XOR U11021 ( .A(n4750), .B(n4751), .Z(n4745) );
  ANDN U11022 ( .B(n4752), .A(n4753), .Z(n4750) );
  AND U11023 ( .A(a[53]), .B(b[61]), .Z(n4749) );
  XOR U11024 ( .A(n4754), .B(n4379), .Z(n4380) );
  XOR U11025 ( .A(n4755), .B(n4756), .Z(n4379) );
  AND U11026 ( .A(n4757), .B(n4758), .Z(n4755) );
  AND U11027 ( .A(a[54]), .B(b[60]), .Z(n4754) );
  XOR U11028 ( .A(n4759), .B(n4384), .Z(n4386) );
  XOR U11029 ( .A(n4760), .B(n4761), .Z(n4384) );
  AND U11030 ( .A(n4762), .B(n4763), .Z(n4760) );
  AND U11031 ( .A(a[55]), .B(b[59]), .Z(n4759) );
  XOR U11032 ( .A(n4764), .B(n4389), .Z(n4391) );
  XOR U11033 ( .A(n4765), .B(n4766), .Z(n4389) );
  AND U11034 ( .A(n4767), .B(n4768), .Z(n4765) );
  AND U11035 ( .A(a[56]), .B(b[58]), .Z(n4764) );
  XOR U11036 ( .A(n4769), .B(n4394), .Z(n4396) );
  XOR U11037 ( .A(n4770), .B(n4771), .Z(n4394) );
  AND U11038 ( .A(n4772), .B(n4773), .Z(n4770) );
  AND U11039 ( .A(a[57]), .B(b[57]), .Z(n4769) );
  XOR U11040 ( .A(n4774), .B(n4399), .Z(n4401) );
  XOR U11041 ( .A(n4775), .B(n4776), .Z(n4399) );
  AND U11042 ( .A(n4777), .B(n4778), .Z(n4775) );
  AND U11043 ( .A(b[56]), .B(a[58]), .Z(n4774) );
  XOR U11044 ( .A(n4779), .B(n4404), .Z(n4406) );
  XOR U11045 ( .A(n4780), .B(n4781), .Z(n4404) );
  AND U11046 ( .A(n4782), .B(n4783), .Z(n4780) );
  AND U11047 ( .A(b[55]), .B(a[59]), .Z(n4779) );
  XOR U11048 ( .A(n4784), .B(n4409), .Z(n4411) );
  XOR U11049 ( .A(n4785), .B(n4786), .Z(n4409) );
  AND U11050 ( .A(n4787), .B(n4788), .Z(n4785) );
  AND U11051 ( .A(b[54]), .B(a[60]), .Z(n4784) );
  XOR U11052 ( .A(n4789), .B(n4414), .Z(n4416) );
  XOR U11053 ( .A(n4790), .B(n4791), .Z(n4414) );
  AND U11054 ( .A(n4792), .B(n4793), .Z(n4790) );
  AND U11055 ( .A(b[53]), .B(a[61]), .Z(n4789) );
  XOR U11056 ( .A(n4794), .B(n4419), .Z(n4421) );
  XOR U11057 ( .A(n4795), .B(n4796), .Z(n4419) );
  AND U11058 ( .A(n4797), .B(n4798), .Z(n4795) );
  AND U11059 ( .A(b[52]), .B(a[62]), .Z(n4794) );
  XOR U11060 ( .A(n4799), .B(n4424), .Z(n4426) );
  XOR U11061 ( .A(n4800), .B(n4801), .Z(n4424) );
  AND U11062 ( .A(n4802), .B(n4803), .Z(n4800) );
  AND U11063 ( .A(b[51]), .B(a[63]), .Z(n4799) );
  XOR U11064 ( .A(n4804), .B(n4429), .Z(n4431) );
  XOR U11065 ( .A(n4805), .B(n4806), .Z(n4429) );
  AND U11066 ( .A(n4807), .B(n4808), .Z(n4805) );
  AND U11067 ( .A(b[50]), .B(a[64]), .Z(n4804) );
  XOR U11068 ( .A(n4809), .B(n4434), .Z(n4436) );
  XOR U11069 ( .A(n4810), .B(n4811), .Z(n4434) );
  AND U11070 ( .A(n4812), .B(n4813), .Z(n4810) );
  AND U11071 ( .A(b[49]), .B(a[65]), .Z(n4809) );
  XOR U11072 ( .A(n4814), .B(n4439), .Z(n4441) );
  XOR U11073 ( .A(n4815), .B(n4816), .Z(n4439) );
  AND U11074 ( .A(n4817), .B(n4818), .Z(n4815) );
  AND U11075 ( .A(b[48]), .B(a[66]), .Z(n4814) );
  XOR U11076 ( .A(n4819), .B(n4444), .Z(n4446) );
  XOR U11077 ( .A(n4820), .B(n4821), .Z(n4444) );
  AND U11078 ( .A(n4822), .B(n4823), .Z(n4820) );
  AND U11079 ( .A(b[47]), .B(a[67]), .Z(n4819) );
  XOR U11080 ( .A(n4824), .B(n4449), .Z(n4451) );
  XOR U11081 ( .A(n4825), .B(n4826), .Z(n4449) );
  AND U11082 ( .A(n4827), .B(n4828), .Z(n4825) );
  AND U11083 ( .A(b[46]), .B(a[68]), .Z(n4824) );
  XOR U11084 ( .A(n4829), .B(n4830), .Z(n4453) );
  AND U11085 ( .A(n4831), .B(n4832), .Z(n4829) );
  XOR U11086 ( .A(n4833), .B(n4458), .Z(n4460) );
  XOR U11087 ( .A(n4834), .B(n4835), .Z(n4458) );
  AND U11088 ( .A(n4836), .B(n4837), .Z(n4834) );
  AND U11089 ( .A(b[45]), .B(a[69]), .Z(n4833) );
  XOR U11090 ( .A(n4838), .B(n4463), .Z(n4465) );
  XOR U11091 ( .A(n4839), .B(n4840), .Z(n4463) );
  AND U11092 ( .A(n4841), .B(n4842), .Z(n4839) );
  AND U11093 ( .A(b[43]), .B(a[71]), .Z(n4838) );
  XOR U11094 ( .A(n4843), .B(n4468), .Z(n4470) );
  XOR U11095 ( .A(n4844), .B(n4845), .Z(n4468) );
  AND U11096 ( .A(n4846), .B(n4847), .Z(n4844) );
  AND U11097 ( .A(b[42]), .B(a[72]), .Z(n4843) );
  XOR U11098 ( .A(n4848), .B(n4473), .Z(n4475) );
  XOR U11099 ( .A(n4849), .B(n4850), .Z(n4473) );
  AND U11100 ( .A(n4851), .B(n4852), .Z(n4849) );
  AND U11101 ( .A(b[41]), .B(a[73]), .Z(n4848) );
  XOR U11102 ( .A(n4853), .B(n4478), .Z(n4480) );
  XOR U11103 ( .A(n4854), .B(n4855), .Z(n4478) );
  AND U11104 ( .A(n4856), .B(n4857), .Z(n4854) );
  AND U11105 ( .A(b[40]), .B(a[74]), .Z(n4853) );
  XOR U11106 ( .A(n4858), .B(n4859), .Z(n4482) );
  AND U11107 ( .A(n4860), .B(n4861), .Z(n4858) );
  XOR U11108 ( .A(n4862), .B(n4487), .Z(n4489) );
  XOR U11109 ( .A(n4863), .B(n4864), .Z(n4487) );
  AND U11110 ( .A(n4865), .B(n4866), .Z(n4863) );
  AND U11111 ( .A(b[39]), .B(a[75]), .Z(n4862) );
  XOR U11112 ( .A(n4867), .B(n4492), .Z(n4494) );
  XOR U11113 ( .A(n4868), .B(n4869), .Z(n4492) );
  AND U11114 ( .A(n4870), .B(n4871), .Z(n4868) );
  AND U11115 ( .A(b[37]), .B(a[77]), .Z(n4867) );
  XOR U11116 ( .A(n4872), .B(n4497), .Z(n4499) );
  XOR U11117 ( .A(n4873), .B(n4874), .Z(n4497) );
  AND U11118 ( .A(n4875), .B(n4876), .Z(n4873) );
  AND U11119 ( .A(b[36]), .B(a[78]), .Z(n4872) );
  XOR U11120 ( .A(n4877), .B(n4502), .Z(n4504) );
  XOR U11121 ( .A(n4878), .B(n4879), .Z(n4502) );
  AND U11122 ( .A(n4880), .B(n4881), .Z(n4878) );
  AND U11123 ( .A(b[35]), .B(a[79]), .Z(n4877) );
  XOR U11124 ( .A(n4882), .B(n4507), .Z(n4509) );
  XOR U11125 ( .A(n4883), .B(n4884), .Z(n4507) );
  AND U11126 ( .A(n4885), .B(n4886), .Z(n4883) );
  AND U11127 ( .A(b[34]), .B(a[80]), .Z(n4882) );
  XOR U11128 ( .A(n4887), .B(n4888), .Z(n4511) );
  AND U11129 ( .A(n4889), .B(n4890), .Z(n4887) );
  XOR U11130 ( .A(n4891), .B(n4516), .Z(n4518) );
  XOR U11131 ( .A(n4892), .B(n4893), .Z(n4516) );
  AND U11132 ( .A(n4894), .B(n4895), .Z(n4892) );
  AND U11133 ( .A(b[33]), .B(a[81]), .Z(n4891) );
  XOR U11134 ( .A(n4896), .B(n4521), .Z(n4523) );
  XOR U11135 ( .A(n4897), .B(n4898), .Z(n4521) );
  AND U11136 ( .A(n4899), .B(n4900), .Z(n4897) );
  AND U11137 ( .A(b[31]), .B(a[83]), .Z(n4896) );
  XOR U11138 ( .A(n4901), .B(n4526), .Z(n4528) );
  XOR U11139 ( .A(n4902), .B(n4903), .Z(n4526) );
  AND U11140 ( .A(n4904), .B(n4905), .Z(n4902) );
  AND U11141 ( .A(b[30]), .B(a[84]), .Z(n4901) );
  XOR U11142 ( .A(n4906), .B(n4531), .Z(n4533) );
  XOR U11143 ( .A(n4907), .B(n4908), .Z(n4531) );
  AND U11144 ( .A(n4909), .B(n4910), .Z(n4907) );
  AND U11145 ( .A(b[29]), .B(a[85]), .Z(n4906) );
  XOR U11146 ( .A(n4911), .B(n4536), .Z(n4538) );
  XOR U11147 ( .A(n4912), .B(n4913), .Z(n4536) );
  AND U11148 ( .A(n4914), .B(n4915), .Z(n4912) );
  AND U11149 ( .A(b[28]), .B(a[86]), .Z(n4911) );
  XOR U11150 ( .A(n4916), .B(n4917), .Z(n4540) );
  AND U11151 ( .A(n4918), .B(n4919), .Z(n4916) );
  XOR U11152 ( .A(n4920), .B(n4545), .Z(n4547) );
  XOR U11153 ( .A(n4921), .B(n4922), .Z(n4545) );
  AND U11154 ( .A(n4923), .B(n4924), .Z(n4921) );
  AND U11155 ( .A(b[27]), .B(a[87]), .Z(n4920) );
  XOR U11156 ( .A(n4925), .B(n4550), .Z(n4552) );
  XOR U11157 ( .A(n4926), .B(n4927), .Z(n4550) );
  AND U11158 ( .A(n4928), .B(n4929), .Z(n4926) );
  AND U11159 ( .A(b[25]), .B(a[89]), .Z(n4925) );
  XOR U11160 ( .A(n4930), .B(n4555), .Z(n4557) );
  XOR U11161 ( .A(n4931), .B(n4932), .Z(n4555) );
  AND U11162 ( .A(n4933), .B(n4934), .Z(n4931) );
  AND U11163 ( .A(b[24]), .B(a[90]), .Z(n4930) );
  XOR U11164 ( .A(n4935), .B(n4560), .Z(n4562) );
  XOR U11165 ( .A(n4936), .B(n4937), .Z(n4560) );
  AND U11166 ( .A(n4938), .B(n4939), .Z(n4936) );
  AND U11167 ( .A(b[23]), .B(a[91]), .Z(n4935) );
  XOR U11168 ( .A(n4940), .B(n4565), .Z(n4567) );
  XOR U11169 ( .A(n4941), .B(n4942), .Z(n4565) );
  AND U11170 ( .A(n4943), .B(n4944), .Z(n4941) );
  AND U11171 ( .A(b[22]), .B(a[92]), .Z(n4940) );
  XOR U11172 ( .A(n4945), .B(n4946), .Z(n4569) );
  AND U11173 ( .A(n4947), .B(n4948), .Z(n4945) );
  XOR U11174 ( .A(n4949), .B(n4574), .Z(n4576) );
  XOR U11175 ( .A(n4950), .B(n4951), .Z(n4574) );
  AND U11176 ( .A(n4952), .B(n4953), .Z(n4950) );
  AND U11177 ( .A(b[21]), .B(a[93]), .Z(n4949) );
  XOR U11178 ( .A(n4954), .B(n4579), .Z(n4581) );
  XOR U11179 ( .A(n4955), .B(n4956), .Z(n4579) );
  AND U11180 ( .A(n4957), .B(n4958), .Z(n4955) );
  AND U11181 ( .A(b[19]), .B(a[95]), .Z(n4954) );
  XOR U11182 ( .A(n4959), .B(n4584), .Z(n4586) );
  XOR U11183 ( .A(n4960), .B(n4961), .Z(n4584) );
  AND U11184 ( .A(n4962), .B(n4963), .Z(n4960) );
  AND U11185 ( .A(b[18]), .B(a[96]), .Z(n4959) );
  XOR U11186 ( .A(n4964), .B(n4589), .Z(n4591) );
  XOR U11187 ( .A(n4965), .B(n4966), .Z(n4589) );
  AND U11188 ( .A(n4967), .B(n4968), .Z(n4965) );
  AND U11189 ( .A(b[17]), .B(a[97]), .Z(n4964) );
  XOR U11190 ( .A(n4969), .B(n4594), .Z(n4596) );
  XOR U11191 ( .A(n4970), .B(n4971), .Z(n4594) );
  AND U11192 ( .A(n4972), .B(n4973), .Z(n4970) );
  AND U11193 ( .A(b[16]), .B(a[98]), .Z(n4969) );
  XOR U11194 ( .A(n4974), .B(n4975), .Z(n4598) );
  AND U11195 ( .A(n4976), .B(n4977), .Z(n4974) );
  XOR U11196 ( .A(n4978), .B(n4603), .Z(n4605) );
  XOR U11197 ( .A(n4979), .B(n4980), .Z(n4603) );
  AND U11198 ( .A(n4981), .B(n4982), .Z(n4979) );
  AND U11199 ( .A(b[15]), .B(a[99]), .Z(n4978) );
  XOR U11200 ( .A(n4983), .B(n4608), .Z(n4610) );
  XOR U11201 ( .A(n4984), .B(n4985), .Z(n4608) );
  AND U11202 ( .A(n4986), .B(n4987), .Z(n4984) );
  AND U11203 ( .A(b[13]), .B(a[101]), .Z(n4983) );
  XOR U11204 ( .A(n4988), .B(n4613), .Z(n4615) );
  XOR U11205 ( .A(n4989), .B(n4990), .Z(n4613) );
  AND U11206 ( .A(n4991), .B(n4992), .Z(n4989) );
  AND U11207 ( .A(b[12]), .B(a[102]), .Z(n4988) );
  XOR U11208 ( .A(n4993), .B(n4618), .Z(n4620) );
  XOR U11209 ( .A(n4994), .B(n4995), .Z(n4618) );
  AND U11210 ( .A(n4996), .B(n4997), .Z(n4994) );
  AND U11211 ( .A(b[11]), .B(a[103]), .Z(n4993) );
  XOR U11212 ( .A(n4998), .B(n4623), .Z(n4625) );
  XOR U11213 ( .A(n4999), .B(n5000), .Z(n4623) );
  AND U11214 ( .A(n5001), .B(n5002), .Z(n4999) );
  AND U11215 ( .A(b[10]), .B(a[104]), .Z(n4998) );
  XOR U11216 ( .A(n5003), .B(n5004), .Z(n4627) );
  AND U11217 ( .A(n5005), .B(n5006), .Z(n5003) );
  XOR U11218 ( .A(n5007), .B(n4632), .Z(n4634) );
  XOR U11219 ( .A(n5008), .B(n5009), .Z(n4632) );
  AND U11220 ( .A(n5010), .B(n5011), .Z(n5008) );
  AND U11221 ( .A(b[9]), .B(a[105]), .Z(n5007) );
  XOR U11222 ( .A(n5012), .B(n4637), .Z(n4639) );
  XOR U11223 ( .A(n5013), .B(n5014), .Z(n4637) );
  AND U11224 ( .A(n5015), .B(n5016), .Z(n5013) );
  AND U11225 ( .A(b[7]), .B(a[107]), .Z(n5012) );
  XOR U11226 ( .A(n5017), .B(n4642), .Z(n4644) );
  XOR U11227 ( .A(n5018), .B(n5019), .Z(n4642) );
  AND U11228 ( .A(n5020), .B(n5021), .Z(n5018) );
  AND U11229 ( .A(b[6]), .B(a[108]), .Z(n5017) );
  XOR U11230 ( .A(n5022), .B(n4647), .Z(n4649) );
  XOR U11231 ( .A(n5023), .B(n5024), .Z(n4647) );
  AND U11232 ( .A(n5025), .B(n5026), .Z(n5023) );
  AND U11233 ( .A(b[5]), .B(a[109]), .Z(n5022) );
  XOR U11234 ( .A(n5027), .B(n4652), .Z(n4654) );
  XOR U11235 ( .A(n5028), .B(n5029), .Z(n4652) );
  AND U11236 ( .A(n5030), .B(n5031), .Z(n5028) );
  AND U11237 ( .A(b[4]), .B(a[110]), .Z(n5027) );
  XOR U11238 ( .A(n5032), .B(n5033), .Z(n4666) );
  NAND U11239 ( .A(n5034), .B(n5035), .Z(n5033) );
  XOR U11240 ( .A(n5036), .B(n4657), .Z(n4659) );
  XNOR U11241 ( .A(n5037), .B(n5038), .Z(n4657) );
  ANDN U11242 ( .B(n5039), .A(n5040), .Z(n5037) );
  AND U11243 ( .A(b[3]), .B(a[111]), .Z(n5036) );
  XNOR U11244 ( .A(n5041), .B(n5042), .Z(swire[113]) );
  XOR U11245 ( .A(n4676), .B(n5043), .Z(n5042) );
  NAND U11246 ( .A(a[113]), .B(b[0]), .Z(n4675) );
  XOR U11247 ( .A(n5044), .B(n5045), .Z(n5034) );
  NAND U11248 ( .A(b[1]), .B(a[112]), .Z(n5045) );
  XNOR U11249 ( .A(n5044), .B(n5040), .Z(n5046) );
  XOR U11250 ( .A(n5047), .B(n5038), .Z(n5040) );
  AND U11251 ( .A(b[2]), .B(a[111]), .Z(n5047) );
  IV U11252 ( .A(n5032), .Z(n5044) );
  ANDN U11253 ( .B(n5048), .A(n5049), .Z(n5032) );
  XOR U11254 ( .A(n5038), .B(n5030), .Z(n5050) );
  XNOR U11255 ( .A(n5029), .B(n5025), .Z(n5051) );
  XNOR U11256 ( .A(n5024), .B(n5020), .Z(n5052) );
  XNOR U11257 ( .A(n5019), .B(n5015), .Z(n5053) );
  XNOR U11258 ( .A(n5006), .B(n5005), .Z(n5054) );
  XOR U11259 ( .A(n5055), .B(n5004), .Z(n5005) );
  AND U11260 ( .A(b[7]), .B(a[106]), .Z(n5055) );
  XNOR U11261 ( .A(n5004), .B(n5010), .Z(n5056) );
  XNOR U11262 ( .A(n5009), .B(n5001), .Z(n5057) );
  XNOR U11263 ( .A(n5000), .B(n4996), .Z(n5058) );
  XNOR U11264 ( .A(n4995), .B(n4991), .Z(n5059) );
  XNOR U11265 ( .A(n4990), .B(n4986), .Z(n5060) );
  XNOR U11266 ( .A(n4977), .B(n4976), .Z(n5061) );
  XOR U11267 ( .A(n5062), .B(n4975), .Z(n4976) );
  AND U11268 ( .A(b[13]), .B(a[100]), .Z(n5062) );
  XNOR U11269 ( .A(n4975), .B(n4981), .Z(n5063) );
  XNOR U11270 ( .A(n4980), .B(n4972), .Z(n5064) );
  XNOR U11271 ( .A(n4971), .B(n4967), .Z(n5065) );
  XNOR U11272 ( .A(n4966), .B(n4962), .Z(n5066) );
  XNOR U11273 ( .A(n4961), .B(n4957), .Z(n5067) );
  XNOR U11274 ( .A(n4948), .B(n4947), .Z(n5068) );
  XOR U11275 ( .A(n5069), .B(n4946), .Z(n4947) );
  AND U11276 ( .A(b[19]), .B(a[94]), .Z(n5069) );
  XNOR U11277 ( .A(n4946), .B(n4952), .Z(n5070) );
  XNOR U11278 ( .A(n4951), .B(n4943), .Z(n5071) );
  XNOR U11279 ( .A(n4942), .B(n4938), .Z(n5072) );
  XNOR U11280 ( .A(n4937), .B(n4933), .Z(n5073) );
  XNOR U11281 ( .A(n4932), .B(n4928), .Z(n5074) );
  XNOR U11282 ( .A(n4919), .B(n4918), .Z(n5075) );
  XOR U11283 ( .A(n5076), .B(n4917), .Z(n4918) );
  AND U11284 ( .A(b[25]), .B(a[88]), .Z(n5076) );
  XNOR U11285 ( .A(n4917), .B(n4923), .Z(n5077) );
  XNOR U11286 ( .A(n4922), .B(n4914), .Z(n5078) );
  XNOR U11287 ( .A(n4913), .B(n4909), .Z(n5079) );
  XNOR U11288 ( .A(n4908), .B(n4904), .Z(n5080) );
  XNOR U11289 ( .A(n4903), .B(n4899), .Z(n5081) );
  XNOR U11290 ( .A(n4890), .B(n4889), .Z(n5082) );
  XOR U11291 ( .A(n5083), .B(n4888), .Z(n4889) );
  AND U11292 ( .A(b[31]), .B(a[82]), .Z(n5083) );
  XNOR U11293 ( .A(n4888), .B(n4894), .Z(n5084) );
  XNOR U11294 ( .A(n4893), .B(n4885), .Z(n5085) );
  XNOR U11295 ( .A(n4884), .B(n4880), .Z(n5086) );
  XNOR U11296 ( .A(n4879), .B(n4875), .Z(n5087) );
  XNOR U11297 ( .A(n4874), .B(n4870), .Z(n5088) );
  XNOR U11298 ( .A(n4861), .B(n4860), .Z(n5089) );
  XOR U11299 ( .A(n5090), .B(n4859), .Z(n4860) );
  AND U11300 ( .A(b[37]), .B(a[76]), .Z(n5090) );
  XNOR U11301 ( .A(n4859), .B(n4865), .Z(n5091) );
  XNOR U11302 ( .A(n4864), .B(n4856), .Z(n5092) );
  XNOR U11303 ( .A(n4855), .B(n4851), .Z(n5093) );
  XNOR U11304 ( .A(n4850), .B(n4846), .Z(n5094) );
  XNOR U11305 ( .A(n4845), .B(n4841), .Z(n5095) );
  XNOR U11306 ( .A(n4832), .B(n4831), .Z(n5096) );
  XOR U11307 ( .A(n5097), .B(n4830), .Z(n4831) );
  AND U11308 ( .A(b[43]), .B(a[70]), .Z(n5097) );
  XNOR U11309 ( .A(n4830), .B(n4836), .Z(n5098) );
  XNOR U11310 ( .A(n4835), .B(n4827), .Z(n5099) );
  XNOR U11311 ( .A(n4826), .B(n4822), .Z(n5100) );
  XNOR U11312 ( .A(n4821), .B(n4817), .Z(n5101) );
  XNOR U11313 ( .A(n4816), .B(n4812), .Z(n5102) );
  XNOR U11314 ( .A(n4811), .B(n4807), .Z(n5103) );
  XNOR U11315 ( .A(n4806), .B(n4802), .Z(n5104) );
  XNOR U11316 ( .A(n4801), .B(n4797), .Z(n5105) );
  XNOR U11317 ( .A(n4796), .B(n4792), .Z(n5106) );
  XNOR U11318 ( .A(n4791), .B(n4787), .Z(n5107) );
  XNOR U11319 ( .A(n4786), .B(n4782), .Z(n5108) );
  XNOR U11320 ( .A(n4781), .B(n4777), .Z(n5109) );
  XNOR U11321 ( .A(n4776), .B(n4772), .Z(n5110) );
  XNOR U11322 ( .A(n4771), .B(n4767), .Z(n5111) );
  XNOR U11323 ( .A(n4766), .B(n4762), .Z(n5112) );
  XNOR U11324 ( .A(n4761), .B(n4757), .Z(n5113) );
  XOR U11325 ( .A(n4756), .B(n4753), .Z(n5114) );
  XOR U11326 ( .A(n5115), .B(n5116), .Z(n4753) );
  XOR U11327 ( .A(n4751), .B(n5117), .Z(n5116) );
  XOR U11328 ( .A(n5118), .B(n5119), .Z(n5117) );
  XOR U11329 ( .A(n5120), .B(n5121), .Z(n5119) );
  NAND U11330 ( .A(a[51]), .B(b[62]), .Z(n5121) );
  AND U11331 ( .A(a[50]), .B(b[63]), .Z(n5120) );
  XOR U11332 ( .A(n5122), .B(n5118), .Z(n5115) );
  XOR U11333 ( .A(n5123), .B(n5124), .Z(n5118) );
  ANDN U11334 ( .B(n5125), .A(n5126), .Z(n5123) );
  AND U11335 ( .A(a[52]), .B(b[61]), .Z(n5122) );
  XOR U11336 ( .A(n5127), .B(n4751), .Z(n4752) );
  XOR U11337 ( .A(n5128), .B(n5129), .Z(n4751) );
  AND U11338 ( .A(n5130), .B(n5131), .Z(n5128) );
  AND U11339 ( .A(a[53]), .B(b[60]), .Z(n5127) );
  XOR U11340 ( .A(n5132), .B(n4756), .Z(n4758) );
  XOR U11341 ( .A(n5133), .B(n5134), .Z(n4756) );
  AND U11342 ( .A(n5135), .B(n5136), .Z(n5133) );
  AND U11343 ( .A(a[54]), .B(b[59]), .Z(n5132) );
  XOR U11344 ( .A(n5137), .B(n4761), .Z(n4763) );
  XOR U11345 ( .A(n5138), .B(n5139), .Z(n4761) );
  AND U11346 ( .A(n5140), .B(n5141), .Z(n5138) );
  AND U11347 ( .A(a[55]), .B(b[58]), .Z(n5137) );
  XOR U11348 ( .A(n5142), .B(n4766), .Z(n4768) );
  XOR U11349 ( .A(n5143), .B(n5144), .Z(n4766) );
  AND U11350 ( .A(n5145), .B(n5146), .Z(n5143) );
  AND U11351 ( .A(a[56]), .B(b[57]), .Z(n5142) );
  XOR U11352 ( .A(n5147), .B(n4771), .Z(n4773) );
  XOR U11353 ( .A(n5148), .B(n5149), .Z(n4771) );
  AND U11354 ( .A(n5150), .B(n5151), .Z(n5148) );
  AND U11355 ( .A(b[56]), .B(a[57]), .Z(n5147) );
  XOR U11356 ( .A(n5152), .B(n4776), .Z(n4778) );
  XOR U11357 ( .A(n5153), .B(n5154), .Z(n4776) );
  AND U11358 ( .A(n5155), .B(n5156), .Z(n5153) );
  AND U11359 ( .A(b[55]), .B(a[58]), .Z(n5152) );
  XOR U11360 ( .A(n5157), .B(n4781), .Z(n4783) );
  XOR U11361 ( .A(n5158), .B(n5159), .Z(n4781) );
  AND U11362 ( .A(n5160), .B(n5161), .Z(n5158) );
  AND U11363 ( .A(b[54]), .B(a[59]), .Z(n5157) );
  XOR U11364 ( .A(n5162), .B(n4786), .Z(n4788) );
  XOR U11365 ( .A(n5163), .B(n5164), .Z(n4786) );
  AND U11366 ( .A(n5165), .B(n5166), .Z(n5163) );
  AND U11367 ( .A(b[53]), .B(a[60]), .Z(n5162) );
  XOR U11368 ( .A(n5167), .B(n4791), .Z(n4793) );
  XOR U11369 ( .A(n5168), .B(n5169), .Z(n4791) );
  AND U11370 ( .A(n5170), .B(n5171), .Z(n5168) );
  AND U11371 ( .A(b[52]), .B(a[61]), .Z(n5167) );
  XOR U11372 ( .A(n5172), .B(n4796), .Z(n4798) );
  XOR U11373 ( .A(n5173), .B(n5174), .Z(n4796) );
  AND U11374 ( .A(n5175), .B(n5176), .Z(n5173) );
  AND U11375 ( .A(b[51]), .B(a[62]), .Z(n5172) );
  XOR U11376 ( .A(n5177), .B(n4801), .Z(n4803) );
  XOR U11377 ( .A(n5178), .B(n5179), .Z(n4801) );
  AND U11378 ( .A(n5180), .B(n5181), .Z(n5178) );
  AND U11379 ( .A(b[50]), .B(a[63]), .Z(n5177) );
  XOR U11380 ( .A(n5182), .B(n4806), .Z(n4808) );
  XOR U11381 ( .A(n5183), .B(n5184), .Z(n4806) );
  AND U11382 ( .A(n5185), .B(n5186), .Z(n5183) );
  AND U11383 ( .A(b[49]), .B(a[64]), .Z(n5182) );
  XOR U11384 ( .A(n5187), .B(n4811), .Z(n4813) );
  XOR U11385 ( .A(n5188), .B(n5189), .Z(n4811) );
  AND U11386 ( .A(n5190), .B(n5191), .Z(n5188) );
  AND U11387 ( .A(b[48]), .B(a[65]), .Z(n5187) );
  XOR U11388 ( .A(n5192), .B(n4816), .Z(n4818) );
  XOR U11389 ( .A(n5193), .B(n5194), .Z(n4816) );
  AND U11390 ( .A(n5195), .B(n5196), .Z(n5193) );
  AND U11391 ( .A(b[47]), .B(a[66]), .Z(n5192) );
  XOR U11392 ( .A(n5197), .B(n4821), .Z(n4823) );
  XOR U11393 ( .A(n5198), .B(n5199), .Z(n4821) );
  AND U11394 ( .A(n5200), .B(n5201), .Z(n5198) );
  AND U11395 ( .A(b[46]), .B(a[67]), .Z(n5197) );
  XOR U11396 ( .A(n5202), .B(n4826), .Z(n4828) );
  XOR U11397 ( .A(n5203), .B(n5204), .Z(n4826) );
  AND U11398 ( .A(n5205), .B(n5206), .Z(n5203) );
  AND U11399 ( .A(b[45]), .B(a[68]), .Z(n5202) );
  XOR U11400 ( .A(n5207), .B(n5208), .Z(n4830) );
  AND U11401 ( .A(n5209), .B(n5210), .Z(n5207) );
  XOR U11402 ( .A(n5211), .B(n4835), .Z(n4837) );
  XOR U11403 ( .A(n5212), .B(n5213), .Z(n4835) );
  AND U11404 ( .A(n5214), .B(n5215), .Z(n5212) );
  AND U11405 ( .A(b[44]), .B(a[69]), .Z(n5211) );
  XOR U11406 ( .A(n5216), .B(n4840), .Z(n4842) );
  XOR U11407 ( .A(n5217), .B(n5218), .Z(n4840) );
  AND U11408 ( .A(n5219), .B(n5220), .Z(n5217) );
  AND U11409 ( .A(b[42]), .B(a[71]), .Z(n5216) );
  XOR U11410 ( .A(n5221), .B(n4845), .Z(n4847) );
  XOR U11411 ( .A(n5222), .B(n5223), .Z(n4845) );
  AND U11412 ( .A(n5224), .B(n5225), .Z(n5222) );
  AND U11413 ( .A(b[41]), .B(a[72]), .Z(n5221) );
  XOR U11414 ( .A(n5226), .B(n4850), .Z(n4852) );
  XOR U11415 ( .A(n5227), .B(n5228), .Z(n4850) );
  AND U11416 ( .A(n5229), .B(n5230), .Z(n5227) );
  AND U11417 ( .A(b[40]), .B(a[73]), .Z(n5226) );
  XOR U11418 ( .A(n5231), .B(n4855), .Z(n4857) );
  XOR U11419 ( .A(n5232), .B(n5233), .Z(n4855) );
  AND U11420 ( .A(n5234), .B(n5235), .Z(n5232) );
  AND U11421 ( .A(b[39]), .B(a[74]), .Z(n5231) );
  XOR U11422 ( .A(n5236), .B(n5237), .Z(n4859) );
  AND U11423 ( .A(n5238), .B(n5239), .Z(n5236) );
  XOR U11424 ( .A(n5240), .B(n4864), .Z(n4866) );
  XOR U11425 ( .A(n5241), .B(n5242), .Z(n4864) );
  AND U11426 ( .A(n5243), .B(n5244), .Z(n5241) );
  AND U11427 ( .A(b[38]), .B(a[75]), .Z(n5240) );
  XOR U11428 ( .A(n5245), .B(n4869), .Z(n4871) );
  XOR U11429 ( .A(n5246), .B(n5247), .Z(n4869) );
  AND U11430 ( .A(n5248), .B(n5249), .Z(n5246) );
  AND U11431 ( .A(b[36]), .B(a[77]), .Z(n5245) );
  XOR U11432 ( .A(n5250), .B(n4874), .Z(n4876) );
  XOR U11433 ( .A(n5251), .B(n5252), .Z(n4874) );
  AND U11434 ( .A(n5253), .B(n5254), .Z(n5251) );
  AND U11435 ( .A(b[35]), .B(a[78]), .Z(n5250) );
  XOR U11436 ( .A(n5255), .B(n4879), .Z(n4881) );
  XOR U11437 ( .A(n5256), .B(n5257), .Z(n4879) );
  AND U11438 ( .A(n5258), .B(n5259), .Z(n5256) );
  AND U11439 ( .A(b[34]), .B(a[79]), .Z(n5255) );
  XOR U11440 ( .A(n5260), .B(n4884), .Z(n4886) );
  XOR U11441 ( .A(n5261), .B(n5262), .Z(n4884) );
  AND U11442 ( .A(n5263), .B(n5264), .Z(n5261) );
  AND U11443 ( .A(b[33]), .B(a[80]), .Z(n5260) );
  XOR U11444 ( .A(n5265), .B(n5266), .Z(n4888) );
  AND U11445 ( .A(n5267), .B(n5268), .Z(n5265) );
  XOR U11446 ( .A(n5269), .B(n4893), .Z(n4895) );
  XOR U11447 ( .A(n5270), .B(n5271), .Z(n4893) );
  AND U11448 ( .A(n5272), .B(n5273), .Z(n5270) );
  AND U11449 ( .A(b[32]), .B(a[81]), .Z(n5269) );
  XOR U11450 ( .A(n5274), .B(n4898), .Z(n4900) );
  XOR U11451 ( .A(n5275), .B(n5276), .Z(n4898) );
  AND U11452 ( .A(n5277), .B(n5278), .Z(n5275) );
  AND U11453 ( .A(b[30]), .B(a[83]), .Z(n5274) );
  XOR U11454 ( .A(n5279), .B(n4903), .Z(n4905) );
  XOR U11455 ( .A(n5280), .B(n5281), .Z(n4903) );
  AND U11456 ( .A(n5282), .B(n5283), .Z(n5280) );
  AND U11457 ( .A(b[29]), .B(a[84]), .Z(n5279) );
  XOR U11458 ( .A(n5284), .B(n4908), .Z(n4910) );
  XOR U11459 ( .A(n5285), .B(n5286), .Z(n4908) );
  AND U11460 ( .A(n5287), .B(n5288), .Z(n5285) );
  AND U11461 ( .A(b[28]), .B(a[85]), .Z(n5284) );
  XOR U11462 ( .A(n5289), .B(n4913), .Z(n4915) );
  XOR U11463 ( .A(n5290), .B(n5291), .Z(n4913) );
  AND U11464 ( .A(n5292), .B(n5293), .Z(n5290) );
  AND U11465 ( .A(b[27]), .B(a[86]), .Z(n5289) );
  XOR U11466 ( .A(n5294), .B(n5295), .Z(n4917) );
  AND U11467 ( .A(n5296), .B(n5297), .Z(n5294) );
  XOR U11468 ( .A(n5298), .B(n4922), .Z(n4924) );
  XOR U11469 ( .A(n5299), .B(n5300), .Z(n4922) );
  AND U11470 ( .A(n5301), .B(n5302), .Z(n5299) );
  AND U11471 ( .A(b[26]), .B(a[87]), .Z(n5298) );
  XOR U11472 ( .A(n5303), .B(n4927), .Z(n4929) );
  XOR U11473 ( .A(n5304), .B(n5305), .Z(n4927) );
  AND U11474 ( .A(n5306), .B(n5307), .Z(n5304) );
  AND U11475 ( .A(b[24]), .B(a[89]), .Z(n5303) );
  XOR U11476 ( .A(n5308), .B(n4932), .Z(n4934) );
  XOR U11477 ( .A(n5309), .B(n5310), .Z(n4932) );
  AND U11478 ( .A(n5311), .B(n5312), .Z(n5309) );
  AND U11479 ( .A(b[23]), .B(a[90]), .Z(n5308) );
  XOR U11480 ( .A(n5313), .B(n4937), .Z(n4939) );
  XOR U11481 ( .A(n5314), .B(n5315), .Z(n4937) );
  AND U11482 ( .A(n5316), .B(n5317), .Z(n5314) );
  AND U11483 ( .A(b[22]), .B(a[91]), .Z(n5313) );
  XOR U11484 ( .A(n5318), .B(n4942), .Z(n4944) );
  XOR U11485 ( .A(n5319), .B(n5320), .Z(n4942) );
  AND U11486 ( .A(n5321), .B(n5322), .Z(n5319) );
  AND U11487 ( .A(b[21]), .B(a[92]), .Z(n5318) );
  XOR U11488 ( .A(n5323), .B(n5324), .Z(n4946) );
  AND U11489 ( .A(n5325), .B(n5326), .Z(n5323) );
  XOR U11490 ( .A(n5327), .B(n4951), .Z(n4953) );
  XOR U11491 ( .A(n5328), .B(n5329), .Z(n4951) );
  AND U11492 ( .A(n5330), .B(n5331), .Z(n5328) );
  AND U11493 ( .A(b[20]), .B(a[93]), .Z(n5327) );
  XOR U11494 ( .A(n5332), .B(n4956), .Z(n4958) );
  XOR U11495 ( .A(n5333), .B(n5334), .Z(n4956) );
  AND U11496 ( .A(n5335), .B(n5336), .Z(n5333) );
  AND U11497 ( .A(b[18]), .B(a[95]), .Z(n5332) );
  XOR U11498 ( .A(n5337), .B(n4961), .Z(n4963) );
  XOR U11499 ( .A(n5338), .B(n5339), .Z(n4961) );
  AND U11500 ( .A(n5340), .B(n5341), .Z(n5338) );
  AND U11501 ( .A(b[17]), .B(a[96]), .Z(n5337) );
  XOR U11502 ( .A(n5342), .B(n4966), .Z(n4968) );
  XOR U11503 ( .A(n5343), .B(n5344), .Z(n4966) );
  AND U11504 ( .A(n5345), .B(n5346), .Z(n5343) );
  AND U11505 ( .A(b[16]), .B(a[97]), .Z(n5342) );
  XOR U11506 ( .A(n5347), .B(n4971), .Z(n4973) );
  XOR U11507 ( .A(n5348), .B(n5349), .Z(n4971) );
  AND U11508 ( .A(n5350), .B(n5351), .Z(n5348) );
  AND U11509 ( .A(b[15]), .B(a[98]), .Z(n5347) );
  XOR U11510 ( .A(n5352), .B(n5353), .Z(n4975) );
  AND U11511 ( .A(n5354), .B(n5355), .Z(n5352) );
  XOR U11512 ( .A(n5356), .B(n4980), .Z(n4982) );
  XOR U11513 ( .A(n5357), .B(n5358), .Z(n4980) );
  AND U11514 ( .A(n5359), .B(n5360), .Z(n5357) );
  AND U11515 ( .A(b[14]), .B(a[99]), .Z(n5356) );
  XOR U11516 ( .A(n5361), .B(n4985), .Z(n4987) );
  XOR U11517 ( .A(n5362), .B(n5363), .Z(n4985) );
  AND U11518 ( .A(n5364), .B(n5365), .Z(n5362) );
  AND U11519 ( .A(b[12]), .B(a[101]), .Z(n5361) );
  XOR U11520 ( .A(n5366), .B(n4990), .Z(n4992) );
  XOR U11521 ( .A(n5367), .B(n5368), .Z(n4990) );
  AND U11522 ( .A(n5369), .B(n5370), .Z(n5367) );
  AND U11523 ( .A(b[11]), .B(a[102]), .Z(n5366) );
  XOR U11524 ( .A(n5371), .B(n4995), .Z(n4997) );
  XOR U11525 ( .A(n5372), .B(n5373), .Z(n4995) );
  AND U11526 ( .A(n5374), .B(n5375), .Z(n5372) );
  AND U11527 ( .A(b[10]), .B(a[103]), .Z(n5371) );
  XOR U11528 ( .A(n5376), .B(n5000), .Z(n5002) );
  XOR U11529 ( .A(n5377), .B(n5378), .Z(n5000) );
  AND U11530 ( .A(n5379), .B(n5380), .Z(n5377) );
  AND U11531 ( .A(b[9]), .B(a[104]), .Z(n5376) );
  XOR U11532 ( .A(n5381), .B(n5382), .Z(n5004) );
  AND U11533 ( .A(n5383), .B(n5384), .Z(n5381) );
  XOR U11534 ( .A(n5385), .B(n5009), .Z(n5011) );
  XOR U11535 ( .A(n5386), .B(n5387), .Z(n5009) );
  AND U11536 ( .A(n5388), .B(n5389), .Z(n5386) );
  AND U11537 ( .A(b[8]), .B(a[105]), .Z(n5385) );
  XOR U11538 ( .A(n5390), .B(n5014), .Z(n5016) );
  XOR U11539 ( .A(n5391), .B(n5392), .Z(n5014) );
  AND U11540 ( .A(n5393), .B(n5394), .Z(n5391) );
  AND U11541 ( .A(b[6]), .B(a[107]), .Z(n5390) );
  XOR U11542 ( .A(n5395), .B(n5019), .Z(n5021) );
  XOR U11543 ( .A(n5396), .B(n5397), .Z(n5019) );
  AND U11544 ( .A(n5398), .B(n5399), .Z(n5396) );
  AND U11545 ( .A(b[5]), .B(a[108]), .Z(n5395) );
  XOR U11546 ( .A(n5400), .B(n5024), .Z(n5026) );
  XOR U11547 ( .A(n5401), .B(n5402), .Z(n5024) );
  AND U11548 ( .A(n5403), .B(n5404), .Z(n5401) );
  AND U11549 ( .A(b[4]), .B(a[109]), .Z(n5400) );
  XOR U11550 ( .A(n5405), .B(n5406), .Z(n5038) );
  NANDN U11551 ( .A(n5407), .B(n5408), .Z(n5406) );
  XOR U11552 ( .A(n5409), .B(n5029), .Z(n5031) );
  XNOR U11553 ( .A(n5410), .B(n5411), .Z(n5029) );
  AND U11554 ( .A(n5412), .B(n5413), .Z(n5410) );
  AND U11555 ( .A(b[3]), .B(a[110]), .Z(n5409) );
  XNOR U11556 ( .A(n5414), .B(n5415), .Z(swire[112]) );
  XOR U11557 ( .A(n5048), .B(n5416), .Z(n5415) );
  NAND U11558 ( .A(a[112]), .B(b[0]), .Z(n5049) );
  XNOR U11559 ( .A(n5408), .B(n5407), .Z(n5048) );
  XOR U11560 ( .A(n5405), .B(n5417), .Z(n5407) );
  NAND U11561 ( .A(b[1]), .B(a[111]), .Z(n5417) );
  XNOR U11562 ( .A(n5413), .B(n5418), .Z(n5408) );
  XNOR U11563 ( .A(n5405), .B(n5412), .Z(n5418) );
  XNOR U11564 ( .A(n5419), .B(n5411), .Z(n5412) );
  AND U11565 ( .A(b[2]), .B(a[110]), .Z(n5419) );
  ANDN U11566 ( .B(n5420), .A(n5421), .Z(n5405) );
  XOR U11567 ( .A(n5411), .B(n5403), .Z(n5422) );
  XNOR U11568 ( .A(n5402), .B(n5398), .Z(n5423) );
  XNOR U11569 ( .A(n5397), .B(n5393), .Z(n5424) );
  XNOR U11570 ( .A(n5384), .B(n5383), .Z(n5425) );
  XOR U11571 ( .A(n5426), .B(n5382), .Z(n5383) );
  AND U11572 ( .A(b[6]), .B(a[106]), .Z(n5426) );
  XNOR U11573 ( .A(n5382), .B(n5388), .Z(n5427) );
  XNOR U11574 ( .A(n5387), .B(n5379), .Z(n5428) );
  XNOR U11575 ( .A(n5378), .B(n5374), .Z(n5429) );
  XNOR U11576 ( .A(n5373), .B(n5369), .Z(n5430) );
  XNOR U11577 ( .A(n5368), .B(n5364), .Z(n5431) );
  XNOR U11578 ( .A(n5355), .B(n5354), .Z(n5432) );
  XOR U11579 ( .A(n5433), .B(n5353), .Z(n5354) );
  AND U11580 ( .A(b[12]), .B(a[100]), .Z(n5433) );
  XNOR U11581 ( .A(n5353), .B(n5359), .Z(n5434) );
  XNOR U11582 ( .A(n5358), .B(n5350), .Z(n5435) );
  XNOR U11583 ( .A(n5349), .B(n5345), .Z(n5436) );
  XNOR U11584 ( .A(n5344), .B(n5340), .Z(n5437) );
  XNOR U11585 ( .A(n5339), .B(n5335), .Z(n5438) );
  XNOR U11586 ( .A(n5326), .B(n5325), .Z(n5439) );
  XOR U11587 ( .A(n5440), .B(n5324), .Z(n5325) );
  AND U11588 ( .A(b[18]), .B(a[94]), .Z(n5440) );
  XNOR U11589 ( .A(n5324), .B(n5330), .Z(n5441) );
  XNOR U11590 ( .A(n5329), .B(n5321), .Z(n5442) );
  XNOR U11591 ( .A(n5320), .B(n5316), .Z(n5443) );
  XNOR U11592 ( .A(n5315), .B(n5311), .Z(n5444) );
  XNOR U11593 ( .A(n5310), .B(n5306), .Z(n5445) );
  XNOR U11594 ( .A(n5297), .B(n5296), .Z(n5446) );
  XOR U11595 ( .A(n5447), .B(n5295), .Z(n5296) );
  AND U11596 ( .A(b[24]), .B(a[88]), .Z(n5447) );
  XNOR U11597 ( .A(n5295), .B(n5301), .Z(n5448) );
  XNOR U11598 ( .A(n5300), .B(n5292), .Z(n5449) );
  XNOR U11599 ( .A(n5291), .B(n5287), .Z(n5450) );
  XNOR U11600 ( .A(n5286), .B(n5282), .Z(n5451) );
  XNOR U11601 ( .A(n5281), .B(n5277), .Z(n5452) );
  XNOR U11602 ( .A(n5268), .B(n5267), .Z(n5453) );
  XOR U11603 ( .A(n5454), .B(n5266), .Z(n5267) );
  AND U11604 ( .A(b[30]), .B(a[82]), .Z(n5454) );
  XNOR U11605 ( .A(n5266), .B(n5272), .Z(n5455) );
  XNOR U11606 ( .A(n5271), .B(n5263), .Z(n5456) );
  XNOR U11607 ( .A(n5262), .B(n5258), .Z(n5457) );
  XNOR U11608 ( .A(n5257), .B(n5253), .Z(n5458) );
  XNOR U11609 ( .A(n5252), .B(n5248), .Z(n5459) );
  XNOR U11610 ( .A(n5239), .B(n5238), .Z(n5460) );
  XOR U11611 ( .A(n5461), .B(n5237), .Z(n5238) );
  AND U11612 ( .A(b[36]), .B(a[76]), .Z(n5461) );
  XNOR U11613 ( .A(n5237), .B(n5243), .Z(n5462) );
  XNOR U11614 ( .A(n5242), .B(n5234), .Z(n5463) );
  XNOR U11615 ( .A(n5233), .B(n5229), .Z(n5464) );
  XNOR U11616 ( .A(n5228), .B(n5224), .Z(n5465) );
  XNOR U11617 ( .A(n5223), .B(n5219), .Z(n5466) );
  XNOR U11618 ( .A(n5210), .B(n5209), .Z(n5467) );
  XOR U11619 ( .A(n5468), .B(n5208), .Z(n5209) );
  AND U11620 ( .A(b[42]), .B(a[70]), .Z(n5468) );
  XNOR U11621 ( .A(n5208), .B(n5214), .Z(n5469) );
  XNOR U11622 ( .A(n5213), .B(n5205), .Z(n5470) );
  XNOR U11623 ( .A(n5204), .B(n5200), .Z(n5471) );
  XNOR U11624 ( .A(n5199), .B(n5195), .Z(n5472) );
  XNOR U11625 ( .A(n5194), .B(n5190), .Z(n5473) );
  XNOR U11626 ( .A(n5189), .B(n5185), .Z(n5474) );
  XNOR U11627 ( .A(n5184), .B(n5180), .Z(n5475) );
  XNOR U11628 ( .A(n5179), .B(n5175), .Z(n5476) );
  XNOR U11629 ( .A(n5174), .B(n5170), .Z(n5477) );
  XNOR U11630 ( .A(n5169), .B(n5165), .Z(n5478) );
  XNOR U11631 ( .A(n5164), .B(n5160), .Z(n5479) );
  XNOR U11632 ( .A(n5159), .B(n5155), .Z(n5480) );
  XNOR U11633 ( .A(n5154), .B(n5150), .Z(n5481) );
  XNOR U11634 ( .A(n5149), .B(n5145), .Z(n5482) );
  XNOR U11635 ( .A(n5144), .B(n5140), .Z(n5483) );
  XNOR U11636 ( .A(n5139), .B(n5135), .Z(n5484) );
  XNOR U11637 ( .A(n5134), .B(n5130), .Z(n5485) );
  XOR U11638 ( .A(n5129), .B(n5126), .Z(n5486) );
  XOR U11639 ( .A(n5487), .B(n5488), .Z(n5126) );
  XOR U11640 ( .A(n5124), .B(n5489), .Z(n5488) );
  XOR U11641 ( .A(n5490), .B(n5491), .Z(n5489) );
  XOR U11642 ( .A(n5492), .B(n5493), .Z(n5491) );
  NAND U11643 ( .A(a[50]), .B(b[62]), .Z(n5493) );
  AND U11644 ( .A(a[49]), .B(b[63]), .Z(n5492) );
  XOR U11645 ( .A(n5494), .B(n5490), .Z(n5487) );
  XOR U11646 ( .A(n5495), .B(n5496), .Z(n5490) );
  ANDN U11647 ( .B(n5497), .A(n5498), .Z(n5495) );
  AND U11648 ( .A(a[51]), .B(b[61]), .Z(n5494) );
  XOR U11649 ( .A(n5499), .B(n5124), .Z(n5125) );
  XOR U11650 ( .A(n5500), .B(n5501), .Z(n5124) );
  AND U11651 ( .A(n5502), .B(n5503), .Z(n5500) );
  AND U11652 ( .A(a[52]), .B(b[60]), .Z(n5499) );
  XOR U11653 ( .A(n5504), .B(n5129), .Z(n5131) );
  XOR U11654 ( .A(n5505), .B(n5506), .Z(n5129) );
  AND U11655 ( .A(n5507), .B(n5508), .Z(n5505) );
  AND U11656 ( .A(a[53]), .B(b[59]), .Z(n5504) );
  XOR U11657 ( .A(n5509), .B(n5134), .Z(n5136) );
  XOR U11658 ( .A(n5510), .B(n5511), .Z(n5134) );
  AND U11659 ( .A(n5512), .B(n5513), .Z(n5510) );
  AND U11660 ( .A(a[54]), .B(b[58]), .Z(n5509) );
  XOR U11661 ( .A(n5514), .B(n5139), .Z(n5141) );
  XOR U11662 ( .A(n5515), .B(n5516), .Z(n5139) );
  AND U11663 ( .A(n5517), .B(n5518), .Z(n5515) );
  AND U11664 ( .A(a[55]), .B(b[57]), .Z(n5514) );
  XOR U11665 ( .A(n5519), .B(n5144), .Z(n5146) );
  XOR U11666 ( .A(n5520), .B(n5521), .Z(n5144) );
  AND U11667 ( .A(n5522), .B(n5523), .Z(n5520) );
  AND U11668 ( .A(a[56]), .B(b[56]), .Z(n5519) );
  XOR U11669 ( .A(n5524), .B(n5149), .Z(n5151) );
  XOR U11670 ( .A(n5525), .B(n5526), .Z(n5149) );
  AND U11671 ( .A(n5527), .B(n5528), .Z(n5525) );
  AND U11672 ( .A(b[55]), .B(a[57]), .Z(n5524) );
  XOR U11673 ( .A(n5529), .B(n5154), .Z(n5156) );
  XOR U11674 ( .A(n5530), .B(n5531), .Z(n5154) );
  AND U11675 ( .A(n5532), .B(n5533), .Z(n5530) );
  AND U11676 ( .A(b[54]), .B(a[58]), .Z(n5529) );
  XOR U11677 ( .A(n5534), .B(n5159), .Z(n5161) );
  XOR U11678 ( .A(n5535), .B(n5536), .Z(n5159) );
  AND U11679 ( .A(n5537), .B(n5538), .Z(n5535) );
  AND U11680 ( .A(b[53]), .B(a[59]), .Z(n5534) );
  XOR U11681 ( .A(n5539), .B(n5164), .Z(n5166) );
  XOR U11682 ( .A(n5540), .B(n5541), .Z(n5164) );
  AND U11683 ( .A(n5542), .B(n5543), .Z(n5540) );
  AND U11684 ( .A(b[52]), .B(a[60]), .Z(n5539) );
  XOR U11685 ( .A(n5544), .B(n5169), .Z(n5171) );
  XOR U11686 ( .A(n5545), .B(n5546), .Z(n5169) );
  AND U11687 ( .A(n5547), .B(n5548), .Z(n5545) );
  AND U11688 ( .A(b[51]), .B(a[61]), .Z(n5544) );
  XOR U11689 ( .A(n5549), .B(n5174), .Z(n5176) );
  XOR U11690 ( .A(n5550), .B(n5551), .Z(n5174) );
  AND U11691 ( .A(n5552), .B(n5553), .Z(n5550) );
  AND U11692 ( .A(b[50]), .B(a[62]), .Z(n5549) );
  XOR U11693 ( .A(n5554), .B(n5179), .Z(n5181) );
  XOR U11694 ( .A(n5555), .B(n5556), .Z(n5179) );
  AND U11695 ( .A(n5557), .B(n5558), .Z(n5555) );
  AND U11696 ( .A(b[49]), .B(a[63]), .Z(n5554) );
  XOR U11697 ( .A(n5559), .B(n5184), .Z(n5186) );
  XOR U11698 ( .A(n5560), .B(n5561), .Z(n5184) );
  AND U11699 ( .A(n5562), .B(n5563), .Z(n5560) );
  AND U11700 ( .A(b[48]), .B(a[64]), .Z(n5559) );
  XOR U11701 ( .A(n5564), .B(n5189), .Z(n5191) );
  XOR U11702 ( .A(n5565), .B(n5566), .Z(n5189) );
  AND U11703 ( .A(n5567), .B(n5568), .Z(n5565) );
  AND U11704 ( .A(b[47]), .B(a[65]), .Z(n5564) );
  XOR U11705 ( .A(n5569), .B(n5194), .Z(n5196) );
  XOR U11706 ( .A(n5570), .B(n5571), .Z(n5194) );
  AND U11707 ( .A(n5572), .B(n5573), .Z(n5570) );
  AND U11708 ( .A(b[46]), .B(a[66]), .Z(n5569) );
  XOR U11709 ( .A(n5574), .B(n5199), .Z(n5201) );
  XOR U11710 ( .A(n5575), .B(n5576), .Z(n5199) );
  AND U11711 ( .A(n5577), .B(n5578), .Z(n5575) );
  AND U11712 ( .A(b[45]), .B(a[67]), .Z(n5574) );
  XOR U11713 ( .A(n5579), .B(n5204), .Z(n5206) );
  XOR U11714 ( .A(n5580), .B(n5581), .Z(n5204) );
  AND U11715 ( .A(n5582), .B(n5583), .Z(n5580) );
  AND U11716 ( .A(b[44]), .B(a[68]), .Z(n5579) );
  XOR U11717 ( .A(n5584), .B(n5585), .Z(n5208) );
  AND U11718 ( .A(n5586), .B(n5587), .Z(n5584) );
  XOR U11719 ( .A(n5588), .B(n5213), .Z(n5215) );
  XOR U11720 ( .A(n5589), .B(n5590), .Z(n5213) );
  AND U11721 ( .A(n5591), .B(n5592), .Z(n5589) );
  AND U11722 ( .A(b[43]), .B(a[69]), .Z(n5588) );
  XOR U11723 ( .A(n5593), .B(n5218), .Z(n5220) );
  XOR U11724 ( .A(n5594), .B(n5595), .Z(n5218) );
  AND U11725 ( .A(n5596), .B(n5597), .Z(n5594) );
  AND U11726 ( .A(b[41]), .B(a[71]), .Z(n5593) );
  XOR U11727 ( .A(n5598), .B(n5223), .Z(n5225) );
  XOR U11728 ( .A(n5599), .B(n5600), .Z(n5223) );
  AND U11729 ( .A(n5601), .B(n5602), .Z(n5599) );
  AND U11730 ( .A(b[40]), .B(a[72]), .Z(n5598) );
  XOR U11731 ( .A(n5603), .B(n5228), .Z(n5230) );
  XOR U11732 ( .A(n5604), .B(n5605), .Z(n5228) );
  AND U11733 ( .A(n5606), .B(n5607), .Z(n5604) );
  AND U11734 ( .A(b[39]), .B(a[73]), .Z(n5603) );
  XOR U11735 ( .A(n5608), .B(n5233), .Z(n5235) );
  XOR U11736 ( .A(n5609), .B(n5610), .Z(n5233) );
  AND U11737 ( .A(n5611), .B(n5612), .Z(n5609) );
  AND U11738 ( .A(b[38]), .B(a[74]), .Z(n5608) );
  XOR U11739 ( .A(n5613), .B(n5614), .Z(n5237) );
  AND U11740 ( .A(n5615), .B(n5616), .Z(n5613) );
  XOR U11741 ( .A(n5617), .B(n5242), .Z(n5244) );
  XOR U11742 ( .A(n5618), .B(n5619), .Z(n5242) );
  AND U11743 ( .A(n5620), .B(n5621), .Z(n5618) );
  AND U11744 ( .A(b[37]), .B(a[75]), .Z(n5617) );
  XOR U11745 ( .A(n5622), .B(n5247), .Z(n5249) );
  XOR U11746 ( .A(n5623), .B(n5624), .Z(n5247) );
  AND U11747 ( .A(n5625), .B(n5626), .Z(n5623) );
  AND U11748 ( .A(b[35]), .B(a[77]), .Z(n5622) );
  XOR U11749 ( .A(n5627), .B(n5252), .Z(n5254) );
  XOR U11750 ( .A(n5628), .B(n5629), .Z(n5252) );
  AND U11751 ( .A(n5630), .B(n5631), .Z(n5628) );
  AND U11752 ( .A(b[34]), .B(a[78]), .Z(n5627) );
  XOR U11753 ( .A(n5632), .B(n5257), .Z(n5259) );
  XOR U11754 ( .A(n5633), .B(n5634), .Z(n5257) );
  AND U11755 ( .A(n5635), .B(n5636), .Z(n5633) );
  AND U11756 ( .A(b[33]), .B(a[79]), .Z(n5632) );
  XOR U11757 ( .A(n5637), .B(n5262), .Z(n5264) );
  XOR U11758 ( .A(n5638), .B(n5639), .Z(n5262) );
  AND U11759 ( .A(n5640), .B(n5641), .Z(n5638) );
  AND U11760 ( .A(b[32]), .B(a[80]), .Z(n5637) );
  XOR U11761 ( .A(n5642), .B(n5643), .Z(n5266) );
  AND U11762 ( .A(n5644), .B(n5645), .Z(n5642) );
  XOR U11763 ( .A(n5646), .B(n5271), .Z(n5273) );
  XOR U11764 ( .A(n5647), .B(n5648), .Z(n5271) );
  AND U11765 ( .A(n5649), .B(n5650), .Z(n5647) );
  AND U11766 ( .A(b[31]), .B(a[81]), .Z(n5646) );
  XOR U11767 ( .A(n5651), .B(n5276), .Z(n5278) );
  XOR U11768 ( .A(n5652), .B(n5653), .Z(n5276) );
  AND U11769 ( .A(n5654), .B(n5655), .Z(n5652) );
  AND U11770 ( .A(b[29]), .B(a[83]), .Z(n5651) );
  XOR U11771 ( .A(n5656), .B(n5281), .Z(n5283) );
  XOR U11772 ( .A(n5657), .B(n5658), .Z(n5281) );
  AND U11773 ( .A(n5659), .B(n5660), .Z(n5657) );
  AND U11774 ( .A(b[28]), .B(a[84]), .Z(n5656) );
  XOR U11775 ( .A(n5661), .B(n5286), .Z(n5288) );
  XOR U11776 ( .A(n5662), .B(n5663), .Z(n5286) );
  AND U11777 ( .A(n5664), .B(n5665), .Z(n5662) );
  AND U11778 ( .A(b[27]), .B(a[85]), .Z(n5661) );
  XOR U11779 ( .A(n5666), .B(n5291), .Z(n5293) );
  XOR U11780 ( .A(n5667), .B(n5668), .Z(n5291) );
  AND U11781 ( .A(n5669), .B(n5670), .Z(n5667) );
  AND U11782 ( .A(b[26]), .B(a[86]), .Z(n5666) );
  XOR U11783 ( .A(n5671), .B(n5672), .Z(n5295) );
  AND U11784 ( .A(n5673), .B(n5674), .Z(n5671) );
  XOR U11785 ( .A(n5675), .B(n5300), .Z(n5302) );
  XOR U11786 ( .A(n5676), .B(n5677), .Z(n5300) );
  AND U11787 ( .A(n5678), .B(n5679), .Z(n5676) );
  AND U11788 ( .A(b[25]), .B(a[87]), .Z(n5675) );
  XOR U11789 ( .A(n5680), .B(n5305), .Z(n5307) );
  XOR U11790 ( .A(n5681), .B(n5682), .Z(n5305) );
  AND U11791 ( .A(n5683), .B(n5684), .Z(n5681) );
  AND U11792 ( .A(b[23]), .B(a[89]), .Z(n5680) );
  XOR U11793 ( .A(n5685), .B(n5310), .Z(n5312) );
  XOR U11794 ( .A(n5686), .B(n5687), .Z(n5310) );
  AND U11795 ( .A(n5688), .B(n5689), .Z(n5686) );
  AND U11796 ( .A(b[22]), .B(a[90]), .Z(n5685) );
  XOR U11797 ( .A(n5690), .B(n5315), .Z(n5317) );
  XOR U11798 ( .A(n5691), .B(n5692), .Z(n5315) );
  AND U11799 ( .A(n5693), .B(n5694), .Z(n5691) );
  AND U11800 ( .A(b[21]), .B(a[91]), .Z(n5690) );
  XOR U11801 ( .A(n5695), .B(n5320), .Z(n5322) );
  XOR U11802 ( .A(n5696), .B(n5697), .Z(n5320) );
  AND U11803 ( .A(n5698), .B(n5699), .Z(n5696) );
  AND U11804 ( .A(b[20]), .B(a[92]), .Z(n5695) );
  XOR U11805 ( .A(n5700), .B(n5701), .Z(n5324) );
  AND U11806 ( .A(n5702), .B(n5703), .Z(n5700) );
  XOR U11807 ( .A(n5704), .B(n5329), .Z(n5331) );
  XOR U11808 ( .A(n5705), .B(n5706), .Z(n5329) );
  AND U11809 ( .A(n5707), .B(n5708), .Z(n5705) );
  AND U11810 ( .A(b[19]), .B(a[93]), .Z(n5704) );
  XOR U11811 ( .A(n5709), .B(n5334), .Z(n5336) );
  XOR U11812 ( .A(n5710), .B(n5711), .Z(n5334) );
  AND U11813 ( .A(n5712), .B(n5713), .Z(n5710) );
  AND U11814 ( .A(b[17]), .B(a[95]), .Z(n5709) );
  XOR U11815 ( .A(n5714), .B(n5339), .Z(n5341) );
  XOR U11816 ( .A(n5715), .B(n5716), .Z(n5339) );
  AND U11817 ( .A(n5717), .B(n5718), .Z(n5715) );
  AND U11818 ( .A(b[16]), .B(a[96]), .Z(n5714) );
  XOR U11819 ( .A(n5719), .B(n5344), .Z(n5346) );
  XOR U11820 ( .A(n5720), .B(n5721), .Z(n5344) );
  AND U11821 ( .A(n5722), .B(n5723), .Z(n5720) );
  AND U11822 ( .A(b[15]), .B(a[97]), .Z(n5719) );
  XOR U11823 ( .A(n5724), .B(n5349), .Z(n5351) );
  XOR U11824 ( .A(n5725), .B(n5726), .Z(n5349) );
  AND U11825 ( .A(n5727), .B(n5728), .Z(n5725) );
  AND U11826 ( .A(b[14]), .B(a[98]), .Z(n5724) );
  XOR U11827 ( .A(n5729), .B(n5730), .Z(n5353) );
  AND U11828 ( .A(n5731), .B(n5732), .Z(n5729) );
  XOR U11829 ( .A(n5733), .B(n5358), .Z(n5360) );
  XOR U11830 ( .A(n5734), .B(n5735), .Z(n5358) );
  AND U11831 ( .A(n5736), .B(n5737), .Z(n5734) );
  AND U11832 ( .A(b[13]), .B(a[99]), .Z(n5733) );
  XOR U11833 ( .A(n5738), .B(n5363), .Z(n5365) );
  XOR U11834 ( .A(n5739), .B(n5740), .Z(n5363) );
  AND U11835 ( .A(n5741), .B(n5742), .Z(n5739) );
  AND U11836 ( .A(b[11]), .B(a[101]), .Z(n5738) );
  XOR U11837 ( .A(n5743), .B(n5368), .Z(n5370) );
  XOR U11838 ( .A(n5744), .B(n5745), .Z(n5368) );
  AND U11839 ( .A(n5746), .B(n5747), .Z(n5744) );
  AND U11840 ( .A(b[10]), .B(a[102]), .Z(n5743) );
  XOR U11841 ( .A(n5748), .B(n5373), .Z(n5375) );
  XOR U11842 ( .A(n5749), .B(n5750), .Z(n5373) );
  AND U11843 ( .A(n5751), .B(n5752), .Z(n5749) );
  AND U11844 ( .A(b[9]), .B(a[103]), .Z(n5748) );
  XOR U11845 ( .A(n5753), .B(n5378), .Z(n5380) );
  XOR U11846 ( .A(n5754), .B(n5755), .Z(n5378) );
  AND U11847 ( .A(n5756), .B(n5757), .Z(n5754) );
  AND U11848 ( .A(b[8]), .B(a[104]), .Z(n5753) );
  XOR U11849 ( .A(n5758), .B(n5759), .Z(n5382) );
  AND U11850 ( .A(n5760), .B(n5761), .Z(n5758) );
  XOR U11851 ( .A(n5762), .B(n5387), .Z(n5389) );
  XOR U11852 ( .A(n5763), .B(n5764), .Z(n5387) );
  AND U11853 ( .A(n5765), .B(n5766), .Z(n5763) );
  AND U11854 ( .A(b[7]), .B(a[105]), .Z(n5762) );
  XOR U11855 ( .A(n5767), .B(n5392), .Z(n5394) );
  XOR U11856 ( .A(n5768), .B(n5769), .Z(n5392) );
  AND U11857 ( .A(n5770), .B(n5771), .Z(n5768) );
  AND U11858 ( .A(b[5]), .B(a[107]), .Z(n5767) );
  XOR U11859 ( .A(n5772), .B(n5397), .Z(n5399) );
  XOR U11860 ( .A(n5773), .B(n5774), .Z(n5397) );
  AND U11861 ( .A(n5775), .B(n5776), .Z(n5773) );
  AND U11862 ( .A(b[4]), .B(a[108]), .Z(n5772) );
  XNOR U11863 ( .A(n5777), .B(n5778), .Z(n5411) );
  NANDN U11864 ( .A(n5779), .B(n5780), .Z(n5778) );
  XOR U11865 ( .A(n5781), .B(n5402), .Z(n5404) );
  XNOR U11866 ( .A(n5782), .B(n5783), .Z(n5402) );
  AND U11867 ( .A(n5784), .B(n5785), .Z(n5782) );
  AND U11868 ( .A(b[3]), .B(a[109]), .Z(n5781) );
  XNOR U11869 ( .A(n5786), .B(n5787), .Z(swire[111]) );
  XOR U11870 ( .A(n5420), .B(n5788), .Z(n5787) );
  NAND U11871 ( .A(a[111]), .B(b[0]), .Z(n5421) );
  XNOR U11872 ( .A(n5779), .B(n5780), .Z(n5420) );
  XOR U11873 ( .A(n5777), .B(n5789), .Z(n5780) );
  NAND U11874 ( .A(b[1]), .B(a[110]), .Z(n5789) );
  XOR U11875 ( .A(n5785), .B(n5790), .Z(n5779) );
  XOR U11876 ( .A(n5777), .B(n5784), .Z(n5790) );
  XNOR U11877 ( .A(n5791), .B(n5783), .Z(n5784) );
  AND U11878 ( .A(b[2]), .B(a[109]), .Z(n5791) );
  NANDN U11879 ( .A(n5792), .B(n5793), .Z(n5777) );
  XOR U11880 ( .A(n5783), .B(n5775), .Z(n5794) );
  XNOR U11881 ( .A(n5774), .B(n5770), .Z(n5795) );
  XNOR U11882 ( .A(n5761), .B(n5760), .Z(n5796) );
  XOR U11883 ( .A(n5797), .B(n5759), .Z(n5760) );
  AND U11884 ( .A(b[5]), .B(a[106]), .Z(n5797) );
  XNOR U11885 ( .A(n5759), .B(n5765), .Z(n5798) );
  XNOR U11886 ( .A(n5764), .B(n5756), .Z(n5799) );
  XNOR U11887 ( .A(n5755), .B(n5751), .Z(n5800) );
  XNOR U11888 ( .A(n5750), .B(n5746), .Z(n5801) );
  XNOR U11889 ( .A(n5745), .B(n5741), .Z(n5802) );
  XNOR U11890 ( .A(n5732), .B(n5731), .Z(n5803) );
  XOR U11891 ( .A(n5804), .B(n5730), .Z(n5731) );
  AND U11892 ( .A(b[11]), .B(a[100]), .Z(n5804) );
  XNOR U11893 ( .A(n5730), .B(n5736), .Z(n5805) );
  XNOR U11894 ( .A(n5735), .B(n5727), .Z(n5806) );
  XNOR U11895 ( .A(n5726), .B(n5722), .Z(n5807) );
  XNOR U11896 ( .A(n5721), .B(n5717), .Z(n5808) );
  XNOR U11897 ( .A(n5716), .B(n5712), .Z(n5809) );
  XNOR U11898 ( .A(n5703), .B(n5702), .Z(n5810) );
  XOR U11899 ( .A(n5811), .B(n5701), .Z(n5702) );
  AND U11900 ( .A(b[17]), .B(a[94]), .Z(n5811) );
  XNOR U11901 ( .A(n5701), .B(n5707), .Z(n5812) );
  XNOR U11902 ( .A(n5706), .B(n5698), .Z(n5813) );
  XNOR U11903 ( .A(n5697), .B(n5693), .Z(n5814) );
  XNOR U11904 ( .A(n5692), .B(n5688), .Z(n5815) );
  XNOR U11905 ( .A(n5687), .B(n5683), .Z(n5816) );
  XNOR U11906 ( .A(n5674), .B(n5673), .Z(n5817) );
  XOR U11907 ( .A(n5818), .B(n5672), .Z(n5673) );
  AND U11908 ( .A(b[23]), .B(a[88]), .Z(n5818) );
  XNOR U11909 ( .A(n5672), .B(n5678), .Z(n5819) );
  XNOR U11910 ( .A(n5677), .B(n5669), .Z(n5820) );
  XNOR U11911 ( .A(n5668), .B(n5664), .Z(n5821) );
  XNOR U11912 ( .A(n5663), .B(n5659), .Z(n5822) );
  XNOR U11913 ( .A(n5658), .B(n5654), .Z(n5823) );
  XNOR U11914 ( .A(n5645), .B(n5644), .Z(n5824) );
  XOR U11915 ( .A(n5825), .B(n5643), .Z(n5644) );
  AND U11916 ( .A(b[29]), .B(a[82]), .Z(n5825) );
  XNOR U11917 ( .A(n5643), .B(n5649), .Z(n5826) );
  XNOR U11918 ( .A(n5648), .B(n5640), .Z(n5827) );
  XNOR U11919 ( .A(n5639), .B(n5635), .Z(n5828) );
  XNOR U11920 ( .A(n5634), .B(n5630), .Z(n5829) );
  XNOR U11921 ( .A(n5629), .B(n5625), .Z(n5830) );
  XNOR U11922 ( .A(n5616), .B(n5615), .Z(n5831) );
  XOR U11923 ( .A(n5832), .B(n5614), .Z(n5615) );
  AND U11924 ( .A(b[35]), .B(a[76]), .Z(n5832) );
  XNOR U11925 ( .A(n5614), .B(n5620), .Z(n5833) );
  XNOR U11926 ( .A(n5619), .B(n5611), .Z(n5834) );
  XNOR U11927 ( .A(n5610), .B(n5606), .Z(n5835) );
  XNOR U11928 ( .A(n5605), .B(n5601), .Z(n5836) );
  XNOR U11929 ( .A(n5600), .B(n5596), .Z(n5837) );
  XNOR U11930 ( .A(n5587), .B(n5586), .Z(n5838) );
  XOR U11931 ( .A(n5839), .B(n5585), .Z(n5586) );
  AND U11932 ( .A(b[41]), .B(a[70]), .Z(n5839) );
  XNOR U11933 ( .A(n5585), .B(n5591), .Z(n5840) );
  XNOR U11934 ( .A(n5590), .B(n5582), .Z(n5841) );
  XNOR U11935 ( .A(n5581), .B(n5577), .Z(n5842) );
  XNOR U11936 ( .A(n5576), .B(n5572), .Z(n5843) );
  XNOR U11937 ( .A(n5571), .B(n5567), .Z(n5844) );
  XNOR U11938 ( .A(n5566), .B(n5562), .Z(n5845) );
  XNOR U11939 ( .A(n5561), .B(n5557), .Z(n5846) );
  XNOR U11940 ( .A(n5556), .B(n5552), .Z(n5847) );
  XNOR U11941 ( .A(n5551), .B(n5547), .Z(n5848) );
  XNOR U11942 ( .A(n5546), .B(n5542), .Z(n5849) );
  XNOR U11943 ( .A(n5541), .B(n5537), .Z(n5850) );
  XNOR U11944 ( .A(n5536), .B(n5532), .Z(n5851) );
  XNOR U11945 ( .A(n5531), .B(n5527), .Z(n5852) );
  XNOR U11946 ( .A(n5526), .B(n5522), .Z(n5853) );
  XNOR U11947 ( .A(n5521), .B(n5517), .Z(n5854) );
  XNOR U11948 ( .A(n5516), .B(n5512), .Z(n5855) );
  XNOR U11949 ( .A(n5511), .B(n5507), .Z(n5856) );
  XNOR U11950 ( .A(n5506), .B(n5502), .Z(n5857) );
  XOR U11951 ( .A(n5501), .B(n5498), .Z(n5858) );
  XOR U11952 ( .A(n5859), .B(n5860), .Z(n5498) );
  XOR U11953 ( .A(n5496), .B(n5861), .Z(n5860) );
  XOR U11954 ( .A(n5862), .B(n5863), .Z(n5861) );
  XOR U11955 ( .A(n5864), .B(n5865), .Z(n5863) );
  NAND U11956 ( .A(a[49]), .B(b[62]), .Z(n5865) );
  AND U11957 ( .A(a[48]), .B(b[63]), .Z(n5864) );
  XOR U11958 ( .A(n5866), .B(n5862), .Z(n5859) );
  XOR U11959 ( .A(n5867), .B(n5868), .Z(n5862) );
  ANDN U11960 ( .B(n5869), .A(n5870), .Z(n5867) );
  AND U11961 ( .A(a[50]), .B(b[61]), .Z(n5866) );
  XOR U11962 ( .A(n5871), .B(n5496), .Z(n5497) );
  XOR U11963 ( .A(n5872), .B(n5873), .Z(n5496) );
  AND U11964 ( .A(n5874), .B(n5875), .Z(n5872) );
  AND U11965 ( .A(a[51]), .B(b[60]), .Z(n5871) );
  XOR U11966 ( .A(n5876), .B(n5501), .Z(n5503) );
  XOR U11967 ( .A(n5877), .B(n5878), .Z(n5501) );
  AND U11968 ( .A(n5879), .B(n5880), .Z(n5877) );
  AND U11969 ( .A(a[52]), .B(b[59]), .Z(n5876) );
  XOR U11970 ( .A(n5881), .B(n5506), .Z(n5508) );
  XOR U11971 ( .A(n5882), .B(n5883), .Z(n5506) );
  AND U11972 ( .A(n5884), .B(n5885), .Z(n5882) );
  AND U11973 ( .A(a[53]), .B(b[58]), .Z(n5881) );
  XOR U11974 ( .A(n5886), .B(n5511), .Z(n5513) );
  XOR U11975 ( .A(n5887), .B(n5888), .Z(n5511) );
  AND U11976 ( .A(n5889), .B(n5890), .Z(n5887) );
  AND U11977 ( .A(a[54]), .B(b[57]), .Z(n5886) );
  XOR U11978 ( .A(n5891), .B(n5516), .Z(n5518) );
  XOR U11979 ( .A(n5892), .B(n5893), .Z(n5516) );
  AND U11980 ( .A(n5894), .B(n5895), .Z(n5892) );
  AND U11981 ( .A(a[55]), .B(b[56]), .Z(n5891) );
  XOR U11982 ( .A(n5896), .B(n5521), .Z(n5523) );
  XOR U11983 ( .A(n5897), .B(n5898), .Z(n5521) );
  AND U11984 ( .A(n5899), .B(n5900), .Z(n5897) );
  AND U11985 ( .A(b[55]), .B(a[56]), .Z(n5896) );
  XOR U11986 ( .A(n5901), .B(n5526), .Z(n5528) );
  XOR U11987 ( .A(n5902), .B(n5903), .Z(n5526) );
  AND U11988 ( .A(n5904), .B(n5905), .Z(n5902) );
  AND U11989 ( .A(b[54]), .B(a[57]), .Z(n5901) );
  XOR U11990 ( .A(n5906), .B(n5531), .Z(n5533) );
  XOR U11991 ( .A(n5907), .B(n5908), .Z(n5531) );
  AND U11992 ( .A(n5909), .B(n5910), .Z(n5907) );
  AND U11993 ( .A(b[53]), .B(a[58]), .Z(n5906) );
  XOR U11994 ( .A(n5911), .B(n5536), .Z(n5538) );
  XOR U11995 ( .A(n5912), .B(n5913), .Z(n5536) );
  AND U11996 ( .A(n5914), .B(n5915), .Z(n5912) );
  AND U11997 ( .A(b[52]), .B(a[59]), .Z(n5911) );
  XOR U11998 ( .A(n5916), .B(n5541), .Z(n5543) );
  XOR U11999 ( .A(n5917), .B(n5918), .Z(n5541) );
  AND U12000 ( .A(n5919), .B(n5920), .Z(n5917) );
  AND U12001 ( .A(b[51]), .B(a[60]), .Z(n5916) );
  XOR U12002 ( .A(n5921), .B(n5546), .Z(n5548) );
  XOR U12003 ( .A(n5922), .B(n5923), .Z(n5546) );
  AND U12004 ( .A(n5924), .B(n5925), .Z(n5922) );
  AND U12005 ( .A(b[50]), .B(a[61]), .Z(n5921) );
  XOR U12006 ( .A(n5926), .B(n5551), .Z(n5553) );
  XOR U12007 ( .A(n5927), .B(n5928), .Z(n5551) );
  AND U12008 ( .A(n5929), .B(n5930), .Z(n5927) );
  AND U12009 ( .A(b[49]), .B(a[62]), .Z(n5926) );
  XOR U12010 ( .A(n5931), .B(n5556), .Z(n5558) );
  XOR U12011 ( .A(n5932), .B(n5933), .Z(n5556) );
  AND U12012 ( .A(n5934), .B(n5935), .Z(n5932) );
  AND U12013 ( .A(b[48]), .B(a[63]), .Z(n5931) );
  XOR U12014 ( .A(n5936), .B(n5561), .Z(n5563) );
  XOR U12015 ( .A(n5937), .B(n5938), .Z(n5561) );
  AND U12016 ( .A(n5939), .B(n5940), .Z(n5937) );
  AND U12017 ( .A(b[47]), .B(a[64]), .Z(n5936) );
  XOR U12018 ( .A(n5941), .B(n5566), .Z(n5568) );
  XOR U12019 ( .A(n5942), .B(n5943), .Z(n5566) );
  AND U12020 ( .A(n5944), .B(n5945), .Z(n5942) );
  AND U12021 ( .A(b[46]), .B(a[65]), .Z(n5941) );
  XOR U12022 ( .A(n5946), .B(n5571), .Z(n5573) );
  XOR U12023 ( .A(n5947), .B(n5948), .Z(n5571) );
  AND U12024 ( .A(n5949), .B(n5950), .Z(n5947) );
  AND U12025 ( .A(b[45]), .B(a[66]), .Z(n5946) );
  XOR U12026 ( .A(n5951), .B(n5576), .Z(n5578) );
  XOR U12027 ( .A(n5952), .B(n5953), .Z(n5576) );
  AND U12028 ( .A(n5954), .B(n5955), .Z(n5952) );
  AND U12029 ( .A(b[44]), .B(a[67]), .Z(n5951) );
  XOR U12030 ( .A(n5956), .B(n5581), .Z(n5583) );
  XOR U12031 ( .A(n5957), .B(n5958), .Z(n5581) );
  AND U12032 ( .A(n5959), .B(n5960), .Z(n5957) );
  AND U12033 ( .A(b[43]), .B(a[68]), .Z(n5956) );
  XOR U12034 ( .A(n5961), .B(n5962), .Z(n5585) );
  AND U12035 ( .A(n5963), .B(n5964), .Z(n5961) );
  XOR U12036 ( .A(n5965), .B(n5590), .Z(n5592) );
  XOR U12037 ( .A(n5966), .B(n5967), .Z(n5590) );
  AND U12038 ( .A(n5968), .B(n5969), .Z(n5966) );
  AND U12039 ( .A(b[42]), .B(a[69]), .Z(n5965) );
  XOR U12040 ( .A(n5970), .B(n5595), .Z(n5597) );
  XOR U12041 ( .A(n5971), .B(n5972), .Z(n5595) );
  AND U12042 ( .A(n5973), .B(n5974), .Z(n5971) );
  AND U12043 ( .A(b[40]), .B(a[71]), .Z(n5970) );
  XOR U12044 ( .A(n5975), .B(n5600), .Z(n5602) );
  XOR U12045 ( .A(n5976), .B(n5977), .Z(n5600) );
  AND U12046 ( .A(n5978), .B(n5979), .Z(n5976) );
  AND U12047 ( .A(b[39]), .B(a[72]), .Z(n5975) );
  XOR U12048 ( .A(n5980), .B(n5605), .Z(n5607) );
  XOR U12049 ( .A(n5981), .B(n5982), .Z(n5605) );
  AND U12050 ( .A(n5983), .B(n5984), .Z(n5981) );
  AND U12051 ( .A(b[38]), .B(a[73]), .Z(n5980) );
  XOR U12052 ( .A(n5985), .B(n5610), .Z(n5612) );
  XOR U12053 ( .A(n5986), .B(n5987), .Z(n5610) );
  AND U12054 ( .A(n5988), .B(n5989), .Z(n5986) );
  AND U12055 ( .A(b[37]), .B(a[74]), .Z(n5985) );
  XOR U12056 ( .A(n5990), .B(n5991), .Z(n5614) );
  AND U12057 ( .A(n5992), .B(n5993), .Z(n5990) );
  XOR U12058 ( .A(n5994), .B(n5619), .Z(n5621) );
  XOR U12059 ( .A(n5995), .B(n5996), .Z(n5619) );
  AND U12060 ( .A(n5997), .B(n5998), .Z(n5995) );
  AND U12061 ( .A(b[36]), .B(a[75]), .Z(n5994) );
  XOR U12062 ( .A(n5999), .B(n5624), .Z(n5626) );
  XOR U12063 ( .A(n6000), .B(n6001), .Z(n5624) );
  AND U12064 ( .A(n6002), .B(n6003), .Z(n6000) );
  AND U12065 ( .A(b[34]), .B(a[77]), .Z(n5999) );
  XOR U12066 ( .A(n6004), .B(n5629), .Z(n5631) );
  XOR U12067 ( .A(n6005), .B(n6006), .Z(n5629) );
  AND U12068 ( .A(n6007), .B(n6008), .Z(n6005) );
  AND U12069 ( .A(b[33]), .B(a[78]), .Z(n6004) );
  XOR U12070 ( .A(n6009), .B(n5634), .Z(n5636) );
  XOR U12071 ( .A(n6010), .B(n6011), .Z(n5634) );
  AND U12072 ( .A(n6012), .B(n6013), .Z(n6010) );
  AND U12073 ( .A(b[32]), .B(a[79]), .Z(n6009) );
  XOR U12074 ( .A(n6014), .B(n5639), .Z(n5641) );
  XOR U12075 ( .A(n6015), .B(n6016), .Z(n5639) );
  AND U12076 ( .A(n6017), .B(n6018), .Z(n6015) );
  AND U12077 ( .A(b[31]), .B(a[80]), .Z(n6014) );
  XOR U12078 ( .A(n6019), .B(n6020), .Z(n5643) );
  AND U12079 ( .A(n6021), .B(n6022), .Z(n6019) );
  XOR U12080 ( .A(n6023), .B(n5648), .Z(n5650) );
  XOR U12081 ( .A(n6024), .B(n6025), .Z(n5648) );
  AND U12082 ( .A(n6026), .B(n6027), .Z(n6024) );
  AND U12083 ( .A(b[30]), .B(a[81]), .Z(n6023) );
  XOR U12084 ( .A(n6028), .B(n5653), .Z(n5655) );
  XOR U12085 ( .A(n6029), .B(n6030), .Z(n5653) );
  AND U12086 ( .A(n6031), .B(n6032), .Z(n6029) );
  AND U12087 ( .A(b[28]), .B(a[83]), .Z(n6028) );
  XOR U12088 ( .A(n6033), .B(n5658), .Z(n5660) );
  XOR U12089 ( .A(n6034), .B(n6035), .Z(n5658) );
  AND U12090 ( .A(n6036), .B(n6037), .Z(n6034) );
  AND U12091 ( .A(b[27]), .B(a[84]), .Z(n6033) );
  XOR U12092 ( .A(n6038), .B(n5663), .Z(n5665) );
  XOR U12093 ( .A(n6039), .B(n6040), .Z(n5663) );
  AND U12094 ( .A(n6041), .B(n6042), .Z(n6039) );
  AND U12095 ( .A(b[26]), .B(a[85]), .Z(n6038) );
  XOR U12096 ( .A(n6043), .B(n5668), .Z(n5670) );
  XOR U12097 ( .A(n6044), .B(n6045), .Z(n5668) );
  AND U12098 ( .A(n6046), .B(n6047), .Z(n6044) );
  AND U12099 ( .A(b[25]), .B(a[86]), .Z(n6043) );
  XOR U12100 ( .A(n6048), .B(n6049), .Z(n5672) );
  AND U12101 ( .A(n6050), .B(n6051), .Z(n6048) );
  XOR U12102 ( .A(n6052), .B(n5677), .Z(n5679) );
  XOR U12103 ( .A(n6053), .B(n6054), .Z(n5677) );
  AND U12104 ( .A(n6055), .B(n6056), .Z(n6053) );
  AND U12105 ( .A(b[24]), .B(a[87]), .Z(n6052) );
  XOR U12106 ( .A(n6057), .B(n5682), .Z(n5684) );
  XOR U12107 ( .A(n6058), .B(n6059), .Z(n5682) );
  AND U12108 ( .A(n6060), .B(n6061), .Z(n6058) );
  AND U12109 ( .A(b[22]), .B(a[89]), .Z(n6057) );
  XOR U12110 ( .A(n6062), .B(n5687), .Z(n5689) );
  XOR U12111 ( .A(n6063), .B(n6064), .Z(n5687) );
  AND U12112 ( .A(n6065), .B(n6066), .Z(n6063) );
  AND U12113 ( .A(b[21]), .B(a[90]), .Z(n6062) );
  XOR U12114 ( .A(n6067), .B(n5692), .Z(n5694) );
  XOR U12115 ( .A(n6068), .B(n6069), .Z(n5692) );
  AND U12116 ( .A(n6070), .B(n6071), .Z(n6068) );
  AND U12117 ( .A(b[20]), .B(a[91]), .Z(n6067) );
  XOR U12118 ( .A(n6072), .B(n5697), .Z(n5699) );
  XOR U12119 ( .A(n6073), .B(n6074), .Z(n5697) );
  AND U12120 ( .A(n6075), .B(n6076), .Z(n6073) );
  AND U12121 ( .A(b[19]), .B(a[92]), .Z(n6072) );
  XOR U12122 ( .A(n6077), .B(n6078), .Z(n5701) );
  AND U12123 ( .A(n6079), .B(n6080), .Z(n6077) );
  XOR U12124 ( .A(n6081), .B(n5706), .Z(n5708) );
  XOR U12125 ( .A(n6082), .B(n6083), .Z(n5706) );
  AND U12126 ( .A(n6084), .B(n6085), .Z(n6082) );
  AND U12127 ( .A(b[18]), .B(a[93]), .Z(n6081) );
  XOR U12128 ( .A(n6086), .B(n5711), .Z(n5713) );
  XOR U12129 ( .A(n6087), .B(n6088), .Z(n5711) );
  AND U12130 ( .A(n6089), .B(n6090), .Z(n6087) );
  AND U12131 ( .A(b[16]), .B(a[95]), .Z(n6086) );
  XOR U12132 ( .A(n6091), .B(n5716), .Z(n5718) );
  XOR U12133 ( .A(n6092), .B(n6093), .Z(n5716) );
  AND U12134 ( .A(n6094), .B(n6095), .Z(n6092) );
  AND U12135 ( .A(b[15]), .B(a[96]), .Z(n6091) );
  XOR U12136 ( .A(n6096), .B(n5721), .Z(n5723) );
  XOR U12137 ( .A(n6097), .B(n6098), .Z(n5721) );
  AND U12138 ( .A(n6099), .B(n6100), .Z(n6097) );
  AND U12139 ( .A(b[14]), .B(a[97]), .Z(n6096) );
  XOR U12140 ( .A(n6101), .B(n5726), .Z(n5728) );
  XOR U12141 ( .A(n6102), .B(n6103), .Z(n5726) );
  AND U12142 ( .A(n6104), .B(n6105), .Z(n6102) );
  AND U12143 ( .A(b[13]), .B(a[98]), .Z(n6101) );
  XOR U12144 ( .A(n6106), .B(n6107), .Z(n5730) );
  AND U12145 ( .A(n6108), .B(n6109), .Z(n6106) );
  XOR U12146 ( .A(n6110), .B(n5735), .Z(n5737) );
  XOR U12147 ( .A(n6111), .B(n6112), .Z(n5735) );
  AND U12148 ( .A(n6113), .B(n6114), .Z(n6111) );
  AND U12149 ( .A(b[12]), .B(a[99]), .Z(n6110) );
  XOR U12150 ( .A(n6115), .B(n5740), .Z(n5742) );
  XOR U12151 ( .A(n6116), .B(n6117), .Z(n5740) );
  AND U12152 ( .A(n6118), .B(n6119), .Z(n6116) );
  AND U12153 ( .A(b[10]), .B(a[101]), .Z(n6115) );
  XOR U12154 ( .A(n6120), .B(n5745), .Z(n5747) );
  XOR U12155 ( .A(n6121), .B(n6122), .Z(n5745) );
  AND U12156 ( .A(n6123), .B(n6124), .Z(n6121) );
  AND U12157 ( .A(b[9]), .B(a[102]), .Z(n6120) );
  XOR U12158 ( .A(n6125), .B(n5750), .Z(n5752) );
  XOR U12159 ( .A(n6126), .B(n6127), .Z(n5750) );
  AND U12160 ( .A(n6128), .B(n6129), .Z(n6126) );
  AND U12161 ( .A(b[8]), .B(a[103]), .Z(n6125) );
  XOR U12162 ( .A(n6130), .B(n5755), .Z(n5757) );
  XOR U12163 ( .A(n6131), .B(n6132), .Z(n5755) );
  AND U12164 ( .A(n6133), .B(n6134), .Z(n6131) );
  AND U12165 ( .A(b[7]), .B(a[104]), .Z(n6130) );
  XOR U12166 ( .A(n6135), .B(n6136), .Z(n5759) );
  AND U12167 ( .A(n6137), .B(n6138), .Z(n6135) );
  XOR U12168 ( .A(n6139), .B(n5764), .Z(n5766) );
  XOR U12169 ( .A(n6140), .B(n6141), .Z(n5764) );
  AND U12170 ( .A(n6142), .B(n6143), .Z(n6140) );
  AND U12171 ( .A(b[6]), .B(a[105]), .Z(n6139) );
  XOR U12172 ( .A(n6144), .B(n5769), .Z(n5771) );
  XOR U12173 ( .A(n6145), .B(n6146), .Z(n5769) );
  AND U12174 ( .A(n6147), .B(n6148), .Z(n6145) );
  AND U12175 ( .A(b[4]), .B(a[107]), .Z(n6144) );
  XNOR U12176 ( .A(n6149), .B(n6150), .Z(n5783) );
  NANDN U12177 ( .A(n6151), .B(n6152), .Z(n6150) );
  XOR U12178 ( .A(n6153), .B(n5774), .Z(n5776) );
  XNOR U12179 ( .A(n6154), .B(n6155), .Z(n5774) );
  AND U12180 ( .A(n6156), .B(n6157), .Z(n6154) );
  AND U12181 ( .A(b[3]), .B(a[108]), .Z(n6153) );
  XNOR U12182 ( .A(n6158), .B(n6159), .Z(swire[110]) );
  XOR U12183 ( .A(n5793), .B(n6160), .Z(n6159) );
  NAND U12184 ( .A(a[110]), .B(b[0]), .Z(n5792) );
  XNOR U12185 ( .A(n6151), .B(n6152), .Z(n5793) );
  XOR U12186 ( .A(n6149), .B(n6161), .Z(n6152) );
  NAND U12187 ( .A(b[1]), .B(a[109]), .Z(n6161) );
  XOR U12188 ( .A(n6157), .B(n6162), .Z(n6151) );
  XOR U12189 ( .A(n6149), .B(n6156), .Z(n6162) );
  XNOR U12190 ( .A(n6163), .B(n6155), .Z(n6156) );
  AND U12191 ( .A(b[2]), .B(a[108]), .Z(n6163) );
  NANDN U12192 ( .A(n6164), .B(n6165), .Z(n6149) );
  XOR U12193 ( .A(n6155), .B(n6147), .Z(n6166) );
  XNOR U12194 ( .A(n6138), .B(n6137), .Z(n6167) );
  XOR U12195 ( .A(n6168), .B(n6136), .Z(n6137) );
  AND U12196 ( .A(b[4]), .B(a[106]), .Z(n6168) );
  XNOR U12197 ( .A(n6136), .B(n6142), .Z(n6169) );
  XNOR U12198 ( .A(n6141), .B(n6133), .Z(n6170) );
  XNOR U12199 ( .A(n6132), .B(n6128), .Z(n6171) );
  XNOR U12200 ( .A(n6127), .B(n6123), .Z(n6172) );
  XNOR U12201 ( .A(n6122), .B(n6118), .Z(n6173) );
  XNOR U12202 ( .A(n6109), .B(n6108), .Z(n6174) );
  XOR U12203 ( .A(n6175), .B(n6107), .Z(n6108) );
  AND U12204 ( .A(b[10]), .B(a[100]), .Z(n6175) );
  XNOR U12205 ( .A(n6107), .B(n6113), .Z(n6176) );
  XNOR U12206 ( .A(n6112), .B(n6104), .Z(n6177) );
  XNOR U12207 ( .A(n6103), .B(n6099), .Z(n6178) );
  XNOR U12208 ( .A(n6098), .B(n6094), .Z(n6179) );
  XNOR U12209 ( .A(n6093), .B(n6089), .Z(n6180) );
  XNOR U12210 ( .A(n6080), .B(n6079), .Z(n6181) );
  XOR U12211 ( .A(n6182), .B(n6078), .Z(n6079) );
  AND U12212 ( .A(b[16]), .B(a[94]), .Z(n6182) );
  XNOR U12213 ( .A(n6078), .B(n6084), .Z(n6183) );
  XNOR U12214 ( .A(n6083), .B(n6075), .Z(n6184) );
  XNOR U12215 ( .A(n6074), .B(n6070), .Z(n6185) );
  XNOR U12216 ( .A(n6069), .B(n6065), .Z(n6186) );
  XNOR U12217 ( .A(n6064), .B(n6060), .Z(n6187) );
  XNOR U12218 ( .A(n6051), .B(n6050), .Z(n6188) );
  XOR U12219 ( .A(n6189), .B(n6049), .Z(n6050) );
  AND U12220 ( .A(b[22]), .B(a[88]), .Z(n6189) );
  XNOR U12221 ( .A(n6049), .B(n6055), .Z(n6190) );
  XNOR U12222 ( .A(n6054), .B(n6046), .Z(n6191) );
  XNOR U12223 ( .A(n6045), .B(n6041), .Z(n6192) );
  XNOR U12224 ( .A(n6040), .B(n6036), .Z(n6193) );
  XNOR U12225 ( .A(n6035), .B(n6031), .Z(n6194) );
  XNOR U12226 ( .A(n6022), .B(n6021), .Z(n6195) );
  XOR U12227 ( .A(n6196), .B(n6020), .Z(n6021) );
  AND U12228 ( .A(b[28]), .B(a[82]), .Z(n6196) );
  XNOR U12229 ( .A(n6020), .B(n6026), .Z(n6197) );
  XNOR U12230 ( .A(n6025), .B(n6017), .Z(n6198) );
  XNOR U12231 ( .A(n6016), .B(n6012), .Z(n6199) );
  XNOR U12232 ( .A(n6011), .B(n6007), .Z(n6200) );
  XNOR U12233 ( .A(n6006), .B(n6002), .Z(n6201) );
  XNOR U12234 ( .A(n5993), .B(n5992), .Z(n6202) );
  XOR U12235 ( .A(n6203), .B(n5991), .Z(n5992) );
  AND U12236 ( .A(b[34]), .B(a[76]), .Z(n6203) );
  XNOR U12237 ( .A(n5991), .B(n5997), .Z(n6204) );
  XNOR U12238 ( .A(n5996), .B(n5988), .Z(n6205) );
  XNOR U12239 ( .A(n5987), .B(n5983), .Z(n6206) );
  XNOR U12240 ( .A(n5982), .B(n5978), .Z(n6207) );
  XNOR U12241 ( .A(n5977), .B(n5973), .Z(n6208) );
  XNOR U12242 ( .A(n5964), .B(n5963), .Z(n6209) );
  XOR U12243 ( .A(n6210), .B(n5962), .Z(n5963) );
  AND U12244 ( .A(b[40]), .B(a[70]), .Z(n6210) );
  XNOR U12245 ( .A(n5962), .B(n5968), .Z(n6211) );
  XNOR U12246 ( .A(n5967), .B(n5959), .Z(n6212) );
  XNOR U12247 ( .A(n5958), .B(n5954), .Z(n6213) );
  XNOR U12248 ( .A(n5953), .B(n5949), .Z(n6214) );
  XNOR U12249 ( .A(n5948), .B(n5944), .Z(n6215) );
  XNOR U12250 ( .A(n5943), .B(n5939), .Z(n6216) );
  XNOR U12251 ( .A(n5938), .B(n5934), .Z(n6217) );
  XNOR U12252 ( .A(n5933), .B(n5929), .Z(n6218) );
  XNOR U12253 ( .A(n5928), .B(n5924), .Z(n6219) );
  XNOR U12254 ( .A(n5923), .B(n5919), .Z(n6220) );
  XNOR U12255 ( .A(n5918), .B(n5914), .Z(n6221) );
  XNOR U12256 ( .A(n5913), .B(n5909), .Z(n6222) );
  XNOR U12257 ( .A(n5908), .B(n5904), .Z(n6223) );
  XNOR U12258 ( .A(n5903), .B(n5899), .Z(n6224) );
  XNOR U12259 ( .A(n5898), .B(n5894), .Z(n6225) );
  XNOR U12260 ( .A(n5893), .B(n5889), .Z(n6226) );
  XNOR U12261 ( .A(n5888), .B(n5884), .Z(n6227) );
  XNOR U12262 ( .A(n5883), .B(n5879), .Z(n6228) );
  XNOR U12263 ( .A(n5878), .B(n5874), .Z(n6229) );
  XOR U12264 ( .A(n5873), .B(n5870), .Z(n6230) );
  XOR U12265 ( .A(n6231), .B(n6232), .Z(n5870) );
  XOR U12266 ( .A(n5868), .B(n6233), .Z(n6232) );
  XOR U12267 ( .A(n6234), .B(n6235), .Z(n6233) );
  XOR U12268 ( .A(n6236), .B(n6237), .Z(n6235) );
  NAND U12269 ( .A(a[48]), .B(b[62]), .Z(n6237) );
  AND U12270 ( .A(a[47]), .B(b[63]), .Z(n6236) );
  XOR U12271 ( .A(n6238), .B(n6234), .Z(n6231) );
  XOR U12272 ( .A(n6239), .B(n6240), .Z(n6234) );
  ANDN U12273 ( .B(n6241), .A(n6242), .Z(n6239) );
  AND U12274 ( .A(a[49]), .B(b[61]), .Z(n6238) );
  XOR U12275 ( .A(n6243), .B(n5868), .Z(n5869) );
  XOR U12276 ( .A(n6244), .B(n6245), .Z(n5868) );
  AND U12277 ( .A(n6246), .B(n6247), .Z(n6244) );
  AND U12278 ( .A(a[50]), .B(b[60]), .Z(n6243) );
  XOR U12279 ( .A(n6248), .B(n5873), .Z(n5875) );
  XOR U12280 ( .A(n6249), .B(n6250), .Z(n5873) );
  AND U12281 ( .A(n6251), .B(n6252), .Z(n6249) );
  AND U12282 ( .A(a[51]), .B(b[59]), .Z(n6248) );
  XOR U12283 ( .A(n6253), .B(n5878), .Z(n5880) );
  XOR U12284 ( .A(n6254), .B(n6255), .Z(n5878) );
  AND U12285 ( .A(n6256), .B(n6257), .Z(n6254) );
  AND U12286 ( .A(a[52]), .B(b[58]), .Z(n6253) );
  XOR U12287 ( .A(n6258), .B(n5883), .Z(n5885) );
  XOR U12288 ( .A(n6259), .B(n6260), .Z(n5883) );
  AND U12289 ( .A(n6261), .B(n6262), .Z(n6259) );
  AND U12290 ( .A(a[53]), .B(b[57]), .Z(n6258) );
  XOR U12291 ( .A(n6263), .B(n5888), .Z(n5890) );
  XOR U12292 ( .A(n6264), .B(n6265), .Z(n5888) );
  AND U12293 ( .A(n6266), .B(n6267), .Z(n6264) );
  AND U12294 ( .A(a[54]), .B(b[56]), .Z(n6263) );
  XOR U12295 ( .A(n6268), .B(n5893), .Z(n5895) );
  XOR U12296 ( .A(n6269), .B(n6270), .Z(n5893) );
  AND U12297 ( .A(n6271), .B(n6272), .Z(n6269) );
  AND U12298 ( .A(a[55]), .B(b[55]), .Z(n6268) );
  XOR U12299 ( .A(n6273), .B(n5898), .Z(n5900) );
  XOR U12300 ( .A(n6274), .B(n6275), .Z(n5898) );
  AND U12301 ( .A(n6276), .B(n6277), .Z(n6274) );
  AND U12302 ( .A(b[54]), .B(a[56]), .Z(n6273) );
  XOR U12303 ( .A(n6278), .B(n5903), .Z(n5905) );
  XOR U12304 ( .A(n6279), .B(n6280), .Z(n5903) );
  AND U12305 ( .A(n6281), .B(n6282), .Z(n6279) );
  AND U12306 ( .A(b[53]), .B(a[57]), .Z(n6278) );
  XOR U12307 ( .A(n6283), .B(n5908), .Z(n5910) );
  XOR U12308 ( .A(n6284), .B(n6285), .Z(n5908) );
  AND U12309 ( .A(n6286), .B(n6287), .Z(n6284) );
  AND U12310 ( .A(b[52]), .B(a[58]), .Z(n6283) );
  XOR U12311 ( .A(n6288), .B(n5913), .Z(n5915) );
  XOR U12312 ( .A(n6289), .B(n6290), .Z(n5913) );
  AND U12313 ( .A(n6291), .B(n6292), .Z(n6289) );
  AND U12314 ( .A(b[51]), .B(a[59]), .Z(n6288) );
  XOR U12315 ( .A(n6293), .B(n5918), .Z(n5920) );
  XOR U12316 ( .A(n6294), .B(n6295), .Z(n5918) );
  AND U12317 ( .A(n6296), .B(n6297), .Z(n6294) );
  AND U12318 ( .A(b[50]), .B(a[60]), .Z(n6293) );
  XOR U12319 ( .A(n6298), .B(n5923), .Z(n5925) );
  XOR U12320 ( .A(n6299), .B(n6300), .Z(n5923) );
  AND U12321 ( .A(n6301), .B(n6302), .Z(n6299) );
  AND U12322 ( .A(b[49]), .B(a[61]), .Z(n6298) );
  XOR U12323 ( .A(n6303), .B(n5928), .Z(n5930) );
  XOR U12324 ( .A(n6304), .B(n6305), .Z(n5928) );
  AND U12325 ( .A(n6306), .B(n6307), .Z(n6304) );
  AND U12326 ( .A(b[48]), .B(a[62]), .Z(n6303) );
  XOR U12327 ( .A(n6308), .B(n5933), .Z(n5935) );
  XOR U12328 ( .A(n6309), .B(n6310), .Z(n5933) );
  AND U12329 ( .A(n6311), .B(n6312), .Z(n6309) );
  AND U12330 ( .A(b[47]), .B(a[63]), .Z(n6308) );
  XOR U12331 ( .A(n6313), .B(n5938), .Z(n5940) );
  XOR U12332 ( .A(n6314), .B(n6315), .Z(n5938) );
  AND U12333 ( .A(n6316), .B(n6317), .Z(n6314) );
  AND U12334 ( .A(b[46]), .B(a[64]), .Z(n6313) );
  XOR U12335 ( .A(n6318), .B(n5943), .Z(n5945) );
  XOR U12336 ( .A(n6319), .B(n6320), .Z(n5943) );
  AND U12337 ( .A(n6321), .B(n6322), .Z(n6319) );
  AND U12338 ( .A(b[45]), .B(a[65]), .Z(n6318) );
  XOR U12339 ( .A(n6323), .B(n5948), .Z(n5950) );
  XOR U12340 ( .A(n6324), .B(n6325), .Z(n5948) );
  AND U12341 ( .A(n6326), .B(n6327), .Z(n6324) );
  AND U12342 ( .A(b[44]), .B(a[66]), .Z(n6323) );
  XOR U12343 ( .A(n6328), .B(n5953), .Z(n5955) );
  XOR U12344 ( .A(n6329), .B(n6330), .Z(n5953) );
  AND U12345 ( .A(n6331), .B(n6332), .Z(n6329) );
  AND U12346 ( .A(b[43]), .B(a[67]), .Z(n6328) );
  XOR U12347 ( .A(n6333), .B(n5958), .Z(n5960) );
  XOR U12348 ( .A(n6334), .B(n6335), .Z(n5958) );
  AND U12349 ( .A(n6336), .B(n6337), .Z(n6334) );
  AND U12350 ( .A(b[42]), .B(a[68]), .Z(n6333) );
  XOR U12351 ( .A(n6338), .B(n6339), .Z(n5962) );
  AND U12352 ( .A(n6340), .B(n6341), .Z(n6338) );
  XOR U12353 ( .A(n6342), .B(n5967), .Z(n5969) );
  XOR U12354 ( .A(n6343), .B(n6344), .Z(n5967) );
  AND U12355 ( .A(n6345), .B(n6346), .Z(n6343) );
  AND U12356 ( .A(b[41]), .B(a[69]), .Z(n6342) );
  XOR U12357 ( .A(n6347), .B(n5972), .Z(n5974) );
  XOR U12358 ( .A(n6348), .B(n6349), .Z(n5972) );
  AND U12359 ( .A(n6350), .B(n6351), .Z(n6348) );
  AND U12360 ( .A(b[39]), .B(a[71]), .Z(n6347) );
  XOR U12361 ( .A(n6352), .B(n5977), .Z(n5979) );
  XOR U12362 ( .A(n6353), .B(n6354), .Z(n5977) );
  AND U12363 ( .A(n6355), .B(n6356), .Z(n6353) );
  AND U12364 ( .A(b[38]), .B(a[72]), .Z(n6352) );
  XOR U12365 ( .A(n6357), .B(n5982), .Z(n5984) );
  XOR U12366 ( .A(n6358), .B(n6359), .Z(n5982) );
  AND U12367 ( .A(n6360), .B(n6361), .Z(n6358) );
  AND U12368 ( .A(b[37]), .B(a[73]), .Z(n6357) );
  XOR U12369 ( .A(n6362), .B(n5987), .Z(n5989) );
  XOR U12370 ( .A(n6363), .B(n6364), .Z(n5987) );
  AND U12371 ( .A(n6365), .B(n6366), .Z(n6363) );
  AND U12372 ( .A(b[36]), .B(a[74]), .Z(n6362) );
  XOR U12373 ( .A(n6367), .B(n6368), .Z(n5991) );
  AND U12374 ( .A(n6369), .B(n6370), .Z(n6367) );
  XOR U12375 ( .A(n6371), .B(n5996), .Z(n5998) );
  XOR U12376 ( .A(n6372), .B(n6373), .Z(n5996) );
  AND U12377 ( .A(n6374), .B(n6375), .Z(n6372) );
  AND U12378 ( .A(b[35]), .B(a[75]), .Z(n6371) );
  XOR U12379 ( .A(n6376), .B(n6001), .Z(n6003) );
  XOR U12380 ( .A(n6377), .B(n6378), .Z(n6001) );
  AND U12381 ( .A(n6379), .B(n6380), .Z(n6377) );
  AND U12382 ( .A(b[33]), .B(a[77]), .Z(n6376) );
  XOR U12383 ( .A(n6381), .B(n6006), .Z(n6008) );
  XOR U12384 ( .A(n6382), .B(n6383), .Z(n6006) );
  AND U12385 ( .A(n6384), .B(n6385), .Z(n6382) );
  AND U12386 ( .A(b[32]), .B(a[78]), .Z(n6381) );
  XOR U12387 ( .A(n6386), .B(n6011), .Z(n6013) );
  XOR U12388 ( .A(n6387), .B(n6388), .Z(n6011) );
  AND U12389 ( .A(n6389), .B(n6390), .Z(n6387) );
  AND U12390 ( .A(b[31]), .B(a[79]), .Z(n6386) );
  XOR U12391 ( .A(n6391), .B(n6016), .Z(n6018) );
  XOR U12392 ( .A(n6392), .B(n6393), .Z(n6016) );
  AND U12393 ( .A(n6394), .B(n6395), .Z(n6392) );
  AND U12394 ( .A(b[30]), .B(a[80]), .Z(n6391) );
  XOR U12395 ( .A(n6396), .B(n6397), .Z(n6020) );
  AND U12396 ( .A(n6398), .B(n6399), .Z(n6396) );
  XOR U12397 ( .A(n6400), .B(n6025), .Z(n6027) );
  XOR U12398 ( .A(n6401), .B(n6402), .Z(n6025) );
  AND U12399 ( .A(n6403), .B(n6404), .Z(n6401) );
  AND U12400 ( .A(b[29]), .B(a[81]), .Z(n6400) );
  XOR U12401 ( .A(n6405), .B(n6030), .Z(n6032) );
  XOR U12402 ( .A(n6406), .B(n6407), .Z(n6030) );
  AND U12403 ( .A(n6408), .B(n6409), .Z(n6406) );
  AND U12404 ( .A(b[27]), .B(a[83]), .Z(n6405) );
  XOR U12405 ( .A(n6410), .B(n6035), .Z(n6037) );
  XOR U12406 ( .A(n6411), .B(n6412), .Z(n6035) );
  AND U12407 ( .A(n6413), .B(n6414), .Z(n6411) );
  AND U12408 ( .A(b[26]), .B(a[84]), .Z(n6410) );
  XOR U12409 ( .A(n6415), .B(n6040), .Z(n6042) );
  XOR U12410 ( .A(n6416), .B(n6417), .Z(n6040) );
  AND U12411 ( .A(n6418), .B(n6419), .Z(n6416) );
  AND U12412 ( .A(b[25]), .B(a[85]), .Z(n6415) );
  XOR U12413 ( .A(n6420), .B(n6045), .Z(n6047) );
  XOR U12414 ( .A(n6421), .B(n6422), .Z(n6045) );
  AND U12415 ( .A(n6423), .B(n6424), .Z(n6421) );
  AND U12416 ( .A(b[24]), .B(a[86]), .Z(n6420) );
  XOR U12417 ( .A(n6425), .B(n6426), .Z(n6049) );
  AND U12418 ( .A(n6427), .B(n6428), .Z(n6425) );
  XOR U12419 ( .A(n6429), .B(n6054), .Z(n6056) );
  XOR U12420 ( .A(n6430), .B(n6431), .Z(n6054) );
  AND U12421 ( .A(n6432), .B(n6433), .Z(n6430) );
  AND U12422 ( .A(b[23]), .B(a[87]), .Z(n6429) );
  XOR U12423 ( .A(n6434), .B(n6059), .Z(n6061) );
  XOR U12424 ( .A(n6435), .B(n6436), .Z(n6059) );
  AND U12425 ( .A(n6437), .B(n6438), .Z(n6435) );
  AND U12426 ( .A(b[21]), .B(a[89]), .Z(n6434) );
  XOR U12427 ( .A(n6439), .B(n6064), .Z(n6066) );
  XOR U12428 ( .A(n6440), .B(n6441), .Z(n6064) );
  AND U12429 ( .A(n6442), .B(n6443), .Z(n6440) );
  AND U12430 ( .A(b[20]), .B(a[90]), .Z(n6439) );
  XOR U12431 ( .A(n6444), .B(n6069), .Z(n6071) );
  XOR U12432 ( .A(n6445), .B(n6446), .Z(n6069) );
  AND U12433 ( .A(n6447), .B(n6448), .Z(n6445) );
  AND U12434 ( .A(b[19]), .B(a[91]), .Z(n6444) );
  XOR U12435 ( .A(n6449), .B(n6074), .Z(n6076) );
  XOR U12436 ( .A(n6450), .B(n6451), .Z(n6074) );
  AND U12437 ( .A(n6452), .B(n6453), .Z(n6450) );
  AND U12438 ( .A(b[18]), .B(a[92]), .Z(n6449) );
  XOR U12439 ( .A(n6454), .B(n6455), .Z(n6078) );
  AND U12440 ( .A(n6456), .B(n6457), .Z(n6454) );
  XOR U12441 ( .A(n6458), .B(n6083), .Z(n6085) );
  XOR U12442 ( .A(n6459), .B(n6460), .Z(n6083) );
  AND U12443 ( .A(n6461), .B(n6462), .Z(n6459) );
  AND U12444 ( .A(b[17]), .B(a[93]), .Z(n6458) );
  XOR U12445 ( .A(n6463), .B(n6088), .Z(n6090) );
  XOR U12446 ( .A(n6464), .B(n6465), .Z(n6088) );
  AND U12447 ( .A(n6466), .B(n6467), .Z(n6464) );
  AND U12448 ( .A(b[15]), .B(a[95]), .Z(n6463) );
  XOR U12449 ( .A(n6468), .B(n6093), .Z(n6095) );
  XOR U12450 ( .A(n6469), .B(n6470), .Z(n6093) );
  AND U12451 ( .A(n6471), .B(n6472), .Z(n6469) );
  AND U12452 ( .A(b[14]), .B(a[96]), .Z(n6468) );
  XOR U12453 ( .A(n6473), .B(n6098), .Z(n6100) );
  XOR U12454 ( .A(n6474), .B(n6475), .Z(n6098) );
  AND U12455 ( .A(n6476), .B(n6477), .Z(n6474) );
  AND U12456 ( .A(b[13]), .B(a[97]), .Z(n6473) );
  XOR U12457 ( .A(n6478), .B(n6103), .Z(n6105) );
  XOR U12458 ( .A(n6479), .B(n6480), .Z(n6103) );
  AND U12459 ( .A(n6481), .B(n6482), .Z(n6479) );
  AND U12460 ( .A(b[12]), .B(a[98]), .Z(n6478) );
  XOR U12461 ( .A(n6483), .B(n6484), .Z(n6107) );
  AND U12462 ( .A(n6485), .B(n6486), .Z(n6483) );
  XOR U12463 ( .A(n6487), .B(n6112), .Z(n6114) );
  XOR U12464 ( .A(n6488), .B(n6489), .Z(n6112) );
  AND U12465 ( .A(n6490), .B(n6491), .Z(n6488) );
  AND U12466 ( .A(b[11]), .B(a[99]), .Z(n6487) );
  XOR U12467 ( .A(n6492), .B(n6117), .Z(n6119) );
  XOR U12468 ( .A(n6493), .B(n6494), .Z(n6117) );
  AND U12469 ( .A(n6495), .B(n6496), .Z(n6493) );
  AND U12470 ( .A(b[9]), .B(a[101]), .Z(n6492) );
  XOR U12471 ( .A(n6497), .B(n6122), .Z(n6124) );
  XOR U12472 ( .A(n6498), .B(n6499), .Z(n6122) );
  AND U12473 ( .A(n6500), .B(n6501), .Z(n6498) );
  AND U12474 ( .A(b[8]), .B(a[102]), .Z(n6497) );
  XOR U12475 ( .A(n6502), .B(n6127), .Z(n6129) );
  XOR U12476 ( .A(n6503), .B(n6504), .Z(n6127) );
  AND U12477 ( .A(n6505), .B(n6506), .Z(n6503) );
  AND U12478 ( .A(b[7]), .B(a[103]), .Z(n6502) );
  XOR U12479 ( .A(n6507), .B(n6132), .Z(n6134) );
  XOR U12480 ( .A(n6508), .B(n6509), .Z(n6132) );
  AND U12481 ( .A(n6510), .B(n6511), .Z(n6508) );
  AND U12482 ( .A(b[6]), .B(a[104]), .Z(n6507) );
  XOR U12483 ( .A(n6512), .B(n6513), .Z(n6136) );
  AND U12484 ( .A(n6514), .B(n6515), .Z(n6512) );
  XOR U12485 ( .A(n6516), .B(n6141), .Z(n6143) );
  XOR U12486 ( .A(n6517), .B(n6518), .Z(n6141) );
  AND U12487 ( .A(n6519), .B(n6520), .Z(n6517) );
  AND U12488 ( .A(b[5]), .B(a[105]), .Z(n6516) );
  XNOR U12489 ( .A(n6521), .B(n6522), .Z(n6155) );
  NANDN U12490 ( .A(n6523), .B(n6524), .Z(n6522) );
  XOR U12491 ( .A(n6525), .B(n6146), .Z(n6148) );
  XNOR U12492 ( .A(n6526), .B(n6527), .Z(n6146) );
  ANDN U12493 ( .B(n6528), .A(n6529), .Z(n6526) );
  AND U12494 ( .A(b[3]), .B(a[107]), .Z(n6525) );
  XNOR U12495 ( .A(n6530), .B(n6531), .Z(swire[109]) );
  XOR U12496 ( .A(n6165), .B(n6532), .Z(n6531) );
  NAND U12497 ( .A(a[109]), .B(b[0]), .Z(n6164) );
  XNOR U12498 ( .A(n6523), .B(n6524), .Z(n6165) );
  XOR U12499 ( .A(n6521), .B(n6533), .Z(n6524) );
  NAND U12500 ( .A(b[1]), .B(a[108]), .Z(n6533) );
  XNOR U12501 ( .A(n6529), .B(n6534), .Z(n6523) );
  XOR U12502 ( .A(n6521), .B(n6528), .Z(n6534) );
  XNOR U12503 ( .A(n6535), .B(n6527), .Z(n6528) );
  AND U12504 ( .A(b[2]), .B(a[107]), .Z(n6535) );
  NANDN U12505 ( .A(n6536), .B(n6537), .Z(n6521) );
  XNOR U12506 ( .A(n6527), .B(n6538), .Z(n6529) );
  XNOR U12507 ( .A(n6515), .B(n6514), .Z(n6538) );
  XOR U12508 ( .A(n6539), .B(n6513), .Z(n6514) );
  AND U12509 ( .A(b[3]), .B(a[106]), .Z(n6539) );
  XNOR U12510 ( .A(n6513), .B(n6519), .Z(n6540) );
  XNOR U12511 ( .A(n6518), .B(n6510), .Z(n6541) );
  XNOR U12512 ( .A(n6509), .B(n6505), .Z(n6542) );
  XNOR U12513 ( .A(n6504), .B(n6500), .Z(n6543) );
  XNOR U12514 ( .A(n6499), .B(n6495), .Z(n6544) );
  XNOR U12515 ( .A(n6486), .B(n6485), .Z(n6545) );
  XOR U12516 ( .A(n6546), .B(n6484), .Z(n6485) );
  AND U12517 ( .A(b[9]), .B(a[100]), .Z(n6546) );
  XNOR U12518 ( .A(n6484), .B(n6490), .Z(n6547) );
  XNOR U12519 ( .A(n6489), .B(n6481), .Z(n6548) );
  XNOR U12520 ( .A(n6480), .B(n6476), .Z(n6549) );
  XNOR U12521 ( .A(n6475), .B(n6471), .Z(n6550) );
  XNOR U12522 ( .A(n6470), .B(n6466), .Z(n6551) );
  XNOR U12523 ( .A(n6457), .B(n6456), .Z(n6552) );
  XOR U12524 ( .A(n6553), .B(n6455), .Z(n6456) );
  AND U12525 ( .A(b[15]), .B(a[94]), .Z(n6553) );
  XNOR U12526 ( .A(n6455), .B(n6461), .Z(n6554) );
  XNOR U12527 ( .A(n6460), .B(n6452), .Z(n6555) );
  XNOR U12528 ( .A(n6451), .B(n6447), .Z(n6556) );
  XNOR U12529 ( .A(n6446), .B(n6442), .Z(n6557) );
  XNOR U12530 ( .A(n6441), .B(n6437), .Z(n6558) );
  XNOR U12531 ( .A(n6428), .B(n6427), .Z(n6559) );
  XOR U12532 ( .A(n6560), .B(n6426), .Z(n6427) );
  AND U12533 ( .A(b[21]), .B(a[88]), .Z(n6560) );
  XNOR U12534 ( .A(n6426), .B(n6432), .Z(n6561) );
  XNOR U12535 ( .A(n6431), .B(n6423), .Z(n6562) );
  XNOR U12536 ( .A(n6422), .B(n6418), .Z(n6563) );
  XNOR U12537 ( .A(n6417), .B(n6413), .Z(n6564) );
  XNOR U12538 ( .A(n6412), .B(n6408), .Z(n6565) );
  XNOR U12539 ( .A(n6399), .B(n6398), .Z(n6566) );
  XOR U12540 ( .A(n6567), .B(n6397), .Z(n6398) );
  AND U12541 ( .A(b[27]), .B(a[82]), .Z(n6567) );
  XNOR U12542 ( .A(n6397), .B(n6403), .Z(n6568) );
  XNOR U12543 ( .A(n6402), .B(n6394), .Z(n6569) );
  XNOR U12544 ( .A(n6393), .B(n6389), .Z(n6570) );
  XNOR U12545 ( .A(n6388), .B(n6384), .Z(n6571) );
  XNOR U12546 ( .A(n6383), .B(n6379), .Z(n6572) );
  XNOR U12547 ( .A(n6370), .B(n6369), .Z(n6573) );
  XOR U12548 ( .A(n6574), .B(n6368), .Z(n6369) );
  AND U12549 ( .A(b[33]), .B(a[76]), .Z(n6574) );
  XNOR U12550 ( .A(n6368), .B(n6374), .Z(n6575) );
  XNOR U12551 ( .A(n6373), .B(n6365), .Z(n6576) );
  XNOR U12552 ( .A(n6364), .B(n6360), .Z(n6577) );
  XNOR U12553 ( .A(n6359), .B(n6355), .Z(n6578) );
  XNOR U12554 ( .A(n6354), .B(n6350), .Z(n6579) );
  XNOR U12555 ( .A(n6341), .B(n6340), .Z(n6580) );
  XOR U12556 ( .A(n6581), .B(n6339), .Z(n6340) );
  AND U12557 ( .A(b[39]), .B(a[70]), .Z(n6581) );
  XNOR U12558 ( .A(n6339), .B(n6345), .Z(n6582) );
  XNOR U12559 ( .A(n6344), .B(n6336), .Z(n6583) );
  XNOR U12560 ( .A(n6335), .B(n6331), .Z(n6584) );
  XNOR U12561 ( .A(n6330), .B(n6326), .Z(n6585) );
  XNOR U12562 ( .A(n6325), .B(n6321), .Z(n6586) );
  XNOR U12563 ( .A(n6320), .B(n6316), .Z(n6587) );
  XNOR U12564 ( .A(n6315), .B(n6311), .Z(n6588) );
  XNOR U12565 ( .A(n6310), .B(n6306), .Z(n6589) );
  XNOR U12566 ( .A(n6305), .B(n6301), .Z(n6590) );
  XNOR U12567 ( .A(n6300), .B(n6296), .Z(n6591) );
  XNOR U12568 ( .A(n6295), .B(n6291), .Z(n6592) );
  XNOR U12569 ( .A(n6290), .B(n6286), .Z(n6593) );
  XNOR U12570 ( .A(n6285), .B(n6281), .Z(n6594) );
  XNOR U12571 ( .A(n6280), .B(n6276), .Z(n6595) );
  XNOR U12572 ( .A(n6275), .B(n6271), .Z(n6596) );
  XNOR U12573 ( .A(n6270), .B(n6266), .Z(n6597) );
  XNOR U12574 ( .A(n6265), .B(n6261), .Z(n6598) );
  XNOR U12575 ( .A(n6260), .B(n6256), .Z(n6599) );
  XNOR U12576 ( .A(n6255), .B(n6251), .Z(n6600) );
  XNOR U12577 ( .A(n6250), .B(n6246), .Z(n6601) );
  XOR U12578 ( .A(n6245), .B(n6242), .Z(n6602) );
  XOR U12579 ( .A(n6603), .B(n6604), .Z(n6242) );
  XOR U12580 ( .A(n6240), .B(n6605), .Z(n6604) );
  XOR U12581 ( .A(n6606), .B(n6607), .Z(n6605) );
  XOR U12582 ( .A(n6608), .B(n6609), .Z(n6607) );
  NAND U12583 ( .A(a[47]), .B(b[62]), .Z(n6609) );
  AND U12584 ( .A(a[46]), .B(b[63]), .Z(n6608) );
  XOR U12585 ( .A(n6610), .B(n6606), .Z(n6603) );
  XOR U12586 ( .A(n6611), .B(n6612), .Z(n6606) );
  ANDN U12587 ( .B(n6613), .A(n6614), .Z(n6611) );
  AND U12588 ( .A(a[48]), .B(b[61]), .Z(n6610) );
  XOR U12589 ( .A(n6615), .B(n6240), .Z(n6241) );
  XOR U12590 ( .A(n6616), .B(n6617), .Z(n6240) );
  AND U12591 ( .A(n6618), .B(n6619), .Z(n6616) );
  AND U12592 ( .A(a[49]), .B(b[60]), .Z(n6615) );
  XOR U12593 ( .A(n6620), .B(n6245), .Z(n6247) );
  XOR U12594 ( .A(n6621), .B(n6622), .Z(n6245) );
  AND U12595 ( .A(n6623), .B(n6624), .Z(n6621) );
  AND U12596 ( .A(a[50]), .B(b[59]), .Z(n6620) );
  XOR U12597 ( .A(n6625), .B(n6250), .Z(n6252) );
  XOR U12598 ( .A(n6626), .B(n6627), .Z(n6250) );
  AND U12599 ( .A(n6628), .B(n6629), .Z(n6626) );
  AND U12600 ( .A(a[51]), .B(b[58]), .Z(n6625) );
  XOR U12601 ( .A(n6630), .B(n6255), .Z(n6257) );
  XOR U12602 ( .A(n6631), .B(n6632), .Z(n6255) );
  AND U12603 ( .A(n6633), .B(n6634), .Z(n6631) );
  AND U12604 ( .A(a[52]), .B(b[57]), .Z(n6630) );
  XOR U12605 ( .A(n6635), .B(n6260), .Z(n6262) );
  XOR U12606 ( .A(n6636), .B(n6637), .Z(n6260) );
  AND U12607 ( .A(n6638), .B(n6639), .Z(n6636) );
  AND U12608 ( .A(a[53]), .B(b[56]), .Z(n6635) );
  XOR U12609 ( .A(n6640), .B(n6265), .Z(n6267) );
  XOR U12610 ( .A(n6641), .B(n6642), .Z(n6265) );
  AND U12611 ( .A(n6643), .B(n6644), .Z(n6641) );
  AND U12612 ( .A(a[54]), .B(b[55]), .Z(n6640) );
  XOR U12613 ( .A(n6645), .B(n6270), .Z(n6272) );
  XOR U12614 ( .A(n6646), .B(n6647), .Z(n6270) );
  AND U12615 ( .A(n6648), .B(n6649), .Z(n6646) );
  AND U12616 ( .A(b[54]), .B(a[55]), .Z(n6645) );
  XOR U12617 ( .A(n6650), .B(n6275), .Z(n6277) );
  XOR U12618 ( .A(n6651), .B(n6652), .Z(n6275) );
  AND U12619 ( .A(n6653), .B(n6654), .Z(n6651) );
  AND U12620 ( .A(b[53]), .B(a[56]), .Z(n6650) );
  XOR U12621 ( .A(n6655), .B(n6280), .Z(n6282) );
  XOR U12622 ( .A(n6656), .B(n6657), .Z(n6280) );
  AND U12623 ( .A(n6658), .B(n6659), .Z(n6656) );
  AND U12624 ( .A(b[52]), .B(a[57]), .Z(n6655) );
  XOR U12625 ( .A(n6660), .B(n6285), .Z(n6287) );
  XOR U12626 ( .A(n6661), .B(n6662), .Z(n6285) );
  AND U12627 ( .A(n6663), .B(n6664), .Z(n6661) );
  AND U12628 ( .A(b[51]), .B(a[58]), .Z(n6660) );
  XOR U12629 ( .A(n6665), .B(n6290), .Z(n6292) );
  XOR U12630 ( .A(n6666), .B(n6667), .Z(n6290) );
  AND U12631 ( .A(n6668), .B(n6669), .Z(n6666) );
  AND U12632 ( .A(b[50]), .B(a[59]), .Z(n6665) );
  XOR U12633 ( .A(n6670), .B(n6295), .Z(n6297) );
  XOR U12634 ( .A(n6671), .B(n6672), .Z(n6295) );
  AND U12635 ( .A(n6673), .B(n6674), .Z(n6671) );
  AND U12636 ( .A(b[49]), .B(a[60]), .Z(n6670) );
  XOR U12637 ( .A(n6675), .B(n6300), .Z(n6302) );
  XOR U12638 ( .A(n6676), .B(n6677), .Z(n6300) );
  AND U12639 ( .A(n6678), .B(n6679), .Z(n6676) );
  AND U12640 ( .A(b[48]), .B(a[61]), .Z(n6675) );
  XOR U12641 ( .A(n6680), .B(n6305), .Z(n6307) );
  XOR U12642 ( .A(n6681), .B(n6682), .Z(n6305) );
  AND U12643 ( .A(n6683), .B(n6684), .Z(n6681) );
  AND U12644 ( .A(b[47]), .B(a[62]), .Z(n6680) );
  XOR U12645 ( .A(n6685), .B(n6310), .Z(n6312) );
  XOR U12646 ( .A(n6686), .B(n6687), .Z(n6310) );
  AND U12647 ( .A(n6688), .B(n6689), .Z(n6686) );
  AND U12648 ( .A(b[46]), .B(a[63]), .Z(n6685) );
  XOR U12649 ( .A(n6690), .B(n6315), .Z(n6317) );
  XOR U12650 ( .A(n6691), .B(n6692), .Z(n6315) );
  AND U12651 ( .A(n6693), .B(n6694), .Z(n6691) );
  AND U12652 ( .A(b[45]), .B(a[64]), .Z(n6690) );
  XOR U12653 ( .A(n6695), .B(n6320), .Z(n6322) );
  XOR U12654 ( .A(n6696), .B(n6697), .Z(n6320) );
  AND U12655 ( .A(n6698), .B(n6699), .Z(n6696) );
  AND U12656 ( .A(b[44]), .B(a[65]), .Z(n6695) );
  XOR U12657 ( .A(n6700), .B(n6325), .Z(n6327) );
  XOR U12658 ( .A(n6701), .B(n6702), .Z(n6325) );
  AND U12659 ( .A(n6703), .B(n6704), .Z(n6701) );
  AND U12660 ( .A(b[43]), .B(a[66]), .Z(n6700) );
  XOR U12661 ( .A(n6705), .B(n6330), .Z(n6332) );
  XOR U12662 ( .A(n6706), .B(n6707), .Z(n6330) );
  AND U12663 ( .A(n6708), .B(n6709), .Z(n6706) );
  AND U12664 ( .A(b[42]), .B(a[67]), .Z(n6705) );
  XOR U12665 ( .A(n6710), .B(n6335), .Z(n6337) );
  XOR U12666 ( .A(n6711), .B(n6712), .Z(n6335) );
  AND U12667 ( .A(n6713), .B(n6714), .Z(n6711) );
  AND U12668 ( .A(b[41]), .B(a[68]), .Z(n6710) );
  XOR U12669 ( .A(n6715), .B(n6716), .Z(n6339) );
  AND U12670 ( .A(n6717), .B(n6718), .Z(n6715) );
  XOR U12671 ( .A(n6719), .B(n6344), .Z(n6346) );
  XOR U12672 ( .A(n6720), .B(n6721), .Z(n6344) );
  AND U12673 ( .A(n6722), .B(n6723), .Z(n6720) );
  AND U12674 ( .A(b[40]), .B(a[69]), .Z(n6719) );
  XOR U12675 ( .A(n6724), .B(n6349), .Z(n6351) );
  XOR U12676 ( .A(n6725), .B(n6726), .Z(n6349) );
  AND U12677 ( .A(n6727), .B(n6728), .Z(n6725) );
  AND U12678 ( .A(b[38]), .B(a[71]), .Z(n6724) );
  XOR U12679 ( .A(n6729), .B(n6354), .Z(n6356) );
  XOR U12680 ( .A(n6730), .B(n6731), .Z(n6354) );
  AND U12681 ( .A(n6732), .B(n6733), .Z(n6730) );
  AND U12682 ( .A(b[37]), .B(a[72]), .Z(n6729) );
  XOR U12683 ( .A(n6734), .B(n6359), .Z(n6361) );
  XOR U12684 ( .A(n6735), .B(n6736), .Z(n6359) );
  AND U12685 ( .A(n6737), .B(n6738), .Z(n6735) );
  AND U12686 ( .A(b[36]), .B(a[73]), .Z(n6734) );
  XOR U12687 ( .A(n6739), .B(n6364), .Z(n6366) );
  XOR U12688 ( .A(n6740), .B(n6741), .Z(n6364) );
  AND U12689 ( .A(n6742), .B(n6743), .Z(n6740) );
  AND U12690 ( .A(b[35]), .B(a[74]), .Z(n6739) );
  XOR U12691 ( .A(n6744), .B(n6745), .Z(n6368) );
  AND U12692 ( .A(n6746), .B(n6747), .Z(n6744) );
  XOR U12693 ( .A(n6748), .B(n6373), .Z(n6375) );
  XOR U12694 ( .A(n6749), .B(n6750), .Z(n6373) );
  AND U12695 ( .A(n6751), .B(n6752), .Z(n6749) );
  AND U12696 ( .A(b[34]), .B(a[75]), .Z(n6748) );
  XOR U12697 ( .A(n6753), .B(n6378), .Z(n6380) );
  XOR U12698 ( .A(n6754), .B(n6755), .Z(n6378) );
  AND U12699 ( .A(n6756), .B(n6757), .Z(n6754) );
  AND U12700 ( .A(b[32]), .B(a[77]), .Z(n6753) );
  XOR U12701 ( .A(n6758), .B(n6383), .Z(n6385) );
  XOR U12702 ( .A(n6759), .B(n6760), .Z(n6383) );
  AND U12703 ( .A(n6761), .B(n6762), .Z(n6759) );
  AND U12704 ( .A(b[31]), .B(a[78]), .Z(n6758) );
  XOR U12705 ( .A(n6763), .B(n6388), .Z(n6390) );
  XOR U12706 ( .A(n6764), .B(n6765), .Z(n6388) );
  AND U12707 ( .A(n6766), .B(n6767), .Z(n6764) );
  AND U12708 ( .A(b[30]), .B(a[79]), .Z(n6763) );
  XOR U12709 ( .A(n6768), .B(n6393), .Z(n6395) );
  XOR U12710 ( .A(n6769), .B(n6770), .Z(n6393) );
  AND U12711 ( .A(n6771), .B(n6772), .Z(n6769) );
  AND U12712 ( .A(b[29]), .B(a[80]), .Z(n6768) );
  XOR U12713 ( .A(n6773), .B(n6774), .Z(n6397) );
  AND U12714 ( .A(n6775), .B(n6776), .Z(n6773) );
  XOR U12715 ( .A(n6777), .B(n6402), .Z(n6404) );
  XOR U12716 ( .A(n6778), .B(n6779), .Z(n6402) );
  AND U12717 ( .A(n6780), .B(n6781), .Z(n6778) );
  AND U12718 ( .A(b[28]), .B(a[81]), .Z(n6777) );
  XOR U12719 ( .A(n6782), .B(n6407), .Z(n6409) );
  XOR U12720 ( .A(n6783), .B(n6784), .Z(n6407) );
  AND U12721 ( .A(n6785), .B(n6786), .Z(n6783) );
  AND U12722 ( .A(b[26]), .B(a[83]), .Z(n6782) );
  XOR U12723 ( .A(n6787), .B(n6412), .Z(n6414) );
  XOR U12724 ( .A(n6788), .B(n6789), .Z(n6412) );
  AND U12725 ( .A(n6790), .B(n6791), .Z(n6788) );
  AND U12726 ( .A(b[25]), .B(a[84]), .Z(n6787) );
  XOR U12727 ( .A(n6792), .B(n6417), .Z(n6419) );
  XOR U12728 ( .A(n6793), .B(n6794), .Z(n6417) );
  AND U12729 ( .A(n6795), .B(n6796), .Z(n6793) );
  AND U12730 ( .A(b[24]), .B(a[85]), .Z(n6792) );
  XOR U12731 ( .A(n6797), .B(n6422), .Z(n6424) );
  XOR U12732 ( .A(n6798), .B(n6799), .Z(n6422) );
  AND U12733 ( .A(n6800), .B(n6801), .Z(n6798) );
  AND U12734 ( .A(b[23]), .B(a[86]), .Z(n6797) );
  XOR U12735 ( .A(n6802), .B(n6803), .Z(n6426) );
  AND U12736 ( .A(n6804), .B(n6805), .Z(n6802) );
  XOR U12737 ( .A(n6806), .B(n6431), .Z(n6433) );
  XOR U12738 ( .A(n6807), .B(n6808), .Z(n6431) );
  AND U12739 ( .A(n6809), .B(n6810), .Z(n6807) );
  AND U12740 ( .A(b[22]), .B(a[87]), .Z(n6806) );
  XOR U12741 ( .A(n6811), .B(n6436), .Z(n6438) );
  XOR U12742 ( .A(n6812), .B(n6813), .Z(n6436) );
  AND U12743 ( .A(n6814), .B(n6815), .Z(n6812) );
  AND U12744 ( .A(b[20]), .B(a[89]), .Z(n6811) );
  XOR U12745 ( .A(n6816), .B(n6441), .Z(n6443) );
  XOR U12746 ( .A(n6817), .B(n6818), .Z(n6441) );
  AND U12747 ( .A(n6819), .B(n6820), .Z(n6817) );
  AND U12748 ( .A(b[19]), .B(a[90]), .Z(n6816) );
  XOR U12749 ( .A(n6821), .B(n6446), .Z(n6448) );
  XOR U12750 ( .A(n6822), .B(n6823), .Z(n6446) );
  AND U12751 ( .A(n6824), .B(n6825), .Z(n6822) );
  AND U12752 ( .A(b[18]), .B(a[91]), .Z(n6821) );
  XOR U12753 ( .A(n6826), .B(n6451), .Z(n6453) );
  XOR U12754 ( .A(n6827), .B(n6828), .Z(n6451) );
  AND U12755 ( .A(n6829), .B(n6830), .Z(n6827) );
  AND U12756 ( .A(b[17]), .B(a[92]), .Z(n6826) );
  XOR U12757 ( .A(n6831), .B(n6832), .Z(n6455) );
  AND U12758 ( .A(n6833), .B(n6834), .Z(n6831) );
  XOR U12759 ( .A(n6835), .B(n6460), .Z(n6462) );
  XOR U12760 ( .A(n6836), .B(n6837), .Z(n6460) );
  AND U12761 ( .A(n6838), .B(n6839), .Z(n6836) );
  AND U12762 ( .A(b[16]), .B(a[93]), .Z(n6835) );
  XOR U12763 ( .A(n6840), .B(n6465), .Z(n6467) );
  XOR U12764 ( .A(n6841), .B(n6842), .Z(n6465) );
  AND U12765 ( .A(n6843), .B(n6844), .Z(n6841) );
  AND U12766 ( .A(b[14]), .B(a[95]), .Z(n6840) );
  XOR U12767 ( .A(n6845), .B(n6470), .Z(n6472) );
  XOR U12768 ( .A(n6846), .B(n6847), .Z(n6470) );
  AND U12769 ( .A(n6848), .B(n6849), .Z(n6846) );
  AND U12770 ( .A(b[13]), .B(a[96]), .Z(n6845) );
  XOR U12771 ( .A(n6850), .B(n6475), .Z(n6477) );
  XOR U12772 ( .A(n6851), .B(n6852), .Z(n6475) );
  AND U12773 ( .A(n6853), .B(n6854), .Z(n6851) );
  AND U12774 ( .A(b[12]), .B(a[97]), .Z(n6850) );
  XOR U12775 ( .A(n6855), .B(n6480), .Z(n6482) );
  XOR U12776 ( .A(n6856), .B(n6857), .Z(n6480) );
  AND U12777 ( .A(n6858), .B(n6859), .Z(n6856) );
  AND U12778 ( .A(b[11]), .B(a[98]), .Z(n6855) );
  XOR U12779 ( .A(n6860), .B(n6861), .Z(n6484) );
  AND U12780 ( .A(n6862), .B(n6863), .Z(n6860) );
  XOR U12781 ( .A(n6864), .B(n6489), .Z(n6491) );
  XOR U12782 ( .A(n6865), .B(n6866), .Z(n6489) );
  AND U12783 ( .A(n6867), .B(n6868), .Z(n6865) );
  AND U12784 ( .A(b[10]), .B(a[99]), .Z(n6864) );
  XOR U12785 ( .A(n6869), .B(n6494), .Z(n6496) );
  XOR U12786 ( .A(n6870), .B(n6871), .Z(n6494) );
  AND U12787 ( .A(n6872), .B(n6873), .Z(n6870) );
  AND U12788 ( .A(b[8]), .B(a[101]), .Z(n6869) );
  XOR U12789 ( .A(n6874), .B(n6499), .Z(n6501) );
  XOR U12790 ( .A(n6875), .B(n6876), .Z(n6499) );
  AND U12791 ( .A(n6877), .B(n6878), .Z(n6875) );
  AND U12792 ( .A(b[7]), .B(a[102]), .Z(n6874) );
  XOR U12793 ( .A(n6879), .B(n6504), .Z(n6506) );
  XOR U12794 ( .A(n6880), .B(n6881), .Z(n6504) );
  AND U12795 ( .A(n6882), .B(n6883), .Z(n6880) );
  AND U12796 ( .A(b[6]), .B(a[103]), .Z(n6879) );
  XOR U12797 ( .A(n6884), .B(n6509), .Z(n6511) );
  XOR U12798 ( .A(n6885), .B(n6886), .Z(n6509) );
  AND U12799 ( .A(n6887), .B(n6888), .Z(n6885) );
  AND U12800 ( .A(b[5]), .B(a[104]), .Z(n6884) );
  XOR U12801 ( .A(n6889), .B(n6890), .Z(n6513) );
  AND U12802 ( .A(n6891), .B(n6892), .Z(n6889) );
  XOR U12803 ( .A(n6893), .B(n6518), .Z(n6520) );
  XOR U12804 ( .A(n6894), .B(n6895), .Z(n6518) );
  AND U12805 ( .A(n6896), .B(n6897), .Z(n6894) );
  AND U12806 ( .A(b[4]), .B(a[105]), .Z(n6893) );
  XNOR U12807 ( .A(n6898), .B(n6899), .Z(n6527) );
  NAND U12808 ( .A(n6900), .B(n6901), .Z(n6899) );
  XNOR U12809 ( .A(n6902), .B(n6903), .Z(swire[108]) );
  XOR U12810 ( .A(n6537), .B(n6904), .Z(n6903) );
  NAND U12811 ( .A(a[108]), .B(b[0]), .Z(n6536) );
  XOR U12812 ( .A(n6900), .B(n6901), .Z(n6537) );
  XOR U12813 ( .A(n6898), .B(n6905), .Z(n6901) );
  NAND U12814 ( .A(b[1]), .B(a[107]), .Z(n6905) );
  XOR U12815 ( .A(n6898), .B(n6891), .Z(n6906) );
  XNOR U12816 ( .A(n6890), .B(n6896), .Z(n6907) );
  XNOR U12817 ( .A(n6895), .B(n6887), .Z(n6908) );
  XNOR U12818 ( .A(n6886), .B(n6882), .Z(n6909) );
  XNOR U12819 ( .A(n6881), .B(n6877), .Z(n6910) );
  XNOR U12820 ( .A(n6876), .B(n6872), .Z(n6911) );
  XNOR U12821 ( .A(n6863), .B(n6862), .Z(n6912) );
  XOR U12822 ( .A(n6913), .B(n6861), .Z(n6862) );
  AND U12823 ( .A(b[8]), .B(a[100]), .Z(n6913) );
  XNOR U12824 ( .A(n6861), .B(n6867), .Z(n6914) );
  XNOR U12825 ( .A(n6866), .B(n6858), .Z(n6915) );
  XNOR U12826 ( .A(n6857), .B(n6853), .Z(n6916) );
  XNOR U12827 ( .A(n6852), .B(n6848), .Z(n6917) );
  XNOR U12828 ( .A(n6847), .B(n6843), .Z(n6918) );
  XNOR U12829 ( .A(n6834), .B(n6833), .Z(n6919) );
  XOR U12830 ( .A(n6920), .B(n6832), .Z(n6833) );
  AND U12831 ( .A(b[14]), .B(a[94]), .Z(n6920) );
  XNOR U12832 ( .A(n6832), .B(n6838), .Z(n6921) );
  XNOR U12833 ( .A(n6837), .B(n6829), .Z(n6922) );
  XNOR U12834 ( .A(n6828), .B(n6824), .Z(n6923) );
  XNOR U12835 ( .A(n6823), .B(n6819), .Z(n6924) );
  XNOR U12836 ( .A(n6818), .B(n6814), .Z(n6925) );
  XNOR U12837 ( .A(n6805), .B(n6804), .Z(n6926) );
  XOR U12838 ( .A(n6927), .B(n6803), .Z(n6804) );
  AND U12839 ( .A(b[20]), .B(a[88]), .Z(n6927) );
  XNOR U12840 ( .A(n6803), .B(n6809), .Z(n6928) );
  XNOR U12841 ( .A(n6808), .B(n6800), .Z(n6929) );
  XNOR U12842 ( .A(n6799), .B(n6795), .Z(n6930) );
  XNOR U12843 ( .A(n6794), .B(n6790), .Z(n6931) );
  XNOR U12844 ( .A(n6789), .B(n6785), .Z(n6932) );
  XNOR U12845 ( .A(n6776), .B(n6775), .Z(n6933) );
  XOR U12846 ( .A(n6934), .B(n6774), .Z(n6775) );
  AND U12847 ( .A(b[26]), .B(a[82]), .Z(n6934) );
  XNOR U12848 ( .A(n6774), .B(n6780), .Z(n6935) );
  XNOR U12849 ( .A(n6779), .B(n6771), .Z(n6936) );
  XNOR U12850 ( .A(n6770), .B(n6766), .Z(n6937) );
  XNOR U12851 ( .A(n6765), .B(n6761), .Z(n6938) );
  XNOR U12852 ( .A(n6760), .B(n6756), .Z(n6939) );
  XNOR U12853 ( .A(n6747), .B(n6746), .Z(n6940) );
  XOR U12854 ( .A(n6941), .B(n6745), .Z(n6746) );
  AND U12855 ( .A(b[32]), .B(a[76]), .Z(n6941) );
  XNOR U12856 ( .A(n6745), .B(n6751), .Z(n6942) );
  XNOR U12857 ( .A(n6750), .B(n6742), .Z(n6943) );
  XNOR U12858 ( .A(n6741), .B(n6737), .Z(n6944) );
  XNOR U12859 ( .A(n6736), .B(n6732), .Z(n6945) );
  XNOR U12860 ( .A(n6731), .B(n6727), .Z(n6946) );
  XNOR U12861 ( .A(n6718), .B(n6717), .Z(n6947) );
  XOR U12862 ( .A(n6948), .B(n6716), .Z(n6717) );
  AND U12863 ( .A(b[38]), .B(a[70]), .Z(n6948) );
  XNOR U12864 ( .A(n6716), .B(n6722), .Z(n6949) );
  XNOR U12865 ( .A(n6721), .B(n6713), .Z(n6950) );
  XNOR U12866 ( .A(n6712), .B(n6708), .Z(n6951) );
  XNOR U12867 ( .A(n6707), .B(n6703), .Z(n6952) );
  XNOR U12868 ( .A(n6702), .B(n6698), .Z(n6953) );
  XNOR U12869 ( .A(n6697), .B(n6693), .Z(n6954) );
  XNOR U12870 ( .A(n6692), .B(n6688), .Z(n6955) );
  XNOR U12871 ( .A(n6687), .B(n6683), .Z(n6956) );
  XNOR U12872 ( .A(n6682), .B(n6678), .Z(n6957) );
  XNOR U12873 ( .A(n6677), .B(n6673), .Z(n6958) );
  XNOR U12874 ( .A(n6672), .B(n6668), .Z(n6959) );
  XNOR U12875 ( .A(n6667), .B(n6663), .Z(n6960) );
  XNOR U12876 ( .A(n6662), .B(n6658), .Z(n6961) );
  XNOR U12877 ( .A(n6657), .B(n6653), .Z(n6962) );
  XNOR U12878 ( .A(n6652), .B(n6648), .Z(n6963) );
  XNOR U12879 ( .A(n6647), .B(n6643), .Z(n6964) );
  XNOR U12880 ( .A(n6642), .B(n6638), .Z(n6965) );
  XNOR U12881 ( .A(n6637), .B(n6633), .Z(n6966) );
  XNOR U12882 ( .A(n6632), .B(n6628), .Z(n6967) );
  XNOR U12883 ( .A(n6627), .B(n6623), .Z(n6968) );
  XNOR U12884 ( .A(n6622), .B(n6618), .Z(n6969) );
  XOR U12885 ( .A(n6617), .B(n6614), .Z(n6970) );
  XOR U12886 ( .A(n6971), .B(n6972), .Z(n6614) );
  XOR U12887 ( .A(n6612), .B(n6973), .Z(n6972) );
  XOR U12888 ( .A(n6974), .B(n6975), .Z(n6973) );
  XOR U12889 ( .A(n6976), .B(n6977), .Z(n6975) );
  NAND U12890 ( .A(a[46]), .B(b[62]), .Z(n6977) );
  AND U12891 ( .A(a[45]), .B(b[63]), .Z(n6976) );
  XOR U12892 ( .A(n6978), .B(n6974), .Z(n6971) );
  XOR U12893 ( .A(n6979), .B(n6980), .Z(n6974) );
  ANDN U12894 ( .B(n6981), .A(n6982), .Z(n6979) );
  AND U12895 ( .A(a[47]), .B(b[61]), .Z(n6978) );
  XOR U12896 ( .A(n6983), .B(n6612), .Z(n6613) );
  XOR U12897 ( .A(n6984), .B(n6985), .Z(n6612) );
  AND U12898 ( .A(n6986), .B(n6987), .Z(n6984) );
  AND U12899 ( .A(a[48]), .B(b[60]), .Z(n6983) );
  XOR U12900 ( .A(n6988), .B(n6617), .Z(n6619) );
  XOR U12901 ( .A(n6989), .B(n6990), .Z(n6617) );
  AND U12902 ( .A(n6991), .B(n6992), .Z(n6989) );
  AND U12903 ( .A(a[49]), .B(b[59]), .Z(n6988) );
  XOR U12904 ( .A(n6993), .B(n6622), .Z(n6624) );
  XOR U12905 ( .A(n6994), .B(n6995), .Z(n6622) );
  AND U12906 ( .A(n6996), .B(n6997), .Z(n6994) );
  AND U12907 ( .A(a[50]), .B(b[58]), .Z(n6993) );
  XOR U12908 ( .A(n6998), .B(n6627), .Z(n6629) );
  XOR U12909 ( .A(n6999), .B(n7000), .Z(n6627) );
  AND U12910 ( .A(n7001), .B(n7002), .Z(n6999) );
  AND U12911 ( .A(a[51]), .B(b[57]), .Z(n6998) );
  XOR U12912 ( .A(n7003), .B(n6632), .Z(n6634) );
  XOR U12913 ( .A(n7004), .B(n7005), .Z(n6632) );
  AND U12914 ( .A(n7006), .B(n7007), .Z(n7004) );
  AND U12915 ( .A(a[52]), .B(b[56]), .Z(n7003) );
  XOR U12916 ( .A(n7008), .B(n6637), .Z(n6639) );
  XOR U12917 ( .A(n7009), .B(n7010), .Z(n6637) );
  AND U12918 ( .A(n7011), .B(n7012), .Z(n7009) );
  AND U12919 ( .A(a[53]), .B(b[55]), .Z(n7008) );
  XOR U12920 ( .A(n7013), .B(n6642), .Z(n6644) );
  XOR U12921 ( .A(n7014), .B(n7015), .Z(n6642) );
  AND U12922 ( .A(n7016), .B(n7017), .Z(n7014) );
  AND U12923 ( .A(a[54]), .B(b[54]), .Z(n7013) );
  XOR U12924 ( .A(n7018), .B(n6647), .Z(n6649) );
  XOR U12925 ( .A(n7019), .B(n7020), .Z(n6647) );
  AND U12926 ( .A(n7021), .B(n7022), .Z(n7019) );
  AND U12927 ( .A(b[53]), .B(a[55]), .Z(n7018) );
  XOR U12928 ( .A(n7023), .B(n6652), .Z(n6654) );
  XOR U12929 ( .A(n7024), .B(n7025), .Z(n6652) );
  AND U12930 ( .A(n7026), .B(n7027), .Z(n7024) );
  AND U12931 ( .A(b[52]), .B(a[56]), .Z(n7023) );
  XOR U12932 ( .A(n7028), .B(n6657), .Z(n6659) );
  XOR U12933 ( .A(n7029), .B(n7030), .Z(n6657) );
  AND U12934 ( .A(n7031), .B(n7032), .Z(n7029) );
  AND U12935 ( .A(b[51]), .B(a[57]), .Z(n7028) );
  XOR U12936 ( .A(n7033), .B(n6662), .Z(n6664) );
  XOR U12937 ( .A(n7034), .B(n7035), .Z(n6662) );
  AND U12938 ( .A(n7036), .B(n7037), .Z(n7034) );
  AND U12939 ( .A(b[50]), .B(a[58]), .Z(n7033) );
  XOR U12940 ( .A(n7038), .B(n6667), .Z(n6669) );
  XOR U12941 ( .A(n7039), .B(n7040), .Z(n6667) );
  AND U12942 ( .A(n7041), .B(n7042), .Z(n7039) );
  AND U12943 ( .A(b[49]), .B(a[59]), .Z(n7038) );
  XOR U12944 ( .A(n7043), .B(n6672), .Z(n6674) );
  XOR U12945 ( .A(n7044), .B(n7045), .Z(n6672) );
  AND U12946 ( .A(n7046), .B(n7047), .Z(n7044) );
  AND U12947 ( .A(b[48]), .B(a[60]), .Z(n7043) );
  XOR U12948 ( .A(n7048), .B(n6677), .Z(n6679) );
  XOR U12949 ( .A(n7049), .B(n7050), .Z(n6677) );
  AND U12950 ( .A(n7051), .B(n7052), .Z(n7049) );
  AND U12951 ( .A(b[47]), .B(a[61]), .Z(n7048) );
  XOR U12952 ( .A(n7053), .B(n6682), .Z(n6684) );
  XOR U12953 ( .A(n7054), .B(n7055), .Z(n6682) );
  AND U12954 ( .A(n7056), .B(n7057), .Z(n7054) );
  AND U12955 ( .A(b[46]), .B(a[62]), .Z(n7053) );
  XOR U12956 ( .A(n7058), .B(n6687), .Z(n6689) );
  XOR U12957 ( .A(n7059), .B(n7060), .Z(n6687) );
  AND U12958 ( .A(n7061), .B(n7062), .Z(n7059) );
  AND U12959 ( .A(b[45]), .B(a[63]), .Z(n7058) );
  XOR U12960 ( .A(n7063), .B(n6692), .Z(n6694) );
  XOR U12961 ( .A(n7064), .B(n7065), .Z(n6692) );
  AND U12962 ( .A(n7066), .B(n7067), .Z(n7064) );
  AND U12963 ( .A(b[44]), .B(a[64]), .Z(n7063) );
  XOR U12964 ( .A(n7068), .B(n6697), .Z(n6699) );
  XOR U12965 ( .A(n7069), .B(n7070), .Z(n6697) );
  AND U12966 ( .A(n7071), .B(n7072), .Z(n7069) );
  AND U12967 ( .A(b[43]), .B(a[65]), .Z(n7068) );
  XOR U12968 ( .A(n7073), .B(n6702), .Z(n6704) );
  XOR U12969 ( .A(n7074), .B(n7075), .Z(n6702) );
  AND U12970 ( .A(n7076), .B(n7077), .Z(n7074) );
  AND U12971 ( .A(b[42]), .B(a[66]), .Z(n7073) );
  XOR U12972 ( .A(n7078), .B(n6707), .Z(n6709) );
  XOR U12973 ( .A(n7079), .B(n7080), .Z(n6707) );
  AND U12974 ( .A(n7081), .B(n7082), .Z(n7079) );
  AND U12975 ( .A(b[41]), .B(a[67]), .Z(n7078) );
  XOR U12976 ( .A(n7083), .B(n6712), .Z(n6714) );
  XOR U12977 ( .A(n7084), .B(n7085), .Z(n6712) );
  AND U12978 ( .A(n7086), .B(n7087), .Z(n7084) );
  AND U12979 ( .A(b[40]), .B(a[68]), .Z(n7083) );
  XOR U12980 ( .A(n7088), .B(n7089), .Z(n6716) );
  AND U12981 ( .A(n7090), .B(n7091), .Z(n7088) );
  XOR U12982 ( .A(n7092), .B(n6721), .Z(n6723) );
  XOR U12983 ( .A(n7093), .B(n7094), .Z(n6721) );
  AND U12984 ( .A(n7095), .B(n7096), .Z(n7093) );
  AND U12985 ( .A(b[39]), .B(a[69]), .Z(n7092) );
  XOR U12986 ( .A(n7097), .B(n6726), .Z(n6728) );
  XOR U12987 ( .A(n7098), .B(n7099), .Z(n6726) );
  AND U12988 ( .A(n7100), .B(n7101), .Z(n7098) );
  AND U12989 ( .A(b[37]), .B(a[71]), .Z(n7097) );
  XOR U12990 ( .A(n7102), .B(n6731), .Z(n6733) );
  XOR U12991 ( .A(n7103), .B(n7104), .Z(n6731) );
  AND U12992 ( .A(n7105), .B(n7106), .Z(n7103) );
  AND U12993 ( .A(b[36]), .B(a[72]), .Z(n7102) );
  XOR U12994 ( .A(n7107), .B(n6736), .Z(n6738) );
  XOR U12995 ( .A(n7108), .B(n7109), .Z(n6736) );
  AND U12996 ( .A(n7110), .B(n7111), .Z(n7108) );
  AND U12997 ( .A(b[35]), .B(a[73]), .Z(n7107) );
  XOR U12998 ( .A(n7112), .B(n6741), .Z(n6743) );
  XOR U12999 ( .A(n7113), .B(n7114), .Z(n6741) );
  AND U13000 ( .A(n7115), .B(n7116), .Z(n7113) );
  AND U13001 ( .A(b[34]), .B(a[74]), .Z(n7112) );
  XOR U13002 ( .A(n7117), .B(n7118), .Z(n6745) );
  AND U13003 ( .A(n7119), .B(n7120), .Z(n7117) );
  XOR U13004 ( .A(n7121), .B(n6750), .Z(n6752) );
  XOR U13005 ( .A(n7122), .B(n7123), .Z(n6750) );
  AND U13006 ( .A(n7124), .B(n7125), .Z(n7122) );
  AND U13007 ( .A(b[33]), .B(a[75]), .Z(n7121) );
  XOR U13008 ( .A(n7126), .B(n6755), .Z(n6757) );
  XOR U13009 ( .A(n7127), .B(n7128), .Z(n6755) );
  AND U13010 ( .A(n7129), .B(n7130), .Z(n7127) );
  AND U13011 ( .A(b[31]), .B(a[77]), .Z(n7126) );
  XOR U13012 ( .A(n7131), .B(n6760), .Z(n6762) );
  XOR U13013 ( .A(n7132), .B(n7133), .Z(n6760) );
  AND U13014 ( .A(n7134), .B(n7135), .Z(n7132) );
  AND U13015 ( .A(b[30]), .B(a[78]), .Z(n7131) );
  XOR U13016 ( .A(n7136), .B(n6765), .Z(n6767) );
  XOR U13017 ( .A(n7137), .B(n7138), .Z(n6765) );
  AND U13018 ( .A(n7139), .B(n7140), .Z(n7137) );
  AND U13019 ( .A(b[29]), .B(a[79]), .Z(n7136) );
  XOR U13020 ( .A(n7141), .B(n6770), .Z(n6772) );
  XOR U13021 ( .A(n7142), .B(n7143), .Z(n6770) );
  AND U13022 ( .A(n7144), .B(n7145), .Z(n7142) );
  AND U13023 ( .A(b[28]), .B(a[80]), .Z(n7141) );
  XOR U13024 ( .A(n7146), .B(n7147), .Z(n6774) );
  AND U13025 ( .A(n7148), .B(n7149), .Z(n7146) );
  XOR U13026 ( .A(n7150), .B(n6779), .Z(n6781) );
  XOR U13027 ( .A(n7151), .B(n7152), .Z(n6779) );
  AND U13028 ( .A(n7153), .B(n7154), .Z(n7151) );
  AND U13029 ( .A(b[27]), .B(a[81]), .Z(n7150) );
  XOR U13030 ( .A(n7155), .B(n6784), .Z(n6786) );
  XOR U13031 ( .A(n7156), .B(n7157), .Z(n6784) );
  AND U13032 ( .A(n7158), .B(n7159), .Z(n7156) );
  AND U13033 ( .A(b[25]), .B(a[83]), .Z(n7155) );
  XOR U13034 ( .A(n7160), .B(n6789), .Z(n6791) );
  XOR U13035 ( .A(n7161), .B(n7162), .Z(n6789) );
  AND U13036 ( .A(n7163), .B(n7164), .Z(n7161) );
  AND U13037 ( .A(b[24]), .B(a[84]), .Z(n7160) );
  XOR U13038 ( .A(n7165), .B(n6794), .Z(n6796) );
  XOR U13039 ( .A(n7166), .B(n7167), .Z(n6794) );
  AND U13040 ( .A(n7168), .B(n7169), .Z(n7166) );
  AND U13041 ( .A(b[23]), .B(a[85]), .Z(n7165) );
  XOR U13042 ( .A(n7170), .B(n6799), .Z(n6801) );
  XOR U13043 ( .A(n7171), .B(n7172), .Z(n6799) );
  AND U13044 ( .A(n7173), .B(n7174), .Z(n7171) );
  AND U13045 ( .A(b[22]), .B(a[86]), .Z(n7170) );
  XOR U13046 ( .A(n7175), .B(n7176), .Z(n6803) );
  AND U13047 ( .A(n7177), .B(n7178), .Z(n7175) );
  XOR U13048 ( .A(n7179), .B(n6808), .Z(n6810) );
  XOR U13049 ( .A(n7180), .B(n7181), .Z(n6808) );
  AND U13050 ( .A(n7182), .B(n7183), .Z(n7180) );
  AND U13051 ( .A(b[21]), .B(a[87]), .Z(n7179) );
  XOR U13052 ( .A(n7184), .B(n6813), .Z(n6815) );
  XOR U13053 ( .A(n7185), .B(n7186), .Z(n6813) );
  AND U13054 ( .A(n7187), .B(n7188), .Z(n7185) );
  AND U13055 ( .A(b[19]), .B(a[89]), .Z(n7184) );
  XOR U13056 ( .A(n7189), .B(n6818), .Z(n6820) );
  XOR U13057 ( .A(n7190), .B(n7191), .Z(n6818) );
  AND U13058 ( .A(n7192), .B(n7193), .Z(n7190) );
  AND U13059 ( .A(b[18]), .B(a[90]), .Z(n7189) );
  XOR U13060 ( .A(n7194), .B(n6823), .Z(n6825) );
  XOR U13061 ( .A(n7195), .B(n7196), .Z(n6823) );
  AND U13062 ( .A(n7197), .B(n7198), .Z(n7195) );
  AND U13063 ( .A(b[17]), .B(a[91]), .Z(n7194) );
  XOR U13064 ( .A(n7199), .B(n6828), .Z(n6830) );
  XOR U13065 ( .A(n7200), .B(n7201), .Z(n6828) );
  AND U13066 ( .A(n7202), .B(n7203), .Z(n7200) );
  AND U13067 ( .A(b[16]), .B(a[92]), .Z(n7199) );
  XOR U13068 ( .A(n7204), .B(n7205), .Z(n6832) );
  AND U13069 ( .A(n7206), .B(n7207), .Z(n7204) );
  XOR U13070 ( .A(n7208), .B(n6837), .Z(n6839) );
  XOR U13071 ( .A(n7209), .B(n7210), .Z(n6837) );
  AND U13072 ( .A(n7211), .B(n7212), .Z(n7209) );
  AND U13073 ( .A(b[15]), .B(a[93]), .Z(n7208) );
  XOR U13074 ( .A(n7213), .B(n6842), .Z(n6844) );
  XOR U13075 ( .A(n7214), .B(n7215), .Z(n6842) );
  AND U13076 ( .A(n7216), .B(n7217), .Z(n7214) );
  AND U13077 ( .A(b[13]), .B(a[95]), .Z(n7213) );
  XOR U13078 ( .A(n7218), .B(n6847), .Z(n6849) );
  XOR U13079 ( .A(n7219), .B(n7220), .Z(n6847) );
  AND U13080 ( .A(n7221), .B(n7222), .Z(n7219) );
  AND U13081 ( .A(b[12]), .B(a[96]), .Z(n7218) );
  XOR U13082 ( .A(n7223), .B(n6852), .Z(n6854) );
  XOR U13083 ( .A(n7224), .B(n7225), .Z(n6852) );
  AND U13084 ( .A(n7226), .B(n7227), .Z(n7224) );
  AND U13085 ( .A(b[11]), .B(a[97]), .Z(n7223) );
  XOR U13086 ( .A(n7228), .B(n6857), .Z(n6859) );
  XOR U13087 ( .A(n7229), .B(n7230), .Z(n6857) );
  AND U13088 ( .A(n7231), .B(n7232), .Z(n7229) );
  AND U13089 ( .A(b[10]), .B(a[98]), .Z(n7228) );
  XOR U13090 ( .A(n7233), .B(n7234), .Z(n6861) );
  AND U13091 ( .A(n7235), .B(n7236), .Z(n7233) );
  XOR U13092 ( .A(n7237), .B(n6866), .Z(n6868) );
  XOR U13093 ( .A(n7238), .B(n7239), .Z(n6866) );
  AND U13094 ( .A(n7240), .B(n7241), .Z(n7238) );
  AND U13095 ( .A(b[9]), .B(a[99]), .Z(n7237) );
  XOR U13096 ( .A(n7242), .B(n6871), .Z(n6873) );
  XOR U13097 ( .A(n7243), .B(n7244), .Z(n6871) );
  AND U13098 ( .A(n7245), .B(n7246), .Z(n7243) );
  AND U13099 ( .A(b[7]), .B(a[101]), .Z(n7242) );
  XOR U13100 ( .A(n7247), .B(n6876), .Z(n6878) );
  XOR U13101 ( .A(n7248), .B(n7249), .Z(n6876) );
  AND U13102 ( .A(n7250), .B(n7251), .Z(n7248) );
  AND U13103 ( .A(b[6]), .B(a[102]), .Z(n7247) );
  XOR U13104 ( .A(n7252), .B(n6881), .Z(n6883) );
  XOR U13105 ( .A(n7253), .B(n7254), .Z(n6881) );
  AND U13106 ( .A(n7255), .B(n7256), .Z(n7253) );
  AND U13107 ( .A(b[5]), .B(a[103]), .Z(n7252) );
  XOR U13108 ( .A(n7257), .B(n6886), .Z(n6888) );
  XOR U13109 ( .A(n7258), .B(n7259), .Z(n6886) );
  AND U13110 ( .A(n7260), .B(n7261), .Z(n7258) );
  AND U13111 ( .A(b[4]), .B(a[104]), .Z(n7257) );
  XOR U13112 ( .A(n7262), .B(n6895), .Z(n6897) );
  XNOR U13113 ( .A(n7263), .B(n7264), .Z(n6895) );
  ANDN U13114 ( .B(n7265), .A(n7266), .Z(n7263) );
  AND U13115 ( .A(b[3]), .B(a[105]), .Z(n7262) );
  NANDN U13116 ( .A(n7267), .B(n7268), .Z(n6898) );
  XOR U13117 ( .A(n7269), .B(n6890), .Z(n6892) );
  XNOR U13118 ( .A(n7270), .B(n7271), .Z(n6890) );
  OR U13119 ( .A(n7272), .B(n7273), .Z(n7271) );
  AND U13120 ( .A(b[2]), .B(a[106]), .Z(n7269) );
  XNOR U13121 ( .A(n7274), .B(n7275), .Z(swire[107]) );
  XOR U13122 ( .A(n7268), .B(n7276), .Z(n7275) );
  NAND U13123 ( .A(a[107]), .B(b[0]), .Z(n7267) );
  XOR U13124 ( .A(n7273), .B(n7272), .Z(n7268) );
  XOR U13125 ( .A(n7270), .B(n7277), .Z(n7272) );
  NAND U13126 ( .A(b[1]), .B(a[106]), .Z(n7277) );
  XOR U13127 ( .A(n7270), .B(n7266), .Z(n7278) );
  XOR U13128 ( .A(n7279), .B(n7264), .Z(n7266) );
  AND U13129 ( .A(b[2]), .B(a[105]), .Z(n7279) );
  ANDN U13130 ( .B(n7280), .A(n7281), .Z(n7270) );
  XOR U13131 ( .A(n7264), .B(n7260), .Z(n7282) );
  XNOR U13132 ( .A(n7259), .B(n7255), .Z(n7283) );
  XNOR U13133 ( .A(n7254), .B(n7250), .Z(n7284) );
  XNOR U13134 ( .A(n7249), .B(n7245), .Z(n7285) );
  XNOR U13135 ( .A(n7236), .B(n7235), .Z(n7286) );
  XOR U13136 ( .A(n7287), .B(n7234), .Z(n7235) );
  AND U13137 ( .A(b[7]), .B(a[100]), .Z(n7287) );
  XNOR U13138 ( .A(n7234), .B(n7240), .Z(n7288) );
  XNOR U13139 ( .A(n7239), .B(n7231), .Z(n7289) );
  XNOR U13140 ( .A(n7230), .B(n7226), .Z(n7290) );
  XNOR U13141 ( .A(n7225), .B(n7221), .Z(n7291) );
  XNOR U13142 ( .A(n7220), .B(n7216), .Z(n7292) );
  XNOR U13143 ( .A(n7207), .B(n7206), .Z(n7293) );
  XOR U13144 ( .A(n7294), .B(n7205), .Z(n7206) );
  AND U13145 ( .A(b[13]), .B(a[94]), .Z(n7294) );
  XNOR U13146 ( .A(n7205), .B(n7211), .Z(n7295) );
  XNOR U13147 ( .A(n7210), .B(n7202), .Z(n7296) );
  XNOR U13148 ( .A(n7201), .B(n7197), .Z(n7297) );
  XNOR U13149 ( .A(n7196), .B(n7192), .Z(n7298) );
  XNOR U13150 ( .A(n7191), .B(n7187), .Z(n7299) );
  XNOR U13151 ( .A(n7178), .B(n7177), .Z(n7300) );
  XOR U13152 ( .A(n7301), .B(n7176), .Z(n7177) );
  AND U13153 ( .A(b[19]), .B(a[88]), .Z(n7301) );
  XNOR U13154 ( .A(n7176), .B(n7182), .Z(n7302) );
  XNOR U13155 ( .A(n7181), .B(n7173), .Z(n7303) );
  XNOR U13156 ( .A(n7172), .B(n7168), .Z(n7304) );
  XNOR U13157 ( .A(n7167), .B(n7163), .Z(n7305) );
  XNOR U13158 ( .A(n7162), .B(n7158), .Z(n7306) );
  XNOR U13159 ( .A(n7149), .B(n7148), .Z(n7307) );
  XOR U13160 ( .A(n7308), .B(n7147), .Z(n7148) );
  AND U13161 ( .A(b[25]), .B(a[82]), .Z(n7308) );
  XNOR U13162 ( .A(n7147), .B(n7153), .Z(n7309) );
  XNOR U13163 ( .A(n7152), .B(n7144), .Z(n7310) );
  XNOR U13164 ( .A(n7143), .B(n7139), .Z(n7311) );
  XNOR U13165 ( .A(n7138), .B(n7134), .Z(n7312) );
  XNOR U13166 ( .A(n7133), .B(n7129), .Z(n7313) );
  XNOR U13167 ( .A(n7120), .B(n7119), .Z(n7314) );
  XOR U13168 ( .A(n7315), .B(n7118), .Z(n7119) );
  AND U13169 ( .A(b[31]), .B(a[76]), .Z(n7315) );
  XNOR U13170 ( .A(n7118), .B(n7124), .Z(n7316) );
  XNOR U13171 ( .A(n7123), .B(n7115), .Z(n7317) );
  XNOR U13172 ( .A(n7114), .B(n7110), .Z(n7318) );
  XNOR U13173 ( .A(n7109), .B(n7105), .Z(n7319) );
  XNOR U13174 ( .A(n7104), .B(n7100), .Z(n7320) );
  XNOR U13175 ( .A(n7091), .B(n7090), .Z(n7321) );
  XOR U13176 ( .A(n7322), .B(n7089), .Z(n7090) );
  AND U13177 ( .A(b[37]), .B(a[70]), .Z(n7322) );
  XNOR U13178 ( .A(n7089), .B(n7095), .Z(n7323) );
  XNOR U13179 ( .A(n7094), .B(n7086), .Z(n7324) );
  XNOR U13180 ( .A(n7085), .B(n7081), .Z(n7325) );
  XNOR U13181 ( .A(n7080), .B(n7076), .Z(n7326) );
  XNOR U13182 ( .A(n7075), .B(n7071), .Z(n7327) );
  XNOR U13183 ( .A(n7070), .B(n7066), .Z(n7328) );
  XNOR U13184 ( .A(n7065), .B(n7061), .Z(n7329) );
  XNOR U13185 ( .A(n7060), .B(n7056), .Z(n7330) );
  XNOR U13186 ( .A(n7055), .B(n7051), .Z(n7331) );
  XNOR U13187 ( .A(n7050), .B(n7046), .Z(n7332) );
  XNOR U13188 ( .A(n7045), .B(n7041), .Z(n7333) );
  XNOR U13189 ( .A(n7040), .B(n7036), .Z(n7334) );
  XNOR U13190 ( .A(n7035), .B(n7031), .Z(n7335) );
  XNOR U13191 ( .A(n7030), .B(n7026), .Z(n7336) );
  XNOR U13192 ( .A(n7025), .B(n7021), .Z(n7337) );
  XNOR U13193 ( .A(n7020), .B(n7016), .Z(n7338) );
  XNOR U13194 ( .A(n7015), .B(n7011), .Z(n7339) );
  XNOR U13195 ( .A(n7010), .B(n7006), .Z(n7340) );
  XNOR U13196 ( .A(n7005), .B(n7001), .Z(n7341) );
  XNOR U13197 ( .A(n7000), .B(n6996), .Z(n7342) );
  XNOR U13198 ( .A(n6995), .B(n6991), .Z(n7343) );
  XNOR U13199 ( .A(n6990), .B(n6986), .Z(n7344) );
  XOR U13200 ( .A(n6985), .B(n6982), .Z(n7345) );
  XOR U13201 ( .A(n7346), .B(n7347), .Z(n6982) );
  XOR U13202 ( .A(n6980), .B(n7348), .Z(n7347) );
  XOR U13203 ( .A(n7349), .B(n7350), .Z(n7348) );
  XOR U13204 ( .A(n7351), .B(n7352), .Z(n7350) );
  NAND U13205 ( .A(a[45]), .B(b[62]), .Z(n7352) );
  AND U13206 ( .A(a[44]), .B(b[63]), .Z(n7351) );
  XOR U13207 ( .A(n7353), .B(n7349), .Z(n7346) );
  XOR U13208 ( .A(n7354), .B(n7355), .Z(n7349) );
  ANDN U13209 ( .B(n7356), .A(n7357), .Z(n7354) );
  AND U13210 ( .A(a[46]), .B(b[61]), .Z(n7353) );
  XOR U13211 ( .A(n7358), .B(n6980), .Z(n6981) );
  XOR U13212 ( .A(n7359), .B(n7360), .Z(n6980) );
  AND U13213 ( .A(n7361), .B(n7362), .Z(n7359) );
  AND U13214 ( .A(a[47]), .B(b[60]), .Z(n7358) );
  XOR U13215 ( .A(n7363), .B(n6985), .Z(n6987) );
  XOR U13216 ( .A(n7364), .B(n7365), .Z(n6985) );
  AND U13217 ( .A(n7366), .B(n7367), .Z(n7364) );
  AND U13218 ( .A(a[48]), .B(b[59]), .Z(n7363) );
  XOR U13219 ( .A(n7368), .B(n6990), .Z(n6992) );
  XOR U13220 ( .A(n7369), .B(n7370), .Z(n6990) );
  AND U13221 ( .A(n7371), .B(n7372), .Z(n7369) );
  AND U13222 ( .A(a[49]), .B(b[58]), .Z(n7368) );
  XOR U13223 ( .A(n7373), .B(n6995), .Z(n6997) );
  XOR U13224 ( .A(n7374), .B(n7375), .Z(n6995) );
  AND U13225 ( .A(n7376), .B(n7377), .Z(n7374) );
  AND U13226 ( .A(a[50]), .B(b[57]), .Z(n7373) );
  XOR U13227 ( .A(n7378), .B(n7000), .Z(n7002) );
  XOR U13228 ( .A(n7379), .B(n7380), .Z(n7000) );
  AND U13229 ( .A(n7381), .B(n7382), .Z(n7379) );
  AND U13230 ( .A(a[51]), .B(b[56]), .Z(n7378) );
  XOR U13231 ( .A(n7383), .B(n7005), .Z(n7007) );
  XOR U13232 ( .A(n7384), .B(n7385), .Z(n7005) );
  AND U13233 ( .A(n7386), .B(n7387), .Z(n7384) );
  AND U13234 ( .A(a[52]), .B(b[55]), .Z(n7383) );
  XOR U13235 ( .A(n7388), .B(n7010), .Z(n7012) );
  XOR U13236 ( .A(n7389), .B(n7390), .Z(n7010) );
  AND U13237 ( .A(n7391), .B(n7392), .Z(n7389) );
  AND U13238 ( .A(a[53]), .B(b[54]), .Z(n7388) );
  XOR U13239 ( .A(n7393), .B(n7015), .Z(n7017) );
  XOR U13240 ( .A(n7394), .B(n7395), .Z(n7015) );
  AND U13241 ( .A(n7396), .B(n7397), .Z(n7394) );
  AND U13242 ( .A(b[53]), .B(a[54]), .Z(n7393) );
  XOR U13243 ( .A(n7398), .B(n7020), .Z(n7022) );
  XOR U13244 ( .A(n7399), .B(n7400), .Z(n7020) );
  AND U13245 ( .A(n7401), .B(n7402), .Z(n7399) );
  AND U13246 ( .A(b[52]), .B(a[55]), .Z(n7398) );
  XOR U13247 ( .A(n7403), .B(n7025), .Z(n7027) );
  XOR U13248 ( .A(n7404), .B(n7405), .Z(n7025) );
  AND U13249 ( .A(n7406), .B(n7407), .Z(n7404) );
  AND U13250 ( .A(b[51]), .B(a[56]), .Z(n7403) );
  XOR U13251 ( .A(n7408), .B(n7030), .Z(n7032) );
  XOR U13252 ( .A(n7409), .B(n7410), .Z(n7030) );
  AND U13253 ( .A(n7411), .B(n7412), .Z(n7409) );
  AND U13254 ( .A(b[50]), .B(a[57]), .Z(n7408) );
  XOR U13255 ( .A(n7413), .B(n7035), .Z(n7037) );
  XOR U13256 ( .A(n7414), .B(n7415), .Z(n7035) );
  AND U13257 ( .A(n7416), .B(n7417), .Z(n7414) );
  AND U13258 ( .A(b[49]), .B(a[58]), .Z(n7413) );
  XOR U13259 ( .A(n7418), .B(n7040), .Z(n7042) );
  XOR U13260 ( .A(n7419), .B(n7420), .Z(n7040) );
  AND U13261 ( .A(n7421), .B(n7422), .Z(n7419) );
  AND U13262 ( .A(b[48]), .B(a[59]), .Z(n7418) );
  XOR U13263 ( .A(n7423), .B(n7045), .Z(n7047) );
  XOR U13264 ( .A(n7424), .B(n7425), .Z(n7045) );
  AND U13265 ( .A(n7426), .B(n7427), .Z(n7424) );
  AND U13266 ( .A(b[47]), .B(a[60]), .Z(n7423) );
  XOR U13267 ( .A(n7428), .B(n7050), .Z(n7052) );
  XOR U13268 ( .A(n7429), .B(n7430), .Z(n7050) );
  AND U13269 ( .A(n7431), .B(n7432), .Z(n7429) );
  AND U13270 ( .A(b[46]), .B(a[61]), .Z(n7428) );
  XOR U13271 ( .A(n7433), .B(n7055), .Z(n7057) );
  XOR U13272 ( .A(n7434), .B(n7435), .Z(n7055) );
  AND U13273 ( .A(n7436), .B(n7437), .Z(n7434) );
  AND U13274 ( .A(b[45]), .B(a[62]), .Z(n7433) );
  XOR U13275 ( .A(n7438), .B(n7060), .Z(n7062) );
  XOR U13276 ( .A(n7439), .B(n7440), .Z(n7060) );
  AND U13277 ( .A(n7441), .B(n7442), .Z(n7439) );
  AND U13278 ( .A(b[44]), .B(a[63]), .Z(n7438) );
  XOR U13279 ( .A(n7443), .B(n7065), .Z(n7067) );
  XOR U13280 ( .A(n7444), .B(n7445), .Z(n7065) );
  AND U13281 ( .A(n7446), .B(n7447), .Z(n7444) );
  AND U13282 ( .A(b[43]), .B(a[64]), .Z(n7443) );
  XOR U13283 ( .A(n7448), .B(n7070), .Z(n7072) );
  XOR U13284 ( .A(n7449), .B(n7450), .Z(n7070) );
  AND U13285 ( .A(n7451), .B(n7452), .Z(n7449) );
  AND U13286 ( .A(b[42]), .B(a[65]), .Z(n7448) );
  XOR U13287 ( .A(n7453), .B(n7075), .Z(n7077) );
  XOR U13288 ( .A(n7454), .B(n7455), .Z(n7075) );
  AND U13289 ( .A(n7456), .B(n7457), .Z(n7454) );
  AND U13290 ( .A(b[41]), .B(a[66]), .Z(n7453) );
  XOR U13291 ( .A(n7458), .B(n7080), .Z(n7082) );
  XOR U13292 ( .A(n7459), .B(n7460), .Z(n7080) );
  AND U13293 ( .A(n7461), .B(n7462), .Z(n7459) );
  AND U13294 ( .A(b[40]), .B(a[67]), .Z(n7458) );
  XOR U13295 ( .A(n7463), .B(n7085), .Z(n7087) );
  XOR U13296 ( .A(n7464), .B(n7465), .Z(n7085) );
  AND U13297 ( .A(n7466), .B(n7467), .Z(n7464) );
  AND U13298 ( .A(b[39]), .B(a[68]), .Z(n7463) );
  XOR U13299 ( .A(n7468), .B(n7469), .Z(n7089) );
  AND U13300 ( .A(n7470), .B(n7471), .Z(n7468) );
  XOR U13301 ( .A(n7472), .B(n7094), .Z(n7096) );
  XOR U13302 ( .A(n7473), .B(n7474), .Z(n7094) );
  AND U13303 ( .A(n7475), .B(n7476), .Z(n7473) );
  AND U13304 ( .A(b[38]), .B(a[69]), .Z(n7472) );
  XOR U13305 ( .A(n7477), .B(n7099), .Z(n7101) );
  XOR U13306 ( .A(n7478), .B(n7479), .Z(n7099) );
  AND U13307 ( .A(n7480), .B(n7481), .Z(n7478) );
  AND U13308 ( .A(b[36]), .B(a[71]), .Z(n7477) );
  XOR U13309 ( .A(n7482), .B(n7104), .Z(n7106) );
  XOR U13310 ( .A(n7483), .B(n7484), .Z(n7104) );
  AND U13311 ( .A(n7485), .B(n7486), .Z(n7483) );
  AND U13312 ( .A(b[35]), .B(a[72]), .Z(n7482) );
  XOR U13313 ( .A(n7487), .B(n7109), .Z(n7111) );
  XOR U13314 ( .A(n7488), .B(n7489), .Z(n7109) );
  AND U13315 ( .A(n7490), .B(n7491), .Z(n7488) );
  AND U13316 ( .A(b[34]), .B(a[73]), .Z(n7487) );
  XOR U13317 ( .A(n7492), .B(n7114), .Z(n7116) );
  XOR U13318 ( .A(n7493), .B(n7494), .Z(n7114) );
  AND U13319 ( .A(n7495), .B(n7496), .Z(n7493) );
  AND U13320 ( .A(b[33]), .B(a[74]), .Z(n7492) );
  XOR U13321 ( .A(n7497), .B(n7498), .Z(n7118) );
  AND U13322 ( .A(n7499), .B(n7500), .Z(n7497) );
  XOR U13323 ( .A(n7501), .B(n7123), .Z(n7125) );
  XOR U13324 ( .A(n7502), .B(n7503), .Z(n7123) );
  AND U13325 ( .A(n7504), .B(n7505), .Z(n7502) );
  AND U13326 ( .A(b[32]), .B(a[75]), .Z(n7501) );
  XOR U13327 ( .A(n7506), .B(n7128), .Z(n7130) );
  XOR U13328 ( .A(n7507), .B(n7508), .Z(n7128) );
  AND U13329 ( .A(n7509), .B(n7510), .Z(n7507) );
  AND U13330 ( .A(b[30]), .B(a[77]), .Z(n7506) );
  XOR U13331 ( .A(n7511), .B(n7133), .Z(n7135) );
  XOR U13332 ( .A(n7512), .B(n7513), .Z(n7133) );
  AND U13333 ( .A(n7514), .B(n7515), .Z(n7512) );
  AND U13334 ( .A(b[29]), .B(a[78]), .Z(n7511) );
  XOR U13335 ( .A(n7516), .B(n7138), .Z(n7140) );
  XOR U13336 ( .A(n7517), .B(n7518), .Z(n7138) );
  AND U13337 ( .A(n7519), .B(n7520), .Z(n7517) );
  AND U13338 ( .A(b[28]), .B(a[79]), .Z(n7516) );
  XOR U13339 ( .A(n7521), .B(n7143), .Z(n7145) );
  XOR U13340 ( .A(n7522), .B(n7523), .Z(n7143) );
  AND U13341 ( .A(n7524), .B(n7525), .Z(n7522) );
  AND U13342 ( .A(b[27]), .B(a[80]), .Z(n7521) );
  XOR U13343 ( .A(n7526), .B(n7527), .Z(n7147) );
  AND U13344 ( .A(n7528), .B(n7529), .Z(n7526) );
  XOR U13345 ( .A(n7530), .B(n7152), .Z(n7154) );
  XOR U13346 ( .A(n7531), .B(n7532), .Z(n7152) );
  AND U13347 ( .A(n7533), .B(n7534), .Z(n7531) );
  AND U13348 ( .A(b[26]), .B(a[81]), .Z(n7530) );
  XOR U13349 ( .A(n7535), .B(n7157), .Z(n7159) );
  XOR U13350 ( .A(n7536), .B(n7537), .Z(n7157) );
  AND U13351 ( .A(n7538), .B(n7539), .Z(n7536) );
  AND U13352 ( .A(b[24]), .B(a[83]), .Z(n7535) );
  XOR U13353 ( .A(n7540), .B(n7162), .Z(n7164) );
  XOR U13354 ( .A(n7541), .B(n7542), .Z(n7162) );
  AND U13355 ( .A(n7543), .B(n7544), .Z(n7541) );
  AND U13356 ( .A(b[23]), .B(a[84]), .Z(n7540) );
  XOR U13357 ( .A(n7545), .B(n7167), .Z(n7169) );
  XOR U13358 ( .A(n7546), .B(n7547), .Z(n7167) );
  AND U13359 ( .A(n7548), .B(n7549), .Z(n7546) );
  AND U13360 ( .A(b[22]), .B(a[85]), .Z(n7545) );
  XOR U13361 ( .A(n7550), .B(n7172), .Z(n7174) );
  XOR U13362 ( .A(n7551), .B(n7552), .Z(n7172) );
  AND U13363 ( .A(n7553), .B(n7554), .Z(n7551) );
  AND U13364 ( .A(b[21]), .B(a[86]), .Z(n7550) );
  XOR U13365 ( .A(n7555), .B(n7556), .Z(n7176) );
  AND U13366 ( .A(n7557), .B(n7558), .Z(n7555) );
  XOR U13367 ( .A(n7559), .B(n7181), .Z(n7183) );
  XOR U13368 ( .A(n7560), .B(n7561), .Z(n7181) );
  AND U13369 ( .A(n7562), .B(n7563), .Z(n7560) );
  AND U13370 ( .A(b[20]), .B(a[87]), .Z(n7559) );
  XOR U13371 ( .A(n7564), .B(n7186), .Z(n7188) );
  XOR U13372 ( .A(n7565), .B(n7566), .Z(n7186) );
  AND U13373 ( .A(n7567), .B(n7568), .Z(n7565) );
  AND U13374 ( .A(b[18]), .B(a[89]), .Z(n7564) );
  XOR U13375 ( .A(n7569), .B(n7191), .Z(n7193) );
  XOR U13376 ( .A(n7570), .B(n7571), .Z(n7191) );
  AND U13377 ( .A(n7572), .B(n7573), .Z(n7570) );
  AND U13378 ( .A(b[17]), .B(a[90]), .Z(n7569) );
  XOR U13379 ( .A(n7574), .B(n7196), .Z(n7198) );
  XOR U13380 ( .A(n7575), .B(n7576), .Z(n7196) );
  AND U13381 ( .A(n7577), .B(n7578), .Z(n7575) );
  AND U13382 ( .A(b[16]), .B(a[91]), .Z(n7574) );
  XOR U13383 ( .A(n7579), .B(n7201), .Z(n7203) );
  XOR U13384 ( .A(n7580), .B(n7581), .Z(n7201) );
  AND U13385 ( .A(n7582), .B(n7583), .Z(n7580) );
  AND U13386 ( .A(b[15]), .B(a[92]), .Z(n7579) );
  XOR U13387 ( .A(n7584), .B(n7585), .Z(n7205) );
  AND U13388 ( .A(n7586), .B(n7587), .Z(n7584) );
  XOR U13389 ( .A(n7588), .B(n7210), .Z(n7212) );
  XOR U13390 ( .A(n7589), .B(n7590), .Z(n7210) );
  AND U13391 ( .A(n7591), .B(n7592), .Z(n7589) );
  AND U13392 ( .A(b[14]), .B(a[93]), .Z(n7588) );
  XOR U13393 ( .A(n7593), .B(n7215), .Z(n7217) );
  XOR U13394 ( .A(n7594), .B(n7595), .Z(n7215) );
  AND U13395 ( .A(n7596), .B(n7597), .Z(n7594) );
  AND U13396 ( .A(b[12]), .B(a[95]), .Z(n7593) );
  XOR U13397 ( .A(n7598), .B(n7220), .Z(n7222) );
  XOR U13398 ( .A(n7599), .B(n7600), .Z(n7220) );
  AND U13399 ( .A(n7601), .B(n7602), .Z(n7599) );
  AND U13400 ( .A(b[11]), .B(a[96]), .Z(n7598) );
  XOR U13401 ( .A(n7603), .B(n7225), .Z(n7227) );
  XOR U13402 ( .A(n7604), .B(n7605), .Z(n7225) );
  AND U13403 ( .A(n7606), .B(n7607), .Z(n7604) );
  AND U13404 ( .A(b[10]), .B(a[97]), .Z(n7603) );
  XOR U13405 ( .A(n7608), .B(n7230), .Z(n7232) );
  XOR U13406 ( .A(n7609), .B(n7610), .Z(n7230) );
  AND U13407 ( .A(n7611), .B(n7612), .Z(n7609) );
  AND U13408 ( .A(b[9]), .B(a[98]), .Z(n7608) );
  XOR U13409 ( .A(n7613), .B(n7614), .Z(n7234) );
  AND U13410 ( .A(n7615), .B(n7616), .Z(n7613) );
  XOR U13411 ( .A(n7617), .B(n7239), .Z(n7241) );
  XOR U13412 ( .A(n7618), .B(n7619), .Z(n7239) );
  AND U13413 ( .A(n7620), .B(n7621), .Z(n7618) );
  AND U13414 ( .A(b[8]), .B(a[99]), .Z(n7617) );
  XOR U13415 ( .A(n7622), .B(n7244), .Z(n7246) );
  XOR U13416 ( .A(n7623), .B(n7624), .Z(n7244) );
  AND U13417 ( .A(n7625), .B(n7626), .Z(n7623) );
  AND U13418 ( .A(b[6]), .B(a[101]), .Z(n7622) );
  XOR U13419 ( .A(n7627), .B(n7249), .Z(n7251) );
  XOR U13420 ( .A(n7628), .B(n7629), .Z(n7249) );
  AND U13421 ( .A(n7630), .B(n7631), .Z(n7628) );
  AND U13422 ( .A(b[5]), .B(a[102]), .Z(n7627) );
  XOR U13423 ( .A(n7632), .B(n7254), .Z(n7256) );
  XOR U13424 ( .A(n7633), .B(n7634), .Z(n7254) );
  AND U13425 ( .A(n7635), .B(n7636), .Z(n7633) );
  AND U13426 ( .A(b[4]), .B(a[103]), .Z(n7632) );
  XNOR U13427 ( .A(n7637), .B(n7638), .Z(n7264) );
  NANDN U13428 ( .A(n7639), .B(n7640), .Z(n7638) );
  XOR U13429 ( .A(n7641), .B(n7259), .Z(n7261) );
  XNOR U13430 ( .A(n7642), .B(n7643), .Z(n7259) );
  AND U13431 ( .A(n7644), .B(n7645), .Z(n7642) );
  AND U13432 ( .A(b[3]), .B(a[104]), .Z(n7641) );
  XOR U13433 ( .A(n7646), .B(n7647), .Z(swire[106]) );
  XOR U13434 ( .A(n7281), .B(n7280), .Z(n7648) );
  XNOR U13435 ( .A(n7639), .B(n7640), .Z(n7280) );
  XOR U13436 ( .A(n7637), .B(n7649), .Z(n7640) );
  NAND U13437 ( .A(b[1]), .B(a[105]), .Z(n7649) );
  XOR U13438 ( .A(n7645), .B(n7650), .Z(n7639) );
  XOR U13439 ( .A(n7637), .B(n7644), .Z(n7650) );
  XNOR U13440 ( .A(n7651), .B(n7643), .Z(n7644) );
  AND U13441 ( .A(b[2]), .B(a[104]), .Z(n7651) );
  NANDN U13442 ( .A(n7652), .B(n7653), .Z(n7637) );
  XOR U13443 ( .A(n7643), .B(n7635), .Z(n7654) );
  XNOR U13444 ( .A(n7634), .B(n7630), .Z(n7655) );
  XNOR U13445 ( .A(n7629), .B(n7625), .Z(n7656) );
  XNOR U13446 ( .A(n7616), .B(n7615), .Z(n7657) );
  XOR U13447 ( .A(n7658), .B(n7614), .Z(n7615) );
  AND U13448 ( .A(b[6]), .B(a[100]), .Z(n7658) );
  XNOR U13449 ( .A(n7614), .B(n7620), .Z(n7659) );
  XNOR U13450 ( .A(n7619), .B(n7611), .Z(n7660) );
  XNOR U13451 ( .A(n7610), .B(n7606), .Z(n7661) );
  XNOR U13452 ( .A(n7605), .B(n7601), .Z(n7662) );
  XNOR U13453 ( .A(n7600), .B(n7596), .Z(n7663) );
  XNOR U13454 ( .A(n7587), .B(n7586), .Z(n7664) );
  XOR U13455 ( .A(n7665), .B(n7585), .Z(n7586) );
  AND U13456 ( .A(b[12]), .B(a[94]), .Z(n7665) );
  XNOR U13457 ( .A(n7585), .B(n7591), .Z(n7666) );
  XNOR U13458 ( .A(n7590), .B(n7582), .Z(n7667) );
  XNOR U13459 ( .A(n7581), .B(n7577), .Z(n7668) );
  XNOR U13460 ( .A(n7576), .B(n7572), .Z(n7669) );
  XNOR U13461 ( .A(n7571), .B(n7567), .Z(n7670) );
  XNOR U13462 ( .A(n7558), .B(n7557), .Z(n7671) );
  XOR U13463 ( .A(n7672), .B(n7556), .Z(n7557) );
  AND U13464 ( .A(b[18]), .B(a[88]), .Z(n7672) );
  XNOR U13465 ( .A(n7556), .B(n7562), .Z(n7673) );
  XNOR U13466 ( .A(n7561), .B(n7553), .Z(n7674) );
  XNOR U13467 ( .A(n7552), .B(n7548), .Z(n7675) );
  XNOR U13468 ( .A(n7547), .B(n7543), .Z(n7676) );
  XNOR U13469 ( .A(n7542), .B(n7538), .Z(n7677) );
  XNOR U13470 ( .A(n7529), .B(n7528), .Z(n7678) );
  XOR U13471 ( .A(n7679), .B(n7527), .Z(n7528) );
  AND U13472 ( .A(b[24]), .B(a[82]), .Z(n7679) );
  XNOR U13473 ( .A(n7527), .B(n7533), .Z(n7680) );
  XNOR U13474 ( .A(n7532), .B(n7524), .Z(n7681) );
  XNOR U13475 ( .A(n7523), .B(n7519), .Z(n7682) );
  XNOR U13476 ( .A(n7518), .B(n7514), .Z(n7683) );
  XNOR U13477 ( .A(n7513), .B(n7509), .Z(n7684) );
  XNOR U13478 ( .A(n7500), .B(n7499), .Z(n7685) );
  XOR U13479 ( .A(n7686), .B(n7498), .Z(n7499) );
  AND U13480 ( .A(b[30]), .B(a[76]), .Z(n7686) );
  XNOR U13481 ( .A(n7498), .B(n7504), .Z(n7687) );
  XNOR U13482 ( .A(n7503), .B(n7495), .Z(n7688) );
  XNOR U13483 ( .A(n7494), .B(n7490), .Z(n7689) );
  XNOR U13484 ( .A(n7489), .B(n7485), .Z(n7690) );
  XNOR U13485 ( .A(n7484), .B(n7480), .Z(n7691) );
  XNOR U13486 ( .A(n7471), .B(n7470), .Z(n7692) );
  XOR U13487 ( .A(n7693), .B(n7469), .Z(n7470) );
  AND U13488 ( .A(b[36]), .B(a[70]), .Z(n7693) );
  XNOR U13489 ( .A(n7469), .B(n7475), .Z(n7694) );
  XNOR U13490 ( .A(n7474), .B(n7466), .Z(n7695) );
  XNOR U13491 ( .A(n7465), .B(n7461), .Z(n7696) );
  XNOR U13492 ( .A(n7460), .B(n7456), .Z(n7697) );
  XNOR U13493 ( .A(n7455), .B(n7451), .Z(n7698) );
  XNOR U13494 ( .A(n7450), .B(n7446), .Z(n7699) );
  XNOR U13495 ( .A(n7445), .B(n7441), .Z(n7700) );
  XNOR U13496 ( .A(n7440), .B(n7436), .Z(n7701) );
  XNOR U13497 ( .A(n7435), .B(n7431), .Z(n7702) );
  XNOR U13498 ( .A(n7430), .B(n7426), .Z(n7703) );
  XNOR U13499 ( .A(n7425), .B(n7421), .Z(n7704) );
  XNOR U13500 ( .A(n7420), .B(n7416), .Z(n7705) );
  XNOR U13501 ( .A(n7415), .B(n7411), .Z(n7706) );
  XNOR U13502 ( .A(n7410), .B(n7406), .Z(n7707) );
  XNOR U13503 ( .A(n7405), .B(n7401), .Z(n7708) );
  XNOR U13504 ( .A(n7400), .B(n7396), .Z(n7709) );
  XNOR U13505 ( .A(n7395), .B(n7391), .Z(n7710) );
  XNOR U13506 ( .A(n7390), .B(n7386), .Z(n7711) );
  XNOR U13507 ( .A(n7385), .B(n7381), .Z(n7712) );
  XNOR U13508 ( .A(n7380), .B(n7376), .Z(n7713) );
  XNOR U13509 ( .A(n7375), .B(n7371), .Z(n7714) );
  XNOR U13510 ( .A(n7370), .B(n7366), .Z(n7715) );
  XNOR U13511 ( .A(n7365), .B(n7361), .Z(n7716) );
  XOR U13512 ( .A(n7360), .B(n7357), .Z(n7717) );
  XOR U13513 ( .A(n7718), .B(n7719), .Z(n7357) );
  XOR U13514 ( .A(n7355), .B(n7720), .Z(n7719) );
  XOR U13515 ( .A(n7721), .B(n7722), .Z(n7720) );
  XOR U13516 ( .A(n7723), .B(n7724), .Z(n7722) );
  NAND U13517 ( .A(a[44]), .B(b[62]), .Z(n7724) );
  AND U13518 ( .A(a[43]), .B(b[63]), .Z(n7723) );
  XOR U13519 ( .A(n7725), .B(n7721), .Z(n7718) );
  XOR U13520 ( .A(n7726), .B(n7727), .Z(n7721) );
  ANDN U13521 ( .B(n7728), .A(n7729), .Z(n7726) );
  AND U13522 ( .A(a[45]), .B(b[61]), .Z(n7725) );
  XOR U13523 ( .A(n7730), .B(n7355), .Z(n7356) );
  XOR U13524 ( .A(n7731), .B(n7732), .Z(n7355) );
  AND U13525 ( .A(n7733), .B(n7734), .Z(n7731) );
  AND U13526 ( .A(a[46]), .B(b[60]), .Z(n7730) );
  XOR U13527 ( .A(n7735), .B(n7360), .Z(n7362) );
  XOR U13528 ( .A(n7736), .B(n7737), .Z(n7360) );
  AND U13529 ( .A(n7738), .B(n7739), .Z(n7736) );
  AND U13530 ( .A(a[47]), .B(b[59]), .Z(n7735) );
  XOR U13531 ( .A(n7740), .B(n7365), .Z(n7367) );
  XOR U13532 ( .A(n7741), .B(n7742), .Z(n7365) );
  AND U13533 ( .A(n7743), .B(n7744), .Z(n7741) );
  AND U13534 ( .A(a[48]), .B(b[58]), .Z(n7740) );
  XOR U13535 ( .A(n7745), .B(n7370), .Z(n7372) );
  XOR U13536 ( .A(n7746), .B(n7747), .Z(n7370) );
  AND U13537 ( .A(n7748), .B(n7749), .Z(n7746) );
  AND U13538 ( .A(a[49]), .B(b[57]), .Z(n7745) );
  XOR U13539 ( .A(n7750), .B(n7375), .Z(n7377) );
  XOR U13540 ( .A(n7751), .B(n7752), .Z(n7375) );
  AND U13541 ( .A(n7753), .B(n7754), .Z(n7751) );
  AND U13542 ( .A(a[50]), .B(b[56]), .Z(n7750) );
  XOR U13543 ( .A(n7755), .B(n7380), .Z(n7382) );
  XOR U13544 ( .A(n7756), .B(n7757), .Z(n7380) );
  AND U13545 ( .A(n7758), .B(n7759), .Z(n7756) );
  AND U13546 ( .A(a[51]), .B(b[55]), .Z(n7755) );
  XOR U13547 ( .A(n7760), .B(n7385), .Z(n7387) );
  XOR U13548 ( .A(n7761), .B(n7762), .Z(n7385) );
  AND U13549 ( .A(n7763), .B(n7764), .Z(n7761) );
  AND U13550 ( .A(a[52]), .B(b[54]), .Z(n7760) );
  XOR U13551 ( .A(n7765), .B(n7390), .Z(n7392) );
  XOR U13552 ( .A(n7766), .B(n7767), .Z(n7390) );
  AND U13553 ( .A(n7768), .B(n7769), .Z(n7766) );
  AND U13554 ( .A(a[53]), .B(b[53]), .Z(n7765) );
  XOR U13555 ( .A(n7770), .B(n7395), .Z(n7397) );
  XOR U13556 ( .A(n7771), .B(n7772), .Z(n7395) );
  AND U13557 ( .A(n7773), .B(n7774), .Z(n7771) );
  AND U13558 ( .A(b[52]), .B(a[54]), .Z(n7770) );
  XOR U13559 ( .A(n7775), .B(n7400), .Z(n7402) );
  XOR U13560 ( .A(n7776), .B(n7777), .Z(n7400) );
  AND U13561 ( .A(n7778), .B(n7779), .Z(n7776) );
  AND U13562 ( .A(b[51]), .B(a[55]), .Z(n7775) );
  XOR U13563 ( .A(n7780), .B(n7405), .Z(n7407) );
  XOR U13564 ( .A(n7781), .B(n7782), .Z(n7405) );
  AND U13565 ( .A(n7783), .B(n7784), .Z(n7781) );
  AND U13566 ( .A(b[50]), .B(a[56]), .Z(n7780) );
  XOR U13567 ( .A(n7785), .B(n7410), .Z(n7412) );
  XOR U13568 ( .A(n7786), .B(n7787), .Z(n7410) );
  AND U13569 ( .A(n7788), .B(n7789), .Z(n7786) );
  AND U13570 ( .A(b[49]), .B(a[57]), .Z(n7785) );
  XOR U13571 ( .A(n7790), .B(n7415), .Z(n7417) );
  XOR U13572 ( .A(n7791), .B(n7792), .Z(n7415) );
  AND U13573 ( .A(n7793), .B(n7794), .Z(n7791) );
  AND U13574 ( .A(b[48]), .B(a[58]), .Z(n7790) );
  XOR U13575 ( .A(n7795), .B(n7420), .Z(n7422) );
  XOR U13576 ( .A(n7796), .B(n7797), .Z(n7420) );
  AND U13577 ( .A(n7798), .B(n7799), .Z(n7796) );
  AND U13578 ( .A(b[47]), .B(a[59]), .Z(n7795) );
  XOR U13579 ( .A(n7800), .B(n7425), .Z(n7427) );
  XOR U13580 ( .A(n7801), .B(n7802), .Z(n7425) );
  AND U13581 ( .A(n7803), .B(n7804), .Z(n7801) );
  AND U13582 ( .A(b[46]), .B(a[60]), .Z(n7800) );
  XOR U13583 ( .A(n7805), .B(n7430), .Z(n7432) );
  XOR U13584 ( .A(n7806), .B(n7807), .Z(n7430) );
  AND U13585 ( .A(n7808), .B(n7809), .Z(n7806) );
  AND U13586 ( .A(b[45]), .B(a[61]), .Z(n7805) );
  XOR U13587 ( .A(n7810), .B(n7435), .Z(n7437) );
  XOR U13588 ( .A(n7811), .B(n7812), .Z(n7435) );
  AND U13589 ( .A(n7813), .B(n7814), .Z(n7811) );
  AND U13590 ( .A(b[44]), .B(a[62]), .Z(n7810) );
  XOR U13591 ( .A(n7815), .B(n7440), .Z(n7442) );
  XOR U13592 ( .A(n7816), .B(n7817), .Z(n7440) );
  AND U13593 ( .A(n7818), .B(n7819), .Z(n7816) );
  AND U13594 ( .A(b[43]), .B(a[63]), .Z(n7815) );
  XOR U13595 ( .A(n7820), .B(n7445), .Z(n7447) );
  XOR U13596 ( .A(n7821), .B(n7822), .Z(n7445) );
  AND U13597 ( .A(n7823), .B(n7824), .Z(n7821) );
  AND U13598 ( .A(b[42]), .B(a[64]), .Z(n7820) );
  XOR U13599 ( .A(n7825), .B(n7450), .Z(n7452) );
  XOR U13600 ( .A(n7826), .B(n7827), .Z(n7450) );
  AND U13601 ( .A(n7828), .B(n7829), .Z(n7826) );
  AND U13602 ( .A(b[41]), .B(a[65]), .Z(n7825) );
  XOR U13603 ( .A(n7830), .B(n7455), .Z(n7457) );
  XOR U13604 ( .A(n7831), .B(n7832), .Z(n7455) );
  AND U13605 ( .A(n7833), .B(n7834), .Z(n7831) );
  AND U13606 ( .A(b[40]), .B(a[66]), .Z(n7830) );
  XOR U13607 ( .A(n7835), .B(n7460), .Z(n7462) );
  XOR U13608 ( .A(n7836), .B(n7837), .Z(n7460) );
  AND U13609 ( .A(n7838), .B(n7839), .Z(n7836) );
  AND U13610 ( .A(b[39]), .B(a[67]), .Z(n7835) );
  XOR U13611 ( .A(n7840), .B(n7465), .Z(n7467) );
  XOR U13612 ( .A(n7841), .B(n7842), .Z(n7465) );
  AND U13613 ( .A(n7843), .B(n7844), .Z(n7841) );
  AND U13614 ( .A(b[38]), .B(a[68]), .Z(n7840) );
  XOR U13615 ( .A(n7845), .B(n7846), .Z(n7469) );
  AND U13616 ( .A(n7847), .B(n7848), .Z(n7845) );
  XOR U13617 ( .A(n7849), .B(n7474), .Z(n7476) );
  XOR U13618 ( .A(n7850), .B(n7851), .Z(n7474) );
  AND U13619 ( .A(n7852), .B(n7853), .Z(n7850) );
  AND U13620 ( .A(b[37]), .B(a[69]), .Z(n7849) );
  XOR U13621 ( .A(n7854), .B(n7479), .Z(n7481) );
  XOR U13622 ( .A(n7855), .B(n7856), .Z(n7479) );
  AND U13623 ( .A(n7857), .B(n7858), .Z(n7855) );
  AND U13624 ( .A(b[35]), .B(a[71]), .Z(n7854) );
  XOR U13625 ( .A(n7859), .B(n7484), .Z(n7486) );
  XOR U13626 ( .A(n7860), .B(n7861), .Z(n7484) );
  AND U13627 ( .A(n7862), .B(n7863), .Z(n7860) );
  AND U13628 ( .A(b[34]), .B(a[72]), .Z(n7859) );
  XOR U13629 ( .A(n7864), .B(n7489), .Z(n7491) );
  XOR U13630 ( .A(n7865), .B(n7866), .Z(n7489) );
  AND U13631 ( .A(n7867), .B(n7868), .Z(n7865) );
  AND U13632 ( .A(b[33]), .B(a[73]), .Z(n7864) );
  XOR U13633 ( .A(n7869), .B(n7494), .Z(n7496) );
  XOR U13634 ( .A(n7870), .B(n7871), .Z(n7494) );
  AND U13635 ( .A(n7872), .B(n7873), .Z(n7870) );
  AND U13636 ( .A(b[32]), .B(a[74]), .Z(n7869) );
  XOR U13637 ( .A(n7874), .B(n7875), .Z(n7498) );
  AND U13638 ( .A(n7876), .B(n7877), .Z(n7874) );
  XOR U13639 ( .A(n7878), .B(n7503), .Z(n7505) );
  XOR U13640 ( .A(n7879), .B(n7880), .Z(n7503) );
  AND U13641 ( .A(n7881), .B(n7882), .Z(n7879) );
  AND U13642 ( .A(b[31]), .B(a[75]), .Z(n7878) );
  XOR U13643 ( .A(n7883), .B(n7508), .Z(n7510) );
  XOR U13644 ( .A(n7884), .B(n7885), .Z(n7508) );
  AND U13645 ( .A(n7886), .B(n7887), .Z(n7884) );
  AND U13646 ( .A(b[29]), .B(a[77]), .Z(n7883) );
  XOR U13647 ( .A(n7888), .B(n7513), .Z(n7515) );
  XOR U13648 ( .A(n7889), .B(n7890), .Z(n7513) );
  AND U13649 ( .A(n7891), .B(n7892), .Z(n7889) );
  AND U13650 ( .A(b[28]), .B(a[78]), .Z(n7888) );
  XOR U13651 ( .A(n7893), .B(n7518), .Z(n7520) );
  XOR U13652 ( .A(n7894), .B(n7895), .Z(n7518) );
  AND U13653 ( .A(n7896), .B(n7897), .Z(n7894) );
  AND U13654 ( .A(b[27]), .B(a[79]), .Z(n7893) );
  XOR U13655 ( .A(n7898), .B(n7523), .Z(n7525) );
  XOR U13656 ( .A(n7899), .B(n7900), .Z(n7523) );
  AND U13657 ( .A(n7901), .B(n7902), .Z(n7899) );
  AND U13658 ( .A(b[26]), .B(a[80]), .Z(n7898) );
  XOR U13659 ( .A(n7903), .B(n7904), .Z(n7527) );
  AND U13660 ( .A(n7905), .B(n7906), .Z(n7903) );
  XOR U13661 ( .A(n7907), .B(n7532), .Z(n7534) );
  XOR U13662 ( .A(n7908), .B(n7909), .Z(n7532) );
  AND U13663 ( .A(n7910), .B(n7911), .Z(n7908) );
  AND U13664 ( .A(b[25]), .B(a[81]), .Z(n7907) );
  XOR U13665 ( .A(n7912), .B(n7537), .Z(n7539) );
  XOR U13666 ( .A(n7913), .B(n7914), .Z(n7537) );
  AND U13667 ( .A(n7915), .B(n7916), .Z(n7913) );
  AND U13668 ( .A(b[23]), .B(a[83]), .Z(n7912) );
  XOR U13669 ( .A(n7917), .B(n7542), .Z(n7544) );
  XOR U13670 ( .A(n7918), .B(n7919), .Z(n7542) );
  AND U13671 ( .A(n7920), .B(n7921), .Z(n7918) );
  AND U13672 ( .A(b[22]), .B(a[84]), .Z(n7917) );
  XOR U13673 ( .A(n7922), .B(n7547), .Z(n7549) );
  XOR U13674 ( .A(n7923), .B(n7924), .Z(n7547) );
  AND U13675 ( .A(n7925), .B(n7926), .Z(n7923) );
  AND U13676 ( .A(b[21]), .B(a[85]), .Z(n7922) );
  XOR U13677 ( .A(n7927), .B(n7552), .Z(n7554) );
  XOR U13678 ( .A(n7928), .B(n7929), .Z(n7552) );
  AND U13679 ( .A(n7930), .B(n7931), .Z(n7928) );
  AND U13680 ( .A(b[20]), .B(a[86]), .Z(n7927) );
  XOR U13681 ( .A(n7932), .B(n7933), .Z(n7556) );
  AND U13682 ( .A(n7934), .B(n7935), .Z(n7932) );
  XOR U13683 ( .A(n7936), .B(n7561), .Z(n7563) );
  XOR U13684 ( .A(n7937), .B(n7938), .Z(n7561) );
  AND U13685 ( .A(n7939), .B(n7940), .Z(n7937) );
  AND U13686 ( .A(b[19]), .B(a[87]), .Z(n7936) );
  XOR U13687 ( .A(n7941), .B(n7566), .Z(n7568) );
  XOR U13688 ( .A(n7942), .B(n7943), .Z(n7566) );
  AND U13689 ( .A(n7944), .B(n7945), .Z(n7942) );
  AND U13690 ( .A(b[17]), .B(a[89]), .Z(n7941) );
  XOR U13691 ( .A(n7946), .B(n7571), .Z(n7573) );
  XOR U13692 ( .A(n7947), .B(n7948), .Z(n7571) );
  AND U13693 ( .A(n7949), .B(n7950), .Z(n7947) );
  AND U13694 ( .A(b[16]), .B(a[90]), .Z(n7946) );
  XOR U13695 ( .A(n7951), .B(n7576), .Z(n7578) );
  XOR U13696 ( .A(n7952), .B(n7953), .Z(n7576) );
  AND U13697 ( .A(n7954), .B(n7955), .Z(n7952) );
  AND U13698 ( .A(b[15]), .B(a[91]), .Z(n7951) );
  XOR U13699 ( .A(n7956), .B(n7581), .Z(n7583) );
  XOR U13700 ( .A(n7957), .B(n7958), .Z(n7581) );
  AND U13701 ( .A(n7959), .B(n7960), .Z(n7957) );
  AND U13702 ( .A(b[14]), .B(a[92]), .Z(n7956) );
  XOR U13703 ( .A(n7961), .B(n7962), .Z(n7585) );
  AND U13704 ( .A(n7963), .B(n7964), .Z(n7961) );
  XOR U13705 ( .A(n7965), .B(n7590), .Z(n7592) );
  XOR U13706 ( .A(n7966), .B(n7967), .Z(n7590) );
  AND U13707 ( .A(n7968), .B(n7969), .Z(n7966) );
  AND U13708 ( .A(b[13]), .B(a[93]), .Z(n7965) );
  XOR U13709 ( .A(n7970), .B(n7595), .Z(n7597) );
  XOR U13710 ( .A(n7971), .B(n7972), .Z(n7595) );
  AND U13711 ( .A(n7973), .B(n7974), .Z(n7971) );
  AND U13712 ( .A(b[11]), .B(a[95]), .Z(n7970) );
  XOR U13713 ( .A(n7975), .B(n7600), .Z(n7602) );
  XOR U13714 ( .A(n7976), .B(n7977), .Z(n7600) );
  AND U13715 ( .A(n7978), .B(n7979), .Z(n7976) );
  AND U13716 ( .A(b[10]), .B(a[96]), .Z(n7975) );
  XOR U13717 ( .A(n7980), .B(n7605), .Z(n7607) );
  XOR U13718 ( .A(n7981), .B(n7982), .Z(n7605) );
  AND U13719 ( .A(n7983), .B(n7984), .Z(n7981) );
  AND U13720 ( .A(b[9]), .B(a[97]), .Z(n7980) );
  XOR U13721 ( .A(n7985), .B(n7610), .Z(n7612) );
  XOR U13722 ( .A(n7986), .B(n7987), .Z(n7610) );
  AND U13723 ( .A(n7988), .B(n7989), .Z(n7986) );
  AND U13724 ( .A(b[8]), .B(a[98]), .Z(n7985) );
  XOR U13725 ( .A(n7990), .B(n7991), .Z(n7614) );
  AND U13726 ( .A(n7992), .B(n7993), .Z(n7990) );
  XOR U13727 ( .A(n7994), .B(n7619), .Z(n7621) );
  XOR U13728 ( .A(n7995), .B(n7996), .Z(n7619) );
  AND U13729 ( .A(n7997), .B(n7998), .Z(n7995) );
  AND U13730 ( .A(b[7]), .B(a[99]), .Z(n7994) );
  XOR U13731 ( .A(n7999), .B(n7624), .Z(n7626) );
  XOR U13732 ( .A(n8000), .B(n8001), .Z(n7624) );
  AND U13733 ( .A(n8002), .B(n8003), .Z(n8000) );
  AND U13734 ( .A(b[5]), .B(a[101]), .Z(n7999) );
  XOR U13735 ( .A(n8004), .B(n7629), .Z(n7631) );
  XOR U13736 ( .A(n8005), .B(n8006), .Z(n7629) );
  AND U13737 ( .A(n8007), .B(n8008), .Z(n8005) );
  AND U13738 ( .A(b[4]), .B(a[102]), .Z(n8004) );
  XNOR U13739 ( .A(n8009), .B(n8010), .Z(n7643) );
  NANDN U13740 ( .A(n8011), .B(n8012), .Z(n8010) );
  XOR U13741 ( .A(n8013), .B(n7634), .Z(n7636) );
  XNOR U13742 ( .A(n8014), .B(n8015), .Z(n7634) );
  AND U13743 ( .A(n8016), .B(n8017), .Z(n8014) );
  AND U13744 ( .A(b[3]), .B(a[103]), .Z(n8013) );
  NAND U13745 ( .A(a[106]), .B(b[0]), .Z(n7281) );
  XOR U13746 ( .A(n8018), .B(n8019), .Z(swire[105]) );
  XOR U13747 ( .A(n7652), .B(n7653), .Z(n8020) );
  XNOR U13748 ( .A(n8011), .B(n8012), .Z(n7653) );
  XOR U13749 ( .A(n8009), .B(n8021), .Z(n8012) );
  NAND U13750 ( .A(b[1]), .B(a[104]), .Z(n8021) );
  XOR U13751 ( .A(n8017), .B(n8022), .Z(n8011) );
  XOR U13752 ( .A(n8009), .B(n8016), .Z(n8022) );
  XNOR U13753 ( .A(n8023), .B(n8015), .Z(n8016) );
  AND U13754 ( .A(b[2]), .B(a[103]), .Z(n8023) );
  NANDN U13755 ( .A(n8024), .B(n8025), .Z(n8009) );
  XOR U13756 ( .A(n8015), .B(n8007), .Z(n8026) );
  XNOR U13757 ( .A(n8006), .B(n8002), .Z(n8027) );
  XNOR U13758 ( .A(n7993), .B(n7992), .Z(n8028) );
  XOR U13759 ( .A(n8029), .B(n7991), .Z(n7992) );
  AND U13760 ( .A(b[5]), .B(a[100]), .Z(n8029) );
  XNOR U13761 ( .A(n7991), .B(n7997), .Z(n8030) );
  XNOR U13762 ( .A(n7996), .B(n7988), .Z(n8031) );
  XNOR U13763 ( .A(n7987), .B(n7983), .Z(n8032) );
  XNOR U13764 ( .A(n7982), .B(n7978), .Z(n8033) );
  XNOR U13765 ( .A(n7977), .B(n7973), .Z(n8034) );
  XNOR U13766 ( .A(n7964), .B(n7963), .Z(n8035) );
  XOR U13767 ( .A(n8036), .B(n7962), .Z(n7963) );
  AND U13768 ( .A(b[11]), .B(a[94]), .Z(n8036) );
  XNOR U13769 ( .A(n7962), .B(n7968), .Z(n8037) );
  XNOR U13770 ( .A(n7967), .B(n7959), .Z(n8038) );
  XNOR U13771 ( .A(n7958), .B(n7954), .Z(n8039) );
  XNOR U13772 ( .A(n7953), .B(n7949), .Z(n8040) );
  XNOR U13773 ( .A(n7948), .B(n7944), .Z(n8041) );
  XNOR U13774 ( .A(n7935), .B(n7934), .Z(n8042) );
  XOR U13775 ( .A(n8043), .B(n7933), .Z(n7934) );
  AND U13776 ( .A(b[17]), .B(a[88]), .Z(n8043) );
  XNOR U13777 ( .A(n7933), .B(n7939), .Z(n8044) );
  XNOR U13778 ( .A(n7938), .B(n7930), .Z(n8045) );
  XNOR U13779 ( .A(n7929), .B(n7925), .Z(n8046) );
  XNOR U13780 ( .A(n7924), .B(n7920), .Z(n8047) );
  XNOR U13781 ( .A(n7919), .B(n7915), .Z(n8048) );
  XNOR U13782 ( .A(n7906), .B(n7905), .Z(n8049) );
  XOR U13783 ( .A(n8050), .B(n7904), .Z(n7905) );
  AND U13784 ( .A(b[23]), .B(a[82]), .Z(n8050) );
  XNOR U13785 ( .A(n7904), .B(n7910), .Z(n8051) );
  XNOR U13786 ( .A(n7909), .B(n7901), .Z(n8052) );
  XNOR U13787 ( .A(n7900), .B(n7896), .Z(n8053) );
  XNOR U13788 ( .A(n7895), .B(n7891), .Z(n8054) );
  XNOR U13789 ( .A(n7890), .B(n7886), .Z(n8055) );
  XNOR U13790 ( .A(n7877), .B(n7876), .Z(n8056) );
  XOR U13791 ( .A(n8057), .B(n7875), .Z(n7876) );
  AND U13792 ( .A(b[29]), .B(a[76]), .Z(n8057) );
  XNOR U13793 ( .A(n7875), .B(n7881), .Z(n8058) );
  XNOR U13794 ( .A(n7880), .B(n7872), .Z(n8059) );
  XNOR U13795 ( .A(n7871), .B(n7867), .Z(n8060) );
  XNOR U13796 ( .A(n7866), .B(n7862), .Z(n8061) );
  XNOR U13797 ( .A(n7861), .B(n7857), .Z(n8062) );
  XNOR U13798 ( .A(n7848), .B(n7847), .Z(n8063) );
  XOR U13799 ( .A(n8064), .B(n7846), .Z(n7847) );
  AND U13800 ( .A(b[35]), .B(a[70]), .Z(n8064) );
  XNOR U13801 ( .A(n7846), .B(n7852), .Z(n8065) );
  XNOR U13802 ( .A(n7851), .B(n7843), .Z(n8066) );
  XNOR U13803 ( .A(n7842), .B(n7838), .Z(n8067) );
  XNOR U13804 ( .A(n7837), .B(n7833), .Z(n8068) );
  XNOR U13805 ( .A(n7832), .B(n7828), .Z(n8069) );
  XNOR U13806 ( .A(n7827), .B(n7823), .Z(n8070) );
  XNOR U13807 ( .A(n7822), .B(n7818), .Z(n8071) );
  XNOR U13808 ( .A(n7817), .B(n7813), .Z(n8072) );
  XNOR U13809 ( .A(n7812), .B(n7808), .Z(n8073) );
  XNOR U13810 ( .A(n7807), .B(n7803), .Z(n8074) );
  XNOR U13811 ( .A(n7802), .B(n7798), .Z(n8075) );
  XNOR U13812 ( .A(n7797), .B(n7793), .Z(n8076) );
  XNOR U13813 ( .A(n7792), .B(n7788), .Z(n8077) );
  XNOR U13814 ( .A(n7787), .B(n7783), .Z(n8078) );
  XNOR U13815 ( .A(n7782), .B(n7778), .Z(n8079) );
  XNOR U13816 ( .A(n7777), .B(n7773), .Z(n8080) );
  XNOR U13817 ( .A(n7772), .B(n7768), .Z(n8081) );
  XNOR U13818 ( .A(n7767), .B(n7763), .Z(n8082) );
  XNOR U13819 ( .A(n7762), .B(n7758), .Z(n8083) );
  XNOR U13820 ( .A(n7757), .B(n7753), .Z(n8084) );
  XNOR U13821 ( .A(n7752), .B(n7748), .Z(n8085) );
  XNOR U13822 ( .A(n7747), .B(n7743), .Z(n8086) );
  XNOR U13823 ( .A(n7742), .B(n7738), .Z(n8087) );
  XNOR U13824 ( .A(n7737), .B(n7733), .Z(n8088) );
  XOR U13825 ( .A(n7732), .B(n7729), .Z(n8089) );
  XOR U13826 ( .A(n8090), .B(n8091), .Z(n7729) );
  XOR U13827 ( .A(n7727), .B(n8092), .Z(n8091) );
  XOR U13828 ( .A(n8093), .B(n8094), .Z(n8092) );
  XOR U13829 ( .A(n8095), .B(n8096), .Z(n8094) );
  NAND U13830 ( .A(a[43]), .B(b[62]), .Z(n8096) );
  AND U13831 ( .A(a[42]), .B(b[63]), .Z(n8095) );
  XOR U13832 ( .A(n8097), .B(n8093), .Z(n8090) );
  XOR U13833 ( .A(n8098), .B(n8099), .Z(n8093) );
  ANDN U13834 ( .B(n8100), .A(n8101), .Z(n8098) );
  AND U13835 ( .A(a[44]), .B(b[61]), .Z(n8097) );
  XOR U13836 ( .A(n8102), .B(n7727), .Z(n7728) );
  XOR U13837 ( .A(n8103), .B(n8104), .Z(n7727) );
  AND U13838 ( .A(n8105), .B(n8106), .Z(n8103) );
  AND U13839 ( .A(a[45]), .B(b[60]), .Z(n8102) );
  XOR U13840 ( .A(n8107), .B(n7732), .Z(n7734) );
  XOR U13841 ( .A(n8108), .B(n8109), .Z(n7732) );
  AND U13842 ( .A(n8110), .B(n8111), .Z(n8108) );
  AND U13843 ( .A(a[46]), .B(b[59]), .Z(n8107) );
  XOR U13844 ( .A(n8112), .B(n7737), .Z(n7739) );
  XOR U13845 ( .A(n8113), .B(n8114), .Z(n7737) );
  AND U13846 ( .A(n8115), .B(n8116), .Z(n8113) );
  AND U13847 ( .A(a[47]), .B(b[58]), .Z(n8112) );
  XOR U13848 ( .A(n8117), .B(n7742), .Z(n7744) );
  XOR U13849 ( .A(n8118), .B(n8119), .Z(n7742) );
  AND U13850 ( .A(n8120), .B(n8121), .Z(n8118) );
  AND U13851 ( .A(a[48]), .B(b[57]), .Z(n8117) );
  XOR U13852 ( .A(n8122), .B(n7747), .Z(n7749) );
  XOR U13853 ( .A(n8123), .B(n8124), .Z(n7747) );
  AND U13854 ( .A(n8125), .B(n8126), .Z(n8123) );
  AND U13855 ( .A(a[49]), .B(b[56]), .Z(n8122) );
  XOR U13856 ( .A(n8127), .B(n7752), .Z(n7754) );
  XOR U13857 ( .A(n8128), .B(n8129), .Z(n7752) );
  AND U13858 ( .A(n8130), .B(n8131), .Z(n8128) );
  AND U13859 ( .A(a[50]), .B(b[55]), .Z(n8127) );
  XOR U13860 ( .A(n8132), .B(n7757), .Z(n7759) );
  XOR U13861 ( .A(n8133), .B(n8134), .Z(n7757) );
  AND U13862 ( .A(n8135), .B(n8136), .Z(n8133) );
  AND U13863 ( .A(a[51]), .B(b[54]), .Z(n8132) );
  XOR U13864 ( .A(n8137), .B(n7762), .Z(n7764) );
  XOR U13865 ( .A(n8138), .B(n8139), .Z(n7762) );
  AND U13866 ( .A(n8140), .B(n8141), .Z(n8138) );
  AND U13867 ( .A(a[52]), .B(b[53]), .Z(n8137) );
  XOR U13868 ( .A(n8142), .B(n7767), .Z(n7769) );
  XOR U13869 ( .A(n8143), .B(n8144), .Z(n7767) );
  AND U13870 ( .A(n8145), .B(n8146), .Z(n8143) );
  AND U13871 ( .A(b[52]), .B(a[53]), .Z(n8142) );
  XOR U13872 ( .A(n8147), .B(n7772), .Z(n7774) );
  XOR U13873 ( .A(n8148), .B(n8149), .Z(n7772) );
  AND U13874 ( .A(n8150), .B(n8151), .Z(n8148) );
  AND U13875 ( .A(b[51]), .B(a[54]), .Z(n8147) );
  XOR U13876 ( .A(n8152), .B(n7777), .Z(n7779) );
  XOR U13877 ( .A(n8153), .B(n8154), .Z(n7777) );
  AND U13878 ( .A(n8155), .B(n8156), .Z(n8153) );
  AND U13879 ( .A(b[50]), .B(a[55]), .Z(n8152) );
  XOR U13880 ( .A(n8157), .B(n7782), .Z(n7784) );
  XOR U13881 ( .A(n8158), .B(n8159), .Z(n7782) );
  AND U13882 ( .A(n8160), .B(n8161), .Z(n8158) );
  AND U13883 ( .A(b[49]), .B(a[56]), .Z(n8157) );
  XOR U13884 ( .A(n8162), .B(n7787), .Z(n7789) );
  XOR U13885 ( .A(n8163), .B(n8164), .Z(n7787) );
  AND U13886 ( .A(n8165), .B(n8166), .Z(n8163) );
  AND U13887 ( .A(b[48]), .B(a[57]), .Z(n8162) );
  XOR U13888 ( .A(n8167), .B(n7792), .Z(n7794) );
  XOR U13889 ( .A(n8168), .B(n8169), .Z(n7792) );
  AND U13890 ( .A(n8170), .B(n8171), .Z(n8168) );
  AND U13891 ( .A(b[47]), .B(a[58]), .Z(n8167) );
  XOR U13892 ( .A(n8172), .B(n7797), .Z(n7799) );
  XOR U13893 ( .A(n8173), .B(n8174), .Z(n7797) );
  AND U13894 ( .A(n8175), .B(n8176), .Z(n8173) );
  AND U13895 ( .A(b[46]), .B(a[59]), .Z(n8172) );
  XOR U13896 ( .A(n8177), .B(n7802), .Z(n7804) );
  XOR U13897 ( .A(n8178), .B(n8179), .Z(n7802) );
  AND U13898 ( .A(n8180), .B(n8181), .Z(n8178) );
  AND U13899 ( .A(b[45]), .B(a[60]), .Z(n8177) );
  XOR U13900 ( .A(n8182), .B(n7807), .Z(n7809) );
  XOR U13901 ( .A(n8183), .B(n8184), .Z(n7807) );
  AND U13902 ( .A(n8185), .B(n8186), .Z(n8183) );
  AND U13903 ( .A(b[44]), .B(a[61]), .Z(n8182) );
  XOR U13904 ( .A(n8187), .B(n7812), .Z(n7814) );
  XOR U13905 ( .A(n8188), .B(n8189), .Z(n7812) );
  AND U13906 ( .A(n8190), .B(n8191), .Z(n8188) );
  AND U13907 ( .A(b[43]), .B(a[62]), .Z(n8187) );
  XOR U13908 ( .A(n8192), .B(n7817), .Z(n7819) );
  XOR U13909 ( .A(n8193), .B(n8194), .Z(n7817) );
  AND U13910 ( .A(n8195), .B(n8196), .Z(n8193) );
  AND U13911 ( .A(b[42]), .B(a[63]), .Z(n8192) );
  XOR U13912 ( .A(n8197), .B(n7822), .Z(n7824) );
  XOR U13913 ( .A(n8198), .B(n8199), .Z(n7822) );
  AND U13914 ( .A(n8200), .B(n8201), .Z(n8198) );
  AND U13915 ( .A(b[41]), .B(a[64]), .Z(n8197) );
  XOR U13916 ( .A(n8202), .B(n7827), .Z(n7829) );
  XOR U13917 ( .A(n8203), .B(n8204), .Z(n7827) );
  AND U13918 ( .A(n8205), .B(n8206), .Z(n8203) );
  AND U13919 ( .A(b[40]), .B(a[65]), .Z(n8202) );
  XOR U13920 ( .A(n8207), .B(n7832), .Z(n7834) );
  XOR U13921 ( .A(n8208), .B(n8209), .Z(n7832) );
  AND U13922 ( .A(n8210), .B(n8211), .Z(n8208) );
  AND U13923 ( .A(b[39]), .B(a[66]), .Z(n8207) );
  XOR U13924 ( .A(n8212), .B(n7837), .Z(n7839) );
  XOR U13925 ( .A(n8213), .B(n8214), .Z(n7837) );
  AND U13926 ( .A(n8215), .B(n8216), .Z(n8213) );
  AND U13927 ( .A(b[38]), .B(a[67]), .Z(n8212) );
  XOR U13928 ( .A(n8217), .B(n7842), .Z(n7844) );
  XOR U13929 ( .A(n8218), .B(n8219), .Z(n7842) );
  AND U13930 ( .A(n8220), .B(n8221), .Z(n8218) );
  AND U13931 ( .A(b[37]), .B(a[68]), .Z(n8217) );
  XOR U13932 ( .A(n8222), .B(n8223), .Z(n7846) );
  AND U13933 ( .A(n8224), .B(n8225), .Z(n8222) );
  XOR U13934 ( .A(n8226), .B(n7851), .Z(n7853) );
  XOR U13935 ( .A(n8227), .B(n8228), .Z(n7851) );
  AND U13936 ( .A(n8229), .B(n8230), .Z(n8227) );
  AND U13937 ( .A(b[36]), .B(a[69]), .Z(n8226) );
  XOR U13938 ( .A(n8231), .B(n7856), .Z(n7858) );
  XOR U13939 ( .A(n8232), .B(n8233), .Z(n7856) );
  AND U13940 ( .A(n8234), .B(n8235), .Z(n8232) );
  AND U13941 ( .A(b[34]), .B(a[71]), .Z(n8231) );
  XOR U13942 ( .A(n8236), .B(n7861), .Z(n7863) );
  XOR U13943 ( .A(n8237), .B(n8238), .Z(n7861) );
  AND U13944 ( .A(n8239), .B(n8240), .Z(n8237) );
  AND U13945 ( .A(b[33]), .B(a[72]), .Z(n8236) );
  XOR U13946 ( .A(n8241), .B(n7866), .Z(n7868) );
  XOR U13947 ( .A(n8242), .B(n8243), .Z(n7866) );
  AND U13948 ( .A(n8244), .B(n8245), .Z(n8242) );
  AND U13949 ( .A(b[32]), .B(a[73]), .Z(n8241) );
  XOR U13950 ( .A(n8246), .B(n7871), .Z(n7873) );
  XOR U13951 ( .A(n8247), .B(n8248), .Z(n7871) );
  AND U13952 ( .A(n8249), .B(n8250), .Z(n8247) );
  AND U13953 ( .A(b[31]), .B(a[74]), .Z(n8246) );
  XOR U13954 ( .A(n8251), .B(n8252), .Z(n7875) );
  AND U13955 ( .A(n8253), .B(n8254), .Z(n8251) );
  XOR U13956 ( .A(n8255), .B(n7880), .Z(n7882) );
  XOR U13957 ( .A(n8256), .B(n8257), .Z(n7880) );
  AND U13958 ( .A(n8258), .B(n8259), .Z(n8256) );
  AND U13959 ( .A(b[30]), .B(a[75]), .Z(n8255) );
  XOR U13960 ( .A(n8260), .B(n7885), .Z(n7887) );
  XOR U13961 ( .A(n8261), .B(n8262), .Z(n7885) );
  AND U13962 ( .A(n8263), .B(n8264), .Z(n8261) );
  AND U13963 ( .A(b[28]), .B(a[77]), .Z(n8260) );
  XOR U13964 ( .A(n8265), .B(n7890), .Z(n7892) );
  XOR U13965 ( .A(n8266), .B(n8267), .Z(n7890) );
  AND U13966 ( .A(n8268), .B(n8269), .Z(n8266) );
  AND U13967 ( .A(b[27]), .B(a[78]), .Z(n8265) );
  XOR U13968 ( .A(n8270), .B(n7895), .Z(n7897) );
  XOR U13969 ( .A(n8271), .B(n8272), .Z(n7895) );
  AND U13970 ( .A(n8273), .B(n8274), .Z(n8271) );
  AND U13971 ( .A(b[26]), .B(a[79]), .Z(n8270) );
  XOR U13972 ( .A(n8275), .B(n7900), .Z(n7902) );
  XOR U13973 ( .A(n8276), .B(n8277), .Z(n7900) );
  AND U13974 ( .A(n8278), .B(n8279), .Z(n8276) );
  AND U13975 ( .A(b[25]), .B(a[80]), .Z(n8275) );
  XOR U13976 ( .A(n8280), .B(n8281), .Z(n7904) );
  AND U13977 ( .A(n8282), .B(n8283), .Z(n8280) );
  XOR U13978 ( .A(n8284), .B(n7909), .Z(n7911) );
  XOR U13979 ( .A(n8285), .B(n8286), .Z(n7909) );
  AND U13980 ( .A(n8287), .B(n8288), .Z(n8285) );
  AND U13981 ( .A(b[24]), .B(a[81]), .Z(n8284) );
  XOR U13982 ( .A(n8289), .B(n7914), .Z(n7916) );
  XOR U13983 ( .A(n8290), .B(n8291), .Z(n7914) );
  AND U13984 ( .A(n8292), .B(n8293), .Z(n8290) );
  AND U13985 ( .A(b[22]), .B(a[83]), .Z(n8289) );
  XOR U13986 ( .A(n8294), .B(n7919), .Z(n7921) );
  XOR U13987 ( .A(n8295), .B(n8296), .Z(n7919) );
  AND U13988 ( .A(n8297), .B(n8298), .Z(n8295) );
  AND U13989 ( .A(b[21]), .B(a[84]), .Z(n8294) );
  XOR U13990 ( .A(n8299), .B(n7924), .Z(n7926) );
  XOR U13991 ( .A(n8300), .B(n8301), .Z(n7924) );
  AND U13992 ( .A(n8302), .B(n8303), .Z(n8300) );
  AND U13993 ( .A(b[20]), .B(a[85]), .Z(n8299) );
  XOR U13994 ( .A(n8304), .B(n7929), .Z(n7931) );
  XOR U13995 ( .A(n8305), .B(n8306), .Z(n7929) );
  AND U13996 ( .A(n8307), .B(n8308), .Z(n8305) );
  AND U13997 ( .A(b[19]), .B(a[86]), .Z(n8304) );
  XOR U13998 ( .A(n8309), .B(n8310), .Z(n7933) );
  AND U13999 ( .A(n8311), .B(n8312), .Z(n8309) );
  XOR U14000 ( .A(n8313), .B(n7938), .Z(n7940) );
  XOR U14001 ( .A(n8314), .B(n8315), .Z(n7938) );
  AND U14002 ( .A(n8316), .B(n8317), .Z(n8314) );
  AND U14003 ( .A(b[18]), .B(a[87]), .Z(n8313) );
  XOR U14004 ( .A(n8318), .B(n7943), .Z(n7945) );
  XOR U14005 ( .A(n8319), .B(n8320), .Z(n7943) );
  AND U14006 ( .A(n8321), .B(n8322), .Z(n8319) );
  AND U14007 ( .A(b[16]), .B(a[89]), .Z(n8318) );
  XOR U14008 ( .A(n8323), .B(n7948), .Z(n7950) );
  XOR U14009 ( .A(n8324), .B(n8325), .Z(n7948) );
  AND U14010 ( .A(n8326), .B(n8327), .Z(n8324) );
  AND U14011 ( .A(b[15]), .B(a[90]), .Z(n8323) );
  XOR U14012 ( .A(n8328), .B(n7953), .Z(n7955) );
  XOR U14013 ( .A(n8329), .B(n8330), .Z(n7953) );
  AND U14014 ( .A(n8331), .B(n8332), .Z(n8329) );
  AND U14015 ( .A(b[14]), .B(a[91]), .Z(n8328) );
  XOR U14016 ( .A(n8333), .B(n7958), .Z(n7960) );
  XOR U14017 ( .A(n8334), .B(n8335), .Z(n7958) );
  AND U14018 ( .A(n8336), .B(n8337), .Z(n8334) );
  AND U14019 ( .A(b[13]), .B(a[92]), .Z(n8333) );
  XOR U14020 ( .A(n8338), .B(n8339), .Z(n7962) );
  AND U14021 ( .A(n8340), .B(n8341), .Z(n8338) );
  XOR U14022 ( .A(n8342), .B(n7967), .Z(n7969) );
  XOR U14023 ( .A(n8343), .B(n8344), .Z(n7967) );
  AND U14024 ( .A(n8345), .B(n8346), .Z(n8343) );
  AND U14025 ( .A(b[12]), .B(a[93]), .Z(n8342) );
  XOR U14026 ( .A(n8347), .B(n7972), .Z(n7974) );
  XOR U14027 ( .A(n8348), .B(n8349), .Z(n7972) );
  AND U14028 ( .A(n8350), .B(n8351), .Z(n8348) );
  AND U14029 ( .A(b[10]), .B(a[95]), .Z(n8347) );
  XOR U14030 ( .A(n8352), .B(n7977), .Z(n7979) );
  XOR U14031 ( .A(n8353), .B(n8354), .Z(n7977) );
  AND U14032 ( .A(n8355), .B(n8356), .Z(n8353) );
  AND U14033 ( .A(b[9]), .B(a[96]), .Z(n8352) );
  XOR U14034 ( .A(n8357), .B(n7982), .Z(n7984) );
  XOR U14035 ( .A(n8358), .B(n8359), .Z(n7982) );
  AND U14036 ( .A(n8360), .B(n8361), .Z(n8358) );
  AND U14037 ( .A(b[8]), .B(a[97]), .Z(n8357) );
  XOR U14038 ( .A(n8362), .B(n7987), .Z(n7989) );
  XOR U14039 ( .A(n8363), .B(n8364), .Z(n7987) );
  AND U14040 ( .A(n8365), .B(n8366), .Z(n8363) );
  AND U14041 ( .A(b[7]), .B(a[98]), .Z(n8362) );
  XOR U14042 ( .A(n8367), .B(n8368), .Z(n7991) );
  AND U14043 ( .A(n8369), .B(n8370), .Z(n8367) );
  XOR U14044 ( .A(n8371), .B(n7996), .Z(n7998) );
  XOR U14045 ( .A(n8372), .B(n8373), .Z(n7996) );
  AND U14046 ( .A(n8374), .B(n8375), .Z(n8372) );
  AND U14047 ( .A(b[6]), .B(a[99]), .Z(n8371) );
  XOR U14048 ( .A(n8376), .B(n8001), .Z(n8003) );
  XOR U14049 ( .A(n8377), .B(n8378), .Z(n8001) );
  AND U14050 ( .A(n8379), .B(n8380), .Z(n8377) );
  AND U14051 ( .A(b[4]), .B(a[101]), .Z(n8376) );
  XNOR U14052 ( .A(n8381), .B(n8382), .Z(n8015) );
  NANDN U14053 ( .A(n8383), .B(n8384), .Z(n8382) );
  XOR U14054 ( .A(n8385), .B(n8006), .Z(n8008) );
  XNOR U14055 ( .A(n8386), .B(n8387), .Z(n8006) );
  AND U14056 ( .A(n8388), .B(n8389), .Z(n8386) );
  AND U14057 ( .A(b[3]), .B(a[102]), .Z(n8385) );
  NAND U14058 ( .A(a[105]), .B(b[0]), .Z(n7652) );
  XOR U14059 ( .A(n8390), .B(n8391), .Z(swire[104]) );
  XOR U14060 ( .A(n8024), .B(n8025), .Z(n8392) );
  XNOR U14061 ( .A(n8383), .B(n8384), .Z(n8025) );
  XOR U14062 ( .A(n8381), .B(n8393), .Z(n8384) );
  NAND U14063 ( .A(b[1]), .B(a[103]), .Z(n8393) );
  XOR U14064 ( .A(n8389), .B(n8394), .Z(n8383) );
  XOR U14065 ( .A(n8381), .B(n8388), .Z(n8394) );
  XNOR U14066 ( .A(n8395), .B(n8387), .Z(n8388) );
  AND U14067 ( .A(b[2]), .B(a[102]), .Z(n8395) );
  NANDN U14068 ( .A(n8396), .B(n8397), .Z(n8381) );
  XOR U14069 ( .A(n8387), .B(n8379), .Z(n8398) );
  XNOR U14070 ( .A(n8370), .B(n8369), .Z(n8399) );
  XOR U14071 ( .A(n8400), .B(n8368), .Z(n8369) );
  AND U14072 ( .A(b[4]), .B(a[100]), .Z(n8400) );
  XNOR U14073 ( .A(n8368), .B(n8374), .Z(n8401) );
  XNOR U14074 ( .A(n8373), .B(n8365), .Z(n8402) );
  XNOR U14075 ( .A(n8364), .B(n8360), .Z(n8403) );
  XNOR U14076 ( .A(n8359), .B(n8355), .Z(n8404) );
  XNOR U14077 ( .A(n8354), .B(n8350), .Z(n8405) );
  XNOR U14078 ( .A(n8341), .B(n8340), .Z(n8406) );
  XOR U14079 ( .A(n8407), .B(n8339), .Z(n8340) );
  AND U14080 ( .A(b[10]), .B(a[94]), .Z(n8407) );
  XNOR U14081 ( .A(n8339), .B(n8345), .Z(n8408) );
  XNOR U14082 ( .A(n8344), .B(n8336), .Z(n8409) );
  XNOR U14083 ( .A(n8335), .B(n8331), .Z(n8410) );
  XNOR U14084 ( .A(n8330), .B(n8326), .Z(n8411) );
  XNOR U14085 ( .A(n8325), .B(n8321), .Z(n8412) );
  XNOR U14086 ( .A(n8312), .B(n8311), .Z(n8413) );
  XOR U14087 ( .A(n8414), .B(n8310), .Z(n8311) );
  AND U14088 ( .A(b[16]), .B(a[88]), .Z(n8414) );
  XNOR U14089 ( .A(n8310), .B(n8316), .Z(n8415) );
  XNOR U14090 ( .A(n8315), .B(n8307), .Z(n8416) );
  XNOR U14091 ( .A(n8306), .B(n8302), .Z(n8417) );
  XNOR U14092 ( .A(n8301), .B(n8297), .Z(n8418) );
  XNOR U14093 ( .A(n8296), .B(n8292), .Z(n8419) );
  XNOR U14094 ( .A(n8283), .B(n8282), .Z(n8420) );
  XOR U14095 ( .A(n8421), .B(n8281), .Z(n8282) );
  AND U14096 ( .A(b[22]), .B(a[82]), .Z(n8421) );
  XNOR U14097 ( .A(n8281), .B(n8287), .Z(n8422) );
  XNOR U14098 ( .A(n8286), .B(n8278), .Z(n8423) );
  XNOR U14099 ( .A(n8277), .B(n8273), .Z(n8424) );
  XNOR U14100 ( .A(n8272), .B(n8268), .Z(n8425) );
  XNOR U14101 ( .A(n8267), .B(n8263), .Z(n8426) );
  XNOR U14102 ( .A(n8254), .B(n8253), .Z(n8427) );
  XOR U14103 ( .A(n8428), .B(n8252), .Z(n8253) );
  AND U14104 ( .A(b[28]), .B(a[76]), .Z(n8428) );
  XNOR U14105 ( .A(n8252), .B(n8258), .Z(n8429) );
  XNOR U14106 ( .A(n8257), .B(n8249), .Z(n8430) );
  XNOR U14107 ( .A(n8248), .B(n8244), .Z(n8431) );
  XNOR U14108 ( .A(n8243), .B(n8239), .Z(n8432) );
  XNOR U14109 ( .A(n8238), .B(n8234), .Z(n8433) );
  XNOR U14110 ( .A(n8225), .B(n8224), .Z(n8434) );
  XOR U14111 ( .A(n8435), .B(n8223), .Z(n8224) );
  AND U14112 ( .A(b[34]), .B(a[70]), .Z(n8435) );
  XNOR U14113 ( .A(n8223), .B(n8229), .Z(n8436) );
  XNOR U14114 ( .A(n8228), .B(n8220), .Z(n8437) );
  XNOR U14115 ( .A(n8219), .B(n8215), .Z(n8438) );
  XNOR U14116 ( .A(n8214), .B(n8210), .Z(n8439) );
  XNOR U14117 ( .A(n8209), .B(n8205), .Z(n8440) );
  XNOR U14118 ( .A(n8204), .B(n8200), .Z(n8441) );
  XNOR U14119 ( .A(n8199), .B(n8195), .Z(n8442) );
  XNOR U14120 ( .A(n8194), .B(n8190), .Z(n8443) );
  XNOR U14121 ( .A(n8189), .B(n8185), .Z(n8444) );
  XNOR U14122 ( .A(n8184), .B(n8180), .Z(n8445) );
  XNOR U14123 ( .A(n8179), .B(n8175), .Z(n8446) );
  XNOR U14124 ( .A(n8174), .B(n8170), .Z(n8447) );
  XNOR U14125 ( .A(n8169), .B(n8165), .Z(n8448) );
  XNOR U14126 ( .A(n8164), .B(n8160), .Z(n8449) );
  XNOR U14127 ( .A(n8159), .B(n8155), .Z(n8450) );
  XNOR U14128 ( .A(n8154), .B(n8150), .Z(n8451) );
  XNOR U14129 ( .A(n8149), .B(n8145), .Z(n8452) );
  XNOR U14130 ( .A(n8144), .B(n8140), .Z(n8453) );
  XNOR U14131 ( .A(n8139), .B(n8135), .Z(n8454) );
  XNOR U14132 ( .A(n8134), .B(n8130), .Z(n8455) );
  XNOR U14133 ( .A(n8129), .B(n8125), .Z(n8456) );
  XNOR U14134 ( .A(n8124), .B(n8120), .Z(n8457) );
  XNOR U14135 ( .A(n8119), .B(n8115), .Z(n8458) );
  XNOR U14136 ( .A(n8114), .B(n8110), .Z(n8459) );
  XNOR U14137 ( .A(n8109), .B(n8105), .Z(n8460) );
  XOR U14138 ( .A(n8104), .B(n8101), .Z(n8461) );
  XOR U14139 ( .A(n8462), .B(n8463), .Z(n8101) );
  XOR U14140 ( .A(n8099), .B(n8464), .Z(n8463) );
  XOR U14141 ( .A(n8465), .B(n8466), .Z(n8464) );
  XOR U14142 ( .A(n8467), .B(n8468), .Z(n8466) );
  NAND U14143 ( .A(a[42]), .B(b[62]), .Z(n8468) );
  AND U14144 ( .A(a[41]), .B(b[63]), .Z(n8467) );
  XOR U14145 ( .A(n8469), .B(n8465), .Z(n8462) );
  XOR U14146 ( .A(n8470), .B(n8471), .Z(n8465) );
  ANDN U14147 ( .B(n8472), .A(n8473), .Z(n8470) );
  AND U14148 ( .A(a[43]), .B(b[61]), .Z(n8469) );
  XOR U14149 ( .A(n8474), .B(n8099), .Z(n8100) );
  XOR U14150 ( .A(n8475), .B(n8476), .Z(n8099) );
  AND U14151 ( .A(n8477), .B(n8478), .Z(n8475) );
  AND U14152 ( .A(a[44]), .B(b[60]), .Z(n8474) );
  XOR U14153 ( .A(n8479), .B(n8104), .Z(n8106) );
  XOR U14154 ( .A(n8480), .B(n8481), .Z(n8104) );
  AND U14155 ( .A(n8482), .B(n8483), .Z(n8480) );
  AND U14156 ( .A(a[45]), .B(b[59]), .Z(n8479) );
  XOR U14157 ( .A(n8484), .B(n8109), .Z(n8111) );
  XOR U14158 ( .A(n8485), .B(n8486), .Z(n8109) );
  AND U14159 ( .A(n8487), .B(n8488), .Z(n8485) );
  AND U14160 ( .A(a[46]), .B(b[58]), .Z(n8484) );
  XOR U14161 ( .A(n8489), .B(n8114), .Z(n8116) );
  XOR U14162 ( .A(n8490), .B(n8491), .Z(n8114) );
  AND U14163 ( .A(n8492), .B(n8493), .Z(n8490) );
  AND U14164 ( .A(a[47]), .B(b[57]), .Z(n8489) );
  XOR U14165 ( .A(n8494), .B(n8119), .Z(n8121) );
  XOR U14166 ( .A(n8495), .B(n8496), .Z(n8119) );
  AND U14167 ( .A(n8497), .B(n8498), .Z(n8495) );
  AND U14168 ( .A(a[48]), .B(b[56]), .Z(n8494) );
  XOR U14169 ( .A(n8499), .B(n8124), .Z(n8126) );
  XOR U14170 ( .A(n8500), .B(n8501), .Z(n8124) );
  AND U14171 ( .A(n8502), .B(n8503), .Z(n8500) );
  AND U14172 ( .A(a[49]), .B(b[55]), .Z(n8499) );
  XOR U14173 ( .A(n8504), .B(n8129), .Z(n8131) );
  XOR U14174 ( .A(n8505), .B(n8506), .Z(n8129) );
  AND U14175 ( .A(n8507), .B(n8508), .Z(n8505) );
  AND U14176 ( .A(a[50]), .B(b[54]), .Z(n8504) );
  XOR U14177 ( .A(n8509), .B(n8134), .Z(n8136) );
  XOR U14178 ( .A(n8510), .B(n8511), .Z(n8134) );
  AND U14179 ( .A(n8512), .B(n8513), .Z(n8510) );
  AND U14180 ( .A(a[51]), .B(b[53]), .Z(n8509) );
  XOR U14181 ( .A(n8514), .B(n8139), .Z(n8141) );
  XOR U14182 ( .A(n8515), .B(n8516), .Z(n8139) );
  AND U14183 ( .A(n8517), .B(n8518), .Z(n8515) );
  AND U14184 ( .A(a[52]), .B(b[52]), .Z(n8514) );
  XOR U14185 ( .A(n8519), .B(n8144), .Z(n8146) );
  XOR U14186 ( .A(n8520), .B(n8521), .Z(n8144) );
  AND U14187 ( .A(n8522), .B(n8523), .Z(n8520) );
  AND U14188 ( .A(b[51]), .B(a[53]), .Z(n8519) );
  XOR U14189 ( .A(n8524), .B(n8149), .Z(n8151) );
  XOR U14190 ( .A(n8525), .B(n8526), .Z(n8149) );
  AND U14191 ( .A(n8527), .B(n8528), .Z(n8525) );
  AND U14192 ( .A(b[50]), .B(a[54]), .Z(n8524) );
  XOR U14193 ( .A(n8529), .B(n8154), .Z(n8156) );
  XOR U14194 ( .A(n8530), .B(n8531), .Z(n8154) );
  AND U14195 ( .A(n8532), .B(n8533), .Z(n8530) );
  AND U14196 ( .A(b[49]), .B(a[55]), .Z(n8529) );
  XOR U14197 ( .A(n8534), .B(n8159), .Z(n8161) );
  XOR U14198 ( .A(n8535), .B(n8536), .Z(n8159) );
  AND U14199 ( .A(n8537), .B(n8538), .Z(n8535) );
  AND U14200 ( .A(b[48]), .B(a[56]), .Z(n8534) );
  XOR U14201 ( .A(n8539), .B(n8164), .Z(n8166) );
  XOR U14202 ( .A(n8540), .B(n8541), .Z(n8164) );
  AND U14203 ( .A(n8542), .B(n8543), .Z(n8540) );
  AND U14204 ( .A(b[47]), .B(a[57]), .Z(n8539) );
  XOR U14205 ( .A(n8544), .B(n8169), .Z(n8171) );
  XOR U14206 ( .A(n8545), .B(n8546), .Z(n8169) );
  AND U14207 ( .A(n8547), .B(n8548), .Z(n8545) );
  AND U14208 ( .A(b[46]), .B(a[58]), .Z(n8544) );
  XOR U14209 ( .A(n8549), .B(n8174), .Z(n8176) );
  XOR U14210 ( .A(n8550), .B(n8551), .Z(n8174) );
  AND U14211 ( .A(n8552), .B(n8553), .Z(n8550) );
  AND U14212 ( .A(b[45]), .B(a[59]), .Z(n8549) );
  XOR U14213 ( .A(n8554), .B(n8179), .Z(n8181) );
  XOR U14214 ( .A(n8555), .B(n8556), .Z(n8179) );
  AND U14215 ( .A(n8557), .B(n8558), .Z(n8555) );
  AND U14216 ( .A(b[44]), .B(a[60]), .Z(n8554) );
  XOR U14217 ( .A(n8559), .B(n8184), .Z(n8186) );
  XOR U14218 ( .A(n8560), .B(n8561), .Z(n8184) );
  AND U14219 ( .A(n8562), .B(n8563), .Z(n8560) );
  AND U14220 ( .A(b[43]), .B(a[61]), .Z(n8559) );
  XOR U14221 ( .A(n8564), .B(n8189), .Z(n8191) );
  XOR U14222 ( .A(n8565), .B(n8566), .Z(n8189) );
  AND U14223 ( .A(n8567), .B(n8568), .Z(n8565) );
  AND U14224 ( .A(b[42]), .B(a[62]), .Z(n8564) );
  XOR U14225 ( .A(n8569), .B(n8194), .Z(n8196) );
  XOR U14226 ( .A(n8570), .B(n8571), .Z(n8194) );
  AND U14227 ( .A(n8572), .B(n8573), .Z(n8570) );
  AND U14228 ( .A(b[41]), .B(a[63]), .Z(n8569) );
  XOR U14229 ( .A(n8574), .B(n8199), .Z(n8201) );
  XOR U14230 ( .A(n8575), .B(n8576), .Z(n8199) );
  AND U14231 ( .A(n8577), .B(n8578), .Z(n8575) );
  AND U14232 ( .A(b[40]), .B(a[64]), .Z(n8574) );
  XOR U14233 ( .A(n8579), .B(n8204), .Z(n8206) );
  XOR U14234 ( .A(n8580), .B(n8581), .Z(n8204) );
  AND U14235 ( .A(n8582), .B(n8583), .Z(n8580) );
  AND U14236 ( .A(b[39]), .B(a[65]), .Z(n8579) );
  XOR U14237 ( .A(n8584), .B(n8209), .Z(n8211) );
  XOR U14238 ( .A(n8585), .B(n8586), .Z(n8209) );
  AND U14239 ( .A(n8587), .B(n8588), .Z(n8585) );
  AND U14240 ( .A(b[38]), .B(a[66]), .Z(n8584) );
  XOR U14241 ( .A(n8589), .B(n8214), .Z(n8216) );
  XOR U14242 ( .A(n8590), .B(n8591), .Z(n8214) );
  AND U14243 ( .A(n8592), .B(n8593), .Z(n8590) );
  AND U14244 ( .A(b[37]), .B(a[67]), .Z(n8589) );
  XOR U14245 ( .A(n8594), .B(n8219), .Z(n8221) );
  XOR U14246 ( .A(n8595), .B(n8596), .Z(n8219) );
  AND U14247 ( .A(n8597), .B(n8598), .Z(n8595) );
  AND U14248 ( .A(b[36]), .B(a[68]), .Z(n8594) );
  XOR U14249 ( .A(n8599), .B(n8600), .Z(n8223) );
  AND U14250 ( .A(n8601), .B(n8602), .Z(n8599) );
  XOR U14251 ( .A(n8603), .B(n8228), .Z(n8230) );
  XOR U14252 ( .A(n8604), .B(n8605), .Z(n8228) );
  AND U14253 ( .A(n8606), .B(n8607), .Z(n8604) );
  AND U14254 ( .A(b[35]), .B(a[69]), .Z(n8603) );
  XOR U14255 ( .A(n8608), .B(n8233), .Z(n8235) );
  XOR U14256 ( .A(n8609), .B(n8610), .Z(n8233) );
  AND U14257 ( .A(n8611), .B(n8612), .Z(n8609) );
  AND U14258 ( .A(b[33]), .B(a[71]), .Z(n8608) );
  XOR U14259 ( .A(n8613), .B(n8238), .Z(n8240) );
  XOR U14260 ( .A(n8614), .B(n8615), .Z(n8238) );
  AND U14261 ( .A(n8616), .B(n8617), .Z(n8614) );
  AND U14262 ( .A(b[32]), .B(a[72]), .Z(n8613) );
  XOR U14263 ( .A(n8618), .B(n8243), .Z(n8245) );
  XOR U14264 ( .A(n8619), .B(n8620), .Z(n8243) );
  AND U14265 ( .A(n8621), .B(n8622), .Z(n8619) );
  AND U14266 ( .A(b[31]), .B(a[73]), .Z(n8618) );
  XOR U14267 ( .A(n8623), .B(n8248), .Z(n8250) );
  XOR U14268 ( .A(n8624), .B(n8625), .Z(n8248) );
  AND U14269 ( .A(n8626), .B(n8627), .Z(n8624) );
  AND U14270 ( .A(b[30]), .B(a[74]), .Z(n8623) );
  XOR U14271 ( .A(n8628), .B(n8629), .Z(n8252) );
  AND U14272 ( .A(n8630), .B(n8631), .Z(n8628) );
  XOR U14273 ( .A(n8632), .B(n8257), .Z(n8259) );
  XOR U14274 ( .A(n8633), .B(n8634), .Z(n8257) );
  AND U14275 ( .A(n8635), .B(n8636), .Z(n8633) );
  AND U14276 ( .A(b[29]), .B(a[75]), .Z(n8632) );
  XOR U14277 ( .A(n8637), .B(n8262), .Z(n8264) );
  XOR U14278 ( .A(n8638), .B(n8639), .Z(n8262) );
  AND U14279 ( .A(n8640), .B(n8641), .Z(n8638) );
  AND U14280 ( .A(b[27]), .B(a[77]), .Z(n8637) );
  XOR U14281 ( .A(n8642), .B(n8267), .Z(n8269) );
  XOR U14282 ( .A(n8643), .B(n8644), .Z(n8267) );
  AND U14283 ( .A(n8645), .B(n8646), .Z(n8643) );
  AND U14284 ( .A(b[26]), .B(a[78]), .Z(n8642) );
  XOR U14285 ( .A(n8647), .B(n8272), .Z(n8274) );
  XOR U14286 ( .A(n8648), .B(n8649), .Z(n8272) );
  AND U14287 ( .A(n8650), .B(n8651), .Z(n8648) );
  AND U14288 ( .A(b[25]), .B(a[79]), .Z(n8647) );
  XOR U14289 ( .A(n8652), .B(n8277), .Z(n8279) );
  XOR U14290 ( .A(n8653), .B(n8654), .Z(n8277) );
  AND U14291 ( .A(n8655), .B(n8656), .Z(n8653) );
  AND U14292 ( .A(b[24]), .B(a[80]), .Z(n8652) );
  XOR U14293 ( .A(n8657), .B(n8658), .Z(n8281) );
  AND U14294 ( .A(n8659), .B(n8660), .Z(n8657) );
  XOR U14295 ( .A(n8661), .B(n8286), .Z(n8288) );
  XOR U14296 ( .A(n8662), .B(n8663), .Z(n8286) );
  AND U14297 ( .A(n8664), .B(n8665), .Z(n8662) );
  AND U14298 ( .A(b[23]), .B(a[81]), .Z(n8661) );
  XOR U14299 ( .A(n8666), .B(n8291), .Z(n8293) );
  XOR U14300 ( .A(n8667), .B(n8668), .Z(n8291) );
  AND U14301 ( .A(n8669), .B(n8670), .Z(n8667) );
  AND U14302 ( .A(b[21]), .B(a[83]), .Z(n8666) );
  XOR U14303 ( .A(n8671), .B(n8296), .Z(n8298) );
  XOR U14304 ( .A(n8672), .B(n8673), .Z(n8296) );
  AND U14305 ( .A(n8674), .B(n8675), .Z(n8672) );
  AND U14306 ( .A(b[20]), .B(a[84]), .Z(n8671) );
  XOR U14307 ( .A(n8676), .B(n8301), .Z(n8303) );
  XOR U14308 ( .A(n8677), .B(n8678), .Z(n8301) );
  AND U14309 ( .A(n8679), .B(n8680), .Z(n8677) );
  AND U14310 ( .A(b[19]), .B(a[85]), .Z(n8676) );
  XOR U14311 ( .A(n8681), .B(n8306), .Z(n8308) );
  XOR U14312 ( .A(n8682), .B(n8683), .Z(n8306) );
  AND U14313 ( .A(n8684), .B(n8685), .Z(n8682) );
  AND U14314 ( .A(b[18]), .B(a[86]), .Z(n8681) );
  XOR U14315 ( .A(n8686), .B(n8687), .Z(n8310) );
  AND U14316 ( .A(n8688), .B(n8689), .Z(n8686) );
  XOR U14317 ( .A(n8690), .B(n8315), .Z(n8317) );
  XOR U14318 ( .A(n8691), .B(n8692), .Z(n8315) );
  AND U14319 ( .A(n8693), .B(n8694), .Z(n8691) );
  AND U14320 ( .A(b[17]), .B(a[87]), .Z(n8690) );
  XOR U14321 ( .A(n8695), .B(n8320), .Z(n8322) );
  XOR U14322 ( .A(n8696), .B(n8697), .Z(n8320) );
  AND U14323 ( .A(n8698), .B(n8699), .Z(n8696) );
  AND U14324 ( .A(b[15]), .B(a[89]), .Z(n8695) );
  XOR U14325 ( .A(n8700), .B(n8325), .Z(n8327) );
  XOR U14326 ( .A(n8701), .B(n8702), .Z(n8325) );
  AND U14327 ( .A(n8703), .B(n8704), .Z(n8701) );
  AND U14328 ( .A(b[14]), .B(a[90]), .Z(n8700) );
  XOR U14329 ( .A(n8705), .B(n8330), .Z(n8332) );
  XOR U14330 ( .A(n8706), .B(n8707), .Z(n8330) );
  AND U14331 ( .A(n8708), .B(n8709), .Z(n8706) );
  AND U14332 ( .A(b[13]), .B(a[91]), .Z(n8705) );
  XOR U14333 ( .A(n8710), .B(n8335), .Z(n8337) );
  XOR U14334 ( .A(n8711), .B(n8712), .Z(n8335) );
  AND U14335 ( .A(n8713), .B(n8714), .Z(n8711) );
  AND U14336 ( .A(b[12]), .B(a[92]), .Z(n8710) );
  XOR U14337 ( .A(n8715), .B(n8716), .Z(n8339) );
  AND U14338 ( .A(n8717), .B(n8718), .Z(n8715) );
  XOR U14339 ( .A(n8719), .B(n8344), .Z(n8346) );
  XOR U14340 ( .A(n8720), .B(n8721), .Z(n8344) );
  AND U14341 ( .A(n8722), .B(n8723), .Z(n8720) );
  AND U14342 ( .A(b[11]), .B(a[93]), .Z(n8719) );
  XOR U14343 ( .A(n8724), .B(n8349), .Z(n8351) );
  XOR U14344 ( .A(n8725), .B(n8726), .Z(n8349) );
  AND U14345 ( .A(n8727), .B(n8728), .Z(n8725) );
  AND U14346 ( .A(b[9]), .B(a[95]), .Z(n8724) );
  XOR U14347 ( .A(n8729), .B(n8354), .Z(n8356) );
  XOR U14348 ( .A(n8730), .B(n8731), .Z(n8354) );
  AND U14349 ( .A(n8732), .B(n8733), .Z(n8730) );
  AND U14350 ( .A(b[8]), .B(a[96]), .Z(n8729) );
  XOR U14351 ( .A(n8734), .B(n8359), .Z(n8361) );
  XOR U14352 ( .A(n8735), .B(n8736), .Z(n8359) );
  AND U14353 ( .A(n8737), .B(n8738), .Z(n8735) );
  AND U14354 ( .A(b[7]), .B(a[97]), .Z(n8734) );
  XOR U14355 ( .A(n8739), .B(n8364), .Z(n8366) );
  XOR U14356 ( .A(n8740), .B(n8741), .Z(n8364) );
  AND U14357 ( .A(n8742), .B(n8743), .Z(n8740) );
  AND U14358 ( .A(b[6]), .B(a[98]), .Z(n8739) );
  XOR U14359 ( .A(n8744), .B(n8745), .Z(n8368) );
  AND U14360 ( .A(n8746), .B(n8747), .Z(n8744) );
  XOR U14361 ( .A(n8748), .B(n8373), .Z(n8375) );
  XOR U14362 ( .A(n8749), .B(n8750), .Z(n8373) );
  AND U14363 ( .A(n8751), .B(n8752), .Z(n8749) );
  AND U14364 ( .A(b[5]), .B(a[99]), .Z(n8748) );
  XNOR U14365 ( .A(n8753), .B(n8754), .Z(n8387) );
  NANDN U14366 ( .A(n8755), .B(n8756), .Z(n8754) );
  XOR U14367 ( .A(n8757), .B(n8378), .Z(n8380) );
  XNOR U14368 ( .A(n8758), .B(n8759), .Z(n8378) );
  ANDN U14369 ( .B(n8760), .A(n8761), .Z(n8758) );
  AND U14370 ( .A(b[3]), .B(a[101]), .Z(n8757) );
  NAND U14371 ( .A(a[104]), .B(b[0]), .Z(n8024) );
  XOR U14372 ( .A(n8762), .B(n8763), .Z(swire[103]) );
  XOR U14373 ( .A(n8396), .B(n8397), .Z(n8764) );
  XNOR U14374 ( .A(n8755), .B(n8756), .Z(n8397) );
  XOR U14375 ( .A(n8753), .B(n8765), .Z(n8756) );
  NAND U14376 ( .A(b[1]), .B(a[102]), .Z(n8765) );
  XNOR U14377 ( .A(n8761), .B(n8766), .Z(n8755) );
  XOR U14378 ( .A(n8753), .B(n8760), .Z(n8766) );
  XNOR U14379 ( .A(n8767), .B(n8759), .Z(n8760) );
  AND U14380 ( .A(b[2]), .B(a[101]), .Z(n8767) );
  NANDN U14381 ( .A(n8768), .B(n8769), .Z(n8753) );
  XNOR U14382 ( .A(n8759), .B(n8770), .Z(n8761) );
  XNOR U14383 ( .A(n8747), .B(n8746), .Z(n8770) );
  XOR U14384 ( .A(n8771), .B(n8745), .Z(n8746) );
  AND U14385 ( .A(b[3]), .B(a[100]), .Z(n8771) );
  XNOR U14386 ( .A(n8745), .B(n8751), .Z(n8772) );
  XNOR U14387 ( .A(n8750), .B(n8742), .Z(n8773) );
  XNOR U14388 ( .A(n8741), .B(n8737), .Z(n8774) );
  XNOR U14389 ( .A(n8736), .B(n8732), .Z(n8775) );
  XNOR U14390 ( .A(n8731), .B(n8727), .Z(n8776) );
  XNOR U14391 ( .A(n8718), .B(n8717), .Z(n8777) );
  XOR U14392 ( .A(n8778), .B(n8716), .Z(n8717) );
  AND U14393 ( .A(b[9]), .B(a[94]), .Z(n8778) );
  XNOR U14394 ( .A(n8716), .B(n8722), .Z(n8779) );
  XNOR U14395 ( .A(n8721), .B(n8713), .Z(n8780) );
  XNOR U14396 ( .A(n8712), .B(n8708), .Z(n8781) );
  XNOR U14397 ( .A(n8707), .B(n8703), .Z(n8782) );
  XNOR U14398 ( .A(n8702), .B(n8698), .Z(n8783) );
  XNOR U14399 ( .A(n8689), .B(n8688), .Z(n8784) );
  XOR U14400 ( .A(n8785), .B(n8687), .Z(n8688) );
  AND U14401 ( .A(b[15]), .B(a[88]), .Z(n8785) );
  XNOR U14402 ( .A(n8687), .B(n8693), .Z(n8786) );
  XNOR U14403 ( .A(n8692), .B(n8684), .Z(n8787) );
  XNOR U14404 ( .A(n8683), .B(n8679), .Z(n8788) );
  XNOR U14405 ( .A(n8678), .B(n8674), .Z(n8789) );
  XNOR U14406 ( .A(n8673), .B(n8669), .Z(n8790) );
  XNOR U14407 ( .A(n8660), .B(n8659), .Z(n8791) );
  XOR U14408 ( .A(n8792), .B(n8658), .Z(n8659) );
  AND U14409 ( .A(b[21]), .B(a[82]), .Z(n8792) );
  XNOR U14410 ( .A(n8658), .B(n8664), .Z(n8793) );
  XNOR U14411 ( .A(n8663), .B(n8655), .Z(n8794) );
  XNOR U14412 ( .A(n8654), .B(n8650), .Z(n8795) );
  XNOR U14413 ( .A(n8649), .B(n8645), .Z(n8796) );
  XNOR U14414 ( .A(n8644), .B(n8640), .Z(n8797) );
  XNOR U14415 ( .A(n8631), .B(n8630), .Z(n8798) );
  XOR U14416 ( .A(n8799), .B(n8629), .Z(n8630) );
  AND U14417 ( .A(b[27]), .B(a[76]), .Z(n8799) );
  XNOR U14418 ( .A(n8629), .B(n8635), .Z(n8800) );
  XNOR U14419 ( .A(n8634), .B(n8626), .Z(n8801) );
  XNOR U14420 ( .A(n8625), .B(n8621), .Z(n8802) );
  XNOR U14421 ( .A(n8620), .B(n8616), .Z(n8803) );
  XNOR U14422 ( .A(n8615), .B(n8611), .Z(n8804) );
  XNOR U14423 ( .A(n8602), .B(n8601), .Z(n8805) );
  XOR U14424 ( .A(n8806), .B(n8600), .Z(n8601) );
  AND U14425 ( .A(b[33]), .B(a[70]), .Z(n8806) );
  XNOR U14426 ( .A(n8600), .B(n8606), .Z(n8807) );
  XNOR U14427 ( .A(n8605), .B(n8597), .Z(n8808) );
  XNOR U14428 ( .A(n8596), .B(n8592), .Z(n8809) );
  XNOR U14429 ( .A(n8591), .B(n8587), .Z(n8810) );
  XNOR U14430 ( .A(n8586), .B(n8582), .Z(n8811) );
  XNOR U14431 ( .A(n8581), .B(n8577), .Z(n8812) );
  XNOR U14432 ( .A(n8576), .B(n8572), .Z(n8813) );
  XNOR U14433 ( .A(n8571), .B(n8567), .Z(n8814) );
  XNOR U14434 ( .A(n8566), .B(n8562), .Z(n8815) );
  XNOR U14435 ( .A(n8561), .B(n8557), .Z(n8816) );
  XNOR U14436 ( .A(n8556), .B(n8552), .Z(n8817) );
  XNOR U14437 ( .A(n8551), .B(n8547), .Z(n8818) );
  XNOR U14438 ( .A(n8546), .B(n8542), .Z(n8819) );
  XNOR U14439 ( .A(n8541), .B(n8537), .Z(n8820) );
  XNOR U14440 ( .A(n8536), .B(n8532), .Z(n8821) );
  XNOR U14441 ( .A(n8531), .B(n8527), .Z(n8822) );
  XNOR U14442 ( .A(n8526), .B(n8522), .Z(n8823) );
  XNOR U14443 ( .A(n8521), .B(n8517), .Z(n8824) );
  XNOR U14444 ( .A(n8516), .B(n8512), .Z(n8825) );
  XNOR U14445 ( .A(n8511), .B(n8507), .Z(n8826) );
  XNOR U14446 ( .A(n8506), .B(n8502), .Z(n8827) );
  XNOR U14447 ( .A(n8501), .B(n8497), .Z(n8828) );
  XNOR U14448 ( .A(n8496), .B(n8492), .Z(n8829) );
  XNOR U14449 ( .A(n8491), .B(n8487), .Z(n8830) );
  XNOR U14450 ( .A(n8486), .B(n8482), .Z(n8831) );
  XNOR U14451 ( .A(n8481), .B(n8477), .Z(n8832) );
  XOR U14452 ( .A(n8476), .B(n8473), .Z(n8833) );
  XOR U14453 ( .A(n8834), .B(n8835), .Z(n8473) );
  XOR U14454 ( .A(n8471), .B(n8836), .Z(n8835) );
  XOR U14455 ( .A(n8837), .B(n8838), .Z(n8836) );
  XOR U14456 ( .A(n8839), .B(n8840), .Z(n8838) );
  NAND U14457 ( .A(a[41]), .B(b[62]), .Z(n8840) );
  AND U14458 ( .A(a[40]), .B(b[63]), .Z(n8839) );
  XOR U14459 ( .A(n8841), .B(n8837), .Z(n8834) );
  XOR U14460 ( .A(n8842), .B(n8843), .Z(n8837) );
  ANDN U14461 ( .B(n8844), .A(n8845), .Z(n8842) );
  AND U14462 ( .A(a[42]), .B(b[61]), .Z(n8841) );
  XOR U14463 ( .A(n8846), .B(n8471), .Z(n8472) );
  XOR U14464 ( .A(n8847), .B(n8848), .Z(n8471) );
  AND U14465 ( .A(n8849), .B(n8850), .Z(n8847) );
  AND U14466 ( .A(a[43]), .B(b[60]), .Z(n8846) );
  XOR U14467 ( .A(n8851), .B(n8476), .Z(n8478) );
  XOR U14468 ( .A(n8852), .B(n8853), .Z(n8476) );
  AND U14469 ( .A(n8854), .B(n8855), .Z(n8852) );
  AND U14470 ( .A(a[44]), .B(b[59]), .Z(n8851) );
  XOR U14471 ( .A(n8856), .B(n8481), .Z(n8483) );
  XOR U14472 ( .A(n8857), .B(n8858), .Z(n8481) );
  AND U14473 ( .A(n8859), .B(n8860), .Z(n8857) );
  AND U14474 ( .A(a[45]), .B(b[58]), .Z(n8856) );
  XOR U14475 ( .A(n8861), .B(n8486), .Z(n8488) );
  XOR U14476 ( .A(n8862), .B(n8863), .Z(n8486) );
  AND U14477 ( .A(n8864), .B(n8865), .Z(n8862) );
  AND U14478 ( .A(a[46]), .B(b[57]), .Z(n8861) );
  XOR U14479 ( .A(n8866), .B(n8491), .Z(n8493) );
  XOR U14480 ( .A(n8867), .B(n8868), .Z(n8491) );
  AND U14481 ( .A(n8869), .B(n8870), .Z(n8867) );
  AND U14482 ( .A(a[47]), .B(b[56]), .Z(n8866) );
  XOR U14483 ( .A(n8871), .B(n8496), .Z(n8498) );
  XOR U14484 ( .A(n8872), .B(n8873), .Z(n8496) );
  AND U14485 ( .A(n8874), .B(n8875), .Z(n8872) );
  AND U14486 ( .A(a[48]), .B(b[55]), .Z(n8871) );
  XOR U14487 ( .A(n8876), .B(n8501), .Z(n8503) );
  XOR U14488 ( .A(n8877), .B(n8878), .Z(n8501) );
  AND U14489 ( .A(n8879), .B(n8880), .Z(n8877) );
  AND U14490 ( .A(a[49]), .B(b[54]), .Z(n8876) );
  XOR U14491 ( .A(n8881), .B(n8506), .Z(n8508) );
  XOR U14492 ( .A(n8882), .B(n8883), .Z(n8506) );
  AND U14493 ( .A(n8884), .B(n8885), .Z(n8882) );
  AND U14494 ( .A(a[50]), .B(b[53]), .Z(n8881) );
  XOR U14495 ( .A(n8886), .B(n8511), .Z(n8513) );
  XOR U14496 ( .A(n8887), .B(n8888), .Z(n8511) );
  AND U14497 ( .A(n8889), .B(n8890), .Z(n8887) );
  AND U14498 ( .A(a[51]), .B(b[52]), .Z(n8886) );
  XOR U14499 ( .A(n8891), .B(n8516), .Z(n8518) );
  XOR U14500 ( .A(n8892), .B(n8893), .Z(n8516) );
  AND U14501 ( .A(n8894), .B(n8895), .Z(n8892) );
  AND U14502 ( .A(b[51]), .B(a[52]), .Z(n8891) );
  XOR U14503 ( .A(n8896), .B(n8521), .Z(n8523) );
  XOR U14504 ( .A(n8897), .B(n8898), .Z(n8521) );
  AND U14505 ( .A(n8899), .B(n8900), .Z(n8897) );
  AND U14506 ( .A(b[50]), .B(a[53]), .Z(n8896) );
  XOR U14507 ( .A(n8901), .B(n8526), .Z(n8528) );
  XOR U14508 ( .A(n8902), .B(n8903), .Z(n8526) );
  AND U14509 ( .A(n8904), .B(n8905), .Z(n8902) );
  AND U14510 ( .A(b[49]), .B(a[54]), .Z(n8901) );
  XOR U14511 ( .A(n8906), .B(n8531), .Z(n8533) );
  XOR U14512 ( .A(n8907), .B(n8908), .Z(n8531) );
  AND U14513 ( .A(n8909), .B(n8910), .Z(n8907) );
  AND U14514 ( .A(b[48]), .B(a[55]), .Z(n8906) );
  XOR U14515 ( .A(n8911), .B(n8536), .Z(n8538) );
  XOR U14516 ( .A(n8912), .B(n8913), .Z(n8536) );
  AND U14517 ( .A(n8914), .B(n8915), .Z(n8912) );
  AND U14518 ( .A(b[47]), .B(a[56]), .Z(n8911) );
  XOR U14519 ( .A(n8916), .B(n8541), .Z(n8543) );
  XOR U14520 ( .A(n8917), .B(n8918), .Z(n8541) );
  AND U14521 ( .A(n8919), .B(n8920), .Z(n8917) );
  AND U14522 ( .A(b[46]), .B(a[57]), .Z(n8916) );
  XOR U14523 ( .A(n8921), .B(n8546), .Z(n8548) );
  XOR U14524 ( .A(n8922), .B(n8923), .Z(n8546) );
  AND U14525 ( .A(n8924), .B(n8925), .Z(n8922) );
  AND U14526 ( .A(b[45]), .B(a[58]), .Z(n8921) );
  XOR U14527 ( .A(n8926), .B(n8551), .Z(n8553) );
  XOR U14528 ( .A(n8927), .B(n8928), .Z(n8551) );
  AND U14529 ( .A(n8929), .B(n8930), .Z(n8927) );
  AND U14530 ( .A(b[44]), .B(a[59]), .Z(n8926) );
  XOR U14531 ( .A(n8931), .B(n8556), .Z(n8558) );
  XOR U14532 ( .A(n8932), .B(n8933), .Z(n8556) );
  AND U14533 ( .A(n8934), .B(n8935), .Z(n8932) );
  AND U14534 ( .A(b[43]), .B(a[60]), .Z(n8931) );
  XOR U14535 ( .A(n8936), .B(n8561), .Z(n8563) );
  XOR U14536 ( .A(n8937), .B(n8938), .Z(n8561) );
  AND U14537 ( .A(n8939), .B(n8940), .Z(n8937) );
  AND U14538 ( .A(b[42]), .B(a[61]), .Z(n8936) );
  XOR U14539 ( .A(n8941), .B(n8566), .Z(n8568) );
  XOR U14540 ( .A(n8942), .B(n8943), .Z(n8566) );
  AND U14541 ( .A(n8944), .B(n8945), .Z(n8942) );
  AND U14542 ( .A(b[41]), .B(a[62]), .Z(n8941) );
  XOR U14543 ( .A(n8946), .B(n8571), .Z(n8573) );
  XOR U14544 ( .A(n8947), .B(n8948), .Z(n8571) );
  AND U14545 ( .A(n8949), .B(n8950), .Z(n8947) );
  AND U14546 ( .A(b[40]), .B(a[63]), .Z(n8946) );
  XOR U14547 ( .A(n8951), .B(n8576), .Z(n8578) );
  XOR U14548 ( .A(n8952), .B(n8953), .Z(n8576) );
  AND U14549 ( .A(n8954), .B(n8955), .Z(n8952) );
  AND U14550 ( .A(b[39]), .B(a[64]), .Z(n8951) );
  XOR U14551 ( .A(n8956), .B(n8581), .Z(n8583) );
  XOR U14552 ( .A(n8957), .B(n8958), .Z(n8581) );
  AND U14553 ( .A(n8959), .B(n8960), .Z(n8957) );
  AND U14554 ( .A(b[38]), .B(a[65]), .Z(n8956) );
  XOR U14555 ( .A(n8961), .B(n8586), .Z(n8588) );
  XOR U14556 ( .A(n8962), .B(n8963), .Z(n8586) );
  AND U14557 ( .A(n8964), .B(n8965), .Z(n8962) );
  AND U14558 ( .A(b[37]), .B(a[66]), .Z(n8961) );
  XOR U14559 ( .A(n8966), .B(n8591), .Z(n8593) );
  XOR U14560 ( .A(n8967), .B(n8968), .Z(n8591) );
  AND U14561 ( .A(n8969), .B(n8970), .Z(n8967) );
  AND U14562 ( .A(b[36]), .B(a[67]), .Z(n8966) );
  XOR U14563 ( .A(n8971), .B(n8596), .Z(n8598) );
  XOR U14564 ( .A(n8972), .B(n8973), .Z(n8596) );
  AND U14565 ( .A(n8974), .B(n8975), .Z(n8972) );
  AND U14566 ( .A(b[35]), .B(a[68]), .Z(n8971) );
  XOR U14567 ( .A(n8976), .B(n8977), .Z(n8600) );
  AND U14568 ( .A(n8978), .B(n8979), .Z(n8976) );
  XOR U14569 ( .A(n8980), .B(n8605), .Z(n8607) );
  XOR U14570 ( .A(n8981), .B(n8982), .Z(n8605) );
  AND U14571 ( .A(n8983), .B(n8984), .Z(n8981) );
  AND U14572 ( .A(b[34]), .B(a[69]), .Z(n8980) );
  XOR U14573 ( .A(n8985), .B(n8610), .Z(n8612) );
  XOR U14574 ( .A(n8986), .B(n8987), .Z(n8610) );
  AND U14575 ( .A(n8988), .B(n8989), .Z(n8986) );
  AND U14576 ( .A(b[32]), .B(a[71]), .Z(n8985) );
  XOR U14577 ( .A(n8990), .B(n8615), .Z(n8617) );
  XOR U14578 ( .A(n8991), .B(n8992), .Z(n8615) );
  AND U14579 ( .A(n8993), .B(n8994), .Z(n8991) );
  AND U14580 ( .A(b[31]), .B(a[72]), .Z(n8990) );
  XOR U14581 ( .A(n8995), .B(n8620), .Z(n8622) );
  XOR U14582 ( .A(n8996), .B(n8997), .Z(n8620) );
  AND U14583 ( .A(n8998), .B(n8999), .Z(n8996) );
  AND U14584 ( .A(b[30]), .B(a[73]), .Z(n8995) );
  XOR U14585 ( .A(n9000), .B(n8625), .Z(n8627) );
  XOR U14586 ( .A(n9001), .B(n9002), .Z(n8625) );
  AND U14587 ( .A(n9003), .B(n9004), .Z(n9001) );
  AND U14588 ( .A(b[29]), .B(a[74]), .Z(n9000) );
  XOR U14589 ( .A(n9005), .B(n9006), .Z(n8629) );
  AND U14590 ( .A(n9007), .B(n9008), .Z(n9005) );
  XOR U14591 ( .A(n9009), .B(n8634), .Z(n8636) );
  XOR U14592 ( .A(n9010), .B(n9011), .Z(n8634) );
  AND U14593 ( .A(n9012), .B(n9013), .Z(n9010) );
  AND U14594 ( .A(b[28]), .B(a[75]), .Z(n9009) );
  XOR U14595 ( .A(n9014), .B(n8639), .Z(n8641) );
  XOR U14596 ( .A(n9015), .B(n9016), .Z(n8639) );
  AND U14597 ( .A(n9017), .B(n9018), .Z(n9015) );
  AND U14598 ( .A(b[26]), .B(a[77]), .Z(n9014) );
  XOR U14599 ( .A(n9019), .B(n8644), .Z(n8646) );
  XOR U14600 ( .A(n9020), .B(n9021), .Z(n8644) );
  AND U14601 ( .A(n9022), .B(n9023), .Z(n9020) );
  AND U14602 ( .A(b[25]), .B(a[78]), .Z(n9019) );
  XOR U14603 ( .A(n9024), .B(n8649), .Z(n8651) );
  XOR U14604 ( .A(n9025), .B(n9026), .Z(n8649) );
  AND U14605 ( .A(n9027), .B(n9028), .Z(n9025) );
  AND U14606 ( .A(b[24]), .B(a[79]), .Z(n9024) );
  XOR U14607 ( .A(n9029), .B(n8654), .Z(n8656) );
  XOR U14608 ( .A(n9030), .B(n9031), .Z(n8654) );
  AND U14609 ( .A(n9032), .B(n9033), .Z(n9030) );
  AND U14610 ( .A(b[23]), .B(a[80]), .Z(n9029) );
  XOR U14611 ( .A(n9034), .B(n9035), .Z(n8658) );
  AND U14612 ( .A(n9036), .B(n9037), .Z(n9034) );
  XOR U14613 ( .A(n9038), .B(n8663), .Z(n8665) );
  XOR U14614 ( .A(n9039), .B(n9040), .Z(n8663) );
  AND U14615 ( .A(n9041), .B(n9042), .Z(n9039) );
  AND U14616 ( .A(b[22]), .B(a[81]), .Z(n9038) );
  XOR U14617 ( .A(n9043), .B(n8668), .Z(n8670) );
  XOR U14618 ( .A(n9044), .B(n9045), .Z(n8668) );
  AND U14619 ( .A(n9046), .B(n9047), .Z(n9044) );
  AND U14620 ( .A(b[20]), .B(a[83]), .Z(n9043) );
  XOR U14621 ( .A(n9048), .B(n8673), .Z(n8675) );
  XOR U14622 ( .A(n9049), .B(n9050), .Z(n8673) );
  AND U14623 ( .A(n9051), .B(n9052), .Z(n9049) );
  AND U14624 ( .A(b[19]), .B(a[84]), .Z(n9048) );
  XOR U14625 ( .A(n9053), .B(n8678), .Z(n8680) );
  XOR U14626 ( .A(n9054), .B(n9055), .Z(n8678) );
  AND U14627 ( .A(n9056), .B(n9057), .Z(n9054) );
  AND U14628 ( .A(b[18]), .B(a[85]), .Z(n9053) );
  XOR U14629 ( .A(n9058), .B(n8683), .Z(n8685) );
  XOR U14630 ( .A(n9059), .B(n9060), .Z(n8683) );
  AND U14631 ( .A(n9061), .B(n9062), .Z(n9059) );
  AND U14632 ( .A(b[17]), .B(a[86]), .Z(n9058) );
  XOR U14633 ( .A(n9063), .B(n9064), .Z(n8687) );
  AND U14634 ( .A(n9065), .B(n9066), .Z(n9063) );
  XOR U14635 ( .A(n9067), .B(n8692), .Z(n8694) );
  XOR U14636 ( .A(n9068), .B(n9069), .Z(n8692) );
  AND U14637 ( .A(n9070), .B(n9071), .Z(n9068) );
  AND U14638 ( .A(b[16]), .B(a[87]), .Z(n9067) );
  XOR U14639 ( .A(n9072), .B(n8697), .Z(n8699) );
  XOR U14640 ( .A(n9073), .B(n9074), .Z(n8697) );
  AND U14641 ( .A(n9075), .B(n9076), .Z(n9073) );
  AND U14642 ( .A(b[14]), .B(a[89]), .Z(n9072) );
  XOR U14643 ( .A(n9077), .B(n8702), .Z(n8704) );
  XOR U14644 ( .A(n9078), .B(n9079), .Z(n8702) );
  AND U14645 ( .A(n9080), .B(n9081), .Z(n9078) );
  AND U14646 ( .A(b[13]), .B(a[90]), .Z(n9077) );
  XOR U14647 ( .A(n9082), .B(n8707), .Z(n8709) );
  XOR U14648 ( .A(n9083), .B(n9084), .Z(n8707) );
  AND U14649 ( .A(n9085), .B(n9086), .Z(n9083) );
  AND U14650 ( .A(b[12]), .B(a[91]), .Z(n9082) );
  XOR U14651 ( .A(n9087), .B(n8712), .Z(n8714) );
  XOR U14652 ( .A(n9088), .B(n9089), .Z(n8712) );
  AND U14653 ( .A(n9090), .B(n9091), .Z(n9088) );
  AND U14654 ( .A(b[11]), .B(a[92]), .Z(n9087) );
  XOR U14655 ( .A(n9092), .B(n9093), .Z(n8716) );
  AND U14656 ( .A(n9094), .B(n9095), .Z(n9092) );
  XOR U14657 ( .A(n9096), .B(n8721), .Z(n8723) );
  XOR U14658 ( .A(n9097), .B(n9098), .Z(n8721) );
  AND U14659 ( .A(n9099), .B(n9100), .Z(n9097) );
  AND U14660 ( .A(b[10]), .B(a[93]), .Z(n9096) );
  XOR U14661 ( .A(n9101), .B(n8726), .Z(n8728) );
  XOR U14662 ( .A(n9102), .B(n9103), .Z(n8726) );
  AND U14663 ( .A(n9104), .B(n9105), .Z(n9102) );
  AND U14664 ( .A(b[8]), .B(a[95]), .Z(n9101) );
  XOR U14665 ( .A(n9106), .B(n8731), .Z(n8733) );
  XOR U14666 ( .A(n9107), .B(n9108), .Z(n8731) );
  AND U14667 ( .A(n9109), .B(n9110), .Z(n9107) );
  AND U14668 ( .A(b[7]), .B(a[96]), .Z(n9106) );
  XOR U14669 ( .A(n9111), .B(n8736), .Z(n8738) );
  XOR U14670 ( .A(n9112), .B(n9113), .Z(n8736) );
  AND U14671 ( .A(n9114), .B(n9115), .Z(n9112) );
  AND U14672 ( .A(b[6]), .B(a[97]), .Z(n9111) );
  XOR U14673 ( .A(n9116), .B(n8741), .Z(n8743) );
  XOR U14674 ( .A(n9117), .B(n9118), .Z(n8741) );
  AND U14675 ( .A(n9119), .B(n9120), .Z(n9117) );
  AND U14676 ( .A(b[5]), .B(a[98]), .Z(n9116) );
  XOR U14677 ( .A(n9121), .B(n9122), .Z(n8745) );
  AND U14678 ( .A(n9123), .B(n9124), .Z(n9121) );
  XOR U14679 ( .A(n9125), .B(n8750), .Z(n8752) );
  XOR U14680 ( .A(n9126), .B(n9127), .Z(n8750) );
  AND U14681 ( .A(n9128), .B(n9129), .Z(n9126) );
  AND U14682 ( .A(b[4]), .B(a[99]), .Z(n9125) );
  XNOR U14683 ( .A(n9130), .B(n9131), .Z(n8759) );
  NAND U14684 ( .A(n9132), .B(n9133), .Z(n9131) );
  NAND U14685 ( .A(a[103]), .B(b[0]), .Z(n8396) );
  XOR U14686 ( .A(n9134), .B(n9135), .Z(swire[102]) );
  XOR U14687 ( .A(n8768), .B(n8769), .Z(n9136) );
  XOR U14688 ( .A(n9132), .B(n9133), .Z(n8769) );
  XOR U14689 ( .A(n9130), .B(n9137), .Z(n9133) );
  NAND U14690 ( .A(b[1]), .B(a[101]), .Z(n9137) );
  XOR U14691 ( .A(n9130), .B(n9123), .Z(n9138) );
  XNOR U14692 ( .A(n9122), .B(n9128), .Z(n9139) );
  XNOR U14693 ( .A(n9127), .B(n9119), .Z(n9140) );
  XNOR U14694 ( .A(n9118), .B(n9114), .Z(n9141) );
  XNOR U14695 ( .A(n9113), .B(n9109), .Z(n9142) );
  XNOR U14696 ( .A(n9108), .B(n9104), .Z(n9143) );
  XNOR U14697 ( .A(n9095), .B(n9094), .Z(n9144) );
  XOR U14698 ( .A(n9145), .B(n9093), .Z(n9094) );
  AND U14699 ( .A(b[8]), .B(a[94]), .Z(n9145) );
  XNOR U14700 ( .A(n9093), .B(n9099), .Z(n9146) );
  XNOR U14701 ( .A(n9098), .B(n9090), .Z(n9147) );
  XNOR U14702 ( .A(n9089), .B(n9085), .Z(n9148) );
  XNOR U14703 ( .A(n9084), .B(n9080), .Z(n9149) );
  XNOR U14704 ( .A(n9079), .B(n9075), .Z(n9150) );
  XNOR U14705 ( .A(n9066), .B(n9065), .Z(n9151) );
  XOR U14706 ( .A(n9152), .B(n9064), .Z(n9065) );
  AND U14707 ( .A(b[14]), .B(a[88]), .Z(n9152) );
  XNOR U14708 ( .A(n9064), .B(n9070), .Z(n9153) );
  XNOR U14709 ( .A(n9069), .B(n9061), .Z(n9154) );
  XNOR U14710 ( .A(n9060), .B(n9056), .Z(n9155) );
  XNOR U14711 ( .A(n9055), .B(n9051), .Z(n9156) );
  XNOR U14712 ( .A(n9050), .B(n9046), .Z(n9157) );
  XNOR U14713 ( .A(n9037), .B(n9036), .Z(n9158) );
  XOR U14714 ( .A(n9159), .B(n9035), .Z(n9036) );
  AND U14715 ( .A(b[20]), .B(a[82]), .Z(n9159) );
  XNOR U14716 ( .A(n9035), .B(n9041), .Z(n9160) );
  XNOR U14717 ( .A(n9040), .B(n9032), .Z(n9161) );
  XNOR U14718 ( .A(n9031), .B(n9027), .Z(n9162) );
  XNOR U14719 ( .A(n9026), .B(n9022), .Z(n9163) );
  XNOR U14720 ( .A(n9021), .B(n9017), .Z(n9164) );
  XNOR U14721 ( .A(n9008), .B(n9007), .Z(n9165) );
  XOR U14722 ( .A(n9166), .B(n9006), .Z(n9007) );
  AND U14723 ( .A(b[26]), .B(a[76]), .Z(n9166) );
  XNOR U14724 ( .A(n9006), .B(n9012), .Z(n9167) );
  XNOR U14725 ( .A(n9011), .B(n9003), .Z(n9168) );
  XNOR U14726 ( .A(n9002), .B(n8998), .Z(n9169) );
  XNOR U14727 ( .A(n8997), .B(n8993), .Z(n9170) );
  XNOR U14728 ( .A(n8992), .B(n8988), .Z(n9171) );
  XNOR U14729 ( .A(n8979), .B(n8978), .Z(n9172) );
  XOR U14730 ( .A(n9173), .B(n8977), .Z(n8978) );
  AND U14731 ( .A(b[32]), .B(a[70]), .Z(n9173) );
  XNOR U14732 ( .A(n8977), .B(n8983), .Z(n9174) );
  XNOR U14733 ( .A(n8982), .B(n8974), .Z(n9175) );
  XNOR U14734 ( .A(n8973), .B(n8969), .Z(n9176) );
  XNOR U14735 ( .A(n8968), .B(n8964), .Z(n9177) );
  XNOR U14736 ( .A(n8963), .B(n8959), .Z(n9178) );
  XNOR U14737 ( .A(n8958), .B(n8954), .Z(n9179) );
  XNOR U14738 ( .A(n8953), .B(n8949), .Z(n9180) );
  XNOR U14739 ( .A(n8948), .B(n8944), .Z(n9181) );
  XNOR U14740 ( .A(n8943), .B(n8939), .Z(n9182) );
  XNOR U14741 ( .A(n8938), .B(n8934), .Z(n9183) );
  XNOR U14742 ( .A(n8933), .B(n8929), .Z(n9184) );
  XNOR U14743 ( .A(n8928), .B(n8924), .Z(n9185) );
  XNOR U14744 ( .A(n8923), .B(n8919), .Z(n9186) );
  XNOR U14745 ( .A(n8918), .B(n8914), .Z(n9187) );
  XNOR U14746 ( .A(n8913), .B(n8909), .Z(n9188) );
  XNOR U14747 ( .A(n8908), .B(n8904), .Z(n9189) );
  XNOR U14748 ( .A(n8903), .B(n8899), .Z(n9190) );
  XNOR U14749 ( .A(n8898), .B(n8894), .Z(n9191) );
  XNOR U14750 ( .A(n8893), .B(n8889), .Z(n9192) );
  XNOR U14751 ( .A(n8888), .B(n8884), .Z(n9193) );
  XNOR U14752 ( .A(n8883), .B(n8879), .Z(n9194) );
  XNOR U14753 ( .A(n8878), .B(n8874), .Z(n9195) );
  XNOR U14754 ( .A(n8873), .B(n8869), .Z(n9196) );
  XNOR U14755 ( .A(n8868), .B(n8864), .Z(n9197) );
  XNOR U14756 ( .A(n8863), .B(n8859), .Z(n9198) );
  XNOR U14757 ( .A(n8858), .B(n8854), .Z(n9199) );
  XNOR U14758 ( .A(n8853), .B(n8849), .Z(n9200) );
  XOR U14759 ( .A(n8848), .B(n8845), .Z(n9201) );
  XOR U14760 ( .A(n9202), .B(n9203), .Z(n8845) );
  XOR U14761 ( .A(n8843), .B(n9204), .Z(n9203) );
  XOR U14762 ( .A(n9205), .B(n9206), .Z(n9204) );
  XOR U14763 ( .A(n9207), .B(n9208), .Z(n9206) );
  NAND U14764 ( .A(a[40]), .B(b[62]), .Z(n9208) );
  AND U14765 ( .A(a[39]), .B(b[63]), .Z(n9207) );
  XOR U14766 ( .A(n9209), .B(n9205), .Z(n9202) );
  XOR U14767 ( .A(n9210), .B(n9211), .Z(n9205) );
  ANDN U14768 ( .B(n9212), .A(n9213), .Z(n9210) );
  AND U14769 ( .A(a[41]), .B(b[61]), .Z(n9209) );
  XOR U14770 ( .A(n9214), .B(n8843), .Z(n8844) );
  XOR U14771 ( .A(n9215), .B(n9216), .Z(n8843) );
  AND U14772 ( .A(n9217), .B(n9218), .Z(n9215) );
  AND U14773 ( .A(a[42]), .B(b[60]), .Z(n9214) );
  XOR U14774 ( .A(n9219), .B(n8848), .Z(n8850) );
  XOR U14775 ( .A(n9220), .B(n9221), .Z(n8848) );
  AND U14776 ( .A(n9222), .B(n9223), .Z(n9220) );
  AND U14777 ( .A(a[43]), .B(b[59]), .Z(n9219) );
  XOR U14778 ( .A(n9224), .B(n8853), .Z(n8855) );
  XOR U14779 ( .A(n9225), .B(n9226), .Z(n8853) );
  AND U14780 ( .A(n9227), .B(n9228), .Z(n9225) );
  AND U14781 ( .A(a[44]), .B(b[58]), .Z(n9224) );
  XOR U14782 ( .A(n9229), .B(n8858), .Z(n8860) );
  XOR U14783 ( .A(n9230), .B(n9231), .Z(n8858) );
  AND U14784 ( .A(n9232), .B(n9233), .Z(n9230) );
  AND U14785 ( .A(a[45]), .B(b[57]), .Z(n9229) );
  XOR U14786 ( .A(n9234), .B(n8863), .Z(n8865) );
  XOR U14787 ( .A(n9235), .B(n9236), .Z(n8863) );
  AND U14788 ( .A(n9237), .B(n9238), .Z(n9235) );
  AND U14789 ( .A(a[46]), .B(b[56]), .Z(n9234) );
  XOR U14790 ( .A(n9239), .B(n8868), .Z(n8870) );
  XOR U14791 ( .A(n9240), .B(n9241), .Z(n8868) );
  AND U14792 ( .A(n9242), .B(n9243), .Z(n9240) );
  AND U14793 ( .A(a[47]), .B(b[55]), .Z(n9239) );
  XOR U14794 ( .A(n9244), .B(n8873), .Z(n8875) );
  XOR U14795 ( .A(n9245), .B(n9246), .Z(n8873) );
  AND U14796 ( .A(n9247), .B(n9248), .Z(n9245) );
  AND U14797 ( .A(a[48]), .B(b[54]), .Z(n9244) );
  XOR U14798 ( .A(n9249), .B(n8878), .Z(n8880) );
  XOR U14799 ( .A(n9250), .B(n9251), .Z(n8878) );
  AND U14800 ( .A(n9252), .B(n9253), .Z(n9250) );
  AND U14801 ( .A(a[49]), .B(b[53]), .Z(n9249) );
  XOR U14802 ( .A(n9254), .B(n8883), .Z(n8885) );
  XOR U14803 ( .A(n9255), .B(n9256), .Z(n8883) );
  AND U14804 ( .A(n9257), .B(n9258), .Z(n9255) );
  AND U14805 ( .A(a[50]), .B(b[52]), .Z(n9254) );
  XOR U14806 ( .A(n9259), .B(n8888), .Z(n8890) );
  XOR U14807 ( .A(n9260), .B(n9261), .Z(n8888) );
  AND U14808 ( .A(n9262), .B(n9263), .Z(n9260) );
  AND U14809 ( .A(a[51]), .B(b[51]), .Z(n9259) );
  XOR U14810 ( .A(n9264), .B(n8893), .Z(n8895) );
  XOR U14811 ( .A(n9265), .B(n9266), .Z(n8893) );
  AND U14812 ( .A(n9267), .B(n9268), .Z(n9265) );
  AND U14813 ( .A(b[50]), .B(a[52]), .Z(n9264) );
  XOR U14814 ( .A(n9269), .B(n8898), .Z(n8900) );
  XOR U14815 ( .A(n9270), .B(n9271), .Z(n8898) );
  AND U14816 ( .A(n9272), .B(n9273), .Z(n9270) );
  AND U14817 ( .A(b[49]), .B(a[53]), .Z(n9269) );
  XOR U14818 ( .A(n9274), .B(n8903), .Z(n8905) );
  XOR U14819 ( .A(n9275), .B(n9276), .Z(n8903) );
  AND U14820 ( .A(n9277), .B(n9278), .Z(n9275) );
  AND U14821 ( .A(b[48]), .B(a[54]), .Z(n9274) );
  XOR U14822 ( .A(n9279), .B(n8908), .Z(n8910) );
  XOR U14823 ( .A(n9280), .B(n9281), .Z(n8908) );
  AND U14824 ( .A(n9282), .B(n9283), .Z(n9280) );
  AND U14825 ( .A(b[47]), .B(a[55]), .Z(n9279) );
  XOR U14826 ( .A(n9284), .B(n8913), .Z(n8915) );
  XOR U14827 ( .A(n9285), .B(n9286), .Z(n8913) );
  AND U14828 ( .A(n9287), .B(n9288), .Z(n9285) );
  AND U14829 ( .A(b[46]), .B(a[56]), .Z(n9284) );
  XOR U14830 ( .A(n9289), .B(n8918), .Z(n8920) );
  XOR U14831 ( .A(n9290), .B(n9291), .Z(n8918) );
  AND U14832 ( .A(n9292), .B(n9293), .Z(n9290) );
  AND U14833 ( .A(b[45]), .B(a[57]), .Z(n9289) );
  XOR U14834 ( .A(n9294), .B(n8923), .Z(n8925) );
  XOR U14835 ( .A(n9295), .B(n9296), .Z(n8923) );
  AND U14836 ( .A(n9297), .B(n9298), .Z(n9295) );
  AND U14837 ( .A(b[44]), .B(a[58]), .Z(n9294) );
  XOR U14838 ( .A(n9299), .B(n8928), .Z(n8930) );
  XOR U14839 ( .A(n9300), .B(n9301), .Z(n8928) );
  AND U14840 ( .A(n9302), .B(n9303), .Z(n9300) );
  AND U14841 ( .A(b[43]), .B(a[59]), .Z(n9299) );
  XOR U14842 ( .A(n9304), .B(n8933), .Z(n8935) );
  XOR U14843 ( .A(n9305), .B(n9306), .Z(n8933) );
  AND U14844 ( .A(n9307), .B(n9308), .Z(n9305) );
  AND U14845 ( .A(b[42]), .B(a[60]), .Z(n9304) );
  XOR U14846 ( .A(n9309), .B(n8938), .Z(n8940) );
  XOR U14847 ( .A(n9310), .B(n9311), .Z(n8938) );
  AND U14848 ( .A(n9312), .B(n9313), .Z(n9310) );
  AND U14849 ( .A(b[41]), .B(a[61]), .Z(n9309) );
  XOR U14850 ( .A(n9314), .B(n8943), .Z(n8945) );
  XOR U14851 ( .A(n9315), .B(n9316), .Z(n8943) );
  AND U14852 ( .A(n9317), .B(n9318), .Z(n9315) );
  AND U14853 ( .A(b[40]), .B(a[62]), .Z(n9314) );
  XOR U14854 ( .A(n9319), .B(n8948), .Z(n8950) );
  XOR U14855 ( .A(n9320), .B(n9321), .Z(n8948) );
  AND U14856 ( .A(n9322), .B(n9323), .Z(n9320) );
  AND U14857 ( .A(b[39]), .B(a[63]), .Z(n9319) );
  XOR U14858 ( .A(n9324), .B(n8953), .Z(n8955) );
  XOR U14859 ( .A(n9325), .B(n9326), .Z(n8953) );
  AND U14860 ( .A(n9327), .B(n9328), .Z(n9325) );
  AND U14861 ( .A(b[38]), .B(a[64]), .Z(n9324) );
  XOR U14862 ( .A(n9329), .B(n8958), .Z(n8960) );
  XOR U14863 ( .A(n9330), .B(n9331), .Z(n8958) );
  AND U14864 ( .A(n9332), .B(n9333), .Z(n9330) );
  AND U14865 ( .A(b[37]), .B(a[65]), .Z(n9329) );
  XOR U14866 ( .A(n9334), .B(n8963), .Z(n8965) );
  XOR U14867 ( .A(n9335), .B(n9336), .Z(n8963) );
  AND U14868 ( .A(n9337), .B(n9338), .Z(n9335) );
  AND U14869 ( .A(b[36]), .B(a[66]), .Z(n9334) );
  XOR U14870 ( .A(n9339), .B(n8968), .Z(n8970) );
  XOR U14871 ( .A(n9340), .B(n9341), .Z(n8968) );
  AND U14872 ( .A(n9342), .B(n9343), .Z(n9340) );
  AND U14873 ( .A(b[35]), .B(a[67]), .Z(n9339) );
  XOR U14874 ( .A(n9344), .B(n8973), .Z(n8975) );
  XOR U14875 ( .A(n9345), .B(n9346), .Z(n8973) );
  AND U14876 ( .A(n9347), .B(n9348), .Z(n9345) );
  AND U14877 ( .A(b[34]), .B(a[68]), .Z(n9344) );
  XOR U14878 ( .A(n9349), .B(n9350), .Z(n8977) );
  AND U14879 ( .A(n9351), .B(n9352), .Z(n9349) );
  XOR U14880 ( .A(n9353), .B(n8982), .Z(n8984) );
  XOR U14881 ( .A(n9354), .B(n9355), .Z(n8982) );
  AND U14882 ( .A(n9356), .B(n9357), .Z(n9354) );
  AND U14883 ( .A(b[33]), .B(a[69]), .Z(n9353) );
  XOR U14884 ( .A(n9358), .B(n8987), .Z(n8989) );
  XOR U14885 ( .A(n9359), .B(n9360), .Z(n8987) );
  AND U14886 ( .A(n9361), .B(n9362), .Z(n9359) );
  AND U14887 ( .A(b[31]), .B(a[71]), .Z(n9358) );
  XOR U14888 ( .A(n9363), .B(n8992), .Z(n8994) );
  XOR U14889 ( .A(n9364), .B(n9365), .Z(n8992) );
  AND U14890 ( .A(n9366), .B(n9367), .Z(n9364) );
  AND U14891 ( .A(b[30]), .B(a[72]), .Z(n9363) );
  XOR U14892 ( .A(n9368), .B(n8997), .Z(n8999) );
  XOR U14893 ( .A(n9369), .B(n9370), .Z(n8997) );
  AND U14894 ( .A(n9371), .B(n9372), .Z(n9369) );
  AND U14895 ( .A(b[29]), .B(a[73]), .Z(n9368) );
  XOR U14896 ( .A(n9373), .B(n9002), .Z(n9004) );
  XOR U14897 ( .A(n9374), .B(n9375), .Z(n9002) );
  AND U14898 ( .A(n9376), .B(n9377), .Z(n9374) );
  AND U14899 ( .A(b[28]), .B(a[74]), .Z(n9373) );
  XOR U14900 ( .A(n9378), .B(n9379), .Z(n9006) );
  AND U14901 ( .A(n9380), .B(n9381), .Z(n9378) );
  XOR U14902 ( .A(n9382), .B(n9011), .Z(n9013) );
  XOR U14903 ( .A(n9383), .B(n9384), .Z(n9011) );
  AND U14904 ( .A(n9385), .B(n9386), .Z(n9383) );
  AND U14905 ( .A(b[27]), .B(a[75]), .Z(n9382) );
  XOR U14906 ( .A(n9387), .B(n9016), .Z(n9018) );
  XOR U14907 ( .A(n9388), .B(n9389), .Z(n9016) );
  AND U14908 ( .A(n9390), .B(n9391), .Z(n9388) );
  AND U14909 ( .A(b[25]), .B(a[77]), .Z(n9387) );
  XOR U14910 ( .A(n9392), .B(n9021), .Z(n9023) );
  XOR U14911 ( .A(n9393), .B(n9394), .Z(n9021) );
  AND U14912 ( .A(n9395), .B(n9396), .Z(n9393) );
  AND U14913 ( .A(b[24]), .B(a[78]), .Z(n9392) );
  XOR U14914 ( .A(n9397), .B(n9026), .Z(n9028) );
  XOR U14915 ( .A(n9398), .B(n9399), .Z(n9026) );
  AND U14916 ( .A(n9400), .B(n9401), .Z(n9398) );
  AND U14917 ( .A(b[23]), .B(a[79]), .Z(n9397) );
  XOR U14918 ( .A(n9402), .B(n9031), .Z(n9033) );
  XOR U14919 ( .A(n9403), .B(n9404), .Z(n9031) );
  AND U14920 ( .A(n9405), .B(n9406), .Z(n9403) );
  AND U14921 ( .A(b[22]), .B(a[80]), .Z(n9402) );
  XOR U14922 ( .A(n9407), .B(n9408), .Z(n9035) );
  AND U14923 ( .A(n9409), .B(n9410), .Z(n9407) );
  XOR U14924 ( .A(n9411), .B(n9040), .Z(n9042) );
  XOR U14925 ( .A(n9412), .B(n9413), .Z(n9040) );
  AND U14926 ( .A(n9414), .B(n9415), .Z(n9412) );
  AND U14927 ( .A(b[21]), .B(a[81]), .Z(n9411) );
  XOR U14928 ( .A(n9416), .B(n9045), .Z(n9047) );
  XOR U14929 ( .A(n9417), .B(n9418), .Z(n9045) );
  AND U14930 ( .A(n9419), .B(n9420), .Z(n9417) );
  AND U14931 ( .A(b[19]), .B(a[83]), .Z(n9416) );
  XOR U14932 ( .A(n9421), .B(n9050), .Z(n9052) );
  XOR U14933 ( .A(n9422), .B(n9423), .Z(n9050) );
  AND U14934 ( .A(n9424), .B(n9425), .Z(n9422) );
  AND U14935 ( .A(b[18]), .B(a[84]), .Z(n9421) );
  XOR U14936 ( .A(n9426), .B(n9055), .Z(n9057) );
  XOR U14937 ( .A(n9427), .B(n9428), .Z(n9055) );
  AND U14938 ( .A(n9429), .B(n9430), .Z(n9427) );
  AND U14939 ( .A(b[17]), .B(a[85]), .Z(n9426) );
  XOR U14940 ( .A(n9431), .B(n9060), .Z(n9062) );
  XOR U14941 ( .A(n9432), .B(n9433), .Z(n9060) );
  AND U14942 ( .A(n9434), .B(n9435), .Z(n9432) );
  AND U14943 ( .A(b[16]), .B(a[86]), .Z(n9431) );
  XOR U14944 ( .A(n9436), .B(n9437), .Z(n9064) );
  AND U14945 ( .A(n9438), .B(n9439), .Z(n9436) );
  XOR U14946 ( .A(n9440), .B(n9069), .Z(n9071) );
  XOR U14947 ( .A(n9441), .B(n9442), .Z(n9069) );
  AND U14948 ( .A(n9443), .B(n9444), .Z(n9441) );
  AND U14949 ( .A(b[15]), .B(a[87]), .Z(n9440) );
  XOR U14950 ( .A(n9445), .B(n9074), .Z(n9076) );
  XOR U14951 ( .A(n9446), .B(n9447), .Z(n9074) );
  AND U14952 ( .A(n9448), .B(n9449), .Z(n9446) );
  AND U14953 ( .A(b[13]), .B(a[89]), .Z(n9445) );
  XOR U14954 ( .A(n9450), .B(n9079), .Z(n9081) );
  XOR U14955 ( .A(n9451), .B(n9452), .Z(n9079) );
  AND U14956 ( .A(n9453), .B(n9454), .Z(n9451) );
  AND U14957 ( .A(b[12]), .B(a[90]), .Z(n9450) );
  XOR U14958 ( .A(n9455), .B(n9084), .Z(n9086) );
  XOR U14959 ( .A(n9456), .B(n9457), .Z(n9084) );
  AND U14960 ( .A(n9458), .B(n9459), .Z(n9456) );
  AND U14961 ( .A(b[11]), .B(a[91]), .Z(n9455) );
  XOR U14962 ( .A(n9460), .B(n9089), .Z(n9091) );
  XOR U14963 ( .A(n9461), .B(n9462), .Z(n9089) );
  AND U14964 ( .A(n9463), .B(n9464), .Z(n9461) );
  AND U14965 ( .A(b[10]), .B(a[92]), .Z(n9460) );
  XOR U14966 ( .A(n9465), .B(n9466), .Z(n9093) );
  AND U14967 ( .A(n9467), .B(n9468), .Z(n9465) );
  XOR U14968 ( .A(n9469), .B(n9098), .Z(n9100) );
  XOR U14969 ( .A(n9470), .B(n9471), .Z(n9098) );
  AND U14970 ( .A(n9472), .B(n9473), .Z(n9470) );
  AND U14971 ( .A(b[9]), .B(a[93]), .Z(n9469) );
  XOR U14972 ( .A(n9474), .B(n9103), .Z(n9105) );
  XOR U14973 ( .A(n9475), .B(n9476), .Z(n9103) );
  AND U14974 ( .A(n9477), .B(n9478), .Z(n9475) );
  AND U14975 ( .A(b[7]), .B(a[95]), .Z(n9474) );
  XOR U14976 ( .A(n9479), .B(n9108), .Z(n9110) );
  XOR U14977 ( .A(n9480), .B(n9481), .Z(n9108) );
  AND U14978 ( .A(n9482), .B(n9483), .Z(n9480) );
  AND U14979 ( .A(b[6]), .B(a[96]), .Z(n9479) );
  XOR U14980 ( .A(n9484), .B(n9113), .Z(n9115) );
  XOR U14981 ( .A(n9485), .B(n9486), .Z(n9113) );
  AND U14982 ( .A(n9487), .B(n9488), .Z(n9485) );
  AND U14983 ( .A(b[5]), .B(a[97]), .Z(n9484) );
  XOR U14984 ( .A(n9489), .B(n9118), .Z(n9120) );
  XOR U14985 ( .A(n9490), .B(n9491), .Z(n9118) );
  AND U14986 ( .A(n9492), .B(n9493), .Z(n9490) );
  AND U14987 ( .A(b[4]), .B(a[98]), .Z(n9489) );
  XOR U14988 ( .A(n9494), .B(n9127), .Z(n9129) );
  XNOR U14989 ( .A(n9495), .B(n9496), .Z(n9127) );
  ANDN U14990 ( .B(n9497), .A(n9498), .Z(n9495) );
  AND U14991 ( .A(b[3]), .B(a[99]), .Z(n9494) );
  NANDN U14992 ( .A(n9499), .B(n9500), .Z(n9130) );
  XOR U14993 ( .A(n9501), .B(n9122), .Z(n9124) );
  XNOR U14994 ( .A(n9502), .B(n9503), .Z(n9122) );
  OR U14995 ( .A(n9504), .B(n9505), .Z(n9503) );
  AND U14996 ( .A(b[2]), .B(a[100]), .Z(n9501) );
  NAND U14997 ( .A(a[102]), .B(b[0]), .Z(n8768) );
  XOR U14998 ( .A(n9506), .B(n9507), .Z(swire[101]) );
  XOR U14999 ( .A(n9499), .B(n9500), .Z(n9508) );
  XOR U15000 ( .A(n9505), .B(n9504), .Z(n9500) );
  XOR U15001 ( .A(n9502), .B(n9509), .Z(n9504) );
  NAND U15002 ( .A(b[1]), .B(a[100]), .Z(n9509) );
  XOR U15003 ( .A(n9502), .B(n9498), .Z(n9510) );
  XOR U15004 ( .A(n9511), .B(n9496), .Z(n9498) );
  AND U15005 ( .A(b[2]), .B(a[99]), .Z(n9511) );
  ANDN U15006 ( .B(n9512), .A(n9513), .Z(n9502) );
  XOR U15007 ( .A(n9496), .B(n9492), .Z(n9514) );
  XNOR U15008 ( .A(n9491), .B(n9487), .Z(n9515) );
  XNOR U15009 ( .A(n9486), .B(n9482), .Z(n9516) );
  XNOR U15010 ( .A(n9481), .B(n9477), .Z(n9517) );
  XNOR U15011 ( .A(n9468), .B(n9467), .Z(n9518) );
  XOR U15012 ( .A(n9519), .B(n9466), .Z(n9467) );
  AND U15013 ( .A(b[7]), .B(a[94]), .Z(n9519) );
  XNOR U15014 ( .A(n9466), .B(n9472), .Z(n9520) );
  XNOR U15015 ( .A(n9471), .B(n9463), .Z(n9521) );
  XNOR U15016 ( .A(n9462), .B(n9458), .Z(n9522) );
  XNOR U15017 ( .A(n9457), .B(n9453), .Z(n9523) );
  XNOR U15018 ( .A(n9452), .B(n9448), .Z(n9524) );
  XNOR U15019 ( .A(n9439), .B(n9438), .Z(n9525) );
  XOR U15020 ( .A(n9526), .B(n9437), .Z(n9438) );
  AND U15021 ( .A(b[13]), .B(a[88]), .Z(n9526) );
  XNOR U15022 ( .A(n9437), .B(n9443), .Z(n9527) );
  XNOR U15023 ( .A(n9442), .B(n9434), .Z(n9528) );
  XNOR U15024 ( .A(n9433), .B(n9429), .Z(n9529) );
  XNOR U15025 ( .A(n9428), .B(n9424), .Z(n9530) );
  XNOR U15026 ( .A(n9423), .B(n9419), .Z(n9531) );
  XNOR U15027 ( .A(n9410), .B(n9409), .Z(n9532) );
  XOR U15028 ( .A(n9533), .B(n9408), .Z(n9409) );
  AND U15029 ( .A(b[19]), .B(a[82]), .Z(n9533) );
  XNOR U15030 ( .A(n9408), .B(n9414), .Z(n9534) );
  XNOR U15031 ( .A(n9413), .B(n9405), .Z(n9535) );
  XNOR U15032 ( .A(n9404), .B(n9400), .Z(n9536) );
  XNOR U15033 ( .A(n9399), .B(n9395), .Z(n9537) );
  XNOR U15034 ( .A(n9394), .B(n9390), .Z(n9538) );
  XNOR U15035 ( .A(n9381), .B(n9380), .Z(n9539) );
  XOR U15036 ( .A(n9540), .B(n9379), .Z(n9380) );
  AND U15037 ( .A(b[25]), .B(a[76]), .Z(n9540) );
  XNOR U15038 ( .A(n9379), .B(n9385), .Z(n9541) );
  XNOR U15039 ( .A(n9384), .B(n9376), .Z(n9542) );
  XNOR U15040 ( .A(n9375), .B(n9371), .Z(n9543) );
  XNOR U15041 ( .A(n9370), .B(n9366), .Z(n9544) );
  XNOR U15042 ( .A(n9365), .B(n9361), .Z(n9545) );
  XNOR U15043 ( .A(n9352), .B(n9351), .Z(n9546) );
  XOR U15044 ( .A(n9547), .B(n9350), .Z(n9351) );
  AND U15045 ( .A(b[31]), .B(a[70]), .Z(n9547) );
  XNOR U15046 ( .A(n9350), .B(n9356), .Z(n9548) );
  XNOR U15047 ( .A(n9355), .B(n9347), .Z(n9549) );
  XNOR U15048 ( .A(n9346), .B(n9342), .Z(n9550) );
  XNOR U15049 ( .A(n9341), .B(n9337), .Z(n9551) );
  XNOR U15050 ( .A(n9336), .B(n9332), .Z(n9552) );
  XNOR U15051 ( .A(n9331), .B(n9327), .Z(n9553) );
  XNOR U15052 ( .A(n9326), .B(n9322), .Z(n9554) );
  XNOR U15053 ( .A(n9321), .B(n9317), .Z(n9555) );
  XNOR U15054 ( .A(n9316), .B(n9312), .Z(n9556) );
  XNOR U15055 ( .A(n9311), .B(n9307), .Z(n9557) );
  XNOR U15056 ( .A(n9306), .B(n9302), .Z(n9558) );
  XNOR U15057 ( .A(n9301), .B(n9297), .Z(n9559) );
  XNOR U15058 ( .A(n9296), .B(n9292), .Z(n9560) );
  XNOR U15059 ( .A(n9291), .B(n9287), .Z(n9561) );
  XNOR U15060 ( .A(n9286), .B(n9282), .Z(n9562) );
  XNOR U15061 ( .A(n9281), .B(n9277), .Z(n9563) );
  XNOR U15062 ( .A(n9276), .B(n9272), .Z(n9564) );
  XNOR U15063 ( .A(n9271), .B(n9267), .Z(n9565) );
  XNOR U15064 ( .A(n9266), .B(n9262), .Z(n9566) );
  XNOR U15065 ( .A(n9261), .B(n9257), .Z(n9567) );
  XNOR U15066 ( .A(n9256), .B(n9252), .Z(n9568) );
  XNOR U15067 ( .A(n9251), .B(n9247), .Z(n9569) );
  XNOR U15068 ( .A(n9246), .B(n9242), .Z(n9570) );
  XNOR U15069 ( .A(n9241), .B(n9237), .Z(n9571) );
  XNOR U15070 ( .A(n9236), .B(n9232), .Z(n9572) );
  XNOR U15071 ( .A(n9231), .B(n9227), .Z(n9573) );
  XNOR U15072 ( .A(n9226), .B(n9222), .Z(n9574) );
  XNOR U15073 ( .A(n9221), .B(n9217), .Z(n9575) );
  XOR U15074 ( .A(n9216), .B(n9213), .Z(n9576) );
  XOR U15075 ( .A(n9577), .B(n9578), .Z(n9213) );
  XOR U15076 ( .A(n9211), .B(n9579), .Z(n9578) );
  XOR U15077 ( .A(n9580), .B(n9581), .Z(n9579) );
  XOR U15078 ( .A(n9582), .B(n9583), .Z(n9581) );
  NAND U15079 ( .A(a[39]), .B(b[62]), .Z(n9583) );
  AND U15080 ( .A(a[38]), .B(b[63]), .Z(n9582) );
  XOR U15081 ( .A(n9584), .B(n9580), .Z(n9577) );
  XOR U15082 ( .A(n9585), .B(n9586), .Z(n9580) );
  ANDN U15083 ( .B(n9587), .A(n9588), .Z(n9585) );
  AND U15084 ( .A(a[40]), .B(b[61]), .Z(n9584) );
  XOR U15085 ( .A(n9589), .B(n9211), .Z(n9212) );
  XOR U15086 ( .A(n9590), .B(n9591), .Z(n9211) );
  AND U15087 ( .A(n9592), .B(n9593), .Z(n9590) );
  AND U15088 ( .A(a[41]), .B(b[60]), .Z(n9589) );
  XOR U15089 ( .A(n9594), .B(n9216), .Z(n9218) );
  XOR U15090 ( .A(n9595), .B(n9596), .Z(n9216) );
  AND U15091 ( .A(n9597), .B(n9598), .Z(n9595) );
  AND U15092 ( .A(a[42]), .B(b[59]), .Z(n9594) );
  XOR U15093 ( .A(n9599), .B(n9221), .Z(n9223) );
  XOR U15094 ( .A(n9600), .B(n9601), .Z(n9221) );
  AND U15095 ( .A(n9602), .B(n9603), .Z(n9600) );
  AND U15096 ( .A(a[43]), .B(b[58]), .Z(n9599) );
  XOR U15097 ( .A(n9604), .B(n9226), .Z(n9228) );
  XOR U15098 ( .A(n9605), .B(n9606), .Z(n9226) );
  AND U15099 ( .A(n9607), .B(n9608), .Z(n9605) );
  AND U15100 ( .A(a[44]), .B(b[57]), .Z(n9604) );
  XOR U15101 ( .A(n9609), .B(n9231), .Z(n9233) );
  XOR U15102 ( .A(n9610), .B(n9611), .Z(n9231) );
  AND U15103 ( .A(n9612), .B(n9613), .Z(n9610) );
  AND U15104 ( .A(a[45]), .B(b[56]), .Z(n9609) );
  XOR U15105 ( .A(n9614), .B(n9236), .Z(n9238) );
  XOR U15106 ( .A(n9615), .B(n9616), .Z(n9236) );
  AND U15107 ( .A(n9617), .B(n9618), .Z(n9615) );
  AND U15108 ( .A(a[46]), .B(b[55]), .Z(n9614) );
  XOR U15109 ( .A(n9619), .B(n9241), .Z(n9243) );
  XOR U15110 ( .A(n9620), .B(n9621), .Z(n9241) );
  AND U15111 ( .A(n9622), .B(n9623), .Z(n9620) );
  AND U15112 ( .A(a[47]), .B(b[54]), .Z(n9619) );
  XOR U15113 ( .A(n9624), .B(n9246), .Z(n9248) );
  XOR U15114 ( .A(n9625), .B(n9626), .Z(n9246) );
  AND U15115 ( .A(n9627), .B(n9628), .Z(n9625) );
  AND U15116 ( .A(a[48]), .B(b[53]), .Z(n9624) );
  XOR U15117 ( .A(n9629), .B(n9251), .Z(n9253) );
  XOR U15118 ( .A(n9630), .B(n9631), .Z(n9251) );
  AND U15119 ( .A(n9632), .B(n9633), .Z(n9630) );
  AND U15120 ( .A(a[49]), .B(b[52]), .Z(n9629) );
  XOR U15121 ( .A(n9634), .B(n9256), .Z(n9258) );
  XOR U15122 ( .A(n9635), .B(n9636), .Z(n9256) );
  AND U15123 ( .A(n9637), .B(n9638), .Z(n9635) );
  AND U15124 ( .A(a[50]), .B(b[51]), .Z(n9634) );
  XOR U15125 ( .A(n9639), .B(n9261), .Z(n9263) );
  XOR U15126 ( .A(n9640), .B(n9641), .Z(n9261) );
  AND U15127 ( .A(n9642), .B(n9643), .Z(n9640) );
  AND U15128 ( .A(b[50]), .B(a[51]), .Z(n9639) );
  XOR U15129 ( .A(n9644), .B(n9266), .Z(n9268) );
  XOR U15130 ( .A(n9645), .B(n9646), .Z(n9266) );
  AND U15131 ( .A(n9647), .B(n9648), .Z(n9645) );
  AND U15132 ( .A(b[49]), .B(a[52]), .Z(n9644) );
  XOR U15133 ( .A(n9649), .B(n9271), .Z(n9273) );
  XOR U15134 ( .A(n9650), .B(n9651), .Z(n9271) );
  AND U15135 ( .A(n9652), .B(n9653), .Z(n9650) );
  AND U15136 ( .A(b[48]), .B(a[53]), .Z(n9649) );
  XOR U15137 ( .A(n9654), .B(n9276), .Z(n9278) );
  XOR U15138 ( .A(n9655), .B(n9656), .Z(n9276) );
  AND U15139 ( .A(n9657), .B(n9658), .Z(n9655) );
  AND U15140 ( .A(b[47]), .B(a[54]), .Z(n9654) );
  XOR U15141 ( .A(n9659), .B(n9281), .Z(n9283) );
  XOR U15142 ( .A(n9660), .B(n9661), .Z(n9281) );
  AND U15143 ( .A(n9662), .B(n9663), .Z(n9660) );
  AND U15144 ( .A(b[46]), .B(a[55]), .Z(n9659) );
  XOR U15145 ( .A(n9664), .B(n9286), .Z(n9288) );
  XOR U15146 ( .A(n9665), .B(n9666), .Z(n9286) );
  AND U15147 ( .A(n9667), .B(n9668), .Z(n9665) );
  AND U15148 ( .A(b[45]), .B(a[56]), .Z(n9664) );
  XOR U15149 ( .A(n9669), .B(n9291), .Z(n9293) );
  XOR U15150 ( .A(n9670), .B(n9671), .Z(n9291) );
  AND U15151 ( .A(n9672), .B(n9673), .Z(n9670) );
  AND U15152 ( .A(b[44]), .B(a[57]), .Z(n9669) );
  XOR U15153 ( .A(n9674), .B(n9296), .Z(n9298) );
  XOR U15154 ( .A(n9675), .B(n9676), .Z(n9296) );
  AND U15155 ( .A(n9677), .B(n9678), .Z(n9675) );
  AND U15156 ( .A(b[43]), .B(a[58]), .Z(n9674) );
  XOR U15157 ( .A(n9679), .B(n9301), .Z(n9303) );
  XOR U15158 ( .A(n9680), .B(n9681), .Z(n9301) );
  AND U15159 ( .A(n9682), .B(n9683), .Z(n9680) );
  AND U15160 ( .A(b[42]), .B(a[59]), .Z(n9679) );
  XOR U15161 ( .A(n9684), .B(n9306), .Z(n9308) );
  XOR U15162 ( .A(n9685), .B(n9686), .Z(n9306) );
  AND U15163 ( .A(n9687), .B(n9688), .Z(n9685) );
  AND U15164 ( .A(b[41]), .B(a[60]), .Z(n9684) );
  XOR U15165 ( .A(n9689), .B(n9311), .Z(n9313) );
  XOR U15166 ( .A(n9690), .B(n9691), .Z(n9311) );
  AND U15167 ( .A(n9692), .B(n9693), .Z(n9690) );
  AND U15168 ( .A(b[40]), .B(a[61]), .Z(n9689) );
  XOR U15169 ( .A(n9694), .B(n9316), .Z(n9318) );
  XOR U15170 ( .A(n9695), .B(n9696), .Z(n9316) );
  AND U15171 ( .A(n9697), .B(n9698), .Z(n9695) );
  AND U15172 ( .A(b[39]), .B(a[62]), .Z(n9694) );
  XOR U15173 ( .A(n9699), .B(n9321), .Z(n9323) );
  XOR U15174 ( .A(n9700), .B(n9701), .Z(n9321) );
  AND U15175 ( .A(n9702), .B(n9703), .Z(n9700) );
  AND U15176 ( .A(b[38]), .B(a[63]), .Z(n9699) );
  XOR U15177 ( .A(n9704), .B(n9326), .Z(n9328) );
  XOR U15178 ( .A(n9705), .B(n9706), .Z(n9326) );
  AND U15179 ( .A(n9707), .B(n9708), .Z(n9705) );
  AND U15180 ( .A(b[37]), .B(a[64]), .Z(n9704) );
  XOR U15181 ( .A(n9709), .B(n9331), .Z(n9333) );
  XOR U15182 ( .A(n9710), .B(n9711), .Z(n9331) );
  AND U15183 ( .A(n9712), .B(n9713), .Z(n9710) );
  AND U15184 ( .A(b[36]), .B(a[65]), .Z(n9709) );
  XOR U15185 ( .A(n9714), .B(n9336), .Z(n9338) );
  XOR U15186 ( .A(n9715), .B(n9716), .Z(n9336) );
  AND U15187 ( .A(n9717), .B(n9718), .Z(n9715) );
  AND U15188 ( .A(b[35]), .B(a[66]), .Z(n9714) );
  XOR U15189 ( .A(n9719), .B(n9341), .Z(n9343) );
  XOR U15190 ( .A(n9720), .B(n9721), .Z(n9341) );
  AND U15191 ( .A(n9722), .B(n9723), .Z(n9720) );
  AND U15192 ( .A(b[34]), .B(a[67]), .Z(n9719) );
  XOR U15193 ( .A(n9724), .B(n9346), .Z(n9348) );
  XOR U15194 ( .A(n9725), .B(n9726), .Z(n9346) );
  AND U15195 ( .A(n9727), .B(n9728), .Z(n9725) );
  AND U15196 ( .A(b[33]), .B(a[68]), .Z(n9724) );
  XNOR U15197 ( .A(n9729), .B(n9730), .Z(n9350) );
  ANDN U15198 ( .B(n9731), .A(n9732), .Z(n9729) );
  XOR U15199 ( .A(n9733), .B(n9355), .Z(n9357) );
  XOR U15200 ( .A(n9734), .B(n9735), .Z(n9355) );
  AND U15201 ( .A(n9736), .B(n9737), .Z(n9734) );
  AND U15202 ( .A(b[32]), .B(a[69]), .Z(n9733) );
  XOR U15203 ( .A(n9738), .B(n9360), .Z(n9362) );
  XOR U15204 ( .A(n9739), .B(n9740), .Z(n9360) );
  AND U15205 ( .A(n9741), .B(n9742), .Z(n9739) );
  AND U15206 ( .A(b[30]), .B(a[71]), .Z(n9738) );
  XOR U15207 ( .A(n9743), .B(n9365), .Z(n9367) );
  XOR U15208 ( .A(n9744), .B(n9745), .Z(n9365) );
  AND U15209 ( .A(n9746), .B(n9747), .Z(n9744) );
  AND U15210 ( .A(b[29]), .B(a[72]), .Z(n9743) );
  XOR U15211 ( .A(n9748), .B(n9370), .Z(n9372) );
  XOR U15212 ( .A(n9749), .B(n9750), .Z(n9370) );
  AND U15213 ( .A(n9751), .B(n9752), .Z(n9749) );
  AND U15214 ( .A(b[28]), .B(a[73]), .Z(n9748) );
  XOR U15215 ( .A(n9753), .B(n9375), .Z(n9377) );
  XOR U15216 ( .A(n9754), .B(n9755), .Z(n9375) );
  AND U15217 ( .A(n9756), .B(n9757), .Z(n9754) );
  AND U15218 ( .A(b[27]), .B(a[74]), .Z(n9753) );
  XNOR U15219 ( .A(n9758), .B(n9759), .Z(n9379) );
  ANDN U15220 ( .B(n9760), .A(n9761), .Z(n9758) );
  XOR U15221 ( .A(n9762), .B(n9384), .Z(n9386) );
  XOR U15222 ( .A(n9763), .B(n9764), .Z(n9384) );
  AND U15223 ( .A(n9765), .B(n9766), .Z(n9763) );
  AND U15224 ( .A(b[26]), .B(a[75]), .Z(n9762) );
  XOR U15225 ( .A(n9767), .B(n9389), .Z(n9391) );
  XOR U15226 ( .A(n9768), .B(n9769), .Z(n9389) );
  AND U15227 ( .A(n9770), .B(n9771), .Z(n9768) );
  AND U15228 ( .A(b[24]), .B(a[77]), .Z(n9767) );
  XOR U15229 ( .A(n9772), .B(n9394), .Z(n9396) );
  XOR U15230 ( .A(n9773), .B(n9774), .Z(n9394) );
  AND U15231 ( .A(n9775), .B(n9776), .Z(n9773) );
  AND U15232 ( .A(b[23]), .B(a[78]), .Z(n9772) );
  XOR U15233 ( .A(n9777), .B(n9399), .Z(n9401) );
  XOR U15234 ( .A(n9778), .B(n9779), .Z(n9399) );
  AND U15235 ( .A(n9780), .B(n9781), .Z(n9778) );
  AND U15236 ( .A(b[22]), .B(a[79]), .Z(n9777) );
  XOR U15237 ( .A(n9782), .B(n9404), .Z(n9406) );
  XOR U15238 ( .A(n9783), .B(n9784), .Z(n9404) );
  AND U15239 ( .A(n9785), .B(n9786), .Z(n9783) );
  AND U15240 ( .A(b[21]), .B(a[80]), .Z(n9782) );
  XNOR U15241 ( .A(n9787), .B(n9788), .Z(n9408) );
  ANDN U15242 ( .B(n9789), .A(n9790), .Z(n9787) );
  XOR U15243 ( .A(n9791), .B(n9413), .Z(n9415) );
  XOR U15244 ( .A(n9792), .B(n9793), .Z(n9413) );
  AND U15245 ( .A(n9794), .B(n9795), .Z(n9792) );
  AND U15246 ( .A(b[20]), .B(a[81]), .Z(n9791) );
  XOR U15247 ( .A(n9796), .B(n9418), .Z(n9420) );
  XOR U15248 ( .A(n9797), .B(n9798), .Z(n9418) );
  AND U15249 ( .A(n9799), .B(n9800), .Z(n9797) );
  AND U15250 ( .A(b[18]), .B(a[83]), .Z(n9796) );
  XOR U15251 ( .A(n9801), .B(n9423), .Z(n9425) );
  XOR U15252 ( .A(n9802), .B(n9803), .Z(n9423) );
  AND U15253 ( .A(n9804), .B(n9805), .Z(n9802) );
  AND U15254 ( .A(b[17]), .B(a[84]), .Z(n9801) );
  XOR U15255 ( .A(n9806), .B(n9428), .Z(n9430) );
  XOR U15256 ( .A(n9807), .B(n9808), .Z(n9428) );
  AND U15257 ( .A(n9809), .B(n9810), .Z(n9807) );
  AND U15258 ( .A(b[16]), .B(a[85]), .Z(n9806) );
  XOR U15259 ( .A(n9811), .B(n9433), .Z(n9435) );
  XOR U15260 ( .A(n9812), .B(n9813), .Z(n9433) );
  AND U15261 ( .A(n9814), .B(n9815), .Z(n9812) );
  AND U15262 ( .A(b[15]), .B(a[86]), .Z(n9811) );
  XNOR U15263 ( .A(n9816), .B(n9817), .Z(n9437) );
  ANDN U15264 ( .B(n9818), .A(n9819), .Z(n9816) );
  XOR U15265 ( .A(n9820), .B(n9442), .Z(n9444) );
  XOR U15266 ( .A(n9821), .B(n9822), .Z(n9442) );
  AND U15267 ( .A(n9823), .B(n9824), .Z(n9821) );
  AND U15268 ( .A(b[14]), .B(a[87]), .Z(n9820) );
  XOR U15269 ( .A(n9825), .B(n9447), .Z(n9449) );
  XOR U15270 ( .A(n9826), .B(n9827), .Z(n9447) );
  AND U15271 ( .A(n9828), .B(n9829), .Z(n9826) );
  AND U15272 ( .A(b[12]), .B(a[89]), .Z(n9825) );
  XOR U15273 ( .A(n9830), .B(n9452), .Z(n9454) );
  XOR U15274 ( .A(n9831), .B(n9832), .Z(n9452) );
  AND U15275 ( .A(n9833), .B(n9834), .Z(n9831) );
  AND U15276 ( .A(b[11]), .B(a[90]), .Z(n9830) );
  XOR U15277 ( .A(n9835), .B(n9457), .Z(n9459) );
  XOR U15278 ( .A(n9836), .B(n9837), .Z(n9457) );
  AND U15279 ( .A(n9838), .B(n9839), .Z(n9836) );
  AND U15280 ( .A(b[10]), .B(a[91]), .Z(n9835) );
  XOR U15281 ( .A(n9840), .B(n9462), .Z(n9464) );
  XOR U15282 ( .A(n9841), .B(n9842), .Z(n9462) );
  AND U15283 ( .A(n9843), .B(n9844), .Z(n9841) );
  AND U15284 ( .A(b[9]), .B(a[92]), .Z(n9840) );
  XNOR U15285 ( .A(n9845), .B(n9846), .Z(n9466) );
  ANDN U15286 ( .B(n9847), .A(n9848), .Z(n9845) );
  XOR U15287 ( .A(n9849), .B(n9471), .Z(n9473) );
  XOR U15288 ( .A(n9850), .B(n9851), .Z(n9471) );
  AND U15289 ( .A(n9852), .B(n9853), .Z(n9850) );
  AND U15290 ( .A(b[8]), .B(a[93]), .Z(n9849) );
  XOR U15291 ( .A(n9854), .B(n9476), .Z(n9478) );
  XOR U15292 ( .A(n9855), .B(n9856), .Z(n9476) );
  AND U15293 ( .A(n9857), .B(n9858), .Z(n9855) );
  AND U15294 ( .A(b[6]), .B(a[95]), .Z(n9854) );
  XOR U15295 ( .A(n9859), .B(n9481), .Z(n9483) );
  XOR U15296 ( .A(n9860), .B(n9861), .Z(n9481) );
  AND U15297 ( .A(n9862), .B(n9863), .Z(n9860) );
  AND U15298 ( .A(b[5]), .B(a[96]), .Z(n9859) );
  XOR U15299 ( .A(n9864), .B(n9486), .Z(n9488) );
  XOR U15300 ( .A(n9865), .B(n9866), .Z(n9486) );
  AND U15301 ( .A(n9867), .B(n9868), .Z(n9865) );
  AND U15302 ( .A(b[4]), .B(a[97]), .Z(n9864) );
  XNOR U15303 ( .A(n9869), .B(n9870), .Z(n9496) );
  NANDN U15304 ( .A(n9871), .B(n9872), .Z(n9870) );
  XOR U15305 ( .A(n9873), .B(n9491), .Z(n9493) );
  XNOR U15306 ( .A(n9874), .B(n9875), .Z(n9491) );
  AND U15307 ( .A(n9876), .B(n9877), .Z(n9874) );
  AND U15308 ( .A(b[3]), .B(a[98]), .Z(n9873) );
  NAND U15309 ( .A(a[101]), .B(b[0]), .Z(n9499) );
  XOR U15310 ( .A(n9878), .B(n9879), .Z(swire[100]) );
  XOR U15311 ( .A(n9513), .B(n9512), .Z(n9880) );
  XNOR U15312 ( .A(n9871), .B(n9872), .Z(n9512) );
  XOR U15313 ( .A(n9869), .B(n9881), .Z(n9872) );
  NAND U15314 ( .A(b[1]), .B(a[99]), .Z(n9881) );
  XOR U15315 ( .A(n9877), .B(n9882), .Z(n9871) );
  XOR U15316 ( .A(n9869), .B(n9876), .Z(n9882) );
  XNOR U15317 ( .A(n9883), .B(n9875), .Z(n9876) );
  AND U15318 ( .A(b[2]), .B(a[98]), .Z(n9883) );
  OR U15319 ( .A(n9884), .B(n9885), .Z(n9869) );
  XOR U15320 ( .A(n9875), .B(n9867), .Z(n9886) );
  XNOR U15321 ( .A(n9866), .B(n9862), .Z(n9887) );
  XNOR U15322 ( .A(n9861), .B(n9857), .Z(n9888) );
  XOR U15323 ( .A(n9889), .B(n9890), .Z(n9857) );
  XOR U15324 ( .A(n9847), .B(n9848), .Z(n9890) );
  XOR U15325 ( .A(n9891), .B(n9846), .Z(n9848) );
  AND U15326 ( .A(b[6]), .B(a[94]), .Z(n9891) );
  XOR U15327 ( .A(n9846), .B(n9852), .Z(n9892) );
  XNOR U15328 ( .A(n9851), .B(n9843), .Z(n9893) );
  XNOR U15329 ( .A(n9842), .B(n9838), .Z(n9894) );
  XNOR U15330 ( .A(n9837), .B(n9833), .Z(n9895) );
  XNOR U15331 ( .A(n9832), .B(n9828), .Z(n9896) );
  XOR U15332 ( .A(n9897), .B(n9898), .Z(n9828) );
  XOR U15333 ( .A(n9818), .B(n9819), .Z(n9898) );
  XOR U15334 ( .A(n9899), .B(n9817), .Z(n9819) );
  AND U15335 ( .A(b[12]), .B(a[88]), .Z(n9899) );
  XOR U15336 ( .A(n9817), .B(n9823), .Z(n9900) );
  XNOR U15337 ( .A(n9822), .B(n9814), .Z(n9901) );
  XNOR U15338 ( .A(n9813), .B(n9809), .Z(n9902) );
  XNOR U15339 ( .A(n9808), .B(n9804), .Z(n9903) );
  XNOR U15340 ( .A(n9803), .B(n9799), .Z(n9904) );
  XOR U15341 ( .A(n9905), .B(n9906), .Z(n9799) );
  XOR U15342 ( .A(n9789), .B(n9790), .Z(n9906) );
  XOR U15343 ( .A(n9907), .B(n9788), .Z(n9790) );
  AND U15344 ( .A(b[18]), .B(a[82]), .Z(n9907) );
  XOR U15345 ( .A(n9788), .B(n9794), .Z(n9908) );
  XNOR U15346 ( .A(n9793), .B(n9785), .Z(n9909) );
  XNOR U15347 ( .A(n9784), .B(n9780), .Z(n9910) );
  XNOR U15348 ( .A(n9779), .B(n9775), .Z(n9911) );
  XNOR U15349 ( .A(n9774), .B(n9770), .Z(n9912) );
  XOR U15350 ( .A(n9913), .B(n9914), .Z(n9770) );
  XOR U15351 ( .A(n9760), .B(n9761), .Z(n9914) );
  XOR U15352 ( .A(n9915), .B(n9759), .Z(n9761) );
  AND U15353 ( .A(b[24]), .B(a[76]), .Z(n9915) );
  XOR U15354 ( .A(n9759), .B(n9765), .Z(n9916) );
  XNOR U15355 ( .A(n9764), .B(n9756), .Z(n9917) );
  XNOR U15356 ( .A(n9755), .B(n9751), .Z(n9918) );
  XNOR U15357 ( .A(n9750), .B(n9746), .Z(n9919) );
  XNOR U15358 ( .A(n9745), .B(n9741), .Z(n9920) );
  XOR U15359 ( .A(n9921), .B(n9922), .Z(n9741) );
  XOR U15360 ( .A(n9731), .B(n9732), .Z(n9922) );
  XOR U15361 ( .A(n9923), .B(n9730), .Z(n9732) );
  AND U15362 ( .A(b[30]), .B(a[70]), .Z(n9923) );
  XOR U15363 ( .A(n9730), .B(n9736), .Z(n9924) );
  XNOR U15364 ( .A(n9735), .B(n9727), .Z(n9925) );
  XNOR U15365 ( .A(n9726), .B(n9722), .Z(n9926) );
  XNOR U15366 ( .A(n9721), .B(n9717), .Z(n9927) );
  XNOR U15367 ( .A(n9716), .B(n9712), .Z(n9928) );
  XNOR U15368 ( .A(n9711), .B(n9707), .Z(n9929) );
  XNOR U15369 ( .A(n9706), .B(n9702), .Z(n9930) );
  XNOR U15370 ( .A(n9701), .B(n9697), .Z(n9931) );
  XNOR U15371 ( .A(n9696), .B(n9692), .Z(n9932) );
  XNOR U15372 ( .A(n9691), .B(n9687), .Z(n9933) );
  XNOR U15373 ( .A(n9686), .B(n9682), .Z(n9934) );
  XNOR U15374 ( .A(n9681), .B(n9677), .Z(n9935) );
  XNOR U15375 ( .A(n9676), .B(n9672), .Z(n9936) );
  XNOR U15376 ( .A(n9671), .B(n9667), .Z(n9937) );
  XNOR U15377 ( .A(n9666), .B(n9662), .Z(n9938) );
  XNOR U15378 ( .A(n9661), .B(n9657), .Z(n9939) );
  XNOR U15379 ( .A(n9656), .B(n9652), .Z(n9940) );
  XNOR U15380 ( .A(n9651), .B(n9647), .Z(n9941) );
  XNOR U15381 ( .A(n9646), .B(n9642), .Z(n9942) );
  XNOR U15382 ( .A(n9641), .B(n9637), .Z(n9943) );
  XNOR U15383 ( .A(n9636), .B(n9632), .Z(n9944) );
  XNOR U15384 ( .A(n9631), .B(n9627), .Z(n9945) );
  XNOR U15385 ( .A(n9626), .B(n9622), .Z(n9946) );
  XNOR U15386 ( .A(n9621), .B(n9617), .Z(n9947) );
  XNOR U15387 ( .A(n9616), .B(n9612), .Z(n9948) );
  XNOR U15388 ( .A(n9611), .B(n9607), .Z(n9949) );
  XNOR U15389 ( .A(n9606), .B(n9602), .Z(n9950) );
  XNOR U15390 ( .A(n9601), .B(n9597), .Z(n9951) );
  XNOR U15391 ( .A(n9596), .B(n9592), .Z(n9952) );
  XOR U15392 ( .A(n9591), .B(n9588), .Z(n9953) );
  XOR U15393 ( .A(n9954), .B(n9955), .Z(n9588) );
  XOR U15394 ( .A(n9586), .B(n9956), .Z(n9955) );
  XNOR U15395 ( .A(n9957), .B(n9958), .Z(n9956) );
  XOR U15396 ( .A(n9959), .B(n9960), .Z(n9958) );
  NAND U15397 ( .A(a[38]), .B(b[62]), .Z(n9960) );
  AND U15398 ( .A(a[37]), .B(b[63]), .Z(n9959) );
  XNOR U15399 ( .A(n9961), .B(n9957), .Z(n9954) );
  XNOR U15400 ( .A(n9962), .B(n9963), .Z(n9957) );
  ANDN U15401 ( .B(n9964), .A(n9965), .Z(n9962) );
  AND U15402 ( .A(a[39]), .B(b[61]), .Z(n9961) );
  XOR U15403 ( .A(n9966), .B(n9586), .Z(n9587) );
  XOR U15404 ( .A(n9967), .B(n9968), .Z(n9586) );
  AND U15405 ( .A(n9969), .B(n9970), .Z(n9967) );
  AND U15406 ( .A(a[40]), .B(b[60]), .Z(n9966) );
  XOR U15407 ( .A(n9971), .B(n9591), .Z(n9593) );
  XOR U15408 ( .A(n9972), .B(n9973), .Z(n9591) );
  AND U15409 ( .A(n9974), .B(n9975), .Z(n9972) );
  AND U15410 ( .A(a[41]), .B(b[59]), .Z(n9971) );
  XOR U15411 ( .A(n9976), .B(n9596), .Z(n9598) );
  XOR U15412 ( .A(n9977), .B(n9978), .Z(n9596) );
  AND U15413 ( .A(n9979), .B(n9980), .Z(n9977) );
  AND U15414 ( .A(a[42]), .B(b[58]), .Z(n9976) );
  XOR U15415 ( .A(n9981), .B(n9601), .Z(n9603) );
  XOR U15416 ( .A(n9982), .B(n9983), .Z(n9601) );
  AND U15417 ( .A(n9984), .B(n9985), .Z(n9982) );
  AND U15418 ( .A(a[43]), .B(b[57]), .Z(n9981) );
  XOR U15419 ( .A(n9986), .B(n9606), .Z(n9608) );
  XOR U15420 ( .A(n9987), .B(n9988), .Z(n9606) );
  AND U15421 ( .A(n9989), .B(n9990), .Z(n9987) );
  AND U15422 ( .A(a[44]), .B(b[56]), .Z(n9986) );
  XOR U15423 ( .A(n9991), .B(n9611), .Z(n9613) );
  XOR U15424 ( .A(n9992), .B(n9993), .Z(n9611) );
  AND U15425 ( .A(n9994), .B(n9995), .Z(n9992) );
  AND U15426 ( .A(a[45]), .B(b[55]), .Z(n9991) );
  XOR U15427 ( .A(n9996), .B(n9616), .Z(n9618) );
  XOR U15428 ( .A(n9997), .B(n9998), .Z(n9616) );
  AND U15429 ( .A(n9999), .B(n10000), .Z(n9997) );
  AND U15430 ( .A(a[46]), .B(b[54]), .Z(n9996) );
  XOR U15431 ( .A(n10001), .B(n9621), .Z(n9623) );
  XOR U15432 ( .A(n10002), .B(n10003), .Z(n9621) );
  AND U15433 ( .A(n10004), .B(n10005), .Z(n10002) );
  AND U15434 ( .A(a[47]), .B(b[53]), .Z(n10001) );
  XOR U15435 ( .A(n10006), .B(n9626), .Z(n9628) );
  XOR U15436 ( .A(n10007), .B(n10008), .Z(n9626) );
  AND U15437 ( .A(n10009), .B(n10010), .Z(n10007) );
  AND U15438 ( .A(a[48]), .B(b[52]), .Z(n10006) );
  XOR U15439 ( .A(n10011), .B(n9631), .Z(n9633) );
  XOR U15440 ( .A(n10012), .B(n10013), .Z(n9631) );
  AND U15441 ( .A(n10014), .B(n10015), .Z(n10012) );
  AND U15442 ( .A(a[49]), .B(b[51]), .Z(n10011) );
  XOR U15443 ( .A(n10016), .B(n9636), .Z(n9638) );
  XOR U15444 ( .A(n10017), .B(n10018), .Z(n9636) );
  AND U15445 ( .A(n10019), .B(n10020), .Z(n10017) );
  AND U15446 ( .A(a[50]), .B(b[50]), .Z(n10016) );
  XOR U15447 ( .A(n10021), .B(n9641), .Z(n9643) );
  XOR U15448 ( .A(n10022), .B(n10023), .Z(n9641) );
  AND U15449 ( .A(n10024), .B(n10025), .Z(n10022) );
  AND U15450 ( .A(b[49]), .B(a[51]), .Z(n10021) );
  XOR U15451 ( .A(n10026), .B(n9646), .Z(n9648) );
  XOR U15452 ( .A(n10027), .B(n10028), .Z(n9646) );
  AND U15453 ( .A(n10029), .B(n10030), .Z(n10027) );
  AND U15454 ( .A(b[48]), .B(a[52]), .Z(n10026) );
  XOR U15455 ( .A(n10031), .B(n9651), .Z(n9653) );
  XOR U15456 ( .A(n10032), .B(n10033), .Z(n9651) );
  AND U15457 ( .A(n10034), .B(n10035), .Z(n10032) );
  AND U15458 ( .A(b[47]), .B(a[53]), .Z(n10031) );
  XOR U15459 ( .A(n10036), .B(n9656), .Z(n9658) );
  XOR U15460 ( .A(n10037), .B(n10038), .Z(n9656) );
  AND U15461 ( .A(n10039), .B(n10040), .Z(n10037) );
  AND U15462 ( .A(b[46]), .B(a[54]), .Z(n10036) );
  XOR U15463 ( .A(n10041), .B(n9661), .Z(n9663) );
  XOR U15464 ( .A(n10042), .B(n10043), .Z(n9661) );
  AND U15465 ( .A(n10044), .B(n10045), .Z(n10042) );
  AND U15466 ( .A(b[45]), .B(a[55]), .Z(n10041) );
  XOR U15467 ( .A(n10046), .B(n9666), .Z(n9668) );
  XOR U15468 ( .A(n10047), .B(n10048), .Z(n9666) );
  AND U15469 ( .A(n10049), .B(n10050), .Z(n10047) );
  AND U15470 ( .A(b[44]), .B(a[56]), .Z(n10046) );
  XOR U15471 ( .A(n10051), .B(n9671), .Z(n9673) );
  XOR U15472 ( .A(n10052), .B(n10053), .Z(n9671) );
  AND U15473 ( .A(n10054), .B(n10055), .Z(n10052) );
  AND U15474 ( .A(b[43]), .B(a[57]), .Z(n10051) );
  XOR U15475 ( .A(n10056), .B(n9676), .Z(n9678) );
  XOR U15476 ( .A(n10057), .B(n10058), .Z(n9676) );
  AND U15477 ( .A(n10059), .B(n10060), .Z(n10057) );
  AND U15478 ( .A(b[42]), .B(a[58]), .Z(n10056) );
  XOR U15479 ( .A(n10061), .B(n9681), .Z(n9683) );
  XOR U15480 ( .A(n10062), .B(n10063), .Z(n9681) );
  AND U15481 ( .A(n10064), .B(n10065), .Z(n10062) );
  AND U15482 ( .A(b[41]), .B(a[59]), .Z(n10061) );
  XOR U15483 ( .A(n10066), .B(n9686), .Z(n9688) );
  XOR U15484 ( .A(n10067), .B(n10068), .Z(n9686) );
  AND U15485 ( .A(n10069), .B(n10070), .Z(n10067) );
  AND U15486 ( .A(b[40]), .B(a[60]), .Z(n10066) );
  XOR U15487 ( .A(n10071), .B(n9691), .Z(n9693) );
  XOR U15488 ( .A(n10072), .B(n10073), .Z(n9691) );
  AND U15489 ( .A(n10074), .B(n10075), .Z(n10072) );
  AND U15490 ( .A(b[39]), .B(a[61]), .Z(n10071) );
  XOR U15491 ( .A(n10076), .B(n9696), .Z(n9698) );
  XOR U15492 ( .A(n10077), .B(n10078), .Z(n9696) );
  AND U15493 ( .A(n10079), .B(n10080), .Z(n10077) );
  AND U15494 ( .A(b[38]), .B(a[62]), .Z(n10076) );
  XOR U15495 ( .A(n10081), .B(n9701), .Z(n9703) );
  XOR U15496 ( .A(n10082), .B(n10083), .Z(n9701) );
  AND U15497 ( .A(n10084), .B(n10085), .Z(n10082) );
  AND U15498 ( .A(b[37]), .B(a[63]), .Z(n10081) );
  XOR U15499 ( .A(n10086), .B(n9706), .Z(n9708) );
  XOR U15500 ( .A(n10087), .B(n10088), .Z(n9706) );
  AND U15501 ( .A(n10089), .B(n10090), .Z(n10087) );
  AND U15502 ( .A(b[36]), .B(a[64]), .Z(n10086) );
  XOR U15503 ( .A(n10091), .B(n9711), .Z(n9713) );
  XOR U15504 ( .A(n10092), .B(n10093), .Z(n9711) );
  AND U15505 ( .A(n10094), .B(n10095), .Z(n10092) );
  AND U15506 ( .A(b[35]), .B(a[65]), .Z(n10091) );
  XOR U15507 ( .A(n10096), .B(n9716), .Z(n9718) );
  XOR U15508 ( .A(n10097), .B(n10098), .Z(n9716) );
  AND U15509 ( .A(n10099), .B(n10100), .Z(n10097) );
  AND U15510 ( .A(b[34]), .B(a[66]), .Z(n10096) );
  XOR U15511 ( .A(n10101), .B(n9721), .Z(n9723) );
  XOR U15512 ( .A(n10102), .B(n10103), .Z(n9721) );
  AND U15513 ( .A(n10104), .B(n10105), .Z(n10102) );
  AND U15514 ( .A(b[33]), .B(a[67]), .Z(n10101) );
  XOR U15515 ( .A(n10106), .B(n9726), .Z(n9728) );
  XOR U15516 ( .A(n10107), .B(n10108), .Z(n9726) );
  AND U15517 ( .A(n10109), .B(n10110), .Z(n10107) );
  AND U15518 ( .A(b[32]), .B(a[68]), .Z(n10106) );
  XNOR U15519 ( .A(n10111), .B(n10112), .Z(n9730) );
  AND U15520 ( .A(n10113), .B(n10114), .Z(n10111) );
  XOR U15521 ( .A(n10115), .B(n9735), .Z(n9737) );
  XOR U15522 ( .A(n10116), .B(n10117), .Z(n9735) );
  AND U15523 ( .A(n10118), .B(n10119), .Z(n10116) );
  AND U15524 ( .A(b[31]), .B(a[69]), .Z(n10115) );
  XOR U15525 ( .A(n10120), .B(n9740), .Z(n9742) );
  IV U15526 ( .A(n9921), .Z(n9740) );
  XOR U15527 ( .A(n10121), .B(n10122), .Z(n9921) );
  AND U15528 ( .A(n10123), .B(n10124), .Z(n10121) );
  AND U15529 ( .A(b[29]), .B(a[71]), .Z(n10120) );
  XOR U15530 ( .A(n10125), .B(n9745), .Z(n9747) );
  XOR U15531 ( .A(n10126), .B(n10127), .Z(n9745) );
  AND U15532 ( .A(n10128), .B(n10129), .Z(n10126) );
  AND U15533 ( .A(b[28]), .B(a[72]), .Z(n10125) );
  XOR U15534 ( .A(n10130), .B(n9750), .Z(n9752) );
  XOR U15535 ( .A(n10131), .B(n10132), .Z(n9750) );
  AND U15536 ( .A(n10133), .B(n10134), .Z(n10131) );
  AND U15537 ( .A(b[27]), .B(a[73]), .Z(n10130) );
  XOR U15538 ( .A(n10135), .B(n9755), .Z(n9757) );
  XOR U15539 ( .A(n10136), .B(n10137), .Z(n9755) );
  AND U15540 ( .A(n10138), .B(n10139), .Z(n10136) );
  AND U15541 ( .A(b[26]), .B(a[74]), .Z(n10135) );
  XNOR U15542 ( .A(n10140), .B(n10141), .Z(n9759) );
  AND U15543 ( .A(n10142), .B(n10143), .Z(n10140) );
  XOR U15544 ( .A(n10144), .B(n9764), .Z(n9766) );
  XOR U15545 ( .A(n10145), .B(n10146), .Z(n9764) );
  AND U15546 ( .A(n10147), .B(n10148), .Z(n10145) );
  AND U15547 ( .A(b[25]), .B(a[75]), .Z(n10144) );
  XOR U15548 ( .A(n10149), .B(n9769), .Z(n9771) );
  IV U15549 ( .A(n9913), .Z(n9769) );
  XOR U15550 ( .A(n10150), .B(n10151), .Z(n9913) );
  AND U15551 ( .A(n10152), .B(n10153), .Z(n10150) );
  AND U15552 ( .A(b[23]), .B(a[77]), .Z(n10149) );
  XOR U15553 ( .A(n10154), .B(n9774), .Z(n9776) );
  XOR U15554 ( .A(n10155), .B(n10156), .Z(n9774) );
  AND U15555 ( .A(n10157), .B(n10158), .Z(n10155) );
  AND U15556 ( .A(b[22]), .B(a[78]), .Z(n10154) );
  XOR U15557 ( .A(n10159), .B(n9779), .Z(n9781) );
  XOR U15558 ( .A(n10160), .B(n10161), .Z(n9779) );
  AND U15559 ( .A(n10162), .B(n10163), .Z(n10160) );
  AND U15560 ( .A(b[21]), .B(a[79]), .Z(n10159) );
  XOR U15561 ( .A(n10164), .B(n9784), .Z(n9786) );
  XOR U15562 ( .A(n10165), .B(n10166), .Z(n9784) );
  AND U15563 ( .A(n10167), .B(n10168), .Z(n10165) );
  AND U15564 ( .A(b[20]), .B(a[80]), .Z(n10164) );
  XNOR U15565 ( .A(n10169), .B(n10170), .Z(n9788) );
  AND U15566 ( .A(n10171), .B(n10172), .Z(n10169) );
  XOR U15567 ( .A(n10173), .B(n9793), .Z(n9795) );
  XOR U15568 ( .A(n10174), .B(n10175), .Z(n9793) );
  AND U15569 ( .A(n10176), .B(n10177), .Z(n10174) );
  AND U15570 ( .A(b[19]), .B(a[81]), .Z(n10173) );
  XOR U15571 ( .A(n10178), .B(n9798), .Z(n9800) );
  IV U15572 ( .A(n9905), .Z(n9798) );
  XOR U15573 ( .A(n10179), .B(n10180), .Z(n9905) );
  AND U15574 ( .A(n10181), .B(n10182), .Z(n10179) );
  AND U15575 ( .A(b[17]), .B(a[83]), .Z(n10178) );
  XOR U15576 ( .A(n10183), .B(n9803), .Z(n9805) );
  XOR U15577 ( .A(n10184), .B(n10185), .Z(n9803) );
  AND U15578 ( .A(n10186), .B(n10187), .Z(n10184) );
  AND U15579 ( .A(b[16]), .B(a[84]), .Z(n10183) );
  XOR U15580 ( .A(n10188), .B(n9808), .Z(n9810) );
  XOR U15581 ( .A(n10189), .B(n10190), .Z(n9808) );
  AND U15582 ( .A(n10191), .B(n10192), .Z(n10189) );
  AND U15583 ( .A(b[15]), .B(a[85]), .Z(n10188) );
  XOR U15584 ( .A(n10193), .B(n9813), .Z(n9815) );
  XOR U15585 ( .A(n10194), .B(n10195), .Z(n9813) );
  AND U15586 ( .A(n10196), .B(n10197), .Z(n10194) );
  AND U15587 ( .A(b[14]), .B(a[86]), .Z(n10193) );
  XNOR U15588 ( .A(n10198), .B(n10199), .Z(n9817) );
  AND U15589 ( .A(n10200), .B(n10201), .Z(n10198) );
  XOR U15590 ( .A(n10202), .B(n9822), .Z(n9824) );
  XOR U15591 ( .A(n10203), .B(n10204), .Z(n9822) );
  AND U15592 ( .A(n10205), .B(n10206), .Z(n10203) );
  AND U15593 ( .A(b[13]), .B(a[87]), .Z(n10202) );
  XOR U15594 ( .A(n10207), .B(n9827), .Z(n9829) );
  IV U15595 ( .A(n9897), .Z(n9827) );
  XOR U15596 ( .A(n10208), .B(n10209), .Z(n9897) );
  AND U15597 ( .A(n10210), .B(n10211), .Z(n10208) );
  AND U15598 ( .A(b[11]), .B(a[89]), .Z(n10207) );
  XOR U15599 ( .A(n10212), .B(n9832), .Z(n9834) );
  XOR U15600 ( .A(n10213), .B(n10214), .Z(n9832) );
  AND U15601 ( .A(n10215), .B(n10216), .Z(n10213) );
  AND U15602 ( .A(b[10]), .B(a[90]), .Z(n10212) );
  XOR U15603 ( .A(n10217), .B(n9837), .Z(n9839) );
  XOR U15604 ( .A(n10218), .B(n10219), .Z(n9837) );
  AND U15605 ( .A(n10220), .B(n10221), .Z(n10218) );
  AND U15606 ( .A(b[9]), .B(a[91]), .Z(n10217) );
  XOR U15607 ( .A(n10222), .B(n9842), .Z(n9844) );
  XOR U15608 ( .A(n10223), .B(n10224), .Z(n9842) );
  AND U15609 ( .A(n10225), .B(n10226), .Z(n10223) );
  AND U15610 ( .A(b[8]), .B(a[92]), .Z(n10222) );
  XNOR U15611 ( .A(n10227), .B(n10228), .Z(n9846) );
  AND U15612 ( .A(n10229), .B(n10230), .Z(n10227) );
  XOR U15613 ( .A(n10231), .B(n9851), .Z(n9853) );
  XOR U15614 ( .A(n10232), .B(n10233), .Z(n9851) );
  AND U15615 ( .A(n10234), .B(n10235), .Z(n10232) );
  AND U15616 ( .A(b[7]), .B(a[93]), .Z(n10231) );
  XOR U15617 ( .A(n10236), .B(n9856), .Z(n9858) );
  IV U15618 ( .A(n9889), .Z(n9856) );
  XOR U15619 ( .A(n10237), .B(n10238), .Z(n9889) );
  AND U15620 ( .A(n10239), .B(n10240), .Z(n10237) );
  AND U15621 ( .A(b[5]), .B(a[95]), .Z(n10236) );
  XOR U15622 ( .A(n10241), .B(n9861), .Z(n9863) );
  XOR U15623 ( .A(n10242), .B(n10243), .Z(n9861) );
  AND U15624 ( .A(n10244), .B(n10245), .Z(n10242) );
  AND U15625 ( .A(b[4]), .B(a[96]), .Z(n10241) );
  XNOR U15626 ( .A(n10246), .B(n10247), .Z(n9875) );
  NANDN U15627 ( .A(n10248), .B(n10249), .Z(n10247) );
  XOR U15628 ( .A(n10250), .B(n9866), .Z(n9868) );
  XOR U15629 ( .A(n10251), .B(n10252), .Z(n9866) );
  AND U15630 ( .A(n10253), .B(n10254), .Z(n10251) );
  AND U15631 ( .A(b[3]), .B(a[97]), .Z(n10250) );
  NAND U15632 ( .A(a[100]), .B(b[0]), .Z(n9513) );
  XOR U15633 ( .A(n9885), .B(n10255), .Z(n2) );
  XNOR U15634 ( .A(n9884), .B(n1), .Z(n10255) );
  XOR U15635 ( .A(n10257), .B(n10258), .Z(n4) );
  XNOR U15636 ( .A(n10259), .B(n10256), .Z(n10258) );
  IV U15637 ( .A(n3), .Z(n10256) );
  XNOR U15638 ( .A(n10260), .B(n10261), .Z(n6) );
  XOR U15639 ( .A(n10263), .B(n10264), .Z(n8) );
  XOR U15640 ( .A(n10266), .B(n10267), .Z(n10) );
  XOR U15641 ( .A(n10269), .B(n10270), .Z(n12) );
  XOR U15642 ( .A(n10272), .B(n10273), .Z(n14) );
  XOR U15643 ( .A(n10275), .B(n10276), .Z(n16) );
  XOR U15644 ( .A(n10278), .B(n10279), .Z(n18) );
  XOR U15645 ( .A(n10281), .B(n10282), .Z(n20) );
  XOR U15646 ( .A(n10284), .B(n10285), .Z(n22) );
  XOR U15647 ( .A(n10287), .B(n10288), .Z(n24) );
  XOR U15648 ( .A(n10290), .B(n10291), .Z(n26) );
  XOR U15649 ( .A(n10293), .B(n10294), .Z(n28) );
  XOR U15650 ( .A(n10296), .B(n10297), .Z(n30) );
  XOR U15651 ( .A(n10299), .B(n10300), .Z(n32) );
  XOR U15652 ( .A(n10302), .B(n10303), .Z(n34) );
  XOR U15653 ( .A(n10305), .B(n10306), .Z(n36) );
  XOR U15654 ( .A(n10308), .B(n10309), .Z(n38) );
  XOR U15655 ( .A(n10311), .B(n10312), .Z(n40) );
  XOR U15656 ( .A(n10314), .B(n10315), .Z(n42) );
  XOR U15657 ( .A(n10317), .B(n10318), .Z(n44) );
  XOR U15658 ( .A(n10320), .B(n10321), .Z(n46) );
  XOR U15659 ( .A(n10323), .B(n10324), .Z(n48) );
  XOR U15660 ( .A(n10326), .B(n10327), .Z(n50) );
  XOR U15661 ( .A(n10329), .B(n10330), .Z(n52) );
  XOR U15662 ( .A(n10332), .B(n10333), .Z(n54) );
  XOR U15663 ( .A(n10335), .B(n10336), .Z(n56) );
  XOR U15664 ( .A(n10338), .B(n10339), .Z(n58) );
  XOR U15665 ( .A(n10341), .B(n10342), .Z(n60) );
  XOR U15666 ( .A(n10344), .B(n10345), .Z(n62) );
  XOR U15667 ( .A(n10347), .B(n10348), .Z(n64) );
  XOR U15668 ( .A(n10350), .B(n10351), .Z(n66) );
  XOR U15669 ( .A(n10353), .B(n10354), .Z(n68) );
  XOR U15670 ( .A(n10356), .B(n10357), .Z(n70) );
  XOR U15671 ( .A(n10359), .B(n10360), .Z(n72) );
  XOR U15672 ( .A(n10361), .B(n71), .Z(n10360) );
  XNOR U15673 ( .A(n10362), .B(n10363), .Z(n71) );
  NOR U15674 ( .A(n10364), .B(n10365), .Z(n10362) );
  NAND U15675 ( .A(a[99]), .B(b[0]), .Z(n9884) );
  XOR U15676 ( .A(n10249), .B(n10248), .Z(n9885) );
  XOR U15677 ( .A(n10246), .B(n10253), .Z(n10366) );
  XOR U15678 ( .A(n10244), .B(n10368), .Z(n10367) );
  XOR U15679 ( .A(n10239), .B(n10370), .Z(n10369) );
  XOR U15680 ( .A(n10229), .B(n10238), .Z(n10371) );
  XOR U15681 ( .A(n10234), .B(n10373), .Z(n10372) );
  XOR U15682 ( .A(n10225), .B(n10375), .Z(n10374) );
  XOR U15683 ( .A(n10220), .B(n10377), .Z(n10376) );
  XOR U15684 ( .A(n10215), .B(n10379), .Z(n10378) );
  XOR U15685 ( .A(n10210), .B(n10381), .Z(n10380) );
  XOR U15686 ( .A(n10200), .B(n10209), .Z(n10382) );
  XOR U15687 ( .A(n10205), .B(n10384), .Z(n10383) );
  XOR U15688 ( .A(n10196), .B(n10386), .Z(n10385) );
  XOR U15689 ( .A(n10191), .B(n10388), .Z(n10387) );
  XOR U15690 ( .A(n10186), .B(n10390), .Z(n10389) );
  XOR U15691 ( .A(n10181), .B(n10392), .Z(n10391) );
  XOR U15692 ( .A(n10171), .B(n10180), .Z(n10393) );
  XOR U15693 ( .A(n10176), .B(n10395), .Z(n10394) );
  XOR U15694 ( .A(n10167), .B(n10397), .Z(n10396) );
  XOR U15695 ( .A(n10162), .B(n10399), .Z(n10398) );
  XOR U15696 ( .A(n10157), .B(n10401), .Z(n10400) );
  XOR U15697 ( .A(n10152), .B(n10403), .Z(n10402) );
  XOR U15698 ( .A(n10142), .B(n10151), .Z(n10404) );
  XOR U15699 ( .A(n10147), .B(n10406), .Z(n10405) );
  XOR U15700 ( .A(n10138), .B(n10408), .Z(n10407) );
  XOR U15701 ( .A(n10133), .B(n10410), .Z(n10409) );
  XOR U15702 ( .A(n10128), .B(n10412), .Z(n10411) );
  XOR U15703 ( .A(n10123), .B(n10414), .Z(n10413) );
  XOR U15704 ( .A(n10113), .B(n10122), .Z(n10415) );
  XOR U15705 ( .A(n10118), .B(n10417), .Z(n10416) );
  XOR U15706 ( .A(n10109), .B(n10419), .Z(n10418) );
  XOR U15707 ( .A(n10104), .B(n10421), .Z(n10420) );
  XOR U15708 ( .A(n10099), .B(n10423), .Z(n10422) );
  XOR U15709 ( .A(n10094), .B(n10425), .Z(n10424) );
  XOR U15710 ( .A(n10089), .B(n10427), .Z(n10426) );
  XOR U15711 ( .A(n10084), .B(n10429), .Z(n10428) );
  XOR U15712 ( .A(n10079), .B(n10431), .Z(n10430) );
  XOR U15713 ( .A(n10074), .B(n10433), .Z(n10432) );
  XOR U15714 ( .A(n10069), .B(n10435), .Z(n10434) );
  XOR U15715 ( .A(n10064), .B(n10437), .Z(n10436) );
  XOR U15716 ( .A(n10059), .B(n10439), .Z(n10438) );
  XOR U15717 ( .A(n10054), .B(n10441), .Z(n10440) );
  XOR U15718 ( .A(n10049), .B(n10443), .Z(n10442) );
  XOR U15719 ( .A(n10044), .B(n10445), .Z(n10444) );
  XOR U15720 ( .A(n10039), .B(n10447), .Z(n10446) );
  XOR U15721 ( .A(n10034), .B(n10449), .Z(n10448) );
  XOR U15722 ( .A(n10029), .B(n10451), .Z(n10450) );
  XOR U15723 ( .A(n10024), .B(n10453), .Z(n10452) );
  XOR U15724 ( .A(n10019), .B(n10455), .Z(n10454) );
  XOR U15725 ( .A(n10014), .B(n10457), .Z(n10456) );
  XOR U15726 ( .A(n10009), .B(n10459), .Z(n10458) );
  XOR U15727 ( .A(n10004), .B(n10461), .Z(n10460) );
  XOR U15728 ( .A(n9999), .B(n10463), .Z(n10462) );
  XOR U15729 ( .A(n9994), .B(n10465), .Z(n10464) );
  XOR U15730 ( .A(n9989), .B(n10467), .Z(n10466) );
  XOR U15731 ( .A(n9984), .B(n10469), .Z(n10468) );
  XOR U15732 ( .A(n9979), .B(n10471), .Z(n10470) );
  XOR U15733 ( .A(n9974), .B(n10473), .Z(n10472) );
  XOR U15734 ( .A(n9969), .B(n10475), .Z(n10474) );
  XNOR U15735 ( .A(n9965), .B(n10477), .Z(n10476) );
  XOR U15736 ( .A(n10478), .B(n10479), .Z(n9965) );
  XOR U15737 ( .A(n10480), .B(n10481), .Z(n10479) );
  XNOR U15738 ( .A(n10482), .B(n10483), .Z(n10480) );
  XOR U15739 ( .A(n10484), .B(n10485), .Z(n10483) );
  AND U15740 ( .A(a[36]), .B(b[63]), .Z(n10485) );
  AND U15741 ( .A(a[37]), .B(b[62]), .Z(n10484) );
  XNOR U15742 ( .A(n10486), .B(n10482), .Z(n10478) );
  XNOR U15743 ( .A(n10487), .B(n10488), .Z(n10482) );
  ANDN U15744 ( .B(n10489), .A(n10490), .Z(n10487) );
  AND U15745 ( .A(a[38]), .B(b[61]), .Z(n10486) );
  XOR U15746 ( .A(n10491), .B(n9963), .Z(n9964) );
  IV U15747 ( .A(n10481), .Z(n9963) );
  XOR U15748 ( .A(n10492), .B(n10493), .Z(n10481) );
  AND U15749 ( .A(n10494), .B(n10495), .Z(n10492) );
  AND U15750 ( .A(a[39]), .B(b[60]), .Z(n10491) );
  XOR U15751 ( .A(n10496), .B(n9968), .Z(n9970) );
  IV U15752 ( .A(n10477), .Z(n9968) );
  XOR U15753 ( .A(n10497), .B(n10498), .Z(n10477) );
  AND U15754 ( .A(n10499), .B(n10500), .Z(n10497) );
  AND U15755 ( .A(a[40]), .B(b[59]), .Z(n10496) );
  XOR U15756 ( .A(n10501), .B(n9973), .Z(n9975) );
  IV U15757 ( .A(n10475), .Z(n9973) );
  XOR U15758 ( .A(n10502), .B(n10503), .Z(n10475) );
  AND U15759 ( .A(n10504), .B(n10505), .Z(n10502) );
  AND U15760 ( .A(a[41]), .B(b[58]), .Z(n10501) );
  XOR U15761 ( .A(n10506), .B(n9978), .Z(n9980) );
  IV U15762 ( .A(n10473), .Z(n9978) );
  XOR U15763 ( .A(n10507), .B(n10508), .Z(n10473) );
  AND U15764 ( .A(n10509), .B(n10510), .Z(n10507) );
  AND U15765 ( .A(a[42]), .B(b[57]), .Z(n10506) );
  XOR U15766 ( .A(n10511), .B(n9983), .Z(n9985) );
  IV U15767 ( .A(n10471), .Z(n9983) );
  XOR U15768 ( .A(n10512), .B(n10513), .Z(n10471) );
  AND U15769 ( .A(n10514), .B(n10515), .Z(n10512) );
  AND U15770 ( .A(a[43]), .B(b[56]), .Z(n10511) );
  XOR U15771 ( .A(n10516), .B(n9988), .Z(n9990) );
  IV U15772 ( .A(n10469), .Z(n9988) );
  XOR U15773 ( .A(n10517), .B(n10518), .Z(n10469) );
  AND U15774 ( .A(n10519), .B(n10520), .Z(n10517) );
  AND U15775 ( .A(a[44]), .B(b[55]), .Z(n10516) );
  XOR U15776 ( .A(n10521), .B(n9993), .Z(n9995) );
  IV U15777 ( .A(n10467), .Z(n9993) );
  XOR U15778 ( .A(n10522), .B(n10523), .Z(n10467) );
  AND U15779 ( .A(n10524), .B(n10525), .Z(n10522) );
  AND U15780 ( .A(a[45]), .B(b[54]), .Z(n10521) );
  XOR U15781 ( .A(n10526), .B(n9998), .Z(n10000) );
  IV U15782 ( .A(n10465), .Z(n9998) );
  XOR U15783 ( .A(n10527), .B(n10528), .Z(n10465) );
  AND U15784 ( .A(n10529), .B(n10530), .Z(n10527) );
  AND U15785 ( .A(a[46]), .B(b[53]), .Z(n10526) );
  XOR U15786 ( .A(n10531), .B(n10003), .Z(n10005) );
  IV U15787 ( .A(n10463), .Z(n10003) );
  XOR U15788 ( .A(n10532), .B(n10533), .Z(n10463) );
  AND U15789 ( .A(n10534), .B(n10535), .Z(n10532) );
  AND U15790 ( .A(a[47]), .B(b[52]), .Z(n10531) );
  XOR U15791 ( .A(n10536), .B(n10008), .Z(n10010) );
  IV U15792 ( .A(n10461), .Z(n10008) );
  XOR U15793 ( .A(n10537), .B(n10538), .Z(n10461) );
  AND U15794 ( .A(n10539), .B(n10540), .Z(n10537) );
  AND U15795 ( .A(a[48]), .B(b[51]), .Z(n10536) );
  XOR U15796 ( .A(n10541), .B(n10013), .Z(n10015) );
  IV U15797 ( .A(n10459), .Z(n10013) );
  XOR U15798 ( .A(n10542), .B(n10543), .Z(n10459) );
  AND U15799 ( .A(n10544), .B(n10545), .Z(n10542) );
  AND U15800 ( .A(a[49]), .B(b[50]), .Z(n10541) );
  XOR U15801 ( .A(n10546), .B(n10018), .Z(n10020) );
  IV U15802 ( .A(n10457), .Z(n10018) );
  XOR U15803 ( .A(n10547), .B(n10548), .Z(n10457) );
  AND U15804 ( .A(n10549), .B(n10550), .Z(n10547) );
  AND U15805 ( .A(b[49]), .B(a[50]), .Z(n10546) );
  XOR U15806 ( .A(n10551), .B(n10023), .Z(n10025) );
  IV U15807 ( .A(n10455), .Z(n10023) );
  XOR U15808 ( .A(n10552), .B(n10553), .Z(n10455) );
  AND U15809 ( .A(n10554), .B(n10555), .Z(n10552) );
  AND U15810 ( .A(b[48]), .B(a[51]), .Z(n10551) );
  XOR U15811 ( .A(n10556), .B(n10028), .Z(n10030) );
  IV U15812 ( .A(n10453), .Z(n10028) );
  XOR U15813 ( .A(n10557), .B(n10558), .Z(n10453) );
  AND U15814 ( .A(n10559), .B(n10560), .Z(n10557) );
  AND U15815 ( .A(b[47]), .B(a[52]), .Z(n10556) );
  XOR U15816 ( .A(n10561), .B(n10033), .Z(n10035) );
  IV U15817 ( .A(n10451), .Z(n10033) );
  XOR U15818 ( .A(n10562), .B(n10563), .Z(n10451) );
  AND U15819 ( .A(n10564), .B(n10565), .Z(n10562) );
  AND U15820 ( .A(b[46]), .B(a[53]), .Z(n10561) );
  XOR U15821 ( .A(n10566), .B(n10038), .Z(n10040) );
  IV U15822 ( .A(n10449), .Z(n10038) );
  XOR U15823 ( .A(n10567), .B(n10568), .Z(n10449) );
  AND U15824 ( .A(n10569), .B(n10570), .Z(n10567) );
  AND U15825 ( .A(b[45]), .B(a[54]), .Z(n10566) );
  XOR U15826 ( .A(n10571), .B(n10043), .Z(n10045) );
  IV U15827 ( .A(n10447), .Z(n10043) );
  XOR U15828 ( .A(n10572), .B(n10573), .Z(n10447) );
  AND U15829 ( .A(n10574), .B(n10575), .Z(n10572) );
  AND U15830 ( .A(b[44]), .B(a[55]), .Z(n10571) );
  XOR U15831 ( .A(n10576), .B(n10048), .Z(n10050) );
  IV U15832 ( .A(n10445), .Z(n10048) );
  XOR U15833 ( .A(n10577), .B(n10578), .Z(n10445) );
  AND U15834 ( .A(n10579), .B(n10580), .Z(n10577) );
  AND U15835 ( .A(b[43]), .B(a[56]), .Z(n10576) );
  XOR U15836 ( .A(n10581), .B(n10053), .Z(n10055) );
  IV U15837 ( .A(n10443), .Z(n10053) );
  XOR U15838 ( .A(n10582), .B(n10583), .Z(n10443) );
  AND U15839 ( .A(n10584), .B(n10585), .Z(n10582) );
  AND U15840 ( .A(b[42]), .B(a[57]), .Z(n10581) );
  XOR U15841 ( .A(n10586), .B(n10058), .Z(n10060) );
  IV U15842 ( .A(n10441), .Z(n10058) );
  XOR U15843 ( .A(n10587), .B(n10588), .Z(n10441) );
  AND U15844 ( .A(n10589), .B(n10590), .Z(n10587) );
  AND U15845 ( .A(b[41]), .B(a[58]), .Z(n10586) );
  XOR U15846 ( .A(n10591), .B(n10063), .Z(n10065) );
  IV U15847 ( .A(n10439), .Z(n10063) );
  XOR U15848 ( .A(n10592), .B(n10593), .Z(n10439) );
  AND U15849 ( .A(n10594), .B(n10595), .Z(n10592) );
  AND U15850 ( .A(b[40]), .B(a[59]), .Z(n10591) );
  XOR U15851 ( .A(n10596), .B(n10068), .Z(n10070) );
  IV U15852 ( .A(n10437), .Z(n10068) );
  XOR U15853 ( .A(n10597), .B(n10598), .Z(n10437) );
  AND U15854 ( .A(n10599), .B(n10600), .Z(n10597) );
  AND U15855 ( .A(b[39]), .B(a[60]), .Z(n10596) );
  XOR U15856 ( .A(n10601), .B(n10073), .Z(n10075) );
  IV U15857 ( .A(n10435), .Z(n10073) );
  XOR U15858 ( .A(n10602), .B(n10603), .Z(n10435) );
  AND U15859 ( .A(n10604), .B(n10605), .Z(n10602) );
  AND U15860 ( .A(b[38]), .B(a[61]), .Z(n10601) );
  XOR U15861 ( .A(n10606), .B(n10078), .Z(n10080) );
  IV U15862 ( .A(n10433), .Z(n10078) );
  XOR U15863 ( .A(n10607), .B(n10608), .Z(n10433) );
  AND U15864 ( .A(n10609), .B(n10610), .Z(n10607) );
  AND U15865 ( .A(b[37]), .B(a[62]), .Z(n10606) );
  XOR U15866 ( .A(n10611), .B(n10083), .Z(n10085) );
  IV U15867 ( .A(n10431), .Z(n10083) );
  XOR U15868 ( .A(n10612), .B(n10613), .Z(n10431) );
  AND U15869 ( .A(n10614), .B(n10615), .Z(n10612) );
  AND U15870 ( .A(b[36]), .B(a[63]), .Z(n10611) );
  XOR U15871 ( .A(n10616), .B(n10088), .Z(n10090) );
  IV U15872 ( .A(n10429), .Z(n10088) );
  XOR U15873 ( .A(n10617), .B(n10618), .Z(n10429) );
  AND U15874 ( .A(n10619), .B(n10620), .Z(n10617) );
  AND U15875 ( .A(b[35]), .B(a[64]), .Z(n10616) );
  XOR U15876 ( .A(n10621), .B(n10093), .Z(n10095) );
  IV U15877 ( .A(n10427), .Z(n10093) );
  XOR U15878 ( .A(n10622), .B(n10623), .Z(n10427) );
  AND U15879 ( .A(n10624), .B(n10625), .Z(n10622) );
  AND U15880 ( .A(b[34]), .B(a[65]), .Z(n10621) );
  XOR U15881 ( .A(n10626), .B(n10098), .Z(n10100) );
  IV U15882 ( .A(n10425), .Z(n10098) );
  XOR U15883 ( .A(n10627), .B(n10628), .Z(n10425) );
  AND U15884 ( .A(n10629), .B(n10630), .Z(n10627) );
  AND U15885 ( .A(b[33]), .B(a[66]), .Z(n10626) );
  XOR U15886 ( .A(n10631), .B(n10103), .Z(n10105) );
  IV U15887 ( .A(n10423), .Z(n10103) );
  XOR U15888 ( .A(n10632), .B(n10633), .Z(n10423) );
  AND U15889 ( .A(n10634), .B(n10635), .Z(n10632) );
  AND U15890 ( .A(b[32]), .B(a[67]), .Z(n10631) );
  XOR U15891 ( .A(n10636), .B(n10108), .Z(n10110) );
  IV U15892 ( .A(n10421), .Z(n10108) );
  XOR U15893 ( .A(n10637), .B(n10638), .Z(n10421) );
  AND U15894 ( .A(n10639), .B(n10640), .Z(n10637) );
  AND U15895 ( .A(b[31]), .B(a[68]), .Z(n10636) );
  XOR U15896 ( .A(n10641), .B(n10117), .Z(n10119) );
  IV U15897 ( .A(n10419), .Z(n10117) );
  XOR U15898 ( .A(n10642), .B(n10643), .Z(n10419) );
  AND U15899 ( .A(n10644), .B(n10645), .Z(n10642) );
  AND U15900 ( .A(b[30]), .B(a[69]), .Z(n10641) );
  XOR U15901 ( .A(n10646), .B(n10112), .Z(n10114) );
  IV U15902 ( .A(n10417), .Z(n10112) );
  XOR U15903 ( .A(n10647), .B(n10648), .Z(n10417) );
  AND U15904 ( .A(n10649), .B(n10650), .Z(n10647) );
  AND U15905 ( .A(b[29]), .B(a[70]), .Z(n10646) );
  XOR U15906 ( .A(n10652), .B(n10653), .Z(n10122) );
  AND U15907 ( .A(n10654), .B(n10655), .Z(n10652) );
  AND U15908 ( .A(b[28]), .B(a[71]), .Z(n10651) );
  XOR U15909 ( .A(n10656), .B(n10127), .Z(n10129) );
  IV U15910 ( .A(n10414), .Z(n10127) );
  XOR U15911 ( .A(n10657), .B(n10658), .Z(n10414) );
  AND U15912 ( .A(n10659), .B(n10660), .Z(n10657) );
  AND U15913 ( .A(b[27]), .B(a[72]), .Z(n10656) );
  XOR U15914 ( .A(n10661), .B(n10132), .Z(n10134) );
  IV U15915 ( .A(n10412), .Z(n10132) );
  XOR U15916 ( .A(n10662), .B(n10663), .Z(n10412) );
  AND U15917 ( .A(n10664), .B(n10665), .Z(n10662) );
  AND U15918 ( .A(b[26]), .B(a[73]), .Z(n10661) );
  XOR U15919 ( .A(n10666), .B(n10137), .Z(n10139) );
  IV U15920 ( .A(n10410), .Z(n10137) );
  XOR U15921 ( .A(n10667), .B(n10668), .Z(n10410) );
  AND U15922 ( .A(n10669), .B(n10670), .Z(n10667) );
  AND U15923 ( .A(b[25]), .B(a[74]), .Z(n10666) );
  XOR U15924 ( .A(n10671), .B(n10146), .Z(n10148) );
  IV U15925 ( .A(n10408), .Z(n10146) );
  XOR U15926 ( .A(n10672), .B(n10673), .Z(n10408) );
  AND U15927 ( .A(n10674), .B(n10675), .Z(n10672) );
  AND U15928 ( .A(b[24]), .B(a[75]), .Z(n10671) );
  XOR U15929 ( .A(n10676), .B(n10141), .Z(n10143) );
  IV U15930 ( .A(n10406), .Z(n10141) );
  XOR U15931 ( .A(n10677), .B(n10678), .Z(n10406) );
  AND U15932 ( .A(n10679), .B(n10680), .Z(n10677) );
  AND U15933 ( .A(b[23]), .B(a[76]), .Z(n10676) );
  XOR U15934 ( .A(n10682), .B(n10683), .Z(n10151) );
  AND U15935 ( .A(n10684), .B(n10685), .Z(n10682) );
  AND U15936 ( .A(b[22]), .B(a[77]), .Z(n10681) );
  XOR U15937 ( .A(n10686), .B(n10156), .Z(n10158) );
  IV U15938 ( .A(n10403), .Z(n10156) );
  XOR U15939 ( .A(n10687), .B(n10688), .Z(n10403) );
  AND U15940 ( .A(n10689), .B(n10690), .Z(n10687) );
  AND U15941 ( .A(b[21]), .B(a[78]), .Z(n10686) );
  XOR U15942 ( .A(n10691), .B(n10161), .Z(n10163) );
  IV U15943 ( .A(n10401), .Z(n10161) );
  XOR U15944 ( .A(n10692), .B(n10693), .Z(n10401) );
  AND U15945 ( .A(n10694), .B(n10695), .Z(n10692) );
  AND U15946 ( .A(b[20]), .B(a[79]), .Z(n10691) );
  XOR U15947 ( .A(n10696), .B(n10166), .Z(n10168) );
  IV U15948 ( .A(n10399), .Z(n10166) );
  XOR U15949 ( .A(n10697), .B(n10698), .Z(n10399) );
  AND U15950 ( .A(n10699), .B(n10700), .Z(n10697) );
  AND U15951 ( .A(b[19]), .B(a[80]), .Z(n10696) );
  XOR U15952 ( .A(n10701), .B(n10175), .Z(n10177) );
  IV U15953 ( .A(n10397), .Z(n10175) );
  XOR U15954 ( .A(n10702), .B(n10703), .Z(n10397) );
  AND U15955 ( .A(n10704), .B(n10705), .Z(n10702) );
  AND U15956 ( .A(b[18]), .B(a[81]), .Z(n10701) );
  XOR U15957 ( .A(n10706), .B(n10170), .Z(n10172) );
  IV U15958 ( .A(n10395), .Z(n10170) );
  XOR U15959 ( .A(n10707), .B(n10708), .Z(n10395) );
  AND U15960 ( .A(n10709), .B(n10710), .Z(n10707) );
  AND U15961 ( .A(b[17]), .B(a[82]), .Z(n10706) );
  XOR U15962 ( .A(n10712), .B(n10713), .Z(n10180) );
  AND U15963 ( .A(n10714), .B(n10715), .Z(n10712) );
  AND U15964 ( .A(b[16]), .B(a[83]), .Z(n10711) );
  XOR U15965 ( .A(n10716), .B(n10185), .Z(n10187) );
  IV U15966 ( .A(n10392), .Z(n10185) );
  XOR U15967 ( .A(n10717), .B(n10718), .Z(n10392) );
  AND U15968 ( .A(n10719), .B(n10720), .Z(n10717) );
  AND U15969 ( .A(b[15]), .B(a[84]), .Z(n10716) );
  XOR U15970 ( .A(n10721), .B(n10190), .Z(n10192) );
  IV U15971 ( .A(n10390), .Z(n10190) );
  XOR U15972 ( .A(n10722), .B(n10723), .Z(n10390) );
  AND U15973 ( .A(n10724), .B(n10725), .Z(n10722) );
  AND U15974 ( .A(b[14]), .B(a[85]), .Z(n10721) );
  XOR U15975 ( .A(n10726), .B(n10195), .Z(n10197) );
  IV U15976 ( .A(n10388), .Z(n10195) );
  XOR U15977 ( .A(n10727), .B(n10728), .Z(n10388) );
  AND U15978 ( .A(n10729), .B(n10730), .Z(n10727) );
  AND U15979 ( .A(b[13]), .B(a[86]), .Z(n10726) );
  XOR U15980 ( .A(n10731), .B(n10204), .Z(n10206) );
  IV U15981 ( .A(n10386), .Z(n10204) );
  XOR U15982 ( .A(n10732), .B(n10733), .Z(n10386) );
  AND U15983 ( .A(n10734), .B(n10735), .Z(n10732) );
  AND U15984 ( .A(b[12]), .B(a[87]), .Z(n10731) );
  XOR U15985 ( .A(n10736), .B(n10199), .Z(n10201) );
  IV U15986 ( .A(n10384), .Z(n10199) );
  XOR U15987 ( .A(n10737), .B(n10738), .Z(n10384) );
  AND U15988 ( .A(n10739), .B(n10740), .Z(n10737) );
  AND U15989 ( .A(b[11]), .B(a[88]), .Z(n10736) );
  XOR U15990 ( .A(n10742), .B(n10743), .Z(n10209) );
  AND U15991 ( .A(n10744), .B(n10745), .Z(n10742) );
  AND U15992 ( .A(b[10]), .B(a[89]), .Z(n10741) );
  XOR U15993 ( .A(n10746), .B(n10214), .Z(n10216) );
  IV U15994 ( .A(n10381), .Z(n10214) );
  XOR U15995 ( .A(n10747), .B(n10748), .Z(n10381) );
  AND U15996 ( .A(n10749), .B(n10750), .Z(n10747) );
  AND U15997 ( .A(b[9]), .B(a[90]), .Z(n10746) );
  XOR U15998 ( .A(n10751), .B(n10219), .Z(n10221) );
  IV U15999 ( .A(n10379), .Z(n10219) );
  XOR U16000 ( .A(n10752), .B(n10753), .Z(n10379) );
  AND U16001 ( .A(n10754), .B(n10755), .Z(n10752) );
  AND U16002 ( .A(b[8]), .B(a[91]), .Z(n10751) );
  XOR U16003 ( .A(n10756), .B(n10224), .Z(n10226) );
  IV U16004 ( .A(n10377), .Z(n10224) );
  XOR U16005 ( .A(n10757), .B(n10758), .Z(n10377) );
  AND U16006 ( .A(n10759), .B(n10760), .Z(n10757) );
  AND U16007 ( .A(b[7]), .B(a[92]), .Z(n10756) );
  XOR U16008 ( .A(n10761), .B(n10233), .Z(n10235) );
  IV U16009 ( .A(n10375), .Z(n10233) );
  XOR U16010 ( .A(n10762), .B(n10763), .Z(n10375) );
  AND U16011 ( .A(n10764), .B(n10765), .Z(n10762) );
  AND U16012 ( .A(b[6]), .B(a[93]), .Z(n10761) );
  XOR U16013 ( .A(n10766), .B(n10228), .Z(n10230) );
  IV U16014 ( .A(n10373), .Z(n10228) );
  XOR U16015 ( .A(n10767), .B(n10768), .Z(n10373) );
  AND U16016 ( .A(n10769), .B(n10770), .Z(n10767) );
  AND U16017 ( .A(b[5]), .B(a[94]), .Z(n10766) );
  XOR U16018 ( .A(n10772), .B(n10773), .Z(n10238) );
  AND U16019 ( .A(n10774), .B(n10775), .Z(n10772) );
  AND U16020 ( .A(b[4]), .B(a[95]), .Z(n10771) );
  XOR U16021 ( .A(n10776), .B(n10243), .Z(n10245) );
  IV U16022 ( .A(n10370), .Z(n10243) );
  XOR U16023 ( .A(n10777), .B(n10778), .Z(n10370) );
  AND U16024 ( .A(n10779), .B(n10780), .Z(n10777) );
  AND U16025 ( .A(b[3]), .B(a[96]), .Z(n10776) );
  XOR U16026 ( .A(n10781), .B(n10252), .Z(n10254) );
  IV U16027 ( .A(n10368), .Z(n10252) );
  XNOR U16028 ( .A(n10782), .B(n10783), .Z(n10368) );
  NANDN U16029 ( .A(n10784), .B(n10785), .Z(n10783) );
  AND U16030 ( .A(b[2]), .B(a[97]), .Z(n10781) );
  XOR U16031 ( .A(n10246), .B(n10786), .Z(n10249) );
  NAND U16032 ( .A(b[1]), .B(a[98]), .Z(n10786) );
  OR U16033 ( .A(n10259), .B(n10257), .Z(n10246) );
  XOR U16034 ( .A(n10785), .B(n10784), .Z(n10257) );
  XOR U16035 ( .A(n10782), .B(n10779), .Z(n10787) );
  XOR U16036 ( .A(n10774), .B(n10778), .Z(n10788) );
  XOR U16037 ( .A(n10769), .B(n10773), .Z(n10789) );
  XOR U16038 ( .A(n10764), .B(n10768), .Z(n10790) );
  XOR U16039 ( .A(n10759), .B(n10763), .Z(n10791) );
  XOR U16040 ( .A(n10754), .B(n10758), .Z(n10792) );
  XOR U16041 ( .A(n10749), .B(n10753), .Z(n10793) );
  XOR U16042 ( .A(n10744), .B(n10748), .Z(n10794) );
  XOR U16043 ( .A(n10739), .B(n10743), .Z(n10795) );
  XOR U16044 ( .A(n10734), .B(n10738), .Z(n10796) );
  XOR U16045 ( .A(n10729), .B(n10733), .Z(n10797) );
  XOR U16046 ( .A(n10724), .B(n10728), .Z(n10798) );
  XOR U16047 ( .A(n10719), .B(n10723), .Z(n10799) );
  XOR U16048 ( .A(n10714), .B(n10718), .Z(n10800) );
  XOR U16049 ( .A(n10709), .B(n10713), .Z(n10801) );
  XOR U16050 ( .A(n10704), .B(n10708), .Z(n10802) );
  XOR U16051 ( .A(n10699), .B(n10703), .Z(n10803) );
  XOR U16052 ( .A(n10694), .B(n10698), .Z(n10804) );
  XOR U16053 ( .A(n10689), .B(n10693), .Z(n10805) );
  XOR U16054 ( .A(n10684), .B(n10688), .Z(n10806) );
  XOR U16055 ( .A(n10679), .B(n10683), .Z(n10807) );
  XOR U16056 ( .A(n10674), .B(n10678), .Z(n10808) );
  XOR U16057 ( .A(n10669), .B(n10673), .Z(n10809) );
  XOR U16058 ( .A(n10664), .B(n10668), .Z(n10810) );
  XOR U16059 ( .A(n10659), .B(n10663), .Z(n10811) );
  XOR U16060 ( .A(n10654), .B(n10658), .Z(n10812) );
  XOR U16061 ( .A(n10649), .B(n10653), .Z(n10813) );
  XOR U16062 ( .A(n10644), .B(n10648), .Z(n10814) );
  XOR U16063 ( .A(n10639), .B(n10643), .Z(n10815) );
  XOR U16064 ( .A(n10634), .B(n10638), .Z(n10816) );
  XOR U16065 ( .A(n10629), .B(n10633), .Z(n10817) );
  XOR U16066 ( .A(n10624), .B(n10628), .Z(n10818) );
  XOR U16067 ( .A(n10619), .B(n10623), .Z(n10819) );
  XOR U16068 ( .A(n10614), .B(n10618), .Z(n10820) );
  XOR U16069 ( .A(n10609), .B(n10613), .Z(n10821) );
  XOR U16070 ( .A(n10604), .B(n10608), .Z(n10822) );
  XOR U16071 ( .A(n10599), .B(n10603), .Z(n10823) );
  XOR U16072 ( .A(n10594), .B(n10598), .Z(n10824) );
  XOR U16073 ( .A(n10589), .B(n10593), .Z(n10825) );
  XOR U16074 ( .A(n10584), .B(n10588), .Z(n10826) );
  XOR U16075 ( .A(n10579), .B(n10583), .Z(n10827) );
  XOR U16076 ( .A(n10574), .B(n10578), .Z(n10828) );
  XOR U16077 ( .A(n10569), .B(n10573), .Z(n10829) );
  XOR U16078 ( .A(n10564), .B(n10568), .Z(n10830) );
  XOR U16079 ( .A(n10559), .B(n10563), .Z(n10831) );
  XOR U16080 ( .A(n10554), .B(n10558), .Z(n10832) );
  XOR U16081 ( .A(n10549), .B(n10553), .Z(n10833) );
  XOR U16082 ( .A(n10544), .B(n10548), .Z(n10834) );
  XOR U16083 ( .A(n10539), .B(n10543), .Z(n10835) );
  XOR U16084 ( .A(n10534), .B(n10538), .Z(n10836) );
  XOR U16085 ( .A(n10529), .B(n10533), .Z(n10837) );
  XOR U16086 ( .A(n10524), .B(n10528), .Z(n10838) );
  XOR U16087 ( .A(n10519), .B(n10523), .Z(n10839) );
  XOR U16088 ( .A(n10514), .B(n10518), .Z(n10840) );
  XOR U16089 ( .A(n10509), .B(n10513), .Z(n10841) );
  XOR U16090 ( .A(n10504), .B(n10508), .Z(n10842) );
  XOR U16091 ( .A(n10499), .B(n10503), .Z(n10843) );
  XOR U16092 ( .A(n10494), .B(n10498), .Z(n10844) );
  XNOR U16093 ( .A(n10490), .B(n10493), .Z(n10845) );
  XOR U16094 ( .A(n10846), .B(n10847), .Z(n10490) );
  XOR U16095 ( .A(n10848), .B(n10849), .Z(n10847) );
  XNOR U16096 ( .A(n10850), .B(n10851), .Z(n10848) );
  XOR U16097 ( .A(n10852), .B(n10853), .Z(n10851) );
  AND U16098 ( .A(a[36]), .B(b[62]), .Z(n10853) );
  AND U16099 ( .A(a[35]), .B(b[63]), .Z(n10852) );
  XNOR U16100 ( .A(n10854), .B(n10850), .Z(n10846) );
  XNOR U16101 ( .A(n10855), .B(n10856), .Z(n10850) );
  ANDN U16102 ( .B(n10857), .A(n10858), .Z(n10855) );
  AND U16103 ( .A(a[37]), .B(b[61]), .Z(n10854) );
  XOR U16104 ( .A(n10859), .B(n10488), .Z(n10489) );
  IV U16105 ( .A(n10849), .Z(n10488) );
  XOR U16106 ( .A(n10860), .B(n10861), .Z(n10849) );
  AND U16107 ( .A(n10862), .B(n10863), .Z(n10860) );
  AND U16108 ( .A(a[38]), .B(b[60]), .Z(n10859) );
  XOR U16109 ( .A(n10865), .B(n10866), .Z(n10493) );
  AND U16110 ( .A(n10867), .B(n10868), .Z(n10865) );
  AND U16111 ( .A(a[39]), .B(b[59]), .Z(n10864) );
  XOR U16112 ( .A(n10870), .B(n10871), .Z(n10498) );
  AND U16113 ( .A(n10872), .B(n10873), .Z(n10870) );
  AND U16114 ( .A(a[40]), .B(b[58]), .Z(n10869) );
  XOR U16115 ( .A(n10875), .B(n10876), .Z(n10503) );
  AND U16116 ( .A(n10877), .B(n10878), .Z(n10875) );
  AND U16117 ( .A(a[41]), .B(b[57]), .Z(n10874) );
  XOR U16118 ( .A(n10880), .B(n10881), .Z(n10508) );
  AND U16119 ( .A(n10882), .B(n10883), .Z(n10880) );
  AND U16120 ( .A(a[42]), .B(b[56]), .Z(n10879) );
  XOR U16121 ( .A(n10885), .B(n10886), .Z(n10513) );
  AND U16122 ( .A(n10887), .B(n10888), .Z(n10885) );
  AND U16123 ( .A(a[43]), .B(b[55]), .Z(n10884) );
  XOR U16124 ( .A(n10890), .B(n10891), .Z(n10518) );
  AND U16125 ( .A(n10892), .B(n10893), .Z(n10890) );
  AND U16126 ( .A(a[44]), .B(b[54]), .Z(n10889) );
  XOR U16127 ( .A(n10895), .B(n10896), .Z(n10523) );
  AND U16128 ( .A(n10897), .B(n10898), .Z(n10895) );
  AND U16129 ( .A(a[45]), .B(b[53]), .Z(n10894) );
  XOR U16130 ( .A(n10900), .B(n10901), .Z(n10528) );
  AND U16131 ( .A(n10902), .B(n10903), .Z(n10900) );
  AND U16132 ( .A(a[46]), .B(b[52]), .Z(n10899) );
  XOR U16133 ( .A(n10905), .B(n10906), .Z(n10533) );
  AND U16134 ( .A(n10907), .B(n10908), .Z(n10905) );
  AND U16135 ( .A(a[47]), .B(b[51]), .Z(n10904) );
  XOR U16136 ( .A(n10910), .B(n10911), .Z(n10538) );
  AND U16137 ( .A(n10912), .B(n10913), .Z(n10910) );
  AND U16138 ( .A(a[48]), .B(b[50]), .Z(n10909) );
  XOR U16139 ( .A(n10915), .B(n10916), .Z(n10543) );
  AND U16140 ( .A(n10917), .B(n10918), .Z(n10915) );
  AND U16141 ( .A(a[49]), .B(b[49]), .Z(n10914) );
  XOR U16142 ( .A(n10920), .B(n10921), .Z(n10548) );
  AND U16143 ( .A(n10922), .B(n10923), .Z(n10920) );
  AND U16144 ( .A(b[48]), .B(a[50]), .Z(n10919) );
  XOR U16145 ( .A(n10925), .B(n10926), .Z(n10553) );
  AND U16146 ( .A(n10927), .B(n10928), .Z(n10925) );
  AND U16147 ( .A(b[47]), .B(a[51]), .Z(n10924) );
  XOR U16148 ( .A(n10930), .B(n10931), .Z(n10558) );
  AND U16149 ( .A(n10932), .B(n10933), .Z(n10930) );
  AND U16150 ( .A(b[46]), .B(a[52]), .Z(n10929) );
  XOR U16151 ( .A(n10935), .B(n10936), .Z(n10563) );
  AND U16152 ( .A(n10937), .B(n10938), .Z(n10935) );
  AND U16153 ( .A(b[45]), .B(a[53]), .Z(n10934) );
  XOR U16154 ( .A(n10940), .B(n10941), .Z(n10568) );
  AND U16155 ( .A(n10942), .B(n10943), .Z(n10940) );
  AND U16156 ( .A(b[44]), .B(a[54]), .Z(n10939) );
  XOR U16157 ( .A(n10945), .B(n10946), .Z(n10573) );
  AND U16158 ( .A(n10947), .B(n10948), .Z(n10945) );
  AND U16159 ( .A(b[43]), .B(a[55]), .Z(n10944) );
  XOR U16160 ( .A(n10950), .B(n10951), .Z(n10578) );
  AND U16161 ( .A(n10952), .B(n10953), .Z(n10950) );
  AND U16162 ( .A(b[42]), .B(a[56]), .Z(n10949) );
  XOR U16163 ( .A(n10955), .B(n10956), .Z(n10583) );
  AND U16164 ( .A(n10957), .B(n10958), .Z(n10955) );
  AND U16165 ( .A(b[41]), .B(a[57]), .Z(n10954) );
  XOR U16166 ( .A(n10960), .B(n10961), .Z(n10588) );
  AND U16167 ( .A(n10962), .B(n10963), .Z(n10960) );
  AND U16168 ( .A(b[40]), .B(a[58]), .Z(n10959) );
  XOR U16169 ( .A(n10965), .B(n10966), .Z(n10593) );
  AND U16170 ( .A(n10967), .B(n10968), .Z(n10965) );
  AND U16171 ( .A(b[39]), .B(a[59]), .Z(n10964) );
  XOR U16172 ( .A(n10970), .B(n10971), .Z(n10598) );
  AND U16173 ( .A(n10972), .B(n10973), .Z(n10970) );
  AND U16174 ( .A(b[38]), .B(a[60]), .Z(n10969) );
  XOR U16175 ( .A(n10975), .B(n10976), .Z(n10603) );
  AND U16176 ( .A(n10977), .B(n10978), .Z(n10975) );
  AND U16177 ( .A(b[37]), .B(a[61]), .Z(n10974) );
  XOR U16178 ( .A(n10980), .B(n10981), .Z(n10608) );
  AND U16179 ( .A(n10982), .B(n10983), .Z(n10980) );
  AND U16180 ( .A(b[36]), .B(a[62]), .Z(n10979) );
  XOR U16181 ( .A(n10985), .B(n10986), .Z(n10613) );
  AND U16182 ( .A(n10987), .B(n10988), .Z(n10985) );
  AND U16183 ( .A(b[35]), .B(a[63]), .Z(n10984) );
  XOR U16184 ( .A(n10990), .B(n10991), .Z(n10618) );
  AND U16185 ( .A(n10992), .B(n10993), .Z(n10990) );
  AND U16186 ( .A(b[34]), .B(a[64]), .Z(n10989) );
  XOR U16187 ( .A(n10995), .B(n10996), .Z(n10623) );
  AND U16188 ( .A(n10997), .B(n10998), .Z(n10995) );
  AND U16189 ( .A(b[33]), .B(a[65]), .Z(n10994) );
  XOR U16190 ( .A(n11000), .B(n11001), .Z(n10628) );
  AND U16191 ( .A(n11002), .B(n11003), .Z(n11000) );
  AND U16192 ( .A(b[32]), .B(a[66]), .Z(n10999) );
  XOR U16193 ( .A(n11005), .B(n11006), .Z(n10633) );
  AND U16194 ( .A(n11007), .B(n11008), .Z(n11005) );
  AND U16195 ( .A(b[31]), .B(a[67]), .Z(n11004) );
  XOR U16196 ( .A(n11010), .B(n11011), .Z(n10638) );
  AND U16197 ( .A(n11012), .B(n11013), .Z(n11010) );
  AND U16198 ( .A(b[30]), .B(a[68]), .Z(n11009) );
  XOR U16199 ( .A(n11015), .B(n11016), .Z(n10643) );
  AND U16200 ( .A(n11017), .B(n11018), .Z(n11015) );
  AND U16201 ( .A(b[29]), .B(a[69]), .Z(n11014) );
  XOR U16202 ( .A(n11020), .B(n11021), .Z(n10648) );
  AND U16203 ( .A(n11022), .B(n11023), .Z(n11020) );
  AND U16204 ( .A(b[28]), .B(a[70]), .Z(n11019) );
  XOR U16205 ( .A(n11025), .B(n11026), .Z(n10653) );
  AND U16206 ( .A(n11027), .B(n11028), .Z(n11025) );
  AND U16207 ( .A(b[27]), .B(a[71]), .Z(n11024) );
  XOR U16208 ( .A(n11030), .B(n11031), .Z(n10658) );
  AND U16209 ( .A(n11032), .B(n11033), .Z(n11030) );
  AND U16210 ( .A(b[26]), .B(a[72]), .Z(n11029) );
  XOR U16211 ( .A(n11035), .B(n11036), .Z(n10663) );
  AND U16212 ( .A(n11037), .B(n11038), .Z(n11035) );
  AND U16213 ( .A(b[25]), .B(a[73]), .Z(n11034) );
  XOR U16214 ( .A(n11040), .B(n11041), .Z(n10668) );
  AND U16215 ( .A(n11042), .B(n11043), .Z(n11040) );
  AND U16216 ( .A(b[24]), .B(a[74]), .Z(n11039) );
  XOR U16217 ( .A(n11045), .B(n11046), .Z(n10673) );
  AND U16218 ( .A(n11047), .B(n11048), .Z(n11045) );
  AND U16219 ( .A(b[23]), .B(a[75]), .Z(n11044) );
  XOR U16220 ( .A(n11050), .B(n11051), .Z(n10678) );
  AND U16221 ( .A(n11052), .B(n11053), .Z(n11050) );
  AND U16222 ( .A(b[22]), .B(a[76]), .Z(n11049) );
  XOR U16223 ( .A(n11055), .B(n11056), .Z(n10683) );
  AND U16224 ( .A(n11057), .B(n11058), .Z(n11055) );
  AND U16225 ( .A(b[21]), .B(a[77]), .Z(n11054) );
  XOR U16226 ( .A(n11060), .B(n11061), .Z(n10688) );
  AND U16227 ( .A(n11062), .B(n11063), .Z(n11060) );
  AND U16228 ( .A(b[20]), .B(a[78]), .Z(n11059) );
  XOR U16229 ( .A(n11065), .B(n11066), .Z(n10693) );
  AND U16230 ( .A(n11067), .B(n11068), .Z(n11065) );
  AND U16231 ( .A(b[19]), .B(a[79]), .Z(n11064) );
  XOR U16232 ( .A(n11070), .B(n11071), .Z(n10698) );
  AND U16233 ( .A(n11072), .B(n11073), .Z(n11070) );
  AND U16234 ( .A(b[18]), .B(a[80]), .Z(n11069) );
  XOR U16235 ( .A(n11075), .B(n11076), .Z(n10703) );
  AND U16236 ( .A(n11077), .B(n11078), .Z(n11075) );
  AND U16237 ( .A(b[17]), .B(a[81]), .Z(n11074) );
  XOR U16238 ( .A(n11080), .B(n11081), .Z(n10708) );
  AND U16239 ( .A(n11082), .B(n11083), .Z(n11080) );
  AND U16240 ( .A(b[16]), .B(a[82]), .Z(n11079) );
  XOR U16241 ( .A(n11085), .B(n11086), .Z(n10713) );
  AND U16242 ( .A(n11087), .B(n11088), .Z(n11085) );
  AND U16243 ( .A(b[15]), .B(a[83]), .Z(n11084) );
  XOR U16244 ( .A(n11090), .B(n11091), .Z(n10718) );
  AND U16245 ( .A(n11092), .B(n11093), .Z(n11090) );
  AND U16246 ( .A(b[14]), .B(a[84]), .Z(n11089) );
  XOR U16247 ( .A(n11095), .B(n11096), .Z(n10723) );
  AND U16248 ( .A(n11097), .B(n11098), .Z(n11095) );
  AND U16249 ( .A(b[13]), .B(a[85]), .Z(n11094) );
  XOR U16250 ( .A(n11100), .B(n11101), .Z(n10728) );
  AND U16251 ( .A(n11102), .B(n11103), .Z(n11100) );
  AND U16252 ( .A(b[12]), .B(a[86]), .Z(n11099) );
  XOR U16253 ( .A(n11105), .B(n11106), .Z(n10733) );
  AND U16254 ( .A(n11107), .B(n11108), .Z(n11105) );
  AND U16255 ( .A(b[11]), .B(a[87]), .Z(n11104) );
  XOR U16256 ( .A(n11110), .B(n11111), .Z(n10738) );
  AND U16257 ( .A(n11112), .B(n11113), .Z(n11110) );
  AND U16258 ( .A(b[10]), .B(a[88]), .Z(n11109) );
  XOR U16259 ( .A(n11115), .B(n11116), .Z(n10743) );
  AND U16260 ( .A(n11117), .B(n11118), .Z(n11115) );
  AND U16261 ( .A(b[9]), .B(a[89]), .Z(n11114) );
  XOR U16262 ( .A(n11120), .B(n11121), .Z(n10748) );
  AND U16263 ( .A(n11122), .B(n11123), .Z(n11120) );
  AND U16264 ( .A(b[8]), .B(a[90]), .Z(n11119) );
  XOR U16265 ( .A(n11125), .B(n11126), .Z(n10753) );
  AND U16266 ( .A(n11127), .B(n11128), .Z(n11125) );
  AND U16267 ( .A(b[7]), .B(a[91]), .Z(n11124) );
  XOR U16268 ( .A(n11130), .B(n11131), .Z(n10758) );
  AND U16269 ( .A(n11132), .B(n11133), .Z(n11130) );
  AND U16270 ( .A(b[6]), .B(a[92]), .Z(n11129) );
  XOR U16271 ( .A(n11135), .B(n11136), .Z(n10763) );
  AND U16272 ( .A(n11137), .B(n11138), .Z(n11135) );
  AND U16273 ( .A(b[5]), .B(a[93]), .Z(n11134) );
  XOR U16274 ( .A(n11140), .B(n11141), .Z(n10768) );
  AND U16275 ( .A(n11142), .B(n11143), .Z(n11140) );
  AND U16276 ( .A(b[4]), .B(a[94]), .Z(n11139) );
  XOR U16277 ( .A(n11145), .B(n11146), .Z(n10773) );
  AND U16278 ( .A(n11147), .B(n11148), .Z(n11145) );
  AND U16279 ( .A(b[3]), .B(a[95]), .Z(n11144) );
  XOR U16280 ( .A(n11150), .B(n11151), .Z(n10778) );
  NANDN U16281 ( .A(n11152), .B(n11153), .Z(n11151) );
  AND U16282 ( .A(b[2]), .B(a[96]), .Z(n11149) );
  XOR U16283 ( .A(n10782), .B(n11154), .Z(n10785) );
  NAND U16284 ( .A(b[1]), .B(a[97]), .Z(n11154) );
  OR U16285 ( .A(n10262), .B(n10260), .Z(n10782) );
  XOR U16286 ( .A(n11153), .B(n11152), .Z(n10260) );
  XOR U16287 ( .A(n11156), .B(n11147), .Z(n11155) );
  XOR U16288 ( .A(n11142), .B(n11146), .Z(n11157) );
  XOR U16289 ( .A(n11137), .B(n11141), .Z(n11158) );
  XOR U16290 ( .A(n11132), .B(n11136), .Z(n11159) );
  XOR U16291 ( .A(n11127), .B(n11131), .Z(n11160) );
  XOR U16292 ( .A(n11122), .B(n11126), .Z(n11161) );
  XOR U16293 ( .A(n11117), .B(n11121), .Z(n11162) );
  XOR U16294 ( .A(n11112), .B(n11116), .Z(n11163) );
  XOR U16295 ( .A(n11107), .B(n11111), .Z(n11164) );
  XOR U16296 ( .A(n11102), .B(n11106), .Z(n11165) );
  XOR U16297 ( .A(n11097), .B(n11101), .Z(n11166) );
  XOR U16298 ( .A(n11092), .B(n11096), .Z(n11167) );
  XOR U16299 ( .A(n11087), .B(n11091), .Z(n11168) );
  XOR U16300 ( .A(n11082), .B(n11086), .Z(n11169) );
  XOR U16301 ( .A(n11077), .B(n11081), .Z(n11170) );
  XOR U16302 ( .A(n11072), .B(n11076), .Z(n11171) );
  XOR U16303 ( .A(n11067), .B(n11071), .Z(n11172) );
  XOR U16304 ( .A(n11062), .B(n11066), .Z(n11173) );
  XOR U16305 ( .A(n11057), .B(n11061), .Z(n11174) );
  XOR U16306 ( .A(n11052), .B(n11056), .Z(n11175) );
  XOR U16307 ( .A(n11047), .B(n11051), .Z(n11176) );
  XOR U16308 ( .A(n11042), .B(n11046), .Z(n11177) );
  XOR U16309 ( .A(n11037), .B(n11041), .Z(n11178) );
  XOR U16310 ( .A(n11032), .B(n11036), .Z(n11179) );
  XOR U16311 ( .A(n11027), .B(n11031), .Z(n11180) );
  XOR U16312 ( .A(n11022), .B(n11026), .Z(n11181) );
  XOR U16313 ( .A(n11017), .B(n11021), .Z(n11182) );
  XOR U16314 ( .A(n11012), .B(n11016), .Z(n11183) );
  XOR U16315 ( .A(n11007), .B(n11011), .Z(n11184) );
  XOR U16316 ( .A(n11002), .B(n11006), .Z(n11185) );
  XOR U16317 ( .A(n10997), .B(n11001), .Z(n11186) );
  XOR U16318 ( .A(n10992), .B(n10996), .Z(n11187) );
  XOR U16319 ( .A(n10987), .B(n10991), .Z(n11188) );
  XOR U16320 ( .A(n10982), .B(n10986), .Z(n11189) );
  XOR U16321 ( .A(n10977), .B(n10981), .Z(n11190) );
  XOR U16322 ( .A(n10972), .B(n10976), .Z(n11191) );
  XOR U16323 ( .A(n10967), .B(n10971), .Z(n11192) );
  XOR U16324 ( .A(n10962), .B(n10966), .Z(n11193) );
  XOR U16325 ( .A(n10957), .B(n10961), .Z(n11194) );
  XOR U16326 ( .A(n10952), .B(n10956), .Z(n11195) );
  XOR U16327 ( .A(n10947), .B(n10951), .Z(n11196) );
  XOR U16328 ( .A(n10942), .B(n10946), .Z(n11197) );
  XOR U16329 ( .A(n10937), .B(n10941), .Z(n11198) );
  XOR U16330 ( .A(n10932), .B(n10936), .Z(n11199) );
  XOR U16331 ( .A(n10927), .B(n10931), .Z(n11200) );
  XOR U16332 ( .A(n10922), .B(n10926), .Z(n11201) );
  XOR U16333 ( .A(n10917), .B(n10921), .Z(n11202) );
  XOR U16334 ( .A(n10912), .B(n10916), .Z(n11203) );
  XOR U16335 ( .A(n10907), .B(n10911), .Z(n11204) );
  XOR U16336 ( .A(n10902), .B(n10906), .Z(n11205) );
  XOR U16337 ( .A(n10897), .B(n10901), .Z(n11206) );
  XOR U16338 ( .A(n10892), .B(n10896), .Z(n11207) );
  XOR U16339 ( .A(n10887), .B(n10891), .Z(n11208) );
  XOR U16340 ( .A(n10882), .B(n10886), .Z(n11209) );
  XOR U16341 ( .A(n10877), .B(n10881), .Z(n11210) );
  XOR U16342 ( .A(n10872), .B(n10876), .Z(n11211) );
  XOR U16343 ( .A(n10867), .B(n10871), .Z(n11212) );
  XOR U16344 ( .A(n10862), .B(n10866), .Z(n11213) );
  XNOR U16345 ( .A(n10858), .B(n10861), .Z(n11214) );
  XOR U16346 ( .A(n11215), .B(n11216), .Z(n10858) );
  XOR U16347 ( .A(n11217), .B(n11218), .Z(n11216) );
  XOR U16348 ( .A(n11219), .B(n11220), .Z(n11217) );
  AND U16349 ( .A(a[36]), .B(b[61]), .Z(n11219) );
  XOR U16350 ( .A(n11220), .B(n11221), .Z(n11215) );
  XOR U16351 ( .A(n11222), .B(n11223), .Z(n11221) );
  AND U16352 ( .A(a[35]), .B(b[62]), .Z(n11223) );
  AND U16353 ( .A(a[34]), .B(b[63]), .Z(n11222) );
  XOR U16354 ( .A(n11224), .B(n11225), .Z(n11220) );
  ANDN U16355 ( .B(n11226), .A(n11227), .Z(n11224) );
  XOR U16356 ( .A(n11228), .B(n10856), .Z(n10857) );
  IV U16357 ( .A(n11218), .Z(n10856) );
  XOR U16358 ( .A(n11229), .B(n11230), .Z(n11218) );
  ANDN U16359 ( .B(n11231), .A(n11232), .Z(n11229) );
  AND U16360 ( .A(a[37]), .B(b[60]), .Z(n11228) );
  XOR U16361 ( .A(n11234), .B(n11235), .Z(n10861) );
  AND U16362 ( .A(n11236), .B(n11237), .Z(n11234) );
  AND U16363 ( .A(a[38]), .B(b[59]), .Z(n11233) );
  XOR U16364 ( .A(n11239), .B(n11240), .Z(n10866) );
  AND U16365 ( .A(n11241), .B(n11242), .Z(n11239) );
  AND U16366 ( .A(a[39]), .B(b[58]), .Z(n11238) );
  XOR U16367 ( .A(n11244), .B(n11245), .Z(n10871) );
  AND U16368 ( .A(n11246), .B(n11247), .Z(n11244) );
  AND U16369 ( .A(a[40]), .B(b[57]), .Z(n11243) );
  XOR U16370 ( .A(n11249), .B(n11250), .Z(n10876) );
  AND U16371 ( .A(n11251), .B(n11252), .Z(n11249) );
  AND U16372 ( .A(a[41]), .B(b[56]), .Z(n11248) );
  XOR U16373 ( .A(n11254), .B(n11255), .Z(n10881) );
  AND U16374 ( .A(n11256), .B(n11257), .Z(n11254) );
  AND U16375 ( .A(a[42]), .B(b[55]), .Z(n11253) );
  XOR U16376 ( .A(n11259), .B(n11260), .Z(n10886) );
  AND U16377 ( .A(n11261), .B(n11262), .Z(n11259) );
  AND U16378 ( .A(a[43]), .B(b[54]), .Z(n11258) );
  XOR U16379 ( .A(n11264), .B(n11265), .Z(n10891) );
  AND U16380 ( .A(n11266), .B(n11267), .Z(n11264) );
  AND U16381 ( .A(a[44]), .B(b[53]), .Z(n11263) );
  XOR U16382 ( .A(n11269), .B(n11270), .Z(n10896) );
  AND U16383 ( .A(n11271), .B(n11272), .Z(n11269) );
  AND U16384 ( .A(a[45]), .B(b[52]), .Z(n11268) );
  XOR U16385 ( .A(n11274), .B(n11275), .Z(n10901) );
  AND U16386 ( .A(n11276), .B(n11277), .Z(n11274) );
  AND U16387 ( .A(a[46]), .B(b[51]), .Z(n11273) );
  XOR U16388 ( .A(n11279), .B(n11280), .Z(n10906) );
  AND U16389 ( .A(n11281), .B(n11282), .Z(n11279) );
  AND U16390 ( .A(a[47]), .B(b[50]), .Z(n11278) );
  XOR U16391 ( .A(n11284), .B(n11285), .Z(n10911) );
  AND U16392 ( .A(n11286), .B(n11287), .Z(n11284) );
  AND U16393 ( .A(a[48]), .B(b[49]), .Z(n11283) );
  XOR U16394 ( .A(n11289), .B(n11290), .Z(n10916) );
  AND U16395 ( .A(n11291), .B(n11292), .Z(n11289) );
  AND U16396 ( .A(b[48]), .B(a[49]), .Z(n11288) );
  XOR U16397 ( .A(n11294), .B(n11295), .Z(n10921) );
  AND U16398 ( .A(n11296), .B(n11297), .Z(n11294) );
  AND U16399 ( .A(b[47]), .B(a[50]), .Z(n11293) );
  XOR U16400 ( .A(n11299), .B(n11300), .Z(n10926) );
  AND U16401 ( .A(n11301), .B(n11302), .Z(n11299) );
  AND U16402 ( .A(b[46]), .B(a[51]), .Z(n11298) );
  XOR U16403 ( .A(n11304), .B(n11305), .Z(n10931) );
  AND U16404 ( .A(n11306), .B(n11307), .Z(n11304) );
  AND U16405 ( .A(b[45]), .B(a[52]), .Z(n11303) );
  XOR U16406 ( .A(n11309), .B(n11310), .Z(n10936) );
  AND U16407 ( .A(n11311), .B(n11312), .Z(n11309) );
  AND U16408 ( .A(b[44]), .B(a[53]), .Z(n11308) );
  XOR U16409 ( .A(n11314), .B(n11315), .Z(n10941) );
  AND U16410 ( .A(n11316), .B(n11317), .Z(n11314) );
  AND U16411 ( .A(b[43]), .B(a[54]), .Z(n11313) );
  XOR U16412 ( .A(n11319), .B(n11320), .Z(n10946) );
  AND U16413 ( .A(n11321), .B(n11322), .Z(n11319) );
  AND U16414 ( .A(b[42]), .B(a[55]), .Z(n11318) );
  XOR U16415 ( .A(n11324), .B(n11325), .Z(n10951) );
  AND U16416 ( .A(n11326), .B(n11327), .Z(n11324) );
  AND U16417 ( .A(b[41]), .B(a[56]), .Z(n11323) );
  XOR U16418 ( .A(n11329), .B(n11330), .Z(n10956) );
  AND U16419 ( .A(n11331), .B(n11332), .Z(n11329) );
  AND U16420 ( .A(b[40]), .B(a[57]), .Z(n11328) );
  XOR U16421 ( .A(n11334), .B(n11335), .Z(n10961) );
  AND U16422 ( .A(n11336), .B(n11337), .Z(n11334) );
  AND U16423 ( .A(b[39]), .B(a[58]), .Z(n11333) );
  XOR U16424 ( .A(n11339), .B(n11340), .Z(n10966) );
  AND U16425 ( .A(n11341), .B(n11342), .Z(n11339) );
  AND U16426 ( .A(b[38]), .B(a[59]), .Z(n11338) );
  XOR U16427 ( .A(n11344), .B(n11345), .Z(n10971) );
  AND U16428 ( .A(n11346), .B(n11347), .Z(n11344) );
  AND U16429 ( .A(b[37]), .B(a[60]), .Z(n11343) );
  XOR U16430 ( .A(n11349), .B(n11350), .Z(n10976) );
  AND U16431 ( .A(n11351), .B(n11352), .Z(n11349) );
  AND U16432 ( .A(b[36]), .B(a[61]), .Z(n11348) );
  XOR U16433 ( .A(n11354), .B(n11355), .Z(n10981) );
  AND U16434 ( .A(n11356), .B(n11357), .Z(n11354) );
  AND U16435 ( .A(b[35]), .B(a[62]), .Z(n11353) );
  XOR U16436 ( .A(n11359), .B(n11360), .Z(n10986) );
  AND U16437 ( .A(n11361), .B(n11362), .Z(n11359) );
  AND U16438 ( .A(b[34]), .B(a[63]), .Z(n11358) );
  XOR U16439 ( .A(n11364), .B(n11365), .Z(n10991) );
  AND U16440 ( .A(n11366), .B(n11367), .Z(n11364) );
  AND U16441 ( .A(b[33]), .B(a[64]), .Z(n11363) );
  XOR U16442 ( .A(n11369), .B(n11370), .Z(n10996) );
  AND U16443 ( .A(n11371), .B(n11372), .Z(n11369) );
  AND U16444 ( .A(b[32]), .B(a[65]), .Z(n11368) );
  XOR U16445 ( .A(n11374), .B(n11375), .Z(n11001) );
  AND U16446 ( .A(n11376), .B(n11377), .Z(n11374) );
  AND U16447 ( .A(b[31]), .B(a[66]), .Z(n11373) );
  XOR U16448 ( .A(n11379), .B(n11380), .Z(n11006) );
  AND U16449 ( .A(n11381), .B(n11382), .Z(n11379) );
  AND U16450 ( .A(b[30]), .B(a[67]), .Z(n11378) );
  XOR U16451 ( .A(n11384), .B(n11385), .Z(n11011) );
  AND U16452 ( .A(n11386), .B(n11387), .Z(n11384) );
  AND U16453 ( .A(b[29]), .B(a[68]), .Z(n11383) );
  XOR U16454 ( .A(n11389), .B(n11390), .Z(n11016) );
  AND U16455 ( .A(n11391), .B(n11392), .Z(n11389) );
  AND U16456 ( .A(b[28]), .B(a[69]), .Z(n11388) );
  XOR U16457 ( .A(n11394), .B(n11395), .Z(n11021) );
  AND U16458 ( .A(n11396), .B(n11397), .Z(n11394) );
  AND U16459 ( .A(b[27]), .B(a[70]), .Z(n11393) );
  XOR U16460 ( .A(n11399), .B(n11400), .Z(n11026) );
  AND U16461 ( .A(n11401), .B(n11402), .Z(n11399) );
  AND U16462 ( .A(b[26]), .B(a[71]), .Z(n11398) );
  XOR U16463 ( .A(n11404), .B(n11405), .Z(n11031) );
  AND U16464 ( .A(n11406), .B(n11407), .Z(n11404) );
  AND U16465 ( .A(b[25]), .B(a[72]), .Z(n11403) );
  XOR U16466 ( .A(n11409), .B(n11410), .Z(n11036) );
  AND U16467 ( .A(n11411), .B(n11412), .Z(n11409) );
  AND U16468 ( .A(b[24]), .B(a[73]), .Z(n11408) );
  XOR U16469 ( .A(n11414), .B(n11415), .Z(n11041) );
  AND U16470 ( .A(n11416), .B(n11417), .Z(n11414) );
  AND U16471 ( .A(b[23]), .B(a[74]), .Z(n11413) );
  XOR U16472 ( .A(n11419), .B(n11420), .Z(n11046) );
  AND U16473 ( .A(n11421), .B(n11422), .Z(n11419) );
  AND U16474 ( .A(b[22]), .B(a[75]), .Z(n11418) );
  XOR U16475 ( .A(n11424), .B(n11425), .Z(n11051) );
  AND U16476 ( .A(n11426), .B(n11427), .Z(n11424) );
  AND U16477 ( .A(b[21]), .B(a[76]), .Z(n11423) );
  XOR U16478 ( .A(n11429), .B(n11430), .Z(n11056) );
  AND U16479 ( .A(n11431), .B(n11432), .Z(n11429) );
  AND U16480 ( .A(b[20]), .B(a[77]), .Z(n11428) );
  XOR U16481 ( .A(n11434), .B(n11435), .Z(n11061) );
  AND U16482 ( .A(n11436), .B(n11437), .Z(n11434) );
  AND U16483 ( .A(b[19]), .B(a[78]), .Z(n11433) );
  XOR U16484 ( .A(n11439), .B(n11440), .Z(n11066) );
  AND U16485 ( .A(n11441), .B(n11442), .Z(n11439) );
  AND U16486 ( .A(b[18]), .B(a[79]), .Z(n11438) );
  XOR U16487 ( .A(n11444), .B(n11445), .Z(n11071) );
  AND U16488 ( .A(n11446), .B(n11447), .Z(n11444) );
  AND U16489 ( .A(b[17]), .B(a[80]), .Z(n11443) );
  XOR U16490 ( .A(n11449), .B(n11450), .Z(n11076) );
  AND U16491 ( .A(n11451), .B(n11452), .Z(n11449) );
  AND U16492 ( .A(b[16]), .B(a[81]), .Z(n11448) );
  XOR U16493 ( .A(n11454), .B(n11455), .Z(n11081) );
  AND U16494 ( .A(n11456), .B(n11457), .Z(n11454) );
  AND U16495 ( .A(b[15]), .B(a[82]), .Z(n11453) );
  XOR U16496 ( .A(n11459), .B(n11460), .Z(n11086) );
  AND U16497 ( .A(n11461), .B(n11462), .Z(n11459) );
  AND U16498 ( .A(b[14]), .B(a[83]), .Z(n11458) );
  XOR U16499 ( .A(n11464), .B(n11465), .Z(n11091) );
  AND U16500 ( .A(n11466), .B(n11467), .Z(n11464) );
  AND U16501 ( .A(b[13]), .B(a[84]), .Z(n11463) );
  XOR U16502 ( .A(n11469), .B(n11470), .Z(n11096) );
  AND U16503 ( .A(n11471), .B(n11472), .Z(n11469) );
  AND U16504 ( .A(b[12]), .B(a[85]), .Z(n11468) );
  XOR U16505 ( .A(n11474), .B(n11475), .Z(n11101) );
  AND U16506 ( .A(n11476), .B(n11477), .Z(n11474) );
  AND U16507 ( .A(b[11]), .B(a[86]), .Z(n11473) );
  XOR U16508 ( .A(n11479), .B(n11480), .Z(n11106) );
  AND U16509 ( .A(n11481), .B(n11482), .Z(n11479) );
  AND U16510 ( .A(b[10]), .B(a[87]), .Z(n11478) );
  XOR U16511 ( .A(n11484), .B(n11485), .Z(n11111) );
  AND U16512 ( .A(n11486), .B(n11487), .Z(n11484) );
  AND U16513 ( .A(b[9]), .B(a[88]), .Z(n11483) );
  XOR U16514 ( .A(n11489), .B(n11490), .Z(n11116) );
  AND U16515 ( .A(n11491), .B(n11492), .Z(n11489) );
  AND U16516 ( .A(b[8]), .B(a[89]), .Z(n11488) );
  XOR U16517 ( .A(n11494), .B(n11495), .Z(n11121) );
  AND U16518 ( .A(n11496), .B(n11497), .Z(n11494) );
  AND U16519 ( .A(b[7]), .B(a[90]), .Z(n11493) );
  XOR U16520 ( .A(n11499), .B(n11500), .Z(n11126) );
  AND U16521 ( .A(n11501), .B(n11502), .Z(n11499) );
  AND U16522 ( .A(b[6]), .B(a[91]), .Z(n11498) );
  XOR U16523 ( .A(n11504), .B(n11505), .Z(n11131) );
  AND U16524 ( .A(n11506), .B(n11507), .Z(n11504) );
  AND U16525 ( .A(b[5]), .B(a[92]), .Z(n11503) );
  XOR U16526 ( .A(n11509), .B(n11510), .Z(n11136) );
  AND U16527 ( .A(n11511), .B(n11512), .Z(n11509) );
  AND U16528 ( .A(b[4]), .B(a[93]), .Z(n11508) );
  XOR U16529 ( .A(n11514), .B(n11515), .Z(n11141) );
  AND U16530 ( .A(n11516), .B(n11517), .Z(n11514) );
  AND U16531 ( .A(b[3]), .B(a[94]), .Z(n11513) );
  IV U16532 ( .A(n11150), .Z(n11156) );
  XOR U16533 ( .A(n11519), .B(n11520), .Z(n11146) );
  OR U16534 ( .A(n11521), .B(n11522), .Z(n11520) );
  AND U16535 ( .A(b[2]), .B(a[95]), .Z(n11518) );
  XNOR U16536 ( .A(n11150), .B(n11523), .Z(n11153) );
  NAND U16537 ( .A(b[1]), .B(a[96]), .Z(n11523) );
  ANDN U16538 ( .B(n10263), .A(n10265), .Z(n11150) );
  NAND U16539 ( .A(a[96]), .B(b[0]), .Z(n10265) );
  XOR U16540 ( .A(n11521), .B(n11522), .Z(n10263) );
  XOR U16541 ( .A(n11525), .B(n11516), .Z(n11524) );
  XOR U16542 ( .A(n11511), .B(n11515), .Z(n11526) );
  XOR U16543 ( .A(n11506), .B(n11510), .Z(n11527) );
  XOR U16544 ( .A(n11501), .B(n11505), .Z(n11528) );
  XOR U16545 ( .A(n11496), .B(n11500), .Z(n11529) );
  XOR U16546 ( .A(n11491), .B(n11495), .Z(n11530) );
  XOR U16547 ( .A(n11486), .B(n11490), .Z(n11531) );
  XOR U16548 ( .A(n11481), .B(n11485), .Z(n11532) );
  XOR U16549 ( .A(n11476), .B(n11480), .Z(n11533) );
  XOR U16550 ( .A(n11471), .B(n11475), .Z(n11534) );
  XOR U16551 ( .A(n11466), .B(n11470), .Z(n11535) );
  XOR U16552 ( .A(n11461), .B(n11465), .Z(n11536) );
  XOR U16553 ( .A(n11456), .B(n11460), .Z(n11537) );
  XOR U16554 ( .A(n11451), .B(n11455), .Z(n11538) );
  XOR U16555 ( .A(n11446), .B(n11450), .Z(n11539) );
  XOR U16556 ( .A(n11441), .B(n11445), .Z(n11540) );
  XOR U16557 ( .A(n11436), .B(n11440), .Z(n11541) );
  XOR U16558 ( .A(n11431), .B(n11435), .Z(n11542) );
  XOR U16559 ( .A(n11426), .B(n11430), .Z(n11543) );
  XOR U16560 ( .A(n11421), .B(n11425), .Z(n11544) );
  XOR U16561 ( .A(n11416), .B(n11420), .Z(n11545) );
  XOR U16562 ( .A(n11411), .B(n11415), .Z(n11546) );
  XOR U16563 ( .A(n11406), .B(n11410), .Z(n11547) );
  XOR U16564 ( .A(n11401), .B(n11405), .Z(n11548) );
  XOR U16565 ( .A(n11396), .B(n11400), .Z(n11549) );
  XOR U16566 ( .A(n11391), .B(n11395), .Z(n11550) );
  XOR U16567 ( .A(n11386), .B(n11390), .Z(n11551) );
  XOR U16568 ( .A(n11381), .B(n11385), .Z(n11552) );
  XOR U16569 ( .A(n11376), .B(n11380), .Z(n11553) );
  XOR U16570 ( .A(n11371), .B(n11375), .Z(n11554) );
  XOR U16571 ( .A(n11366), .B(n11370), .Z(n11555) );
  XOR U16572 ( .A(n11361), .B(n11365), .Z(n11556) );
  XOR U16573 ( .A(n11356), .B(n11360), .Z(n11557) );
  XOR U16574 ( .A(n11351), .B(n11355), .Z(n11558) );
  XOR U16575 ( .A(n11346), .B(n11350), .Z(n11559) );
  XOR U16576 ( .A(n11341), .B(n11345), .Z(n11560) );
  XOR U16577 ( .A(n11336), .B(n11340), .Z(n11561) );
  XOR U16578 ( .A(n11331), .B(n11335), .Z(n11562) );
  XOR U16579 ( .A(n11326), .B(n11330), .Z(n11563) );
  XOR U16580 ( .A(n11321), .B(n11325), .Z(n11564) );
  XOR U16581 ( .A(n11316), .B(n11320), .Z(n11565) );
  XOR U16582 ( .A(n11311), .B(n11315), .Z(n11566) );
  XOR U16583 ( .A(n11306), .B(n11310), .Z(n11567) );
  XOR U16584 ( .A(n11301), .B(n11305), .Z(n11568) );
  XOR U16585 ( .A(n11296), .B(n11300), .Z(n11569) );
  XOR U16586 ( .A(n11291), .B(n11295), .Z(n11570) );
  XOR U16587 ( .A(n11286), .B(n11290), .Z(n11571) );
  XOR U16588 ( .A(n11281), .B(n11285), .Z(n11572) );
  XOR U16589 ( .A(n11276), .B(n11280), .Z(n11573) );
  XOR U16590 ( .A(n11271), .B(n11275), .Z(n11574) );
  XOR U16591 ( .A(n11266), .B(n11270), .Z(n11575) );
  XOR U16592 ( .A(n11261), .B(n11265), .Z(n11576) );
  XOR U16593 ( .A(n11256), .B(n11260), .Z(n11577) );
  XOR U16594 ( .A(n11251), .B(n11255), .Z(n11578) );
  XOR U16595 ( .A(n11246), .B(n11250), .Z(n11579) );
  XOR U16596 ( .A(n11241), .B(n11245), .Z(n11580) );
  XOR U16597 ( .A(n11236), .B(n11240), .Z(n11581) );
  XNOR U16598 ( .A(n11232), .B(n11235), .Z(n11582) );
  XNOR U16599 ( .A(n11227), .B(n11583), .Z(n11232) );
  XOR U16600 ( .A(n11226), .B(n11230), .Z(n11583) );
  XOR U16601 ( .A(n11584), .B(n11225), .Z(n11226) );
  AND U16602 ( .A(a[36]), .B(b[60]), .Z(n11584) );
  XOR U16603 ( .A(n11585), .B(n11586), .Z(n11227) );
  XOR U16604 ( .A(n11225), .B(n11587), .Z(n11586) );
  XOR U16605 ( .A(n11588), .B(n11589), .Z(n11587) );
  XOR U16606 ( .A(n11590), .B(n11591), .Z(n11589) );
  NAND U16607 ( .A(a[34]), .B(b[62]), .Z(n11591) );
  AND U16608 ( .A(a[33]), .B(b[63]), .Z(n11590) );
  XOR U16609 ( .A(n11592), .B(n11593), .Z(n11225) );
  AND U16610 ( .A(n11594), .B(n11595), .Z(n11592) );
  XOR U16611 ( .A(n11596), .B(n11588), .Z(n11585) );
  XOR U16612 ( .A(n11597), .B(n11598), .Z(n11588) );
  ANDN U16613 ( .B(n11599), .A(n11600), .Z(n11597) );
  AND U16614 ( .A(a[35]), .B(b[61]), .Z(n11596) );
  XOR U16615 ( .A(n11602), .B(n11603), .Z(n11230) );
  AND U16616 ( .A(n11604), .B(n11605), .Z(n11602) );
  AND U16617 ( .A(a[37]), .B(b[59]), .Z(n11601) );
  XOR U16618 ( .A(n11607), .B(n11608), .Z(n11235) );
  AND U16619 ( .A(n11609), .B(n11610), .Z(n11607) );
  AND U16620 ( .A(a[38]), .B(b[58]), .Z(n11606) );
  XOR U16621 ( .A(n11612), .B(n11613), .Z(n11240) );
  AND U16622 ( .A(n11614), .B(n11615), .Z(n11612) );
  AND U16623 ( .A(a[39]), .B(b[57]), .Z(n11611) );
  XOR U16624 ( .A(n11617), .B(n11618), .Z(n11245) );
  AND U16625 ( .A(n11619), .B(n11620), .Z(n11617) );
  AND U16626 ( .A(a[40]), .B(b[56]), .Z(n11616) );
  XOR U16627 ( .A(n11622), .B(n11623), .Z(n11250) );
  AND U16628 ( .A(n11624), .B(n11625), .Z(n11622) );
  AND U16629 ( .A(a[41]), .B(b[55]), .Z(n11621) );
  XOR U16630 ( .A(n11627), .B(n11628), .Z(n11255) );
  AND U16631 ( .A(n11629), .B(n11630), .Z(n11627) );
  AND U16632 ( .A(a[42]), .B(b[54]), .Z(n11626) );
  XOR U16633 ( .A(n11632), .B(n11633), .Z(n11260) );
  AND U16634 ( .A(n11634), .B(n11635), .Z(n11632) );
  AND U16635 ( .A(a[43]), .B(b[53]), .Z(n11631) );
  XOR U16636 ( .A(n11637), .B(n11638), .Z(n11265) );
  AND U16637 ( .A(n11639), .B(n11640), .Z(n11637) );
  AND U16638 ( .A(a[44]), .B(b[52]), .Z(n11636) );
  XOR U16639 ( .A(n11642), .B(n11643), .Z(n11270) );
  AND U16640 ( .A(n11644), .B(n11645), .Z(n11642) );
  AND U16641 ( .A(a[45]), .B(b[51]), .Z(n11641) );
  XOR U16642 ( .A(n11647), .B(n11648), .Z(n11275) );
  AND U16643 ( .A(n11649), .B(n11650), .Z(n11647) );
  AND U16644 ( .A(a[46]), .B(b[50]), .Z(n11646) );
  XOR U16645 ( .A(n11652), .B(n11653), .Z(n11280) );
  AND U16646 ( .A(n11654), .B(n11655), .Z(n11652) );
  AND U16647 ( .A(a[47]), .B(b[49]), .Z(n11651) );
  XOR U16648 ( .A(n11657), .B(n11658), .Z(n11285) );
  AND U16649 ( .A(n11659), .B(n11660), .Z(n11657) );
  AND U16650 ( .A(a[48]), .B(b[48]), .Z(n11656) );
  XOR U16651 ( .A(n11662), .B(n11663), .Z(n11290) );
  AND U16652 ( .A(n11664), .B(n11665), .Z(n11662) );
  AND U16653 ( .A(b[47]), .B(a[49]), .Z(n11661) );
  XOR U16654 ( .A(n11667), .B(n11668), .Z(n11295) );
  AND U16655 ( .A(n11669), .B(n11670), .Z(n11667) );
  AND U16656 ( .A(b[46]), .B(a[50]), .Z(n11666) );
  XOR U16657 ( .A(n11672), .B(n11673), .Z(n11300) );
  AND U16658 ( .A(n11674), .B(n11675), .Z(n11672) );
  AND U16659 ( .A(b[45]), .B(a[51]), .Z(n11671) );
  XOR U16660 ( .A(n11677), .B(n11678), .Z(n11305) );
  AND U16661 ( .A(n11679), .B(n11680), .Z(n11677) );
  AND U16662 ( .A(b[44]), .B(a[52]), .Z(n11676) );
  XOR U16663 ( .A(n11682), .B(n11683), .Z(n11310) );
  AND U16664 ( .A(n11684), .B(n11685), .Z(n11682) );
  AND U16665 ( .A(b[43]), .B(a[53]), .Z(n11681) );
  XOR U16666 ( .A(n11687), .B(n11688), .Z(n11315) );
  AND U16667 ( .A(n11689), .B(n11690), .Z(n11687) );
  AND U16668 ( .A(b[42]), .B(a[54]), .Z(n11686) );
  XOR U16669 ( .A(n11692), .B(n11693), .Z(n11320) );
  AND U16670 ( .A(n11694), .B(n11695), .Z(n11692) );
  AND U16671 ( .A(b[41]), .B(a[55]), .Z(n11691) );
  XOR U16672 ( .A(n11697), .B(n11698), .Z(n11325) );
  AND U16673 ( .A(n11699), .B(n11700), .Z(n11697) );
  AND U16674 ( .A(b[40]), .B(a[56]), .Z(n11696) );
  XOR U16675 ( .A(n11702), .B(n11703), .Z(n11330) );
  AND U16676 ( .A(n11704), .B(n11705), .Z(n11702) );
  AND U16677 ( .A(b[39]), .B(a[57]), .Z(n11701) );
  XOR U16678 ( .A(n11707), .B(n11708), .Z(n11335) );
  AND U16679 ( .A(n11709), .B(n11710), .Z(n11707) );
  AND U16680 ( .A(b[38]), .B(a[58]), .Z(n11706) );
  XOR U16681 ( .A(n11712), .B(n11713), .Z(n11340) );
  AND U16682 ( .A(n11714), .B(n11715), .Z(n11712) );
  AND U16683 ( .A(b[37]), .B(a[59]), .Z(n11711) );
  XOR U16684 ( .A(n11717), .B(n11718), .Z(n11345) );
  AND U16685 ( .A(n11719), .B(n11720), .Z(n11717) );
  AND U16686 ( .A(b[36]), .B(a[60]), .Z(n11716) );
  XOR U16687 ( .A(n11722), .B(n11723), .Z(n11350) );
  AND U16688 ( .A(n11724), .B(n11725), .Z(n11722) );
  AND U16689 ( .A(b[35]), .B(a[61]), .Z(n11721) );
  XOR U16690 ( .A(n11727), .B(n11728), .Z(n11355) );
  AND U16691 ( .A(n11729), .B(n11730), .Z(n11727) );
  AND U16692 ( .A(b[34]), .B(a[62]), .Z(n11726) );
  XOR U16693 ( .A(n11732), .B(n11733), .Z(n11360) );
  AND U16694 ( .A(n11734), .B(n11735), .Z(n11732) );
  AND U16695 ( .A(b[33]), .B(a[63]), .Z(n11731) );
  XOR U16696 ( .A(n11737), .B(n11738), .Z(n11365) );
  AND U16697 ( .A(n11739), .B(n11740), .Z(n11737) );
  AND U16698 ( .A(b[32]), .B(a[64]), .Z(n11736) );
  XOR U16699 ( .A(n11742), .B(n11743), .Z(n11370) );
  AND U16700 ( .A(n11744), .B(n11745), .Z(n11742) );
  AND U16701 ( .A(b[31]), .B(a[65]), .Z(n11741) );
  XOR U16702 ( .A(n11747), .B(n11748), .Z(n11375) );
  AND U16703 ( .A(n11749), .B(n11750), .Z(n11747) );
  AND U16704 ( .A(b[30]), .B(a[66]), .Z(n11746) );
  XOR U16705 ( .A(n11752), .B(n11753), .Z(n11380) );
  AND U16706 ( .A(n11754), .B(n11755), .Z(n11752) );
  AND U16707 ( .A(b[29]), .B(a[67]), .Z(n11751) );
  XOR U16708 ( .A(n11757), .B(n11758), .Z(n11385) );
  AND U16709 ( .A(n11759), .B(n11760), .Z(n11757) );
  AND U16710 ( .A(b[28]), .B(a[68]), .Z(n11756) );
  XOR U16711 ( .A(n11762), .B(n11763), .Z(n11390) );
  AND U16712 ( .A(n11764), .B(n11765), .Z(n11762) );
  AND U16713 ( .A(b[27]), .B(a[69]), .Z(n11761) );
  XOR U16714 ( .A(n11767), .B(n11768), .Z(n11395) );
  AND U16715 ( .A(n11769), .B(n11770), .Z(n11767) );
  AND U16716 ( .A(b[26]), .B(a[70]), .Z(n11766) );
  XOR U16717 ( .A(n11772), .B(n11773), .Z(n11400) );
  AND U16718 ( .A(n11774), .B(n11775), .Z(n11772) );
  AND U16719 ( .A(b[25]), .B(a[71]), .Z(n11771) );
  XOR U16720 ( .A(n11777), .B(n11778), .Z(n11405) );
  AND U16721 ( .A(n11779), .B(n11780), .Z(n11777) );
  AND U16722 ( .A(b[24]), .B(a[72]), .Z(n11776) );
  XOR U16723 ( .A(n11782), .B(n11783), .Z(n11410) );
  AND U16724 ( .A(n11784), .B(n11785), .Z(n11782) );
  AND U16725 ( .A(b[23]), .B(a[73]), .Z(n11781) );
  XOR U16726 ( .A(n11787), .B(n11788), .Z(n11415) );
  AND U16727 ( .A(n11789), .B(n11790), .Z(n11787) );
  AND U16728 ( .A(b[22]), .B(a[74]), .Z(n11786) );
  XOR U16729 ( .A(n11792), .B(n11793), .Z(n11420) );
  AND U16730 ( .A(n11794), .B(n11795), .Z(n11792) );
  AND U16731 ( .A(b[21]), .B(a[75]), .Z(n11791) );
  XOR U16732 ( .A(n11797), .B(n11798), .Z(n11425) );
  AND U16733 ( .A(n11799), .B(n11800), .Z(n11797) );
  AND U16734 ( .A(b[20]), .B(a[76]), .Z(n11796) );
  XOR U16735 ( .A(n11802), .B(n11803), .Z(n11430) );
  AND U16736 ( .A(n11804), .B(n11805), .Z(n11802) );
  AND U16737 ( .A(b[19]), .B(a[77]), .Z(n11801) );
  XOR U16738 ( .A(n11807), .B(n11808), .Z(n11435) );
  AND U16739 ( .A(n11809), .B(n11810), .Z(n11807) );
  AND U16740 ( .A(b[18]), .B(a[78]), .Z(n11806) );
  XOR U16741 ( .A(n11812), .B(n11813), .Z(n11440) );
  AND U16742 ( .A(n11814), .B(n11815), .Z(n11812) );
  AND U16743 ( .A(b[17]), .B(a[79]), .Z(n11811) );
  XOR U16744 ( .A(n11817), .B(n11818), .Z(n11445) );
  AND U16745 ( .A(n11819), .B(n11820), .Z(n11817) );
  AND U16746 ( .A(b[16]), .B(a[80]), .Z(n11816) );
  XOR U16747 ( .A(n11822), .B(n11823), .Z(n11450) );
  AND U16748 ( .A(n11824), .B(n11825), .Z(n11822) );
  AND U16749 ( .A(b[15]), .B(a[81]), .Z(n11821) );
  XOR U16750 ( .A(n11827), .B(n11828), .Z(n11455) );
  AND U16751 ( .A(n11829), .B(n11830), .Z(n11827) );
  AND U16752 ( .A(b[14]), .B(a[82]), .Z(n11826) );
  XOR U16753 ( .A(n11832), .B(n11833), .Z(n11460) );
  AND U16754 ( .A(n11834), .B(n11835), .Z(n11832) );
  AND U16755 ( .A(b[13]), .B(a[83]), .Z(n11831) );
  XOR U16756 ( .A(n11837), .B(n11838), .Z(n11465) );
  AND U16757 ( .A(n11839), .B(n11840), .Z(n11837) );
  AND U16758 ( .A(b[12]), .B(a[84]), .Z(n11836) );
  XOR U16759 ( .A(n11842), .B(n11843), .Z(n11470) );
  AND U16760 ( .A(n11844), .B(n11845), .Z(n11842) );
  AND U16761 ( .A(b[11]), .B(a[85]), .Z(n11841) );
  XOR U16762 ( .A(n11847), .B(n11848), .Z(n11475) );
  AND U16763 ( .A(n11849), .B(n11850), .Z(n11847) );
  AND U16764 ( .A(b[10]), .B(a[86]), .Z(n11846) );
  XOR U16765 ( .A(n11852), .B(n11853), .Z(n11480) );
  AND U16766 ( .A(n11854), .B(n11855), .Z(n11852) );
  AND U16767 ( .A(b[9]), .B(a[87]), .Z(n11851) );
  XOR U16768 ( .A(n11857), .B(n11858), .Z(n11485) );
  AND U16769 ( .A(n11859), .B(n11860), .Z(n11857) );
  AND U16770 ( .A(b[8]), .B(a[88]), .Z(n11856) );
  XOR U16771 ( .A(n11862), .B(n11863), .Z(n11490) );
  AND U16772 ( .A(n11864), .B(n11865), .Z(n11862) );
  AND U16773 ( .A(b[7]), .B(a[89]), .Z(n11861) );
  XOR U16774 ( .A(n11867), .B(n11868), .Z(n11495) );
  AND U16775 ( .A(n11869), .B(n11870), .Z(n11867) );
  AND U16776 ( .A(b[6]), .B(a[90]), .Z(n11866) );
  XOR U16777 ( .A(n11872), .B(n11873), .Z(n11500) );
  AND U16778 ( .A(n11874), .B(n11875), .Z(n11872) );
  AND U16779 ( .A(b[5]), .B(a[91]), .Z(n11871) );
  XOR U16780 ( .A(n11877), .B(n11878), .Z(n11505) );
  AND U16781 ( .A(n11879), .B(n11880), .Z(n11877) );
  AND U16782 ( .A(b[4]), .B(a[92]), .Z(n11876) );
  XOR U16783 ( .A(n11882), .B(n11883), .Z(n11510) );
  AND U16784 ( .A(n11884), .B(n11885), .Z(n11882) );
  AND U16785 ( .A(b[3]), .B(a[93]), .Z(n11881) );
  XOR U16786 ( .A(n11887), .B(n11888), .Z(n11515) );
  OR U16787 ( .A(n11889), .B(n11890), .Z(n11888) );
  AND U16788 ( .A(b[2]), .B(a[94]), .Z(n11886) );
  XNOR U16789 ( .A(n11525), .B(n11891), .Z(n11521) );
  NAND U16790 ( .A(b[1]), .B(a[95]), .Z(n11891) );
  IV U16791 ( .A(n11519), .Z(n11525) );
  ANDN U16792 ( .B(n10266), .A(n10268), .Z(n11519) );
  NAND U16793 ( .A(a[95]), .B(b[0]), .Z(n10268) );
  XOR U16794 ( .A(n11889), .B(n11890), .Z(n10266) );
  XOR U16795 ( .A(n11893), .B(n11884), .Z(n11892) );
  XOR U16796 ( .A(n11879), .B(n11883), .Z(n11894) );
  XOR U16797 ( .A(n11874), .B(n11878), .Z(n11895) );
  XOR U16798 ( .A(n11869), .B(n11873), .Z(n11896) );
  XOR U16799 ( .A(n11864), .B(n11868), .Z(n11897) );
  XOR U16800 ( .A(n11859), .B(n11863), .Z(n11898) );
  XOR U16801 ( .A(n11854), .B(n11858), .Z(n11899) );
  XOR U16802 ( .A(n11849), .B(n11853), .Z(n11900) );
  XOR U16803 ( .A(n11844), .B(n11848), .Z(n11901) );
  XOR U16804 ( .A(n11839), .B(n11843), .Z(n11902) );
  XOR U16805 ( .A(n11834), .B(n11838), .Z(n11903) );
  XOR U16806 ( .A(n11829), .B(n11833), .Z(n11904) );
  XOR U16807 ( .A(n11824), .B(n11828), .Z(n11905) );
  XOR U16808 ( .A(n11819), .B(n11823), .Z(n11906) );
  XOR U16809 ( .A(n11814), .B(n11818), .Z(n11907) );
  XOR U16810 ( .A(n11809), .B(n11813), .Z(n11908) );
  XOR U16811 ( .A(n11804), .B(n11808), .Z(n11909) );
  XOR U16812 ( .A(n11799), .B(n11803), .Z(n11910) );
  XOR U16813 ( .A(n11794), .B(n11798), .Z(n11911) );
  XOR U16814 ( .A(n11789), .B(n11793), .Z(n11912) );
  XOR U16815 ( .A(n11784), .B(n11788), .Z(n11913) );
  XOR U16816 ( .A(n11779), .B(n11783), .Z(n11914) );
  XOR U16817 ( .A(n11774), .B(n11778), .Z(n11915) );
  XOR U16818 ( .A(n11769), .B(n11773), .Z(n11916) );
  XOR U16819 ( .A(n11764), .B(n11768), .Z(n11917) );
  XOR U16820 ( .A(n11759), .B(n11763), .Z(n11918) );
  XOR U16821 ( .A(n11754), .B(n11758), .Z(n11919) );
  XOR U16822 ( .A(n11749), .B(n11753), .Z(n11920) );
  XOR U16823 ( .A(n11744), .B(n11748), .Z(n11921) );
  XOR U16824 ( .A(n11739), .B(n11743), .Z(n11922) );
  XOR U16825 ( .A(n11734), .B(n11738), .Z(n11923) );
  XOR U16826 ( .A(n11729), .B(n11733), .Z(n11924) );
  XOR U16827 ( .A(n11724), .B(n11728), .Z(n11925) );
  XOR U16828 ( .A(n11719), .B(n11723), .Z(n11926) );
  XOR U16829 ( .A(n11714), .B(n11718), .Z(n11927) );
  XOR U16830 ( .A(n11709), .B(n11713), .Z(n11928) );
  XOR U16831 ( .A(n11704), .B(n11708), .Z(n11929) );
  XOR U16832 ( .A(n11699), .B(n11703), .Z(n11930) );
  XOR U16833 ( .A(n11694), .B(n11698), .Z(n11931) );
  XOR U16834 ( .A(n11689), .B(n11693), .Z(n11932) );
  XOR U16835 ( .A(n11684), .B(n11688), .Z(n11933) );
  XOR U16836 ( .A(n11679), .B(n11683), .Z(n11934) );
  XOR U16837 ( .A(n11674), .B(n11678), .Z(n11935) );
  XOR U16838 ( .A(n11669), .B(n11673), .Z(n11936) );
  XOR U16839 ( .A(n11664), .B(n11668), .Z(n11937) );
  XOR U16840 ( .A(n11659), .B(n11663), .Z(n11938) );
  XOR U16841 ( .A(n11654), .B(n11658), .Z(n11939) );
  XOR U16842 ( .A(n11649), .B(n11653), .Z(n11940) );
  XOR U16843 ( .A(n11644), .B(n11648), .Z(n11941) );
  XOR U16844 ( .A(n11639), .B(n11643), .Z(n11942) );
  XOR U16845 ( .A(n11634), .B(n11638), .Z(n11943) );
  XOR U16846 ( .A(n11629), .B(n11633), .Z(n11944) );
  XOR U16847 ( .A(n11624), .B(n11628), .Z(n11945) );
  XOR U16848 ( .A(n11619), .B(n11623), .Z(n11946) );
  XOR U16849 ( .A(n11614), .B(n11618), .Z(n11947) );
  XOR U16850 ( .A(n11609), .B(n11613), .Z(n11948) );
  XOR U16851 ( .A(n11604), .B(n11608), .Z(n11949) );
  XOR U16852 ( .A(n11594), .B(n11603), .Z(n11950) );
  XOR U16853 ( .A(n11951), .B(n11593), .Z(n11594) );
  AND U16854 ( .A(a[36]), .B(b[59]), .Z(n11951) );
  XOR U16855 ( .A(n11593), .B(n11600), .Z(n11952) );
  XOR U16856 ( .A(n11953), .B(n11954), .Z(n11600) );
  XOR U16857 ( .A(n11598), .B(n11955), .Z(n11954) );
  XOR U16858 ( .A(n11956), .B(n11957), .Z(n11955) );
  XOR U16859 ( .A(n11958), .B(n11959), .Z(n11957) );
  NAND U16860 ( .A(a[33]), .B(b[62]), .Z(n11959) );
  AND U16861 ( .A(a[32]), .B(b[63]), .Z(n11958) );
  XOR U16862 ( .A(n11960), .B(n11956), .Z(n11953) );
  XOR U16863 ( .A(n11961), .B(n11962), .Z(n11956) );
  ANDN U16864 ( .B(n11963), .A(n11964), .Z(n11961) );
  AND U16865 ( .A(a[34]), .B(b[61]), .Z(n11960) );
  XOR U16866 ( .A(n11965), .B(n11966), .Z(n11593) );
  AND U16867 ( .A(n11967), .B(n11968), .Z(n11965) );
  XOR U16868 ( .A(n11969), .B(n11598), .Z(n11599) );
  XOR U16869 ( .A(n11970), .B(n11971), .Z(n11598) );
  AND U16870 ( .A(n11972), .B(n11973), .Z(n11970) );
  AND U16871 ( .A(a[35]), .B(b[60]), .Z(n11969) );
  XOR U16872 ( .A(n11975), .B(n11976), .Z(n11603) );
  AND U16873 ( .A(n11977), .B(n11978), .Z(n11975) );
  AND U16874 ( .A(a[37]), .B(b[58]), .Z(n11974) );
  XOR U16875 ( .A(n11980), .B(n11981), .Z(n11608) );
  AND U16876 ( .A(n11982), .B(n11983), .Z(n11980) );
  AND U16877 ( .A(a[38]), .B(b[57]), .Z(n11979) );
  XOR U16878 ( .A(n11985), .B(n11986), .Z(n11613) );
  AND U16879 ( .A(n11987), .B(n11988), .Z(n11985) );
  AND U16880 ( .A(a[39]), .B(b[56]), .Z(n11984) );
  XOR U16881 ( .A(n11990), .B(n11991), .Z(n11618) );
  AND U16882 ( .A(n11992), .B(n11993), .Z(n11990) );
  AND U16883 ( .A(a[40]), .B(b[55]), .Z(n11989) );
  XOR U16884 ( .A(n11995), .B(n11996), .Z(n11623) );
  AND U16885 ( .A(n11997), .B(n11998), .Z(n11995) );
  AND U16886 ( .A(a[41]), .B(b[54]), .Z(n11994) );
  XOR U16887 ( .A(n12000), .B(n12001), .Z(n11628) );
  AND U16888 ( .A(n12002), .B(n12003), .Z(n12000) );
  AND U16889 ( .A(a[42]), .B(b[53]), .Z(n11999) );
  XOR U16890 ( .A(n12005), .B(n12006), .Z(n11633) );
  AND U16891 ( .A(n12007), .B(n12008), .Z(n12005) );
  AND U16892 ( .A(a[43]), .B(b[52]), .Z(n12004) );
  XOR U16893 ( .A(n12010), .B(n12011), .Z(n11638) );
  AND U16894 ( .A(n12012), .B(n12013), .Z(n12010) );
  AND U16895 ( .A(a[44]), .B(b[51]), .Z(n12009) );
  XOR U16896 ( .A(n12015), .B(n12016), .Z(n11643) );
  AND U16897 ( .A(n12017), .B(n12018), .Z(n12015) );
  AND U16898 ( .A(a[45]), .B(b[50]), .Z(n12014) );
  XOR U16899 ( .A(n12020), .B(n12021), .Z(n11648) );
  AND U16900 ( .A(n12022), .B(n12023), .Z(n12020) );
  AND U16901 ( .A(a[46]), .B(b[49]), .Z(n12019) );
  XOR U16902 ( .A(n12025), .B(n12026), .Z(n11653) );
  AND U16903 ( .A(n12027), .B(n12028), .Z(n12025) );
  AND U16904 ( .A(a[47]), .B(b[48]), .Z(n12024) );
  XOR U16905 ( .A(n12030), .B(n12031), .Z(n11658) );
  AND U16906 ( .A(n12032), .B(n12033), .Z(n12030) );
  AND U16907 ( .A(b[47]), .B(a[48]), .Z(n12029) );
  XOR U16908 ( .A(n12035), .B(n12036), .Z(n11663) );
  AND U16909 ( .A(n12037), .B(n12038), .Z(n12035) );
  AND U16910 ( .A(b[46]), .B(a[49]), .Z(n12034) );
  XOR U16911 ( .A(n12040), .B(n12041), .Z(n11668) );
  AND U16912 ( .A(n12042), .B(n12043), .Z(n12040) );
  AND U16913 ( .A(b[45]), .B(a[50]), .Z(n12039) );
  XOR U16914 ( .A(n12045), .B(n12046), .Z(n11673) );
  AND U16915 ( .A(n12047), .B(n12048), .Z(n12045) );
  AND U16916 ( .A(b[44]), .B(a[51]), .Z(n12044) );
  XOR U16917 ( .A(n12050), .B(n12051), .Z(n11678) );
  AND U16918 ( .A(n12052), .B(n12053), .Z(n12050) );
  AND U16919 ( .A(b[43]), .B(a[52]), .Z(n12049) );
  XOR U16920 ( .A(n12055), .B(n12056), .Z(n11683) );
  AND U16921 ( .A(n12057), .B(n12058), .Z(n12055) );
  AND U16922 ( .A(b[42]), .B(a[53]), .Z(n12054) );
  XOR U16923 ( .A(n12060), .B(n12061), .Z(n11688) );
  AND U16924 ( .A(n12062), .B(n12063), .Z(n12060) );
  AND U16925 ( .A(b[41]), .B(a[54]), .Z(n12059) );
  XOR U16926 ( .A(n12065), .B(n12066), .Z(n11693) );
  AND U16927 ( .A(n12067), .B(n12068), .Z(n12065) );
  AND U16928 ( .A(b[40]), .B(a[55]), .Z(n12064) );
  XOR U16929 ( .A(n12070), .B(n12071), .Z(n11698) );
  AND U16930 ( .A(n12072), .B(n12073), .Z(n12070) );
  AND U16931 ( .A(b[39]), .B(a[56]), .Z(n12069) );
  XOR U16932 ( .A(n12075), .B(n12076), .Z(n11703) );
  AND U16933 ( .A(n12077), .B(n12078), .Z(n12075) );
  AND U16934 ( .A(b[38]), .B(a[57]), .Z(n12074) );
  XOR U16935 ( .A(n12080), .B(n12081), .Z(n11708) );
  AND U16936 ( .A(n12082), .B(n12083), .Z(n12080) );
  AND U16937 ( .A(b[37]), .B(a[58]), .Z(n12079) );
  XOR U16938 ( .A(n12085), .B(n12086), .Z(n11713) );
  AND U16939 ( .A(n12087), .B(n12088), .Z(n12085) );
  AND U16940 ( .A(b[36]), .B(a[59]), .Z(n12084) );
  XOR U16941 ( .A(n12090), .B(n12091), .Z(n11718) );
  AND U16942 ( .A(n12092), .B(n12093), .Z(n12090) );
  AND U16943 ( .A(b[35]), .B(a[60]), .Z(n12089) );
  XOR U16944 ( .A(n12095), .B(n12096), .Z(n11723) );
  AND U16945 ( .A(n12097), .B(n12098), .Z(n12095) );
  AND U16946 ( .A(b[34]), .B(a[61]), .Z(n12094) );
  XOR U16947 ( .A(n12100), .B(n12101), .Z(n11728) );
  AND U16948 ( .A(n12102), .B(n12103), .Z(n12100) );
  AND U16949 ( .A(b[33]), .B(a[62]), .Z(n12099) );
  XOR U16950 ( .A(n12105), .B(n12106), .Z(n11733) );
  AND U16951 ( .A(n12107), .B(n12108), .Z(n12105) );
  AND U16952 ( .A(b[32]), .B(a[63]), .Z(n12104) );
  XOR U16953 ( .A(n12110), .B(n12111), .Z(n11738) );
  AND U16954 ( .A(n12112), .B(n12113), .Z(n12110) );
  AND U16955 ( .A(b[31]), .B(a[64]), .Z(n12109) );
  XOR U16956 ( .A(n12115), .B(n12116), .Z(n11743) );
  AND U16957 ( .A(n12117), .B(n12118), .Z(n12115) );
  AND U16958 ( .A(b[30]), .B(a[65]), .Z(n12114) );
  XOR U16959 ( .A(n12120), .B(n12121), .Z(n11748) );
  AND U16960 ( .A(n12122), .B(n12123), .Z(n12120) );
  AND U16961 ( .A(b[29]), .B(a[66]), .Z(n12119) );
  XOR U16962 ( .A(n12125), .B(n12126), .Z(n11753) );
  AND U16963 ( .A(n12127), .B(n12128), .Z(n12125) );
  AND U16964 ( .A(b[28]), .B(a[67]), .Z(n12124) );
  XOR U16965 ( .A(n12130), .B(n12131), .Z(n11758) );
  AND U16966 ( .A(n12132), .B(n12133), .Z(n12130) );
  AND U16967 ( .A(b[27]), .B(a[68]), .Z(n12129) );
  XOR U16968 ( .A(n12135), .B(n12136), .Z(n11763) );
  AND U16969 ( .A(n12137), .B(n12138), .Z(n12135) );
  AND U16970 ( .A(b[26]), .B(a[69]), .Z(n12134) );
  XOR U16971 ( .A(n12140), .B(n12141), .Z(n11768) );
  AND U16972 ( .A(n12142), .B(n12143), .Z(n12140) );
  AND U16973 ( .A(b[25]), .B(a[70]), .Z(n12139) );
  XOR U16974 ( .A(n12145), .B(n12146), .Z(n11773) );
  AND U16975 ( .A(n12147), .B(n12148), .Z(n12145) );
  AND U16976 ( .A(b[24]), .B(a[71]), .Z(n12144) );
  XOR U16977 ( .A(n12150), .B(n12151), .Z(n11778) );
  AND U16978 ( .A(n12152), .B(n12153), .Z(n12150) );
  AND U16979 ( .A(b[23]), .B(a[72]), .Z(n12149) );
  XOR U16980 ( .A(n12155), .B(n12156), .Z(n11783) );
  AND U16981 ( .A(n12157), .B(n12158), .Z(n12155) );
  AND U16982 ( .A(b[22]), .B(a[73]), .Z(n12154) );
  XOR U16983 ( .A(n12160), .B(n12161), .Z(n11788) );
  AND U16984 ( .A(n12162), .B(n12163), .Z(n12160) );
  AND U16985 ( .A(b[21]), .B(a[74]), .Z(n12159) );
  XOR U16986 ( .A(n12165), .B(n12166), .Z(n11793) );
  AND U16987 ( .A(n12167), .B(n12168), .Z(n12165) );
  AND U16988 ( .A(b[20]), .B(a[75]), .Z(n12164) );
  XOR U16989 ( .A(n12170), .B(n12171), .Z(n11798) );
  AND U16990 ( .A(n12172), .B(n12173), .Z(n12170) );
  AND U16991 ( .A(b[19]), .B(a[76]), .Z(n12169) );
  XOR U16992 ( .A(n12175), .B(n12176), .Z(n11803) );
  AND U16993 ( .A(n12177), .B(n12178), .Z(n12175) );
  AND U16994 ( .A(b[18]), .B(a[77]), .Z(n12174) );
  XOR U16995 ( .A(n12180), .B(n12181), .Z(n11808) );
  AND U16996 ( .A(n12182), .B(n12183), .Z(n12180) );
  AND U16997 ( .A(b[17]), .B(a[78]), .Z(n12179) );
  XOR U16998 ( .A(n12185), .B(n12186), .Z(n11813) );
  AND U16999 ( .A(n12187), .B(n12188), .Z(n12185) );
  AND U17000 ( .A(b[16]), .B(a[79]), .Z(n12184) );
  XOR U17001 ( .A(n12190), .B(n12191), .Z(n11818) );
  AND U17002 ( .A(n12192), .B(n12193), .Z(n12190) );
  AND U17003 ( .A(b[15]), .B(a[80]), .Z(n12189) );
  XOR U17004 ( .A(n12195), .B(n12196), .Z(n11823) );
  AND U17005 ( .A(n12197), .B(n12198), .Z(n12195) );
  AND U17006 ( .A(b[14]), .B(a[81]), .Z(n12194) );
  XOR U17007 ( .A(n12200), .B(n12201), .Z(n11828) );
  AND U17008 ( .A(n12202), .B(n12203), .Z(n12200) );
  AND U17009 ( .A(b[13]), .B(a[82]), .Z(n12199) );
  XOR U17010 ( .A(n12205), .B(n12206), .Z(n11833) );
  AND U17011 ( .A(n12207), .B(n12208), .Z(n12205) );
  AND U17012 ( .A(b[12]), .B(a[83]), .Z(n12204) );
  XOR U17013 ( .A(n12210), .B(n12211), .Z(n11838) );
  AND U17014 ( .A(n12212), .B(n12213), .Z(n12210) );
  AND U17015 ( .A(b[11]), .B(a[84]), .Z(n12209) );
  XOR U17016 ( .A(n12215), .B(n12216), .Z(n11843) );
  AND U17017 ( .A(n12217), .B(n12218), .Z(n12215) );
  AND U17018 ( .A(b[10]), .B(a[85]), .Z(n12214) );
  XOR U17019 ( .A(n12220), .B(n12221), .Z(n11848) );
  AND U17020 ( .A(n12222), .B(n12223), .Z(n12220) );
  AND U17021 ( .A(b[9]), .B(a[86]), .Z(n12219) );
  XOR U17022 ( .A(n12225), .B(n12226), .Z(n11853) );
  AND U17023 ( .A(n12227), .B(n12228), .Z(n12225) );
  AND U17024 ( .A(b[8]), .B(a[87]), .Z(n12224) );
  XOR U17025 ( .A(n12230), .B(n12231), .Z(n11858) );
  AND U17026 ( .A(n12232), .B(n12233), .Z(n12230) );
  AND U17027 ( .A(b[7]), .B(a[88]), .Z(n12229) );
  XOR U17028 ( .A(n12235), .B(n12236), .Z(n11863) );
  AND U17029 ( .A(n12237), .B(n12238), .Z(n12235) );
  AND U17030 ( .A(b[6]), .B(a[89]), .Z(n12234) );
  XOR U17031 ( .A(n12240), .B(n12241), .Z(n11868) );
  AND U17032 ( .A(n12242), .B(n12243), .Z(n12240) );
  AND U17033 ( .A(b[5]), .B(a[90]), .Z(n12239) );
  XOR U17034 ( .A(n12245), .B(n12246), .Z(n11873) );
  AND U17035 ( .A(n12247), .B(n12248), .Z(n12245) );
  AND U17036 ( .A(b[4]), .B(a[91]), .Z(n12244) );
  XOR U17037 ( .A(n12250), .B(n12251), .Z(n11878) );
  AND U17038 ( .A(n12252), .B(n12253), .Z(n12250) );
  AND U17039 ( .A(b[3]), .B(a[92]), .Z(n12249) );
  XOR U17040 ( .A(n12255), .B(n12256), .Z(n11883) );
  OR U17041 ( .A(n12257), .B(n12258), .Z(n12256) );
  AND U17042 ( .A(b[2]), .B(a[93]), .Z(n12254) );
  XNOR U17043 ( .A(n11893), .B(n12259), .Z(n11889) );
  NAND U17044 ( .A(b[1]), .B(a[94]), .Z(n12259) );
  IV U17045 ( .A(n11887), .Z(n11893) );
  ANDN U17046 ( .B(n10269), .A(n10271), .Z(n11887) );
  NAND U17047 ( .A(a[94]), .B(b[0]), .Z(n10271) );
  XOR U17048 ( .A(n12257), .B(n12258), .Z(n10269) );
  XOR U17049 ( .A(n12261), .B(n12252), .Z(n12260) );
  XOR U17050 ( .A(n12247), .B(n12251), .Z(n12262) );
  XOR U17051 ( .A(n12242), .B(n12246), .Z(n12263) );
  XOR U17052 ( .A(n12237), .B(n12241), .Z(n12264) );
  XOR U17053 ( .A(n12232), .B(n12236), .Z(n12265) );
  XOR U17054 ( .A(n12227), .B(n12231), .Z(n12266) );
  XOR U17055 ( .A(n12222), .B(n12226), .Z(n12267) );
  XOR U17056 ( .A(n12217), .B(n12221), .Z(n12268) );
  XOR U17057 ( .A(n12212), .B(n12216), .Z(n12269) );
  XOR U17058 ( .A(n12207), .B(n12211), .Z(n12270) );
  XOR U17059 ( .A(n12202), .B(n12206), .Z(n12271) );
  XOR U17060 ( .A(n12197), .B(n12201), .Z(n12272) );
  XOR U17061 ( .A(n12192), .B(n12196), .Z(n12273) );
  XOR U17062 ( .A(n12187), .B(n12191), .Z(n12274) );
  XOR U17063 ( .A(n12182), .B(n12186), .Z(n12275) );
  XOR U17064 ( .A(n12177), .B(n12181), .Z(n12276) );
  XOR U17065 ( .A(n12172), .B(n12176), .Z(n12277) );
  XOR U17066 ( .A(n12167), .B(n12171), .Z(n12278) );
  XOR U17067 ( .A(n12162), .B(n12166), .Z(n12279) );
  XOR U17068 ( .A(n12157), .B(n12161), .Z(n12280) );
  XOR U17069 ( .A(n12152), .B(n12156), .Z(n12281) );
  XOR U17070 ( .A(n12147), .B(n12151), .Z(n12282) );
  XOR U17071 ( .A(n12142), .B(n12146), .Z(n12283) );
  XOR U17072 ( .A(n12137), .B(n12141), .Z(n12284) );
  XOR U17073 ( .A(n12132), .B(n12136), .Z(n12285) );
  XOR U17074 ( .A(n12127), .B(n12131), .Z(n12286) );
  XOR U17075 ( .A(n12122), .B(n12126), .Z(n12287) );
  XOR U17076 ( .A(n12117), .B(n12121), .Z(n12288) );
  XOR U17077 ( .A(n12112), .B(n12116), .Z(n12289) );
  XOR U17078 ( .A(n12107), .B(n12111), .Z(n12290) );
  XOR U17079 ( .A(n12102), .B(n12106), .Z(n12291) );
  XOR U17080 ( .A(n12097), .B(n12101), .Z(n12292) );
  XOR U17081 ( .A(n12092), .B(n12096), .Z(n12293) );
  XOR U17082 ( .A(n12087), .B(n12091), .Z(n12294) );
  XOR U17083 ( .A(n12082), .B(n12086), .Z(n12295) );
  XOR U17084 ( .A(n12077), .B(n12081), .Z(n12296) );
  XOR U17085 ( .A(n12072), .B(n12076), .Z(n12297) );
  XOR U17086 ( .A(n12067), .B(n12071), .Z(n12298) );
  XOR U17087 ( .A(n12062), .B(n12066), .Z(n12299) );
  XOR U17088 ( .A(n12057), .B(n12061), .Z(n12300) );
  XOR U17089 ( .A(n12052), .B(n12056), .Z(n12301) );
  XOR U17090 ( .A(n12047), .B(n12051), .Z(n12302) );
  XOR U17091 ( .A(n12042), .B(n12046), .Z(n12303) );
  XOR U17092 ( .A(n12037), .B(n12041), .Z(n12304) );
  XOR U17093 ( .A(n12032), .B(n12036), .Z(n12305) );
  XOR U17094 ( .A(n12027), .B(n12031), .Z(n12306) );
  XOR U17095 ( .A(n12022), .B(n12026), .Z(n12307) );
  XOR U17096 ( .A(n12017), .B(n12021), .Z(n12308) );
  XOR U17097 ( .A(n12012), .B(n12016), .Z(n12309) );
  XOR U17098 ( .A(n12007), .B(n12011), .Z(n12310) );
  XOR U17099 ( .A(n12002), .B(n12006), .Z(n12311) );
  XOR U17100 ( .A(n11997), .B(n12001), .Z(n12312) );
  XOR U17101 ( .A(n11992), .B(n11996), .Z(n12313) );
  XOR U17102 ( .A(n11987), .B(n11991), .Z(n12314) );
  XOR U17103 ( .A(n11982), .B(n11986), .Z(n12315) );
  XOR U17104 ( .A(n11977), .B(n11981), .Z(n12316) );
  XOR U17105 ( .A(n11967), .B(n11976), .Z(n12317) );
  XOR U17106 ( .A(n12318), .B(n11966), .Z(n11967) );
  AND U17107 ( .A(a[36]), .B(b[58]), .Z(n12318) );
  XNOR U17108 ( .A(n11966), .B(n11972), .Z(n12319) );
  XOR U17109 ( .A(n11971), .B(n11964), .Z(n12320) );
  XOR U17110 ( .A(n12321), .B(n12322), .Z(n11964) );
  XOR U17111 ( .A(n11962), .B(n12323), .Z(n12322) );
  XOR U17112 ( .A(n12324), .B(n12325), .Z(n12323) );
  XOR U17113 ( .A(n12326), .B(n12327), .Z(n12325) );
  NAND U17114 ( .A(a[32]), .B(b[62]), .Z(n12327) );
  AND U17115 ( .A(a[31]), .B(b[63]), .Z(n12326) );
  XOR U17116 ( .A(n12328), .B(n12324), .Z(n12321) );
  XOR U17117 ( .A(n12329), .B(n12330), .Z(n12324) );
  ANDN U17118 ( .B(n12331), .A(n12332), .Z(n12329) );
  AND U17119 ( .A(a[33]), .B(b[61]), .Z(n12328) );
  XOR U17120 ( .A(n12333), .B(n11962), .Z(n11963) );
  XOR U17121 ( .A(n12334), .B(n12335), .Z(n11962) );
  AND U17122 ( .A(n12336), .B(n12337), .Z(n12334) );
  AND U17123 ( .A(a[34]), .B(b[60]), .Z(n12333) );
  XOR U17124 ( .A(n12338), .B(n12339), .Z(n11966) );
  AND U17125 ( .A(n12340), .B(n12341), .Z(n12338) );
  XOR U17126 ( .A(n12342), .B(n11971), .Z(n11973) );
  XOR U17127 ( .A(n12343), .B(n12344), .Z(n11971) );
  AND U17128 ( .A(n12345), .B(n12346), .Z(n12343) );
  AND U17129 ( .A(a[35]), .B(b[59]), .Z(n12342) );
  XOR U17130 ( .A(n12348), .B(n12349), .Z(n11976) );
  AND U17131 ( .A(n12350), .B(n12351), .Z(n12348) );
  AND U17132 ( .A(a[37]), .B(b[57]), .Z(n12347) );
  XOR U17133 ( .A(n12353), .B(n12354), .Z(n11981) );
  AND U17134 ( .A(n12355), .B(n12356), .Z(n12353) );
  AND U17135 ( .A(a[38]), .B(b[56]), .Z(n12352) );
  XOR U17136 ( .A(n12358), .B(n12359), .Z(n11986) );
  AND U17137 ( .A(n12360), .B(n12361), .Z(n12358) );
  AND U17138 ( .A(a[39]), .B(b[55]), .Z(n12357) );
  XOR U17139 ( .A(n12363), .B(n12364), .Z(n11991) );
  AND U17140 ( .A(n12365), .B(n12366), .Z(n12363) );
  AND U17141 ( .A(a[40]), .B(b[54]), .Z(n12362) );
  XOR U17142 ( .A(n12368), .B(n12369), .Z(n11996) );
  AND U17143 ( .A(n12370), .B(n12371), .Z(n12368) );
  AND U17144 ( .A(a[41]), .B(b[53]), .Z(n12367) );
  XOR U17145 ( .A(n12373), .B(n12374), .Z(n12001) );
  AND U17146 ( .A(n12375), .B(n12376), .Z(n12373) );
  AND U17147 ( .A(a[42]), .B(b[52]), .Z(n12372) );
  XOR U17148 ( .A(n12378), .B(n12379), .Z(n12006) );
  AND U17149 ( .A(n12380), .B(n12381), .Z(n12378) );
  AND U17150 ( .A(a[43]), .B(b[51]), .Z(n12377) );
  XOR U17151 ( .A(n12383), .B(n12384), .Z(n12011) );
  AND U17152 ( .A(n12385), .B(n12386), .Z(n12383) );
  AND U17153 ( .A(a[44]), .B(b[50]), .Z(n12382) );
  XOR U17154 ( .A(n12388), .B(n12389), .Z(n12016) );
  AND U17155 ( .A(n12390), .B(n12391), .Z(n12388) );
  AND U17156 ( .A(a[45]), .B(b[49]), .Z(n12387) );
  XOR U17157 ( .A(n12393), .B(n12394), .Z(n12021) );
  AND U17158 ( .A(n12395), .B(n12396), .Z(n12393) );
  AND U17159 ( .A(a[46]), .B(b[48]), .Z(n12392) );
  XOR U17160 ( .A(n12398), .B(n12399), .Z(n12026) );
  AND U17161 ( .A(n12400), .B(n12401), .Z(n12398) );
  AND U17162 ( .A(a[47]), .B(b[47]), .Z(n12397) );
  XOR U17163 ( .A(n12403), .B(n12404), .Z(n12031) );
  AND U17164 ( .A(n12405), .B(n12406), .Z(n12403) );
  AND U17165 ( .A(b[46]), .B(a[48]), .Z(n12402) );
  XOR U17166 ( .A(n12408), .B(n12409), .Z(n12036) );
  AND U17167 ( .A(n12410), .B(n12411), .Z(n12408) );
  AND U17168 ( .A(b[45]), .B(a[49]), .Z(n12407) );
  XOR U17169 ( .A(n12413), .B(n12414), .Z(n12041) );
  AND U17170 ( .A(n12415), .B(n12416), .Z(n12413) );
  AND U17171 ( .A(b[44]), .B(a[50]), .Z(n12412) );
  XOR U17172 ( .A(n12418), .B(n12419), .Z(n12046) );
  AND U17173 ( .A(n12420), .B(n12421), .Z(n12418) );
  AND U17174 ( .A(b[43]), .B(a[51]), .Z(n12417) );
  XOR U17175 ( .A(n12423), .B(n12424), .Z(n12051) );
  AND U17176 ( .A(n12425), .B(n12426), .Z(n12423) );
  AND U17177 ( .A(b[42]), .B(a[52]), .Z(n12422) );
  XOR U17178 ( .A(n12428), .B(n12429), .Z(n12056) );
  AND U17179 ( .A(n12430), .B(n12431), .Z(n12428) );
  AND U17180 ( .A(b[41]), .B(a[53]), .Z(n12427) );
  XOR U17181 ( .A(n12433), .B(n12434), .Z(n12061) );
  AND U17182 ( .A(n12435), .B(n12436), .Z(n12433) );
  AND U17183 ( .A(b[40]), .B(a[54]), .Z(n12432) );
  XOR U17184 ( .A(n12438), .B(n12439), .Z(n12066) );
  AND U17185 ( .A(n12440), .B(n12441), .Z(n12438) );
  AND U17186 ( .A(b[39]), .B(a[55]), .Z(n12437) );
  XOR U17187 ( .A(n12443), .B(n12444), .Z(n12071) );
  AND U17188 ( .A(n12445), .B(n12446), .Z(n12443) );
  AND U17189 ( .A(b[38]), .B(a[56]), .Z(n12442) );
  XOR U17190 ( .A(n12448), .B(n12449), .Z(n12076) );
  AND U17191 ( .A(n12450), .B(n12451), .Z(n12448) );
  AND U17192 ( .A(b[37]), .B(a[57]), .Z(n12447) );
  XOR U17193 ( .A(n12453), .B(n12454), .Z(n12081) );
  AND U17194 ( .A(n12455), .B(n12456), .Z(n12453) );
  AND U17195 ( .A(b[36]), .B(a[58]), .Z(n12452) );
  XOR U17196 ( .A(n12458), .B(n12459), .Z(n12086) );
  AND U17197 ( .A(n12460), .B(n12461), .Z(n12458) );
  AND U17198 ( .A(b[35]), .B(a[59]), .Z(n12457) );
  XOR U17199 ( .A(n12463), .B(n12464), .Z(n12091) );
  AND U17200 ( .A(n12465), .B(n12466), .Z(n12463) );
  AND U17201 ( .A(b[34]), .B(a[60]), .Z(n12462) );
  XOR U17202 ( .A(n12468), .B(n12469), .Z(n12096) );
  AND U17203 ( .A(n12470), .B(n12471), .Z(n12468) );
  AND U17204 ( .A(b[33]), .B(a[61]), .Z(n12467) );
  XOR U17205 ( .A(n12473), .B(n12474), .Z(n12101) );
  AND U17206 ( .A(n12475), .B(n12476), .Z(n12473) );
  AND U17207 ( .A(b[32]), .B(a[62]), .Z(n12472) );
  XOR U17208 ( .A(n12478), .B(n12479), .Z(n12106) );
  AND U17209 ( .A(n12480), .B(n12481), .Z(n12478) );
  AND U17210 ( .A(b[31]), .B(a[63]), .Z(n12477) );
  XOR U17211 ( .A(n12483), .B(n12484), .Z(n12111) );
  AND U17212 ( .A(n12485), .B(n12486), .Z(n12483) );
  AND U17213 ( .A(b[30]), .B(a[64]), .Z(n12482) );
  XOR U17214 ( .A(n12488), .B(n12489), .Z(n12116) );
  AND U17215 ( .A(n12490), .B(n12491), .Z(n12488) );
  AND U17216 ( .A(b[29]), .B(a[65]), .Z(n12487) );
  XOR U17217 ( .A(n12493), .B(n12494), .Z(n12121) );
  AND U17218 ( .A(n12495), .B(n12496), .Z(n12493) );
  AND U17219 ( .A(b[28]), .B(a[66]), .Z(n12492) );
  XOR U17220 ( .A(n12498), .B(n12499), .Z(n12126) );
  AND U17221 ( .A(n12500), .B(n12501), .Z(n12498) );
  AND U17222 ( .A(b[27]), .B(a[67]), .Z(n12497) );
  XOR U17223 ( .A(n12503), .B(n12504), .Z(n12131) );
  AND U17224 ( .A(n12505), .B(n12506), .Z(n12503) );
  AND U17225 ( .A(b[26]), .B(a[68]), .Z(n12502) );
  XOR U17226 ( .A(n12508), .B(n12509), .Z(n12136) );
  AND U17227 ( .A(n12510), .B(n12511), .Z(n12508) );
  AND U17228 ( .A(b[25]), .B(a[69]), .Z(n12507) );
  XOR U17229 ( .A(n12513), .B(n12514), .Z(n12141) );
  AND U17230 ( .A(n12515), .B(n12516), .Z(n12513) );
  AND U17231 ( .A(b[24]), .B(a[70]), .Z(n12512) );
  XOR U17232 ( .A(n12518), .B(n12519), .Z(n12146) );
  AND U17233 ( .A(n12520), .B(n12521), .Z(n12518) );
  AND U17234 ( .A(b[23]), .B(a[71]), .Z(n12517) );
  XOR U17235 ( .A(n12523), .B(n12524), .Z(n12151) );
  AND U17236 ( .A(n12525), .B(n12526), .Z(n12523) );
  AND U17237 ( .A(b[22]), .B(a[72]), .Z(n12522) );
  XOR U17238 ( .A(n12528), .B(n12529), .Z(n12156) );
  AND U17239 ( .A(n12530), .B(n12531), .Z(n12528) );
  AND U17240 ( .A(b[21]), .B(a[73]), .Z(n12527) );
  XOR U17241 ( .A(n12533), .B(n12534), .Z(n12161) );
  AND U17242 ( .A(n12535), .B(n12536), .Z(n12533) );
  AND U17243 ( .A(b[20]), .B(a[74]), .Z(n12532) );
  XOR U17244 ( .A(n12538), .B(n12539), .Z(n12166) );
  AND U17245 ( .A(n12540), .B(n12541), .Z(n12538) );
  AND U17246 ( .A(b[19]), .B(a[75]), .Z(n12537) );
  XOR U17247 ( .A(n12543), .B(n12544), .Z(n12171) );
  AND U17248 ( .A(n12545), .B(n12546), .Z(n12543) );
  AND U17249 ( .A(b[18]), .B(a[76]), .Z(n12542) );
  XOR U17250 ( .A(n12548), .B(n12549), .Z(n12176) );
  AND U17251 ( .A(n12550), .B(n12551), .Z(n12548) );
  AND U17252 ( .A(b[17]), .B(a[77]), .Z(n12547) );
  XOR U17253 ( .A(n12553), .B(n12554), .Z(n12181) );
  AND U17254 ( .A(n12555), .B(n12556), .Z(n12553) );
  AND U17255 ( .A(b[16]), .B(a[78]), .Z(n12552) );
  XOR U17256 ( .A(n12558), .B(n12559), .Z(n12186) );
  AND U17257 ( .A(n12560), .B(n12561), .Z(n12558) );
  AND U17258 ( .A(b[15]), .B(a[79]), .Z(n12557) );
  XOR U17259 ( .A(n12563), .B(n12564), .Z(n12191) );
  AND U17260 ( .A(n12565), .B(n12566), .Z(n12563) );
  AND U17261 ( .A(b[14]), .B(a[80]), .Z(n12562) );
  XOR U17262 ( .A(n12568), .B(n12569), .Z(n12196) );
  AND U17263 ( .A(n12570), .B(n12571), .Z(n12568) );
  AND U17264 ( .A(b[13]), .B(a[81]), .Z(n12567) );
  XOR U17265 ( .A(n12573), .B(n12574), .Z(n12201) );
  AND U17266 ( .A(n12575), .B(n12576), .Z(n12573) );
  AND U17267 ( .A(b[12]), .B(a[82]), .Z(n12572) );
  XOR U17268 ( .A(n12578), .B(n12579), .Z(n12206) );
  AND U17269 ( .A(n12580), .B(n12581), .Z(n12578) );
  AND U17270 ( .A(b[11]), .B(a[83]), .Z(n12577) );
  XOR U17271 ( .A(n12583), .B(n12584), .Z(n12211) );
  AND U17272 ( .A(n12585), .B(n12586), .Z(n12583) );
  AND U17273 ( .A(b[10]), .B(a[84]), .Z(n12582) );
  XOR U17274 ( .A(n12588), .B(n12589), .Z(n12216) );
  AND U17275 ( .A(n12590), .B(n12591), .Z(n12588) );
  AND U17276 ( .A(b[9]), .B(a[85]), .Z(n12587) );
  XOR U17277 ( .A(n12593), .B(n12594), .Z(n12221) );
  AND U17278 ( .A(n12595), .B(n12596), .Z(n12593) );
  AND U17279 ( .A(b[8]), .B(a[86]), .Z(n12592) );
  XOR U17280 ( .A(n12598), .B(n12599), .Z(n12226) );
  AND U17281 ( .A(n12600), .B(n12601), .Z(n12598) );
  AND U17282 ( .A(b[7]), .B(a[87]), .Z(n12597) );
  XOR U17283 ( .A(n12603), .B(n12604), .Z(n12231) );
  AND U17284 ( .A(n12605), .B(n12606), .Z(n12603) );
  AND U17285 ( .A(b[6]), .B(a[88]), .Z(n12602) );
  XOR U17286 ( .A(n12608), .B(n12609), .Z(n12236) );
  AND U17287 ( .A(n12610), .B(n12611), .Z(n12608) );
  AND U17288 ( .A(b[5]), .B(a[89]), .Z(n12607) );
  XOR U17289 ( .A(n12613), .B(n12614), .Z(n12241) );
  AND U17290 ( .A(n12615), .B(n12616), .Z(n12613) );
  AND U17291 ( .A(b[4]), .B(a[90]), .Z(n12612) );
  XOR U17292 ( .A(n12618), .B(n12619), .Z(n12246) );
  AND U17293 ( .A(n12620), .B(n12621), .Z(n12618) );
  AND U17294 ( .A(b[3]), .B(a[91]), .Z(n12617) );
  XOR U17295 ( .A(n12623), .B(n12624), .Z(n12251) );
  OR U17296 ( .A(n12625), .B(n12626), .Z(n12624) );
  AND U17297 ( .A(b[2]), .B(a[92]), .Z(n12622) );
  XNOR U17298 ( .A(n12261), .B(n12627), .Z(n12257) );
  NAND U17299 ( .A(b[1]), .B(a[93]), .Z(n12627) );
  IV U17300 ( .A(n12255), .Z(n12261) );
  ANDN U17301 ( .B(n10272), .A(n10274), .Z(n12255) );
  NAND U17302 ( .A(a[93]), .B(b[0]), .Z(n10274) );
  XOR U17303 ( .A(n12625), .B(n12626), .Z(n10272) );
  XOR U17304 ( .A(n12629), .B(n12620), .Z(n12628) );
  XOR U17305 ( .A(n12615), .B(n12619), .Z(n12630) );
  XOR U17306 ( .A(n12610), .B(n12614), .Z(n12631) );
  XOR U17307 ( .A(n12605), .B(n12609), .Z(n12632) );
  XOR U17308 ( .A(n12600), .B(n12604), .Z(n12633) );
  XOR U17309 ( .A(n12595), .B(n12599), .Z(n12634) );
  XOR U17310 ( .A(n12590), .B(n12594), .Z(n12635) );
  XOR U17311 ( .A(n12585), .B(n12589), .Z(n12636) );
  XOR U17312 ( .A(n12580), .B(n12584), .Z(n12637) );
  XOR U17313 ( .A(n12575), .B(n12579), .Z(n12638) );
  XOR U17314 ( .A(n12570), .B(n12574), .Z(n12639) );
  XOR U17315 ( .A(n12565), .B(n12569), .Z(n12640) );
  XOR U17316 ( .A(n12560), .B(n12564), .Z(n12641) );
  XOR U17317 ( .A(n12555), .B(n12559), .Z(n12642) );
  XOR U17318 ( .A(n12550), .B(n12554), .Z(n12643) );
  XOR U17319 ( .A(n12545), .B(n12549), .Z(n12644) );
  XOR U17320 ( .A(n12540), .B(n12544), .Z(n12645) );
  XOR U17321 ( .A(n12535), .B(n12539), .Z(n12646) );
  XOR U17322 ( .A(n12530), .B(n12534), .Z(n12647) );
  XOR U17323 ( .A(n12525), .B(n12529), .Z(n12648) );
  XOR U17324 ( .A(n12520), .B(n12524), .Z(n12649) );
  XOR U17325 ( .A(n12515), .B(n12519), .Z(n12650) );
  XOR U17326 ( .A(n12510), .B(n12514), .Z(n12651) );
  XOR U17327 ( .A(n12505), .B(n12509), .Z(n12652) );
  XOR U17328 ( .A(n12500), .B(n12504), .Z(n12653) );
  XOR U17329 ( .A(n12495), .B(n12499), .Z(n12654) );
  XOR U17330 ( .A(n12490), .B(n12494), .Z(n12655) );
  XOR U17331 ( .A(n12485), .B(n12489), .Z(n12656) );
  XOR U17332 ( .A(n12480), .B(n12484), .Z(n12657) );
  XOR U17333 ( .A(n12475), .B(n12479), .Z(n12658) );
  XOR U17334 ( .A(n12470), .B(n12474), .Z(n12659) );
  XOR U17335 ( .A(n12465), .B(n12469), .Z(n12660) );
  XOR U17336 ( .A(n12460), .B(n12464), .Z(n12661) );
  XOR U17337 ( .A(n12455), .B(n12459), .Z(n12662) );
  XOR U17338 ( .A(n12450), .B(n12454), .Z(n12663) );
  XOR U17339 ( .A(n12445), .B(n12449), .Z(n12664) );
  XOR U17340 ( .A(n12440), .B(n12444), .Z(n12665) );
  XOR U17341 ( .A(n12435), .B(n12439), .Z(n12666) );
  XOR U17342 ( .A(n12430), .B(n12434), .Z(n12667) );
  XOR U17343 ( .A(n12425), .B(n12429), .Z(n12668) );
  XOR U17344 ( .A(n12420), .B(n12424), .Z(n12669) );
  XOR U17345 ( .A(n12415), .B(n12419), .Z(n12670) );
  XOR U17346 ( .A(n12410), .B(n12414), .Z(n12671) );
  XOR U17347 ( .A(n12405), .B(n12409), .Z(n12672) );
  XOR U17348 ( .A(n12400), .B(n12404), .Z(n12673) );
  XOR U17349 ( .A(n12395), .B(n12399), .Z(n12674) );
  XOR U17350 ( .A(n12390), .B(n12394), .Z(n12675) );
  XOR U17351 ( .A(n12385), .B(n12389), .Z(n12676) );
  XOR U17352 ( .A(n12380), .B(n12384), .Z(n12677) );
  XOR U17353 ( .A(n12375), .B(n12379), .Z(n12678) );
  XOR U17354 ( .A(n12370), .B(n12374), .Z(n12679) );
  XOR U17355 ( .A(n12365), .B(n12369), .Z(n12680) );
  XOR U17356 ( .A(n12360), .B(n12364), .Z(n12681) );
  XOR U17357 ( .A(n12355), .B(n12359), .Z(n12682) );
  XOR U17358 ( .A(n12350), .B(n12354), .Z(n12683) );
  XOR U17359 ( .A(n12340), .B(n12349), .Z(n12684) );
  XOR U17360 ( .A(n12685), .B(n12339), .Z(n12340) );
  AND U17361 ( .A(a[36]), .B(b[57]), .Z(n12685) );
  XNOR U17362 ( .A(n12339), .B(n12345), .Z(n12686) );
  XNOR U17363 ( .A(n12344), .B(n12336), .Z(n12687) );
  XOR U17364 ( .A(n12335), .B(n12332), .Z(n12688) );
  XOR U17365 ( .A(n12689), .B(n12690), .Z(n12332) );
  XOR U17366 ( .A(n12330), .B(n12691), .Z(n12690) );
  XOR U17367 ( .A(n12692), .B(n12693), .Z(n12691) );
  XOR U17368 ( .A(n12694), .B(n12695), .Z(n12693) );
  NAND U17369 ( .A(a[31]), .B(b[62]), .Z(n12695) );
  AND U17370 ( .A(a[30]), .B(b[63]), .Z(n12694) );
  XOR U17371 ( .A(n12696), .B(n12692), .Z(n12689) );
  XOR U17372 ( .A(n12697), .B(n12698), .Z(n12692) );
  ANDN U17373 ( .B(n12699), .A(n12700), .Z(n12697) );
  AND U17374 ( .A(a[32]), .B(b[61]), .Z(n12696) );
  XOR U17375 ( .A(n12701), .B(n12330), .Z(n12331) );
  XOR U17376 ( .A(n12702), .B(n12703), .Z(n12330) );
  AND U17377 ( .A(n12704), .B(n12705), .Z(n12702) );
  AND U17378 ( .A(a[33]), .B(b[60]), .Z(n12701) );
  XOR U17379 ( .A(n12706), .B(n12335), .Z(n12337) );
  XOR U17380 ( .A(n12707), .B(n12708), .Z(n12335) );
  AND U17381 ( .A(n12709), .B(n12710), .Z(n12707) );
  AND U17382 ( .A(a[34]), .B(b[59]), .Z(n12706) );
  XOR U17383 ( .A(n12711), .B(n12712), .Z(n12339) );
  AND U17384 ( .A(n12713), .B(n12714), .Z(n12711) );
  XOR U17385 ( .A(n12715), .B(n12344), .Z(n12346) );
  XOR U17386 ( .A(n12716), .B(n12717), .Z(n12344) );
  AND U17387 ( .A(n12718), .B(n12719), .Z(n12716) );
  AND U17388 ( .A(a[35]), .B(b[58]), .Z(n12715) );
  XOR U17389 ( .A(n12721), .B(n12722), .Z(n12349) );
  AND U17390 ( .A(n12723), .B(n12724), .Z(n12721) );
  AND U17391 ( .A(a[37]), .B(b[56]), .Z(n12720) );
  XOR U17392 ( .A(n12726), .B(n12727), .Z(n12354) );
  AND U17393 ( .A(n12728), .B(n12729), .Z(n12726) );
  AND U17394 ( .A(a[38]), .B(b[55]), .Z(n12725) );
  XOR U17395 ( .A(n12731), .B(n12732), .Z(n12359) );
  AND U17396 ( .A(n12733), .B(n12734), .Z(n12731) );
  AND U17397 ( .A(a[39]), .B(b[54]), .Z(n12730) );
  XOR U17398 ( .A(n12736), .B(n12737), .Z(n12364) );
  AND U17399 ( .A(n12738), .B(n12739), .Z(n12736) );
  AND U17400 ( .A(a[40]), .B(b[53]), .Z(n12735) );
  XOR U17401 ( .A(n12741), .B(n12742), .Z(n12369) );
  AND U17402 ( .A(n12743), .B(n12744), .Z(n12741) );
  AND U17403 ( .A(a[41]), .B(b[52]), .Z(n12740) );
  XOR U17404 ( .A(n12746), .B(n12747), .Z(n12374) );
  AND U17405 ( .A(n12748), .B(n12749), .Z(n12746) );
  AND U17406 ( .A(a[42]), .B(b[51]), .Z(n12745) );
  XOR U17407 ( .A(n12751), .B(n12752), .Z(n12379) );
  AND U17408 ( .A(n12753), .B(n12754), .Z(n12751) );
  AND U17409 ( .A(a[43]), .B(b[50]), .Z(n12750) );
  XOR U17410 ( .A(n12756), .B(n12757), .Z(n12384) );
  AND U17411 ( .A(n12758), .B(n12759), .Z(n12756) );
  AND U17412 ( .A(a[44]), .B(b[49]), .Z(n12755) );
  XOR U17413 ( .A(n12761), .B(n12762), .Z(n12389) );
  AND U17414 ( .A(n12763), .B(n12764), .Z(n12761) );
  AND U17415 ( .A(a[45]), .B(b[48]), .Z(n12760) );
  XOR U17416 ( .A(n12766), .B(n12767), .Z(n12394) );
  AND U17417 ( .A(n12768), .B(n12769), .Z(n12766) );
  AND U17418 ( .A(a[46]), .B(b[47]), .Z(n12765) );
  XOR U17419 ( .A(n12771), .B(n12772), .Z(n12399) );
  AND U17420 ( .A(n12773), .B(n12774), .Z(n12771) );
  AND U17421 ( .A(b[46]), .B(a[47]), .Z(n12770) );
  XOR U17422 ( .A(n12776), .B(n12777), .Z(n12404) );
  AND U17423 ( .A(n12778), .B(n12779), .Z(n12776) );
  AND U17424 ( .A(b[45]), .B(a[48]), .Z(n12775) );
  XOR U17425 ( .A(n12781), .B(n12782), .Z(n12409) );
  AND U17426 ( .A(n12783), .B(n12784), .Z(n12781) );
  AND U17427 ( .A(b[44]), .B(a[49]), .Z(n12780) );
  XOR U17428 ( .A(n12786), .B(n12787), .Z(n12414) );
  AND U17429 ( .A(n12788), .B(n12789), .Z(n12786) );
  AND U17430 ( .A(b[43]), .B(a[50]), .Z(n12785) );
  XOR U17431 ( .A(n12791), .B(n12792), .Z(n12419) );
  AND U17432 ( .A(n12793), .B(n12794), .Z(n12791) );
  AND U17433 ( .A(b[42]), .B(a[51]), .Z(n12790) );
  XOR U17434 ( .A(n12796), .B(n12797), .Z(n12424) );
  AND U17435 ( .A(n12798), .B(n12799), .Z(n12796) );
  AND U17436 ( .A(b[41]), .B(a[52]), .Z(n12795) );
  XOR U17437 ( .A(n12801), .B(n12802), .Z(n12429) );
  AND U17438 ( .A(n12803), .B(n12804), .Z(n12801) );
  AND U17439 ( .A(b[40]), .B(a[53]), .Z(n12800) );
  XOR U17440 ( .A(n12806), .B(n12807), .Z(n12434) );
  AND U17441 ( .A(n12808), .B(n12809), .Z(n12806) );
  AND U17442 ( .A(b[39]), .B(a[54]), .Z(n12805) );
  XOR U17443 ( .A(n12811), .B(n12812), .Z(n12439) );
  AND U17444 ( .A(n12813), .B(n12814), .Z(n12811) );
  AND U17445 ( .A(b[38]), .B(a[55]), .Z(n12810) );
  XOR U17446 ( .A(n12816), .B(n12817), .Z(n12444) );
  AND U17447 ( .A(n12818), .B(n12819), .Z(n12816) );
  AND U17448 ( .A(b[37]), .B(a[56]), .Z(n12815) );
  XOR U17449 ( .A(n12821), .B(n12822), .Z(n12449) );
  AND U17450 ( .A(n12823), .B(n12824), .Z(n12821) );
  AND U17451 ( .A(b[36]), .B(a[57]), .Z(n12820) );
  XOR U17452 ( .A(n12826), .B(n12827), .Z(n12454) );
  AND U17453 ( .A(n12828), .B(n12829), .Z(n12826) );
  AND U17454 ( .A(b[35]), .B(a[58]), .Z(n12825) );
  XOR U17455 ( .A(n12831), .B(n12832), .Z(n12459) );
  AND U17456 ( .A(n12833), .B(n12834), .Z(n12831) );
  AND U17457 ( .A(b[34]), .B(a[59]), .Z(n12830) );
  XOR U17458 ( .A(n12836), .B(n12837), .Z(n12464) );
  AND U17459 ( .A(n12838), .B(n12839), .Z(n12836) );
  AND U17460 ( .A(b[33]), .B(a[60]), .Z(n12835) );
  XOR U17461 ( .A(n12841), .B(n12842), .Z(n12469) );
  AND U17462 ( .A(n12843), .B(n12844), .Z(n12841) );
  AND U17463 ( .A(b[32]), .B(a[61]), .Z(n12840) );
  XOR U17464 ( .A(n12846), .B(n12847), .Z(n12474) );
  AND U17465 ( .A(n12848), .B(n12849), .Z(n12846) );
  AND U17466 ( .A(b[31]), .B(a[62]), .Z(n12845) );
  XOR U17467 ( .A(n12851), .B(n12852), .Z(n12479) );
  AND U17468 ( .A(n12853), .B(n12854), .Z(n12851) );
  AND U17469 ( .A(b[30]), .B(a[63]), .Z(n12850) );
  XOR U17470 ( .A(n12856), .B(n12857), .Z(n12484) );
  AND U17471 ( .A(n12858), .B(n12859), .Z(n12856) );
  AND U17472 ( .A(b[29]), .B(a[64]), .Z(n12855) );
  XOR U17473 ( .A(n12861), .B(n12862), .Z(n12489) );
  AND U17474 ( .A(n12863), .B(n12864), .Z(n12861) );
  AND U17475 ( .A(b[28]), .B(a[65]), .Z(n12860) );
  XOR U17476 ( .A(n12866), .B(n12867), .Z(n12494) );
  AND U17477 ( .A(n12868), .B(n12869), .Z(n12866) );
  AND U17478 ( .A(b[27]), .B(a[66]), .Z(n12865) );
  XOR U17479 ( .A(n12871), .B(n12872), .Z(n12499) );
  AND U17480 ( .A(n12873), .B(n12874), .Z(n12871) );
  AND U17481 ( .A(b[26]), .B(a[67]), .Z(n12870) );
  XOR U17482 ( .A(n12876), .B(n12877), .Z(n12504) );
  AND U17483 ( .A(n12878), .B(n12879), .Z(n12876) );
  AND U17484 ( .A(b[25]), .B(a[68]), .Z(n12875) );
  XOR U17485 ( .A(n12881), .B(n12882), .Z(n12509) );
  AND U17486 ( .A(n12883), .B(n12884), .Z(n12881) );
  AND U17487 ( .A(b[24]), .B(a[69]), .Z(n12880) );
  XOR U17488 ( .A(n12886), .B(n12887), .Z(n12514) );
  AND U17489 ( .A(n12888), .B(n12889), .Z(n12886) );
  AND U17490 ( .A(b[23]), .B(a[70]), .Z(n12885) );
  XOR U17491 ( .A(n12891), .B(n12892), .Z(n12519) );
  AND U17492 ( .A(n12893), .B(n12894), .Z(n12891) );
  AND U17493 ( .A(b[22]), .B(a[71]), .Z(n12890) );
  XOR U17494 ( .A(n12896), .B(n12897), .Z(n12524) );
  AND U17495 ( .A(n12898), .B(n12899), .Z(n12896) );
  AND U17496 ( .A(b[21]), .B(a[72]), .Z(n12895) );
  XOR U17497 ( .A(n12901), .B(n12902), .Z(n12529) );
  AND U17498 ( .A(n12903), .B(n12904), .Z(n12901) );
  AND U17499 ( .A(b[20]), .B(a[73]), .Z(n12900) );
  XOR U17500 ( .A(n12906), .B(n12907), .Z(n12534) );
  AND U17501 ( .A(n12908), .B(n12909), .Z(n12906) );
  AND U17502 ( .A(b[19]), .B(a[74]), .Z(n12905) );
  XOR U17503 ( .A(n12911), .B(n12912), .Z(n12539) );
  AND U17504 ( .A(n12913), .B(n12914), .Z(n12911) );
  AND U17505 ( .A(b[18]), .B(a[75]), .Z(n12910) );
  XOR U17506 ( .A(n12916), .B(n12917), .Z(n12544) );
  AND U17507 ( .A(n12918), .B(n12919), .Z(n12916) );
  AND U17508 ( .A(b[17]), .B(a[76]), .Z(n12915) );
  XOR U17509 ( .A(n12921), .B(n12922), .Z(n12549) );
  AND U17510 ( .A(n12923), .B(n12924), .Z(n12921) );
  AND U17511 ( .A(b[16]), .B(a[77]), .Z(n12920) );
  XOR U17512 ( .A(n12926), .B(n12927), .Z(n12554) );
  AND U17513 ( .A(n12928), .B(n12929), .Z(n12926) );
  AND U17514 ( .A(b[15]), .B(a[78]), .Z(n12925) );
  XOR U17515 ( .A(n12931), .B(n12932), .Z(n12559) );
  AND U17516 ( .A(n12933), .B(n12934), .Z(n12931) );
  AND U17517 ( .A(b[14]), .B(a[79]), .Z(n12930) );
  XOR U17518 ( .A(n12936), .B(n12937), .Z(n12564) );
  AND U17519 ( .A(n12938), .B(n12939), .Z(n12936) );
  AND U17520 ( .A(b[13]), .B(a[80]), .Z(n12935) );
  XOR U17521 ( .A(n12941), .B(n12942), .Z(n12569) );
  AND U17522 ( .A(n12943), .B(n12944), .Z(n12941) );
  AND U17523 ( .A(b[12]), .B(a[81]), .Z(n12940) );
  XOR U17524 ( .A(n12946), .B(n12947), .Z(n12574) );
  AND U17525 ( .A(n12948), .B(n12949), .Z(n12946) );
  AND U17526 ( .A(b[11]), .B(a[82]), .Z(n12945) );
  XOR U17527 ( .A(n12951), .B(n12952), .Z(n12579) );
  AND U17528 ( .A(n12953), .B(n12954), .Z(n12951) );
  AND U17529 ( .A(b[10]), .B(a[83]), .Z(n12950) );
  XOR U17530 ( .A(n12956), .B(n12957), .Z(n12584) );
  AND U17531 ( .A(n12958), .B(n12959), .Z(n12956) );
  AND U17532 ( .A(b[9]), .B(a[84]), .Z(n12955) );
  XOR U17533 ( .A(n12961), .B(n12962), .Z(n12589) );
  AND U17534 ( .A(n12963), .B(n12964), .Z(n12961) );
  AND U17535 ( .A(b[8]), .B(a[85]), .Z(n12960) );
  XOR U17536 ( .A(n12966), .B(n12967), .Z(n12594) );
  AND U17537 ( .A(n12968), .B(n12969), .Z(n12966) );
  AND U17538 ( .A(b[7]), .B(a[86]), .Z(n12965) );
  XOR U17539 ( .A(n12971), .B(n12972), .Z(n12599) );
  AND U17540 ( .A(n12973), .B(n12974), .Z(n12971) );
  AND U17541 ( .A(b[6]), .B(a[87]), .Z(n12970) );
  XOR U17542 ( .A(n12976), .B(n12977), .Z(n12604) );
  AND U17543 ( .A(n12978), .B(n12979), .Z(n12976) );
  AND U17544 ( .A(b[5]), .B(a[88]), .Z(n12975) );
  XOR U17545 ( .A(n12981), .B(n12982), .Z(n12609) );
  AND U17546 ( .A(n12983), .B(n12984), .Z(n12981) );
  AND U17547 ( .A(b[4]), .B(a[89]), .Z(n12980) );
  XOR U17548 ( .A(n12986), .B(n12987), .Z(n12614) );
  AND U17549 ( .A(n12988), .B(n12989), .Z(n12986) );
  AND U17550 ( .A(b[3]), .B(a[90]), .Z(n12985) );
  XOR U17551 ( .A(n12991), .B(n12992), .Z(n12619) );
  OR U17552 ( .A(n12993), .B(n12994), .Z(n12992) );
  AND U17553 ( .A(b[2]), .B(a[91]), .Z(n12990) );
  XNOR U17554 ( .A(n12629), .B(n12995), .Z(n12625) );
  NAND U17555 ( .A(b[1]), .B(a[92]), .Z(n12995) );
  IV U17556 ( .A(n12623), .Z(n12629) );
  ANDN U17557 ( .B(n10275), .A(n10277), .Z(n12623) );
  NAND U17558 ( .A(a[92]), .B(b[0]), .Z(n10277) );
  XOR U17559 ( .A(n12993), .B(n12994), .Z(n10275) );
  XOR U17560 ( .A(n12997), .B(n12988), .Z(n12996) );
  XOR U17561 ( .A(n12983), .B(n12987), .Z(n12998) );
  XOR U17562 ( .A(n12978), .B(n12982), .Z(n12999) );
  XOR U17563 ( .A(n12973), .B(n12977), .Z(n13000) );
  XOR U17564 ( .A(n12968), .B(n12972), .Z(n13001) );
  XOR U17565 ( .A(n12963), .B(n12967), .Z(n13002) );
  XOR U17566 ( .A(n12958), .B(n12962), .Z(n13003) );
  XOR U17567 ( .A(n12953), .B(n12957), .Z(n13004) );
  XOR U17568 ( .A(n12948), .B(n12952), .Z(n13005) );
  XOR U17569 ( .A(n12943), .B(n12947), .Z(n13006) );
  XOR U17570 ( .A(n12938), .B(n12942), .Z(n13007) );
  XOR U17571 ( .A(n12933), .B(n12937), .Z(n13008) );
  XOR U17572 ( .A(n12928), .B(n12932), .Z(n13009) );
  XOR U17573 ( .A(n12923), .B(n12927), .Z(n13010) );
  XOR U17574 ( .A(n12918), .B(n12922), .Z(n13011) );
  XOR U17575 ( .A(n12913), .B(n12917), .Z(n13012) );
  XOR U17576 ( .A(n12908), .B(n12912), .Z(n13013) );
  XOR U17577 ( .A(n12903), .B(n12907), .Z(n13014) );
  XOR U17578 ( .A(n12898), .B(n12902), .Z(n13015) );
  XOR U17579 ( .A(n12893), .B(n12897), .Z(n13016) );
  XOR U17580 ( .A(n12888), .B(n12892), .Z(n13017) );
  XOR U17581 ( .A(n12883), .B(n12887), .Z(n13018) );
  XOR U17582 ( .A(n12878), .B(n12882), .Z(n13019) );
  XOR U17583 ( .A(n12873), .B(n12877), .Z(n13020) );
  XOR U17584 ( .A(n12868), .B(n12872), .Z(n13021) );
  XOR U17585 ( .A(n12863), .B(n12867), .Z(n13022) );
  XOR U17586 ( .A(n12858), .B(n12862), .Z(n13023) );
  XOR U17587 ( .A(n12853), .B(n12857), .Z(n13024) );
  XOR U17588 ( .A(n12848), .B(n12852), .Z(n13025) );
  XOR U17589 ( .A(n12843), .B(n12847), .Z(n13026) );
  XOR U17590 ( .A(n12838), .B(n12842), .Z(n13027) );
  XOR U17591 ( .A(n12833), .B(n12837), .Z(n13028) );
  XOR U17592 ( .A(n12828), .B(n12832), .Z(n13029) );
  XOR U17593 ( .A(n12823), .B(n12827), .Z(n13030) );
  XOR U17594 ( .A(n12818), .B(n12822), .Z(n13031) );
  XOR U17595 ( .A(n12813), .B(n12817), .Z(n13032) );
  XOR U17596 ( .A(n12808), .B(n12812), .Z(n13033) );
  XOR U17597 ( .A(n12803), .B(n12807), .Z(n13034) );
  XOR U17598 ( .A(n12798), .B(n12802), .Z(n13035) );
  XOR U17599 ( .A(n12793), .B(n12797), .Z(n13036) );
  XOR U17600 ( .A(n12788), .B(n12792), .Z(n13037) );
  XOR U17601 ( .A(n12783), .B(n12787), .Z(n13038) );
  XOR U17602 ( .A(n12778), .B(n12782), .Z(n13039) );
  XOR U17603 ( .A(n12773), .B(n12777), .Z(n13040) );
  XOR U17604 ( .A(n12768), .B(n12772), .Z(n13041) );
  XOR U17605 ( .A(n12763), .B(n12767), .Z(n13042) );
  XOR U17606 ( .A(n12758), .B(n12762), .Z(n13043) );
  XOR U17607 ( .A(n12753), .B(n12757), .Z(n13044) );
  XOR U17608 ( .A(n12748), .B(n12752), .Z(n13045) );
  XOR U17609 ( .A(n12743), .B(n12747), .Z(n13046) );
  XOR U17610 ( .A(n12738), .B(n12742), .Z(n13047) );
  XOR U17611 ( .A(n12733), .B(n12737), .Z(n13048) );
  XOR U17612 ( .A(n12728), .B(n12732), .Z(n13049) );
  XOR U17613 ( .A(n12723), .B(n12727), .Z(n13050) );
  XOR U17614 ( .A(n12713), .B(n12722), .Z(n13051) );
  XOR U17615 ( .A(n13052), .B(n12712), .Z(n12713) );
  AND U17616 ( .A(a[36]), .B(b[56]), .Z(n13052) );
  XNOR U17617 ( .A(n12712), .B(n12718), .Z(n13053) );
  XNOR U17618 ( .A(n12717), .B(n12709), .Z(n13054) );
  XNOR U17619 ( .A(n12708), .B(n12704), .Z(n13055) );
  XOR U17620 ( .A(n12703), .B(n12700), .Z(n13056) );
  XOR U17621 ( .A(n13057), .B(n13058), .Z(n12700) );
  XOR U17622 ( .A(n12698), .B(n13059), .Z(n13058) );
  XOR U17623 ( .A(n13060), .B(n13061), .Z(n13059) );
  XOR U17624 ( .A(n13062), .B(n13063), .Z(n13061) );
  NAND U17625 ( .A(a[30]), .B(b[62]), .Z(n13063) );
  AND U17626 ( .A(a[29]), .B(b[63]), .Z(n13062) );
  XOR U17627 ( .A(n13064), .B(n13060), .Z(n13057) );
  XOR U17628 ( .A(n13065), .B(n13066), .Z(n13060) );
  ANDN U17629 ( .B(n13067), .A(n13068), .Z(n13065) );
  AND U17630 ( .A(a[31]), .B(b[61]), .Z(n13064) );
  XOR U17631 ( .A(n13069), .B(n12698), .Z(n12699) );
  XOR U17632 ( .A(n13070), .B(n13071), .Z(n12698) );
  AND U17633 ( .A(n13072), .B(n13073), .Z(n13070) );
  AND U17634 ( .A(a[32]), .B(b[60]), .Z(n13069) );
  XOR U17635 ( .A(n13074), .B(n12703), .Z(n12705) );
  XOR U17636 ( .A(n13075), .B(n13076), .Z(n12703) );
  AND U17637 ( .A(n13077), .B(n13078), .Z(n13075) );
  AND U17638 ( .A(a[33]), .B(b[59]), .Z(n13074) );
  XOR U17639 ( .A(n13079), .B(n12708), .Z(n12710) );
  XOR U17640 ( .A(n13080), .B(n13081), .Z(n12708) );
  AND U17641 ( .A(n13082), .B(n13083), .Z(n13080) );
  AND U17642 ( .A(a[34]), .B(b[58]), .Z(n13079) );
  XOR U17643 ( .A(n13084), .B(n13085), .Z(n12712) );
  AND U17644 ( .A(n13086), .B(n13087), .Z(n13084) );
  XOR U17645 ( .A(n13088), .B(n12717), .Z(n12719) );
  XOR U17646 ( .A(n13089), .B(n13090), .Z(n12717) );
  AND U17647 ( .A(n13091), .B(n13092), .Z(n13089) );
  AND U17648 ( .A(a[35]), .B(b[57]), .Z(n13088) );
  XOR U17649 ( .A(n13094), .B(n13095), .Z(n12722) );
  AND U17650 ( .A(n13096), .B(n13097), .Z(n13094) );
  AND U17651 ( .A(a[37]), .B(b[55]), .Z(n13093) );
  XOR U17652 ( .A(n13099), .B(n13100), .Z(n12727) );
  AND U17653 ( .A(n13101), .B(n13102), .Z(n13099) );
  AND U17654 ( .A(a[38]), .B(b[54]), .Z(n13098) );
  XOR U17655 ( .A(n13104), .B(n13105), .Z(n12732) );
  AND U17656 ( .A(n13106), .B(n13107), .Z(n13104) );
  AND U17657 ( .A(a[39]), .B(b[53]), .Z(n13103) );
  XOR U17658 ( .A(n13109), .B(n13110), .Z(n12737) );
  AND U17659 ( .A(n13111), .B(n13112), .Z(n13109) );
  AND U17660 ( .A(a[40]), .B(b[52]), .Z(n13108) );
  XOR U17661 ( .A(n13114), .B(n13115), .Z(n12742) );
  AND U17662 ( .A(n13116), .B(n13117), .Z(n13114) );
  AND U17663 ( .A(a[41]), .B(b[51]), .Z(n13113) );
  XOR U17664 ( .A(n13119), .B(n13120), .Z(n12747) );
  AND U17665 ( .A(n13121), .B(n13122), .Z(n13119) );
  AND U17666 ( .A(a[42]), .B(b[50]), .Z(n13118) );
  XOR U17667 ( .A(n13124), .B(n13125), .Z(n12752) );
  AND U17668 ( .A(n13126), .B(n13127), .Z(n13124) );
  AND U17669 ( .A(a[43]), .B(b[49]), .Z(n13123) );
  XOR U17670 ( .A(n13129), .B(n13130), .Z(n12757) );
  AND U17671 ( .A(n13131), .B(n13132), .Z(n13129) );
  AND U17672 ( .A(a[44]), .B(b[48]), .Z(n13128) );
  XOR U17673 ( .A(n13134), .B(n13135), .Z(n12762) );
  AND U17674 ( .A(n13136), .B(n13137), .Z(n13134) );
  AND U17675 ( .A(a[45]), .B(b[47]), .Z(n13133) );
  XOR U17676 ( .A(n13139), .B(n13140), .Z(n12767) );
  AND U17677 ( .A(n13141), .B(n13142), .Z(n13139) );
  AND U17678 ( .A(a[46]), .B(b[46]), .Z(n13138) );
  XOR U17679 ( .A(n13144), .B(n13145), .Z(n12772) );
  AND U17680 ( .A(n13146), .B(n13147), .Z(n13144) );
  AND U17681 ( .A(b[45]), .B(a[47]), .Z(n13143) );
  XOR U17682 ( .A(n13149), .B(n13150), .Z(n12777) );
  AND U17683 ( .A(n13151), .B(n13152), .Z(n13149) );
  AND U17684 ( .A(b[44]), .B(a[48]), .Z(n13148) );
  XOR U17685 ( .A(n13154), .B(n13155), .Z(n12782) );
  AND U17686 ( .A(n13156), .B(n13157), .Z(n13154) );
  AND U17687 ( .A(b[43]), .B(a[49]), .Z(n13153) );
  XOR U17688 ( .A(n13159), .B(n13160), .Z(n12787) );
  AND U17689 ( .A(n13161), .B(n13162), .Z(n13159) );
  AND U17690 ( .A(b[42]), .B(a[50]), .Z(n13158) );
  XOR U17691 ( .A(n13164), .B(n13165), .Z(n12792) );
  AND U17692 ( .A(n13166), .B(n13167), .Z(n13164) );
  AND U17693 ( .A(b[41]), .B(a[51]), .Z(n13163) );
  XOR U17694 ( .A(n13169), .B(n13170), .Z(n12797) );
  AND U17695 ( .A(n13171), .B(n13172), .Z(n13169) );
  AND U17696 ( .A(b[40]), .B(a[52]), .Z(n13168) );
  XOR U17697 ( .A(n13174), .B(n13175), .Z(n12802) );
  AND U17698 ( .A(n13176), .B(n13177), .Z(n13174) );
  AND U17699 ( .A(b[39]), .B(a[53]), .Z(n13173) );
  XOR U17700 ( .A(n13179), .B(n13180), .Z(n12807) );
  AND U17701 ( .A(n13181), .B(n13182), .Z(n13179) );
  AND U17702 ( .A(b[38]), .B(a[54]), .Z(n13178) );
  XOR U17703 ( .A(n13184), .B(n13185), .Z(n12812) );
  AND U17704 ( .A(n13186), .B(n13187), .Z(n13184) );
  AND U17705 ( .A(b[37]), .B(a[55]), .Z(n13183) );
  XOR U17706 ( .A(n13189), .B(n13190), .Z(n12817) );
  AND U17707 ( .A(n13191), .B(n13192), .Z(n13189) );
  AND U17708 ( .A(b[36]), .B(a[56]), .Z(n13188) );
  XOR U17709 ( .A(n13194), .B(n13195), .Z(n12822) );
  AND U17710 ( .A(n13196), .B(n13197), .Z(n13194) );
  AND U17711 ( .A(b[35]), .B(a[57]), .Z(n13193) );
  XOR U17712 ( .A(n13199), .B(n13200), .Z(n12827) );
  AND U17713 ( .A(n13201), .B(n13202), .Z(n13199) );
  AND U17714 ( .A(b[34]), .B(a[58]), .Z(n13198) );
  XOR U17715 ( .A(n13204), .B(n13205), .Z(n12832) );
  AND U17716 ( .A(n13206), .B(n13207), .Z(n13204) );
  AND U17717 ( .A(b[33]), .B(a[59]), .Z(n13203) );
  XOR U17718 ( .A(n13209), .B(n13210), .Z(n12837) );
  AND U17719 ( .A(n13211), .B(n13212), .Z(n13209) );
  AND U17720 ( .A(b[32]), .B(a[60]), .Z(n13208) );
  XOR U17721 ( .A(n13214), .B(n13215), .Z(n12842) );
  AND U17722 ( .A(n13216), .B(n13217), .Z(n13214) );
  AND U17723 ( .A(b[31]), .B(a[61]), .Z(n13213) );
  XOR U17724 ( .A(n13219), .B(n13220), .Z(n12847) );
  AND U17725 ( .A(n13221), .B(n13222), .Z(n13219) );
  AND U17726 ( .A(b[30]), .B(a[62]), .Z(n13218) );
  XOR U17727 ( .A(n13224), .B(n13225), .Z(n12852) );
  AND U17728 ( .A(n13226), .B(n13227), .Z(n13224) );
  AND U17729 ( .A(b[29]), .B(a[63]), .Z(n13223) );
  XOR U17730 ( .A(n13229), .B(n13230), .Z(n12857) );
  AND U17731 ( .A(n13231), .B(n13232), .Z(n13229) );
  AND U17732 ( .A(b[28]), .B(a[64]), .Z(n13228) );
  XOR U17733 ( .A(n13234), .B(n13235), .Z(n12862) );
  AND U17734 ( .A(n13236), .B(n13237), .Z(n13234) );
  AND U17735 ( .A(b[27]), .B(a[65]), .Z(n13233) );
  XOR U17736 ( .A(n13239), .B(n13240), .Z(n12867) );
  AND U17737 ( .A(n13241), .B(n13242), .Z(n13239) );
  AND U17738 ( .A(b[26]), .B(a[66]), .Z(n13238) );
  XOR U17739 ( .A(n13244), .B(n13245), .Z(n12872) );
  AND U17740 ( .A(n13246), .B(n13247), .Z(n13244) );
  AND U17741 ( .A(b[25]), .B(a[67]), .Z(n13243) );
  XOR U17742 ( .A(n13249), .B(n13250), .Z(n12877) );
  AND U17743 ( .A(n13251), .B(n13252), .Z(n13249) );
  AND U17744 ( .A(b[24]), .B(a[68]), .Z(n13248) );
  XOR U17745 ( .A(n13254), .B(n13255), .Z(n12882) );
  AND U17746 ( .A(n13256), .B(n13257), .Z(n13254) );
  AND U17747 ( .A(b[23]), .B(a[69]), .Z(n13253) );
  XOR U17748 ( .A(n13259), .B(n13260), .Z(n12887) );
  AND U17749 ( .A(n13261), .B(n13262), .Z(n13259) );
  AND U17750 ( .A(b[22]), .B(a[70]), .Z(n13258) );
  XOR U17751 ( .A(n13264), .B(n13265), .Z(n12892) );
  AND U17752 ( .A(n13266), .B(n13267), .Z(n13264) );
  AND U17753 ( .A(b[21]), .B(a[71]), .Z(n13263) );
  XOR U17754 ( .A(n13269), .B(n13270), .Z(n12897) );
  AND U17755 ( .A(n13271), .B(n13272), .Z(n13269) );
  AND U17756 ( .A(b[20]), .B(a[72]), .Z(n13268) );
  XOR U17757 ( .A(n13274), .B(n13275), .Z(n12902) );
  AND U17758 ( .A(n13276), .B(n13277), .Z(n13274) );
  AND U17759 ( .A(b[19]), .B(a[73]), .Z(n13273) );
  XOR U17760 ( .A(n13279), .B(n13280), .Z(n12907) );
  AND U17761 ( .A(n13281), .B(n13282), .Z(n13279) );
  AND U17762 ( .A(b[18]), .B(a[74]), .Z(n13278) );
  XOR U17763 ( .A(n13284), .B(n13285), .Z(n12912) );
  AND U17764 ( .A(n13286), .B(n13287), .Z(n13284) );
  AND U17765 ( .A(b[17]), .B(a[75]), .Z(n13283) );
  XOR U17766 ( .A(n13289), .B(n13290), .Z(n12917) );
  AND U17767 ( .A(n13291), .B(n13292), .Z(n13289) );
  AND U17768 ( .A(b[16]), .B(a[76]), .Z(n13288) );
  XOR U17769 ( .A(n13294), .B(n13295), .Z(n12922) );
  AND U17770 ( .A(n13296), .B(n13297), .Z(n13294) );
  AND U17771 ( .A(b[15]), .B(a[77]), .Z(n13293) );
  XOR U17772 ( .A(n13299), .B(n13300), .Z(n12927) );
  AND U17773 ( .A(n13301), .B(n13302), .Z(n13299) );
  AND U17774 ( .A(b[14]), .B(a[78]), .Z(n13298) );
  XOR U17775 ( .A(n13304), .B(n13305), .Z(n12932) );
  AND U17776 ( .A(n13306), .B(n13307), .Z(n13304) );
  AND U17777 ( .A(b[13]), .B(a[79]), .Z(n13303) );
  XOR U17778 ( .A(n13309), .B(n13310), .Z(n12937) );
  AND U17779 ( .A(n13311), .B(n13312), .Z(n13309) );
  AND U17780 ( .A(b[12]), .B(a[80]), .Z(n13308) );
  XOR U17781 ( .A(n13314), .B(n13315), .Z(n12942) );
  AND U17782 ( .A(n13316), .B(n13317), .Z(n13314) );
  AND U17783 ( .A(b[11]), .B(a[81]), .Z(n13313) );
  XOR U17784 ( .A(n13319), .B(n13320), .Z(n12947) );
  AND U17785 ( .A(n13321), .B(n13322), .Z(n13319) );
  AND U17786 ( .A(b[10]), .B(a[82]), .Z(n13318) );
  XOR U17787 ( .A(n13324), .B(n13325), .Z(n12952) );
  AND U17788 ( .A(n13326), .B(n13327), .Z(n13324) );
  AND U17789 ( .A(b[9]), .B(a[83]), .Z(n13323) );
  XOR U17790 ( .A(n13329), .B(n13330), .Z(n12957) );
  AND U17791 ( .A(n13331), .B(n13332), .Z(n13329) );
  AND U17792 ( .A(b[8]), .B(a[84]), .Z(n13328) );
  XOR U17793 ( .A(n13334), .B(n13335), .Z(n12962) );
  AND U17794 ( .A(n13336), .B(n13337), .Z(n13334) );
  AND U17795 ( .A(b[7]), .B(a[85]), .Z(n13333) );
  XOR U17796 ( .A(n13339), .B(n13340), .Z(n12967) );
  AND U17797 ( .A(n13341), .B(n13342), .Z(n13339) );
  AND U17798 ( .A(b[6]), .B(a[86]), .Z(n13338) );
  XOR U17799 ( .A(n13344), .B(n13345), .Z(n12972) );
  AND U17800 ( .A(n13346), .B(n13347), .Z(n13344) );
  AND U17801 ( .A(b[5]), .B(a[87]), .Z(n13343) );
  XOR U17802 ( .A(n13349), .B(n13350), .Z(n12977) );
  AND U17803 ( .A(n13351), .B(n13352), .Z(n13349) );
  AND U17804 ( .A(b[4]), .B(a[88]), .Z(n13348) );
  XOR U17805 ( .A(n13354), .B(n13355), .Z(n12982) );
  AND U17806 ( .A(n13356), .B(n13357), .Z(n13354) );
  AND U17807 ( .A(b[3]), .B(a[89]), .Z(n13353) );
  XOR U17808 ( .A(n13359), .B(n13360), .Z(n12987) );
  OR U17809 ( .A(n13361), .B(n13362), .Z(n13360) );
  AND U17810 ( .A(b[2]), .B(a[90]), .Z(n13358) );
  XNOR U17811 ( .A(n12997), .B(n13363), .Z(n12993) );
  NAND U17812 ( .A(b[1]), .B(a[91]), .Z(n13363) );
  IV U17813 ( .A(n12991), .Z(n12997) );
  ANDN U17814 ( .B(n10278), .A(n10280), .Z(n12991) );
  NAND U17815 ( .A(a[91]), .B(b[0]), .Z(n10280) );
  XOR U17816 ( .A(n13361), .B(n13362), .Z(n10278) );
  XOR U17817 ( .A(n13365), .B(n13356), .Z(n13364) );
  XOR U17818 ( .A(n13351), .B(n13355), .Z(n13366) );
  XOR U17819 ( .A(n13346), .B(n13350), .Z(n13367) );
  XOR U17820 ( .A(n13341), .B(n13345), .Z(n13368) );
  XOR U17821 ( .A(n13336), .B(n13340), .Z(n13369) );
  XOR U17822 ( .A(n13331), .B(n13335), .Z(n13370) );
  XOR U17823 ( .A(n13326), .B(n13330), .Z(n13371) );
  XOR U17824 ( .A(n13321), .B(n13325), .Z(n13372) );
  XOR U17825 ( .A(n13316), .B(n13320), .Z(n13373) );
  XOR U17826 ( .A(n13311), .B(n13315), .Z(n13374) );
  XOR U17827 ( .A(n13306), .B(n13310), .Z(n13375) );
  XOR U17828 ( .A(n13301), .B(n13305), .Z(n13376) );
  XOR U17829 ( .A(n13296), .B(n13300), .Z(n13377) );
  XOR U17830 ( .A(n13291), .B(n13295), .Z(n13378) );
  XOR U17831 ( .A(n13286), .B(n13290), .Z(n13379) );
  XOR U17832 ( .A(n13281), .B(n13285), .Z(n13380) );
  XOR U17833 ( .A(n13276), .B(n13280), .Z(n13381) );
  XOR U17834 ( .A(n13271), .B(n13275), .Z(n13382) );
  XOR U17835 ( .A(n13266), .B(n13270), .Z(n13383) );
  XOR U17836 ( .A(n13261), .B(n13265), .Z(n13384) );
  XOR U17837 ( .A(n13256), .B(n13260), .Z(n13385) );
  XOR U17838 ( .A(n13251), .B(n13255), .Z(n13386) );
  XOR U17839 ( .A(n13246), .B(n13250), .Z(n13387) );
  XOR U17840 ( .A(n13241), .B(n13245), .Z(n13388) );
  XOR U17841 ( .A(n13236), .B(n13240), .Z(n13389) );
  XOR U17842 ( .A(n13231), .B(n13235), .Z(n13390) );
  XOR U17843 ( .A(n13226), .B(n13230), .Z(n13391) );
  XOR U17844 ( .A(n13221), .B(n13225), .Z(n13392) );
  XOR U17845 ( .A(n13216), .B(n13220), .Z(n13393) );
  XOR U17846 ( .A(n13211), .B(n13215), .Z(n13394) );
  XOR U17847 ( .A(n13206), .B(n13210), .Z(n13395) );
  XOR U17848 ( .A(n13201), .B(n13205), .Z(n13396) );
  XOR U17849 ( .A(n13196), .B(n13200), .Z(n13397) );
  XOR U17850 ( .A(n13191), .B(n13195), .Z(n13398) );
  XOR U17851 ( .A(n13186), .B(n13190), .Z(n13399) );
  XOR U17852 ( .A(n13181), .B(n13185), .Z(n13400) );
  XOR U17853 ( .A(n13176), .B(n13180), .Z(n13401) );
  XOR U17854 ( .A(n13171), .B(n13175), .Z(n13402) );
  XOR U17855 ( .A(n13166), .B(n13170), .Z(n13403) );
  XOR U17856 ( .A(n13161), .B(n13165), .Z(n13404) );
  XOR U17857 ( .A(n13156), .B(n13160), .Z(n13405) );
  XOR U17858 ( .A(n13151), .B(n13155), .Z(n13406) );
  XOR U17859 ( .A(n13146), .B(n13150), .Z(n13407) );
  XOR U17860 ( .A(n13141), .B(n13145), .Z(n13408) );
  XOR U17861 ( .A(n13136), .B(n13140), .Z(n13409) );
  XOR U17862 ( .A(n13131), .B(n13135), .Z(n13410) );
  XOR U17863 ( .A(n13126), .B(n13130), .Z(n13411) );
  XOR U17864 ( .A(n13121), .B(n13125), .Z(n13412) );
  XOR U17865 ( .A(n13116), .B(n13120), .Z(n13413) );
  XOR U17866 ( .A(n13111), .B(n13115), .Z(n13414) );
  XOR U17867 ( .A(n13106), .B(n13110), .Z(n13415) );
  XOR U17868 ( .A(n13101), .B(n13105), .Z(n13416) );
  XOR U17869 ( .A(n13096), .B(n13100), .Z(n13417) );
  XOR U17870 ( .A(n13086), .B(n13095), .Z(n13418) );
  XOR U17871 ( .A(n13419), .B(n13085), .Z(n13086) );
  AND U17872 ( .A(a[36]), .B(b[55]), .Z(n13419) );
  XNOR U17873 ( .A(n13085), .B(n13091), .Z(n13420) );
  XNOR U17874 ( .A(n13090), .B(n13082), .Z(n13421) );
  XNOR U17875 ( .A(n13081), .B(n13077), .Z(n13422) );
  XNOR U17876 ( .A(n13076), .B(n13072), .Z(n13423) );
  XOR U17877 ( .A(n13071), .B(n13068), .Z(n13424) );
  XOR U17878 ( .A(n13425), .B(n13426), .Z(n13068) );
  XOR U17879 ( .A(n13066), .B(n13427), .Z(n13426) );
  XOR U17880 ( .A(n13428), .B(n13429), .Z(n13427) );
  XOR U17881 ( .A(n13430), .B(n13431), .Z(n13429) );
  NAND U17882 ( .A(a[29]), .B(b[62]), .Z(n13431) );
  AND U17883 ( .A(a[28]), .B(b[63]), .Z(n13430) );
  XOR U17884 ( .A(n13432), .B(n13428), .Z(n13425) );
  XOR U17885 ( .A(n13433), .B(n13434), .Z(n13428) );
  ANDN U17886 ( .B(n13435), .A(n13436), .Z(n13433) );
  AND U17887 ( .A(a[30]), .B(b[61]), .Z(n13432) );
  XOR U17888 ( .A(n13437), .B(n13066), .Z(n13067) );
  XOR U17889 ( .A(n13438), .B(n13439), .Z(n13066) );
  AND U17890 ( .A(n13440), .B(n13441), .Z(n13438) );
  AND U17891 ( .A(a[31]), .B(b[60]), .Z(n13437) );
  XOR U17892 ( .A(n13442), .B(n13071), .Z(n13073) );
  XOR U17893 ( .A(n13443), .B(n13444), .Z(n13071) );
  AND U17894 ( .A(n13445), .B(n13446), .Z(n13443) );
  AND U17895 ( .A(a[32]), .B(b[59]), .Z(n13442) );
  XOR U17896 ( .A(n13447), .B(n13076), .Z(n13078) );
  XOR U17897 ( .A(n13448), .B(n13449), .Z(n13076) );
  AND U17898 ( .A(n13450), .B(n13451), .Z(n13448) );
  AND U17899 ( .A(a[33]), .B(b[58]), .Z(n13447) );
  XOR U17900 ( .A(n13452), .B(n13081), .Z(n13083) );
  XOR U17901 ( .A(n13453), .B(n13454), .Z(n13081) );
  AND U17902 ( .A(n13455), .B(n13456), .Z(n13453) );
  AND U17903 ( .A(a[34]), .B(b[57]), .Z(n13452) );
  XOR U17904 ( .A(n13457), .B(n13458), .Z(n13085) );
  AND U17905 ( .A(n13459), .B(n13460), .Z(n13457) );
  XOR U17906 ( .A(n13461), .B(n13090), .Z(n13092) );
  XOR U17907 ( .A(n13462), .B(n13463), .Z(n13090) );
  AND U17908 ( .A(n13464), .B(n13465), .Z(n13462) );
  AND U17909 ( .A(a[35]), .B(b[56]), .Z(n13461) );
  XOR U17910 ( .A(n13467), .B(n13468), .Z(n13095) );
  AND U17911 ( .A(n13469), .B(n13470), .Z(n13467) );
  AND U17912 ( .A(a[37]), .B(b[54]), .Z(n13466) );
  XOR U17913 ( .A(n13472), .B(n13473), .Z(n13100) );
  AND U17914 ( .A(n13474), .B(n13475), .Z(n13472) );
  AND U17915 ( .A(a[38]), .B(b[53]), .Z(n13471) );
  XOR U17916 ( .A(n13477), .B(n13478), .Z(n13105) );
  AND U17917 ( .A(n13479), .B(n13480), .Z(n13477) );
  AND U17918 ( .A(a[39]), .B(b[52]), .Z(n13476) );
  XOR U17919 ( .A(n13482), .B(n13483), .Z(n13110) );
  AND U17920 ( .A(n13484), .B(n13485), .Z(n13482) );
  AND U17921 ( .A(a[40]), .B(b[51]), .Z(n13481) );
  XOR U17922 ( .A(n13487), .B(n13488), .Z(n13115) );
  AND U17923 ( .A(n13489), .B(n13490), .Z(n13487) );
  AND U17924 ( .A(a[41]), .B(b[50]), .Z(n13486) );
  XOR U17925 ( .A(n13492), .B(n13493), .Z(n13120) );
  AND U17926 ( .A(n13494), .B(n13495), .Z(n13492) );
  AND U17927 ( .A(a[42]), .B(b[49]), .Z(n13491) );
  XOR U17928 ( .A(n13497), .B(n13498), .Z(n13125) );
  AND U17929 ( .A(n13499), .B(n13500), .Z(n13497) );
  AND U17930 ( .A(a[43]), .B(b[48]), .Z(n13496) );
  XOR U17931 ( .A(n13502), .B(n13503), .Z(n13130) );
  AND U17932 ( .A(n13504), .B(n13505), .Z(n13502) );
  AND U17933 ( .A(a[44]), .B(b[47]), .Z(n13501) );
  XOR U17934 ( .A(n13507), .B(n13508), .Z(n13135) );
  AND U17935 ( .A(n13509), .B(n13510), .Z(n13507) );
  AND U17936 ( .A(a[45]), .B(b[46]), .Z(n13506) );
  XOR U17937 ( .A(n13512), .B(n13513), .Z(n13140) );
  AND U17938 ( .A(n13514), .B(n13515), .Z(n13512) );
  AND U17939 ( .A(b[45]), .B(a[46]), .Z(n13511) );
  XOR U17940 ( .A(n13517), .B(n13518), .Z(n13145) );
  AND U17941 ( .A(n13519), .B(n13520), .Z(n13517) );
  AND U17942 ( .A(b[44]), .B(a[47]), .Z(n13516) );
  XOR U17943 ( .A(n13522), .B(n13523), .Z(n13150) );
  AND U17944 ( .A(n13524), .B(n13525), .Z(n13522) );
  AND U17945 ( .A(b[43]), .B(a[48]), .Z(n13521) );
  XOR U17946 ( .A(n13527), .B(n13528), .Z(n13155) );
  AND U17947 ( .A(n13529), .B(n13530), .Z(n13527) );
  AND U17948 ( .A(b[42]), .B(a[49]), .Z(n13526) );
  XOR U17949 ( .A(n13532), .B(n13533), .Z(n13160) );
  AND U17950 ( .A(n13534), .B(n13535), .Z(n13532) );
  AND U17951 ( .A(b[41]), .B(a[50]), .Z(n13531) );
  XOR U17952 ( .A(n13537), .B(n13538), .Z(n13165) );
  AND U17953 ( .A(n13539), .B(n13540), .Z(n13537) );
  AND U17954 ( .A(b[40]), .B(a[51]), .Z(n13536) );
  XOR U17955 ( .A(n13542), .B(n13543), .Z(n13170) );
  AND U17956 ( .A(n13544), .B(n13545), .Z(n13542) );
  AND U17957 ( .A(b[39]), .B(a[52]), .Z(n13541) );
  XOR U17958 ( .A(n13547), .B(n13548), .Z(n13175) );
  AND U17959 ( .A(n13549), .B(n13550), .Z(n13547) );
  AND U17960 ( .A(b[38]), .B(a[53]), .Z(n13546) );
  XOR U17961 ( .A(n13552), .B(n13553), .Z(n13180) );
  AND U17962 ( .A(n13554), .B(n13555), .Z(n13552) );
  AND U17963 ( .A(b[37]), .B(a[54]), .Z(n13551) );
  XOR U17964 ( .A(n13557), .B(n13558), .Z(n13185) );
  AND U17965 ( .A(n13559), .B(n13560), .Z(n13557) );
  AND U17966 ( .A(b[36]), .B(a[55]), .Z(n13556) );
  XOR U17967 ( .A(n13562), .B(n13563), .Z(n13190) );
  AND U17968 ( .A(n13564), .B(n13565), .Z(n13562) );
  AND U17969 ( .A(b[35]), .B(a[56]), .Z(n13561) );
  XOR U17970 ( .A(n13567), .B(n13568), .Z(n13195) );
  AND U17971 ( .A(n13569), .B(n13570), .Z(n13567) );
  AND U17972 ( .A(b[34]), .B(a[57]), .Z(n13566) );
  XOR U17973 ( .A(n13572), .B(n13573), .Z(n13200) );
  AND U17974 ( .A(n13574), .B(n13575), .Z(n13572) );
  AND U17975 ( .A(b[33]), .B(a[58]), .Z(n13571) );
  XOR U17976 ( .A(n13577), .B(n13578), .Z(n13205) );
  AND U17977 ( .A(n13579), .B(n13580), .Z(n13577) );
  AND U17978 ( .A(b[32]), .B(a[59]), .Z(n13576) );
  XOR U17979 ( .A(n13582), .B(n13583), .Z(n13210) );
  AND U17980 ( .A(n13584), .B(n13585), .Z(n13582) );
  AND U17981 ( .A(b[31]), .B(a[60]), .Z(n13581) );
  XOR U17982 ( .A(n13587), .B(n13588), .Z(n13215) );
  AND U17983 ( .A(n13589), .B(n13590), .Z(n13587) );
  AND U17984 ( .A(b[30]), .B(a[61]), .Z(n13586) );
  XOR U17985 ( .A(n13592), .B(n13593), .Z(n13220) );
  AND U17986 ( .A(n13594), .B(n13595), .Z(n13592) );
  AND U17987 ( .A(b[29]), .B(a[62]), .Z(n13591) );
  XOR U17988 ( .A(n13597), .B(n13598), .Z(n13225) );
  AND U17989 ( .A(n13599), .B(n13600), .Z(n13597) );
  AND U17990 ( .A(b[28]), .B(a[63]), .Z(n13596) );
  XOR U17991 ( .A(n13602), .B(n13603), .Z(n13230) );
  AND U17992 ( .A(n13604), .B(n13605), .Z(n13602) );
  AND U17993 ( .A(b[27]), .B(a[64]), .Z(n13601) );
  XOR U17994 ( .A(n13607), .B(n13608), .Z(n13235) );
  AND U17995 ( .A(n13609), .B(n13610), .Z(n13607) );
  AND U17996 ( .A(b[26]), .B(a[65]), .Z(n13606) );
  XOR U17997 ( .A(n13612), .B(n13613), .Z(n13240) );
  AND U17998 ( .A(n13614), .B(n13615), .Z(n13612) );
  AND U17999 ( .A(b[25]), .B(a[66]), .Z(n13611) );
  XOR U18000 ( .A(n13617), .B(n13618), .Z(n13245) );
  AND U18001 ( .A(n13619), .B(n13620), .Z(n13617) );
  AND U18002 ( .A(b[24]), .B(a[67]), .Z(n13616) );
  XOR U18003 ( .A(n13622), .B(n13623), .Z(n13250) );
  AND U18004 ( .A(n13624), .B(n13625), .Z(n13622) );
  AND U18005 ( .A(b[23]), .B(a[68]), .Z(n13621) );
  XOR U18006 ( .A(n13627), .B(n13628), .Z(n13255) );
  AND U18007 ( .A(n13629), .B(n13630), .Z(n13627) );
  AND U18008 ( .A(b[22]), .B(a[69]), .Z(n13626) );
  XOR U18009 ( .A(n13632), .B(n13633), .Z(n13260) );
  AND U18010 ( .A(n13634), .B(n13635), .Z(n13632) );
  AND U18011 ( .A(b[21]), .B(a[70]), .Z(n13631) );
  XOR U18012 ( .A(n13637), .B(n13638), .Z(n13265) );
  AND U18013 ( .A(n13639), .B(n13640), .Z(n13637) );
  AND U18014 ( .A(b[20]), .B(a[71]), .Z(n13636) );
  XOR U18015 ( .A(n13642), .B(n13643), .Z(n13270) );
  AND U18016 ( .A(n13644), .B(n13645), .Z(n13642) );
  AND U18017 ( .A(b[19]), .B(a[72]), .Z(n13641) );
  XOR U18018 ( .A(n13647), .B(n13648), .Z(n13275) );
  AND U18019 ( .A(n13649), .B(n13650), .Z(n13647) );
  AND U18020 ( .A(b[18]), .B(a[73]), .Z(n13646) );
  XOR U18021 ( .A(n13652), .B(n13653), .Z(n13280) );
  AND U18022 ( .A(n13654), .B(n13655), .Z(n13652) );
  AND U18023 ( .A(b[17]), .B(a[74]), .Z(n13651) );
  XOR U18024 ( .A(n13657), .B(n13658), .Z(n13285) );
  AND U18025 ( .A(n13659), .B(n13660), .Z(n13657) );
  AND U18026 ( .A(b[16]), .B(a[75]), .Z(n13656) );
  XOR U18027 ( .A(n13662), .B(n13663), .Z(n13290) );
  AND U18028 ( .A(n13664), .B(n13665), .Z(n13662) );
  AND U18029 ( .A(b[15]), .B(a[76]), .Z(n13661) );
  XOR U18030 ( .A(n13667), .B(n13668), .Z(n13295) );
  AND U18031 ( .A(n13669), .B(n13670), .Z(n13667) );
  AND U18032 ( .A(b[14]), .B(a[77]), .Z(n13666) );
  XOR U18033 ( .A(n13672), .B(n13673), .Z(n13300) );
  AND U18034 ( .A(n13674), .B(n13675), .Z(n13672) );
  AND U18035 ( .A(b[13]), .B(a[78]), .Z(n13671) );
  XOR U18036 ( .A(n13677), .B(n13678), .Z(n13305) );
  AND U18037 ( .A(n13679), .B(n13680), .Z(n13677) );
  AND U18038 ( .A(b[12]), .B(a[79]), .Z(n13676) );
  XOR U18039 ( .A(n13682), .B(n13683), .Z(n13310) );
  AND U18040 ( .A(n13684), .B(n13685), .Z(n13682) );
  AND U18041 ( .A(b[11]), .B(a[80]), .Z(n13681) );
  XOR U18042 ( .A(n13687), .B(n13688), .Z(n13315) );
  AND U18043 ( .A(n13689), .B(n13690), .Z(n13687) );
  AND U18044 ( .A(b[10]), .B(a[81]), .Z(n13686) );
  XOR U18045 ( .A(n13692), .B(n13693), .Z(n13320) );
  AND U18046 ( .A(n13694), .B(n13695), .Z(n13692) );
  AND U18047 ( .A(b[9]), .B(a[82]), .Z(n13691) );
  XOR U18048 ( .A(n13697), .B(n13698), .Z(n13325) );
  AND U18049 ( .A(n13699), .B(n13700), .Z(n13697) );
  AND U18050 ( .A(b[8]), .B(a[83]), .Z(n13696) );
  XOR U18051 ( .A(n13702), .B(n13703), .Z(n13330) );
  AND U18052 ( .A(n13704), .B(n13705), .Z(n13702) );
  AND U18053 ( .A(b[7]), .B(a[84]), .Z(n13701) );
  XOR U18054 ( .A(n13707), .B(n13708), .Z(n13335) );
  AND U18055 ( .A(n13709), .B(n13710), .Z(n13707) );
  AND U18056 ( .A(b[6]), .B(a[85]), .Z(n13706) );
  XOR U18057 ( .A(n13712), .B(n13713), .Z(n13340) );
  AND U18058 ( .A(n13714), .B(n13715), .Z(n13712) );
  AND U18059 ( .A(b[5]), .B(a[86]), .Z(n13711) );
  XOR U18060 ( .A(n13717), .B(n13718), .Z(n13345) );
  AND U18061 ( .A(n13719), .B(n13720), .Z(n13717) );
  AND U18062 ( .A(b[4]), .B(a[87]), .Z(n13716) );
  XOR U18063 ( .A(n13722), .B(n13723), .Z(n13350) );
  AND U18064 ( .A(n13724), .B(n13725), .Z(n13722) );
  AND U18065 ( .A(b[3]), .B(a[88]), .Z(n13721) );
  XOR U18066 ( .A(n13727), .B(n13728), .Z(n13355) );
  OR U18067 ( .A(n13729), .B(n13730), .Z(n13728) );
  AND U18068 ( .A(b[2]), .B(a[89]), .Z(n13726) );
  XNOR U18069 ( .A(n13365), .B(n13731), .Z(n13361) );
  NAND U18070 ( .A(b[1]), .B(a[90]), .Z(n13731) );
  IV U18071 ( .A(n13359), .Z(n13365) );
  ANDN U18072 ( .B(n10281), .A(n10283), .Z(n13359) );
  NAND U18073 ( .A(a[90]), .B(b[0]), .Z(n10283) );
  XOR U18074 ( .A(n13729), .B(n13730), .Z(n10281) );
  XOR U18075 ( .A(n13733), .B(n13724), .Z(n13732) );
  XOR U18076 ( .A(n13719), .B(n13723), .Z(n13734) );
  XOR U18077 ( .A(n13714), .B(n13718), .Z(n13735) );
  XOR U18078 ( .A(n13709), .B(n13713), .Z(n13736) );
  XOR U18079 ( .A(n13704), .B(n13708), .Z(n13737) );
  XOR U18080 ( .A(n13699), .B(n13703), .Z(n13738) );
  XOR U18081 ( .A(n13694), .B(n13698), .Z(n13739) );
  XOR U18082 ( .A(n13689), .B(n13693), .Z(n13740) );
  XOR U18083 ( .A(n13684), .B(n13688), .Z(n13741) );
  XOR U18084 ( .A(n13679), .B(n13683), .Z(n13742) );
  XOR U18085 ( .A(n13674), .B(n13678), .Z(n13743) );
  XOR U18086 ( .A(n13669), .B(n13673), .Z(n13744) );
  XOR U18087 ( .A(n13664), .B(n13668), .Z(n13745) );
  XOR U18088 ( .A(n13659), .B(n13663), .Z(n13746) );
  XOR U18089 ( .A(n13654), .B(n13658), .Z(n13747) );
  XOR U18090 ( .A(n13649), .B(n13653), .Z(n13748) );
  XOR U18091 ( .A(n13644), .B(n13648), .Z(n13749) );
  XOR U18092 ( .A(n13639), .B(n13643), .Z(n13750) );
  XOR U18093 ( .A(n13634), .B(n13638), .Z(n13751) );
  XOR U18094 ( .A(n13629), .B(n13633), .Z(n13752) );
  XOR U18095 ( .A(n13624), .B(n13628), .Z(n13753) );
  XOR U18096 ( .A(n13619), .B(n13623), .Z(n13754) );
  XOR U18097 ( .A(n13614), .B(n13618), .Z(n13755) );
  XOR U18098 ( .A(n13609), .B(n13613), .Z(n13756) );
  XOR U18099 ( .A(n13604), .B(n13608), .Z(n13757) );
  XOR U18100 ( .A(n13599), .B(n13603), .Z(n13758) );
  XOR U18101 ( .A(n13594), .B(n13598), .Z(n13759) );
  XOR U18102 ( .A(n13589), .B(n13593), .Z(n13760) );
  XOR U18103 ( .A(n13584), .B(n13588), .Z(n13761) );
  XOR U18104 ( .A(n13579), .B(n13583), .Z(n13762) );
  XOR U18105 ( .A(n13574), .B(n13578), .Z(n13763) );
  XOR U18106 ( .A(n13569), .B(n13573), .Z(n13764) );
  XOR U18107 ( .A(n13564), .B(n13568), .Z(n13765) );
  XOR U18108 ( .A(n13559), .B(n13563), .Z(n13766) );
  XOR U18109 ( .A(n13554), .B(n13558), .Z(n13767) );
  XOR U18110 ( .A(n13549), .B(n13553), .Z(n13768) );
  XOR U18111 ( .A(n13544), .B(n13548), .Z(n13769) );
  XOR U18112 ( .A(n13539), .B(n13543), .Z(n13770) );
  XOR U18113 ( .A(n13534), .B(n13538), .Z(n13771) );
  XOR U18114 ( .A(n13529), .B(n13533), .Z(n13772) );
  XOR U18115 ( .A(n13524), .B(n13528), .Z(n13773) );
  XOR U18116 ( .A(n13519), .B(n13523), .Z(n13774) );
  XOR U18117 ( .A(n13514), .B(n13518), .Z(n13775) );
  XOR U18118 ( .A(n13509), .B(n13513), .Z(n13776) );
  XOR U18119 ( .A(n13504), .B(n13508), .Z(n13777) );
  XOR U18120 ( .A(n13499), .B(n13503), .Z(n13778) );
  XOR U18121 ( .A(n13494), .B(n13498), .Z(n13779) );
  XOR U18122 ( .A(n13489), .B(n13493), .Z(n13780) );
  XOR U18123 ( .A(n13484), .B(n13488), .Z(n13781) );
  XOR U18124 ( .A(n13479), .B(n13483), .Z(n13782) );
  XOR U18125 ( .A(n13474), .B(n13478), .Z(n13783) );
  XOR U18126 ( .A(n13469), .B(n13473), .Z(n13784) );
  XOR U18127 ( .A(n13459), .B(n13468), .Z(n13785) );
  XOR U18128 ( .A(n13786), .B(n13458), .Z(n13459) );
  AND U18129 ( .A(a[36]), .B(b[54]), .Z(n13786) );
  XNOR U18130 ( .A(n13458), .B(n13464), .Z(n13787) );
  XNOR U18131 ( .A(n13463), .B(n13455), .Z(n13788) );
  XNOR U18132 ( .A(n13454), .B(n13450), .Z(n13789) );
  XNOR U18133 ( .A(n13449), .B(n13445), .Z(n13790) );
  XNOR U18134 ( .A(n13444), .B(n13440), .Z(n13791) );
  XOR U18135 ( .A(n13439), .B(n13436), .Z(n13792) );
  XOR U18136 ( .A(n13793), .B(n13794), .Z(n13436) );
  XOR U18137 ( .A(n13434), .B(n13795), .Z(n13794) );
  XOR U18138 ( .A(n13796), .B(n13797), .Z(n13795) );
  XOR U18139 ( .A(n13798), .B(n13799), .Z(n13797) );
  NAND U18140 ( .A(a[28]), .B(b[62]), .Z(n13799) );
  AND U18141 ( .A(a[27]), .B(b[63]), .Z(n13798) );
  XOR U18142 ( .A(n13800), .B(n13796), .Z(n13793) );
  XOR U18143 ( .A(n13801), .B(n13802), .Z(n13796) );
  ANDN U18144 ( .B(n13803), .A(n13804), .Z(n13801) );
  AND U18145 ( .A(a[29]), .B(b[61]), .Z(n13800) );
  XOR U18146 ( .A(n13805), .B(n13434), .Z(n13435) );
  XOR U18147 ( .A(n13806), .B(n13807), .Z(n13434) );
  AND U18148 ( .A(n13808), .B(n13809), .Z(n13806) );
  AND U18149 ( .A(a[30]), .B(b[60]), .Z(n13805) );
  XOR U18150 ( .A(n13810), .B(n13439), .Z(n13441) );
  XOR U18151 ( .A(n13811), .B(n13812), .Z(n13439) );
  AND U18152 ( .A(n13813), .B(n13814), .Z(n13811) );
  AND U18153 ( .A(a[31]), .B(b[59]), .Z(n13810) );
  XOR U18154 ( .A(n13815), .B(n13444), .Z(n13446) );
  XOR U18155 ( .A(n13816), .B(n13817), .Z(n13444) );
  AND U18156 ( .A(n13818), .B(n13819), .Z(n13816) );
  AND U18157 ( .A(a[32]), .B(b[58]), .Z(n13815) );
  XOR U18158 ( .A(n13820), .B(n13449), .Z(n13451) );
  XOR U18159 ( .A(n13821), .B(n13822), .Z(n13449) );
  AND U18160 ( .A(n13823), .B(n13824), .Z(n13821) );
  AND U18161 ( .A(a[33]), .B(b[57]), .Z(n13820) );
  XOR U18162 ( .A(n13825), .B(n13454), .Z(n13456) );
  XOR U18163 ( .A(n13826), .B(n13827), .Z(n13454) );
  AND U18164 ( .A(n13828), .B(n13829), .Z(n13826) );
  AND U18165 ( .A(a[34]), .B(b[56]), .Z(n13825) );
  XOR U18166 ( .A(n13830), .B(n13831), .Z(n13458) );
  AND U18167 ( .A(n13832), .B(n13833), .Z(n13830) );
  XOR U18168 ( .A(n13834), .B(n13463), .Z(n13465) );
  XOR U18169 ( .A(n13835), .B(n13836), .Z(n13463) );
  AND U18170 ( .A(n13837), .B(n13838), .Z(n13835) );
  AND U18171 ( .A(a[35]), .B(b[55]), .Z(n13834) );
  XOR U18172 ( .A(n13840), .B(n13841), .Z(n13468) );
  AND U18173 ( .A(n13842), .B(n13843), .Z(n13840) );
  AND U18174 ( .A(a[37]), .B(b[53]), .Z(n13839) );
  XOR U18175 ( .A(n13845), .B(n13846), .Z(n13473) );
  AND U18176 ( .A(n13847), .B(n13848), .Z(n13845) );
  AND U18177 ( .A(a[38]), .B(b[52]), .Z(n13844) );
  XOR U18178 ( .A(n13850), .B(n13851), .Z(n13478) );
  AND U18179 ( .A(n13852), .B(n13853), .Z(n13850) );
  AND U18180 ( .A(a[39]), .B(b[51]), .Z(n13849) );
  XOR U18181 ( .A(n13855), .B(n13856), .Z(n13483) );
  AND U18182 ( .A(n13857), .B(n13858), .Z(n13855) );
  AND U18183 ( .A(a[40]), .B(b[50]), .Z(n13854) );
  XOR U18184 ( .A(n13860), .B(n13861), .Z(n13488) );
  AND U18185 ( .A(n13862), .B(n13863), .Z(n13860) );
  AND U18186 ( .A(a[41]), .B(b[49]), .Z(n13859) );
  XOR U18187 ( .A(n13865), .B(n13866), .Z(n13493) );
  AND U18188 ( .A(n13867), .B(n13868), .Z(n13865) );
  AND U18189 ( .A(a[42]), .B(b[48]), .Z(n13864) );
  XOR U18190 ( .A(n13870), .B(n13871), .Z(n13498) );
  AND U18191 ( .A(n13872), .B(n13873), .Z(n13870) );
  AND U18192 ( .A(a[43]), .B(b[47]), .Z(n13869) );
  XOR U18193 ( .A(n13875), .B(n13876), .Z(n13503) );
  AND U18194 ( .A(n13877), .B(n13878), .Z(n13875) );
  AND U18195 ( .A(a[44]), .B(b[46]), .Z(n13874) );
  XOR U18196 ( .A(n13880), .B(n13881), .Z(n13508) );
  AND U18197 ( .A(n13882), .B(n13883), .Z(n13880) );
  AND U18198 ( .A(a[45]), .B(b[45]), .Z(n13879) );
  XOR U18199 ( .A(n13885), .B(n13886), .Z(n13513) );
  AND U18200 ( .A(n13887), .B(n13888), .Z(n13885) );
  AND U18201 ( .A(b[44]), .B(a[46]), .Z(n13884) );
  XOR U18202 ( .A(n13890), .B(n13891), .Z(n13518) );
  AND U18203 ( .A(n13892), .B(n13893), .Z(n13890) );
  AND U18204 ( .A(b[43]), .B(a[47]), .Z(n13889) );
  XOR U18205 ( .A(n13895), .B(n13896), .Z(n13523) );
  AND U18206 ( .A(n13897), .B(n13898), .Z(n13895) );
  AND U18207 ( .A(b[42]), .B(a[48]), .Z(n13894) );
  XOR U18208 ( .A(n13900), .B(n13901), .Z(n13528) );
  AND U18209 ( .A(n13902), .B(n13903), .Z(n13900) );
  AND U18210 ( .A(b[41]), .B(a[49]), .Z(n13899) );
  XOR U18211 ( .A(n13905), .B(n13906), .Z(n13533) );
  AND U18212 ( .A(n13907), .B(n13908), .Z(n13905) );
  AND U18213 ( .A(b[40]), .B(a[50]), .Z(n13904) );
  XOR U18214 ( .A(n13910), .B(n13911), .Z(n13538) );
  AND U18215 ( .A(n13912), .B(n13913), .Z(n13910) );
  AND U18216 ( .A(b[39]), .B(a[51]), .Z(n13909) );
  XOR U18217 ( .A(n13915), .B(n13916), .Z(n13543) );
  AND U18218 ( .A(n13917), .B(n13918), .Z(n13915) );
  AND U18219 ( .A(b[38]), .B(a[52]), .Z(n13914) );
  XOR U18220 ( .A(n13920), .B(n13921), .Z(n13548) );
  AND U18221 ( .A(n13922), .B(n13923), .Z(n13920) );
  AND U18222 ( .A(b[37]), .B(a[53]), .Z(n13919) );
  XOR U18223 ( .A(n13925), .B(n13926), .Z(n13553) );
  AND U18224 ( .A(n13927), .B(n13928), .Z(n13925) );
  AND U18225 ( .A(b[36]), .B(a[54]), .Z(n13924) );
  XOR U18226 ( .A(n13930), .B(n13931), .Z(n13558) );
  AND U18227 ( .A(n13932), .B(n13933), .Z(n13930) );
  AND U18228 ( .A(b[35]), .B(a[55]), .Z(n13929) );
  XOR U18229 ( .A(n13935), .B(n13936), .Z(n13563) );
  AND U18230 ( .A(n13937), .B(n13938), .Z(n13935) );
  AND U18231 ( .A(b[34]), .B(a[56]), .Z(n13934) );
  XOR U18232 ( .A(n13940), .B(n13941), .Z(n13568) );
  AND U18233 ( .A(n13942), .B(n13943), .Z(n13940) );
  AND U18234 ( .A(b[33]), .B(a[57]), .Z(n13939) );
  XOR U18235 ( .A(n13945), .B(n13946), .Z(n13573) );
  AND U18236 ( .A(n13947), .B(n13948), .Z(n13945) );
  AND U18237 ( .A(b[32]), .B(a[58]), .Z(n13944) );
  XOR U18238 ( .A(n13950), .B(n13951), .Z(n13578) );
  AND U18239 ( .A(n13952), .B(n13953), .Z(n13950) );
  AND U18240 ( .A(b[31]), .B(a[59]), .Z(n13949) );
  XOR U18241 ( .A(n13955), .B(n13956), .Z(n13583) );
  AND U18242 ( .A(n13957), .B(n13958), .Z(n13955) );
  AND U18243 ( .A(b[30]), .B(a[60]), .Z(n13954) );
  XOR U18244 ( .A(n13960), .B(n13961), .Z(n13588) );
  AND U18245 ( .A(n13962), .B(n13963), .Z(n13960) );
  AND U18246 ( .A(b[29]), .B(a[61]), .Z(n13959) );
  XOR U18247 ( .A(n13965), .B(n13966), .Z(n13593) );
  AND U18248 ( .A(n13967), .B(n13968), .Z(n13965) );
  AND U18249 ( .A(b[28]), .B(a[62]), .Z(n13964) );
  XOR U18250 ( .A(n13970), .B(n13971), .Z(n13598) );
  AND U18251 ( .A(n13972), .B(n13973), .Z(n13970) );
  AND U18252 ( .A(b[27]), .B(a[63]), .Z(n13969) );
  XOR U18253 ( .A(n13975), .B(n13976), .Z(n13603) );
  AND U18254 ( .A(n13977), .B(n13978), .Z(n13975) );
  AND U18255 ( .A(b[26]), .B(a[64]), .Z(n13974) );
  XOR U18256 ( .A(n13980), .B(n13981), .Z(n13608) );
  AND U18257 ( .A(n13982), .B(n13983), .Z(n13980) );
  AND U18258 ( .A(b[25]), .B(a[65]), .Z(n13979) );
  XOR U18259 ( .A(n13985), .B(n13986), .Z(n13613) );
  AND U18260 ( .A(n13987), .B(n13988), .Z(n13985) );
  AND U18261 ( .A(b[24]), .B(a[66]), .Z(n13984) );
  XOR U18262 ( .A(n13990), .B(n13991), .Z(n13618) );
  AND U18263 ( .A(n13992), .B(n13993), .Z(n13990) );
  AND U18264 ( .A(b[23]), .B(a[67]), .Z(n13989) );
  XOR U18265 ( .A(n13995), .B(n13996), .Z(n13623) );
  AND U18266 ( .A(n13997), .B(n13998), .Z(n13995) );
  AND U18267 ( .A(b[22]), .B(a[68]), .Z(n13994) );
  XOR U18268 ( .A(n14000), .B(n14001), .Z(n13628) );
  AND U18269 ( .A(n14002), .B(n14003), .Z(n14000) );
  AND U18270 ( .A(b[21]), .B(a[69]), .Z(n13999) );
  XOR U18271 ( .A(n14005), .B(n14006), .Z(n13633) );
  AND U18272 ( .A(n14007), .B(n14008), .Z(n14005) );
  AND U18273 ( .A(b[20]), .B(a[70]), .Z(n14004) );
  XOR U18274 ( .A(n14010), .B(n14011), .Z(n13638) );
  AND U18275 ( .A(n14012), .B(n14013), .Z(n14010) );
  AND U18276 ( .A(b[19]), .B(a[71]), .Z(n14009) );
  XOR U18277 ( .A(n14015), .B(n14016), .Z(n13643) );
  AND U18278 ( .A(n14017), .B(n14018), .Z(n14015) );
  AND U18279 ( .A(b[18]), .B(a[72]), .Z(n14014) );
  XOR U18280 ( .A(n14020), .B(n14021), .Z(n13648) );
  AND U18281 ( .A(n14022), .B(n14023), .Z(n14020) );
  AND U18282 ( .A(b[17]), .B(a[73]), .Z(n14019) );
  XOR U18283 ( .A(n14025), .B(n14026), .Z(n13653) );
  AND U18284 ( .A(n14027), .B(n14028), .Z(n14025) );
  AND U18285 ( .A(b[16]), .B(a[74]), .Z(n14024) );
  XOR U18286 ( .A(n14030), .B(n14031), .Z(n13658) );
  AND U18287 ( .A(n14032), .B(n14033), .Z(n14030) );
  AND U18288 ( .A(b[15]), .B(a[75]), .Z(n14029) );
  XOR U18289 ( .A(n14035), .B(n14036), .Z(n13663) );
  AND U18290 ( .A(n14037), .B(n14038), .Z(n14035) );
  AND U18291 ( .A(b[14]), .B(a[76]), .Z(n14034) );
  XOR U18292 ( .A(n14040), .B(n14041), .Z(n13668) );
  AND U18293 ( .A(n14042), .B(n14043), .Z(n14040) );
  AND U18294 ( .A(b[13]), .B(a[77]), .Z(n14039) );
  XOR U18295 ( .A(n14045), .B(n14046), .Z(n13673) );
  AND U18296 ( .A(n14047), .B(n14048), .Z(n14045) );
  AND U18297 ( .A(b[12]), .B(a[78]), .Z(n14044) );
  XOR U18298 ( .A(n14050), .B(n14051), .Z(n13678) );
  AND U18299 ( .A(n14052), .B(n14053), .Z(n14050) );
  AND U18300 ( .A(b[11]), .B(a[79]), .Z(n14049) );
  XOR U18301 ( .A(n14055), .B(n14056), .Z(n13683) );
  AND U18302 ( .A(n14057), .B(n14058), .Z(n14055) );
  AND U18303 ( .A(b[10]), .B(a[80]), .Z(n14054) );
  XOR U18304 ( .A(n14060), .B(n14061), .Z(n13688) );
  AND U18305 ( .A(n14062), .B(n14063), .Z(n14060) );
  AND U18306 ( .A(b[9]), .B(a[81]), .Z(n14059) );
  XOR U18307 ( .A(n14065), .B(n14066), .Z(n13693) );
  AND U18308 ( .A(n14067), .B(n14068), .Z(n14065) );
  AND U18309 ( .A(b[8]), .B(a[82]), .Z(n14064) );
  XOR U18310 ( .A(n14070), .B(n14071), .Z(n13698) );
  AND U18311 ( .A(n14072), .B(n14073), .Z(n14070) );
  AND U18312 ( .A(b[7]), .B(a[83]), .Z(n14069) );
  XOR U18313 ( .A(n14075), .B(n14076), .Z(n13703) );
  AND U18314 ( .A(n14077), .B(n14078), .Z(n14075) );
  AND U18315 ( .A(b[6]), .B(a[84]), .Z(n14074) );
  XOR U18316 ( .A(n14080), .B(n14081), .Z(n13708) );
  AND U18317 ( .A(n14082), .B(n14083), .Z(n14080) );
  AND U18318 ( .A(b[5]), .B(a[85]), .Z(n14079) );
  XOR U18319 ( .A(n14085), .B(n14086), .Z(n13713) );
  AND U18320 ( .A(n14087), .B(n14088), .Z(n14085) );
  AND U18321 ( .A(b[4]), .B(a[86]), .Z(n14084) );
  XOR U18322 ( .A(n14090), .B(n14091), .Z(n13718) );
  AND U18323 ( .A(n14092), .B(n14093), .Z(n14090) );
  AND U18324 ( .A(b[3]), .B(a[87]), .Z(n14089) );
  XOR U18325 ( .A(n14095), .B(n14096), .Z(n13723) );
  OR U18326 ( .A(n14097), .B(n14098), .Z(n14096) );
  AND U18327 ( .A(b[2]), .B(a[88]), .Z(n14094) );
  XNOR U18328 ( .A(n13733), .B(n14099), .Z(n13729) );
  NAND U18329 ( .A(b[1]), .B(a[89]), .Z(n14099) );
  IV U18330 ( .A(n13727), .Z(n13733) );
  ANDN U18331 ( .B(n10284), .A(n10286), .Z(n13727) );
  NAND U18332 ( .A(a[89]), .B(b[0]), .Z(n10286) );
  XOR U18333 ( .A(n14097), .B(n14098), .Z(n10284) );
  XOR U18334 ( .A(n14101), .B(n14092), .Z(n14100) );
  XOR U18335 ( .A(n14087), .B(n14091), .Z(n14102) );
  XOR U18336 ( .A(n14082), .B(n14086), .Z(n14103) );
  XOR U18337 ( .A(n14077), .B(n14081), .Z(n14104) );
  XOR U18338 ( .A(n14072), .B(n14076), .Z(n14105) );
  XOR U18339 ( .A(n14067), .B(n14071), .Z(n14106) );
  XOR U18340 ( .A(n14062), .B(n14066), .Z(n14107) );
  XOR U18341 ( .A(n14057), .B(n14061), .Z(n14108) );
  XOR U18342 ( .A(n14052), .B(n14056), .Z(n14109) );
  XOR U18343 ( .A(n14047), .B(n14051), .Z(n14110) );
  XOR U18344 ( .A(n14042), .B(n14046), .Z(n14111) );
  XOR U18345 ( .A(n14037), .B(n14041), .Z(n14112) );
  XOR U18346 ( .A(n14032), .B(n14036), .Z(n14113) );
  XOR U18347 ( .A(n14027), .B(n14031), .Z(n14114) );
  XOR U18348 ( .A(n14022), .B(n14026), .Z(n14115) );
  XOR U18349 ( .A(n14017), .B(n14021), .Z(n14116) );
  XOR U18350 ( .A(n14012), .B(n14016), .Z(n14117) );
  XOR U18351 ( .A(n14007), .B(n14011), .Z(n14118) );
  XOR U18352 ( .A(n14002), .B(n14006), .Z(n14119) );
  XOR U18353 ( .A(n13997), .B(n14001), .Z(n14120) );
  XOR U18354 ( .A(n13992), .B(n13996), .Z(n14121) );
  XOR U18355 ( .A(n13987), .B(n13991), .Z(n14122) );
  XOR U18356 ( .A(n13982), .B(n13986), .Z(n14123) );
  XOR U18357 ( .A(n13977), .B(n13981), .Z(n14124) );
  XOR U18358 ( .A(n13972), .B(n13976), .Z(n14125) );
  XOR U18359 ( .A(n13967), .B(n13971), .Z(n14126) );
  XOR U18360 ( .A(n13962), .B(n13966), .Z(n14127) );
  XOR U18361 ( .A(n13957), .B(n13961), .Z(n14128) );
  XOR U18362 ( .A(n13952), .B(n13956), .Z(n14129) );
  XOR U18363 ( .A(n13947), .B(n13951), .Z(n14130) );
  XOR U18364 ( .A(n13942), .B(n13946), .Z(n14131) );
  XOR U18365 ( .A(n13937), .B(n13941), .Z(n14132) );
  XOR U18366 ( .A(n13932), .B(n13936), .Z(n14133) );
  XOR U18367 ( .A(n13927), .B(n13931), .Z(n14134) );
  XOR U18368 ( .A(n13922), .B(n13926), .Z(n14135) );
  XOR U18369 ( .A(n13917), .B(n13921), .Z(n14136) );
  XOR U18370 ( .A(n13912), .B(n13916), .Z(n14137) );
  XOR U18371 ( .A(n13907), .B(n13911), .Z(n14138) );
  XOR U18372 ( .A(n13902), .B(n13906), .Z(n14139) );
  XOR U18373 ( .A(n13897), .B(n13901), .Z(n14140) );
  XOR U18374 ( .A(n13892), .B(n13896), .Z(n14141) );
  XOR U18375 ( .A(n13887), .B(n13891), .Z(n14142) );
  XOR U18376 ( .A(n13882), .B(n13886), .Z(n14143) );
  XOR U18377 ( .A(n13877), .B(n13881), .Z(n14144) );
  XOR U18378 ( .A(n13872), .B(n13876), .Z(n14145) );
  XOR U18379 ( .A(n13867), .B(n13871), .Z(n14146) );
  XOR U18380 ( .A(n13862), .B(n13866), .Z(n14147) );
  XOR U18381 ( .A(n13857), .B(n13861), .Z(n14148) );
  XOR U18382 ( .A(n13852), .B(n13856), .Z(n14149) );
  XOR U18383 ( .A(n13847), .B(n13851), .Z(n14150) );
  XOR U18384 ( .A(n13842), .B(n13846), .Z(n14151) );
  XOR U18385 ( .A(n13832), .B(n13841), .Z(n14152) );
  XOR U18386 ( .A(n14153), .B(n13831), .Z(n13832) );
  AND U18387 ( .A(a[36]), .B(b[53]), .Z(n14153) );
  XNOR U18388 ( .A(n13831), .B(n13837), .Z(n14154) );
  XNOR U18389 ( .A(n13836), .B(n13828), .Z(n14155) );
  XNOR U18390 ( .A(n13827), .B(n13823), .Z(n14156) );
  XNOR U18391 ( .A(n13822), .B(n13818), .Z(n14157) );
  XNOR U18392 ( .A(n13817), .B(n13813), .Z(n14158) );
  XNOR U18393 ( .A(n13812), .B(n13808), .Z(n14159) );
  XOR U18394 ( .A(n13807), .B(n13804), .Z(n14160) );
  XOR U18395 ( .A(n14161), .B(n14162), .Z(n13804) );
  XOR U18396 ( .A(n13802), .B(n14163), .Z(n14162) );
  XOR U18397 ( .A(n14164), .B(n14165), .Z(n14163) );
  XOR U18398 ( .A(n14166), .B(n14167), .Z(n14165) );
  NAND U18399 ( .A(a[27]), .B(b[62]), .Z(n14167) );
  AND U18400 ( .A(a[26]), .B(b[63]), .Z(n14166) );
  XOR U18401 ( .A(n14168), .B(n14164), .Z(n14161) );
  XOR U18402 ( .A(n14169), .B(n14170), .Z(n14164) );
  ANDN U18403 ( .B(n14171), .A(n14172), .Z(n14169) );
  AND U18404 ( .A(a[28]), .B(b[61]), .Z(n14168) );
  XOR U18405 ( .A(n14173), .B(n13802), .Z(n13803) );
  XOR U18406 ( .A(n14174), .B(n14175), .Z(n13802) );
  AND U18407 ( .A(n14176), .B(n14177), .Z(n14174) );
  AND U18408 ( .A(a[29]), .B(b[60]), .Z(n14173) );
  XOR U18409 ( .A(n14178), .B(n13807), .Z(n13809) );
  XOR U18410 ( .A(n14179), .B(n14180), .Z(n13807) );
  AND U18411 ( .A(n14181), .B(n14182), .Z(n14179) );
  AND U18412 ( .A(a[30]), .B(b[59]), .Z(n14178) );
  XOR U18413 ( .A(n14183), .B(n13812), .Z(n13814) );
  XOR U18414 ( .A(n14184), .B(n14185), .Z(n13812) );
  AND U18415 ( .A(n14186), .B(n14187), .Z(n14184) );
  AND U18416 ( .A(a[31]), .B(b[58]), .Z(n14183) );
  XOR U18417 ( .A(n14188), .B(n13817), .Z(n13819) );
  XOR U18418 ( .A(n14189), .B(n14190), .Z(n13817) );
  AND U18419 ( .A(n14191), .B(n14192), .Z(n14189) );
  AND U18420 ( .A(a[32]), .B(b[57]), .Z(n14188) );
  XOR U18421 ( .A(n14193), .B(n13822), .Z(n13824) );
  XOR U18422 ( .A(n14194), .B(n14195), .Z(n13822) );
  AND U18423 ( .A(n14196), .B(n14197), .Z(n14194) );
  AND U18424 ( .A(a[33]), .B(b[56]), .Z(n14193) );
  XOR U18425 ( .A(n14198), .B(n13827), .Z(n13829) );
  XOR U18426 ( .A(n14199), .B(n14200), .Z(n13827) );
  AND U18427 ( .A(n14201), .B(n14202), .Z(n14199) );
  AND U18428 ( .A(a[34]), .B(b[55]), .Z(n14198) );
  XOR U18429 ( .A(n14203), .B(n14204), .Z(n13831) );
  AND U18430 ( .A(n14205), .B(n14206), .Z(n14203) );
  XOR U18431 ( .A(n14207), .B(n13836), .Z(n13838) );
  XOR U18432 ( .A(n14208), .B(n14209), .Z(n13836) );
  AND U18433 ( .A(n14210), .B(n14211), .Z(n14208) );
  AND U18434 ( .A(a[35]), .B(b[54]), .Z(n14207) );
  XOR U18435 ( .A(n14213), .B(n14214), .Z(n13841) );
  AND U18436 ( .A(n14215), .B(n14216), .Z(n14213) );
  AND U18437 ( .A(a[37]), .B(b[52]), .Z(n14212) );
  XOR U18438 ( .A(n14218), .B(n14219), .Z(n13846) );
  AND U18439 ( .A(n14220), .B(n14221), .Z(n14218) );
  AND U18440 ( .A(a[38]), .B(b[51]), .Z(n14217) );
  XOR U18441 ( .A(n14223), .B(n14224), .Z(n13851) );
  AND U18442 ( .A(n14225), .B(n14226), .Z(n14223) );
  AND U18443 ( .A(a[39]), .B(b[50]), .Z(n14222) );
  XOR U18444 ( .A(n14228), .B(n14229), .Z(n13856) );
  AND U18445 ( .A(n14230), .B(n14231), .Z(n14228) );
  AND U18446 ( .A(a[40]), .B(b[49]), .Z(n14227) );
  XOR U18447 ( .A(n14233), .B(n14234), .Z(n13861) );
  AND U18448 ( .A(n14235), .B(n14236), .Z(n14233) );
  AND U18449 ( .A(a[41]), .B(b[48]), .Z(n14232) );
  XOR U18450 ( .A(n14238), .B(n14239), .Z(n13866) );
  AND U18451 ( .A(n14240), .B(n14241), .Z(n14238) );
  AND U18452 ( .A(a[42]), .B(b[47]), .Z(n14237) );
  XOR U18453 ( .A(n14243), .B(n14244), .Z(n13871) );
  AND U18454 ( .A(n14245), .B(n14246), .Z(n14243) );
  AND U18455 ( .A(a[43]), .B(b[46]), .Z(n14242) );
  XOR U18456 ( .A(n14248), .B(n14249), .Z(n13876) );
  AND U18457 ( .A(n14250), .B(n14251), .Z(n14248) );
  AND U18458 ( .A(a[44]), .B(b[45]), .Z(n14247) );
  XOR U18459 ( .A(n14253), .B(n14254), .Z(n13881) );
  AND U18460 ( .A(n14255), .B(n14256), .Z(n14253) );
  AND U18461 ( .A(b[44]), .B(a[45]), .Z(n14252) );
  XOR U18462 ( .A(n14258), .B(n14259), .Z(n13886) );
  AND U18463 ( .A(n14260), .B(n14261), .Z(n14258) );
  AND U18464 ( .A(b[43]), .B(a[46]), .Z(n14257) );
  XOR U18465 ( .A(n14263), .B(n14264), .Z(n13891) );
  AND U18466 ( .A(n14265), .B(n14266), .Z(n14263) );
  AND U18467 ( .A(b[42]), .B(a[47]), .Z(n14262) );
  XOR U18468 ( .A(n14268), .B(n14269), .Z(n13896) );
  AND U18469 ( .A(n14270), .B(n14271), .Z(n14268) );
  AND U18470 ( .A(b[41]), .B(a[48]), .Z(n14267) );
  XOR U18471 ( .A(n14273), .B(n14274), .Z(n13901) );
  AND U18472 ( .A(n14275), .B(n14276), .Z(n14273) );
  AND U18473 ( .A(b[40]), .B(a[49]), .Z(n14272) );
  XOR U18474 ( .A(n14278), .B(n14279), .Z(n13906) );
  AND U18475 ( .A(n14280), .B(n14281), .Z(n14278) );
  AND U18476 ( .A(b[39]), .B(a[50]), .Z(n14277) );
  XOR U18477 ( .A(n14283), .B(n14284), .Z(n13911) );
  AND U18478 ( .A(n14285), .B(n14286), .Z(n14283) );
  AND U18479 ( .A(b[38]), .B(a[51]), .Z(n14282) );
  XOR U18480 ( .A(n14288), .B(n14289), .Z(n13916) );
  AND U18481 ( .A(n14290), .B(n14291), .Z(n14288) );
  AND U18482 ( .A(b[37]), .B(a[52]), .Z(n14287) );
  XOR U18483 ( .A(n14293), .B(n14294), .Z(n13921) );
  AND U18484 ( .A(n14295), .B(n14296), .Z(n14293) );
  AND U18485 ( .A(b[36]), .B(a[53]), .Z(n14292) );
  XOR U18486 ( .A(n14298), .B(n14299), .Z(n13926) );
  AND U18487 ( .A(n14300), .B(n14301), .Z(n14298) );
  AND U18488 ( .A(b[35]), .B(a[54]), .Z(n14297) );
  XOR U18489 ( .A(n14303), .B(n14304), .Z(n13931) );
  AND U18490 ( .A(n14305), .B(n14306), .Z(n14303) );
  AND U18491 ( .A(b[34]), .B(a[55]), .Z(n14302) );
  XOR U18492 ( .A(n14308), .B(n14309), .Z(n13936) );
  AND U18493 ( .A(n14310), .B(n14311), .Z(n14308) );
  AND U18494 ( .A(b[33]), .B(a[56]), .Z(n14307) );
  XOR U18495 ( .A(n14313), .B(n14314), .Z(n13941) );
  AND U18496 ( .A(n14315), .B(n14316), .Z(n14313) );
  AND U18497 ( .A(b[32]), .B(a[57]), .Z(n14312) );
  XOR U18498 ( .A(n14318), .B(n14319), .Z(n13946) );
  AND U18499 ( .A(n14320), .B(n14321), .Z(n14318) );
  AND U18500 ( .A(b[31]), .B(a[58]), .Z(n14317) );
  XOR U18501 ( .A(n14323), .B(n14324), .Z(n13951) );
  AND U18502 ( .A(n14325), .B(n14326), .Z(n14323) );
  AND U18503 ( .A(b[30]), .B(a[59]), .Z(n14322) );
  XOR U18504 ( .A(n14328), .B(n14329), .Z(n13956) );
  AND U18505 ( .A(n14330), .B(n14331), .Z(n14328) );
  AND U18506 ( .A(b[29]), .B(a[60]), .Z(n14327) );
  XOR U18507 ( .A(n14333), .B(n14334), .Z(n13961) );
  AND U18508 ( .A(n14335), .B(n14336), .Z(n14333) );
  AND U18509 ( .A(b[28]), .B(a[61]), .Z(n14332) );
  XOR U18510 ( .A(n14338), .B(n14339), .Z(n13966) );
  AND U18511 ( .A(n14340), .B(n14341), .Z(n14338) );
  AND U18512 ( .A(b[27]), .B(a[62]), .Z(n14337) );
  XOR U18513 ( .A(n14343), .B(n14344), .Z(n13971) );
  AND U18514 ( .A(n14345), .B(n14346), .Z(n14343) );
  AND U18515 ( .A(b[26]), .B(a[63]), .Z(n14342) );
  XOR U18516 ( .A(n14348), .B(n14349), .Z(n13976) );
  AND U18517 ( .A(n14350), .B(n14351), .Z(n14348) );
  AND U18518 ( .A(b[25]), .B(a[64]), .Z(n14347) );
  XOR U18519 ( .A(n14353), .B(n14354), .Z(n13981) );
  AND U18520 ( .A(n14355), .B(n14356), .Z(n14353) );
  AND U18521 ( .A(b[24]), .B(a[65]), .Z(n14352) );
  XOR U18522 ( .A(n14358), .B(n14359), .Z(n13986) );
  AND U18523 ( .A(n14360), .B(n14361), .Z(n14358) );
  AND U18524 ( .A(b[23]), .B(a[66]), .Z(n14357) );
  XOR U18525 ( .A(n14363), .B(n14364), .Z(n13991) );
  AND U18526 ( .A(n14365), .B(n14366), .Z(n14363) );
  AND U18527 ( .A(b[22]), .B(a[67]), .Z(n14362) );
  XOR U18528 ( .A(n14368), .B(n14369), .Z(n13996) );
  AND U18529 ( .A(n14370), .B(n14371), .Z(n14368) );
  AND U18530 ( .A(b[21]), .B(a[68]), .Z(n14367) );
  XOR U18531 ( .A(n14373), .B(n14374), .Z(n14001) );
  AND U18532 ( .A(n14375), .B(n14376), .Z(n14373) );
  AND U18533 ( .A(b[20]), .B(a[69]), .Z(n14372) );
  XOR U18534 ( .A(n14378), .B(n14379), .Z(n14006) );
  AND U18535 ( .A(n14380), .B(n14381), .Z(n14378) );
  AND U18536 ( .A(b[19]), .B(a[70]), .Z(n14377) );
  XOR U18537 ( .A(n14383), .B(n14384), .Z(n14011) );
  AND U18538 ( .A(n14385), .B(n14386), .Z(n14383) );
  AND U18539 ( .A(b[18]), .B(a[71]), .Z(n14382) );
  XOR U18540 ( .A(n14388), .B(n14389), .Z(n14016) );
  AND U18541 ( .A(n14390), .B(n14391), .Z(n14388) );
  AND U18542 ( .A(b[17]), .B(a[72]), .Z(n14387) );
  XOR U18543 ( .A(n14393), .B(n14394), .Z(n14021) );
  AND U18544 ( .A(n14395), .B(n14396), .Z(n14393) );
  AND U18545 ( .A(b[16]), .B(a[73]), .Z(n14392) );
  XOR U18546 ( .A(n14398), .B(n14399), .Z(n14026) );
  AND U18547 ( .A(n14400), .B(n14401), .Z(n14398) );
  AND U18548 ( .A(b[15]), .B(a[74]), .Z(n14397) );
  XOR U18549 ( .A(n14403), .B(n14404), .Z(n14031) );
  AND U18550 ( .A(n14405), .B(n14406), .Z(n14403) );
  AND U18551 ( .A(b[14]), .B(a[75]), .Z(n14402) );
  XOR U18552 ( .A(n14408), .B(n14409), .Z(n14036) );
  AND U18553 ( .A(n14410), .B(n14411), .Z(n14408) );
  AND U18554 ( .A(b[13]), .B(a[76]), .Z(n14407) );
  XOR U18555 ( .A(n14413), .B(n14414), .Z(n14041) );
  AND U18556 ( .A(n14415), .B(n14416), .Z(n14413) );
  AND U18557 ( .A(b[12]), .B(a[77]), .Z(n14412) );
  XOR U18558 ( .A(n14418), .B(n14419), .Z(n14046) );
  AND U18559 ( .A(n14420), .B(n14421), .Z(n14418) );
  AND U18560 ( .A(b[11]), .B(a[78]), .Z(n14417) );
  XOR U18561 ( .A(n14423), .B(n14424), .Z(n14051) );
  AND U18562 ( .A(n14425), .B(n14426), .Z(n14423) );
  AND U18563 ( .A(b[10]), .B(a[79]), .Z(n14422) );
  XOR U18564 ( .A(n14428), .B(n14429), .Z(n14056) );
  AND U18565 ( .A(n14430), .B(n14431), .Z(n14428) );
  AND U18566 ( .A(b[9]), .B(a[80]), .Z(n14427) );
  XOR U18567 ( .A(n14433), .B(n14434), .Z(n14061) );
  AND U18568 ( .A(n14435), .B(n14436), .Z(n14433) );
  AND U18569 ( .A(b[8]), .B(a[81]), .Z(n14432) );
  XOR U18570 ( .A(n14438), .B(n14439), .Z(n14066) );
  AND U18571 ( .A(n14440), .B(n14441), .Z(n14438) );
  AND U18572 ( .A(b[7]), .B(a[82]), .Z(n14437) );
  XOR U18573 ( .A(n14443), .B(n14444), .Z(n14071) );
  AND U18574 ( .A(n14445), .B(n14446), .Z(n14443) );
  AND U18575 ( .A(b[6]), .B(a[83]), .Z(n14442) );
  XOR U18576 ( .A(n14448), .B(n14449), .Z(n14076) );
  AND U18577 ( .A(n14450), .B(n14451), .Z(n14448) );
  AND U18578 ( .A(b[5]), .B(a[84]), .Z(n14447) );
  XOR U18579 ( .A(n14453), .B(n14454), .Z(n14081) );
  AND U18580 ( .A(n14455), .B(n14456), .Z(n14453) );
  AND U18581 ( .A(b[4]), .B(a[85]), .Z(n14452) );
  XOR U18582 ( .A(n14458), .B(n14459), .Z(n14086) );
  AND U18583 ( .A(n14460), .B(n14461), .Z(n14458) );
  AND U18584 ( .A(b[3]), .B(a[86]), .Z(n14457) );
  XOR U18585 ( .A(n14463), .B(n14464), .Z(n14091) );
  OR U18586 ( .A(n14465), .B(n14466), .Z(n14464) );
  AND U18587 ( .A(b[2]), .B(a[87]), .Z(n14462) );
  XNOR U18588 ( .A(n14101), .B(n14467), .Z(n14097) );
  NAND U18589 ( .A(b[1]), .B(a[88]), .Z(n14467) );
  IV U18590 ( .A(n14095), .Z(n14101) );
  ANDN U18591 ( .B(n10287), .A(n10289), .Z(n14095) );
  NAND U18592 ( .A(a[88]), .B(b[0]), .Z(n10289) );
  XOR U18593 ( .A(n14465), .B(n14466), .Z(n10287) );
  XOR U18594 ( .A(n14469), .B(n14460), .Z(n14468) );
  XOR U18595 ( .A(n14455), .B(n14459), .Z(n14470) );
  XOR U18596 ( .A(n14450), .B(n14454), .Z(n14471) );
  XOR U18597 ( .A(n14445), .B(n14449), .Z(n14472) );
  XOR U18598 ( .A(n14440), .B(n14444), .Z(n14473) );
  XOR U18599 ( .A(n14435), .B(n14439), .Z(n14474) );
  XOR U18600 ( .A(n14430), .B(n14434), .Z(n14475) );
  XOR U18601 ( .A(n14425), .B(n14429), .Z(n14476) );
  XOR U18602 ( .A(n14420), .B(n14424), .Z(n14477) );
  XOR U18603 ( .A(n14415), .B(n14419), .Z(n14478) );
  XOR U18604 ( .A(n14410), .B(n14414), .Z(n14479) );
  XOR U18605 ( .A(n14405), .B(n14409), .Z(n14480) );
  XOR U18606 ( .A(n14400), .B(n14404), .Z(n14481) );
  XOR U18607 ( .A(n14395), .B(n14399), .Z(n14482) );
  XOR U18608 ( .A(n14390), .B(n14394), .Z(n14483) );
  XOR U18609 ( .A(n14385), .B(n14389), .Z(n14484) );
  XOR U18610 ( .A(n14380), .B(n14384), .Z(n14485) );
  XOR U18611 ( .A(n14375), .B(n14379), .Z(n14486) );
  XOR U18612 ( .A(n14370), .B(n14374), .Z(n14487) );
  XOR U18613 ( .A(n14365), .B(n14369), .Z(n14488) );
  XOR U18614 ( .A(n14360), .B(n14364), .Z(n14489) );
  XOR U18615 ( .A(n14355), .B(n14359), .Z(n14490) );
  XOR U18616 ( .A(n14350), .B(n14354), .Z(n14491) );
  XOR U18617 ( .A(n14345), .B(n14349), .Z(n14492) );
  XOR U18618 ( .A(n14340), .B(n14344), .Z(n14493) );
  XOR U18619 ( .A(n14335), .B(n14339), .Z(n14494) );
  XOR U18620 ( .A(n14330), .B(n14334), .Z(n14495) );
  XOR U18621 ( .A(n14325), .B(n14329), .Z(n14496) );
  XOR U18622 ( .A(n14320), .B(n14324), .Z(n14497) );
  XOR U18623 ( .A(n14315), .B(n14319), .Z(n14498) );
  XOR U18624 ( .A(n14310), .B(n14314), .Z(n14499) );
  XOR U18625 ( .A(n14305), .B(n14309), .Z(n14500) );
  XOR U18626 ( .A(n14300), .B(n14304), .Z(n14501) );
  XOR U18627 ( .A(n14295), .B(n14299), .Z(n14502) );
  XOR U18628 ( .A(n14290), .B(n14294), .Z(n14503) );
  XOR U18629 ( .A(n14285), .B(n14289), .Z(n14504) );
  XOR U18630 ( .A(n14280), .B(n14284), .Z(n14505) );
  XOR U18631 ( .A(n14275), .B(n14279), .Z(n14506) );
  XOR U18632 ( .A(n14270), .B(n14274), .Z(n14507) );
  XOR U18633 ( .A(n14265), .B(n14269), .Z(n14508) );
  XOR U18634 ( .A(n14260), .B(n14264), .Z(n14509) );
  XOR U18635 ( .A(n14255), .B(n14259), .Z(n14510) );
  XOR U18636 ( .A(n14250), .B(n14254), .Z(n14511) );
  XOR U18637 ( .A(n14245), .B(n14249), .Z(n14512) );
  XOR U18638 ( .A(n14240), .B(n14244), .Z(n14513) );
  XOR U18639 ( .A(n14235), .B(n14239), .Z(n14514) );
  XOR U18640 ( .A(n14230), .B(n14234), .Z(n14515) );
  XOR U18641 ( .A(n14225), .B(n14229), .Z(n14516) );
  XOR U18642 ( .A(n14220), .B(n14224), .Z(n14517) );
  XOR U18643 ( .A(n14215), .B(n14219), .Z(n14518) );
  XOR U18644 ( .A(n14205), .B(n14214), .Z(n14519) );
  XOR U18645 ( .A(n14520), .B(n14204), .Z(n14205) );
  AND U18646 ( .A(a[36]), .B(b[52]), .Z(n14520) );
  XNOR U18647 ( .A(n14204), .B(n14210), .Z(n14521) );
  XNOR U18648 ( .A(n14209), .B(n14201), .Z(n14522) );
  XNOR U18649 ( .A(n14200), .B(n14196), .Z(n14523) );
  XNOR U18650 ( .A(n14195), .B(n14191), .Z(n14524) );
  XNOR U18651 ( .A(n14190), .B(n14186), .Z(n14525) );
  XNOR U18652 ( .A(n14185), .B(n14181), .Z(n14526) );
  XNOR U18653 ( .A(n14180), .B(n14176), .Z(n14527) );
  XOR U18654 ( .A(n14175), .B(n14172), .Z(n14528) );
  XOR U18655 ( .A(n14529), .B(n14530), .Z(n14172) );
  XOR U18656 ( .A(n14170), .B(n14531), .Z(n14530) );
  XOR U18657 ( .A(n14532), .B(n14533), .Z(n14531) );
  XOR U18658 ( .A(n14534), .B(n14535), .Z(n14533) );
  NAND U18659 ( .A(a[26]), .B(b[62]), .Z(n14535) );
  AND U18660 ( .A(a[25]), .B(b[63]), .Z(n14534) );
  XOR U18661 ( .A(n14536), .B(n14532), .Z(n14529) );
  XOR U18662 ( .A(n14537), .B(n14538), .Z(n14532) );
  ANDN U18663 ( .B(n14539), .A(n14540), .Z(n14537) );
  AND U18664 ( .A(a[27]), .B(b[61]), .Z(n14536) );
  XOR U18665 ( .A(n14541), .B(n14170), .Z(n14171) );
  XOR U18666 ( .A(n14542), .B(n14543), .Z(n14170) );
  AND U18667 ( .A(n14544), .B(n14545), .Z(n14542) );
  AND U18668 ( .A(a[28]), .B(b[60]), .Z(n14541) );
  XOR U18669 ( .A(n14546), .B(n14175), .Z(n14177) );
  XOR U18670 ( .A(n14547), .B(n14548), .Z(n14175) );
  AND U18671 ( .A(n14549), .B(n14550), .Z(n14547) );
  AND U18672 ( .A(a[29]), .B(b[59]), .Z(n14546) );
  XOR U18673 ( .A(n14551), .B(n14180), .Z(n14182) );
  XOR U18674 ( .A(n14552), .B(n14553), .Z(n14180) );
  AND U18675 ( .A(n14554), .B(n14555), .Z(n14552) );
  AND U18676 ( .A(a[30]), .B(b[58]), .Z(n14551) );
  XOR U18677 ( .A(n14556), .B(n14185), .Z(n14187) );
  XOR U18678 ( .A(n14557), .B(n14558), .Z(n14185) );
  AND U18679 ( .A(n14559), .B(n14560), .Z(n14557) );
  AND U18680 ( .A(a[31]), .B(b[57]), .Z(n14556) );
  XOR U18681 ( .A(n14561), .B(n14190), .Z(n14192) );
  XOR U18682 ( .A(n14562), .B(n14563), .Z(n14190) );
  AND U18683 ( .A(n14564), .B(n14565), .Z(n14562) );
  AND U18684 ( .A(a[32]), .B(b[56]), .Z(n14561) );
  XOR U18685 ( .A(n14566), .B(n14195), .Z(n14197) );
  XOR U18686 ( .A(n14567), .B(n14568), .Z(n14195) );
  AND U18687 ( .A(n14569), .B(n14570), .Z(n14567) );
  AND U18688 ( .A(a[33]), .B(b[55]), .Z(n14566) );
  XOR U18689 ( .A(n14571), .B(n14200), .Z(n14202) );
  XOR U18690 ( .A(n14572), .B(n14573), .Z(n14200) );
  AND U18691 ( .A(n14574), .B(n14575), .Z(n14572) );
  AND U18692 ( .A(a[34]), .B(b[54]), .Z(n14571) );
  XOR U18693 ( .A(n14576), .B(n14577), .Z(n14204) );
  AND U18694 ( .A(n14578), .B(n14579), .Z(n14576) );
  XOR U18695 ( .A(n14580), .B(n14209), .Z(n14211) );
  XOR U18696 ( .A(n14581), .B(n14582), .Z(n14209) );
  AND U18697 ( .A(n14583), .B(n14584), .Z(n14581) );
  AND U18698 ( .A(a[35]), .B(b[53]), .Z(n14580) );
  XOR U18699 ( .A(n14586), .B(n14587), .Z(n14214) );
  AND U18700 ( .A(n14588), .B(n14589), .Z(n14586) );
  AND U18701 ( .A(a[37]), .B(b[51]), .Z(n14585) );
  XOR U18702 ( .A(n14591), .B(n14592), .Z(n14219) );
  AND U18703 ( .A(n14593), .B(n14594), .Z(n14591) );
  AND U18704 ( .A(a[38]), .B(b[50]), .Z(n14590) );
  XOR U18705 ( .A(n14596), .B(n14597), .Z(n14224) );
  AND U18706 ( .A(n14598), .B(n14599), .Z(n14596) );
  AND U18707 ( .A(a[39]), .B(b[49]), .Z(n14595) );
  XOR U18708 ( .A(n14601), .B(n14602), .Z(n14229) );
  AND U18709 ( .A(n14603), .B(n14604), .Z(n14601) );
  AND U18710 ( .A(a[40]), .B(b[48]), .Z(n14600) );
  XOR U18711 ( .A(n14606), .B(n14607), .Z(n14234) );
  AND U18712 ( .A(n14608), .B(n14609), .Z(n14606) );
  AND U18713 ( .A(a[41]), .B(b[47]), .Z(n14605) );
  XOR U18714 ( .A(n14611), .B(n14612), .Z(n14239) );
  AND U18715 ( .A(n14613), .B(n14614), .Z(n14611) );
  AND U18716 ( .A(a[42]), .B(b[46]), .Z(n14610) );
  XOR U18717 ( .A(n14616), .B(n14617), .Z(n14244) );
  AND U18718 ( .A(n14618), .B(n14619), .Z(n14616) );
  AND U18719 ( .A(a[43]), .B(b[45]), .Z(n14615) );
  XOR U18720 ( .A(n14621), .B(n14622), .Z(n14249) );
  AND U18721 ( .A(n14623), .B(n14624), .Z(n14621) );
  AND U18722 ( .A(a[44]), .B(b[44]), .Z(n14620) );
  XOR U18723 ( .A(n14626), .B(n14627), .Z(n14254) );
  AND U18724 ( .A(n14628), .B(n14629), .Z(n14626) );
  AND U18725 ( .A(b[43]), .B(a[45]), .Z(n14625) );
  XOR U18726 ( .A(n14631), .B(n14632), .Z(n14259) );
  AND U18727 ( .A(n14633), .B(n14634), .Z(n14631) );
  AND U18728 ( .A(b[42]), .B(a[46]), .Z(n14630) );
  XOR U18729 ( .A(n14636), .B(n14637), .Z(n14264) );
  AND U18730 ( .A(n14638), .B(n14639), .Z(n14636) );
  AND U18731 ( .A(b[41]), .B(a[47]), .Z(n14635) );
  XOR U18732 ( .A(n14641), .B(n14642), .Z(n14269) );
  AND U18733 ( .A(n14643), .B(n14644), .Z(n14641) );
  AND U18734 ( .A(b[40]), .B(a[48]), .Z(n14640) );
  XOR U18735 ( .A(n14646), .B(n14647), .Z(n14274) );
  AND U18736 ( .A(n14648), .B(n14649), .Z(n14646) );
  AND U18737 ( .A(b[39]), .B(a[49]), .Z(n14645) );
  XOR U18738 ( .A(n14651), .B(n14652), .Z(n14279) );
  AND U18739 ( .A(n14653), .B(n14654), .Z(n14651) );
  AND U18740 ( .A(b[38]), .B(a[50]), .Z(n14650) );
  XOR U18741 ( .A(n14656), .B(n14657), .Z(n14284) );
  AND U18742 ( .A(n14658), .B(n14659), .Z(n14656) );
  AND U18743 ( .A(b[37]), .B(a[51]), .Z(n14655) );
  XOR U18744 ( .A(n14661), .B(n14662), .Z(n14289) );
  AND U18745 ( .A(n14663), .B(n14664), .Z(n14661) );
  AND U18746 ( .A(b[36]), .B(a[52]), .Z(n14660) );
  XOR U18747 ( .A(n14666), .B(n14667), .Z(n14294) );
  AND U18748 ( .A(n14668), .B(n14669), .Z(n14666) );
  AND U18749 ( .A(b[35]), .B(a[53]), .Z(n14665) );
  XOR U18750 ( .A(n14671), .B(n14672), .Z(n14299) );
  AND U18751 ( .A(n14673), .B(n14674), .Z(n14671) );
  AND U18752 ( .A(b[34]), .B(a[54]), .Z(n14670) );
  XOR U18753 ( .A(n14676), .B(n14677), .Z(n14304) );
  AND U18754 ( .A(n14678), .B(n14679), .Z(n14676) );
  AND U18755 ( .A(b[33]), .B(a[55]), .Z(n14675) );
  XOR U18756 ( .A(n14681), .B(n14682), .Z(n14309) );
  AND U18757 ( .A(n14683), .B(n14684), .Z(n14681) );
  AND U18758 ( .A(b[32]), .B(a[56]), .Z(n14680) );
  XOR U18759 ( .A(n14686), .B(n14687), .Z(n14314) );
  AND U18760 ( .A(n14688), .B(n14689), .Z(n14686) );
  AND U18761 ( .A(b[31]), .B(a[57]), .Z(n14685) );
  XOR U18762 ( .A(n14691), .B(n14692), .Z(n14319) );
  AND U18763 ( .A(n14693), .B(n14694), .Z(n14691) );
  AND U18764 ( .A(b[30]), .B(a[58]), .Z(n14690) );
  XOR U18765 ( .A(n14696), .B(n14697), .Z(n14324) );
  AND U18766 ( .A(n14698), .B(n14699), .Z(n14696) );
  AND U18767 ( .A(b[29]), .B(a[59]), .Z(n14695) );
  XOR U18768 ( .A(n14701), .B(n14702), .Z(n14329) );
  AND U18769 ( .A(n14703), .B(n14704), .Z(n14701) );
  AND U18770 ( .A(b[28]), .B(a[60]), .Z(n14700) );
  XOR U18771 ( .A(n14706), .B(n14707), .Z(n14334) );
  AND U18772 ( .A(n14708), .B(n14709), .Z(n14706) );
  AND U18773 ( .A(b[27]), .B(a[61]), .Z(n14705) );
  XOR U18774 ( .A(n14711), .B(n14712), .Z(n14339) );
  AND U18775 ( .A(n14713), .B(n14714), .Z(n14711) );
  AND U18776 ( .A(b[26]), .B(a[62]), .Z(n14710) );
  XOR U18777 ( .A(n14716), .B(n14717), .Z(n14344) );
  AND U18778 ( .A(n14718), .B(n14719), .Z(n14716) );
  AND U18779 ( .A(b[25]), .B(a[63]), .Z(n14715) );
  XOR U18780 ( .A(n14721), .B(n14722), .Z(n14349) );
  AND U18781 ( .A(n14723), .B(n14724), .Z(n14721) );
  AND U18782 ( .A(b[24]), .B(a[64]), .Z(n14720) );
  XOR U18783 ( .A(n14726), .B(n14727), .Z(n14354) );
  AND U18784 ( .A(n14728), .B(n14729), .Z(n14726) );
  AND U18785 ( .A(b[23]), .B(a[65]), .Z(n14725) );
  XOR U18786 ( .A(n14731), .B(n14732), .Z(n14359) );
  AND U18787 ( .A(n14733), .B(n14734), .Z(n14731) );
  AND U18788 ( .A(b[22]), .B(a[66]), .Z(n14730) );
  XOR U18789 ( .A(n14736), .B(n14737), .Z(n14364) );
  AND U18790 ( .A(n14738), .B(n14739), .Z(n14736) );
  AND U18791 ( .A(b[21]), .B(a[67]), .Z(n14735) );
  XOR U18792 ( .A(n14741), .B(n14742), .Z(n14369) );
  AND U18793 ( .A(n14743), .B(n14744), .Z(n14741) );
  AND U18794 ( .A(b[20]), .B(a[68]), .Z(n14740) );
  XOR U18795 ( .A(n14746), .B(n14747), .Z(n14374) );
  AND U18796 ( .A(n14748), .B(n14749), .Z(n14746) );
  AND U18797 ( .A(b[19]), .B(a[69]), .Z(n14745) );
  XOR U18798 ( .A(n14751), .B(n14752), .Z(n14379) );
  AND U18799 ( .A(n14753), .B(n14754), .Z(n14751) );
  AND U18800 ( .A(b[18]), .B(a[70]), .Z(n14750) );
  XOR U18801 ( .A(n14756), .B(n14757), .Z(n14384) );
  AND U18802 ( .A(n14758), .B(n14759), .Z(n14756) );
  AND U18803 ( .A(b[17]), .B(a[71]), .Z(n14755) );
  XOR U18804 ( .A(n14761), .B(n14762), .Z(n14389) );
  AND U18805 ( .A(n14763), .B(n14764), .Z(n14761) );
  AND U18806 ( .A(b[16]), .B(a[72]), .Z(n14760) );
  XOR U18807 ( .A(n14766), .B(n14767), .Z(n14394) );
  AND U18808 ( .A(n14768), .B(n14769), .Z(n14766) );
  AND U18809 ( .A(b[15]), .B(a[73]), .Z(n14765) );
  XOR U18810 ( .A(n14771), .B(n14772), .Z(n14399) );
  AND U18811 ( .A(n14773), .B(n14774), .Z(n14771) );
  AND U18812 ( .A(b[14]), .B(a[74]), .Z(n14770) );
  XOR U18813 ( .A(n14776), .B(n14777), .Z(n14404) );
  AND U18814 ( .A(n14778), .B(n14779), .Z(n14776) );
  AND U18815 ( .A(b[13]), .B(a[75]), .Z(n14775) );
  XOR U18816 ( .A(n14781), .B(n14782), .Z(n14409) );
  AND U18817 ( .A(n14783), .B(n14784), .Z(n14781) );
  AND U18818 ( .A(b[12]), .B(a[76]), .Z(n14780) );
  XOR U18819 ( .A(n14786), .B(n14787), .Z(n14414) );
  AND U18820 ( .A(n14788), .B(n14789), .Z(n14786) );
  AND U18821 ( .A(b[11]), .B(a[77]), .Z(n14785) );
  XOR U18822 ( .A(n14791), .B(n14792), .Z(n14419) );
  AND U18823 ( .A(n14793), .B(n14794), .Z(n14791) );
  AND U18824 ( .A(b[10]), .B(a[78]), .Z(n14790) );
  XOR U18825 ( .A(n14796), .B(n14797), .Z(n14424) );
  AND U18826 ( .A(n14798), .B(n14799), .Z(n14796) );
  AND U18827 ( .A(b[9]), .B(a[79]), .Z(n14795) );
  XOR U18828 ( .A(n14801), .B(n14802), .Z(n14429) );
  AND U18829 ( .A(n14803), .B(n14804), .Z(n14801) );
  AND U18830 ( .A(b[8]), .B(a[80]), .Z(n14800) );
  XOR U18831 ( .A(n14806), .B(n14807), .Z(n14434) );
  AND U18832 ( .A(n14808), .B(n14809), .Z(n14806) );
  AND U18833 ( .A(b[7]), .B(a[81]), .Z(n14805) );
  XOR U18834 ( .A(n14811), .B(n14812), .Z(n14439) );
  AND U18835 ( .A(n14813), .B(n14814), .Z(n14811) );
  AND U18836 ( .A(b[6]), .B(a[82]), .Z(n14810) );
  XOR U18837 ( .A(n14816), .B(n14817), .Z(n14444) );
  AND U18838 ( .A(n14818), .B(n14819), .Z(n14816) );
  AND U18839 ( .A(b[5]), .B(a[83]), .Z(n14815) );
  XOR U18840 ( .A(n14821), .B(n14822), .Z(n14449) );
  AND U18841 ( .A(n14823), .B(n14824), .Z(n14821) );
  AND U18842 ( .A(b[4]), .B(a[84]), .Z(n14820) );
  XOR U18843 ( .A(n14826), .B(n14827), .Z(n14454) );
  AND U18844 ( .A(n14828), .B(n14829), .Z(n14826) );
  AND U18845 ( .A(b[3]), .B(a[85]), .Z(n14825) );
  XOR U18846 ( .A(n14831), .B(n14832), .Z(n14459) );
  OR U18847 ( .A(n14833), .B(n14834), .Z(n14832) );
  AND U18848 ( .A(b[2]), .B(a[86]), .Z(n14830) );
  XNOR U18849 ( .A(n14469), .B(n14835), .Z(n14465) );
  NAND U18850 ( .A(b[1]), .B(a[87]), .Z(n14835) );
  IV U18851 ( .A(n14463), .Z(n14469) );
  ANDN U18852 ( .B(n10290), .A(n10292), .Z(n14463) );
  NAND U18853 ( .A(a[87]), .B(b[0]), .Z(n10292) );
  XOR U18854 ( .A(n14833), .B(n14834), .Z(n10290) );
  XOR U18855 ( .A(n14837), .B(n14828), .Z(n14836) );
  XOR U18856 ( .A(n14823), .B(n14827), .Z(n14838) );
  XOR U18857 ( .A(n14818), .B(n14822), .Z(n14839) );
  XOR U18858 ( .A(n14813), .B(n14817), .Z(n14840) );
  XOR U18859 ( .A(n14808), .B(n14812), .Z(n14841) );
  XOR U18860 ( .A(n14803), .B(n14807), .Z(n14842) );
  XOR U18861 ( .A(n14798), .B(n14802), .Z(n14843) );
  XOR U18862 ( .A(n14793), .B(n14797), .Z(n14844) );
  XOR U18863 ( .A(n14788), .B(n14792), .Z(n14845) );
  XOR U18864 ( .A(n14783), .B(n14787), .Z(n14846) );
  XOR U18865 ( .A(n14778), .B(n14782), .Z(n14847) );
  XOR U18866 ( .A(n14773), .B(n14777), .Z(n14848) );
  XOR U18867 ( .A(n14768), .B(n14772), .Z(n14849) );
  XOR U18868 ( .A(n14763), .B(n14767), .Z(n14850) );
  XOR U18869 ( .A(n14758), .B(n14762), .Z(n14851) );
  XOR U18870 ( .A(n14753), .B(n14757), .Z(n14852) );
  XOR U18871 ( .A(n14748), .B(n14752), .Z(n14853) );
  XOR U18872 ( .A(n14743), .B(n14747), .Z(n14854) );
  XOR U18873 ( .A(n14738), .B(n14742), .Z(n14855) );
  XOR U18874 ( .A(n14733), .B(n14737), .Z(n14856) );
  XOR U18875 ( .A(n14728), .B(n14732), .Z(n14857) );
  XOR U18876 ( .A(n14723), .B(n14727), .Z(n14858) );
  XOR U18877 ( .A(n14718), .B(n14722), .Z(n14859) );
  XOR U18878 ( .A(n14713), .B(n14717), .Z(n14860) );
  XOR U18879 ( .A(n14708), .B(n14712), .Z(n14861) );
  XOR U18880 ( .A(n14703), .B(n14707), .Z(n14862) );
  XOR U18881 ( .A(n14698), .B(n14702), .Z(n14863) );
  XOR U18882 ( .A(n14693), .B(n14697), .Z(n14864) );
  XOR U18883 ( .A(n14688), .B(n14692), .Z(n14865) );
  XOR U18884 ( .A(n14683), .B(n14687), .Z(n14866) );
  XOR U18885 ( .A(n14678), .B(n14682), .Z(n14867) );
  XOR U18886 ( .A(n14673), .B(n14677), .Z(n14868) );
  XOR U18887 ( .A(n14668), .B(n14672), .Z(n14869) );
  XOR U18888 ( .A(n14663), .B(n14667), .Z(n14870) );
  XOR U18889 ( .A(n14658), .B(n14662), .Z(n14871) );
  XOR U18890 ( .A(n14653), .B(n14657), .Z(n14872) );
  XOR U18891 ( .A(n14648), .B(n14652), .Z(n14873) );
  XOR U18892 ( .A(n14643), .B(n14647), .Z(n14874) );
  XOR U18893 ( .A(n14638), .B(n14642), .Z(n14875) );
  XOR U18894 ( .A(n14633), .B(n14637), .Z(n14876) );
  XOR U18895 ( .A(n14628), .B(n14632), .Z(n14877) );
  XOR U18896 ( .A(n14623), .B(n14627), .Z(n14878) );
  XOR U18897 ( .A(n14618), .B(n14622), .Z(n14879) );
  XOR U18898 ( .A(n14613), .B(n14617), .Z(n14880) );
  XOR U18899 ( .A(n14608), .B(n14612), .Z(n14881) );
  XOR U18900 ( .A(n14603), .B(n14607), .Z(n14882) );
  XOR U18901 ( .A(n14598), .B(n14602), .Z(n14883) );
  XOR U18902 ( .A(n14593), .B(n14597), .Z(n14884) );
  XOR U18903 ( .A(n14588), .B(n14592), .Z(n14885) );
  XOR U18904 ( .A(n14578), .B(n14587), .Z(n14886) );
  XOR U18905 ( .A(n14887), .B(n14577), .Z(n14578) );
  AND U18906 ( .A(a[36]), .B(b[51]), .Z(n14887) );
  XNOR U18907 ( .A(n14577), .B(n14583), .Z(n14888) );
  XNOR U18908 ( .A(n14582), .B(n14574), .Z(n14889) );
  XNOR U18909 ( .A(n14573), .B(n14569), .Z(n14890) );
  XNOR U18910 ( .A(n14568), .B(n14564), .Z(n14891) );
  XNOR U18911 ( .A(n14563), .B(n14559), .Z(n14892) );
  XNOR U18912 ( .A(n14558), .B(n14554), .Z(n14893) );
  XNOR U18913 ( .A(n14553), .B(n14549), .Z(n14894) );
  XNOR U18914 ( .A(n14548), .B(n14544), .Z(n14895) );
  XOR U18915 ( .A(n14543), .B(n14540), .Z(n14896) );
  XOR U18916 ( .A(n14897), .B(n14898), .Z(n14540) );
  XOR U18917 ( .A(n14538), .B(n14899), .Z(n14898) );
  XOR U18918 ( .A(n14900), .B(n14901), .Z(n14899) );
  XOR U18919 ( .A(n14902), .B(n14903), .Z(n14901) );
  NAND U18920 ( .A(a[25]), .B(b[62]), .Z(n14903) );
  AND U18921 ( .A(a[24]), .B(b[63]), .Z(n14902) );
  XOR U18922 ( .A(n14904), .B(n14900), .Z(n14897) );
  XOR U18923 ( .A(n14905), .B(n14906), .Z(n14900) );
  ANDN U18924 ( .B(n14907), .A(n14908), .Z(n14905) );
  AND U18925 ( .A(a[26]), .B(b[61]), .Z(n14904) );
  XOR U18926 ( .A(n14909), .B(n14538), .Z(n14539) );
  XOR U18927 ( .A(n14910), .B(n14911), .Z(n14538) );
  AND U18928 ( .A(n14912), .B(n14913), .Z(n14910) );
  AND U18929 ( .A(a[27]), .B(b[60]), .Z(n14909) );
  XOR U18930 ( .A(n14914), .B(n14543), .Z(n14545) );
  XOR U18931 ( .A(n14915), .B(n14916), .Z(n14543) );
  AND U18932 ( .A(n14917), .B(n14918), .Z(n14915) );
  AND U18933 ( .A(a[28]), .B(b[59]), .Z(n14914) );
  XOR U18934 ( .A(n14919), .B(n14548), .Z(n14550) );
  XOR U18935 ( .A(n14920), .B(n14921), .Z(n14548) );
  AND U18936 ( .A(n14922), .B(n14923), .Z(n14920) );
  AND U18937 ( .A(a[29]), .B(b[58]), .Z(n14919) );
  XOR U18938 ( .A(n14924), .B(n14553), .Z(n14555) );
  XOR U18939 ( .A(n14925), .B(n14926), .Z(n14553) );
  AND U18940 ( .A(n14927), .B(n14928), .Z(n14925) );
  AND U18941 ( .A(a[30]), .B(b[57]), .Z(n14924) );
  XOR U18942 ( .A(n14929), .B(n14558), .Z(n14560) );
  XOR U18943 ( .A(n14930), .B(n14931), .Z(n14558) );
  AND U18944 ( .A(n14932), .B(n14933), .Z(n14930) );
  AND U18945 ( .A(a[31]), .B(b[56]), .Z(n14929) );
  XOR U18946 ( .A(n14934), .B(n14563), .Z(n14565) );
  XOR U18947 ( .A(n14935), .B(n14936), .Z(n14563) );
  AND U18948 ( .A(n14937), .B(n14938), .Z(n14935) );
  AND U18949 ( .A(a[32]), .B(b[55]), .Z(n14934) );
  XOR U18950 ( .A(n14939), .B(n14568), .Z(n14570) );
  XOR U18951 ( .A(n14940), .B(n14941), .Z(n14568) );
  AND U18952 ( .A(n14942), .B(n14943), .Z(n14940) );
  AND U18953 ( .A(a[33]), .B(b[54]), .Z(n14939) );
  XOR U18954 ( .A(n14944), .B(n14573), .Z(n14575) );
  XOR U18955 ( .A(n14945), .B(n14946), .Z(n14573) );
  AND U18956 ( .A(n14947), .B(n14948), .Z(n14945) );
  AND U18957 ( .A(a[34]), .B(b[53]), .Z(n14944) );
  XOR U18958 ( .A(n14949), .B(n14950), .Z(n14577) );
  AND U18959 ( .A(n14951), .B(n14952), .Z(n14949) );
  XOR U18960 ( .A(n14953), .B(n14582), .Z(n14584) );
  XOR U18961 ( .A(n14954), .B(n14955), .Z(n14582) );
  AND U18962 ( .A(n14956), .B(n14957), .Z(n14954) );
  AND U18963 ( .A(a[35]), .B(b[52]), .Z(n14953) );
  XOR U18964 ( .A(n14959), .B(n14960), .Z(n14587) );
  AND U18965 ( .A(n14961), .B(n14962), .Z(n14959) );
  AND U18966 ( .A(a[37]), .B(b[50]), .Z(n14958) );
  XOR U18967 ( .A(n14964), .B(n14965), .Z(n14592) );
  AND U18968 ( .A(n14966), .B(n14967), .Z(n14964) );
  AND U18969 ( .A(a[38]), .B(b[49]), .Z(n14963) );
  XOR U18970 ( .A(n14969), .B(n14970), .Z(n14597) );
  AND U18971 ( .A(n14971), .B(n14972), .Z(n14969) );
  AND U18972 ( .A(a[39]), .B(b[48]), .Z(n14968) );
  XOR U18973 ( .A(n14974), .B(n14975), .Z(n14602) );
  AND U18974 ( .A(n14976), .B(n14977), .Z(n14974) );
  AND U18975 ( .A(a[40]), .B(b[47]), .Z(n14973) );
  XOR U18976 ( .A(n14979), .B(n14980), .Z(n14607) );
  AND U18977 ( .A(n14981), .B(n14982), .Z(n14979) );
  AND U18978 ( .A(a[41]), .B(b[46]), .Z(n14978) );
  XOR U18979 ( .A(n14984), .B(n14985), .Z(n14612) );
  AND U18980 ( .A(n14986), .B(n14987), .Z(n14984) );
  AND U18981 ( .A(a[42]), .B(b[45]), .Z(n14983) );
  XOR U18982 ( .A(n14989), .B(n14990), .Z(n14617) );
  AND U18983 ( .A(n14991), .B(n14992), .Z(n14989) );
  AND U18984 ( .A(a[43]), .B(b[44]), .Z(n14988) );
  XOR U18985 ( .A(n14994), .B(n14995), .Z(n14622) );
  AND U18986 ( .A(n14996), .B(n14997), .Z(n14994) );
  AND U18987 ( .A(b[43]), .B(a[44]), .Z(n14993) );
  XOR U18988 ( .A(n14999), .B(n15000), .Z(n14627) );
  AND U18989 ( .A(n15001), .B(n15002), .Z(n14999) );
  AND U18990 ( .A(b[42]), .B(a[45]), .Z(n14998) );
  XOR U18991 ( .A(n15004), .B(n15005), .Z(n14632) );
  AND U18992 ( .A(n15006), .B(n15007), .Z(n15004) );
  AND U18993 ( .A(b[41]), .B(a[46]), .Z(n15003) );
  XOR U18994 ( .A(n15009), .B(n15010), .Z(n14637) );
  AND U18995 ( .A(n15011), .B(n15012), .Z(n15009) );
  AND U18996 ( .A(b[40]), .B(a[47]), .Z(n15008) );
  XOR U18997 ( .A(n15014), .B(n15015), .Z(n14642) );
  AND U18998 ( .A(n15016), .B(n15017), .Z(n15014) );
  AND U18999 ( .A(b[39]), .B(a[48]), .Z(n15013) );
  XOR U19000 ( .A(n15019), .B(n15020), .Z(n14647) );
  AND U19001 ( .A(n15021), .B(n15022), .Z(n15019) );
  AND U19002 ( .A(b[38]), .B(a[49]), .Z(n15018) );
  XOR U19003 ( .A(n15024), .B(n15025), .Z(n14652) );
  AND U19004 ( .A(n15026), .B(n15027), .Z(n15024) );
  AND U19005 ( .A(b[37]), .B(a[50]), .Z(n15023) );
  XOR U19006 ( .A(n15029), .B(n15030), .Z(n14657) );
  AND U19007 ( .A(n15031), .B(n15032), .Z(n15029) );
  AND U19008 ( .A(b[36]), .B(a[51]), .Z(n15028) );
  XOR U19009 ( .A(n15034), .B(n15035), .Z(n14662) );
  AND U19010 ( .A(n15036), .B(n15037), .Z(n15034) );
  AND U19011 ( .A(b[35]), .B(a[52]), .Z(n15033) );
  XOR U19012 ( .A(n15039), .B(n15040), .Z(n14667) );
  AND U19013 ( .A(n15041), .B(n15042), .Z(n15039) );
  AND U19014 ( .A(b[34]), .B(a[53]), .Z(n15038) );
  XOR U19015 ( .A(n15044), .B(n15045), .Z(n14672) );
  AND U19016 ( .A(n15046), .B(n15047), .Z(n15044) );
  AND U19017 ( .A(b[33]), .B(a[54]), .Z(n15043) );
  XOR U19018 ( .A(n15049), .B(n15050), .Z(n14677) );
  AND U19019 ( .A(n15051), .B(n15052), .Z(n15049) );
  AND U19020 ( .A(b[32]), .B(a[55]), .Z(n15048) );
  XOR U19021 ( .A(n15054), .B(n15055), .Z(n14682) );
  AND U19022 ( .A(n15056), .B(n15057), .Z(n15054) );
  AND U19023 ( .A(b[31]), .B(a[56]), .Z(n15053) );
  XOR U19024 ( .A(n15059), .B(n15060), .Z(n14687) );
  AND U19025 ( .A(n15061), .B(n15062), .Z(n15059) );
  AND U19026 ( .A(b[30]), .B(a[57]), .Z(n15058) );
  XOR U19027 ( .A(n15064), .B(n15065), .Z(n14692) );
  AND U19028 ( .A(n15066), .B(n15067), .Z(n15064) );
  AND U19029 ( .A(b[29]), .B(a[58]), .Z(n15063) );
  XOR U19030 ( .A(n15069), .B(n15070), .Z(n14697) );
  AND U19031 ( .A(n15071), .B(n15072), .Z(n15069) );
  AND U19032 ( .A(b[28]), .B(a[59]), .Z(n15068) );
  XOR U19033 ( .A(n15074), .B(n15075), .Z(n14702) );
  AND U19034 ( .A(n15076), .B(n15077), .Z(n15074) );
  AND U19035 ( .A(b[27]), .B(a[60]), .Z(n15073) );
  XOR U19036 ( .A(n15079), .B(n15080), .Z(n14707) );
  AND U19037 ( .A(n15081), .B(n15082), .Z(n15079) );
  AND U19038 ( .A(b[26]), .B(a[61]), .Z(n15078) );
  XOR U19039 ( .A(n15084), .B(n15085), .Z(n14712) );
  AND U19040 ( .A(n15086), .B(n15087), .Z(n15084) );
  AND U19041 ( .A(b[25]), .B(a[62]), .Z(n15083) );
  XOR U19042 ( .A(n15089), .B(n15090), .Z(n14717) );
  AND U19043 ( .A(n15091), .B(n15092), .Z(n15089) );
  AND U19044 ( .A(b[24]), .B(a[63]), .Z(n15088) );
  XOR U19045 ( .A(n15094), .B(n15095), .Z(n14722) );
  AND U19046 ( .A(n15096), .B(n15097), .Z(n15094) );
  AND U19047 ( .A(b[23]), .B(a[64]), .Z(n15093) );
  XOR U19048 ( .A(n15099), .B(n15100), .Z(n14727) );
  AND U19049 ( .A(n15101), .B(n15102), .Z(n15099) );
  AND U19050 ( .A(b[22]), .B(a[65]), .Z(n15098) );
  XOR U19051 ( .A(n15104), .B(n15105), .Z(n14732) );
  AND U19052 ( .A(n15106), .B(n15107), .Z(n15104) );
  AND U19053 ( .A(b[21]), .B(a[66]), .Z(n15103) );
  XOR U19054 ( .A(n15109), .B(n15110), .Z(n14737) );
  AND U19055 ( .A(n15111), .B(n15112), .Z(n15109) );
  AND U19056 ( .A(b[20]), .B(a[67]), .Z(n15108) );
  XOR U19057 ( .A(n15114), .B(n15115), .Z(n14742) );
  AND U19058 ( .A(n15116), .B(n15117), .Z(n15114) );
  AND U19059 ( .A(b[19]), .B(a[68]), .Z(n15113) );
  XOR U19060 ( .A(n15119), .B(n15120), .Z(n14747) );
  AND U19061 ( .A(n15121), .B(n15122), .Z(n15119) );
  AND U19062 ( .A(b[18]), .B(a[69]), .Z(n15118) );
  XOR U19063 ( .A(n15124), .B(n15125), .Z(n14752) );
  AND U19064 ( .A(n15126), .B(n15127), .Z(n15124) );
  AND U19065 ( .A(b[17]), .B(a[70]), .Z(n15123) );
  XOR U19066 ( .A(n15129), .B(n15130), .Z(n14757) );
  AND U19067 ( .A(n15131), .B(n15132), .Z(n15129) );
  AND U19068 ( .A(b[16]), .B(a[71]), .Z(n15128) );
  XOR U19069 ( .A(n15134), .B(n15135), .Z(n14762) );
  AND U19070 ( .A(n15136), .B(n15137), .Z(n15134) );
  AND U19071 ( .A(b[15]), .B(a[72]), .Z(n15133) );
  XOR U19072 ( .A(n15139), .B(n15140), .Z(n14767) );
  AND U19073 ( .A(n15141), .B(n15142), .Z(n15139) );
  AND U19074 ( .A(b[14]), .B(a[73]), .Z(n15138) );
  XOR U19075 ( .A(n15144), .B(n15145), .Z(n14772) );
  AND U19076 ( .A(n15146), .B(n15147), .Z(n15144) );
  AND U19077 ( .A(b[13]), .B(a[74]), .Z(n15143) );
  XOR U19078 ( .A(n15149), .B(n15150), .Z(n14777) );
  AND U19079 ( .A(n15151), .B(n15152), .Z(n15149) );
  AND U19080 ( .A(b[12]), .B(a[75]), .Z(n15148) );
  XOR U19081 ( .A(n15154), .B(n15155), .Z(n14782) );
  AND U19082 ( .A(n15156), .B(n15157), .Z(n15154) );
  AND U19083 ( .A(b[11]), .B(a[76]), .Z(n15153) );
  XOR U19084 ( .A(n15159), .B(n15160), .Z(n14787) );
  AND U19085 ( .A(n15161), .B(n15162), .Z(n15159) );
  AND U19086 ( .A(b[10]), .B(a[77]), .Z(n15158) );
  XOR U19087 ( .A(n15164), .B(n15165), .Z(n14792) );
  AND U19088 ( .A(n15166), .B(n15167), .Z(n15164) );
  AND U19089 ( .A(b[9]), .B(a[78]), .Z(n15163) );
  XOR U19090 ( .A(n15169), .B(n15170), .Z(n14797) );
  AND U19091 ( .A(n15171), .B(n15172), .Z(n15169) );
  AND U19092 ( .A(b[8]), .B(a[79]), .Z(n15168) );
  XOR U19093 ( .A(n15174), .B(n15175), .Z(n14802) );
  AND U19094 ( .A(n15176), .B(n15177), .Z(n15174) );
  AND U19095 ( .A(b[7]), .B(a[80]), .Z(n15173) );
  XOR U19096 ( .A(n15179), .B(n15180), .Z(n14807) );
  AND U19097 ( .A(n15181), .B(n15182), .Z(n15179) );
  AND U19098 ( .A(b[6]), .B(a[81]), .Z(n15178) );
  XOR U19099 ( .A(n15184), .B(n15185), .Z(n14812) );
  AND U19100 ( .A(n15186), .B(n15187), .Z(n15184) );
  AND U19101 ( .A(b[5]), .B(a[82]), .Z(n15183) );
  XOR U19102 ( .A(n15189), .B(n15190), .Z(n14817) );
  AND U19103 ( .A(n15191), .B(n15192), .Z(n15189) );
  AND U19104 ( .A(b[4]), .B(a[83]), .Z(n15188) );
  XOR U19105 ( .A(n15194), .B(n15195), .Z(n14822) );
  AND U19106 ( .A(n15196), .B(n15197), .Z(n15194) );
  AND U19107 ( .A(b[3]), .B(a[84]), .Z(n15193) );
  XOR U19108 ( .A(n15199), .B(n15200), .Z(n14827) );
  OR U19109 ( .A(n15201), .B(n15202), .Z(n15200) );
  AND U19110 ( .A(b[2]), .B(a[85]), .Z(n15198) );
  XNOR U19111 ( .A(n14837), .B(n15203), .Z(n14833) );
  NAND U19112 ( .A(b[1]), .B(a[86]), .Z(n15203) );
  IV U19113 ( .A(n14831), .Z(n14837) );
  ANDN U19114 ( .B(n10293), .A(n10295), .Z(n14831) );
  NAND U19115 ( .A(a[86]), .B(b[0]), .Z(n10295) );
  XOR U19116 ( .A(n15201), .B(n15202), .Z(n10293) );
  XOR U19117 ( .A(n15205), .B(n15196), .Z(n15204) );
  XOR U19118 ( .A(n15191), .B(n15195), .Z(n15206) );
  XOR U19119 ( .A(n15186), .B(n15190), .Z(n15207) );
  XOR U19120 ( .A(n15181), .B(n15185), .Z(n15208) );
  XOR U19121 ( .A(n15176), .B(n15180), .Z(n15209) );
  XOR U19122 ( .A(n15171), .B(n15175), .Z(n15210) );
  XOR U19123 ( .A(n15166), .B(n15170), .Z(n15211) );
  XOR U19124 ( .A(n15161), .B(n15165), .Z(n15212) );
  XOR U19125 ( .A(n15156), .B(n15160), .Z(n15213) );
  XOR U19126 ( .A(n15151), .B(n15155), .Z(n15214) );
  XOR U19127 ( .A(n15146), .B(n15150), .Z(n15215) );
  XOR U19128 ( .A(n15141), .B(n15145), .Z(n15216) );
  XOR U19129 ( .A(n15136), .B(n15140), .Z(n15217) );
  XOR U19130 ( .A(n15131), .B(n15135), .Z(n15218) );
  XOR U19131 ( .A(n15126), .B(n15130), .Z(n15219) );
  XOR U19132 ( .A(n15121), .B(n15125), .Z(n15220) );
  XOR U19133 ( .A(n15116), .B(n15120), .Z(n15221) );
  XOR U19134 ( .A(n15111), .B(n15115), .Z(n15222) );
  XOR U19135 ( .A(n15106), .B(n15110), .Z(n15223) );
  XOR U19136 ( .A(n15101), .B(n15105), .Z(n15224) );
  XOR U19137 ( .A(n15096), .B(n15100), .Z(n15225) );
  XOR U19138 ( .A(n15091), .B(n15095), .Z(n15226) );
  XOR U19139 ( .A(n15086), .B(n15090), .Z(n15227) );
  XOR U19140 ( .A(n15081), .B(n15085), .Z(n15228) );
  XOR U19141 ( .A(n15076), .B(n15080), .Z(n15229) );
  XOR U19142 ( .A(n15071), .B(n15075), .Z(n15230) );
  XOR U19143 ( .A(n15066), .B(n15070), .Z(n15231) );
  XOR U19144 ( .A(n15061), .B(n15065), .Z(n15232) );
  XOR U19145 ( .A(n15056), .B(n15060), .Z(n15233) );
  XOR U19146 ( .A(n15051), .B(n15055), .Z(n15234) );
  XOR U19147 ( .A(n15046), .B(n15050), .Z(n15235) );
  XOR U19148 ( .A(n15041), .B(n15045), .Z(n15236) );
  XOR U19149 ( .A(n15036), .B(n15040), .Z(n15237) );
  XOR U19150 ( .A(n15031), .B(n15035), .Z(n15238) );
  XOR U19151 ( .A(n15026), .B(n15030), .Z(n15239) );
  XOR U19152 ( .A(n15021), .B(n15025), .Z(n15240) );
  XOR U19153 ( .A(n15016), .B(n15020), .Z(n15241) );
  XOR U19154 ( .A(n15011), .B(n15015), .Z(n15242) );
  XOR U19155 ( .A(n15006), .B(n15010), .Z(n15243) );
  XOR U19156 ( .A(n15001), .B(n15005), .Z(n15244) );
  XOR U19157 ( .A(n14996), .B(n15000), .Z(n15245) );
  XOR U19158 ( .A(n14991), .B(n14995), .Z(n15246) );
  XOR U19159 ( .A(n14986), .B(n14990), .Z(n15247) );
  XOR U19160 ( .A(n14981), .B(n14985), .Z(n15248) );
  XOR U19161 ( .A(n14976), .B(n14980), .Z(n15249) );
  XOR U19162 ( .A(n14971), .B(n14975), .Z(n15250) );
  XOR U19163 ( .A(n14966), .B(n14970), .Z(n15251) );
  XOR U19164 ( .A(n14961), .B(n14965), .Z(n15252) );
  XOR U19165 ( .A(n14951), .B(n14960), .Z(n15253) );
  XOR U19166 ( .A(n15254), .B(n14950), .Z(n14951) );
  AND U19167 ( .A(a[36]), .B(b[50]), .Z(n15254) );
  XNOR U19168 ( .A(n14950), .B(n14956), .Z(n15255) );
  XNOR U19169 ( .A(n14955), .B(n14947), .Z(n15256) );
  XNOR U19170 ( .A(n14946), .B(n14942), .Z(n15257) );
  XNOR U19171 ( .A(n14941), .B(n14937), .Z(n15258) );
  XNOR U19172 ( .A(n14936), .B(n14932), .Z(n15259) );
  XNOR U19173 ( .A(n14931), .B(n14927), .Z(n15260) );
  XNOR U19174 ( .A(n14926), .B(n14922), .Z(n15261) );
  XNOR U19175 ( .A(n14921), .B(n14917), .Z(n15262) );
  XNOR U19176 ( .A(n14916), .B(n14912), .Z(n15263) );
  XOR U19177 ( .A(n14911), .B(n14908), .Z(n15264) );
  XOR U19178 ( .A(n15265), .B(n15266), .Z(n14908) );
  XOR U19179 ( .A(n14906), .B(n15267), .Z(n15266) );
  XOR U19180 ( .A(n15268), .B(n15269), .Z(n15267) );
  XOR U19181 ( .A(n15270), .B(n15271), .Z(n15269) );
  NAND U19182 ( .A(a[24]), .B(b[62]), .Z(n15271) );
  AND U19183 ( .A(a[23]), .B(b[63]), .Z(n15270) );
  XOR U19184 ( .A(n15272), .B(n15268), .Z(n15265) );
  XOR U19185 ( .A(n15273), .B(n15274), .Z(n15268) );
  ANDN U19186 ( .B(n15275), .A(n15276), .Z(n15273) );
  AND U19187 ( .A(a[25]), .B(b[61]), .Z(n15272) );
  XOR U19188 ( .A(n15277), .B(n14906), .Z(n14907) );
  XOR U19189 ( .A(n15278), .B(n15279), .Z(n14906) );
  AND U19190 ( .A(n15280), .B(n15281), .Z(n15278) );
  AND U19191 ( .A(a[26]), .B(b[60]), .Z(n15277) );
  XOR U19192 ( .A(n15282), .B(n14911), .Z(n14913) );
  XOR U19193 ( .A(n15283), .B(n15284), .Z(n14911) );
  AND U19194 ( .A(n15285), .B(n15286), .Z(n15283) );
  AND U19195 ( .A(a[27]), .B(b[59]), .Z(n15282) );
  XOR U19196 ( .A(n15287), .B(n14916), .Z(n14918) );
  XOR U19197 ( .A(n15288), .B(n15289), .Z(n14916) );
  AND U19198 ( .A(n15290), .B(n15291), .Z(n15288) );
  AND U19199 ( .A(a[28]), .B(b[58]), .Z(n15287) );
  XOR U19200 ( .A(n15292), .B(n14921), .Z(n14923) );
  XOR U19201 ( .A(n15293), .B(n15294), .Z(n14921) );
  AND U19202 ( .A(n15295), .B(n15296), .Z(n15293) );
  AND U19203 ( .A(a[29]), .B(b[57]), .Z(n15292) );
  XOR U19204 ( .A(n15297), .B(n14926), .Z(n14928) );
  XOR U19205 ( .A(n15298), .B(n15299), .Z(n14926) );
  AND U19206 ( .A(n15300), .B(n15301), .Z(n15298) );
  AND U19207 ( .A(a[30]), .B(b[56]), .Z(n15297) );
  XOR U19208 ( .A(n15302), .B(n14931), .Z(n14933) );
  XOR U19209 ( .A(n15303), .B(n15304), .Z(n14931) );
  AND U19210 ( .A(n15305), .B(n15306), .Z(n15303) );
  AND U19211 ( .A(a[31]), .B(b[55]), .Z(n15302) );
  XOR U19212 ( .A(n15307), .B(n14936), .Z(n14938) );
  XOR U19213 ( .A(n15308), .B(n15309), .Z(n14936) );
  AND U19214 ( .A(n15310), .B(n15311), .Z(n15308) );
  AND U19215 ( .A(a[32]), .B(b[54]), .Z(n15307) );
  XOR U19216 ( .A(n15312), .B(n14941), .Z(n14943) );
  XOR U19217 ( .A(n15313), .B(n15314), .Z(n14941) );
  AND U19218 ( .A(n15315), .B(n15316), .Z(n15313) );
  AND U19219 ( .A(a[33]), .B(b[53]), .Z(n15312) );
  XOR U19220 ( .A(n15317), .B(n14946), .Z(n14948) );
  XOR U19221 ( .A(n15318), .B(n15319), .Z(n14946) );
  AND U19222 ( .A(n15320), .B(n15321), .Z(n15318) );
  AND U19223 ( .A(a[34]), .B(b[52]), .Z(n15317) );
  XOR U19224 ( .A(n15322), .B(n15323), .Z(n14950) );
  AND U19225 ( .A(n15324), .B(n15325), .Z(n15322) );
  XOR U19226 ( .A(n15326), .B(n14955), .Z(n14957) );
  XOR U19227 ( .A(n15327), .B(n15328), .Z(n14955) );
  AND U19228 ( .A(n15329), .B(n15330), .Z(n15327) );
  AND U19229 ( .A(a[35]), .B(b[51]), .Z(n15326) );
  XOR U19230 ( .A(n15332), .B(n15333), .Z(n14960) );
  AND U19231 ( .A(n15334), .B(n15335), .Z(n15332) );
  AND U19232 ( .A(a[37]), .B(b[49]), .Z(n15331) );
  XOR U19233 ( .A(n15337), .B(n15338), .Z(n14965) );
  AND U19234 ( .A(n15339), .B(n15340), .Z(n15337) );
  AND U19235 ( .A(a[38]), .B(b[48]), .Z(n15336) );
  XOR U19236 ( .A(n15342), .B(n15343), .Z(n14970) );
  AND U19237 ( .A(n15344), .B(n15345), .Z(n15342) );
  AND U19238 ( .A(a[39]), .B(b[47]), .Z(n15341) );
  XOR U19239 ( .A(n15347), .B(n15348), .Z(n14975) );
  AND U19240 ( .A(n15349), .B(n15350), .Z(n15347) );
  AND U19241 ( .A(a[40]), .B(b[46]), .Z(n15346) );
  XOR U19242 ( .A(n15352), .B(n15353), .Z(n14980) );
  AND U19243 ( .A(n15354), .B(n15355), .Z(n15352) );
  AND U19244 ( .A(a[41]), .B(b[45]), .Z(n15351) );
  XOR U19245 ( .A(n15357), .B(n15358), .Z(n14985) );
  AND U19246 ( .A(n15359), .B(n15360), .Z(n15357) );
  AND U19247 ( .A(a[42]), .B(b[44]), .Z(n15356) );
  XOR U19248 ( .A(n15362), .B(n15363), .Z(n14990) );
  AND U19249 ( .A(n15364), .B(n15365), .Z(n15362) );
  AND U19250 ( .A(a[43]), .B(b[43]), .Z(n15361) );
  XOR U19251 ( .A(n15367), .B(n15368), .Z(n14995) );
  AND U19252 ( .A(n15369), .B(n15370), .Z(n15367) );
  AND U19253 ( .A(b[42]), .B(a[44]), .Z(n15366) );
  XOR U19254 ( .A(n15372), .B(n15373), .Z(n15000) );
  AND U19255 ( .A(n15374), .B(n15375), .Z(n15372) );
  AND U19256 ( .A(b[41]), .B(a[45]), .Z(n15371) );
  XOR U19257 ( .A(n15377), .B(n15378), .Z(n15005) );
  AND U19258 ( .A(n15379), .B(n15380), .Z(n15377) );
  AND U19259 ( .A(b[40]), .B(a[46]), .Z(n15376) );
  XOR U19260 ( .A(n15382), .B(n15383), .Z(n15010) );
  AND U19261 ( .A(n15384), .B(n15385), .Z(n15382) );
  AND U19262 ( .A(b[39]), .B(a[47]), .Z(n15381) );
  XOR U19263 ( .A(n15387), .B(n15388), .Z(n15015) );
  AND U19264 ( .A(n15389), .B(n15390), .Z(n15387) );
  AND U19265 ( .A(b[38]), .B(a[48]), .Z(n15386) );
  XOR U19266 ( .A(n15392), .B(n15393), .Z(n15020) );
  AND U19267 ( .A(n15394), .B(n15395), .Z(n15392) );
  AND U19268 ( .A(b[37]), .B(a[49]), .Z(n15391) );
  XOR U19269 ( .A(n15397), .B(n15398), .Z(n15025) );
  AND U19270 ( .A(n15399), .B(n15400), .Z(n15397) );
  AND U19271 ( .A(b[36]), .B(a[50]), .Z(n15396) );
  XOR U19272 ( .A(n15402), .B(n15403), .Z(n15030) );
  AND U19273 ( .A(n15404), .B(n15405), .Z(n15402) );
  AND U19274 ( .A(b[35]), .B(a[51]), .Z(n15401) );
  XOR U19275 ( .A(n15407), .B(n15408), .Z(n15035) );
  AND U19276 ( .A(n15409), .B(n15410), .Z(n15407) );
  AND U19277 ( .A(b[34]), .B(a[52]), .Z(n15406) );
  XOR U19278 ( .A(n15412), .B(n15413), .Z(n15040) );
  AND U19279 ( .A(n15414), .B(n15415), .Z(n15412) );
  AND U19280 ( .A(b[33]), .B(a[53]), .Z(n15411) );
  XOR U19281 ( .A(n15417), .B(n15418), .Z(n15045) );
  AND U19282 ( .A(n15419), .B(n15420), .Z(n15417) );
  AND U19283 ( .A(b[32]), .B(a[54]), .Z(n15416) );
  XOR U19284 ( .A(n15422), .B(n15423), .Z(n15050) );
  AND U19285 ( .A(n15424), .B(n15425), .Z(n15422) );
  AND U19286 ( .A(b[31]), .B(a[55]), .Z(n15421) );
  XOR U19287 ( .A(n15427), .B(n15428), .Z(n15055) );
  AND U19288 ( .A(n15429), .B(n15430), .Z(n15427) );
  AND U19289 ( .A(b[30]), .B(a[56]), .Z(n15426) );
  XOR U19290 ( .A(n15432), .B(n15433), .Z(n15060) );
  AND U19291 ( .A(n15434), .B(n15435), .Z(n15432) );
  AND U19292 ( .A(b[29]), .B(a[57]), .Z(n15431) );
  XOR U19293 ( .A(n15437), .B(n15438), .Z(n15065) );
  AND U19294 ( .A(n15439), .B(n15440), .Z(n15437) );
  AND U19295 ( .A(b[28]), .B(a[58]), .Z(n15436) );
  XOR U19296 ( .A(n15442), .B(n15443), .Z(n15070) );
  AND U19297 ( .A(n15444), .B(n15445), .Z(n15442) );
  AND U19298 ( .A(b[27]), .B(a[59]), .Z(n15441) );
  XOR U19299 ( .A(n15447), .B(n15448), .Z(n15075) );
  AND U19300 ( .A(n15449), .B(n15450), .Z(n15447) );
  AND U19301 ( .A(b[26]), .B(a[60]), .Z(n15446) );
  XOR U19302 ( .A(n15452), .B(n15453), .Z(n15080) );
  AND U19303 ( .A(n15454), .B(n15455), .Z(n15452) );
  AND U19304 ( .A(b[25]), .B(a[61]), .Z(n15451) );
  XOR U19305 ( .A(n15457), .B(n15458), .Z(n15085) );
  AND U19306 ( .A(n15459), .B(n15460), .Z(n15457) );
  AND U19307 ( .A(b[24]), .B(a[62]), .Z(n15456) );
  XOR U19308 ( .A(n15462), .B(n15463), .Z(n15090) );
  AND U19309 ( .A(n15464), .B(n15465), .Z(n15462) );
  AND U19310 ( .A(b[23]), .B(a[63]), .Z(n15461) );
  XOR U19311 ( .A(n15467), .B(n15468), .Z(n15095) );
  AND U19312 ( .A(n15469), .B(n15470), .Z(n15467) );
  AND U19313 ( .A(b[22]), .B(a[64]), .Z(n15466) );
  XOR U19314 ( .A(n15472), .B(n15473), .Z(n15100) );
  AND U19315 ( .A(n15474), .B(n15475), .Z(n15472) );
  AND U19316 ( .A(b[21]), .B(a[65]), .Z(n15471) );
  XOR U19317 ( .A(n15477), .B(n15478), .Z(n15105) );
  AND U19318 ( .A(n15479), .B(n15480), .Z(n15477) );
  AND U19319 ( .A(b[20]), .B(a[66]), .Z(n15476) );
  XOR U19320 ( .A(n15482), .B(n15483), .Z(n15110) );
  AND U19321 ( .A(n15484), .B(n15485), .Z(n15482) );
  AND U19322 ( .A(b[19]), .B(a[67]), .Z(n15481) );
  XOR U19323 ( .A(n15487), .B(n15488), .Z(n15115) );
  AND U19324 ( .A(n15489), .B(n15490), .Z(n15487) );
  AND U19325 ( .A(b[18]), .B(a[68]), .Z(n15486) );
  XOR U19326 ( .A(n15492), .B(n15493), .Z(n15120) );
  AND U19327 ( .A(n15494), .B(n15495), .Z(n15492) );
  AND U19328 ( .A(b[17]), .B(a[69]), .Z(n15491) );
  XOR U19329 ( .A(n15497), .B(n15498), .Z(n15125) );
  AND U19330 ( .A(n15499), .B(n15500), .Z(n15497) );
  AND U19331 ( .A(b[16]), .B(a[70]), .Z(n15496) );
  XOR U19332 ( .A(n15502), .B(n15503), .Z(n15130) );
  AND U19333 ( .A(n15504), .B(n15505), .Z(n15502) );
  AND U19334 ( .A(b[15]), .B(a[71]), .Z(n15501) );
  XOR U19335 ( .A(n15507), .B(n15508), .Z(n15135) );
  AND U19336 ( .A(n15509), .B(n15510), .Z(n15507) );
  AND U19337 ( .A(b[14]), .B(a[72]), .Z(n15506) );
  XOR U19338 ( .A(n15512), .B(n15513), .Z(n15140) );
  AND U19339 ( .A(n15514), .B(n15515), .Z(n15512) );
  AND U19340 ( .A(b[13]), .B(a[73]), .Z(n15511) );
  XOR U19341 ( .A(n15517), .B(n15518), .Z(n15145) );
  AND U19342 ( .A(n15519), .B(n15520), .Z(n15517) );
  AND U19343 ( .A(b[12]), .B(a[74]), .Z(n15516) );
  XOR U19344 ( .A(n15522), .B(n15523), .Z(n15150) );
  AND U19345 ( .A(n15524), .B(n15525), .Z(n15522) );
  AND U19346 ( .A(b[11]), .B(a[75]), .Z(n15521) );
  XOR U19347 ( .A(n15527), .B(n15528), .Z(n15155) );
  AND U19348 ( .A(n15529), .B(n15530), .Z(n15527) );
  AND U19349 ( .A(b[10]), .B(a[76]), .Z(n15526) );
  XOR U19350 ( .A(n15532), .B(n15533), .Z(n15160) );
  AND U19351 ( .A(n15534), .B(n15535), .Z(n15532) );
  AND U19352 ( .A(b[9]), .B(a[77]), .Z(n15531) );
  XOR U19353 ( .A(n15537), .B(n15538), .Z(n15165) );
  AND U19354 ( .A(n15539), .B(n15540), .Z(n15537) );
  AND U19355 ( .A(b[8]), .B(a[78]), .Z(n15536) );
  XOR U19356 ( .A(n15542), .B(n15543), .Z(n15170) );
  AND U19357 ( .A(n15544), .B(n15545), .Z(n15542) );
  AND U19358 ( .A(b[7]), .B(a[79]), .Z(n15541) );
  XOR U19359 ( .A(n15547), .B(n15548), .Z(n15175) );
  AND U19360 ( .A(n15549), .B(n15550), .Z(n15547) );
  AND U19361 ( .A(b[6]), .B(a[80]), .Z(n15546) );
  XOR U19362 ( .A(n15552), .B(n15553), .Z(n15180) );
  AND U19363 ( .A(n15554), .B(n15555), .Z(n15552) );
  AND U19364 ( .A(b[5]), .B(a[81]), .Z(n15551) );
  XOR U19365 ( .A(n15557), .B(n15558), .Z(n15185) );
  AND U19366 ( .A(n15559), .B(n15560), .Z(n15557) );
  AND U19367 ( .A(b[4]), .B(a[82]), .Z(n15556) );
  XOR U19368 ( .A(n15562), .B(n15563), .Z(n15190) );
  AND U19369 ( .A(n15564), .B(n15565), .Z(n15562) );
  AND U19370 ( .A(b[3]), .B(a[83]), .Z(n15561) );
  XOR U19371 ( .A(n15567), .B(n15568), .Z(n15195) );
  OR U19372 ( .A(n15569), .B(n15570), .Z(n15568) );
  AND U19373 ( .A(b[2]), .B(a[84]), .Z(n15566) );
  XNOR U19374 ( .A(n15205), .B(n15571), .Z(n15201) );
  NAND U19375 ( .A(b[1]), .B(a[85]), .Z(n15571) );
  IV U19376 ( .A(n15199), .Z(n15205) );
  ANDN U19377 ( .B(n10296), .A(n10298), .Z(n15199) );
  NAND U19378 ( .A(a[85]), .B(b[0]), .Z(n10298) );
  XOR U19379 ( .A(n15569), .B(n15570), .Z(n10296) );
  XOR U19380 ( .A(n15573), .B(n15564), .Z(n15572) );
  XOR U19381 ( .A(n15559), .B(n15563), .Z(n15574) );
  XOR U19382 ( .A(n15554), .B(n15558), .Z(n15575) );
  XOR U19383 ( .A(n15549), .B(n15553), .Z(n15576) );
  XOR U19384 ( .A(n15544), .B(n15548), .Z(n15577) );
  XOR U19385 ( .A(n15539), .B(n15543), .Z(n15578) );
  XOR U19386 ( .A(n15534), .B(n15538), .Z(n15579) );
  XOR U19387 ( .A(n15529), .B(n15533), .Z(n15580) );
  XOR U19388 ( .A(n15524), .B(n15528), .Z(n15581) );
  XOR U19389 ( .A(n15519), .B(n15523), .Z(n15582) );
  XOR U19390 ( .A(n15514), .B(n15518), .Z(n15583) );
  XOR U19391 ( .A(n15509), .B(n15513), .Z(n15584) );
  XOR U19392 ( .A(n15504), .B(n15508), .Z(n15585) );
  XOR U19393 ( .A(n15499), .B(n15503), .Z(n15586) );
  XOR U19394 ( .A(n15494), .B(n15498), .Z(n15587) );
  XOR U19395 ( .A(n15489), .B(n15493), .Z(n15588) );
  XOR U19396 ( .A(n15484), .B(n15488), .Z(n15589) );
  XOR U19397 ( .A(n15479), .B(n15483), .Z(n15590) );
  XOR U19398 ( .A(n15474), .B(n15478), .Z(n15591) );
  XOR U19399 ( .A(n15469), .B(n15473), .Z(n15592) );
  XOR U19400 ( .A(n15464), .B(n15468), .Z(n15593) );
  XOR U19401 ( .A(n15459), .B(n15463), .Z(n15594) );
  XOR U19402 ( .A(n15454), .B(n15458), .Z(n15595) );
  XOR U19403 ( .A(n15449), .B(n15453), .Z(n15596) );
  XOR U19404 ( .A(n15444), .B(n15448), .Z(n15597) );
  XOR U19405 ( .A(n15439), .B(n15443), .Z(n15598) );
  XOR U19406 ( .A(n15434), .B(n15438), .Z(n15599) );
  XOR U19407 ( .A(n15429), .B(n15433), .Z(n15600) );
  XOR U19408 ( .A(n15424), .B(n15428), .Z(n15601) );
  XOR U19409 ( .A(n15419), .B(n15423), .Z(n15602) );
  XOR U19410 ( .A(n15414), .B(n15418), .Z(n15603) );
  XOR U19411 ( .A(n15409), .B(n15413), .Z(n15604) );
  XOR U19412 ( .A(n15404), .B(n15408), .Z(n15605) );
  XOR U19413 ( .A(n15399), .B(n15403), .Z(n15606) );
  XOR U19414 ( .A(n15394), .B(n15398), .Z(n15607) );
  XOR U19415 ( .A(n15389), .B(n15393), .Z(n15608) );
  XOR U19416 ( .A(n15384), .B(n15388), .Z(n15609) );
  XOR U19417 ( .A(n15379), .B(n15383), .Z(n15610) );
  XOR U19418 ( .A(n15374), .B(n15378), .Z(n15611) );
  XOR U19419 ( .A(n15369), .B(n15373), .Z(n15612) );
  XOR U19420 ( .A(n15364), .B(n15368), .Z(n15613) );
  XOR U19421 ( .A(n15359), .B(n15363), .Z(n15614) );
  XOR U19422 ( .A(n15354), .B(n15358), .Z(n15615) );
  XOR U19423 ( .A(n15349), .B(n15353), .Z(n15616) );
  XOR U19424 ( .A(n15344), .B(n15348), .Z(n15617) );
  XOR U19425 ( .A(n15339), .B(n15343), .Z(n15618) );
  XOR U19426 ( .A(n15334), .B(n15338), .Z(n15619) );
  XOR U19427 ( .A(n15324), .B(n15333), .Z(n15620) );
  XOR U19428 ( .A(n15621), .B(n15323), .Z(n15324) );
  AND U19429 ( .A(a[36]), .B(b[49]), .Z(n15621) );
  XNOR U19430 ( .A(n15323), .B(n15329), .Z(n15622) );
  XNOR U19431 ( .A(n15328), .B(n15320), .Z(n15623) );
  XNOR U19432 ( .A(n15319), .B(n15315), .Z(n15624) );
  XNOR U19433 ( .A(n15314), .B(n15310), .Z(n15625) );
  XNOR U19434 ( .A(n15309), .B(n15305), .Z(n15626) );
  XNOR U19435 ( .A(n15304), .B(n15300), .Z(n15627) );
  XNOR U19436 ( .A(n15299), .B(n15295), .Z(n15628) );
  XNOR U19437 ( .A(n15294), .B(n15290), .Z(n15629) );
  XNOR U19438 ( .A(n15289), .B(n15285), .Z(n15630) );
  XNOR U19439 ( .A(n15284), .B(n15280), .Z(n15631) );
  XOR U19440 ( .A(n15279), .B(n15276), .Z(n15632) );
  XOR U19441 ( .A(n15633), .B(n15634), .Z(n15276) );
  XOR U19442 ( .A(n15274), .B(n15635), .Z(n15634) );
  XOR U19443 ( .A(n15636), .B(n15637), .Z(n15635) );
  XOR U19444 ( .A(n15638), .B(n15639), .Z(n15637) );
  NAND U19445 ( .A(a[23]), .B(b[62]), .Z(n15639) );
  AND U19446 ( .A(a[22]), .B(b[63]), .Z(n15638) );
  XOR U19447 ( .A(n15640), .B(n15636), .Z(n15633) );
  XOR U19448 ( .A(n15641), .B(n15642), .Z(n15636) );
  ANDN U19449 ( .B(n15643), .A(n15644), .Z(n15641) );
  AND U19450 ( .A(a[24]), .B(b[61]), .Z(n15640) );
  XOR U19451 ( .A(n15645), .B(n15274), .Z(n15275) );
  XOR U19452 ( .A(n15646), .B(n15647), .Z(n15274) );
  AND U19453 ( .A(n15648), .B(n15649), .Z(n15646) );
  AND U19454 ( .A(a[25]), .B(b[60]), .Z(n15645) );
  XOR U19455 ( .A(n15650), .B(n15279), .Z(n15281) );
  XOR U19456 ( .A(n15651), .B(n15652), .Z(n15279) );
  AND U19457 ( .A(n15653), .B(n15654), .Z(n15651) );
  AND U19458 ( .A(a[26]), .B(b[59]), .Z(n15650) );
  XOR U19459 ( .A(n15655), .B(n15284), .Z(n15286) );
  XOR U19460 ( .A(n15656), .B(n15657), .Z(n15284) );
  AND U19461 ( .A(n15658), .B(n15659), .Z(n15656) );
  AND U19462 ( .A(a[27]), .B(b[58]), .Z(n15655) );
  XOR U19463 ( .A(n15660), .B(n15289), .Z(n15291) );
  XOR U19464 ( .A(n15661), .B(n15662), .Z(n15289) );
  AND U19465 ( .A(n15663), .B(n15664), .Z(n15661) );
  AND U19466 ( .A(a[28]), .B(b[57]), .Z(n15660) );
  XOR U19467 ( .A(n15665), .B(n15294), .Z(n15296) );
  XOR U19468 ( .A(n15666), .B(n15667), .Z(n15294) );
  AND U19469 ( .A(n15668), .B(n15669), .Z(n15666) );
  AND U19470 ( .A(a[29]), .B(b[56]), .Z(n15665) );
  XOR U19471 ( .A(n15670), .B(n15299), .Z(n15301) );
  XOR U19472 ( .A(n15671), .B(n15672), .Z(n15299) );
  AND U19473 ( .A(n15673), .B(n15674), .Z(n15671) );
  AND U19474 ( .A(a[30]), .B(b[55]), .Z(n15670) );
  XOR U19475 ( .A(n15675), .B(n15304), .Z(n15306) );
  XOR U19476 ( .A(n15676), .B(n15677), .Z(n15304) );
  AND U19477 ( .A(n15678), .B(n15679), .Z(n15676) );
  AND U19478 ( .A(a[31]), .B(b[54]), .Z(n15675) );
  XOR U19479 ( .A(n15680), .B(n15309), .Z(n15311) );
  XOR U19480 ( .A(n15681), .B(n15682), .Z(n15309) );
  AND U19481 ( .A(n15683), .B(n15684), .Z(n15681) );
  AND U19482 ( .A(a[32]), .B(b[53]), .Z(n15680) );
  XOR U19483 ( .A(n15685), .B(n15314), .Z(n15316) );
  XOR U19484 ( .A(n15686), .B(n15687), .Z(n15314) );
  AND U19485 ( .A(n15688), .B(n15689), .Z(n15686) );
  AND U19486 ( .A(a[33]), .B(b[52]), .Z(n15685) );
  XOR U19487 ( .A(n15690), .B(n15319), .Z(n15321) );
  XOR U19488 ( .A(n15691), .B(n15692), .Z(n15319) );
  AND U19489 ( .A(n15693), .B(n15694), .Z(n15691) );
  AND U19490 ( .A(a[34]), .B(b[51]), .Z(n15690) );
  XOR U19491 ( .A(n15695), .B(n15696), .Z(n15323) );
  AND U19492 ( .A(n15697), .B(n15698), .Z(n15695) );
  XOR U19493 ( .A(n15699), .B(n15328), .Z(n15330) );
  XOR U19494 ( .A(n15700), .B(n15701), .Z(n15328) );
  AND U19495 ( .A(n15702), .B(n15703), .Z(n15700) );
  AND U19496 ( .A(a[35]), .B(b[50]), .Z(n15699) );
  XOR U19497 ( .A(n15705), .B(n15706), .Z(n15333) );
  AND U19498 ( .A(n15707), .B(n15708), .Z(n15705) );
  AND U19499 ( .A(a[37]), .B(b[48]), .Z(n15704) );
  XOR U19500 ( .A(n15710), .B(n15711), .Z(n15338) );
  AND U19501 ( .A(n15712), .B(n15713), .Z(n15710) );
  AND U19502 ( .A(a[38]), .B(b[47]), .Z(n15709) );
  XOR U19503 ( .A(n15715), .B(n15716), .Z(n15343) );
  AND U19504 ( .A(n15717), .B(n15718), .Z(n15715) );
  AND U19505 ( .A(a[39]), .B(b[46]), .Z(n15714) );
  XOR U19506 ( .A(n15720), .B(n15721), .Z(n15348) );
  AND U19507 ( .A(n15722), .B(n15723), .Z(n15720) );
  AND U19508 ( .A(a[40]), .B(b[45]), .Z(n15719) );
  XOR U19509 ( .A(n15725), .B(n15726), .Z(n15353) );
  AND U19510 ( .A(n15727), .B(n15728), .Z(n15725) );
  AND U19511 ( .A(a[41]), .B(b[44]), .Z(n15724) );
  XOR U19512 ( .A(n15730), .B(n15731), .Z(n15358) );
  AND U19513 ( .A(n15732), .B(n15733), .Z(n15730) );
  AND U19514 ( .A(a[42]), .B(b[43]), .Z(n15729) );
  XOR U19515 ( .A(n15735), .B(n15736), .Z(n15363) );
  AND U19516 ( .A(n15737), .B(n15738), .Z(n15735) );
  AND U19517 ( .A(b[42]), .B(a[43]), .Z(n15734) );
  XOR U19518 ( .A(n15740), .B(n15741), .Z(n15368) );
  AND U19519 ( .A(n15742), .B(n15743), .Z(n15740) );
  AND U19520 ( .A(b[41]), .B(a[44]), .Z(n15739) );
  XOR U19521 ( .A(n15745), .B(n15746), .Z(n15373) );
  AND U19522 ( .A(n15747), .B(n15748), .Z(n15745) );
  AND U19523 ( .A(b[40]), .B(a[45]), .Z(n15744) );
  XOR U19524 ( .A(n15750), .B(n15751), .Z(n15378) );
  AND U19525 ( .A(n15752), .B(n15753), .Z(n15750) );
  AND U19526 ( .A(b[39]), .B(a[46]), .Z(n15749) );
  XOR U19527 ( .A(n15755), .B(n15756), .Z(n15383) );
  AND U19528 ( .A(n15757), .B(n15758), .Z(n15755) );
  AND U19529 ( .A(b[38]), .B(a[47]), .Z(n15754) );
  XOR U19530 ( .A(n15760), .B(n15761), .Z(n15388) );
  AND U19531 ( .A(n15762), .B(n15763), .Z(n15760) );
  AND U19532 ( .A(b[37]), .B(a[48]), .Z(n15759) );
  XOR U19533 ( .A(n15765), .B(n15766), .Z(n15393) );
  AND U19534 ( .A(n15767), .B(n15768), .Z(n15765) );
  AND U19535 ( .A(b[36]), .B(a[49]), .Z(n15764) );
  XOR U19536 ( .A(n15770), .B(n15771), .Z(n15398) );
  AND U19537 ( .A(n15772), .B(n15773), .Z(n15770) );
  AND U19538 ( .A(b[35]), .B(a[50]), .Z(n15769) );
  XOR U19539 ( .A(n15775), .B(n15776), .Z(n15403) );
  AND U19540 ( .A(n15777), .B(n15778), .Z(n15775) );
  AND U19541 ( .A(b[34]), .B(a[51]), .Z(n15774) );
  XOR U19542 ( .A(n15780), .B(n15781), .Z(n15408) );
  AND U19543 ( .A(n15782), .B(n15783), .Z(n15780) );
  AND U19544 ( .A(b[33]), .B(a[52]), .Z(n15779) );
  XOR U19545 ( .A(n15785), .B(n15786), .Z(n15413) );
  AND U19546 ( .A(n15787), .B(n15788), .Z(n15785) );
  AND U19547 ( .A(b[32]), .B(a[53]), .Z(n15784) );
  XOR U19548 ( .A(n15790), .B(n15791), .Z(n15418) );
  AND U19549 ( .A(n15792), .B(n15793), .Z(n15790) );
  AND U19550 ( .A(b[31]), .B(a[54]), .Z(n15789) );
  XOR U19551 ( .A(n15795), .B(n15796), .Z(n15423) );
  AND U19552 ( .A(n15797), .B(n15798), .Z(n15795) );
  AND U19553 ( .A(b[30]), .B(a[55]), .Z(n15794) );
  XOR U19554 ( .A(n15800), .B(n15801), .Z(n15428) );
  AND U19555 ( .A(n15802), .B(n15803), .Z(n15800) );
  AND U19556 ( .A(b[29]), .B(a[56]), .Z(n15799) );
  XOR U19557 ( .A(n15805), .B(n15806), .Z(n15433) );
  AND U19558 ( .A(n15807), .B(n15808), .Z(n15805) );
  AND U19559 ( .A(b[28]), .B(a[57]), .Z(n15804) );
  XOR U19560 ( .A(n15810), .B(n15811), .Z(n15438) );
  AND U19561 ( .A(n15812), .B(n15813), .Z(n15810) );
  AND U19562 ( .A(b[27]), .B(a[58]), .Z(n15809) );
  XOR U19563 ( .A(n15815), .B(n15816), .Z(n15443) );
  AND U19564 ( .A(n15817), .B(n15818), .Z(n15815) );
  AND U19565 ( .A(b[26]), .B(a[59]), .Z(n15814) );
  XOR U19566 ( .A(n15820), .B(n15821), .Z(n15448) );
  AND U19567 ( .A(n15822), .B(n15823), .Z(n15820) );
  AND U19568 ( .A(b[25]), .B(a[60]), .Z(n15819) );
  XOR U19569 ( .A(n15825), .B(n15826), .Z(n15453) );
  AND U19570 ( .A(n15827), .B(n15828), .Z(n15825) );
  AND U19571 ( .A(b[24]), .B(a[61]), .Z(n15824) );
  XOR U19572 ( .A(n15830), .B(n15831), .Z(n15458) );
  AND U19573 ( .A(n15832), .B(n15833), .Z(n15830) );
  AND U19574 ( .A(b[23]), .B(a[62]), .Z(n15829) );
  XOR U19575 ( .A(n15835), .B(n15836), .Z(n15463) );
  AND U19576 ( .A(n15837), .B(n15838), .Z(n15835) );
  AND U19577 ( .A(b[22]), .B(a[63]), .Z(n15834) );
  XOR U19578 ( .A(n15840), .B(n15841), .Z(n15468) );
  AND U19579 ( .A(n15842), .B(n15843), .Z(n15840) );
  AND U19580 ( .A(b[21]), .B(a[64]), .Z(n15839) );
  XOR U19581 ( .A(n15845), .B(n15846), .Z(n15473) );
  AND U19582 ( .A(n15847), .B(n15848), .Z(n15845) );
  AND U19583 ( .A(b[20]), .B(a[65]), .Z(n15844) );
  XOR U19584 ( .A(n15850), .B(n15851), .Z(n15478) );
  AND U19585 ( .A(n15852), .B(n15853), .Z(n15850) );
  AND U19586 ( .A(b[19]), .B(a[66]), .Z(n15849) );
  XOR U19587 ( .A(n15855), .B(n15856), .Z(n15483) );
  AND U19588 ( .A(n15857), .B(n15858), .Z(n15855) );
  AND U19589 ( .A(b[18]), .B(a[67]), .Z(n15854) );
  XOR U19590 ( .A(n15860), .B(n15861), .Z(n15488) );
  AND U19591 ( .A(n15862), .B(n15863), .Z(n15860) );
  AND U19592 ( .A(b[17]), .B(a[68]), .Z(n15859) );
  XOR U19593 ( .A(n15865), .B(n15866), .Z(n15493) );
  AND U19594 ( .A(n15867), .B(n15868), .Z(n15865) );
  AND U19595 ( .A(b[16]), .B(a[69]), .Z(n15864) );
  XOR U19596 ( .A(n15870), .B(n15871), .Z(n15498) );
  AND U19597 ( .A(n15872), .B(n15873), .Z(n15870) );
  AND U19598 ( .A(b[15]), .B(a[70]), .Z(n15869) );
  XOR U19599 ( .A(n15875), .B(n15876), .Z(n15503) );
  AND U19600 ( .A(n15877), .B(n15878), .Z(n15875) );
  AND U19601 ( .A(b[14]), .B(a[71]), .Z(n15874) );
  XOR U19602 ( .A(n15880), .B(n15881), .Z(n15508) );
  AND U19603 ( .A(n15882), .B(n15883), .Z(n15880) );
  AND U19604 ( .A(b[13]), .B(a[72]), .Z(n15879) );
  XOR U19605 ( .A(n15885), .B(n15886), .Z(n15513) );
  AND U19606 ( .A(n15887), .B(n15888), .Z(n15885) );
  AND U19607 ( .A(b[12]), .B(a[73]), .Z(n15884) );
  XOR U19608 ( .A(n15890), .B(n15891), .Z(n15518) );
  AND U19609 ( .A(n15892), .B(n15893), .Z(n15890) );
  AND U19610 ( .A(b[11]), .B(a[74]), .Z(n15889) );
  XOR U19611 ( .A(n15895), .B(n15896), .Z(n15523) );
  AND U19612 ( .A(n15897), .B(n15898), .Z(n15895) );
  AND U19613 ( .A(b[10]), .B(a[75]), .Z(n15894) );
  XOR U19614 ( .A(n15900), .B(n15901), .Z(n15528) );
  AND U19615 ( .A(n15902), .B(n15903), .Z(n15900) );
  AND U19616 ( .A(b[9]), .B(a[76]), .Z(n15899) );
  XOR U19617 ( .A(n15905), .B(n15906), .Z(n15533) );
  AND U19618 ( .A(n15907), .B(n15908), .Z(n15905) );
  AND U19619 ( .A(b[8]), .B(a[77]), .Z(n15904) );
  XOR U19620 ( .A(n15910), .B(n15911), .Z(n15538) );
  AND U19621 ( .A(n15912), .B(n15913), .Z(n15910) );
  AND U19622 ( .A(b[7]), .B(a[78]), .Z(n15909) );
  XOR U19623 ( .A(n15915), .B(n15916), .Z(n15543) );
  AND U19624 ( .A(n15917), .B(n15918), .Z(n15915) );
  AND U19625 ( .A(b[6]), .B(a[79]), .Z(n15914) );
  XOR U19626 ( .A(n15920), .B(n15921), .Z(n15548) );
  AND U19627 ( .A(n15922), .B(n15923), .Z(n15920) );
  AND U19628 ( .A(b[5]), .B(a[80]), .Z(n15919) );
  XOR U19629 ( .A(n15925), .B(n15926), .Z(n15553) );
  AND U19630 ( .A(n15927), .B(n15928), .Z(n15925) );
  AND U19631 ( .A(b[4]), .B(a[81]), .Z(n15924) );
  XOR U19632 ( .A(n15930), .B(n15931), .Z(n15558) );
  AND U19633 ( .A(n15932), .B(n15933), .Z(n15930) );
  AND U19634 ( .A(b[3]), .B(a[82]), .Z(n15929) );
  XOR U19635 ( .A(n15935), .B(n15936), .Z(n15563) );
  OR U19636 ( .A(n15937), .B(n15938), .Z(n15936) );
  AND U19637 ( .A(b[2]), .B(a[83]), .Z(n15934) );
  XNOR U19638 ( .A(n15573), .B(n15939), .Z(n15569) );
  NAND U19639 ( .A(b[1]), .B(a[84]), .Z(n15939) );
  IV U19640 ( .A(n15567), .Z(n15573) );
  ANDN U19641 ( .B(n10299), .A(n10301), .Z(n15567) );
  NAND U19642 ( .A(a[84]), .B(b[0]), .Z(n10301) );
  XOR U19643 ( .A(n15937), .B(n15938), .Z(n10299) );
  XOR U19644 ( .A(n15941), .B(n15932), .Z(n15940) );
  XOR U19645 ( .A(n15927), .B(n15931), .Z(n15942) );
  XOR U19646 ( .A(n15922), .B(n15926), .Z(n15943) );
  XOR U19647 ( .A(n15917), .B(n15921), .Z(n15944) );
  XOR U19648 ( .A(n15912), .B(n15916), .Z(n15945) );
  XOR U19649 ( .A(n15907), .B(n15911), .Z(n15946) );
  XOR U19650 ( .A(n15902), .B(n15906), .Z(n15947) );
  XOR U19651 ( .A(n15897), .B(n15901), .Z(n15948) );
  XOR U19652 ( .A(n15892), .B(n15896), .Z(n15949) );
  XOR U19653 ( .A(n15887), .B(n15891), .Z(n15950) );
  XOR U19654 ( .A(n15882), .B(n15886), .Z(n15951) );
  XOR U19655 ( .A(n15877), .B(n15881), .Z(n15952) );
  XOR U19656 ( .A(n15872), .B(n15876), .Z(n15953) );
  XOR U19657 ( .A(n15867), .B(n15871), .Z(n15954) );
  XOR U19658 ( .A(n15862), .B(n15866), .Z(n15955) );
  XOR U19659 ( .A(n15857), .B(n15861), .Z(n15956) );
  XOR U19660 ( .A(n15852), .B(n15856), .Z(n15957) );
  XOR U19661 ( .A(n15847), .B(n15851), .Z(n15958) );
  XOR U19662 ( .A(n15842), .B(n15846), .Z(n15959) );
  XOR U19663 ( .A(n15837), .B(n15841), .Z(n15960) );
  XOR U19664 ( .A(n15832), .B(n15836), .Z(n15961) );
  XOR U19665 ( .A(n15827), .B(n15831), .Z(n15962) );
  XOR U19666 ( .A(n15822), .B(n15826), .Z(n15963) );
  XOR U19667 ( .A(n15817), .B(n15821), .Z(n15964) );
  XOR U19668 ( .A(n15812), .B(n15816), .Z(n15965) );
  XOR U19669 ( .A(n15807), .B(n15811), .Z(n15966) );
  XOR U19670 ( .A(n15802), .B(n15806), .Z(n15967) );
  XOR U19671 ( .A(n15797), .B(n15801), .Z(n15968) );
  XOR U19672 ( .A(n15792), .B(n15796), .Z(n15969) );
  XOR U19673 ( .A(n15787), .B(n15791), .Z(n15970) );
  XOR U19674 ( .A(n15782), .B(n15786), .Z(n15971) );
  XOR U19675 ( .A(n15777), .B(n15781), .Z(n15972) );
  XOR U19676 ( .A(n15772), .B(n15776), .Z(n15973) );
  XOR U19677 ( .A(n15767), .B(n15771), .Z(n15974) );
  XOR U19678 ( .A(n15762), .B(n15766), .Z(n15975) );
  XOR U19679 ( .A(n15757), .B(n15761), .Z(n15976) );
  XOR U19680 ( .A(n15752), .B(n15756), .Z(n15977) );
  XOR U19681 ( .A(n15747), .B(n15751), .Z(n15978) );
  XOR U19682 ( .A(n15742), .B(n15746), .Z(n15979) );
  XOR U19683 ( .A(n15737), .B(n15741), .Z(n15980) );
  XOR U19684 ( .A(n15732), .B(n15736), .Z(n15981) );
  XOR U19685 ( .A(n15727), .B(n15731), .Z(n15982) );
  XOR U19686 ( .A(n15722), .B(n15726), .Z(n15983) );
  XOR U19687 ( .A(n15717), .B(n15721), .Z(n15984) );
  XOR U19688 ( .A(n15712), .B(n15716), .Z(n15985) );
  XOR U19689 ( .A(n15707), .B(n15711), .Z(n15986) );
  XOR U19690 ( .A(n15697), .B(n15706), .Z(n15987) );
  XOR U19691 ( .A(n15988), .B(n15696), .Z(n15697) );
  AND U19692 ( .A(a[36]), .B(b[48]), .Z(n15988) );
  XNOR U19693 ( .A(n15696), .B(n15702), .Z(n15989) );
  XNOR U19694 ( .A(n15701), .B(n15693), .Z(n15990) );
  XNOR U19695 ( .A(n15692), .B(n15688), .Z(n15991) );
  XNOR U19696 ( .A(n15687), .B(n15683), .Z(n15992) );
  XNOR U19697 ( .A(n15682), .B(n15678), .Z(n15993) );
  XNOR U19698 ( .A(n15677), .B(n15673), .Z(n15994) );
  XNOR U19699 ( .A(n15672), .B(n15668), .Z(n15995) );
  XNOR U19700 ( .A(n15667), .B(n15663), .Z(n15996) );
  XNOR U19701 ( .A(n15662), .B(n15658), .Z(n15997) );
  XNOR U19702 ( .A(n15657), .B(n15653), .Z(n15998) );
  XNOR U19703 ( .A(n15652), .B(n15648), .Z(n15999) );
  XOR U19704 ( .A(n15647), .B(n15644), .Z(n16000) );
  XOR U19705 ( .A(n16001), .B(n16002), .Z(n15644) );
  XOR U19706 ( .A(n15642), .B(n16003), .Z(n16002) );
  XOR U19707 ( .A(n16004), .B(n16005), .Z(n16003) );
  XOR U19708 ( .A(n16006), .B(n16007), .Z(n16005) );
  NAND U19709 ( .A(a[22]), .B(b[62]), .Z(n16007) );
  AND U19710 ( .A(a[21]), .B(b[63]), .Z(n16006) );
  XOR U19711 ( .A(n16008), .B(n16004), .Z(n16001) );
  XOR U19712 ( .A(n16009), .B(n16010), .Z(n16004) );
  ANDN U19713 ( .B(n16011), .A(n16012), .Z(n16009) );
  AND U19714 ( .A(a[23]), .B(b[61]), .Z(n16008) );
  XOR U19715 ( .A(n16013), .B(n15642), .Z(n15643) );
  XOR U19716 ( .A(n16014), .B(n16015), .Z(n15642) );
  AND U19717 ( .A(n16016), .B(n16017), .Z(n16014) );
  AND U19718 ( .A(a[24]), .B(b[60]), .Z(n16013) );
  XOR U19719 ( .A(n16018), .B(n15647), .Z(n15649) );
  XOR U19720 ( .A(n16019), .B(n16020), .Z(n15647) );
  AND U19721 ( .A(n16021), .B(n16022), .Z(n16019) );
  AND U19722 ( .A(a[25]), .B(b[59]), .Z(n16018) );
  XOR U19723 ( .A(n16023), .B(n15652), .Z(n15654) );
  XOR U19724 ( .A(n16024), .B(n16025), .Z(n15652) );
  AND U19725 ( .A(n16026), .B(n16027), .Z(n16024) );
  AND U19726 ( .A(a[26]), .B(b[58]), .Z(n16023) );
  XOR U19727 ( .A(n16028), .B(n15657), .Z(n15659) );
  XOR U19728 ( .A(n16029), .B(n16030), .Z(n15657) );
  AND U19729 ( .A(n16031), .B(n16032), .Z(n16029) );
  AND U19730 ( .A(a[27]), .B(b[57]), .Z(n16028) );
  XOR U19731 ( .A(n16033), .B(n15662), .Z(n15664) );
  XOR U19732 ( .A(n16034), .B(n16035), .Z(n15662) );
  AND U19733 ( .A(n16036), .B(n16037), .Z(n16034) );
  AND U19734 ( .A(a[28]), .B(b[56]), .Z(n16033) );
  XOR U19735 ( .A(n16038), .B(n15667), .Z(n15669) );
  XOR U19736 ( .A(n16039), .B(n16040), .Z(n15667) );
  AND U19737 ( .A(n16041), .B(n16042), .Z(n16039) );
  AND U19738 ( .A(a[29]), .B(b[55]), .Z(n16038) );
  XOR U19739 ( .A(n16043), .B(n15672), .Z(n15674) );
  XOR U19740 ( .A(n16044), .B(n16045), .Z(n15672) );
  AND U19741 ( .A(n16046), .B(n16047), .Z(n16044) );
  AND U19742 ( .A(a[30]), .B(b[54]), .Z(n16043) );
  XOR U19743 ( .A(n16048), .B(n15677), .Z(n15679) );
  XOR U19744 ( .A(n16049), .B(n16050), .Z(n15677) );
  AND U19745 ( .A(n16051), .B(n16052), .Z(n16049) );
  AND U19746 ( .A(a[31]), .B(b[53]), .Z(n16048) );
  XOR U19747 ( .A(n16053), .B(n15682), .Z(n15684) );
  XOR U19748 ( .A(n16054), .B(n16055), .Z(n15682) );
  AND U19749 ( .A(n16056), .B(n16057), .Z(n16054) );
  AND U19750 ( .A(a[32]), .B(b[52]), .Z(n16053) );
  XOR U19751 ( .A(n16058), .B(n15687), .Z(n15689) );
  XOR U19752 ( .A(n16059), .B(n16060), .Z(n15687) );
  AND U19753 ( .A(n16061), .B(n16062), .Z(n16059) );
  AND U19754 ( .A(a[33]), .B(b[51]), .Z(n16058) );
  XOR U19755 ( .A(n16063), .B(n15692), .Z(n15694) );
  XOR U19756 ( .A(n16064), .B(n16065), .Z(n15692) );
  AND U19757 ( .A(n16066), .B(n16067), .Z(n16064) );
  AND U19758 ( .A(a[34]), .B(b[50]), .Z(n16063) );
  XOR U19759 ( .A(n16068), .B(n16069), .Z(n15696) );
  AND U19760 ( .A(n16070), .B(n16071), .Z(n16068) );
  XOR U19761 ( .A(n16072), .B(n15701), .Z(n15703) );
  XOR U19762 ( .A(n16073), .B(n16074), .Z(n15701) );
  AND U19763 ( .A(n16075), .B(n16076), .Z(n16073) );
  AND U19764 ( .A(a[35]), .B(b[49]), .Z(n16072) );
  XOR U19765 ( .A(n16078), .B(n16079), .Z(n15706) );
  AND U19766 ( .A(n16080), .B(n16081), .Z(n16078) );
  AND U19767 ( .A(a[37]), .B(b[47]), .Z(n16077) );
  XOR U19768 ( .A(n16083), .B(n16084), .Z(n15711) );
  AND U19769 ( .A(n16085), .B(n16086), .Z(n16083) );
  AND U19770 ( .A(a[38]), .B(b[46]), .Z(n16082) );
  XOR U19771 ( .A(n16088), .B(n16089), .Z(n15716) );
  AND U19772 ( .A(n16090), .B(n16091), .Z(n16088) );
  AND U19773 ( .A(a[39]), .B(b[45]), .Z(n16087) );
  XOR U19774 ( .A(n16093), .B(n16094), .Z(n15721) );
  AND U19775 ( .A(n16095), .B(n16096), .Z(n16093) );
  AND U19776 ( .A(a[40]), .B(b[44]), .Z(n16092) );
  XOR U19777 ( .A(n16098), .B(n16099), .Z(n15726) );
  AND U19778 ( .A(n16100), .B(n16101), .Z(n16098) );
  AND U19779 ( .A(a[41]), .B(b[43]), .Z(n16097) );
  XOR U19780 ( .A(n16103), .B(n16104), .Z(n15731) );
  AND U19781 ( .A(n16105), .B(n16106), .Z(n16103) );
  AND U19782 ( .A(a[42]), .B(b[42]), .Z(n16102) );
  XOR U19783 ( .A(n16108), .B(n16109), .Z(n15736) );
  AND U19784 ( .A(n16110), .B(n16111), .Z(n16108) );
  AND U19785 ( .A(b[41]), .B(a[43]), .Z(n16107) );
  XOR U19786 ( .A(n16113), .B(n16114), .Z(n15741) );
  AND U19787 ( .A(n16115), .B(n16116), .Z(n16113) );
  AND U19788 ( .A(b[40]), .B(a[44]), .Z(n16112) );
  XOR U19789 ( .A(n16118), .B(n16119), .Z(n15746) );
  AND U19790 ( .A(n16120), .B(n16121), .Z(n16118) );
  AND U19791 ( .A(b[39]), .B(a[45]), .Z(n16117) );
  XOR U19792 ( .A(n16123), .B(n16124), .Z(n15751) );
  AND U19793 ( .A(n16125), .B(n16126), .Z(n16123) );
  AND U19794 ( .A(b[38]), .B(a[46]), .Z(n16122) );
  XOR U19795 ( .A(n16128), .B(n16129), .Z(n15756) );
  AND U19796 ( .A(n16130), .B(n16131), .Z(n16128) );
  AND U19797 ( .A(b[37]), .B(a[47]), .Z(n16127) );
  XOR U19798 ( .A(n16133), .B(n16134), .Z(n15761) );
  AND U19799 ( .A(n16135), .B(n16136), .Z(n16133) );
  AND U19800 ( .A(b[36]), .B(a[48]), .Z(n16132) );
  XOR U19801 ( .A(n16138), .B(n16139), .Z(n15766) );
  AND U19802 ( .A(n16140), .B(n16141), .Z(n16138) );
  AND U19803 ( .A(b[35]), .B(a[49]), .Z(n16137) );
  XOR U19804 ( .A(n16143), .B(n16144), .Z(n15771) );
  AND U19805 ( .A(n16145), .B(n16146), .Z(n16143) );
  AND U19806 ( .A(b[34]), .B(a[50]), .Z(n16142) );
  XOR U19807 ( .A(n16148), .B(n16149), .Z(n15776) );
  AND U19808 ( .A(n16150), .B(n16151), .Z(n16148) );
  AND U19809 ( .A(b[33]), .B(a[51]), .Z(n16147) );
  XOR U19810 ( .A(n16153), .B(n16154), .Z(n15781) );
  AND U19811 ( .A(n16155), .B(n16156), .Z(n16153) );
  AND U19812 ( .A(b[32]), .B(a[52]), .Z(n16152) );
  XOR U19813 ( .A(n16158), .B(n16159), .Z(n15786) );
  AND U19814 ( .A(n16160), .B(n16161), .Z(n16158) );
  AND U19815 ( .A(b[31]), .B(a[53]), .Z(n16157) );
  XOR U19816 ( .A(n16163), .B(n16164), .Z(n15791) );
  AND U19817 ( .A(n16165), .B(n16166), .Z(n16163) );
  AND U19818 ( .A(b[30]), .B(a[54]), .Z(n16162) );
  XOR U19819 ( .A(n16168), .B(n16169), .Z(n15796) );
  AND U19820 ( .A(n16170), .B(n16171), .Z(n16168) );
  AND U19821 ( .A(b[29]), .B(a[55]), .Z(n16167) );
  XOR U19822 ( .A(n16173), .B(n16174), .Z(n15801) );
  AND U19823 ( .A(n16175), .B(n16176), .Z(n16173) );
  AND U19824 ( .A(b[28]), .B(a[56]), .Z(n16172) );
  XOR U19825 ( .A(n16178), .B(n16179), .Z(n15806) );
  AND U19826 ( .A(n16180), .B(n16181), .Z(n16178) );
  AND U19827 ( .A(b[27]), .B(a[57]), .Z(n16177) );
  XOR U19828 ( .A(n16183), .B(n16184), .Z(n15811) );
  AND U19829 ( .A(n16185), .B(n16186), .Z(n16183) );
  AND U19830 ( .A(b[26]), .B(a[58]), .Z(n16182) );
  XOR U19831 ( .A(n16188), .B(n16189), .Z(n15816) );
  AND U19832 ( .A(n16190), .B(n16191), .Z(n16188) );
  AND U19833 ( .A(b[25]), .B(a[59]), .Z(n16187) );
  XOR U19834 ( .A(n16193), .B(n16194), .Z(n15821) );
  AND U19835 ( .A(n16195), .B(n16196), .Z(n16193) );
  AND U19836 ( .A(b[24]), .B(a[60]), .Z(n16192) );
  XOR U19837 ( .A(n16198), .B(n16199), .Z(n15826) );
  AND U19838 ( .A(n16200), .B(n16201), .Z(n16198) );
  AND U19839 ( .A(b[23]), .B(a[61]), .Z(n16197) );
  XOR U19840 ( .A(n16203), .B(n16204), .Z(n15831) );
  AND U19841 ( .A(n16205), .B(n16206), .Z(n16203) );
  AND U19842 ( .A(b[22]), .B(a[62]), .Z(n16202) );
  XOR U19843 ( .A(n16208), .B(n16209), .Z(n15836) );
  AND U19844 ( .A(n16210), .B(n16211), .Z(n16208) );
  AND U19845 ( .A(b[21]), .B(a[63]), .Z(n16207) );
  XOR U19846 ( .A(n16213), .B(n16214), .Z(n15841) );
  AND U19847 ( .A(n16215), .B(n16216), .Z(n16213) );
  AND U19848 ( .A(b[20]), .B(a[64]), .Z(n16212) );
  XOR U19849 ( .A(n16218), .B(n16219), .Z(n15846) );
  AND U19850 ( .A(n16220), .B(n16221), .Z(n16218) );
  AND U19851 ( .A(b[19]), .B(a[65]), .Z(n16217) );
  XOR U19852 ( .A(n16223), .B(n16224), .Z(n15851) );
  AND U19853 ( .A(n16225), .B(n16226), .Z(n16223) );
  AND U19854 ( .A(b[18]), .B(a[66]), .Z(n16222) );
  XOR U19855 ( .A(n16228), .B(n16229), .Z(n15856) );
  AND U19856 ( .A(n16230), .B(n16231), .Z(n16228) );
  AND U19857 ( .A(b[17]), .B(a[67]), .Z(n16227) );
  XOR U19858 ( .A(n16233), .B(n16234), .Z(n15861) );
  AND U19859 ( .A(n16235), .B(n16236), .Z(n16233) );
  AND U19860 ( .A(b[16]), .B(a[68]), .Z(n16232) );
  XOR U19861 ( .A(n16238), .B(n16239), .Z(n15866) );
  AND U19862 ( .A(n16240), .B(n16241), .Z(n16238) );
  AND U19863 ( .A(b[15]), .B(a[69]), .Z(n16237) );
  XOR U19864 ( .A(n16243), .B(n16244), .Z(n15871) );
  AND U19865 ( .A(n16245), .B(n16246), .Z(n16243) );
  AND U19866 ( .A(b[14]), .B(a[70]), .Z(n16242) );
  XOR U19867 ( .A(n16248), .B(n16249), .Z(n15876) );
  AND U19868 ( .A(n16250), .B(n16251), .Z(n16248) );
  AND U19869 ( .A(b[13]), .B(a[71]), .Z(n16247) );
  XOR U19870 ( .A(n16253), .B(n16254), .Z(n15881) );
  AND U19871 ( .A(n16255), .B(n16256), .Z(n16253) );
  AND U19872 ( .A(b[12]), .B(a[72]), .Z(n16252) );
  XOR U19873 ( .A(n16258), .B(n16259), .Z(n15886) );
  AND U19874 ( .A(n16260), .B(n16261), .Z(n16258) );
  AND U19875 ( .A(b[11]), .B(a[73]), .Z(n16257) );
  XOR U19876 ( .A(n16263), .B(n16264), .Z(n15891) );
  AND U19877 ( .A(n16265), .B(n16266), .Z(n16263) );
  AND U19878 ( .A(b[10]), .B(a[74]), .Z(n16262) );
  XOR U19879 ( .A(n16268), .B(n16269), .Z(n15896) );
  AND U19880 ( .A(n16270), .B(n16271), .Z(n16268) );
  AND U19881 ( .A(b[9]), .B(a[75]), .Z(n16267) );
  XOR U19882 ( .A(n16273), .B(n16274), .Z(n15901) );
  AND U19883 ( .A(n16275), .B(n16276), .Z(n16273) );
  AND U19884 ( .A(b[8]), .B(a[76]), .Z(n16272) );
  XOR U19885 ( .A(n16278), .B(n16279), .Z(n15906) );
  AND U19886 ( .A(n16280), .B(n16281), .Z(n16278) );
  AND U19887 ( .A(b[7]), .B(a[77]), .Z(n16277) );
  XOR U19888 ( .A(n16283), .B(n16284), .Z(n15911) );
  AND U19889 ( .A(n16285), .B(n16286), .Z(n16283) );
  AND U19890 ( .A(b[6]), .B(a[78]), .Z(n16282) );
  XOR U19891 ( .A(n16288), .B(n16289), .Z(n15916) );
  AND U19892 ( .A(n16290), .B(n16291), .Z(n16288) );
  AND U19893 ( .A(b[5]), .B(a[79]), .Z(n16287) );
  XOR U19894 ( .A(n16293), .B(n16294), .Z(n15921) );
  AND U19895 ( .A(n16295), .B(n16296), .Z(n16293) );
  AND U19896 ( .A(b[4]), .B(a[80]), .Z(n16292) );
  XOR U19897 ( .A(n16298), .B(n16299), .Z(n15926) );
  AND U19898 ( .A(n16300), .B(n16301), .Z(n16298) );
  AND U19899 ( .A(b[3]), .B(a[81]), .Z(n16297) );
  XOR U19900 ( .A(n16303), .B(n16304), .Z(n15931) );
  OR U19901 ( .A(n16305), .B(n16306), .Z(n16304) );
  AND U19902 ( .A(b[2]), .B(a[82]), .Z(n16302) );
  XNOR U19903 ( .A(n15941), .B(n16307), .Z(n15937) );
  NAND U19904 ( .A(b[1]), .B(a[83]), .Z(n16307) );
  IV U19905 ( .A(n15935), .Z(n15941) );
  ANDN U19906 ( .B(n10302), .A(n10304), .Z(n15935) );
  NAND U19907 ( .A(a[83]), .B(b[0]), .Z(n10304) );
  XOR U19908 ( .A(n16305), .B(n16306), .Z(n10302) );
  XOR U19909 ( .A(n16309), .B(n16300), .Z(n16308) );
  XOR U19910 ( .A(n16295), .B(n16299), .Z(n16310) );
  XOR U19911 ( .A(n16290), .B(n16294), .Z(n16311) );
  XOR U19912 ( .A(n16285), .B(n16289), .Z(n16312) );
  XOR U19913 ( .A(n16280), .B(n16284), .Z(n16313) );
  XOR U19914 ( .A(n16275), .B(n16279), .Z(n16314) );
  XOR U19915 ( .A(n16270), .B(n16274), .Z(n16315) );
  XOR U19916 ( .A(n16265), .B(n16269), .Z(n16316) );
  XOR U19917 ( .A(n16260), .B(n16264), .Z(n16317) );
  XOR U19918 ( .A(n16255), .B(n16259), .Z(n16318) );
  XOR U19919 ( .A(n16250), .B(n16254), .Z(n16319) );
  XOR U19920 ( .A(n16245), .B(n16249), .Z(n16320) );
  XOR U19921 ( .A(n16240), .B(n16244), .Z(n16321) );
  XOR U19922 ( .A(n16235), .B(n16239), .Z(n16322) );
  XOR U19923 ( .A(n16230), .B(n16234), .Z(n16323) );
  XOR U19924 ( .A(n16225), .B(n16229), .Z(n16324) );
  XOR U19925 ( .A(n16220), .B(n16224), .Z(n16325) );
  XOR U19926 ( .A(n16215), .B(n16219), .Z(n16326) );
  XOR U19927 ( .A(n16210), .B(n16214), .Z(n16327) );
  XOR U19928 ( .A(n16205), .B(n16209), .Z(n16328) );
  XOR U19929 ( .A(n16200), .B(n16204), .Z(n16329) );
  XOR U19930 ( .A(n16195), .B(n16199), .Z(n16330) );
  XOR U19931 ( .A(n16190), .B(n16194), .Z(n16331) );
  XOR U19932 ( .A(n16185), .B(n16189), .Z(n16332) );
  XOR U19933 ( .A(n16180), .B(n16184), .Z(n16333) );
  XOR U19934 ( .A(n16175), .B(n16179), .Z(n16334) );
  XOR U19935 ( .A(n16170), .B(n16174), .Z(n16335) );
  XOR U19936 ( .A(n16165), .B(n16169), .Z(n16336) );
  XOR U19937 ( .A(n16160), .B(n16164), .Z(n16337) );
  XOR U19938 ( .A(n16155), .B(n16159), .Z(n16338) );
  XOR U19939 ( .A(n16150), .B(n16154), .Z(n16339) );
  XOR U19940 ( .A(n16145), .B(n16149), .Z(n16340) );
  XOR U19941 ( .A(n16140), .B(n16144), .Z(n16341) );
  XOR U19942 ( .A(n16135), .B(n16139), .Z(n16342) );
  XOR U19943 ( .A(n16130), .B(n16134), .Z(n16343) );
  XOR U19944 ( .A(n16125), .B(n16129), .Z(n16344) );
  XOR U19945 ( .A(n16120), .B(n16124), .Z(n16345) );
  XOR U19946 ( .A(n16115), .B(n16119), .Z(n16346) );
  XOR U19947 ( .A(n16110), .B(n16114), .Z(n16347) );
  XOR U19948 ( .A(n16105), .B(n16109), .Z(n16348) );
  XOR U19949 ( .A(n16100), .B(n16104), .Z(n16349) );
  XOR U19950 ( .A(n16095), .B(n16099), .Z(n16350) );
  XOR U19951 ( .A(n16090), .B(n16094), .Z(n16351) );
  XOR U19952 ( .A(n16085), .B(n16089), .Z(n16352) );
  XOR U19953 ( .A(n16080), .B(n16084), .Z(n16353) );
  XOR U19954 ( .A(n16070), .B(n16079), .Z(n16354) );
  XOR U19955 ( .A(n16355), .B(n16069), .Z(n16070) );
  AND U19956 ( .A(a[36]), .B(b[47]), .Z(n16355) );
  XNOR U19957 ( .A(n16069), .B(n16075), .Z(n16356) );
  XNOR U19958 ( .A(n16074), .B(n16066), .Z(n16357) );
  XNOR U19959 ( .A(n16065), .B(n16061), .Z(n16358) );
  XNOR U19960 ( .A(n16060), .B(n16056), .Z(n16359) );
  XNOR U19961 ( .A(n16055), .B(n16051), .Z(n16360) );
  XNOR U19962 ( .A(n16050), .B(n16046), .Z(n16361) );
  XNOR U19963 ( .A(n16045), .B(n16041), .Z(n16362) );
  XNOR U19964 ( .A(n16040), .B(n16036), .Z(n16363) );
  XNOR U19965 ( .A(n16035), .B(n16031), .Z(n16364) );
  XNOR U19966 ( .A(n16030), .B(n16026), .Z(n16365) );
  XNOR U19967 ( .A(n16025), .B(n16021), .Z(n16366) );
  XNOR U19968 ( .A(n16020), .B(n16016), .Z(n16367) );
  XOR U19969 ( .A(n16015), .B(n16012), .Z(n16368) );
  XOR U19970 ( .A(n16369), .B(n16370), .Z(n16012) );
  XOR U19971 ( .A(n16010), .B(n16371), .Z(n16370) );
  XOR U19972 ( .A(n16372), .B(n16373), .Z(n16371) );
  XOR U19973 ( .A(n16374), .B(n16375), .Z(n16373) );
  NAND U19974 ( .A(a[21]), .B(b[62]), .Z(n16375) );
  AND U19975 ( .A(a[20]), .B(b[63]), .Z(n16374) );
  XOR U19976 ( .A(n16376), .B(n16372), .Z(n16369) );
  XOR U19977 ( .A(n16377), .B(n16378), .Z(n16372) );
  ANDN U19978 ( .B(n16379), .A(n16380), .Z(n16377) );
  AND U19979 ( .A(a[22]), .B(b[61]), .Z(n16376) );
  XOR U19980 ( .A(n16381), .B(n16010), .Z(n16011) );
  XOR U19981 ( .A(n16382), .B(n16383), .Z(n16010) );
  AND U19982 ( .A(n16384), .B(n16385), .Z(n16382) );
  AND U19983 ( .A(a[23]), .B(b[60]), .Z(n16381) );
  XOR U19984 ( .A(n16386), .B(n16015), .Z(n16017) );
  XOR U19985 ( .A(n16387), .B(n16388), .Z(n16015) );
  AND U19986 ( .A(n16389), .B(n16390), .Z(n16387) );
  AND U19987 ( .A(a[24]), .B(b[59]), .Z(n16386) );
  XOR U19988 ( .A(n16391), .B(n16020), .Z(n16022) );
  XOR U19989 ( .A(n16392), .B(n16393), .Z(n16020) );
  AND U19990 ( .A(n16394), .B(n16395), .Z(n16392) );
  AND U19991 ( .A(a[25]), .B(b[58]), .Z(n16391) );
  XOR U19992 ( .A(n16396), .B(n16025), .Z(n16027) );
  XOR U19993 ( .A(n16397), .B(n16398), .Z(n16025) );
  AND U19994 ( .A(n16399), .B(n16400), .Z(n16397) );
  AND U19995 ( .A(a[26]), .B(b[57]), .Z(n16396) );
  XOR U19996 ( .A(n16401), .B(n16030), .Z(n16032) );
  XOR U19997 ( .A(n16402), .B(n16403), .Z(n16030) );
  AND U19998 ( .A(n16404), .B(n16405), .Z(n16402) );
  AND U19999 ( .A(a[27]), .B(b[56]), .Z(n16401) );
  XOR U20000 ( .A(n16406), .B(n16035), .Z(n16037) );
  XOR U20001 ( .A(n16407), .B(n16408), .Z(n16035) );
  AND U20002 ( .A(n16409), .B(n16410), .Z(n16407) );
  AND U20003 ( .A(a[28]), .B(b[55]), .Z(n16406) );
  XOR U20004 ( .A(n16411), .B(n16040), .Z(n16042) );
  XOR U20005 ( .A(n16412), .B(n16413), .Z(n16040) );
  AND U20006 ( .A(n16414), .B(n16415), .Z(n16412) );
  AND U20007 ( .A(a[29]), .B(b[54]), .Z(n16411) );
  XOR U20008 ( .A(n16416), .B(n16045), .Z(n16047) );
  XOR U20009 ( .A(n16417), .B(n16418), .Z(n16045) );
  AND U20010 ( .A(n16419), .B(n16420), .Z(n16417) );
  AND U20011 ( .A(a[30]), .B(b[53]), .Z(n16416) );
  XOR U20012 ( .A(n16421), .B(n16050), .Z(n16052) );
  XOR U20013 ( .A(n16422), .B(n16423), .Z(n16050) );
  AND U20014 ( .A(n16424), .B(n16425), .Z(n16422) );
  AND U20015 ( .A(a[31]), .B(b[52]), .Z(n16421) );
  XOR U20016 ( .A(n16426), .B(n16055), .Z(n16057) );
  XOR U20017 ( .A(n16427), .B(n16428), .Z(n16055) );
  AND U20018 ( .A(n16429), .B(n16430), .Z(n16427) );
  AND U20019 ( .A(a[32]), .B(b[51]), .Z(n16426) );
  XOR U20020 ( .A(n16431), .B(n16060), .Z(n16062) );
  XOR U20021 ( .A(n16432), .B(n16433), .Z(n16060) );
  AND U20022 ( .A(n16434), .B(n16435), .Z(n16432) );
  AND U20023 ( .A(a[33]), .B(b[50]), .Z(n16431) );
  XOR U20024 ( .A(n16436), .B(n16065), .Z(n16067) );
  XOR U20025 ( .A(n16437), .B(n16438), .Z(n16065) );
  AND U20026 ( .A(n16439), .B(n16440), .Z(n16437) );
  AND U20027 ( .A(a[34]), .B(b[49]), .Z(n16436) );
  XOR U20028 ( .A(n16441), .B(n16442), .Z(n16069) );
  AND U20029 ( .A(n16443), .B(n16444), .Z(n16441) );
  XOR U20030 ( .A(n16445), .B(n16074), .Z(n16076) );
  XOR U20031 ( .A(n16446), .B(n16447), .Z(n16074) );
  AND U20032 ( .A(n16448), .B(n16449), .Z(n16446) );
  AND U20033 ( .A(a[35]), .B(b[48]), .Z(n16445) );
  XOR U20034 ( .A(n16451), .B(n16452), .Z(n16079) );
  AND U20035 ( .A(n16453), .B(n16454), .Z(n16451) );
  AND U20036 ( .A(a[37]), .B(b[46]), .Z(n16450) );
  XOR U20037 ( .A(n16456), .B(n16457), .Z(n16084) );
  AND U20038 ( .A(n16458), .B(n16459), .Z(n16456) );
  AND U20039 ( .A(a[38]), .B(b[45]), .Z(n16455) );
  XOR U20040 ( .A(n16461), .B(n16462), .Z(n16089) );
  AND U20041 ( .A(n16463), .B(n16464), .Z(n16461) );
  AND U20042 ( .A(a[39]), .B(b[44]), .Z(n16460) );
  XOR U20043 ( .A(n16466), .B(n16467), .Z(n16094) );
  AND U20044 ( .A(n16468), .B(n16469), .Z(n16466) );
  AND U20045 ( .A(a[40]), .B(b[43]), .Z(n16465) );
  XOR U20046 ( .A(n16471), .B(n16472), .Z(n16099) );
  AND U20047 ( .A(n16473), .B(n16474), .Z(n16471) );
  AND U20048 ( .A(a[41]), .B(b[42]), .Z(n16470) );
  XOR U20049 ( .A(n16476), .B(n16477), .Z(n16104) );
  AND U20050 ( .A(n16478), .B(n16479), .Z(n16476) );
  AND U20051 ( .A(b[41]), .B(a[42]), .Z(n16475) );
  XOR U20052 ( .A(n16481), .B(n16482), .Z(n16109) );
  AND U20053 ( .A(n16483), .B(n16484), .Z(n16481) );
  AND U20054 ( .A(b[40]), .B(a[43]), .Z(n16480) );
  XOR U20055 ( .A(n16486), .B(n16487), .Z(n16114) );
  AND U20056 ( .A(n16488), .B(n16489), .Z(n16486) );
  AND U20057 ( .A(b[39]), .B(a[44]), .Z(n16485) );
  XOR U20058 ( .A(n16491), .B(n16492), .Z(n16119) );
  AND U20059 ( .A(n16493), .B(n16494), .Z(n16491) );
  AND U20060 ( .A(b[38]), .B(a[45]), .Z(n16490) );
  XOR U20061 ( .A(n16496), .B(n16497), .Z(n16124) );
  AND U20062 ( .A(n16498), .B(n16499), .Z(n16496) );
  AND U20063 ( .A(b[37]), .B(a[46]), .Z(n16495) );
  XOR U20064 ( .A(n16501), .B(n16502), .Z(n16129) );
  AND U20065 ( .A(n16503), .B(n16504), .Z(n16501) );
  AND U20066 ( .A(b[36]), .B(a[47]), .Z(n16500) );
  XOR U20067 ( .A(n16506), .B(n16507), .Z(n16134) );
  AND U20068 ( .A(n16508), .B(n16509), .Z(n16506) );
  AND U20069 ( .A(b[35]), .B(a[48]), .Z(n16505) );
  XOR U20070 ( .A(n16511), .B(n16512), .Z(n16139) );
  AND U20071 ( .A(n16513), .B(n16514), .Z(n16511) );
  AND U20072 ( .A(b[34]), .B(a[49]), .Z(n16510) );
  XOR U20073 ( .A(n16516), .B(n16517), .Z(n16144) );
  AND U20074 ( .A(n16518), .B(n16519), .Z(n16516) );
  AND U20075 ( .A(b[33]), .B(a[50]), .Z(n16515) );
  XOR U20076 ( .A(n16521), .B(n16522), .Z(n16149) );
  AND U20077 ( .A(n16523), .B(n16524), .Z(n16521) );
  AND U20078 ( .A(b[32]), .B(a[51]), .Z(n16520) );
  XOR U20079 ( .A(n16526), .B(n16527), .Z(n16154) );
  AND U20080 ( .A(n16528), .B(n16529), .Z(n16526) );
  AND U20081 ( .A(b[31]), .B(a[52]), .Z(n16525) );
  XOR U20082 ( .A(n16531), .B(n16532), .Z(n16159) );
  AND U20083 ( .A(n16533), .B(n16534), .Z(n16531) );
  AND U20084 ( .A(b[30]), .B(a[53]), .Z(n16530) );
  XOR U20085 ( .A(n16536), .B(n16537), .Z(n16164) );
  AND U20086 ( .A(n16538), .B(n16539), .Z(n16536) );
  AND U20087 ( .A(b[29]), .B(a[54]), .Z(n16535) );
  XOR U20088 ( .A(n16541), .B(n16542), .Z(n16169) );
  AND U20089 ( .A(n16543), .B(n16544), .Z(n16541) );
  AND U20090 ( .A(b[28]), .B(a[55]), .Z(n16540) );
  XOR U20091 ( .A(n16546), .B(n16547), .Z(n16174) );
  AND U20092 ( .A(n16548), .B(n16549), .Z(n16546) );
  AND U20093 ( .A(b[27]), .B(a[56]), .Z(n16545) );
  XOR U20094 ( .A(n16551), .B(n16552), .Z(n16179) );
  AND U20095 ( .A(n16553), .B(n16554), .Z(n16551) );
  AND U20096 ( .A(b[26]), .B(a[57]), .Z(n16550) );
  XOR U20097 ( .A(n16556), .B(n16557), .Z(n16184) );
  AND U20098 ( .A(n16558), .B(n16559), .Z(n16556) );
  AND U20099 ( .A(b[25]), .B(a[58]), .Z(n16555) );
  XOR U20100 ( .A(n16561), .B(n16562), .Z(n16189) );
  AND U20101 ( .A(n16563), .B(n16564), .Z(n16561) );
  AND U20102 ( .A(b[24]), .B(a[59]), .Z(n16560) );
  XOR U20103 ( .A(n16566), .B(n16567), .Z(n16194) );
  AND U20104 ( .A(n16568), .B(n16569), .Z(n16566) );
  AND U20105 ( .A(b[23]), .B(a[60]), .Z(n16565) );
  XOR U20106 ( .A(n16571), .B(n16572), .Z(n16199) );
  AND U20107 ( .A(n16573), .B(n16574), .Z(n16571) );
  AND U20108 ( .A(b[22]), .B(a[61]), .Z(n16570) );
  XOR U20109 ( .A(n16576), .B(n16577), .Z(n16204) );
  AND U20110 ( .A(n16578), .B(n16579), .Z(n16576) );
  AND U20111 ( .A(b[21]), .B(a[62]), .Z(n16575) );
  XOR U20112 ( .A(n16581), .B(n16582), .Z(n16209) );
  AND U20113 ( .A(n16583), .B(n16584), .Z(n16581) );
  AND U20114 ( .A(b[20]), .B(a[63]), .Z(n16580) );
  XOR U20115 ( .A(n16586), .B(n16587), .Z(n16214) );
  AND U20116 ( .A(n16588), .B(n16589), .Z(n16586) );
  AND U20117 ( .A(b[19]), .B(a[64]), .Z(n16585) );
  XOR U20118 ( .A(n16591), .B(n16592), .Z(n16219) );
  AND U20119 ( .A(n16593), .B(n16594), .Z(n16591) );
  AND U20120 ( .A(b[18]), .B(a[65]), .Z(n16590) );
  XOR U20121 ( .A(n16596), .B(n16597), .Z(n16224) );
  AND U20122 ( .A(n16598), .B(n16599), .Z(n16596) );
  AND U20123 ( .A(b[17]), .B(a[66]), .Z(n16595) );
  XOR U20124 ( .A(n16601), .B(n16602), .Z(n16229) );
  AND U20125 ( .A(n16603), .B(n16604), .Z(n16601) );
  AND U20126 ( .A(b[16]), .B(a[67]), .Z(n16600) );
  XOR U20127 ( .A(n16606), .B(n16607), .Z(n16234) );
  AND U20128 ( .A(n16608), .B(n16609), .Z(n16606) );
  AND U20129 ( .A(b[15]), .B(a[68]), .Z(n16605) );
  XOR U20130 ( .A(n16611), .B(n16612), .Z(n16239) );
  AND U20131 ( .A(n16613), .B(n16614), .Z(n16611) );
  AND U20132 ( .A(b[14]), .B(a[69]), .Z(n16610) );
  XOR U20133 ( .A(n16616), .B(n16617), .Z(n16244) );
  AND U20134 ( .A(n16618), .B(n16619), .Z(n16616) );
  AND U20135 ( .A(b[13]), .B(a[70]), .Z(n16615) );
  XOR U20136 ( .A(n16621), .B(n16622), .Z(n16249) );
  AND U20137 ( .A(n16623), .B(n16624), .Z(n16621) );
  AND U20138 ( .A(b[12]), .B(a[71]), .Z(n16620) );
  XOR U20139 ( .A(n16626), .B(n16627), .Z(n16254) );
  AND U20140 ( .A(n16628), .B(n16629), .Z(n16626) );
  AND U20141 ( .A(b[11]), .B(a[72]), .Z(n16625) );
  XOR U20142 ( .A(n16631), .B(n16632), .Z(n16259) );
  AND U20143 ( .A(n16633), .B(n16634), .Z(n16631) );
  AND U20144 ( .A(b[10]), .B(a[73]), .Z(n16630) );
  XOR U20145 ( .A(n16636), .B(n16637), .Z(n16264) );
  AND U20146 ( .A(n16638), .B(n16639), .Z(n16636) );
  AND U20147 ( .A(b[9]), .B(a[74]), .Z(n16635) );
  XOR U20148 ( .A(n16641), .B(n16642), .Z(n16269) );
  AND U20149 ( .A(n16643), .B(n16644), .Z(n16641) );
  AND U20150 ( .A(b[8]), .B(a[75]), .Z(n16640) );
  XOR U20151 ( .A(n16646), .B(n16647), .Z(n16274) );
  AND U20152 ( .A(n16648), .B(n16649), .Z(n16646) );
  AND U20153 ( .A(b[7]), .B(a[76]), .Z(n16645) );
  XOR U20154 ( .A(n16651), .B(n16652), .Z(n16279) );
  AND U20155 ( .A(n16653), .B(n16654), .Z(n16651) );
  AND U20156 ( .A(b[6]), .B(a[77]), .Z(n16650) );
  XOR U20157 ( .A(n16656), .B(n16657), .Z(n16284) );
  AND U20158 ( .A(n16658), .B(n16659), .Z(n16656) );
  AND U20159 ( .A(b[5]), .B(a[78]), .Z(n16655) );
  XOR U20160 ( .A(n16661), .B(n16662), .Z(n16289) );
  AND U20161 ( .A(n16663), .B(n16664), .Z(n16661) );
  AND U20162 ( .A(b[4]), .B(a[79]), .Z(n16660) );
  XOR U20163 ( .A(n16666), .B(n16667), .Z(n16294) );
  AND U20164 ( .A(n16668), .B(n16669), .Z(n16666) );
  AND U20165 ( .A(b[3]), .B(a[80]), .Z(n16665) );
  XOR U20166 ( .A(n16671), .B(n16672), .Z(n16299) );
  OR U20167 ( .A(n16673), .B(n16674), .Z(n16672) );
  AND U20168 ( .A(b[2]), .B(a[81]), .Z(n16670) );
  XNOR U20169 ( .A(n16309), .B(n16675), .Z(n16305) );
  NAND U20170 ( .A(b[1]), .B(a[82]), .Z(n16675) );
  IV U20171 ( .A(n16303), .Z(n16309) );
  ANDN U20172 ( .B(n10305), .A(n10307), .Z(n16303) );
  NAND U20173 ( .A(a[82]), .B(b[0]), .Z(n10307) );
  XOR U20174 ( .A(n16673), .B(n16674), .Z(n10305) );
  XOR U20175 ( .A(n16677), .B(n16668), .Z(n16676) );
  XOR U20176 ( .A(n16663), .B(n16667), .Z(n16678) );
  XOR U20177 ( .A(n16658), .B(n16662), .Z(n16679) );
  XOR U20178 ( .A(n16653), .B(n16657), .Z(n16680) );
  XOR U20179 ( .A(n16648), .B(n16652), .Z(n16681) );
  XOR U20180 ( .A(n16643), .B(n16647), .Z(n16682) );
  XOR U20181 ( .A(n16638), .B(n16642), .Z(n16683) );
  XOR U20182 ( .A(n16633), .B(n16637), .Z(n16684) );
  XOR U20183 ( .A(n16628), .B(n16632), .Z(n16685) );
  XOR U20184 ( .A(n16623), .B(n16627), .Z(n16686) );
  XOR U20185 ( .A(n16618), .B(n16622), .Z(n16687) );
  XOR U20186 ( .A(n16613), .B(n16617), .Z(n16688) );
  XOR U20187 ( .A(n16608), .B(n16612), .Z(n16689) );
  XOR U20188 ( .A(n16603), .B(n16607), .Z(n16690) );
  XOR U20189 ( .A(n16598), .B(n16602), .Z(n16691) );
  XOR U20190 ( .A(n16593), .B(n16597), .Z(n16692) );
  XOR U20191 ( .A(n16588), .B(n16592), .Z(n16693) );
  XOR U20192 ( .A(n16583), .B(n16587), .Z(n16694) );
  XOR U20193 ( .A(n16578), .B(n16582), .Z(n16695) );
  XOR U20194 ( .A(n16573), .B(n16577), .Z(n16696) );
  XOR U20195 ( .A(n16568), .B(n16572), .Z(n16697) );
  XOR U20196 ( .A(n16563), .B(n16567), .Z(n16698) );
  XOR U20197 ( .A(n16558), .B(n16562), .Z(n16699) );
  XOR U20198 ( .A(n16553), .B(n16557), .Z(n16700) );
  XOR U20199 ( .A(n16548), .B(n16552), .Z(n16701) );
  XOR U20200 ( .A(n16543), .B(n16547), .Z(n16702) );
  XOR U20201 ( .A(n16538), .B(n16542), .Z(n16703) );
  XOR U20202 ( .A(n16533), .B(n16537), .Z(n16704) );
  XOR U20203 ( .A(n16528), .B(n16532), .Z(n16705) );
  XOR U20204 ( .A(n16523), .B(n16527), .Z(n16706) );
  XOR U20205 ( .A(n16518), .B(n16522), .Z(n16707) );
  XOR U20206 ( .A(n16513), .B(n16517), .Z(n16708) );
  XOR U20207 ( .A(n16508), .B(n16512), .Z(n16709) );
  XOR U20208 ( .A(n16503), .B(n16507), .Z(n16710) );
  XOR U20209 ( .A(n16498), .B(n16502), .Z(n16711) );
  XOR U20210 ( .A(n16493), .B(n16497), .Z(n16712) );
  XOR U20211 ( .A(n16488), .B(n16492), .Z(n16713) );
  XOR U20212 ( .A(n16483), .B(n16487), .Z(n16714) );
  XOR U20213 ( .A(n16478), .B(n16482), .Z(n16715) );
  XOR U20214 ( .A(n16473), .B(n16477), .Z(n16716) );
  XOR U20215 ( .A(n16468), .B(n16472), .Z(n16717) );
  XOR U20216 ( .A(n16463), .B(n16467), .Z(n16718) );
  XOR U20217 ( .A(n16458), .B(n16462), .Z(n16719) );
  XOR U20218 ( .A(n16453), .B(n16457), .Z(n16720) );
  XOR U20219 ( .A(n16443), .B(n16452), .Z(n16721) );
  XOR U20220 ( .A(n16722), .B(n16442), .Z(n16443) );
  AND U20221 ( .A(a[36]), .B(b[46]), .Z(n16722) );
  XNOR U20222 ( .A(n16442), .B(n16448), .Z(n16723) );
  XNOR U20223 ( .A(n16447), .B(n16439), .Z(n16724) );
  XNOR U20224 ( .A(n16438), .B(n16434), .Z(n16725) );
  XNOR U20225 ( .A(n16433), .B(n16429), .Z(n16726) );
  XNOR U20226 ( .A(n16428), .B(n16424), .Z(n16727) );
  XNOR U20227 ( .A(n16423), .B(n16419), .Z(n16728) );
  XNOR U20228 ( .A(n16418), .B(n16414), .Z(n16729) );
  XNOR U20229 ( .A(n16413), .B(n16409), .Z(n16730) );
  XNOR U20230 ( .A(n16408), .B(n16404), .Z(n16731) );
  XNOR U20231 ( .A(n16403), .B(n16399), .Z(n16732) );
  XNOR U20232 ( .A(n16398), .B(n16394), .Z(n16733) );
  XNOR U20233 ( .A(n16393), .B(n16389), .Z(n16734) );
  XNOR U20234 ( .A(n16388), .B(n16384), .Z(n16735) );
  XOR U20235 ( .A(n16383), .B(n16380), .Z(n16736) );
  XOR U20236 ( .A(n16737), .B(n16738), .Z(n16380) );
  XOR U20237 ( .A(n16378), .B(n16739), .Z(n16738) );
  XOR U20238 ( .A(n16740), .B(n16741), .Z(n16739) );
  XOR U20239 ( .A(n16742), .B(n16743), .Z(n16741) );
  NAND U20240 ( .A(a[20]), .B(b[62]), .Z(n16743) );
  AND U20241 ( .A(a[19]), .B(b[63]), .Z(n16742) );
  XOR U20242 ( .A(n16744), .B(n16740), .Z(n16737) );
  XOR U20243 ( .A(n16745), .B(n16746), .Z(n16740) );
  ANDN U20244 ( .B(n16747), .A(n16748), .Z(n16745) );
  AND U20245 ( .A(a[21]), .B(b[61]), .Z(n16744) );
  XOR U20246 ( .A(n16749), .B(n16378), .Z(n16379) );
  XOR U20247 ( .A(n16750), .B(n16751), .Z(n16378) );
  AND U20248 ( .A(n16752), .B(n16753), .Z(n16750) );
  AND U20249 ( .A(a[22]), .B(b[60]), .Z(n16749) );
  XOR U20250 ( .A(n16754), .B(n16383), .Z(n16385) );
  XOR U20251 ( .A(n16755), .B(n16756), .Z(n16383) );
  AND U20252 ( .A(n16757), .B(n16758), .Z(n16755) );
  AND U20253 ( .A(a[23]), .B(b[59]), .Z(n16754) );
  XOR U20254 ( .A(n16759), .B(n16388), .Z(n16390) );
  XOR U20255 ( .A(n16760), .B(n16761), .Z(n16388) );
  AND U20256 ( .A(n16762), .B(n16763), .Z(n16760) );
  AND U20257 ( .A(a[24]), .B(b[58]), .Z(n16759) );
  XOR U20258 ( .A(n16764), .B(n16393), .Z(n16395) );
  XOR U20259 ( .A(n16765), .B(n16766), .Z(n16393) );
  AND U20260 ( .A(n16767), .B(n16768), .Z(n16765) );
  AND U20261 ( .A(a[25]), .B(b[57]), .Z(n16764) );
  XOR U20262 ( .A(n16769), .B(n16398), .Z(n16400) );
  XOR U20263 ( .A(n16770), .B(n16771), .Z(n16398) );
  AND U20264 ( .A(n16772), .B(n16773), .Z(n16770) );
  AND U20265 ( .A(a[26]), .B(b[56]), .Z(n16769) );
  XOR U20266 ( .A(n16774), .B(n16403), .Z(n16405) );
  XOR U20267 ( .A(n16775), .B(n16776), .Z(n16403) );
  AND U20268 ( .A(n16777), .B(n16778), .Z(n16775) );
  AND U20269 ( .A(a[27]), .B(b[55]), .Z(n16774) );
  XOR U20270 ( .A(n16779), .B(n16408), .Z(n16410) );
  XOR U20271 ( .A(n16780), .B(n16781), .Z(n16408) );
  AND U20272 ( .A(n16782), .B(n16783), .Z(n16780) );
  AND U20273 ( .A(a[28]), .B(b[54]), .Z(n16779) );
  XOR U20274 ( .A(n16784), .B(n16413), .Z(n16415) );
  XOR U20275 ( .A(n16785), .B(n16786), .Z(n16413) );
  AND U20276 ( .A(n16787), .B(n16788), .Z(n16785) );
  AND U20277 ( .A(a[29]), .B(b[53]), .Z(n16784) );
  XOR U20278 ( .A(n16789), .B(n16418), .Z(n16420) );
  XOR U20279 ( .A(n16790), .B(n16791), .Z(n16418) );
  AND U20280 ( .A(n16792), .B(n16793), .Z(n16790) );
  AND U20281 ( .A(a[30]), .B(b[52]), .Z(n16789) );
  XOR U20282 ( .A(n16794), .B(n16423), .Z(n16425) );
  XOR U20283 ( .A(n16795), .B(n16796), .Z(n16423) );
  AND U20284 ( .A(n16797), .B(n16798), .Z(n16795) );
  AND U20285 ( .A(a[31]), .B(b[51]), .Z(n16794) );
  XOR U20286 ( .A(n16799), .B(n16428), .Z(n16430) );
  XOR U20287 ( .A(n16800), .B(n16801), .Z(n16428) );
  AND U20288 ( .A(n16802), .B(n16803), .Z(n16800) );
  AND U20289 ( .A(a[32]), .B(b[50]), .Z(n16799) );
  XOR U20290 ( .A(n16804), .B(n16433), .Z(n16435) );
  XOR U20291 ( .A(n16805), .B(n16806), .Z(n16433) );
  AND U20292 ( .A(n16807), .B(n16808), .Z(n16805) );
  AND U20293 ( .A(a[33]), .B(b[49]), .Z(n16804) );
  XOR U20294 ( .A(n16809), .B(n16438), .Z(n16440) );
  XOR U20295 ( .A(n16810), .B(n16811), .Z(n16438) );
  AND U20296 ( .A(n16812), .B(n16813), .Z(n16810) );
  AND U20297 ( .A(a[34]), .B(b[48]), .Z(n16809) );
  XOR U20298 ( .A(n16814), .B(n16815), .Z(n16442) );
  AND U20299 ( .A(n16816), .B(n16817), .Z(n16814) );
  XOR U20300 ( .A(n16818), .B(n16447), .Z(n16449) );
  XOR U20301 ( .A(n16819), .B(n16820), .Z(n16447) );
  AND U20302 ( .A(n16821), .B(n16822), .Z(n16819) );
  AND U20303 ( .A(a[35]), .B(b[47]), .Z(n16818) );
  XOR U20304 ( .A(n16824), .B(n16825), .Z(n16452) );
  AND U20305 ( .A(n16826), .B(n16827), .Z(n16824) );
  AND U20306 ( .A(a[37]), .B(b[45]), .Z(n16823) );
  XOR U20307 ( .A(n16829), .B(n16830), .Z(n16457) );
  AND U20308 ( .A(n16831), .B(n16832), .Z(n16829) );
  AND U20309 ( .A(a[38]), .B(b[44]), .Z(n16828) );
  XOR U20310 ( .A(n16834), .B(n16835), .Z(n16462) );
  AND U20311 ( .A(n16836), .B(n16837), .Z(n16834) );
  AND U20312 ( .A(a[39]), .B(b[43]), .Z(n16833) );
  XOR U20313 ( .A(n16839), .B(n16840), .Z(n16467) );
  AND U20314 ( .A(n16841), .B(n16842), .Z(n16839) );
  AND U20315 ( .A(a[40]), .B(b[42]), .Z(n16838) );
  XOR U20316 ( .A(n16844), .B(n16845), .Z(n16472) );
  AND U20317 ( .A(n16846), .B(n16847), .Z(n16844) );
  AND U20318 ( .A(a[41]), .B(b[41]), .Z(n16843) );
  XOR U20319 ( .A(n16849), .B(n16850), .Z(n16477) );
  AND U20320 ( .A(n16851), .B(n16852), .Z(n16849) );
  AND U20321 ( .A(b[40]), .B(a[42]), .Z(n16848) );
  XOR U20322 ( .A(n16854), .B(n16855), .Z(n16482) );
  AND U20323 ( .A(n16856), .B(n16857), .Z(n16854) );
  AND U20324 ( .A(b[39]), .B(a[43]), .Z(n16853) );
  XOR U20325 ( .A(n16859), .B(n16860), .Z(n16487) );
  AND U20326 ( .A(n16861), .B(n16862), .Z(n16859) );
  AND U20327 ( .A(b[38]), .B(a[44]), .Z(n16858) );
  XOR U20328 ( .A(n16864), .B(n16865), .Z(n16492) );
  AND U20329 ( .A(n16866), .B(n16867), .Z(n16864) );
  AND U20330 ( .A(b[37]), .B(a[45]), .Z(n16863) );
  XOR U20331 ( .A(n16869), .B(n16870), .Z(n16497) );
  AND U20332 ( .A(n16871), .B(n16872), .Z(n16869) );
  AND U20333 ( .A(b[36]), .B(a[46]), .Z(n16868) );
  XOR U20334 ( .A(n16874), .B(n16875), .Z(n16502) );
  AND U20335 ( .A(n16876), .B(n16877), .Z(n16874) );
  AND U20336 ( .A(b[35]), .B(a[47]), .Z(n16873) );
  XOR U20337 ( .A(n16879), .B(n16880), .Z(n16507) );
  AND U20338 ( .A(n16881), .B(n16882), .Z(n16879) );
  AND U20339 ( .A(b[34]), .B(a[48]), .Z(n16878) );
  XOR U20340 ( .A(n16884), .B(n16885), .Z(n16512) );
  AND U20341 ( .A(n16886), .B(n16887), .Z(n16884) );
  AND U20342 ( .A(b[33]), .B(a[49]), .Z(n16883) );
  XOR U20343 ( .A(n16889), .B(n16890), .Z(n16517) );
  AND U20344 ( .A(n16891), .B(n16892), .Z(n16889) );
  AND U20345 ( .A(b[32]), .B(a[50]), .Z(n16888) );
  XOR U20346 ( .A(n16894), .B(n16895), .Z(n16522) );
  AND U20347 ( .A(n16896), .B(n16897), .Z(n16894) );
  AND U20348 ( .A(b[31]), .B(a[51]), .Z(n16893) );
  XOR U20349 ( .A(n16899), .B(n16900), .Z(n16527) );
  AND U20350 ( .A(n16901), .B(n16902), .Z(n16899) );
  AND U20351 ( .A(b[30]), .B(a[52]), .Z(n16898) );
  XOR U20352 ( .A(n16904), .B(n16905), .Z(n16532) );
  AND U20353 ( .A(n16906), .B(n16907), .Z(n16904) );
  AND U20354 ( .A(b[29]), .B(a[53]), .Z(n16903) );
  XOR U20355 ( .A(n16909), .B(n16910), .Z(n16537) );
  AND U20356 ( .A(n16911), .B(n16912), .Z(n16909) );
  AND U20357 ( .A(b[28]), .B(a[54]), .Z(n16908) );
  XOR U20358 ( .A(n16914), .B(n16915), .Z(n16542) );
  AND U20359 ( .A(n16916), .B(n16917), .Z(n16914) );
  AND U20360 ( .A(b[27]), .B(a[55]), .Z(n16913) );
  XOR U20361 ( .A(n16919), .B(n16920), .Z(n16547) );
  AND U20362 ( .A(n16921), .B(n16922), .Z(n16919) );
  AND U20363 ( .A(b[26]), .B(a[56]), .Z(n16918) );
  XOR U20364 ( .A(n16924), .B(n16925), .Z(n16552) );
  AND U20365 ( .A(n16926), .B(n16927), .Z(n16924) );
  AND U20366 ( .A(b[25]), .B(a[57]), .Z(n16923) );
  XOR U20367 ( .A(n16929), .B(n16930), .Z(n16557) );
  AND U20368 ( .A(n16931), .B(n16932), .Z(n16929) );
  AND U20369 ( .A(b[24]), .B(a[58]), .Z(n16928) );
  XOR U20370 ( .A(n16934), .B(n16935), .Z(n16562) );
  AND U20371 ( .A(n16936), .B(n16937), .Z(n16934) );
  AND U20372 ( .A(b[23]), .B(a[59]), .Z(n16933) );
  XOR U20373 ( .A(n16939), .B(n16940), .Z(n16567) );
  AND U20374 ( .A(n16941), .B(n16942), .Z(n16939) );
  AND U20375 ( .A(b[22]), .B(a[60]), .Z(n16938) );
  XOR U20376 ( .A(n16944), .B(n16945), .Z(n16572) );
  AND U20377 ( .A(n16946), .B(n16947), .Z(n16944) );
  AND U20378 ( .A(b[21]), .B(a[61]), .Z(n16943) );
  XOR U20379 ( .A(n16949), .B(n16950), .Z(n16577) );
  AND U20380 ( .A(n16951), .B(n16952), .Z(n16949) );
  AND U20381 ( .A(b[20]), .B(a[62]), .Z(n16948) );
  XOR U20382 ( .A(n16954), .B(n16955), .Z(n16582) );
  AND U20383 ( .A(n16956), .B(n16957), .Z(n16954) );
  AND U20384 ( .A(b[19]), .B(a[63]), .Z(n16953) );
  XOR U20385 ( .A(n16959), .B(n16960), .Z(n16587) );
  AND U20386 ( .A(n16961), .B(n16962), .Z(n16959) );
  AND U20387 ( .A(b[18]), .B(a[64]), .Z(n16958) );
  XOR U20388 ( .A(n16964), .B(n16965), .Z(n16592) );
  AND U20389 ( .A(n16966), .B(n16967), .Z(n16964) );
  AND U20390 ( .A(b[17]), .B(a[65]), .Z(n16963) );
  XOR U20391 ( .A(n16969), .B(n16970), .Z(n16597) );
  AND U20392 ( .A(n16971), .B(n16972), .Z(n16969) );
  AND U20393 ( .A(b[16]), .B(a[66]), .Z(n16968) );
  XOR U20394 ( .A(n16974), .B(n16975), .Z(n16602) );
  AND U20395 ( .A(n16976), .B(n16977), .Z(n16974) );
  AND U20396 ( .A(b[15]), .B(a[67]), .Z(n16973) );
  XOR U20397 ( .A(n16979), .B(n16980), .Z(n16607) );
  AND U20398 ( .A(n16981), .B(n16982), .Z(n16979) );
  AND U20399 ( .A(b[14]), .B(a[68]), .Z(n16978) );
  XOR U20400 ( .A(n16984), .B(n16985), .Z(n16612) );
  AND U20401 ( .A(n16986), .B(n16987), .Z(n16984) );
  AND U20402 ( .A(b[13]), .B(a[69]), .Z(n16983) );
  XOR U20403 ( .A(n16989), .B(n16990), .Z(n16617) );
  AND U20404 ( .A(n16991), .B(n16992), .Z(n16989) );
  AND U20405 ( .A(b[12]), .B(a[70]), .Z(n16988) );
  XOR U20406 ( .A(n16994), .B(n16995), .Z(n16622) );
  AND U20407 ( .A(n16996), .B(n16997), .Z(n16994) );
  AND U20408 ( .A(b[11]), .B(a[71]), .Z(n16993) );
  XOR U20409 ( .A(n16999), .B(n17000), .Z(n16627) );
  AND U20410 ( .A(n17001), .B(n17002), .Z(n16999) );
  AND U20411 ( .A(b[10]), .B(a[72]), .Z(n16998) );
  XOR U20412 ( .A(n17004), .B(n17005), .Z(n16632) );
  AND U20413 ( .A(n17006), .B(n17007), .Z(n17004) );
  AND U20414 ( .A(b[9]), .B(a[73]), .Z(n17003) );
  XOR U20415 ( .A(n17009), .B(n17010), .Z(n16637) );
  AND U20416 ( .A(n17011), .B(n17012), .Z(n17009) );
  AND U20417 ( .A(b[8]), .B(a[74]), .Z(n17008) );
  XOR U20418 ( .A(n17014), .B(n17015), .Z(n16642) );
  AND U20419 ( .A(n17016), .B(n17017), .Z(n17014) );
  AND U20420 ( .A(b[7]), .B(a[75]), .Z(n17013) );
  XOR U20421 ( .A(n17019), .B(n17020), .Z(n16647) );
  AND U20422 ( .A(n17021), .B(n17022), .Z(n17019) );
  AND U20423 ( .A(b[6]), .B(a[76]), .Z(n17018) );
  XOR U20424 ( .A(n17024), .B(n17025), .Z(n16652) );
  AND U20425 ( .A(n17026), .B(n17027), .Z(n17024) );
  AND U20426 ( .A(b[5]), .B(a[77]), .Z(n17023) );
  XOR U20427 ( .A(n17029), .B(n17030), .Z(n16657) );
  AND U20428 ( .A(n17031), .B(n17032), .Z(n17029) );
  AND U20429 ( .A(b[4]), .B(a[78]), .Z(n17028) );
  XOR U20430 ( .A(n17034), .B(n17035), .Z(n16662) );
  AND U20431 ( .A(n17036), .B(n17037), .Z(n17034) );
  AND U20432 ( .A(b[3]), .B(a[79]), .Z(n17033) );
  XOR U20433 ( .A(n17039), .B(n17040), .Z(n16667) );
  OR U20434 ( .A(n17041), .B(n17042), .Z(n17040) );
  AND U20435 ( .A(b[2]), .B(a[80]), .Z(n17038) );
  XNOR U20436 ( .A(n16677), .B(n17043), .Z(n16673) );
  NAND U20437 ( .A(b[1]), .B(a[81]), .Z(n17043) );
  IV U20438 ( .A(n16671), .Z(n16677) );
  ANDN U20439 ( .B(n10308), .A(n10310), .Z(n16671) );
  NAND U20440 ( .A(a[81]), .B(b[0]), .Z(n10310) );
  XOR U20441 ( .A(n17041), .B(n17042), .Z(n10308) );
  XOR U20442 ( .A(n17045), .B(n17036), .Z(n17044) );
  XOR U20443 ( .A(n17031), .B(n17035), .Z(n17046) );
  XOR U20444 ( .A(n17026), .B(n17030), .Z(n17047) );
  XOR U20445 ( .A(n17021), .B(n17025), .Z(n17048) );
  XOR U20446 ( .A(n17016), .B(n17020), .Z(n17049) );
  XOR U20447 ( .A(n17011), .B(n17015), .Z(n17050) );
  XOR U20448 ( .A(n17006), .B(n17010), .Z(n17051) );
  XOR U20449 ( .A(n17001), .B(n17005), .Z(n17052) );
  XOR U20450 ( .A(n16996), .B(n17000), .Z(n17053) );
  XOR U20451 ( .A(n16991), .B(n16995), .Z(n17054) );
  XOR U20452 ( .A(n16986), .B(n16990), .Z(n17055) );
  XOR U20453 ( .A(n16981), .B(n16985), .Z(n17056) );
  XOR U20454 ( .A(n16976), .B(n16980), .Z(n17057) );
  XOR U20455 ( .A(n16971), .B(n16975), .Z(n17058) );
  XOR U20456 ( .A(n16966), .B(n16970), .Z(n17059) );
  XOR U20457 ( .A(n16961), .B(n16965), .Z(n17060) );
  XOR U20458 ( .A(n16956), .B(n16960), .Z(n17061) );
  XOR U20459 ( .A(n16951), .B(n16955), .Z(n17062) );
  XOR U20460 ( .A(n16946), .B(n16950), .Z(n17063) );
  XOR U20461 ( .A(n16941), .B(n16945), .Z(n17064) );
  XOR U20462 ( .A(n16936), .B(n16940), .Z(n17065) );
  XOR U20463 ( .A(n16931), .B(n16935), .Z(n17066) );
  XOR U20464 ( .A(n16926), .B(n16930), .Z(n17067) );
  XOR U20465 ( .A(n16921), .B(n16925), .Z(n17068) );
  XOR U20466 ( .A(n16916), .B(n16920), .Z(n17069) );
  XOR U20467 ( .A(n16911), .B(n16915), .Z(n17070) );
  XOR U20468 ( .A(n16906), .B(n16910), .Z(n17071) );
  XOR U20469 ( .A(n16901), .B(n16905), .Z(n17072) );
  XOR U20470 ( .A(n16896), .B(n16900), .Z(n17073) );
  XOR U20471 ( .A(n16891), .B(n16895), .Z(n17074) );
  XOR U20472 ( .A(n16886), .B(n16890), .Z(n17075) );
  XOR U20473 ( .A(n16881), .B(n16885), .Z(n17076) );
  XOR U20474 ( .A(n16876), .B(n16880), .Z(n17077) );
  XOR U20475 ( .A(n16871), .B(n16875), .Z(n17078) );
  XOR U20476 ( .A(n16866), .B(n16870), .Z(n17079) );
  XOR U20477 ( .A(n16861), .B(n16865), .Z(n17080) );
  XOR U20478 ( .A(n16856), .B(n16860), .Z(n17081) );
  XOR U20479 ( .A(n16851), .B(n16855), .Z(n17082) );
  XOR U20480 ( .A(n16846), .B(n16850), .Z(n17083) );
  XOR U20481 ( .A(n16841), .B(n16845), .Z(n17084) );
  XOR U20482 ( .A(n16836), .B(n16840), .Z(n17085) );
  XOR U20483 ( .A(n16831), .B(n16835), .Z(n17086) );
  XOR U20484 ( .A(n16826), .B(n16830), .Z(n17087) );
  XOR U20485 ( .A(n16816), .B(n16825), .Z(n17088) );
  XOR U20486 ( .A(n17089), .B(n16815), .Z(n16816) );
  AND U20487 ( .A(a[36]), .B(b[45]), .Z(n17089) );
  XNOR U20488 ( .A(n16815), .B(n16821), .Z(n17090) );
  XNOR U20489 ( .A(n16820), .B(n16812), .Z(n17091) );
  XNOR U20490 ( .A(n16811), .B(n16807), .Z(n17092) );
  XNOR U20491 ( .A(n16806), .B(n16802), .Z(n17093) );
  XNOR U20492 ( .A(n16801), .B(n16797), .Z(n17094) );
  XNOR U20493 ( .A(n16796), .B(n16792), .Z(n17095) );
  XNOR U20494 ( .A(n16791), .B(n16787), .Z(n17096) );
  XNOR U20495 ( .A(n16786), .B(n16782), .Z(n17097) );
  XNOR U20496 ( .A(n16781), .B(n16777), .Z(n17098) );
  XNOR U20497 ( .A(n16776), .B(n16772), .Z(n17099) );
  XNOR U20498 ( .A(n16771), .B(n16767), .Z(n17100) );
  XNOR U20499 ( .A(n16766), .B(n16762), .Z(n17101) );
  XNOR U20500 ( .A(n16761), .B(n16757), .Z(n17102) );
  XNOR U20501 ( .A(n16756), .B(n16752), .Z(n17103) );
  XOR U20502 ( .A(n16751), .B(n16748), .Z(n17104) );
  XOR U20503 ( .A(n17105), .B(n17106), .Z(n16748) );
  XOR U20504 ( .A(n16746), .B(n17107), .Z(n17106) );
  XOR U20505 ( .A(n17108), .B(n17109), .Z(n17107) );
  XOR U20506 ( .A(n17110), .B(n17111), .Z(n17109) );
  NAND U20507 ( .A(a[19]), .B(b[62]), .Z(n17111) );
  AND U20508 ( .A(a[18]), .B(b[63]), .Z(n17110) );
  XOR U20509 ( .A(n17112), .B(n17108), .Z(n17105) );
  XOR U20510 ( .A(n17113), .B(n17114), .Z(n17108) );
  ANDN U20511 ( .B(n17115), .A(n17116), .Z(n17113) );
  AND U20512 ( .A(a[20]), .B(b[61]), .Z(n17112) );
  XOR U20513 ( .A(n17117), .B(n16746), .Z(n16747) );
  XOR U20514 ( .A(n17118), .B(n17119), .Z(n16746) );
  AND U20515 ( .A(n17120), .B(n17121), .Z(n17118) );
  AND U20516 ( .A(a[21]), .B(b[60]), .Z(n17117) );
  XOR U20517 ( .A(n17122), .B(n16751), .Z(n16753) );
  XOR U20518 ( .A(n17123), .B(n17124), .Z(n16751) );
  AND U20519 ( .A(n17125), .B(n17126), .Z(n17123) );
  AND U20520 ( .A(a[22]), .B(b[59]), .Z(n17122) );
  XOR U20521 ( .A(n17127), .B(n16756), .Z(n16758) );
  XOR U20522 ( .A(n17128), .B(n17129), .Z(n16756) );
  AND U20523 ( .A(n17130), .B(n17131), .Z(n17128) );
  AND U20524 ( .A(a[23]), .B(b[58]), .Z(n17127) );
  XOR U20525 ( .A(n17132), .B(n16761), .Z(n16763) );
  XOR U20526 ( .A(n17133), .B(n17134), .Z(n16761) );
  AND U20527 ( .A(n17135), .B(n17136), .Z(n17133) );
  AND U20528 ( .A(a[24]), .B(b[57]), .Z(n17132) );
  XOR U20529 ( .A(n17137), .B(n16766), .Z(n16768) );
  XOR U20530 ( .A(n17138), .B(n17139), .Z(n16766) );
  AND U20531 ( .A(n17140), .B(n17141), .Z(n17138) );
  AND U20532 ( .A(a[25]), .B(b[56]), .Z(n17137) );
  XOR U20533 ( .A(n17142), .B(n16771), .Z(n16773) );
  XOR U20534 ( .A(n17143), .B(n17144), .Z(n16771) );
  AND U20535 ( .A(n17145), .B(n17146), .Z(n17143) );
  AND U20536 ( .A(a[26]), .B(b[55]), .Z(n17142) );
  XOR U20537 ( .A(n17147), .B(n16776), .Z(n16778) );
  XOR U20538 ( .A(n17148), .B(n17149), .Z(n16776) );
  AND U20539 ( .A(n17150), .B(n17151), .Z(n17148) );
  AND U20540 ( .A(a[27]), .B(b[54]), .Z(n17147) );
  XOR U20541 ( .A(n17152), .B(n16781), .Z(n16783) );
  XOR U20542 ( .A(n17153), .B(n17154), .Z(n16781) );
  AND U20543 ( .A(n17155), .B(n17156), .Z(n17153) );
  AND U20544 ( .A(a[28]), .B(b[53]), .Z(n17152) );
  XOR U20545 ( .A(n17157), .B(n16786), .Z(n16788) );
  XOR U20546 ( .A(n17158), .B(n17159), .Z(n16786) );
  AND U20547 ( .A(n17160), .B(n17161), .Z(n17158) );
  AND U20548 ( .A(a[29]), .B(b[52]), .Z(n17157) );
  XOR U20549 ( .A(n17162), .B(n16791), .Z(n16793) );
  XOR U20550 ( .A(n17163), .B(n17164), .Z(n16791) );
  AND U20551 ( .A(n17165), .B(n17166), .Z(n17163) );
  AND U20552 ( .A(a[30]), .B(b[51]), .Z(n17162) );
  XOR U20553 ( .A(n17167), .B(n16796), .Z(n16798) );
  XOR U20554 ( .A(n17168), .B(n17169), .Z(n16796) );
  AND U20555 ( .A(n17170), .B(n17171), .Z(n17168) );
  AND U20556 ( .A(a[31]), .B(b[50]), .Z(n17167) );
  XOR U20557 ( .A(n17172), .B(n16801), .Z(n16803) );
  XOR U20558 ( .A(n17173), .B(n17174), .Z(n16801) );
  AND U20559 ( .A(n17175), .B(n17176), .Z(n17173) );
  AND U20560 ( .A(a[32]), .B(b[49]), .Z(n17172) );
  XOR U20561 ( .A(n17177), .B(n16806), .Z(n16808) );
  XOR U20562 ( .A(n17178), .B(n17179), .Z(n16806) );
  AND U20563 ( .A(n17180), .B(n17181), .Z(n17178) );
  AND U20564 ( .A(a[33]), .B(b[48]), .Z(n17177) );
  XOR U20565 ( .A(n17182), .B(n16811), .Z(n16813) );
  XOR U20566 ( .A(n17183), .B(n17184), .Z(n16811) );
  AND U20567 ( .A(n17185), .B(n17186), .Z(n17183) );
  AND U20568 ( .A(a[34]), .B(b[47]), .Z(n17182) );
  XOR U20569 ( .A(n17187), .B(n17188), .Z(n16815) );
  AND U20570 ( .A(n17189), .B(n17190), .Z(n17187) );
  XOR U20571 ( .A(n17191), .B(n16820), .Z(n16822) );
  XOR U20572 ( .A(n17192), .B(n17193), .Z(n16820) );
  AND U20573 ( .A(n17194), .B(n17195), .Z(n17192) );
  AND U20574 ( .A(a[35]), .B(b[46]), .Z(n17191) );
  XOR U20575 ( .A(n17197), .B(n17198), .Z(n16825) );
  AND U20576 ( .A(n17199), .B(n17200), .Z(n17197) );
  AND U20577 ( .A(a[37]), .B(b[44]), .Z(n17196) );
  XOR U20578 ( .A(n17202), .B(n17203), .Z(n16830) );
  AND U20579 ( .A(n17204), .B(n17205), .Z(n17202) );
  AND U20580 ( .A(a[38]), .B(b[43]), .Z(n17201) );
  XOR U20581 ( .A(n17207), .B(n17208), .Z(n16835) );
  AND U20582 ( .A(n17209), .B(n17210), .Z(n17207) );
  AND U20583 ( .A(a[39]), .B(b[42]), .Z(n17206) );
  XOR U20584 ( .A(n17212), .B(n17213), .Z(n16840) );
  AND U20585 ( .A(n17214), .B(n17215), .Z(n17212) );
  AND U20586 ( .A(a[40]), .B(b[41]), .Z(n17211) );
  XOR U20587 ( .A(n17217), .B(n17218), .Z(n16845) );
  AND U20588 ( .A(n17219), .B(n17220), .Z(n17217) );
  AND U20589 ( .A(b[40]), .B(a[41]), .Z(n17216) );
  XOR U20590 ( .A(n17222), .B(n17223), .Z(n16850) );
  AND U20591 ( .A(n17224), .B(n17225), .Z(n17222) );
  AND U20592 ( .A(b[39]), .B(a[42]), .Z(n17221) );
  XOR U20593 ( .A(n17227), .B(n17228), .Z(n16855) );
  AND U20594 ( .A(n17229), .B(n17230), .Z(n17227) );
  AND U20595 ( .A(b[38]), .B(a[43]), .Z(n17226) );
  XOR U20596 ( .A(n17232), .B(n17233), .Z(n16860) );
  AND U20597 ( .A(n17234), .B(n17235), .Z(n17232) );
  AND U20598 ( .A(b[37]), .B(a[44]), .Z(n17231) );
  XOR U20599 ( .A(n17237), .B(n17238), .Z(n16865) );
  AND U20600 ( .A(n17239), .B(n17240), .Z(n17237) );
  AND U20601 ( .A(b[36]), .B(a[45]), .Z(n17236) );
  XOR U20602 ( .A(n17242), .B(n17243), .Z(n16870) );
  AND U20603 ( .A(n17244), .B(n17245), .Z(n17242) );
  AND U20604 ( .A(b[35]), .B(a[46]), .Z(n17241) );
  XOR U20605 ( .A(n17247), .B(n17248), .Z(n16875) );
  AND U20606 ( .A(n17249), .B(n17250), .Z(n17247) );
  AND U20607 ( .A(b[34]), .B(a[47]), .Z(n17246) );
  XOR U20608 ( .A(n17252), .B(n17253), .Z(n16880) );
  AND U20609 ( .A(n17254), .B(n17255), .Z(n17252) );
  AND U20610 ( .A(b[33]), .B(a[48]), .Z(n17251) );
  XOR U20611 ( .A(n17257), .B(n17258), .Z(n16885) );
  AND U20612 ( .A(n17259), .B(n17260), .Z(n17257) );
  AND U20613 ( .A(b[32]), .B(a[49]), .Z(n17256) );
  XOR U20614 ( .A(n17262), .B(n17263), .Z(n16890) );
  AND U20615 ( .A(n17264), .B(n17265), .Z(n17262) );
  AND U20616 ( .A(b[31]), .B(a[50]), .Z(n17261) );
  XOR U20617 ( .A(n17267), .B(n17268), .Z(n16895) );
  AND U20618 ( .A(n17269), .B(n17270), .Z(n17267) );
  AND U20619 ( .A(b[30]), .B(a[51]), .Z(n17266) );
  XOR U20620 ( .A(n17272), .B(n17273), .Z(n16900) );
  AND U20621 ( .A(n17274), .B(n17275), .Z(n17272) );
  AND U20622 ( .A(b[29]), .B(a[52]), .Z(n17271) );
  XOR U20623 ( .A(n17277), .B(n17278), .Z(n16905) );
  AND U20624 ( .A(n17279), .B(n17280), .Z(n17277) );
  AND U20625 ( .A(b[28]), .B(a[53]), .Z(n17276) );
  XOR U20626 ( .A(n17282), .B(n17283), .Z(n16910) );
  AND U20627 ( .A(n17284), .B(n17285), .Z(n17282) );
  AND U20628 ( .A(b[27]), .B(a[54]), .Z(n17281) );
  XOR U20629 ( .A(n17287), .B(n17288), .Z(n16915) );
  AND U20630 ( .A(n17289), .B(n17290), .Z(n17287) );
  AND U20631 ( .A(b[26]), .B(a[55]), .Z(n17286) );
  XOR U20632 ( .A(n17292), .B(n17293), .Z(n16920) );
  AND U20633 ( .A(n17294), .B(n17295), .Z(n17292) );
  AND U20634 ( .A(b[25]), .B(a[56]), .Z(n17291) );
  XOR U20635 ( .A(n17297), .B(n17298), .Z(n16925) );
  AND U20636 ( .A(n17299), .B(n17300), .Z(n17297) );
  AND U20637 ( .A(b[24]), .B(a[57]), .Z(n17296) );
  XOR U20638 ( .A(n17302), .B(n17303), .Z(n16930) );
  AND U20639 ( .A(n17304), .B(n17305), .Z(n17302) );
  AND U20640 ( .A(b[23]), .B(a[58]), .Z(n17301) );
  XOR U20641 ( .A(n17307), .B(n17308), .Z(n16935) );
  AND U20642 ( .A(n17309), .B(n17310), .Z(n17307) );
  AND U20643 ( .A(b[22]), .B(a[59]), .Z(n17306) );
  XOR U20644 ( .A(n17312), .B(n17313), .Z(n16940) );
  AND U20645 ( .A(n17314), .B(n17315), .Z(n17312) );
  AND U20646 ( .A(b[21]), .B(a[60]), .Z(n17311) );
  XOR U20647 ( .A(n17317), .B(n17318), .Z(n16945) );
  AND U20648 ( .A(n17319), .B(n17320), .Z(n17317) );
  AND U20649 ( .A(b[20]), .B(a[61]), .Z(n17316) );
  XOR U20650 ( .A(n17322), .B(n17323), .Z(n16950) );
  AND U20651 ( .A(n17324), .B(n17325), .Z(n17322) );
  AND U20652 ( .A(b[19]), .B(a[62]), .Z(n17321) );
  XOR U20653 ( .A(n17327), .B(n17328), .Z(n16955) );
  AND U20654 ( .A(n17329), .B(n17330), .Z(n17327) );
  AND U20655 ( .A(b[18]), .B(a[63]), .Z(n17326) );
  XOR U20656 ( .A(n17332), .B(n17333), .Z(n16960) );
  AND U20657 ( .A(n17334), .B(n17335), .Z(n17332) );
  AND U20658 ( .A(b[17]), .B(a[64]), .Z(n17331) );
  XOR U20659 ( .A(n17337), .B(n17338), .Z(n16965) );
  AND U20660 ( .A(n17339), .B(n17340), .Z(n17337) );
  AND U20661 ( .A(b[16]), .B(a[65]), .Z(n17336) );
  XOR U20662 ( .A(n17342), .B(n17343), .Z(n16970) );
  AND U20663 ( .A(n17344), .B(n17345), .Z(n17342) );
  AND U20664 ( .A(b[15]), .B(a[66]), .Z(n17341) );
  XOR U20665 ( .A(n17347), .B(n17348), .Z(n16975) );
  AND U20666 ( .A(n17349), .B(n17350), .Z(n17347) );
  AND U20667 ( .A(b[14]), .B(a[67]), .Z(n17346) );
  XOR U20668 ( .A(n17352), .B(n17353), .Z(n16980) );
  AND U20669 ( .A(n17354), .B(n17355), .Z(n17352) );
  AND U20670 ( .A(b[13]), .B(a[68]), .Z(n17351) );
  XOR U20671 ( .A(n17357), .B(n17358), .Z(n16985) );
  AND U20672 ( .A(n17359), .B(n17360), .Z(n17357) );
  AND U20673 ( .A(b[12]), .B(a[69]), .Z(n17356) );
  XOR U20674 ( .A(n17362), .B(n17363), .Z(n16990) );
  AND U20675 ( .A(n17364), .B(n17365), .Z(n17362) );
  AND U20676 ( .A(b[11]), .B(a[70]), .Z(n17361) );
  XOR U20677 ( .A(n17367), .B(n17368), .Z(n16995) );
  AND U20678 ( .A(n17369), .B(n17370), .Z(n17367) );
  AND U20679 ( .A(b[10]), .B(a[71]), .Z(n17366) );
  XOR U20680 ( .A(n17372), .B(n17373), .Z(n17000) );
  AND U20681 ( .A(n17374), .B(n17375), .Z(n17372) );
  AND U20682 ( .A(b[9]), .B(a[72]), .Z(n17371) );
  XOR U20683 ( .A(n17377), .B(n17378), .Z(n17005) );
  AND U20684 ( .A(n17379), .B(n17380), .Z(n17377) );
  AND U20685 ( .A(b[8]), .B(a[73]), .Z(n17376) );
  XOR U20686 ( .A(n17382), .B(n17383), .Z(n17010) );
  AND U20687 ( .A(n17384), .B(n17385), .Z(n17382) );
  AND U20688 ( .A(b[7]), .B(a[74]), .Z(n17381) );
  XOR U20689 ( .A(n17387), .B(n17388), .Z(n17015) );
  AND U20690 ( .A(n17389), .B(n17390), .Z(n17387) );
  AND U20691 ( .A(b[6]), .B(a[75]), .Z(n17386) );
  XOR U20692 ( .A(n17392), .B(n17393), .Z(n17020) );
  AND U20693 ( .A(n17394), .B(n17395), .Z(n17392) );
  AND U20694 ( .A(b[5]), .B(a[76]), .Z(n17391) );
  XOR U20695 ( .A(n17397), .B(n17398), .Z(n17025) );
  AND U20696 ( .A(n17399), .B(n17400), .Z(n17397) );
  AND U20697 ( .A(b[4]), .B(a[77]), .Z(n17396) );
  XOR U20698 ( .A(n17402), .B(n17403), .Z(n17030) );
  AND U20699 ( .A(n17404), .B(n17405), .Z(n17402) );
  AND U20700 ( .A(b[3]), .B(a[78]), .Z(n17401) );
  XOR U20701 ( .A(n17407), .B(n17408), .Z(n17035) );
  OR U20702 ( .A(n17409), .B(n17410), .Z(n17408) );
  AND U20703 ( .A(b[2]), .B(a[79]), .Z(n17406) );
  XNOR U20704 ( .A(n17045), .B(n17411), .Z(n17041) );
  NAND U20705 ( .A(b[1]), .B(a[80]), .Z(n17411) );
  IV U20706 ( .A(n17039), .Z(n17045) );
  ANDN U20707 ( .B(n10311), .A(n10313), .Z(n17039) );
  NAND U20708 ( .A(a[80]), .B(b[0]), .Z(n10313) );
  XOR U20709 ( .A(n17409), .B(n17410), .Z(n10311) );
  XOR U20710 ( .A(n17413), .B(n17404), .Z(n17412) );
  XOR U20711 ( .A(n17399), .B(n17403), .Z(n17414) );
  XOR U20712 ( .A(n17394), .B(n17398), .Z(n17415) );
  XOR U20713 ( .A(n17389), .B(n17393), .Z(n17416) );
  XOR U20714 ( .A(n17384), .B(n17388), .Z(n17417) );
  XOR U20715 ( .A(n17379), .B(n17383), .Z(n17418) );
  XOR U20716 ( .A(n17374), .B(n17378), .Z(n17419) );
  XOR U20717 ( .A(n17369), .B(n17373), .Z(n17420) );
  XOR U20718 ( .A(n17364), .B(n17368), .Z(n17421) );
  XOR U20719 ( .A(n17359), .B(n17363), .Z(n17422) );
  XOR U20720 ( .A(n17354), .B(n17358), .Z(n17423) );
  XOR U20721 ( .A(n17349), .B(n17353), .Z(n17424) );
  XOR U20722 ( .A(n17344), .B(n17348), .Z(n17425) );
  XOR U20723 ( .A(n17339), .B(n17343), .Z(n17426) );
  XOR U20724 ( .A(n17334), .B(n17338), .Z(n17427) );
  XOR U20725 ( .A(n17329), .B(n17333), .Z(n17428) );
  XOR U20726 ( .A(n17324), .B(n17328), .Z(n17429) );
  XOR U20727 ( .A(n17319), .B(n17323), .Z(n17430) );
  XOR U20728 ( .A(n17314), .B(n17318), .Z(n17431) );
  XOR U20729 ( .A(n17309), .B(n17313), .Z(n17432) );
  XOR U20730 ( .A(n17304), .B(n17308), .Z(n17433) );
  XOR U20731 ( .A(n17299), .B(n17303), .Z(n17434) );
  XOR U20732 ( .A(n17294), .B(n17298), .Z(n17435) );
  XOR U20733 ( .A(n17289), .B(n17293), .Z(n17436) );
  XOR U20734 ( .A(n17284), .B(n17288), .Z(n17437) );
  XOR U20735 ( .A(n17279), .B(n17283), .Z(n17438) );
  XOR U20736 ( .A(n17274), .B(n17278), .Z(n17439) );
  XOR U20737 ( .A(n17269), .B(n17273), .Z(n17440) );
  XOR U20738 ( .A(n17264), .B(n17268), .Z(n17441) );
  XOR U20739 ( .A(n17259), .B(n17263), .Z(n17442) );
  XOR U20740 ( .A(n17254), .B(n17258), .Z(n17443) );
  XOR U20741 ( .A(n17249), .B(n17253), .Z(n17444) );
  XOR U20742 ( .A(n17244), .B(n17248), .Z(n17445) );
  XOR U20743 ( .A(n17239), .B(n17243), .Z(n17446) );
  XOR U20744 ( .A(n17234), .B(n17238), .Z(n17447) );
  XOR U20745 ( .A(n17229), .B(n17233), .Z(n17448) );
  XOR U20746 ( .A(n17224), .B(n17228), .Z(n17449) );
  XOR U20747 ( .A(n17219), .B(n17223), .Z(n17450) );
  XOR U20748 ( .A(n17214), .B(n17218), .Z(n17451) );
  XOR U20749 ( .A(n17209), .B(n17213), .Z(n17452) );
  XOR U20750 ( .A(n17204), .B(n17208), .Z(n17453) );
  XOR U20751 ( .A(n17199), .B(n17203), .Z(n17454) );
  XOR U20752 ( .A(n17189), .B(n17198), .Z(n17455) );
  XOR U20753 ( .A(n17456), .B(n17188), .Z(n17189) );
  AND U20754 ( .A(a[36]), .B(b[44]), .Z(n17456) );
  XNOR U20755 ( .A(n17188), .B(n17194), .Z(n17457) );
  XNOR U20756 ( .A(n17193), .B(n17185), .Z(n17458) );
  XNOR U20757 ( .A(n17184), .B(n17180), .Z(n17459) );
  XNOR U20758 ( .A(n17179), .B(n17175), .Z(n17460) );
  XNOR U20759 ( .A(n17174), .B(n17170), .Z(n17461) );
  XNOR U20760 ( .A(n17169), .B(n17165), .Z(n17462) );
  XNOR U20761 ( .A(n17164), .B(n17160), .Z(n17463) );
  XNOR U20762 ( .A(n17159), .B(n17155), .Z(n17464) );
  XNOR U20763 ( .A(n17154), .B(n17150), .Z(n17465) );
  XNOR U20764 ( .A(n17149), .B(n17145), .Z(n17466) );
  XNOR U20765 ( .A(n17144), .B(n17140), .Z(n17467) );
  XNOR U20766 ( .A(n17139), .B(n17135), .Z(n17468) );
  XNOR U20767 ( .A(n17134), .B(n17130), .Z(n17469) );
  XNOR U20768 ( .A(n17129), .B(n17125), .Z(n17470) );
  XNOR U20769 ( .A(n17124), .B(n17120), .Z(n17471) );
  XOR U20770 ( .A(n17119), .B(n17116), .Z(n17472) );
  XOR U20771 ( .A(n17473), .B(n17474), .Z(n17116) );
  XOR U20772 ( .A(n17114), .B(n17475), .Z(n17474) );
  XOR U20773 ( .A(n17476), .B(n17477), .Z(n17475) );
  XOR U20774 ( .A(n17478), .B(n17479), .Z(n17477) );
  NAND U20775 ( .A(a[18]), .B(b[62]), .Z(n17479) );
  AND U20776 ( .A(a[17]), .B(b[63]), .Z(n17478) );
  XOR U20777 ( .A(n17480), .B(n17476), .Z(n17473) );
  XOR U20778 ( .A(n17481), .B(n17482), .Z(n17476) );
  ANDN U20779 ( .B(n17483), .A(n17484), .Z(n17481) );
  AND U20780 ( .A(a[19]), .B(b[61]), .Z(n17480) );
  XOR U20781 ( .A(n17485), .B(n17114), .Z(n17115) );
  XOR U20782 ( .A(n17486), .B(n17487), .Z(n17114) );
  AND U20783 ( .A(n17488), .B(n17489), .Z(n17486) );
  AND U20784 ( .A(a[20]), .B(b[60]), .Z(n17485) );
  XOR U20785 ( .A(n17490), .B(n17119), .Z(n17121) );
  XOR U20786 ( .A(n17491), .B(n17492), .Z(n17119) );
  AND U20787 ( .A(n17493), .B(n17494), .Z(n17491) );
  AND U20788 ( .A(a[21]), .B(b[59]), .Z(n17490) );
  XOR U20789 ( .A(n17495), .B(n17124), .Z(n17126) );
  XOR U20790 ( .A(n17496), .B(n17497), .Z(n17124) );
  AND U20791 ( .A(n17498), .B(n17499), .Z(n17496) );
  AND U20792 ( .A(a[22]), .B(b[58]), .Z(n17495) );
  XOR U20793 ( .A(n17500), .B(n17129), .Z(n17131) );
  XOR U20794 ( .A(n17501), .B(n17502), .Z(n17129) );
  AND U20795 ( .A(n17503), .B(n17504), .Z(n17501) );
  AND U20796 ( .A(a[23]), .B(b[57]), .Z(n17500) );
  XOR U20797 ( .A(n17505), .B(n17134), .Z(n17136) );
  XOR U20798 ( .A(n17506), .B(n17507), .Z(n17134) );
  AND U20799 ( .A(n17508), .B(n17509), .Z(n17506) );
  AND U20800 ( .A(a[24]), .B(b[56]), .Z(n17505) );
  XOR U20801 ( .A(n17510), .B(n17139), .Z(n17141) );
  XOR U20802 ( .A(n17511), .B(n17512), .Z(n17139) );
  AND U20803 ( .A(n17513), .B(n17514), .Z(n17511) );
  AND U20804 ( .A(a[25]), .B(b[55]), .Z(n17510) );
  XOR U20805 ( .A(n17515), .B(n17144), .Z(n17146) );
  XOR U20806 ( .A(n17516), .B(n17517), .Z(n17144) );
  AND U20807 ( .A(n17518), .B(n17519), .Z(n17516) );
  AND U20808 ( .A(a[26]), .B(b[54]), .Z(n17515) );
  XOR U20809 ( .A(n17520), .B(n17149), .Z(n17151) );
  XOR U20810 ( .A(n17521), .B(n17522), .Z(n17149) );
  AND U20811 ( .A(n17523), .B(n17524), .Z(n17521) );
  AND U20812 ( .A(a[27]), .B(b[53]), .Z(n17520) );
  XOR U20813 ( .A(n17525), .B(n17154), .Z(n17156) );
  XOR U20814 ( .A(n17526), .B(n17527), .Z(n17154) );
  AND U20815 ( .A(n17528), .B(n17529), .Z(n17526) );
  AND U20816 ( .A(a[28]), .B(b[52]), .Z(n17525) );
  XOR U20817 ( .A(n17530), .B(n17159), .Z(n17161) );
  XOR U20818 ( .A(n17531), .B(n17532), .Z(n17159) );
  AND U20819 ( .A(n17533), .B(n17534), .Z(n17531) );
  AND U20820 ( .A(a[29]), .B(b[51]), .Z(n17530) );
  XOR U20821 ( .A(n17535), .B(n17164), .Z(n17166) );
  XOR U20822 ( .A(n17536), .B(n17537), .Z(n17164) );
  AND U20823 ( .A(n17538), .B(n17539), .Z(n17536) );
  AND U20824 ( .A(a[30]), .B(b[50]), .Z(n17535) );
  XOR U20825 ( .A(n17540), .B(n17169), .Z(n17171) );
  XOR U20826 ( .A(n17541), .B(n17542), .Z(n17169) );
  AND U20827 ( .A(n17543), .B(n17544), .Z(n17541) );
  AND U20828 ( .A(a[31]), .B(b[49]), .Z(n17540) );
  XOR U20829 ( .A(n17545), .B(n17174), .Z(n17176) );
  XOR U20830 ( .A(n17546), .B(n17547), .Z(n17174) );
  AND U20831 ( .A(n17548), .B(n17549), .Z(n17546) );
  AND U20832 ( .A(a[32]), .B(b[48]), .Z(n17545) );
  XOR U20833 ( .A(n17550), .B(n17179), .Z(n17181) );
  XOR U20834 ( .A(n17551), .B(n17552), .Z(n17179) );
  AND U20835 ( .A(n17553), .B(n17554), .Z(n17551) );
  AND U20836 ( .A(a[33]), .B(b[47]), .Z(n17550) );
  XOR U20837 ( .A(n17555), .B(n17184), .Z(n17186) );
  XOR U20838 ( .A(n17556), .B(n17557), .Z(n17184) );
  AND U20839 ( .A(n17558), .B(n17559), .Z(n17556) );
  AND U20840 ( .A(a[34]), .B(b[46]), .Z(n17555) );
  XOR U20841 ( .A(n17560), .B(n17561), .Z(n17188) );
  AND U20842 ( .A(n17562), .B(n17563), .Z(n17560) );
  XOR U20843 ( .A(n17564), .B(n17193), .Z(n17195) );
  XOR U20844 ( .A(n17565), .B(n17566), .Z(n17193) );
  AND U20845 ( .A(n17567), .B(n17568), .Z(n17565) );
  AND U20846 ( .A(a[35]), .B(b[45]), .Z(n17564) );
  XOR U20847 ( .A(n17570), .B(n17571), .Z(n17198) );
  AND U20848 ( .A(n17572), .B(n17573), .Z(n17570) );
  AND U20849 ( .A(a[37]), .B(b[43]), .Z(n17569) );
  XOR U20850 ( .A(n17575), .B(n17576), .Z(n17203) );
  AND U20851 ( .A(n17577), .B(n17578), .Z(n17575) );
  AND U20852 ( .A(a[38]), .B(b[42]), .Z(n17574) );
  XOR U20853 ( .A(n17580), .B(n17581), .Z(n17208) );
  AND U20854 ( .A(n17582), .B(n17583), .Z(n17580) );
  AND U20855 ( .A(a[39]), .B(b[41]), .Z(n17579) );
  XOR U20856 ( .A(n17585), .B(n17586), .Z(n17213) );
  AND U20857 ( .A(n17587), .B(n17588), .Z(n17585) );
  AND U20858 ( .A(a[40]), .B(b[40]), .Z(n17584) );
  XOR U20859 ( .A(n17590), .B(n17591), .Z(n17218) );
  AND U20860 ( .A(n17592), .B(n17593), .Z(n17590) );
  AND U20861 ( .A(b[39]), .B(a[41]), .Z(n17589) );
  XOR U20862 ( .A(n17595), .B(n17596), .Z(n17223) );
  AND U20863 ( .A(n17597), .B(n17598), .Z(n17595) );
  AND U20864 ( .A(b[38]), .B(a[42]), .Z(n17594) );
  XOR U20865 ( .A(n17600), .B(n17601), .Z(n17228) );
  AND U20866 ( .A(n17602), .B(n17603), .Z(n17600) );
  AND U20867 ( .A(b[37]), .B(a[43]), .Z(n17599) );
  XOR U20868 ( .A(n17605), .B(n17606), .Z(n17233) );
  AND U20869 ( .A(n17607), .B(n17608), .Z(n17605) );
  AND U20870 ( .A(b[36]), .B(a[44]), .Z(n17604) );
  XOR U20871 ( .A(n17610), .B(n17611), .Z(n17238) );
  AND U20872 ( .A(n17612), .B(n17613), .Z(n17610) );
  AND U20873 ( .A(b[35]), .B(a[45]), .Z(n17609) );
  XOR U20874 ( .A(n17615), .B(n17616), .Z(n17243) );
  AND U20875 ( .A(n17617), .B(n17618), .Z(n17615) );
  AND U20876 ( .A(b[34]), .B(a[46]), .Z(n17614) );
  XOR U20877 ( .A(n17620), .B(n17621), .Z(n17248) );
  AND U20878 ( .A(n17622), .B(n17623), .Z(n17620) );
  AND U20879 ( .A(b[33]), .B(a[47]), .Z(n17619) );
  XOR U20880 ( .A(n17625), .B(n17626), .Z(n17253) );
  AND U20881 ( .A(n17627), .B(n17628), .Z(n17625) );
  AND U20882 ( .A(b[32]), .B(a[48]), .Z(n17624) );
  XOR U20883 ( .A(n17630), .B(n17631), .Z(n17258) );
  AND U20884 ( .A(n17632), .B(n17633), .Z(n17630) );
  AND U20885 ( .A(b[31]), .B(a[49]), .Z(n17629) );
  XOR U20886 ( .A(n17635), .B(n17636), .Z(n17263) );
  AND U20887 ( .A(n17637), .B(n17638), .Z(n17635) );
  AND U20888 ( .A(b[30]), .B(a[50]), .Z(n17634) );
  XOR U20889 ( .A(n17640), .B(n17641), .Z(n17268) );
  AND U20890 ( .A(n17642), .B(n17643), .Z(n17640) );
  AND U20891 ( .A(b[29]), .B(a[51]), .Z(n17639) );
  XOR U20892 ( .A(n17645), .B(n17646), .Z(n17273) );
  AND U20893 ( .A(n17647), .B(n17648), .Z(n17645) );
  AND U20894 ( .A(b[28]), .B(a[52]), .Z(n17644) );
  XOR U20895 ( .A(n17650), .B(n17651), .Z(n17278) );
  AND U20896 ( .A(n17652), .B(n17653), .Z(n17650) );
  AND U20897 ( .A(b[27]), .B(a[53]), .Z(n17649) );
  XOR U20898 ( .A(n17655), .B(n17656), .Z(n17283) );
  AND U20899 ( .A(n17657), .B(n17658), .Z(n17655) );
  AND U20900 ( .A(b[26]), .B(a[54]), .Z(n17654) );
  XOR U20901 ( .A(n17660), .B(n17661), .Z(n17288) );
  AND U20902 ( .A(n17662), .B(n17663), .Z(n17660) );
  AND U20903 ( .A(b[25]), .B(a[55]), .Z(n17659) );
  XOR U20904 ( .A(n17665), .B(n17666), .Z(n17293) );
  AND U20905 ( .A(n17667), .B(n17668), .Z(n17665) );
  AND U20906 ( .A(b[24]), .B(a[56]), .Z(n17664) );
  XOR U20907 ( .A(n17670), .B(n17671), .Z(n17298) );
  AND U20908 ( .A(n17672), .B(n17673), .Z(n17670) );
  AND U20909 ( .A(b[23]), .B(a[57]), .Z(n17669) );
  XOR U20910 ( .A(n17675), .B(n17676), .Z(n17303) );
  AND U20911 ( .A(n17677), .B(n17678), .Z(n17675) );
  AND U20912 ( .A(b[22]), .B(a[58]), .Z(n17674) );
  XOR U20913 ( .A(n17680), .B(n17681), .Z(n17308) );
  AND U20914 ( .A(n17682), .B(n17683), .Z(n17680) );
  AND U20915 ( .A(b[21]), .B(a[59]), .Z(n17679) );
  XOR U20916 ( .A(n17685), .B(n17686), .Z(n17313) );
  AND U20917 ( .A(n17687), .B(n17688), .Z(n17685) );
  AND U20918 ( .A(b[20]), .B(a[60]), .Z(n17684) );
  XOR U20919 ( .A(n17690), .B(n17691), .Z(n17318) );
  AND U20920 ( .A(n17692), .B(n17693), .Z(n17690) );
  AND U20921 ( .A(b[19]), .B(a[61]), .Z(n17689) );
  XOR U20922 ( .A(n17695), .B(n17696), .Z(n17323) );
  AND U20923 ( .A(n17697), .B(n17698), .Z(n17695) );
  AND U20924 ( .A(b[18]), .B(a[62]), .Z(n17694) );
  XOR U20925 ( .A(n17700), .B(n17701), .Z(n17328) );
  AND U20926 ( .A(n17702), .B(n17703), .Z(n17700) );
  AND U20927 ( .A(b[17]), .B(a[63]), .Z(n17699) );
  XOR U20928 ( .A(n17705), .B(n17706), .Z(n17333) );
  AND U20929 ( .A(n17707), .B(n17708), .Z(n17705) );
  AND U20930 ( .A(b[16]), .B(a[64]), .Z(n17704) );
  XOR U20931 ( .A(n17710), .B(n17711), .Z(n17338) );
  AND U20932 ( .A(n17712), .B(n17713), .Z(n17710) );
  AND U20933 ( .A(b[15]), .B(a[65]), .Z(n17709) );
  XOR U20934 ( .A(n17715), .B(n17716), .Z(n17343) );
  AND U20935 ( .A(n17717), .B(n17718), .Z(n17715) );
  AND U20936 ( .A(b[14]), .B(a[66]), .Z(n17714) );
  XOR U20937 ( .A(n17720), .B(n17721), .Z(n17348) );
  AND U20938 ( .A(n17722), .B(n17723), .Z(n17720) );
  AND U20939 ( .A(b[13]), .B(a[67]), .Z(n17719) );
  XOR U20940 ( .A(n17725), .B(n17726), .Z(n17353) );
  AND U20941 ( .A(n17727), .B(n17728), .Z(n17725) );
  AND U20942 ( .A(b[12]), .B(a[68]), .Z(n17724) );
  XOR U20943 ( .A(n17730), .B(n17731), .Z(n17358) );
  AND U20944 ( .A(n17732), .B(n17733), .Z(n17730) );
  AND U20945 ( .A(b[11]), .B(a[69]), .Z(n17729) );
  XOR U20946 ( .A(n17735), .B(n17736), .Z(n17363) );
  AND U20947 ( .A(n17737), .B(n17738), .Z(n17735) );
  AND U20948 ( .A(b[10]), .B(a[70]), .Z(n17734) );
  XOR U20949 ( .A(n17740), .B(n17741), .Z(n17368) );
  AND U20950 ( .A(n17742), .B(n17743), .Z(n17740) );
  AND U20951 ( .A(b[9]), .B(a[71]), .Z(n17739) );
  XOR U20952 ( .A(n17745), .B(n17746), .Z(n17373) );
  AND U20953 ( .A(n17747), .B(n17748), .Z(n17745) );
  AND U20954 ( .A(b[8]), .B(a[72]), .Z(n17744) );
  XOR U20955 ( .A(n17750), .B(n17751), .Z(n17378) );
  AND U20956 ( .A(n17752), .B(n17753), .Z(n17750) );
  AND U20957 ( .A(b[7]), .B(a[73]), .Z(n17749) );
  XOR U20958 ( .A(n17755), .B(n17756), .Z(n17383) );
  AND U20959 ( .A(n17757), .B(n17758), .Z(n17755) );
  AND U20960 ( .A(b[6]), .B(a[74]), .Z(n17754) );
  XOR U20961 ( .A(n17760), .B(n17761), .Z(n17388) );
  AND U20962 ( .A(n17762), .B(n17763), .Z(n17760) );
  AND U20963 ( .A(b[5]), .B(a[75]), .Z(n17759) );
  XOR U20964 ( .A(n17765), .B(n17766), .Z(n17393) );
  AND U20965 ( .A(n17767), .B(n17768), .Z(n17765) );
  AND U20966 ( .A(b[4]), .B(a[76]), .Z(n17764) );
  XOR U20967 ( .A(n17770), .B(n17771), .Z(n17398) );
  AND U20968 ( .A(n17772), .B(n17773), .Z(n17770) );
  AND U20969 ( .A(b[3]), .B(a[77]), .Z(n17769) );
  XOR U20970 ( .A(n17775), .B(n17776), .Z(n17403) );
  OR U20971 ( .A(n17777), .B(n17778), .Z(n17776) );
  AND U20972 ( .A(b[2]), .B(a[78]), .Z(n17774) );
  XNOR U20973 ( .A(n17413), .B(n17779), .Z(n17409) );
  NAND U20974 ( .A(b[1]), .B(a[79]), .Z(n17779) );
  IV U20975 ( .A(n17407), .Z(n17413) );
  ANDN U20976 ( .B(n10314), .A(n10316), .Z(n17407) );
  NAND U20977 ( .A(a[79]), .B(b[0]), .Z(n10316) );
  XOR U20978 ( .A(n17777), .B(n17778), .Z(n10314) );
  XOR U20979 ( .A(n17781), .B(n17772), .Z(n17780) );
  XOR U20980 ( .A(n17767), .B(n17771), .Z(n17782) );
  XOR U20981 ( .A(n17762), .B(n17766), .Z(n17783) );
  XOR U20982 ( .A(n17757), .B(n17761), .Z(n17784) );
  XOR U20983 ( .A(n17752), .B(n17756), .Z(n17785) );
  XOR U20984 ( .A(n17747), .B(n17751), .Z(n17786) );
  XOR U20985 ( .A(n17742), .B(n17746), .Z(n17787) );
  XOR U20986 ( .A(n17737), .B(n17741), .Z(n17788) );
  XOR U20987 ( .A(n17732), .B(n17736), .Z(n17789) );
  XOR U20988 ( .A(n17727), .B(n17731), .Z(n17790) );
  XOR U20989 ( .A(n17722), .B(n17726), .Z(n17791) );
  XOR U20990 ( .A(n17717), .B(n17721), .Z(n17792) );
  XOR U20991 ( .A(n17712), .B(n17716), .Z(n17793) );
  XOR U20992 ( .A(n17707), .B(n17711), .Z(n17794) );
  XOR U20993 ( .A(n17702), .B(n17706), .Z(n17795) );
  XOR U20994 ( .A(n17697), .B(n17701), .Z(n17796) );
  XOR U20995 ( .A(n17692), .B(n17696), .Z(n17797) );
  XOR U20996 ( .A(n17687), .B(n17691), .Z(n17798) );
  XOR U20997 ( .A(n17682), .B(n17686), .Z(n17799) );
  XOR U20998 ( .A(n17677), .B(n17681), .Z(n17800) );
  XOR U20999 ( .A(n17672), .B(n17676), .Z(n17801) );
  XOR U21000 ( .A(n17667), .B(n17671), .Z(n17802) );
  XOR U21001 ( .A(n17662), .B(n17666), .Z(n17803) );
  XOR U21002 ( .A(n17657), .B(n17661), .Z(n17804) );
  XOR U21003 ( .A(n17652), .B(n17656), .Z(n17805) );
  XOR U21004 ( .A(n17647), .B(n17651), .Z(n17806) );
  XOR U21005 ( .A(n17642), .B(n17646), .Z(n17807) );
  XOR U21006 ( .A(n17637), .B(n17641), .Z(n17808) );
  XOR U21007 ( .A(n17632), .B(n17636), .Z(n17809) );
  XOR U21008 ( .A(n17627), .B(n17631), .Z(n17810) );
  XOR U21009 ( .A(n17622), .B(n17626), .Z(n17811) );
  XOR U21010 ( .A(n17617), .B(n17621), .Z(n17812) );
  XOR U21011 ( .A(n17612), .B(n17616), .Z(n17813) );
  XOR U21012 ( .A(n17607), .B(n17611), .Z(n17814) );
  XOR U21013 ( .A(n17602), .B(n17606), .Z(n17815) );
  XOR U21014 ( .A(n17597), .B(n17601), .Z(n17816) );
  XOR U21015 ( .A(n17592), .B(n17596), .Z(n17817) );
  XOR U21016 ( .A(n17587), .B(n17591), .Z(n17818) );
  XOR U21017 ( .A(n17582), .B(n17586), .Z(n17819) );
  XOR U21018 ( .A(n17577), .B(n17581), .Z(n17820) );
  XOR U21019 ( .A(n17572), .B(n17576), .Z(n17821) );
  XOR U21020 ( .A(n17562), .B(n17571), .Z(n17822) );
  XOR U21021 ( .A(n17823), .B(n17561), .Z(n17562) );
  AND U21022 ( .A(a[36]), .B(b[43]), .Z(n17823) );
  XNOR U21023 ( .A(n17561), .B(n17567), .Z(n17824) );
  XNOR U21024 ( .A(n17566), .B(n17558), .Z(n17825) );
  XNOR U21025 ( .A(n17557), .B(n17553), .Z(n17826) );
  XNOR U21026 ( .A(n17552), .B(n17548), .Z(n17827) );
  XNOR U21027 ( .A(n17547), .B(n17543), .Z(n17828) );
  XNOR U21028 ( .A(n17542), .B(n17538), .Z(n17829) );
  XNOR U21029 ( .A(n17537), .B(n17533), .Z(n17830) );
  XNOR U21030 ( .A(n17532), .B(n17528), .Z(n17831) );
  XNOR U21031 ( .A(n17527), .B(n17523), .Z(n17832) );
  XNOR U21032 ( .A(n17522), .B(n17518), .Z(n17833) );
  XNOR U21033 ( .A(n17517), .B(n17513), .Z(n17834) );
  XNOR U21034 ( .A(n17512), .B(n17508), .Z(n17835) );
  XNOR U21035 ( .A(n17507), .B(n17503), .Z(n17836) );
  XNOR U21036 ( .A(n17502), .B(n17498), .Z(n17837) );
  XNOR U21037 ( .A(n17497), .B(n17493), .Z(n17838) );
  XNOR U21038 ( .A(n17492), .B(n17488), .Z(n17839) );
  XOR U21039 ( .A(n17487), .B(n17484), .Z(n17840) );
  XOR U21040 ( .A(n17841), .B(n17842), .Z(n17484) );
  XOR U21041 ( .A(n17482), .B(n17843), .Z(n17842) );
  XOR U21042 ( .A(n17844), .B(n17845), .Z(n17843) );
  XOR U21043 ( .A(n17846), .B(n17847), .Z(n17845) );
  NAND U21044 ( .A(a[17]), .B(b[62]), .Z(n17847) );
  AND U21045 ( .A(a[16]), .B(b[63]), .Z(n17846) );
  XOR U21046 ( .A(n17848), .B(n17844), .Z(n17841) );
  XOR U21047 ( .A(n17849), .B(n17850), .Z(n17844) );
  ANDN U21048 ( .B(n17851), .A(n17852), .Z(n17849) );
  AND U21049 ( .A(a[18]), .B(b[61]), .Z(n17848) );
  XOR U21050 ( .A(n17853), .B(n17482), .Z(n17483) );
  XOR U21051 ( .A(n17854), .B(n17855), .Z(n17482) );
  AND U21052 ( .A(n17856), .B(n17857), .Z(n17854) );
  AND U21053 ( .A(a[19]), .B(b[60]), .Z(n17853) );
  XOR U21054 ( .A(n17858), .B(n17487), .Z(n17489) );
  XOR U21055 ( .A(n17859), .B(n17860), .Z(n17487) );
  AND U21056 ( .A(n17861), .B(n17862), .Z(n17859) );
  AND U21057 ( .A(a[20]), .B(b[59]), .Z(n17858) );
  XOR U21058 ( .A(n17863), .B(n17492), .Z(n17494) );
  XOR U21059 ( .A(n17864), .B(n17865), .Z(n17492) );
  AND U21060 ( .A(n17866), .B(n17867), .Z(n17864) );
  AND U21061 ( .A(a[21]), .B(b[58]), .Z(n17863) );
  XOR U21062 ( .A(n17868), .B(n17497), .Z(n17499) );
  XOR U21063 ( .A(n17869), .B(n17870), .Z(n17497) );
  AND U21064 ( .A(n17871), .B(n17872), .Z(n17869) );
  AND U21065 ( .A(a[22]), .B(b[57]), .Z(n17868) );
  XOR U21066 ( .A(n17873), .B(n17502), .Z(n17504) );
  XOR U21067 ( .A(n17874), .B(n17875), .Z(n17502) );
  AND U21068 ( .A(n17876), .B(n17877), .Z(n17874) );
  AND U21069 ( .A(a[23]), .B(b[56]), .Z(n17873) );
  XOR U21070 ( .A(n17878), .B(n17507), .Z(n17509) );
  XOR U21071 ( .A(n17879), .B(n17880), .Z(n17507) );
  AND U21072 ( .A(n17881), .B(n17882), .Z(n17879) );
  AND U21073 ( .A(a[24]), .B(b[55]), .Z(n17878) );
  XOR U21074 ( .A(n17883), .B(n17512), .Z(n17514) );
  XOR U21075 ( .A(n17884), .B(n17885), .Z(n17512) );
  AND U21076 ( .A(n17886), .B(n17887), .Z(n17884) );
  AND U21077 ( .A(a[25]), .B(b[54]), .Z(n17883) );
  XOR U21078 ( .A(n17888), .B(n17517), .Z(n17519) );
  XOR U21079 ( .A(n17889), .B(n17890), .Z(n17517) );
  AND U21080 ( .A(n17891), .B(n17892), .Z(n17889) );
  AND U21081 ( .A(a[26]), .B(b[53]), .Z(n17888) );
  XOR U21082 ( .A(n17893), .B(n17522), .Z(n17524) );
  XOR U21083 ( .A(n17894), .B(n17895), .Z(n17522) );
  AND U21084 ( .A(n17896), .B(n17897), .Z(n17894) );
  AND U21085 ( .A(a[27]), .B(b[52]), .Z(n17893) );
  XOR U21086 ( .A(n17898), .B(n17527), .Z(n17529) );
  XOR U21087 ( .A(n17899), .B(n17900), .Z(n17527) );
  AND U21088 ( .A(n17901), .B(n17902), .Z(n17899) );
  AND U21089 ( .A(a[28]), .B(b[51]), .Z(n17898) );
  XOR U21090 ( .A(n17903), .B(n17532), .Z(n17534) );
  XOR U21091 ( .A(n17904), .B(n17905), .Z(n17532) );
  AND U21092 ( .A(n17906), .B(n17907), .Z(n17904) );
  AND U21093 ( .A(a[29]), .B(b[50]), .Z(n17903) );
  XOR U21094 ( .A(n17908), .B(n17537), .Z(n17539) );
  XOR U21095 ( .A(n17909), .B(n17910), .Z(n17537) );
  AND U21096 ( .A(n17911), .B(n17912), .Z(n17909) );
  AND U21097 ( .A(a[30]), .B(b[49]), .Z(n17908) );
  XOR U21098 ( .A(n17913), .B(n17542), .Z(n17544) );
  XOR U21099 ( .A(n17914), .B(n17915), .Z(n17542) );
  AND U21100 ( .A(n17916), .B(n17917), .Z(n17914) );
  AND U21101 ( .A(a[31]), .B(b[48]), .Z(n17913) );
  XOR U21102 ( .A(n17918), .B(n17547), .Z(n17549) );
  XOR U21103 ( .A(n17919), .B(n17920), .Z(n17547) );
  AND U21104 ( .A(n17921), .B(n17922), .Z(n17919) );
  AND U21105 ( .A(a[32]), .B(b[47]), .Z(n17918) );
  XOR U21106 ( .A(n17923), .B(n17552), .Z(n17554) );
  XOR U21107 ( .A(n17924), .B(n17925), .Z(n17552) );
  AND U21108 ( .A(n17926), .B(n17927), .Z(n17924) );
  AND U21109 ( .A(a[33]), .B(b[46]), .Z(n17923) );
  XOR U21110 ( .A(n17928), .B(n17557), .Z(n17559) );
  XOR U21111 ( .A(n17929), .B(n17930), .Z(n17557) );
  AND U21112 ( .A(n17931), .B(n17932), .Z(n17929) );
  AND U21113 ( .A(a[34]), .B(b[45]), .Z(n17928) );
  XOR U21114 ( .A(n17933), .B(n17934), .Z(n17561) );
  AND U21115 ( .A(n17935), .B(n17936), .Z(n17933) );
  XOR U21116 ( .A(n17937), .B(n17566), .Z(n17568) );
  XOR U21117 ( .A(n17938), .B(n17939), .Z(n17566) );
  AND U21118 ( .A(n17940), .B(n17941), .Z(n17938) );
  AND U21119 ( .A(a[35]), .B(b[44]), .Z(n17937) );
  XOR U21120 ( .A(n17943), .B(n17944), .Z(n17571) );
  AND U21121 ( .A(n17945), .B(n17946), .Z(n17943) );
  AND U21122 ( .A(a[37]), .B(b[42]), .Z(n17942) );
  XOR U21123 ( .A(n17948), .B(n17949), .Z(n17576) );
  AND U21124 ( .A(n17950), .B(n17951), .Z(n17948) );
  AND U21125 ( .A(a[38]), .B(b[41]), .Z(n17947) );
  XOR U21126 ( .A(n17953), .B(n17954), .Z(n17581) );
  AND U21127 ( .A(n17955), .B(n17956), .Z(n17953) );
  AND U21128 ( .A(a[39]), .B(b[40]), .Z(n17952) );
  XOR U21129 ( .A(n17958), .B(n17959), .Z(n17586) );
  AND U21130 ( .A(n17960), .B(n17961), .Z(n17958) );
  AND U21131 ( .A(b[39]), .B(a[40]), .Z(n17957) );
  XOR U21132 ( .A(n17963), .B(n17964), .Z(n17591) );
  AND U21133 ( .A(n17965), .B(n17966), .Z(n17963) );
  AND U21134 ( .A(b[38]), .B(a[41]), .Z(n17962) );
  XOR U21135 ( .A(n17968), .B(n17969), .Z(n17596) );
  AND U21136 ( .A(n17970), .B(n17971), .Z(n17968) );
  AND U21137 ( .A(b[37]), .B(a[42]), .Z(n17967) );
  XOR U21138 ( .A(n17973), .B(n17974), .Z(n17601) );
  AND U21139 ( .A(n17975), .B(n17976), .Z(n17973) );
  AND U21140 ( .A(b[36]), .B(a[43]), .Z(n17972) );
  XOR U21141 ( .A(n17978), .B(n17979), .Z(n17606) );
  AND U21142 ( .A(n17980), .B(n17981), .Z(n17978) );
  AND U21143 ( .A(b[35]), .B(a[44]), .Z(n17977) );
  XOR U21144 ( .A(n17983), .B(n17984), .Z(n17611) );
  AND U21145 ( .A(n17985), .B(n17986), .Z(n17983) );
  AND U21146 ( .A(b[34]), .B(a[45]), .Z(n17982) );
  XOR U21147 ( .A(n17988), .B(n17989), .Z(n17616) );
  AND U21148 ( .A(n17990), .B(n17991), .Z(n17988) );
  AND U21149 ( .A(b[33]), .B(a[46]), .Z(n17987) );
  XOR U21150 ( .A(n17993), .B(n17994), .Z(n17621) );
  AND U21151 ( .A(n17995), .B(n17996), .Z(n17993) );
  AND U21152 ( .A(b[32]), .B(a[47]), .Z(n17992) );
  XOR U21153 ( .A(n17998), .B(n17999), .Z(n17626) );
  AND U21154 ( .A(n18000), .B(n18001), .Z(n17998) );
  AND U21155 ( .A(b[31]), .B(a[48]), .Z(n17997) );
  XOR U21156 ( .A(n18003), .B(n18004), .Z(n17631) );
  AND U21157 ( .A(n18005), .B(n18006), .Z(n18003) );
  AND U21158 ( .A(b[30]), .B(a[49]), .Z(n18002) );
  XOR U21159 ( .A(n18008), .B(n18009), .Z(n17636) );
  AND U21160 ( .A(n18010), .B(n18011), .Z(n18008) );
  AND U21161 ( .A(b[29]), .B(a[50]), .Z(n18007) );
  XOR U21162 ( .A(n18013), .B(n18014), .Z(n17641) );
  AND U21163 ( .A(n18015), .B(n18016), .Z(n18013) );
  AND U21164 ( .A(b[28]), .B(a[51]), .Z(n18012) );
  XOR U21165 ( .A(n18018), .B(n18019), .Z(n17646) );
  AND U21166 ( .A(n18020), .B(n18021), .Z(n18018) );
  AND U21167 ( .A(b[27]), .B(a[52]), .Z(n18017) );
  XOR U21168 ( .A(n18023), .B(n18024), .Z(n17651) );
  AND U21169 ( .A(n18025), .B(n18026), .Z(n18023) );
  AND U21170 ( .A(b[26]), .B(a[53]), .Z(n18022) );
  XOR U21171 ( .A(n18028), .B(n18029), .Z(n17656) );
  AND U21172 ( .A(n18030), .B(n18031), .Z(n18028) );
  AND U21173 ( .A(b[25]), .B(a[54]), .Z(n18027) );
  XOR U21174 ( .A(n18033), .B(n18034), .Z(n17661) );
  AND U21175 ( .A(n18035), .B(n18036), .Z(n18033) );
  AND U21176 ( .A(b[24]), .B(a[55]), .Z(n18032) );
  XOR U21177 ( .A(n18038), .B(n18039), .Z(n17666) );
  AND U21178 ( .A(n18040), .B(n18041), .Z(n18038) );
  AND U21179 ( .A(b[23]), .B(a[56]), .Z(n18037) );
  XOR U21180 ( .A(n18043), .B(n18044), .Z(n17671) );
  AND U21181 ( .A(n18045), .B(n18046), .Z(n18043) );
  AND U21182 ( .A(b[22]), .B(a[57]), .Z(n18042) );
  XOR U21183 ( .A(n18048), .B(n18049), .Z(n17676) );
  AND U21184 ( .A(n18050), .B(n18051), .Z(n18048) );
  AND U21185 ( .A(b[21]), .B(a[58]), .Z(n18047) );
  XOR U21186 ( .A(n18053), .B(n18054), .Z(n17681) );
  AND U21187 ( .A(n18055), .B(n18056), .Z(n18053) );
  AND U21188 ( .A(b[20]), .B(a[59]), .Z(n18052) );
  XOR U21189 ( .A(n18058), .B(n18059), .Z(n17686) );
  AND U21190 ( .A(n18060), .B(n18061), .Z(n18058) );
  AND U21191 ( .A(b[19]), .B(a[60]), .Z(n18057) );
  XOR U21192 ( .A(n18063), .B(n18064), .Z(n17691) );
  AND U21193 ( .A(n18065), .B(n18066), .Z(n18063) );
  AND U21194 ( .A(b[18]), .B(a[61]), .Z(n18062) );
  XOR U21195 ( .A(n18068), .B(n18069), .Z(n17696) );
  AND U21196 ( .A(n18070), .B(n18071), .Z(n18068) );
  AND U21197 ( .A(b[17]), .B(a[62]), .Z(n18067) );
  XOR U21198 ( .A(n18073), .B(n18074), .Z(n17701) );
  AND U21199 ( .A(n18075), .B(n18076), .Z(n18073) );
  AND U21200 ( .A(b[16]), .B(a[63]), .Z(n18072) );
  XOR U21201 ( .A(n18078), .B(n18079), .Z(n17706) );
  AND U21202 ( .A(n18080), .B(n18081), .Z(n18078) );
  AND U21203 ( .A(b[15]), .B(a[64]), .Z(n18077) );
  XOR U21204 ( .A(n18083), .B(n18084), .Z(n17711) );
  AND U21205 ( .A(n18085), .B(n18086), .Z(n18083) );
  AND U21206 ( .A(b[14]), .B(a[65]), .Z(n18082) );
  XOR U21207 ( .A(n18088), .B(n18089), .Z(n17716) );
  AND U21208 ( .A(n18090), .B(n18091), .Z(n18088) );
  AND U21209 ( .A(b[13]), .B(a[66]), .Z(n18087) );
  XOR U21210 ( .A(n18093), .B(n18094), .Z(n17721) );
  AND U21211 ( .A(n18095), .B(n18096), .Z(n18093) );
  AND U21212 ( .A(b[12]), .B(a[67]), .Z(n18092) );
  XOR U21213 ( .A(n18098), .B(n18099), .Z(n17726) );
  AND U21214 ( .A(n18100), .B(n18101), .Z(n18098) );
  AND U21215 ( .A(b[11]), .B(a[68]), .Z(n18097) );
  XOR U21216 ( .A(n18103), .B(n18104), .Z(n17731) );
  AND U21217 ( .A(n18105), .B(n18106), .Z(n18103) );
  AND U21218 ( .A(b[10]), .B(a[69]), .Z(n18102) );
  XOR U21219 ( .A(n18108), .B(n18109), .Z(n17736) );
  AND U21220 ( .A(n18110), .B(n18111), .Z(n18108) );
  AND U21221 ( .A(b[9]), .B(a[70]), .Z(n18107) );
  XOR U21222 ( .A(n18113), .B(n18114), .Z(n17741) );
  AND U21223 ( .A(n18115), .B(n18116), .Z(n18113) );
  AND U21224 ( .A(b[8]), .B(a[71]), .Z(n18112) );
  XOR U21225 ( .A(n18118), .B(n18119), .Z(n17746) );
  AND U21226 ( .A(n18120), .B(n18121), .Z(n18118) );
  AND U21227 ( .A(b[7]), .B(a[72]), .Z(n18117) );
  XOR U21228 ( .A(n18123), .B(n18124), .Z(n17751) );
  AND U21229 ( .A(n18125), .B(n18126), .Z(n18123) );
  AND U21230 ( .A(b[6]), .B(a[73]), .Z(n18122) );
  XOR U21231 ( .A(n18128), .B(n18129), .Z(n17756) );
  AND U21232 ( .A(n18130), .B(n18131), .Z(n18128) );
  AND U21233 ( .A(b[5]), .B(a[74]), .Z(n18127) );
  XOR U21234 ( .A(n18133), .B(n18134), .Z(n17761) );
  AND U21235 ( .A(n18135), .B(n18136), .Z(n18133) );
  AND U21236 ( .A(b[4]), .B(a[75]), .Z(n18132) );
  XOR U21237 ( .A(n18138), .B(n18139), .Z(n17766) );
  AND U21238 ( .A(n18140), .B(n18141), .Z(n18138) );
  AND U21239 ( .A(b[3]), .B(a[76]), .Z(n18137) );
  XOR U21240 ( .A(n18143), .B(n18144), .Z(n17771) );
  OR U21241 ( .A(n18145), .B(n18146), .Z(n18144) );
  AND U21242 ( .A(b[2]), .B(a[77]), .Z(n18142) );
  XNOR U21243 ( .A(n17781), .B(n18147), .Z(n17777) );
  NAND U21244 ( .A(b[1]), .B(a[78]), .Z(n18147) );
  IV U21245 ( .A(n17775), .Z(n17781) );
  ANDN U21246 ( .B(n10317), .A(n10319), .Z(n17775) );
  NAND U21247 ( .A(a[78]), .B(b[0]), .Z(n10319) );
  XOR U21248 ( .A(n18145), .B(n18146), .Z(n10317) );
  XOR U21249 ( .A(n18149), .B(n18140), .Z(n18148) );
  XOR U21250 ( .A(n18135), .B(n18139), .Z(n18150) );
  XOR U21251 ( .A(n18130), .B(n18134), .Z(n18151) );
  XOR U21252 ( .A(n18125), .B(n18129), .Z(n18152) );
  XOR U21253 ( .A(n18120), .B(n18124), .Z(n18153) );
  XOR U21254 ( .A(n18115), .B(n18119), .Z(n18154) );
  XOR U21255 ( .A(n18110), .B(n18114), .Z(n18155) );
  XOR U21256 ( .A(n18105), .B(n18109), .Z(n18156) );
  XOR U21257 ( .A(n18100), .B(n18104), .Z(n18157) );
  XOR U21258 ( .A(n18095), .B(n18099), .Z(n18158) );
  XOR U21259 ( .A(n18090), .B(n18094), .Z(n18159) );
  XOR U21260 ( .A(n18085), .B(n18089), .Z(n18160) );
  XOR U21261 ( .A(n18080), .B(n18084), .Z(n18161) );
  XOR U21262 ( .A(n18075), .B(n18079), .Z(n18162) );
  XOR U21263 ( .A(n18070), .B(n18074), .Z(n18163) );
  XOR U21264 ( .A(n18065), .B(n18069), .Z(n18164) );
  XOR U21265 ( .A(n18060), .B(n18064), .Z(n18165) );
  XOR U21266 ( .A(n18055), .B(n18059), .Z(n18166) );
  XOR U21267 ( .A(n18050), .B(n18054), .Z(n18167) );
  XOR U21268 ( .A(n18045), .B(n18049), .Z(n18168) );
  XOR U21269 ( .A(n18040), .B(n18044), .Z(n18169) );
  XOR U21270 ( .A(n18035), .B(n18039), .Z(n18170) );
  XOR U21271 ( .A(n18030), .B(n18034), .Z(n18171) );
  XOR U21272 ( .A(n18025), .B(n18029), .Z(n18172) );
  XOR U21273 ( .A(n18020), .B(n18024), .Z(n18173) );
  XOR U21274 ( .A(n18015), .B(n18019), .Z(n18174) );
  XOR U21275 ( .A(n18010), .B(n18014), .Z(n18175) );
  XOR U21276 ( .A(n18005), .B(n18009), .Z(n18176) );
  XOR U21277 ( .A(n18000), .B(n18004), .Z(n18177) );
  XOR U21278 ( .A(n17995), .B(n17999), .Z(n18178) );
  XOR U21279 ( .A(n17990), .B(n17994), .Z(n18179) );
  XOR U21280 ( .A(n17985), .B(n17989), .Z(n18180) );
  XOR U21281 ( .A(n17980), .B(n17984), .Z(n18181) );
  XOR U21282 ( .A(n17975), .B(n17979), .Z(n18182) );
  XOR U21283 ( .A(n17970), .B(n17974), .Z(n18183) );
  XOR U21284 ( .A(n17965), .B(n17969), .Z(n18184) );
  XOR U21285 ( .A(n17960), .B(n17964), .Z(n18185) );
  XOR U21286 ( .A(n17955), .B(n17959), .Z(n18186) );
  XOR U21287 ( .A(n17950), .B(n17954), .Z(n18187) );
  XOR U21288 ( .A(n17945), .B(n17949), .Z(n18188) );
  XOR U21289 ( .A(n17935), .B(n17944), .Z(n18189) );
  XOR U21290 ( .A(n18190), .B(n17934), .Z(n17935) );
  AND U21291 ( .A(a[36]), .B(b[42]), .Z(n18190) );
  XNOR U21292 ( .A(n17934), .B(n17940), .Z(n18191) );
  XNOR U21293 ( .A(n17939), .B(n17931), .Z(n18192) );
  XNOR U21294 ( .A(n17930), .B(n17926), .Z(n18193) );
  XNOR U21295 ( .A(n17925), .B(n17921), .Z(n18194) );
  XNOR U21296 ( .A(n17920), .B(n17916), .Z(n18195) );
  XNOR U21297 ( .A(n17915), .B(n17911), .Z(n18196) );
  XNOR U21298 ( .A(n17910), .B(n17906), .Z(n18197) );
  XNOR U21299 ( .A(n17905), .B(n17901), .Z(n18198) );
  XNOR U21300 ( .A(n17900), .B(n17896), .Z(n18199) );
  XNOR U21301 ( .A(n17895), .B(n17891), .Z(n18200) );
  XNOR U21302 ( .A(n17890), .B(n17886), .Z(n18201) );
  XNOR U21303 ( .A(n17885), .B(n17881), .Z(n18202) );
  XNOR U21304 ( .A(n17880), .B(n17876), .Z(n18203) );
  XNOR U21305 ( .A(n17875), .B(n17871), .Z(n18204) );
  XNOR U21306 ( .A(n17870), .B(n17866), .Z(n18205) );
  XNOR U21307 ( .A(n17865), .B(n17861), .Z(n18206) );
  XNOR U21308 ( .A(n17860), .B(n17856), .Z(n18207) );
  XOR U21309 ( .A(n17855), .B(n17852), .Z(n18208) );
  XOR U21310 ( .A(n18209), .B(n18210), .Z(n17852) );
  XOR U21311 ( .A(n17850), .B(n18211), .Z(n18210) );
  XOR U21312 ( .A(n18212), .B(n18213), .Z(n18211) );
  XOR U21313 ( .A(n18214), .B(n18215), .Z(n18213) );
  NAND U21314 ( .A(a[16]), .B(b[62]), .Z(n18215) );
  AND U21315 ( .A(a[15]), .B(b[63]), .Z(n18214) );
  XOR U21316 ( .A(n18216), .B(n18212), .Z(n18209) );
  XOR U21317 ( .A(n18217), .B(n18218), .Z(n18212) );
  ANDN U21318 ( .B(n18219), .A(n18220), .Z(n18217) );
  AND U21319 ( .A(a[17]), .B(b[61]), .Z(n18216) );
  XOR U21320 ( .A(n18221), .B(n17850), .Z(n17851) );
  XOR U21321 ( .A(n18222), .B(n18223), .Z(n17850) );
  AND U21322 ( .A(n18224), .B(n18225), .Z(n18222) );
  AND U21323 ( .A(a[18]), .B(b[60]), .Z(n18221) );
  XOR U21324 ( .A(n18226), .B(n17855), .Z(n17857) );
  XOR U21325 ( .A(n18227), .B(n18228), .Z(n17855) );
  AND U21326 ( .A(n18229), .B(n18230), .Z(n18227) );
  AND U21327 ( .A(a[19]), .B(b[59]), .Z(n18226) );
  XOR U21328 ( .A(n18231), .B(n17860), .Z(n17862) );
  XOR U21329 ( .A(n18232), .B(n18233), .Z(n17860) );
  AND U21330 ( .A(n18234), .B(n18235), .Z(n18232) );
  AND U21331 ( .A(a[20]), .B(b[58]), .Z(n18231) );
  XOR U21332 ( .A(n18236), .B(n17865), .Z(n17867) );
  XOR U21333 ( .A(n18237), .B(n18238), .Z(n17865) );
  AND U21334 ( .A(n18239), .B(n18240), .Z(n18237) );
  AND U21335 ( .A(a[21]), .B(b[57]), .Z(n18236) );
  XOR U21336 ( .A(n18241), .B(n17870), .Z(n17872) );
  XOR U21337 ( .A(n18242), .B(n18243), .Z(n17870) );
  AND U21338 ( .A(n18244), .B(n18245), .Z(n18242) );
  AND U21339 ( .A(a[22]), .B(b[56]), .Z(n18241) );
  XOR U21340 ( .A(n18246), .B(n17875), .Z(n17877) );
  XOR U21341 ( .A(n18247), .B(n18248), .Z(n17875) );
  AND U21342 ( .A(n18249), .B(n18250), .Z(n18247) );
  AND U21343 ( .A(a[23]), .B(b[55]), .Z(n18246) );
  XOR U21344 ( .A(n18251), .B(n17880), .Z(n17882) );
  XOR U21345 ( .A(n18252), .B(n18253), .Z(n17880) );
  AND U21346 ( .A(n18254), .B(n18255), .Z(n18252) );
  AND U21347 ( .A(a[24]), .B(b[54]), .Z(n18251) );
  XOR U21348 ( .A(n18256), .B(n17885), .Z(n17887) );
  XOR U21349 ( .A(n18257), .B(n18258), .Z(n17885) );
  AND U21350 ( .A(n18259), .B(n18260), .Z(n18257) );
  AND U21351 ( .A(a[25]), .B(b[53]), .Z(n18256) );
  XOR U21352 ( .A(n18261), .B(n17890), .Z(n17892) );
  XOR U21353 ( .A(n18262), .B(n18263), .Z(n17890) );
  AND U21354 ( .A(n18264), .B(n18265), .Z(n18262) );
  AND U21355 ( .A(a[26]), .B(b[52]), .Z(n18261) );
  XOR U21356 ( .A(n18266), .B(n17895), .Z(n17897) );
  XOR U21357 ( .A(n18267), .B(n18268), .Z(n17895) );
  AND U21358 ( .A(n18269), .B(n18270), .Z(n18267) );
  AND U21359 ( .A(a[27]), .B(b[51]), .Z(n18266) );
  XOR U21360 ( .A(n18271), .B(n17900), .Z(n17902) );
  XOR U21361 ( .A(n18272), .B(n18273), .Z(n17900) );
  AND U21362 ( .A(n18274), .B(n18275), .Z(n18272) );
  AND U21363 ( .A(a[28]), .B(b[50]), .Z(n18271) );
  XOR U21364 ( .A(n18276), .B(n17905), .Z(n17907) );
  XOR U21365 ( .A(n18277), .B(n18278), .Z(n17905) );
  AND U21366 ( .A(n18279), .B(n18280), .Z(n18277) );
  AND U21367 ( .A(a[29]), .B(b[49]), .Z(n18276) );
  XOR U21368 ( .A(n18281), .B(n17910), .Z(n17912) );
  XOR U21369 ( .A(n18282), .B(n18283), .Z(n17910) );
  AND U21370 ( .A(n18284), .B(n18285), .Z(n18282) );
  AND U21371 ( .A(a[30]), .B(b[48]), .Z(n18281) );
  XOR U21372 ( .A(n18286), .B(n17915), .Z(n17917) );
  XOR U21373 ( .A(n18287), .B(n18288), .Z(n17915) );
  AND U21374 ( .A(n18289), .B(n18290), .Z(n18287) );
  AND U21375 ( .A(a[31]), .B(b[47]), .Z(n18286) );
  XOR U21376 ( .A(n18291), .B(n17920), .Z(n17922) );
  XOR U21377 ( .A(n18292), .B(n18293), .Z(n17920) );
  AND U21378 ( .A(n18294), .B(n18295), .Z(n18292) );
  AND U21379 ( .A(a[32]), .B(b[46]), .Z(n18291) );
  XOR U21380 ( .A(n18296), .B(n17925), .Z(n17927) );
  XOR U21381 ( .A(n18297), .B(n18298), .Z(n17925) );
  AND U21382 ( .A(n18299), .B(n18300), .Z(n18297) );
  AND U21383 ( .A(a[33]), .B(b[45]), .Z(n18296) );
  XOR U21384 ( .A(n18301), .B(n17930), .Z(n17932) );
  XOR U21385 ( .A(n18302), .B(n18303), .Z(n17930) );
  AND U21386 ( .A(n18304), .B(n18305), .Z(n18302) );
  AND U21387 ( .A(a[34]), .B(b[44]), .Z(n18301) );
  XOR U21388 ( .A(n18306), .B(n18307), .Z(n17934) );
  AND U21389 ( .A(n18308), .B(n18309), .Z(n18306) );
  XOR U21390 ( .A(n18310), .B(n17939), .Z(n17941) );
  XOR U21391 ( .A(n18311), .B(n18312), .Z(n17939) );
  AND U21392 ( .A(n18313), .B(n18314), .Z(n18311) );
  AND U21393 ( .A(a[35]), .B(b[43]), .Z(n18310) );
  XOR U21394 ( .A(n18316), .B(n18317), .Z(n17944) );
  AND U21395 ( .A(n18318), .B(n18319), .Z(n18316) );
  AND U21396 ( .A(a[37]), .B(b[41]), .Z(n18315) );
  XOR U21397 ( .A(n18321), .B(n18322), .Z(n17949) );
  AND U21398 ( .A(n18323), .B(n18324), .Z(n18321) );
  AND U21399 ( .A(a[38]), .B(b[40]), .Z(n18320) );
  XOR U21400 ( .A(n18326), .B(n18327), .Z(n17954) );
  AND U21401 ( .A(n18328), .B(n18329), .Z(n18326) );
  AND U21402 ( .A(a[39]), .B(b[39]), .Z(n18325) );
  XOR U21403 ( .A(n18331), .B(n18332), .Z(n17959) );
  AND U21404 ( .A(n18333), .B(n18334), .Z(n18331) );
  AND U21405 ( .A(b[38]), .B(a[40]), .Z(n18330) );
  XOR U21406 ( .A(n18336), .B(n18337), .Z(n17964) );
  AND U21407 ( .A(n18338), .B(n18339), .Z(n18336) );
  AND U21408 ( .A(b[37]), .B(a[41]), .Z(n18335) );
  XOR U21409 ( .A(n18341), .B(n18342), .Z(n17969) );
  AND U21410 ( .A(n18343), .B(n18344), .Z(n18341) );
  AND U21411 ( .A(b[36]), .B(a[42]), .Z(n18340) );
  XOR U21412 ( .A(n18346), .B(n18347), .Z(n17974) );
  AND U21413 ( .A(n18348), .B(n18349), .Z(n18346) );
  AND U21414 ( .A(b[35]), .B(a[43]), .Z(n18345) );
  XOR U21415 ( .A(n18351), .B(n18352), .Z(n17979) );
  AND U21416 ( .A(n18353), .B(n18354), .Z(n18351) );
  AND U21417 ( .A(b[34]), .B(a[44]), .Z(n18350) );
  XOR U21418 ( .A(n18356), .B(n18357), .Z(n17984) );
  AND U21419 ( .A(n18358), .B(n18359), .Z(n18356) );
  AND U21420 ( .A(b[33]), .B(a[45]), .Z(n18355) );
  XOR U21421 ( .A(n18361), .B(n18362), .Z(n17989) );
  AND U21422 ( .A(n18363), .B(n18364), .Z(n18361) );
  AND U21423 ( .A(b[32]), .B(a[46]), .Z(n18360) );
  XOR U21424 ( .A(n18366), .B(n18367), .Z(n17994) );
  AND U21425 ( .A(n18368), .B(n18369), .Z(n18366) );
  AND U21426 ( .A(b[31]), .B(a[47]), .Z(n18365) );
  XOR U21427 ( .A(n18371), .B(n18372), .Z(n17999) );
  AND U21428 ( .A(n18373), .B(n18374), .Z(n18371) );
  AND U21429 ( .A(b[30]), .B(a[48]), .Z(n18370) );
  XOR U21430 ( .A(n18376), .B(n18377), .Z(n18004) );
  AND U21431 ( .A(n18378), .B(n18379), .Z(n18376) );
  AND U21432 ( .A(b[29]), .B(a[49]), .Z(n18375) );
  XOR U21433 ( .A(n18381), .B(n18382), .Z(n18009) );
  AND U21434 ( .A(n18383), .B(n18384), .Z(n18381) );
  AND U21435 ( .A(b[28]), .B(a[50]), .Z(n18380) );
  XOR U21436 ( .A(n18386), .B(n18387), .Z(n18014) );
  AND U21437 ( .A(n18388), .B(n18389), .Z(n18386) );
  AND U21438 ( .A(b[27]), .B(a[51]), .Z(n18385) );
  XOR U21439 ( .A(n18391), .B(n18392), .Z(n18019) );
  AND U21440 ( .A(n18393), .B(n18394), .Z(n18391) );
  AND U21441 ( .A(b[26]), .B(a[52]), .Z(n18390) );
  XOR U21442 ( .A(n18396), .B(n18397), .Z(n18024) );
  AND U21443 ( .A(n18398), .B(n18399), .Z(n18396) );
  AND U21444 ( .A(b[25]), .B(a[53]), .Z(n18395) );
  XOR U21445 ( .A(n18401), .B(n18402), .Z(n18029) );
  AND U21446 ( .A(n18403), .B(n18404), .Z(n18401) );
  AND U21447 ( .A(b[24]), .B(a[54]), .Z(n18400) );
  XOR U21448 ( .A(n18406), .B(n18407), .Z(n18034) );
  AND U21449 ( .A(n18408), .B(n18409), .Z(n18406) );
  AND U21450 ( .A(b[23]), .B(a[55]), .Z(n18405) );
  XOR U21451 ( .A(n18411), .B(n18412), .Z(n18039) );
  AND U21452 ( .A(n18413), .B(n18414), .Z(n18411) );
  AND U21453 ( .A(b[22]), .B(a[56]), .Z(n18410) );
  XOR U21454 ( .A(n18416), .B(n18417), .Z(n18044) );
  AND U21455 ( .A(n18418), .B(n18419), .Z(n18416) );
  AND U21456 ( .A(b[21]), .B(a[57]), .Z(n18415) );
  XOR U21457 ( .A(n18421), .B(n18422), .Z(n18049) );
  AND U21458 ( .A(n18423), .B(n18424), .Z(n18421) );
  AND U21459 ( .A(b[20]), .B(a[58]), .Z(n18420) );
  XOR U21460 ( .A(n18426), .B(n18427), .Z(n18054) );
  AND U21461 ( .A(n18428), .B(n18429), .Z(n18426) );
  AND U21462 ( .A(b[19]), .B(a[59]), .Z(n18425) );
  XOR U21463 ( .A(n18431), .B(n18432), .Z(n18059) );
  AND U21464 ( .A(n18433), .B(n18434), .Z(n18431) );
  AND U21465 ( .A(b[18]), .B(a[60]), .Z(n18430) );
  XOR U21466 ( .A(n18436), .B(n18437), .Z(n18064) );
  AND U21467 ( .A(n18438), .B(n18439), .Z(n18436) );
  AND U21468 ( .A(b[17]), .B(a[61]), .Z(n18435) );
  XOR U21469 ( .A(n18441), .B(n18442), .Z(n18069) );
  AND U21470 ( .A(n18443), .B(n18444), .Z(n18441) );
  AND U21471 ( .A(b[16]), .B(a[62]), .Z(n18440) );
  XOR U21472 ( .A(n18446), .B(n18447), .Z(n18074) );
  AND U21473 ( .A(n18448), .B(n18449), .Z(n18446) );
  AND U21474 ( .A(b[15]), .B(a[63]), .Z(n18445) );
  XOR U21475 ( .A(n18451), .B(n18452), .Z(n18079) );
  AND U21476 ( .A(n18453), .B(n18454), .Z(n18451) );
  AND U21477 ( .A(b[14]), .B(a[64]), .Z(n18450) );
  XOR U21478 ( .A(n18456), .B(n18457), .Z(n18084) );
  AND U21479 ( .A(n18458), .B(n18459), .Z(n18456) );
  AND U21480 ( .A(b[13]), .B(a[65]), .Z(n18455) );
  XOR U21481 ( .A(n18461), .B(n18462), .Z(n18089) );
  AND U21482 ( .A(n18463), .B(n18464), .Z(n18461) );
  AND U21483 ( .A(b[12]), .B(a[66]), .Z(n18460) );
  XOR U21484 ( .A(n18466), .B(n18467), .Z(n18094) );
  AND U21485 ( .A(n18468), .B(n18469), .Z(n18466) );
  AND U21486 ( .A(b[11]), .B(a[67]), .Z(n18465) );
  XOR U21487 ( .A(n18471), .B(n18472), .Z(n18099) );
  AND U21488 ( .A(n18473), .B(n18474), .Z(n18471) );
  AND U21489 ( .A(b[10]), .B(a[68]), .Z(n18470) );
  XOR U21490 ( .A(n18476), .B(n18477), .Z(n18104) );
  AND U21491 ( .A(n18478), .B(n18479), .Z(n18476) );
  AND U21492 ( .A(b[9]), .B(a[69]), .Z(n18475) );
  XOR U21493 ( .A(n18481), .B(n18482), .Z(n18109) );
  AND U21494 ( .A(n18483), .B(n18484), .Z(n18481) );
  AND U21495 ( .A(b[8]), .B(a[70]), .Z(n18480) );
  XOR U21496 ( .A(n18486), .B(n18487), .Z(n18114) );
  AND U21497 ( .A(n18488), .B(n18489), .Z(n18486) );
  AND U21498 ( .A(b[7]), .B(a[71]), .Z(n18485) );
  XOR U21499 ( .A(n18491), .B(n18492), .Z(n18119) );
  AND U21500 ( .A(n18493), .B(n18494), .Z(n18491) );
  AND U21501 ( .A(b[6]), .B(a[72]), .Z(n18490) );
  XOR U21502 ( .A(n18496), .B(n18497), .Z(n18124) );
  AND U21503 ( .A(n18498), .B(n18499), .Z(n18496) );
  AND U21504 ( .A(b[5]), .B(a[73]), .Z(n18495) );
  XOR U21505 ( .A(n18501), .B(n18502), .Z(n18129) );
  AND U21506 ( .A(n18503), .B(n18504), .Z(n18501) );
  AND U21507 ( .A(b[4]), .B(a[74]), .Z(n18500) );
  XOR U21508 ( .A(n18506), .B(n18507), .Z(n18134) );
  AND U21509 ( .A(n18508), .B(n18509), .Z(n18506) );
  AND U21510 ( .A(b[3]), .B(a[75]), .Z(n18505) );
  XOR U21511 ( .A(n18511), .B(n18512), .Z(n18139) );
  OR U21512 ( .A(n18513), .B(n18514), .Z(n18512) );
  AND U21513 ( .A(b[2]), .B(a[76]), .Z(n18510) );
  XNOR U21514 ( .A(n18149), .B(n18515), .Z(n18145) );
  NAND U21515 ( .A(b[1]), .B(a[77]), .Z(n18515) );
  IV U21516 ( .A(n18143), .Z(n18149) );
  ANDN U21517 ( .B(n10320), .A(n10322), .Z(n18143) );
  NAND U21518 ( .A(a[77]), .B(b[0]), .Z(n10322) );
  XOR U21519 ( .A(n18513), .B(n18514), .Z(n10320) );
  XOR U21520 ( .A(n18517), .B(n18508), .Z(n18516) );
  XOR U21521 ( .A(n18503), .B(n18507), .Z(n18518) );
  XOR U21522 ( .A(n18498), .B(n18502), .Z(n18519) );
  XOR U21523 ( .A(n18493), .B(n18497), .Z(n18520) );
  XOR U21524 ( .A(n18488), .B(n18492), .Z(n18521) );
  XOR U21525 ( .A(n18483), .B(n18487), .Z(n18522) );
  XOR U21526 ( .A(n18478), .B(n18482), .Z(n18523) );
  XOR U21527 ( .A(n18473), .B(n18477), .Z(n18524) );
  XOR U21528 ( .A(n18468), .B(n18472), .Z(n18525) );
  XOR U21529 ( .A(n18463), .B(n18467), .Z(n18526) );
  XOR U21530 ( .A(n18458), .B(n18462), .Z(n18527) );
  XOR U21531 ( .A(n18453), .B(n18457), .Z(n18528) );
  XOR U21532 ( .A(n18448), .B(n18452), .Z(n18529) );
  XOR U21533 ( .A(n18443), .B(n18447), .Z(n18530) );
  XOR U21534 ( .A(n18438), .B(n18442), .Z(n18531) );
  XOR U21535 ( .A(n18433), .B(n18437), .Z(n18532) );
  XOR U21536 ( .A(n18428), .B(n18432), .Z(n18533) );
  XOR U21537 ( .A(n18423), .B(n18427), .Z(n18534) );
  XOR U21538 ( .A(n18418), .B(n18422), .Z(n18535) );
  XOR U21539 ( .A(n18413), .B(n18417), .Z(n18536) );
  XOR U21540 ( .A(n18408), .B(n18412), .Z(n18537) );
  XOR U21541 ( .A(n18403), .B(n18407), .Z(n18538) );
  XOR U21542 ( .A(n18398), .B(n18402), .Z(n18539) );
  XOR U21543 ( .A(n18393), .B(n18397), .Z(n18540) );
  XOR U21544 ( .A(n18388), .B(n18392), .Z(n18541) );
  XOR U21545 ( .A(n18383), .B(n18387), .Z(n18542) );
  XOR U21546 ( .A(n18378), .B(n18382), .Z(n18543) );
  XOR U21547 ( .A(n18373), .B(n18377), .Z(n18544) );
  XOR U21548 ( .A(n18368), .B(n18372), .Z(n18545) );
  XOR U21549 ( .A(n18363), .B(n18367), .Z(n18546) );
  XOR U21550 ( .A(n18358), .B(n18362), .Z(n18547) );
  XOR U21551 ( .A(n18353), .B(n18357), .Z(n18548) );
  XOR U21552 ( .A(n18348), .B(n18352), .Z(n18549) );
  XOR U21553 ( .A(n18343), .B(n18347), .Z(n18550) );
  XOR U21554 ( .A(n18338), .B(n18342), .Z(n18551) );
  XOR U21555 ( .A(n18333), .B(n18337), .Z(n18552) );
  XOR U21556 ( .A(n18328), .B(n18332), .Z(n18553) );
  XOR U21557 ( .A(n18323), .B(n18327), .Z(n18554) );
  XOR U21558 ( .A(n18318), .B(n18322), .Z(n18555) );
  XOR U21559 ( .A(n18308), .B(n18317), .Z(n18556) );
  XOR U21560 ( .A(n18557), .B(n18307), .Z(n18308) );
  AND U21561 ( .A(a[36]), .B(b[41]), .Z(n18557) );
  XNOR U21562 ( .A(n18307), .B(n18313), .Z(n18558) );
  XNOR U21563 ( .A(n18312), .B(n18304), .Z(n18559) );
  XNOR U21564 ( .A(n18303), .B(n18299), .Z(n18560) );
  XNOR U21565 ( .A(n18298), .B(n18294), .Z(n18561) );
  XNOR U21566 ( .A(n18293), .B(n18289), .Z(n18562) );
  XNOR U21567 ( .A(n18288), .B(n18284), .Z(n18563) );
  XNOR U21568 ( .A(n18283), .B(n18279), .Z(n18564) );
  XNOR U21569 ( .A(n18278), .B(n18274), .Z(n18565) );
  XNOR U21570 ( .A(n18273), .B(n18269), .Z(n18566) );
  XNOR U21571 ( .A(n18268), .B(n18264), .Z(n18567) );
  XNOR U21572 ( .A(n18263), .B(n18259), .Z(n18568) );
  XNOR U21573 ( .A(n18258), .B(n18254), .Z(n18569) );
  XNOR U21574 ( .A(n18253), .B(n18249), .Z(n18570) );
  XNOR U21575 ( .A(n18248), .B(n18244), .Z(n18571) );
  XNOR U21576 ( .A(n18243), .B(n18239), .Z(n18572) );
  XNOR U21577 ( .A(n18238), .B(n18234), .Z(n18573) );
  XNOR U21578 ( .A(n18233), .B(n18229), .Z(n18574) );
  XNOR U21579 ( .A(n18228), .B(n18224), .Z(n18575) );
  XOR U21580 ( .A(n18223), .B(n18220), .Z(n18576) );
  XOR U21581 ( .A(n18577), .B(n18578), .Z(n18220) );
  XOR U21582 ( .A(n18218), .B(n18579), .Z(n18578) );
  XOR U21583 ( .A(n18580), .B(n18581), .Z(n18579) );
  XOR U21584 ( .A(n18582), .B(n18583), .Z(n18581) );
  NAND U21585 ( .A(a[15]), .B(b[62]), .Z(n18583) );
  AND U21586 ( .A(a[14]), .B(b[63]), .Z(n18582) );
  XOR U21587 ( .A(n18584), .B(n18580), .Z(n18577) );
  XOR U21588 ( .A(n18585), .B(n18586), .Z(n18580) );
  ANDN U21589 ( .B(n18587), .A(n18588), .Z(n18585) );
  AND U21590 ( .A(a[16]), .B(b[61]), .Z(n18584) );
  XOR U21591 ( .A(n18589), .B(n18218), .Z(n18219) );
  XOR U21592 ( .A(n18590), .B(n18591), .Z(n18218) );
  AND U21593 ( .A(n18592), .B(n18593), .Z(n18590) );
  AND U21594 ( .A(a[17]), .B(b[60]), .Z(n18589) );
  XOR U21595 ( .A(n18594), .B(n18223), .Z(n18225) );
  XOR U21596 ( .A(n18595), .B(n18596), .Z(n18223) );
  AND U21597 ( .A(n18597), .B(n18598), .Z(n18595) );
  AND U21598 ( .A(a[18]), .B(b[59]), .Z(n18594) );
  XOR U21599 ( .A(n18599), .B(n18228), .Z(n18230) );
  XOR U21600 ( .A(n18600), .B(n18601), .Z(n18228) );
  AND U21601 ( .A(n18602), .B(n18603), .Z(n18600) );
  AND U21602 ( .A(a[19]), .B(b[58]), .Z(n18599) );
  XOR U21603 ( .A(n18604), .B(n18233), .Z(n18235) );
  XOR U21604 ( .A(n18605), .B(n18606), .Z(n18233) );
  AND U21605 ( .A(n18607), .B(n18608), .Z(n18605) );
  AND U21606 ( .A(a[20]), .B(b[57]), .Z(n18604) );
  XOR U21607 ( .A(n18609), .B(n18238), .Z(n18240) );
  XOR U21608 ( .A(n18610), .B(n18611), .Z(n18238) );
  AND U21609 ( .A(n18612), .B(n18613), .Z(n18610) );
  AND U21610 ( .A(a[21]), .B(b[56]), .Z(n18609) );
  XOR U21611 ( .A(n18614), .B(n18243), .Z(n18245) );
  XOR U21612 ( .A(n18615), .B(n18616), .Z(n18243) );
  AND U21613 ( .A(n18617), .B(n18618), .Z(n18615) );
  AND U21614 ( .A(a[22]), .B(b[55]), .Z(n18614) );
  XOR U21615 ( .A(n18619), .B(n18248), .Z(n18250) );
  XOR U21616 ( .A(n18620), .B(n18621), .Z(n18248) );
  AND U21617 ( .A(n18622), .B(n18623), .Z(n18620) );
  AND U21618 ( .A(a[23]), .B(b[54]), .Z(n18619) );
  XOR U21619 ( .A(n18624), .B(n18253), .Z(n18255) );
  XOR U21620 ( .A(n18625), .B(n18626), .Z(n18253) );
  AND U21621 ( .A(n18627), .B(n18628), .Z(n18625) );
  AND U21622 ( .A(a[24]), .B(b[53]), .Z(n18624) );
  XOR U21623 ( .A(n18629), .B(n18258), .Z(n18260) );
  XOR U21624 ( .A(n18630), .B(n18631), .Z(n18258) );
  AND U21625 ( .A(n18632), .B(n18633), .Z(n18630) );
  AND U21626 ( .A(a[25]), .B(b[52]), .Z(n18629) );
  XOR U21627 ( .A(n18634), .B(n18263), .Z(n18265) );
  XOR U21628 ( .A(n18635), .B(n18636), .Z(n18263) );
  AND U21629 ( .A(n18637), .B(n18638), .Z(n18635) );
  AND U21630 ( .A(a[26]), .B(b[51]), .Z(n18634) );
  XOR U21631 ( .A(n18639), .B(n18268), .Z(n18270) );
  XOR U21632 ( .A(n18640), .B(n18641), .Z(n18268) );
  AND U21633 ( .A(n18642), .B(n18643), .Z(n18640) );
  AND U21634 ( .A(a[27]), .B(b[50]), .Z(n18639) );
  XOR U21635 ( .A(n18644), .B(n18273), .Z(n18275) );
  XOR U21636 ( .A(n18645), .B(n18646), .Z(n18273) );
  AND U21637 ( .A(n18647), .B(n18648), .Z(n18645) );
  AND U21638 ( .A(a[28]), .B(b[49]), .Z(n18644) );
  XOR U21639 ( .A(n18649), .B(n18278), .Z(n18280) );
  XOR U21640 ( .A(n18650), .B(n18651), .Z(n18278) );
  AND U21641 ( .A(n18652), .B(n18653), .Z(n18650) );
  AND U21642 ( .A(a[29]), .B(b[48]), .Z(n18649) );
  XOR U21643 ( .A(n18654), .B(n18283), .Z(n18285) );
  XOR U21644 ( .A(n18655), .B(n18656), .Z(n18283) );
  AND U21645 ( .A(n18657), .B(n18658), .Z(n18655) );
  AND U21646 ( .A(a[30]), .B(b[47]), .Z(n18654) );
  XOR U21647 ( .A(n18659), .B(n18288), .Z(n18290) );
  XOR U21648 ( .A(n18660), .B(n18661), .Z(n18288) );
  AND U21649 ( .A(n18662), .B(n18663), .Z(n18660) );
  AND U21650 ( .A(a[31]), .B(b[46]), .Z(n18659) );
  XOR U21651 ( .A(n18664), .B(n18293), .Z(n18295) );
  XOR U21652 ( .A(n18665), .B(n18666), .Z(n18293) );
  AND U21653 ( .A(n18667), .B(n18668), .Z(n18665) );
  AND U21654 ( .A(a[32]), .B(b[45]), .Z(n18664) );
  XOR U21655 ( .A(n18669), .B(n18298), .Z(n18300) );
  XOR U21656 ( .A(n18670), .B(n18671), .Z(n18298) );
  AND U21657 ( .A(n18672), .B(n18673), .Z(n18670) );
  AND U21658 ( .A(a[33]), .B(b[44]), .Z(n18669) );
  XOR U21659 ( .A(n18674), .B(n18303), .Z(n18305) );
  XOR U21660 ( .A(n18675), .B(n18676), .Z(n18303) );
  AND U21661 ( .A(n18677), .B(n18678), .Z(n18675) );
  AND U21662 ( .A(a[34]), .B(b[43]), .Z(n18674) );
  XOR U21663 ( .A(n18679), .B(n18680), .Z(n18307) );
  AND U21664 ( .A(n18681), .B(n18682), .Z(n18679) );
  XOR U21665 ( .A(n18683), .B(n18312), .Z(n18314) );
  XOR U21666 ( .A(n18684), .B(n18685), .Z(n18312) );
  AND U21667 ( .A(n18686), .B(n18687), .Z(n18684) );
  AND U21668 ( .A(a[35]), .B(b[42]), .Z(n18683) );
  XOR U21669 ( .A(n18689), .B(n18690), .Z(n18317) );
  AND U21670 ( .A(n18691), .B(n18692), .Z(n18689) );
  AND U21671 ( .A(a[37]), .B(b[40]), .Z(n18688) );
  XOR U21672 ( .A(n18694), .B(n18695), .Z(n18322) );
  AND U21673 ( .A(n18696), .B(n18697), .Z(n18694) );
  AND U21674 ( .A(a[38]), .B(b[39]), .Z(n18693) );
  XOR U21675 ( .A(n18699), .B(n18700), .Z(n18327) );
  AND U21676 ( .A(n18701), .B(n18702), .Z(n18699) );
  AND U21677 ( .A(b[38]), .B(a[39]), .Z(n18698) );
  XOR U21678 ( .A(n18704), .B(n18705), .Z(n18332) );
  AND U21679 ( .A(n18706), .B(n18707), .Z(n18704) );
  AND U21680 ( .A(b[37]), .B(a[40]), .Z(n18703) );
  XOR U21681 ( .A(n18709), .B(n18710), .Z(n18337) );
  AND U21682 ( .A(n18711), .B(n18712), .Z(n18709) );
  AND U21683 ( .A(b[36]), .B(a[41]), .Z(n18708) );
  XOR U21684 ( .A(n18714), .B(n18715), .Z(n18342) );
  AND U21685 ( .A(n18716), .B(n18717), .Z(n18714) );
  AND U21686 ( .A(b[35]), .B(a[42]), .Z(n18713) );
  XOR U21687 ( .A(n18719), .B(n18720), .Z(n18347) );
  AND U21688 ( .A(n18721), .B(n18722), .Z(n18719) );
  AND U21689 ( .A(b[34]), .B(a[43]), .Z(n18718) );
  XOR U21690 ( .A(n18724), .B(n18725), .Z(n18352) );
  AND U21691 ( .A(n18726), .B(n18727), .Z(n18724) );
  AND U21692 ( .A(b[33]), .B(a[44]), .Z(n18723) );
  XOR U21693 ( .A(n18729), .B(n18730), .Z(n18357) );
  AND U21694 ( .A(n18731), .B(n18732), .Z(n18729) );
  AND U21695 ( .A(b[32]), .B(a[45]), .Z(n18728) );
  XOR U21696 ( .A(n18734), .B(n18735), .Z(n18362) );
  AND U21697 ( .A(n18736), .B(n18737), .Z(n18734) );
  AND U21698 ( .A(b[31]), .B(a[46]), .Z(n18733) );
  XOR U21699 ( .A(n18739), .B(n18740), .Z(n18367) );
  AND U21700 ( .A(n18741), .B(n18742), .Z(n18739) );
  AND U21701 ( .A(b[30]), .B(a[47]), .Z(n18738) );
  XOR U21702 ( .A(n18744), .B(n18745), .Z(n18372) );
  AND U21703 ( .A(n18746), .B(n18747), .Z(n18744) );
  AND U21704 ( .A(b[29]), .B(a[48]), .Z(n18743) );
  XOR U21705 ( .A(n18749), .B(n18750), .Z(n18377) );
  AND U21706 ( .A(n18751), .B(n18752), .Z(n18749) );
  AND U21707 ( .A(b[28]), .B(a[49]), .Z(n18748) );
  XOR U21708 ( .A(n18754), .B(n18755), .Z(n18382) );
  AND U21709 ( .A(n18756), .B(n18757), .Z(n18754) );
  AND U21710 ( .A(b[27]), .B(a[50]), .Z(n18753) );
  XOR U21711 ( .A(n18759), .B(n18760), .Z(n18387) );
  AND U21712 ( .A(n18761), .B(n18762), .Z(n18759) );
  AND U21713 ( .A(b[26]), .B(a[51]), .Z(n18758) );
  XOR U21714 ( .A(n18764), .B(n18765), .Z(n18392) );
  AND U21715 ( .A(n18766), .B(n18767), .Z(n18764) );
  AND U21716 ( .A(b[25]), .B(a[52]), .Z(n18763) );
  XOR U21717 ( .A(n18769), .B(n18770), .Z(n18397) );
  AND U21718 ( .A(n18771), .B(n18772), .Z(n18769) );
  AND U21719 ( .A(b[24]), .B(a[53]), .Z(n18768) );
  XOR U21720 ( .A(n18774), .B(n18775), .Z(n18402) );
  AND U21721 ( .A(n18776), .B(n18777), .Z(n18774) );
  AND U21722 ( .A(b[23]), .B(a[54]), .Z(n18773) );
  XOR U21723 ( .A(n18779), .B(n18780), .Z(n18407) );
  AND U21724 ( .A(n18781), .B(n18782), .Z(n18779) );
  AND U21725 ( .A(b[22]), .B(a[55]), .Z(n18778) );
  XOR U21726 ( .A(n18784), .B(n18785), .Z(n18412) );
  AND U21727 ( .A(n18786), .B(n18787), .Z(n18784) );
  AND U21728 ( .A(b[21]), .B(a[56]), .Z(n18783) );
  XOR U21729 ( .A(n18789), .B(n18790), .Z(n18417) );
  AND U21730 ( .A(n18791), .B(n18792), .Z(n18789) );
  AND U21731 ( .A(b[20]), .B(a[57]), .Z(n18788) );
  XOR U21732 ( .A(n18794), .B(n18795), .Z(n18422) );
  AND U21733 ( .A(n18796), .B(n18797), .Z(n18794) );
  AND U21734 ( .A(b[19]), .B(a[58]), .Z(n18793) );
  XOR U21735 ( .A(n18799), .B(n18800), .Z(n18427) );
  AND U21736 ( .A(n18801), .B(n18802), .Z(n18799) );
  AND U21737 ( .A(b[18]), .B(a[59]), .Z(n18798) );
  XOR U21738 ( .A(n18804), .B(n18805), .Z(n18432) );
  AND U21739 ( .A(n18806), .B(n18807), .Z(n18804) );
  AND U21740 ( .A(b[17]), .B(a[60]), .Z(n18803) );
  XOR U21741 ( .A(n18809), .B(n18810), .Z(n18437) );
  AND U21742 ( .A(n18811), .B(n18812), .Z(n18809) );
  AND U21743 ( .A(b[16]), .B(a[61]), .Z(n18808) );
  XOR U21744 ( .A(n18814), .B(n18815), .Z(n18442) );
  AND U21745 ( .A(n18816), .B(n18817), .Z(n18814) );
  AND U21746 ( .A(b[15]), .B(a[62]), .Z(n18813) );
  XOR U21747 ( .A(n18819), .B(n18820), .Z(n18447) );
  AND U21748 ( .A(n18821), .B(n18822), .Z(n18819) );
  AND U21749 ( .A(b[14]), .B(a[63]), .Z(n18818) );
  XOR U21750 ( .A(n18824), .B(n18825), .Z(n18452) );
  AND U21751 ( .A(n18826), .B(n18827), .Z(n18824) );
  AND U21752 ( .A(b[13]), .B(a[64]), .Z(n18823) );
  XOR U21753 ( .A(n18829), .B(n18830), .Z(n18457) );
  AND U21754 ( .A(n18831), .B(n18832), .Z(n18829) );
  AND U21755 ( .A(b[12]), .B(a[65]), .Z(n18828) );
  XOR U21756 ( .A(n18834), .B(n18835), .Z(n18462) );
  AND U21757 ( .A(n18836), .B(n18837), .Z(n18834) );
  AND U21758 ( .A(b[11]), .B(a[66]), .Z(n18833) );
  XOR U21759 ( .A(n18839), .B(n18840), .Z(n18467) );
  AND U21760 ( .A(n18841), .B(n18842), .Z(n18839) );
  AND U21761 ( .A(b[10]), .B(a[67]), .Z(n18838) );
  XOR U21762 ( .A(n18844), .B(n18845), .Z(n18472) );
  AND U21763 ( .A(n18846), .B(n18847), .Z(n18844) );
  AND U21764 ( .A(b[9]), .B(a[68]), .Z(n18843) );
  XOR U21765 ( .A(n18849), .B(n18850), .Z(n18477) );
  AND U21766 ( .A(n18851), .B(n18852), .Z(n18849) );
  AND U21767 ( .A(b[8]), .B(a[69]), .Z(n18848) );
  XOR U21768 ( .A(n18854), .B(n18855), .Z(n18482) );
  AND U21769 ( .A(n18856), .B(n18857), .Z(n18854) );
  AND U21770 ( .A(b[7]), .B(a[70]), .Z(n18853) );
  XOR U21771 ( .A(n18859), .B(n18860), .Z(n18487) );
  AND U21772 ( .A(n18861), .B(n18862), .Z(n18859) );
  AND U21773 ( .A(b[6]), .B(a[71]), .Z(n18858) );
  XOR U21774 ( .A(n18864), .B(n18865), .Z(n18492) );
  AND U21775 ( .A(n18866), .B(n18867), .Z(n18864) );
  AND U21776 ( .A(b[5]), .B(a[72]), .Z(n18863) );
  XOR U21777 ( .A(n18869), .B(n18870), .Z(n18497) );
  AND U21778 ( .A(n18871), .B(n18872), .Z(n18869) );
  AND U21779 ( .A(b[4]), .B(a[73]), .Z(n18868) );
  XOR U21780 ( .A(n18874), .B(n18875), .Z(n18502) );
  AND U21781 ( .A(n18876), .B(n18877), .Z(n18874) );
  AND U21782 ( .A(b[3]), .B(a[74]), .Z(n18873) );
  XOR U21783 ( .A(n18879), .B(n18880), .Z(n18507) );
  OR U21784 ( .A(n18881), .B(n18882), .Z(n18880) );
  AND U21785 ( .A(b[2]), .B(a[75]), .Z(n18878) );
  XNOR U21786 ( .A(n18517), .B(n18883), .Z(n18513) );
  NAND U21787 ( .A(b[1]), .B(a[76]), .Z(n18883) );
  IV U21788 ( .A(n18511), .Z(n18517) );
  ANDN U21789 ( .B(n10323), .A(n10325), .Z(n18511) );
  NAND U21790 ( .A(a[76]), .B(b[0]), .Z(n10325) );
  XOR U21791 ( .A(n18881), .B(n18882), .Z(n10323) );
  XOR U21792 ( .A(n18885), .B(n18876), .Z(n18884) );
  XOR U21793 ( .A(n18871), .B(n18875), .Z(n18886) );
  XOR U21794 ( .A(n18866), .B(n18870), .Z(n18887) );
  XOR U21795 ( .A(n18861), .B(n18865), .Z(n18888) );
  XOR U21796 ( .A(n18856), .B(n18860), .Z(n18889) );
  XOR U21797 ( .A(n18851), .B(n18855), .Z(n18890) );
  XOR U21798 ( .A(n18846), .B(n18850), .Z(n18891) );
  XOR U21799 ( .A(n18841), .B(n18845), .Z(n18892) );
  XOR U21800 ( .A(n18836), .B(n18840), .Z(n18893) );
  XOR U21801 ( .A(n18831), .B(n18835), .Z(n18894) );
  XOR U21802 ( .A(n18826), .B(n18830), .Z(n18895) );
  XOR U21803 ( .A(n18821), .B(n18825), .Z(n18896) );
  XOR U21804 ( .A(n18816), .B(n18820), .Z(n18897) );
  XOR U21805 ( .A(n18811), .B(n18815), .Z(n18898) );
  XOR U21806 ( .A(n18806), .B(n18810), .Z(n18899) );
  XOR U21807 ( .A(n18801), .B(n18805), .Z(n18900) );
  XOR U21808 ( .A(n18796), .B(n18800), .Z(n18901) );
  XOR U21809 ( .A(n18791), .B(n18795), .Z(n18902) );
  XOR U21810 ( .A(n18786), .B(n18790), .Z(n18903) );
  XOR U21811 ( .A(n18781), .B(n18785), .Z(n18904) );
  XOR U21812 ( .A(n18776), .B(n18780), .Z(n18905) );
  XOR U21813 ( .A(n18771), .B(n18775), .Z(n18906) );
  XOR U21814 ( .A(n18766), .B(n18770), .Z(n18907) );
  XOR U21815 ( .A(n18761), .B(n18765), .Z(n18908) );
  XOR U21816 ( .A(n18756), .B(n18760), .Z(n18909) );
  XOR U21817 ( .A(n18751), .B(n18755), .Z(n18910) );
  XOR U21818 ( .A(n18746), .B(n18750), .Z(n18911) );
  XOR U21819 ( .A(n18741), .B(n18745), .Z(n18912) );
  XOR U21820 ( .A(n18736), .B(n18740), .Z(n18913) );
  XOR U21821 ( .A(n18731), .B(n18735), .Z(n18914) );
  XOR U21822 ( .A(n18726), .B(n18730), .Z(n18915) );
  XOR U21823 ( .A(n18721), .B(n18725), .Z(n18916) );
  XOR U21824 ( .A(n18716), .B(n18720), .Z(n18917) );
  XOR U21825 ( .A(n18711), .B(n18715), .Z(n18918) );
  XOR U21826 ( .A(n18706), .B(n18710), .Z(n18919) );
  XOR U21827 ( .A(n18701), .B(n18705), .Z(n18920) );
  XOR U21828 ( .A(n18696), .B(n18700), .Z(n18921) );
  XOR U21829 ( .A(n18691), .B(n18695), .Z(n18922) );
  XOR U21830 ( .A(n18681), .B(n18690), .Z(n18923) );
  XOR U21831 ( .A(n18924), .B(n18680), .Z(n18681) );
  AND U21832 ( .A(a[36]), .B(b[40]), .Z(n18924) );
  XNOR U21833 ( .A(n18680), .B(n18686), .Z(n18925) );
  XNOR U21834 ( .A(n18685), .B(n18677), .Z(n18926) );
  XNOR U21835 ( .A(n18676), .B(n18672), .Z(n18927) );
  XNOR U21836 ( .A(n18671), .B(n18667), .Z(n18928) );
  XNOR U21837 ( .A(n18666), .B(n18662), .Z(n18929) );
  XNOR U21838 ( .A(n18661), .B(n18657), .Z(n18930) );
  XNOR U21839 ( .A(n18656), .B(n18652), .Z(n18931) );
  XNOR U21840 ( .A(n18651), .B(n18647), .Z(n18932) );
  XNOR U21841 ( .A(n18646), .B(n18642), .Z(n18933) );
  XNOR U21842 ( .A(n18641), .B(n18637), .Z(n18934) );
  XNOR U21843 ( .A(n18636), .B(n18632), .Z(n18935) );
  XNOR U21844 ( .A(n18631), .B(n18627), .Z(n18936) );
  XNOR U21845 ( .A(n18626), .B(n18622), .Z(n18937) );
  XNOR U21846 ( .A(n18621), .B(n18617), .Z(n18938) );
  XNOR U21847 ( .A(n18616), .B(n18612), .Z(n18939) );
  XNOR U21848 ( .A(n18611), .B(n18607), .Z(n18940) );
  XNOR U21849 ( .A(n18606), .B(n18602), .Z(n18941) );
  XNOR U21850 ( .A(n18601), .B(n18597), .Z(n18942) );
  XNOR U21851 ( .A(n18596), .B(n18592), .Z(n18943) );
  XOR U21852 ( .A(n18591), .B(n18588), .Z(n18944) );
  XOR U21853 ( .A(n18945), .B(n18946), .Z(n18588) );
  XOR U21854 ( .A(n18586), .B(n18947), .Z(n18946) );
  XOR U21855 ( .A(n18948), .B(n18949), .Z(n18947) );
  XOR U21856 ( .A(n18950), .B(n18951), .Z(n18949) );
  NAND U21857 ( .A(a[14]), .B(b[62]), .Z(n18951) );
  AND U21858 ( .A(a[13]), .B(b[63]), .Z(n18950) );
  XOR U21859 ( .A(n18952), .B(n18948), .Z(n18945) );
  XOR U21860 ( .A(n18953), .B(n18954), .Z(n18948) );
  ANDN U21861 ( .B(n18955), .A(n18956), .Z(n18953) );
  AND U21862 ( .A(a[15]), .B(b[61]), .Z(n18952) );
  XOR U21863 ( .A(n18957), .B(n18586), .Z(n18587) );
  XOR U21864 ( .A(n18958), .B(n18959), .Z(n18586) );
  AND U21865 ( .A(n18960), .B(n18961), .Z(n18958) );
  AND U21866 ( .A(a[16]), .B(b[60]), .Z(n18957) );
  XOR U21867 ( .A(n18962), .B(n18591), .Z(n18593) );
  XOR U21868 ( .A(n18963), .B(n18964), .Z(n18591) );
  AND U21869 ( .A(n18965), .B(n18966), .Z(n18963) );
  AND U21870 ( .A(a[17]), .B(b[59]), .Z(n18962) );
  XOR U21871 ( .A(n18967), .B(n18596), .Z(n18598) );
  XOR U21872 ( .A(n18968), .B(n18969), .Z(n18596) );
  AND U21873 ( .A(n18970), .B(n18971), .Z(n18968) );
  AND U21874 ( .A(a[18]), .B(b[58]), .Z(n18967) );
  XOR U21875 ( .A(n18972), .B(n18601), .Z(n18603) );
  XOR U21876 ( .A(n18973), .B(n18974), .Z(n18601) );
  AND U21877 ( .A(n18975), .B(n18976), .Z(n18973) );
  AND U21878 ( .A(a[19]), .B(b[57]), .Z(n18972) );
  XOR U21879 ( .A(n18977), .B(n18606), .Z(n18608) );
  XOR U21880 ( .A(n18978), .B(n18979), .Z(n18606) );
  AND U21881 ( .A(n18980), .B(n18981), .Z(n18978) );
  AND U21882 ( .A(a[20]), .B(b[56]), .Z(n18977) );
  XOR U21883 ( .A(n18982), .B(n18611), .Z(n18613) );
  XOR U21884 ( .A(n18983), .B(n18984), .Z(n18611) );
  AND U21885 ( .A(n18985), .B(n18986), .Z(n18983) );
  AND U21886 ( .A(a[21]), .B(b[55]), .Z(n18982) );
  XOR U21887 ( .A(n18987), .B(n18616), .Z(n18618) );
  XOR U21888 ( .A(n18988), .B(n18989), .Z(n18616) );
  AND U21889 ( .A(n18990), .B(n18991), .Z(n18988) );
  AND U21890 ( .A(a[22]), .B(b[54]), .Z(n18987) );
  XOR U21891 ( .A(n18992), .B(n18621), .Z(n18623) );
  XOR U21892 ( .A(n18993), .B(n18994), .Z(n18621) );
  AND U21893 ( .A(n18995), .B(n18996), .Z(n18993) );
  AND U21894 ( .A(a[23]), .B(b[53]), .Z(n18992) );
  XOR U21895 ( .A(n18997), .B(n18626), .Z(n18628) );
  XOR U21896 ( .A(n18998), .B(n18999), .Z(n18626) );
  AND U21897 ( .A(n19000), .B(n19001), .Z(n18998) );
  AND U21898 ( .A(a[24]), .B(b[52]), .Z(n18997) );
  XOR U21899 ( .A(n19002), .B(n18631), .Z(n18633) );
  XOR U21900 ( .A(n19003), .B(n19004), .Z(n18631) );
  AND U21901 ( .A(n19005), .B(n19006), .Z(n19003) );
  AND U21902 ( .A(a[25]), .B(b[51]), .Z(n19002) );
  XOR U21903 ( .A(n19007), .B(n18636), .Z(n18638) );
  XOR U21904 ( .A(n19008), .B(n19009), .Z(n18636) );
  AND U21905 ( .A(n19010), .B(n19011), .Z(n19008) );
  AND U21906 ( .A(a[26]), .B(b[50]), .Z(n19007) );
  XOR U21907 ( .A(n19012), .B(n18641), .Z(n18643) );
  XOR U21908 ( .A(n19013), .B(n19014), .Z(n18641) );
  AND U21909 ( .A(n19015), .B(n19016), .Z(n19013) );
  AND U21910 ( .A(a[27]), .B(b[49]), .Z(n19012) );
  XOR U21911 ( .A(n19017), .B(n18646), .Z(n18648) );
  XOR U21912 ( .A(n19018), .B(n19019), .Z(n18646) );
  AND U21913 ( .A(n19020), .B(n19021), .Z(n19018) );
  AND U21914 ( .A(a[28]), .B(b[48]), .Z(n19017) );
  XOR U21915 ( .A(n19022), .B(n18651), .Z(n18653) );
  XOR U21916 ( .A(n19023), .B(n19024), .Z(n18651) );
  AND U21917 ( .A(n19025), .B(n19026), .Z(n19023) );
  AND U21918 ( .A(a[29]), .B(b[47]), .Z(n19022) );
  XOR U21919 ( .A(n19027), .B(n18656), .Z(n18658) );
  XOR U21920 ( .A(n19028), .B(n19029), .Z(n18656) );
  AND U21921 ( .A(n19030), .B(n19031), .Z(n19028) );
  AND U21922 ( .A(a[30]), .B(b[46]), .Z(n19027) );
  XOR U21923 ( .A(n19032), .B(n18661), .Z(n18663) );
  XOR U21924 ( .A(n19033), .B(n19034), .Z(n18661) );
  AND U21925 ( .A(n19035), .B(n19036), .Z(n19033) );
  AND U21926 ( .A(a[31]), .B(b[45]), .Z(n19032) );
  XOR U21927 ( .A(n19037), .B(n18666), .Z(n18668) );
  XOR U21928 ( .A(n19038), .B(n19039), .Z(n18666) );
  AND U21929 ( .A(n19040), .B(n19041), .Z(n19038) );
  AND U21930 ( .A(a[32]), .B(b[44]), .Z(n19037) );
  XOR U21931 ( .A(n19042), .B(n18671), .Z(n18673) );
  XOR U21932 ( .A(n19043), .B(n19044), .Z(n18671) );
  AND U21933 ( .A(n19045), .B(n19046), .Z(n19043) );
  AND U21934 ( .A(a[33]), .B(b[43]), .Z(n19042) );
  XOR U21935 ( .A(n19047), .B(n18676), .Z(n18678) );
  XOR U21936 ( .A(n19048), .B(n19049), .Z(n18676) );
  AND U21937 ( .A(n19050), .B(n19051), .Z(n19048) );
  AND U21938 ( .A(a[34]), .B(b[42]), .Z(n19047) );
  XOR U21939 ( .A(n19052), .B(n19053), .Z(n18680) );
  AND U21940 ( .A(n19054), .B(n19055), .Z(n19052) );
  XOR U21941 ( .A(n19056), .B(n18685), .Z(n18687) );
  XOR U21942 ( .A(n19057), .B(n19058), .Z(n18685) );
  AND U21943 ( .A(n19059), .B(n19060), .Z(n19057) );
  AND U21944 ( .A(a[35]), .B(b[41]), .Z(n19056) );
  XOR U21945 ( .A(n19062), .B(n19063), .Z(n18690) );
  AND U21946 ( .A(n19064), .B(n19065), .Z(n19062) );
  AND U21947 ( .A(a[37]), .B(b[39]), .Z(n19061) );
  XOR U21948 ( .A(n19067), .B(n19068), .Z(n18695) );
  AND U21949 ( .A(n19069), .B(n19070), .Z(n19067) );
  AND U21950 ( .A(a[38]), .B(b[38]), .Z(n19066) );
  XOR U21951 ( .A(n19072), .B(n19073), .Z(n18700) );
  AND U21952 ( .A(n19074), .B(n19075), .Z(n19072) );
  AND U21953 ( .A(b[37]), .B(a[39]), .Z(n19071) );
  XOR U21954 ( .A(n19077), .B(n19078), .Z(n18705) );
  AND U21955 ( .A(n19079), .B(n19080), .Z(n19077) );
  AND U21956 ( .A(b[36]), .B(a[40]), .Z(n19076) );
  XOR U21957 ( .A(n19082), .B(n19083), .Z(n18710) );
  AND U21958 ( .A(n19084), .B(n19085), .Z(n19082) );
  AND U21959 ( .A(b[35]), .B(a[41]), .Z(n19081) );
  XOR U21960 ( .A(n19087), .B(n19088), .Z(n18715) );
  AND U21961 ( .A(n19089), .B(n19090), .Z(n19087) );
  AND U21962 ( .A(b[34]), .B(a[42]), .Z(n19086) );
  XOR U21963 ( .A(n19092), .B(n19093), .Z(n18720) );
  AND U21964 ( .A(n19094), .B(n19095), .Z(n19092) );
  AND U21965 ( .A(b[33]), .B(a[43]), .Z(n19091) );
  XOR U21966 ( .A(n19097), .B(n19098), .Z(n18725) );
  AND U21967 ( .A(n19099), .B(n19100), .Z(n19097) );
  AND U21968 ( .A(b[32]), .B(a[44]), .Z(n19096) );
  XOR U21969 ( .A(n19102), .B(n19103), .Z(n18730) );
  AND U21970 ( .A(n19104), .B(n19105), .Z(n19102) );
  AND U21971 ( .A(b[31]), .B(a[45]), .Z(n19101) );
  XOR U21972 ( .A(n19107), .B(n19108), .Z(n18735) );
  AND U21973 ( .A(n19109), .B(n19110), .Z(n19107) );
  AND U21974 ( .A(b[30]), .B(a[46]), .Z(n19106) );
  XOR U21975 ( .A(n19112), .B(n19113), .Z(n18740) );
  AND U21976 ( .A(n19114), .B(n19115), .Z(n19112) );
  AND U21977 ( .A(b[29]), .B(a[47]), .Z(n19111) );
  XOR U21978 ( .A(n19117), .B(n19118), .Z(n18745) );
  AND U21979 ( .A(n19119), .B(n19120), .Z(n19117) );
  AND U21980 ( .A(b[28]), .B(a[48]), .Z(n19116) );
  XOR U21981 ( .A(n19122), .B(n19123), .Z(n18750) );
  AND U21982 ( .A(n19124), .B(n19125), .Z(n19122) );
  AND U21983 ( .A(b[27]), .B(a[49]), .Z(n19121) );
  XOR U21984 ( .A(n19127), .B(n19128), .Z(n18755) );
  AND U21985 ( .A(n19129), .B(n19130), .Z(n19127) );
  AND U21986 ( .A(b[26]), .B(a[50]), .Z(n19126) );
  XOR U21987 ( .A(n19132), .B(n19133), .Z(n18760) );
  AND U21988 ( .A(n19134), .B(n19135), .Z(n19132) );
  AND U21989 ( .A(b[25]), .B(a[51]), .Z(n19131) );
  XOR U21990 ( .A(n19137), .B(n19138), .Z(n18765) );
  AND U21991 ( .A(n19139), .B(n19140), .Z(n19137) );
  AND U21992 ( .A(b[24]), .B(a[52]), .Z(n19136) );
  XOR U21993 ( .A(n19142), .B(n19143), .Z(n18770) );
  AND U21994 ( .A(n19144), .B(n19145), .Z(n19142) );
  AND U21995 ( .A(b[23]), .B(a[53]), .Z(n19141) );
  XOR U21996 ( .A(n19147), .B(n19148), .Z(n18775) );
  AND U21997 ( .A(n19149), .B(n19150), .Z(n19147) );
  AND U21998 ( .A(b[22]), .B(a[54]), .Z(n19146) );
  XOR U21999 ( .A(n19152), .B(n19153), .Z(n18780) );
  AND U22000 ( .A(n19154), .B(n19155), .Z(n19152) );
  AND U22001 ( .A(b[21]), .B(a[55]), .Z(n19151) );
  XOR U22002 ( .A(n19157), .B(n19158), .Z(n18785) );
  AND U22003 ( .A(n19159), .B(n19160), .Z(n19157) );
  AND U22004 ( .A(b[20]), .B(a[56]), .Z(n19156) );
  XOR U22005 ( .A(n19162), .B(n19163), .Z(n18790) );
  AND U22006 ( .A(n19164), .B(n19165), .Z(n19162) );
  AND U22007 ( .A(b[19]), .B(a[57]), .Z(n19161) );
  XOR U22008 ( .A(n19167), .B(n19168), .Z(n18795) );
  AND U22009 ( .A(n19169), .B(n19170), .Z(n19167) );
  AND U22010 ( .A(b[18]), .B(a[58]), .Z(n19166) );
  XOR U22011 ( .A(n19172), .B(n19173), .Z(n18800) );
  AND U22012 ( .A(n19174), .B(n19175), .Z(n19172) );
  AND U22013 ( .A(b[17]), .B(a[59]), .Z(n19171) );
  XOR U22014 ( .A(n19177), .B(n19178), .Z(n18805) );
  AND U22015 ( .A(n19179), .B(n19180), .Z(n19177) );
  AND U22016 ( .A(b[16]), .B(a[60]), .Z(n19176) );
  XOR U22017 ( .A(n19182), .B(n19183), .Z(n18810) );
  AND U22018 ( .A(n19184), .B(n19185), .Z(n19182) );
  AND U22019 ( .A(b[15]), .B(a[61]), .Z(n19181) );
  XOR U22020 ( .A(n19187), .B(n19188), .Z(n18815) );
  AND U22021 ( .A(n19189), .B(n19190), .Z(n19187) );
  AND U22022 ( .A(b[14]), .B(a[62]), .Z(n19186) );
  XOR U22023 ( .A(n19192), .B(n19193), .Z(n18820) );
  AND U22024 ( .A(n19194), .B(n19195), .Z(n19192) );
  AND U22025 ( .A(b[13]), .B(a[63]), .Z(n19191) );
  XOR U22026 ( .A(n19197), .B(n19198), .Z(n18825) );
  AND U22027 ( .A(n19199), .B(n19200), .Z(n19197) );
  AND U22028 ( .A(b[12]), .B(a[64]), .Z(n19196) );
  XOR U22029 ( .A(n19202), .B(n19203), .Z(n18830) );
  AND U22030 ( .A(n19204), .B(n19205), .Z(n19202) );
  AND U22031 ( .A(b[11]), .B(a[65]), .Z(n19201) );
  XOR U22032 ( .A(n19207), .B(n19208), .Z(n18835) );
  AND U22033 ( .A(n19209), .B(n19210), .Z(n19207) );
  AND U22034 ( .A(b[10]), .B(a[66]), .Z(n19206) );
  XOR U22035 ( .A(n19212), .B(n19213), .Z(n18840) );
  AND U22036 ( .A(n19214), .B(n19215), .Z(n19212) );
  AND U22037 ( .A(b[9]), .B(a[67]), .Z(n19211) );
  XOR U22038 ( .A(n19217), .B(n19218), .Z(n18845) );
  AND U22039 ( .A(n19219), .B(n19220), .Z(n19217) );
  AND U22040 ( .A(b[8]), .B(a[68]), .Z(n19216) );
  XOR U22041 ( .A(n19222), .B(n19223), .Z(n18850) );
  AND U22042 ( .A(n19224), .B(n19225), .Z(n19222) );
  AND U22043 ( .A(b[7]), .B(a[69]), .Z(n19221) );
  XOR U22044 ( .A(n19227), .B(n19228), .Z(n18855) );
  AND U22045 ( .A(n19229), .B(n19230), .Z(n19227) );
  AND U22046 ( .A(b[6]), .B(a[70]), .Z(n19226) );
  XOR U22047 ( .A(n19232), .B(n19233), .Z(n18860) );
  AND U22048 ( .A(n19234), .B(n19235), .Z(n19232) );
  AND U22049 ( .A(b[5]), .B(a[71]), .Z(n19231) );
  XOR U22050 ( .A(n19237), .B(n19238), .Z(n18865) );
  AND U22051 ( .A(n19239), .B(n19240), .Z(n19237) );
  AND U22052 ( .A(b[4]), .B(a[72]), .Z(n19236) );
  XOR U22053 ( .A(n19242), .B(n19243), .Z(n18870) );
  AND U22054 ( .A(n19244), .B(n19245), .Z(n19242) );
  AND U22055 ( .A(b[3]), .B(a[73]), .Z(n19241) );
  XOR U22056 ( .A(n19247), .B(n19248), .Z(n18875) );
  OR U22057 ( .A(n19249), .B(n19250), .Z(n19248) );
  AND U22058 ( .A(b[2]), .B(a[74]), .Z(n19246) );
  XNOR U22059 ( .A(n18885), .B(n19251), .Z(n18881) );
  NAND U22060 ( .A(b[1]), .B(a[75]), .Z(n19251) );
  IV U22061 ( .A(n18879), .Z(n18885) );
  ANDN U22062 ( .B(n10326), .A(n10328), .Z(n18879) );
  NAND U22063 ( .A(a[75]), .B(b[0]), .Z(n10328) );
  XOR U22064 ( .A(n19249), .B(n19250), .Z(n10326) );
  XOR U22065 ( .A(n19253), .B(n19244), .Z(n19252) );
  XOR U22066 ( .A(n19239), .B(n19243), .Z(n19254) );
  XOR U22067 ( .A(n19234), .B(n19238), .Z(n19255) );
  XOR U22068 ( .A(n19229), .B(n19233), .Z(n19256) );
  XOR U22069 ( .A(n19224), .B(n19228), .Z(n19257) );
  XOR U22070 ( .A(n19219), .B(n19223), .Z(n19258) );
  XOR U22071 ( .A(n19214), .B(n19218), .Z(n19259) );
  XOR U22072 ( .A(n19209), .B(n19213), .Z(n19260) );
  XOR U22073 ( .A(n19204), .B(n19208), .Z(n19261) );
  XOR U22074 ( .A(n19199), .B(n19203), .Z(n19262) );
  XOR U22075 ( .A(n19194), .B(n19198), .Z(n19263) );
  XOR U22076 ( .A(n19189), .B(n19193), .Z(n19264) );
  XOR U22077 ( .A(n19184), .B(n19188), .Z(n19265) );
  XOR U22078 ( .A(n19179), .B(n19183), .Z(n19266) );
  XOR U22079 ( .A(n19174), .B(n19178), .Z(n19267) );
  XOR U22080 ( .A(n19169), .B(n19173), .Z(n19268) );
  XOR U22081 ( .A(n19164), .B(n19168), .Z(n19269) );
  XOR U22082 ( .A(n19159), .B(n19163), .Z(n19270) );
  XOR U22083 ( .A(n19154), .B(n19158), .Z(n19271) );
  XOR U22084 ( .A(n19149), .B(n19153), .Z(n19272) );
  XOR U22085 ( .A(n19144), .B(n19148), .Z(n19273) );
  XOR U22086 ( .A(n19139), .B(n19143), .Z(n19274) );
  XOR U22087 ( .A(n19134), .B(n19138), .Z(n19275) );
  XOR U22088 ( .A(n19129), .B(n19133), .Z(n19276) );
  XOR U22089 ( .A(n19124), .B(n19128), .Z(n19277) );
  XOR U22090 ( .A(n19119), .B(n19123), .Z(n19278) );
  XOR U22091 ( .A(n19114), .B(n19118), .Z(n19279) );
  XOR U22092 ( .A(n19109), .B(n19113), .Z(n19280) );
  XOR U22093 ( .A(n19104), .B(n19108), .Z(n19281) );
  XOR U22094 ( .A(n19099), .B(n19103), .Z(n19282) );
  XOR U22095 ( .A(n19094), .B(n19098), .Z(n19283) );
  XOR U22096 ( .A(n19089), .B(n19093), .Z(n19284) );
  XOR U22097 ( .A(n19084), .B(n19088), .Z(n19285) );
  XOR U22098 ( .A(n19079), .B(n19083), .Z(n19286) );
  XOR U22099 ( .A(n19074), .B(n19078), .Z(n19287) );
  XOR U22100 ( .A(n19069), .B(n19073), .Z(n19288) );
  XOR U22101 ( .A(n19064), .B(n19068), .Z(n19289) );
  XOR U22102 ( .A(n19054), .B(n19063), .Z(n19290) );
  XOR U22103 ( .A(n19291), .B(n19053), .Z(n19054) );
  AND U22104 ( .A(a[36]), .B(b[39]), .Z(n19291) );
  XNOR U22105 ( .A(n19053), .B(n19059), .Z(n19292) );
  XNOR U22106 ( .A(n19058), .B(n19050), .Z(n19293) );
  XNOR U22107 ( .A(n19049), .B(n19045), .Z(n19294) );
  XNOR U22108 ( .A(n19044), .B(n19040), .Z(n19295) );
  XNOR U22109 ( .A(n19039), .B(n19035), .Z(n19296) );
  XNOR U22110 ( .A(n19034), .B(n19030), .Z(n19297) );
  XNOR U22111 ( .A(n19029), .B(n19025), .Z(n19298) );
  XNOR U22112 ( .A(n19024), .B(n19020), .Z(n19299) );
  XNOR U22113 ( .A(n19019), .B(n19015), .Z(n19300) );
  XNOR U22114 ( .A(n19014), .B(n19010), .Z(n19301) );
  XNOR U22115 ( .A(n19009), .B(n19005), .Z(n19302) );
  XNOR U22116 ( .A(n19004), .B(n19000), .Z(n19303) );
  XNOR U22117 ( .A(n18999), .B(n18995), .Z(n19304) );
  XNOR U22118 ( .A(n18994), .B(n18990), .Z(n19305) );
  XNOR U22119 ( .A(n18989), .B(n18985), .Z(n19306) );
  XNOR U22120 ( .A(n18984), .B(n18980), .Z(n19307) );
  XNOR U22121 ( .A(n18979), .B(n18975), .Z(n19308) );
  XNOR U22122 ( .A(n18974), .B(n18970), .Z(n19309) );
  XNOR U22123 ( .A(n18969), .B(n18965), .Z(n19310) );
  XNOR U22124 ( .A(n18964), .B(n18960), .Z(n19311) );
  XOR U22125 ( .A(n18959), .B(n18956), .Z(n19312) );
  XOR U22126 ( .A(n19313), .B(n19314), .Z(n18956) );
  XOR U22127 ( .A(n18954), .B(n19315), .Z(n19314) );
  XOR U22128 ( .A(n19316), .B(n19317), .Z(n19315) );
  XOR U22129 ( .A(n19318), .B(n19319), .Z(n19317) );
  NAND U22130 ( .A(a[13]), .B(b[62]), .Z(n19319) );
  AND U22131 ( .A(a[12]), .B(b[63]), .Z(n19318) );
  XOR U22132 ( .A(n19320), .B(n19316), .Z(n19313) );
  XOR U22133 ( .A(n19321), .B(n19322), .Z(n19316) );
  ANDN U22134 ( .B(n19323), .A(n19324), .Z(n19321) );
  AND U22135 ( .A(a[14]), .B(b[61]), .Z(n19320) );
  XOR U22136 ( .A(n19325), .B(n18954), .Z(n18955) );
  XOR U22137 ( .A(n19326), .B(n19327), .Z(n18954) );
  AND U22138 ( .A(n19328), .B(n19329), .Z(n19326) );
  AND U22139 ( .A(a[15]), .B(b[60]), .Z(n19325) );
  XOR U22140 ( .A(n19330), .B(n18959), .Z(n18961) );
  XOR U22141 ( .A(n19331), .B(n19332), .Z(n18959) );
  AND U22142 ( .A(n19333), .B(n19334), .Z(n19331) );
  AND U22143 ( .A(a[16]), .B(b[59]), .Z(n19330) );
  XOR U22144 ( .A(n19335), .B(n18964), .Z(n18966) );
  XOR U22145 ( .A(n19336), .B(n19337), .Z(n18964) );
  AND U22146 ( .A(n19338), .B(n19339), .Z(n19336) );
  AND U22147 ( .A(a[17]), .B(b[58]), .Z(n19335) );
  XOR U22148 ( .A(n19340), .B(n18969), .Z(n18971) );
  XOR U22149 ( .A(n19341), .B(n19342), .Z(n18969) );
  AND U22150 ( .A(n19343), .B(n19344), .Z(n19341) );
  AND U22151 ( .A(a[18]), .B(b[57]), .Z(n19340) );
  XOR U22152 ( .A(n19345), .B(n18974), .Z(n18976) );
  XOR U22153 ( .A(n19346), .B(n19347), .Z(n18974) );
  AND U22154 ( .A(n19348), .B(n19349), .Z(n19346) );
  AND U22155 ( .A(a[19]), .B(b[56]), .Z(n19345) );
  XOR U22156 ( .A(n19350), .B(n18979), .Z(n18981) );
  XOR U22157 ( .A(n19351), .B(n19352), .Z(n18979) );
  AND U22158 ( .A(n19353), .B(n19354), .Z(n19351) );
  AND U22159 ( .A(a[20]), .B(b[55]), .Z(n19350) );
  XOR U22160 ( .A(n19355), .B(n18984), .Z(n18986) );
  XOR U22161 ( .A(n19356), .B(n19357), .Z(n18984) );
  AND U22162 ( .A(n19358), .B(n19359), .Z(n19356) );
  AND U22163 ( .A(a[21]), .B(b[54]), .Z(n19355) );
  XOR U22164 ( .A(n19360), .B(n18989), .Z(n18991) );
  XOR U22165 ( .A(n19361), .B(n19362), .Z(n18989) );
  AND U22166 ( .A(n19363), .B(n19364), .Z(n19361) );
  AND U22167 ( .A(a[22]), .B(b[53]), .Z(n19360) );
  XOR U22168 ( .A(n19365), .B(n18994), .Z(n18996) );
  XOR U22169 ( .A(n19366), .B(n19367), .Z(n18994) );
  AND U22170 ( .A(n19368), .B(n19369), .Z(n19366) );
  AND U22171 ( .A(a[23]), .B(b[52]), .Z(n19365) );
  XOR U22172 ( .A(n19370), .B(n18999), .Z(n19001) );
  XOR U22173 ( .A(n19371), .B(n19372), .Z(n18999) );
  AND U22174 ( .A(n19373), .B(n19374), .Z(n19371) );
  AND U22175 ( .A(a[24]), .B(b[51]), .Z(n19370) );
  XOR U22176 ( .A(n19375), .B(n19004), .Z(n19006) );
  XOR U22177 ( .A(n19376), .B(n19377), .Z(n19004) );
  AND U22178 ( .A(n19378), .B(n19379), .Z(n19376) );
  AND U22179 ( .A(a[25]), .B(b[50]), .Z(n19375) );
  XOR U22180 ( .A(n19380), .B(n19009), .Z(n19011) );
  XOR U22181 ( .A(n19381), .B(n19382), .Z(n19009) );
  AND U22182 ( .A(n19383), .B(n19384), .Z(n19381) );
  AND U22183 ( .A(a[26]), .B(b[49]), .Z(n19380) );
  XOR U22184 ( .A(n19385), .B(n19014), .Z(n19016) );
  XOR U22185 ( .A(n19386), .B(n19387), .Z(n19014) );
  AND U22186 ( .A(n19388), .B(n19389), .Z(n19386) );
  AND U22187 ( .A(a[27]), .B(b[48]), .Z(n19385) );
  XOR U22188 ( .A(n19390), .B(n19019), .Z(n19021) );
  XOR U22189 ( .A(n19391), .B(n19392), .Z(n19019) );
  AND U22190 ( .A(n19393), .B(n19394), .Z(n19391) );
  AND U22191 ( .A(a[28]), .B(b[47]), .Z(n19390) );
  XOR U22192 ( .A(n19395), .B(n19024), .Z(n19026) );
  XOR U22193 ( .A(n19396), .B(n19397), .Z(n19024) );
  AND U22194 ( .A(n19398), .B(n19399), .Z(n19396) );
  AND U22195 ( .A(a[29]), .B(b[46]), .Z(n19395) );
  XOR U22196 ( .A(n19400), .B(n19029), .Z(n19031) );
  XOR U22197 ( .A(n19401), .B(n19402), .Z(n19029) );
  AND U22198 ( .A(n19403), .B(n19404), .Z(n19401) );
  AND U22199 ( .A(a[30]), .B(b[45]), .Z(n19400) );
  XOR U22200 ( .A(n19405), .B(n19034), .Z(n19036) );
  XOR U22201 ( .A(n19406), .B(n19407), .Z(n19034) );
  AND U22202 ( .A(n19408), .B(n19409), .Z(n19406) );
  AND U22203 ( .A(a[31]), .B(b[44]), .Z(n19405) );
  XOR U22204 ( .A(n19410), .B(n19039), .Z(n19041) );
  XOR U22205 ( .A(n19411), .B(n19412), .Z(n19039) );
  AND U22206 ( .A(n19413), .B(n19414), .Z(n19411) );
  AND U22207 ( .A(a[32]), .B(b[43]), .Z(n19410) );
  XOR U22208 ( .A(n19415), .B(n19044), .Z(n19046) );
  XOR U22209 ( .A(n19416), .B(n19417), .Z(n19044) );
  AND U22210 ( .A(n19418), .B(n19419), .Z(n19416) );
  AND U22211 ( .A(a[33]), .B(b[42]), .Z(n19415) );
  XOR U22212 ( .A(n19420), .B(n19049), .Z(n19051) );
  XOR U22213 ( .A(n19421), .B(n19422), .Z(n19049) );
  AND U22214 ( .A(n19423), .B(n19424), .Z(n19421) );
  AND U22215 ( .A(a[34]), .B(b[41]), .Z(n19420) );
  XOR U22216 ( .A(n19425), .B(n19426), .Z(n19053) );
  AND U22217 ( .A(n19427), .B(n19428), .Z(n19425) );
  XOR U22218 ( .A(n19429), .B(n19058), .Z(n19060) );
  XOR U22219 ( .A(n19430), .B(n19431), .Z(n19058) );
  AND U22220 ( .A(n19432), .B(n19433), .Z(n19430) );
  AND U22221 ( .A(a[35]), .B(b[40]), .Z(n19429) );
  XOR U22222 ( .A(n19435), .B(n19436), .Z(n19063) );
  AND U22223 ( .A(n19437), .B(n19438), .Z(n19435) );
  AND U22224 ( .A(a[37]), .B(b[38]), .Z(n19434) );
  XOR U22225 ( .A(n19440), .B(n19441), .Z(n19068) );
  AND U22226 ( .A(n19442), .B(n19443), .Z(n19440) );
  AND U22227 ( .A(b[37]), .B(a[38]), .Z(n19439) );
  XOR U22228 ( .A(n19445), .B(n19446), .Z(n19073) );
  AND U22229 ( .A(n19447), .B(n19448), .Z(n19445) );
  AND U22230 ( .A(b[36]), .B(a[39]), .Z(n19444) );
  XOR U22231 ( .A(n19450), .B(n19451), .Z(n19078) );
  AND U22232 ( .A(n19452), .B(n19453), .Z(n19450) );
  AND U22233 ( .A(b[35]), .B(a[40]), .Z(n19449) );
  XOR U22234 ( .A(n19455), .B(n19456), .Z(n19083) );
  AND U22235 ( .A(n19457), .B(n19458), .Z(n19455) );
  AND U22236 ( .A(b[34]), .B(a[41]), .Z(n19454) );
  XOR U22237 ( .A(n19460), .B(n19461), .Z(n19088) );
  AND U22238 ( .A(n19462), .B(n19463), .Z(n19460) );
  AND U22239 ( .A(b[33]), .B(a[42]), .Z(n19459) );
  XOR U22240 ( .A(n19465), .B(n19466), .Z(n19093) );
  AND U22241 ( .A(n19467), .B(n19468), .Z(n19465) );
  AND U22242 ( .A(b[32]), .B(a[43]), .Z(n19464) );
  XOR U22243 ( .A(n19470), .B(n19471), .Z(n19098) );
  AND U22244 ( .A(n19472), .B(n19473), .Z(n19470) );
  AND U22245 ( .A(b[31]), .B(a[44]), .Z(n19469) );
  XOR U22246 ( .A(n19475), .B(n19476), .Z(n19103) );
  AND U22247 ( .A(n19477), .B(n19478), .Z(n19475) );
  AND U22248 ( .A(b[30]), .B(a[45]), .Z(n19474) );
  XOR U22249 ( .A(n19480), .B(n19481), .Z(n19108) );
  AND U22250 ( .A(n19482), .B(n19483), .Z(n19480) );
  AND U22251 ( .A(b[29]), .B(a[46]), .Z(n19479) );
  XOR U22252 ( .A(n19485), .B(n19486), .Z(n19113) );
  AND U22253 ( .A(n19487), .B(n19488), .Z(n19485) );
  AND U22254 ( .A(b[28]), .B(a[47]), .Z(n19484) );
  XOR U22255 ( .A(n19490), .B(n19491), .Z(n19118) );
  AND U22256 ( .A(n19492), .B(n19493), .Z(n19490) );
  AND U22257 ( .A(b[27]), .B(a[48]), .Z(n19489) );
  XOR U22258 ( .A(n19495), .B(n19496), .Z(n19123) );
  AND U22259 ( .A(n19497), .B(n19498), .Z(n19495) );
  AND U22260 ( .A(b[26]), .B(a[49]), .Z(n19494) );
  XOR U22261 ( .A(n19500), .B(n19501), .Z(n19128) );
  AND U22262 ( .A(n19502), .B(n19503), .Z(n19500) );
  AND U22263 ( .A(b[25]), .B(a[50]), .Z(n19499) );
  XOR U22264 ( .A(n19505), .B(n19506), .Z(n19133) );
  AND U22265 ( .A(n19507), .B(n19508), .Z(n19505) );
  AND U22266 ( .A(b[24]), .B(a[51]), .Z(n19504) );
  XOR U22267 ( .A(n19510), .B(n19511), .Z(n19138) );
  AND U22268 ( .A(n19512), .B(n19513), .Z(n19510) );
  AND U22269 ( .A(b[23]), .B(a[52]), .Z(n19509) );
  XOR U22270 ( .A(n19515), .B(n19516), .Z(n19143) );
  AND U22271 ( .A(n19517), .B(n19518), .Z(n19515) );
  AND U22272 ( .A(b[22]), .B(a[53]), .Z(n19514) );
  XOR U22273 ( .A(n19520), .B(n19521), .Z(n19148) );
  AND U22274 ( .A(n19522), .B(n19523), .Z(n19520) );
  AND U22275 ( .A(b[21]), .B(a[54]), .Z(n19519) );
  XOR U22276 ( .A(n19525), .B(n19526), .Z(n19153) );
  AND U22277 ( .A(n19527), .B(n19528), .Z(n19525) );
  AND U22278 ( .A(b[20]), .B(a[55]), .Z(n19524) );
  XOR U22279 ( .A(n19530), .B(n19531), .Z(n19158) );
  AND U22280 ( .A(n19532), .B(n19533), .Z(n19530) );
  AND U22281 ( .A(b[19]), .B(a[56]), .Z(n19529) );
  XOR U22282 ( .A(n19535), .B(n19536), .Z(n19163) );
  AND U22283 ( .A(n19537), .B(n19538), .Z(n19535) );
  AND U22284 ( .A(b[18]), .B(a[57]), .Z(n19534) );
  XOR U22285 ( .A(n19540), .B(n19541), .Z(n19168) );
  AND U22286 ( .A(n19542), .B(n19543), .Z(n19540) );
  AND U22287 ( .A(b[17]), .B(a[58]), .Z(n19539) );
  XOR U22288 ( .A(n19545), .B(n19546), .Z(n19173) );
  AND U22289 ( .A(n19547), .B(n19548), .Z(n19545) );
  AND U22290 ( .A(b[16]), .B(a[59]), .Z(n19544) );
  XOR U22291 ( .A(n19550), .B(n19551), .Z(n19178) );
  AND U22292 ( .A(n19552), .B(n19553), .Z(n19550) );
  AND U22293 ( .A(b[15]), .B(a[60]), .Z(n19549) );
  XOR U22294 ( .A(n19555), .B(n19556), .Z(n19183) );
  AND U22295 ( .A(n19557), .B(n19558), .Z(n19555) );
  AND U22296 ( .A(b[14]), .B(a[61]), .Z(n19554) );
  XOR U22297 ( .A(n19560), .B(n19561), .Z(n19188) );
  AND U22298 ( .A(n19562), .B(n19563), .Z(n19560) );
  AND U22299 ( .A(b[13]), .B(a[62]), .Z(n19559) );
  XOR U22300 ( .A(n19565), .B(n19566), .Z(n19193) );
  AND U22301 ( .A(n19567), .B(n19568), .Z(n19565) );
  AND U22302 ( .A(b[12]), .B(a[63]), .Z(n19564) );
  XOR U22303 ( .A(n19570), .B(n19571), .Z(n19198) );
  AND U22304 ( .A(n19572), .B(n19573), .Z(n19570) );
  AND U22305 ( .A(b[11]), .B(a[64]), .Z(n19569) );
  XOR U22306 ( .A(n19575), .B(n19576), .Z(n19203) );
  AND U22307 ( .A(n19577), .B(n19578), .Z(n19575) );
  AND U22308 ( .A(b[10]), .B(a[65]), .Z(n19574) );
  XOR U22309 ( .A(n19580), .B(n19581), .Z(n19208) );
  AND U22310 ( .A(n19582), .B(n19583), .Z(n19580) );
  AND U22311 ( .A(b[9]), .B(a[66]), .Z(n19579) );
  XOR U22312 ( .A(n19585), .B(n19586), .Z(n19213) );
  AND U22313 ( .A(n19587), .B(n19588), .Z(n19585) );
  AND U22314 ( .A(b[8]), .B(a[67]), .Z(n19584) );
  XOR U22315 ( .A(n19590), .B(n19591), .Z(n19218) );
  AND U22316 ( .A(n19592), .B(n19593), .Z(n19590) );
  AND U22317 ( .A(b[7]), .B(a[68]), .Z(n19589) );
  XOR U22318 ( .A(n19595), .B(n19596), .Z(n19223) );
  AND U22319 ( .A(n19597), .B(n19598), .Z(n19595) );
  AND U22320 ( .A(b[6]), .B(a[69]), .Z(n19594) );
  XOR U22321 ( .A(n19600), .B(n19601), .Z(n19228) );
  AND U22322 ( .A(n19602), .B(n19603), .Z(n19600) );
  AND U22323 ( .A(b[5]), .B(a[70]), .Z(n19599) );
  XOR U22324 ( .A(n19605), .B(n19606), .Z(n19233) );
  AND U22325 ( .A(n19607), .B(n19608), .Z(n19605) );
  AND U22326 ( .A(b[4]), .B(a[71]), .Z(n19604) );
  XOR U22327 ( .A(n19610), .B(n19611), .Z(n19238) );
  AND U22328 ( .A(n19612), .B(n19613), .Z(n19610) );
  AND U22329 ( .A(b[3]), .B(a[72]), .Z(n19609) );
  XOR U22330 ( .A(n19615), .B(n19616), .Z(n19243) );
  OR U22331 ( .A(n19617), .B(n19618), .Z(n19616) );
  AND U22332 ( .A(b[2]), .B(a[73]), .Z(n19614) );
  XNOR U22333 ( .A(n19253), .B(n19619), .Z(n19249) );
  NAND U22334 ( .A(b[1]), .B(a[74]), .Z(n19619) );
  IV U22335 ( .A(n19247), .Z(n19253) );
  ANDN U22336 ( .B(n10329), .A(n10331), .Z(n19247) );
  NAND U22337 ( .A(a[74]), .B(b[0]), .Z(n10331) );
  XOR U22338 ( .A(n19617), .B(n19618), .Z(n10329) );
  XOR U22339 ( .A(n19621), .B(n19612), .Z(n19620) );
  XOR U22340 ( .A(n19607), .B(n19611), .Z(n19622) );
  XOR U22341 ( .A(n19602), .B(n19606), .Z(n19623) );
  XOR U22342 ( .A(n19597), .B(n19601), .Z(n19624) );
  XOR U22343 ( .A(n19592), .B(n19596), .Z(n19625) );
  XOR U22344 ( .A(n19587), .B(n19591), .Z(n19626) );
  XOR U22345 ( .A(n19582), .B(n19586), .Z(n19627) );
  XOR U22346 ( .A(n19577), .B(n19581), .Z(n19628) );
  XOR U22347 ( .A(n19572), .B(n19576), .Z(n19629) );
  XOR U22348 ( .A(n19567), .B(n19571), .Z(n19630) );
  XOR U22349 ( .A(n19562), .B(n19566), .Z(n19631) );
  XOR U22350 ( .A(n19557), .B(n19561), .Z(n19632) );
  XOR U22351 ( .A(n19552), .B(n19556), .Z(n19633) );
  XOR U22352 ( .A(n19547), .B(n19551), .Z(n19634) );
  XOR U22353 ( .A(n19542), .B(n19546), .Z(n19635) );
  XOR U22354 ( .A(n19537), .B(n19541), .Z(n19636) );
  XOR U22355 ( .A(n19532), .B(n19536), .Z(n19637) );
  XOR U22356 ( .A(n19527), .B(n19531), .Z(n19638) );
  XOR U22357 ( .A(n19522), .B(n19526), .Z(n19639) );
  XOR U22358 ( .A(n19517), .B(n19521), .Z(n19640) );
  XOR U22359 ( .A(n19512), .B(n19516), .Z(n19641) );
  XOR U22360 ( .A(n19507), .B(n19511), .Z(n19642) );
  XOR U22361 ( .A(n19502), .B(n19506), .Z(n19643) );
  XOR U22362 ( .A(n19497), .B(n19501), .Z(n19644) );
  XOR U22363 ( .A(n19492), .B(n19496), .Z(n19645) );
  XOR U22364 ( .A(n19487), .B(n19491), .Z(n19646) );
  XOR U22365 ( .A(n19482), .B(n19486), .Z(n19647) );
  XOR U22366 ( .A(n19477), .B(n19481), .Z(n19648) );
  XOR U22367 ( .A(n19472), .B(n19476), .Z(n19649) );
  XOR U22368 ( .A(n19467), .B(n19471), .Z(n19650) );
  XOR U22369 ( .A(n19462), .B(n19466), .Z(n19651) );
  XOR U22370 ( .A(n19457), .B(n19461), .Z(n19652) );
  XOR U22371 ( .A(n19452), .B(n19456), .Z(n19653) );
  XOR U22372 ( .A(n19447), .B(n19451), .Z(n19654) );
  XOR U22373 ( .A(n19442), .B(n19446), .Z(n19655) );
  XOR U22374 ( .A(n19437), .B(n19441), .Z(n19656) );
  XOR U22375 ( .A(n19427), .B(n19436), .Z(n19657) );
  XOR U22376 ( .A(n19658), .B(n19426), .Z(n19427) );
  AND U22377 ( .A(a[36]), .B(b[38]), .Z(n19658) );
  XNOR U22378 ( .A(n19426), .B(n19432), .Z(n19659) );
  XNOR U22379 ( .A(n19431), .B(n19423), .Z(n19660) );
  XNOR U22380 ( .A(n19422), .B(n19418), .Z(n19661) );
  XNOR U22381 ( .A(n19417), .B(n19413), .Z(n19662) );
  XNOR U22382 ( .A(n19412), .B(n19408), .Z(n19663) );
  XNOR U22383 ( .A(n19407), .B(n19403), .Z(n19664) );
  XNOR U22384 ( .A(n19402), .B(n19398), .Z(n19665) );
  XNOR U22385 ( .A(n19397), .B(n19393), .Z(n19666) );
  XNOR U22386 ( .A(n19392), .B(n19388), .Z(n19667) );
  XNOR U22387 ( .A(n19387), .B(n19383), .Z(n19668) );
  XNOR U22388 ( .A(n19382), .B(n19378), .Z(n19669) );
  XNOR U22389 ( .A(n19377), .B(n19373), .Z(n19670) );
  XNOR U22390 ( .A(n19372), .B(n19368), .Z(n19671) );
  XNOR U22391 ( .A(n19367), .B(n19363), .Z(n19672) );
  XNOR U22392 ( .A(n19362), .B(n19358), .Z(n19673) );
  XNOR U22393 ( .A(n19357), .B(n19353), .Z(n19674) );
  XNOR U22394 ( .A(n19352), .B(n19348), .Z(n19675) );
  XNOR U22395 ( .A(n19347), .B(n19343), .Z(n19676) );
  XNOR U22396 ( .A(n19342), .B(n19338), .Z(n19677) );
  XNOR U22397 ( .A(n19337), .B(n19333), .Z(n19678) );
  XNOR U22398 ( .A(n19332), .B(n19328), .Z(n19679) );
  XOR U22399 ( .A(n19327), .B(n19324), .Z(n19680) );
  XOR U22400 ( .A(n19681), .B(n19682), .Z(n19324) );
  XOR U22401 ( .A(n19322), .B(n19683), .Z(n19682) );
  XOR U22402 ( .A(n19684), .B(n19685), .Z(n19683) );
  XOR U22403 ( .A(n19686), .B(n19687), .Z(n19685) );
  NAND U22404 ( .A(a[12]), .B(b[62]), .Z(n19687) );
  AND U22405 ( .A(a[11]), .B(b[63]), .Z(n19686) );
  XOR U22406 ( .A(n19688), .B(n19684), .Z(n19681) );
  XOR U22407 ( .A(n19689), .B(n19690), .Z(n19684) );
  ANDN U22408 ( .B(n19691), .A(n19692), .Z(n19689) );
  AND U22409 ( .A(a[13]), .B(b[61]), .Z(n19688) );
  XOR U22410 ( .A(n19693), .B(n19322), .Z(n19323) );
  XOR U22411 ( .A(n19694), .B(n19695), .Z(n19322) );
  AND U22412 ( .A(n19696), .B(n19697), .Z(n19694) );
  AND U22413 ( .A(a[14]), .B(b[60]), .Z(n19693) );
  XOR U22414 ( .A(n19698), .B(n19327), .Z(n19329) );
  XOR U22415 ( .A(n19699), .B(n19700), .Z(n19327) );
  AND U22416 ( .A(n19701), .B(n19702), .Z(n19699) );
  AND U22417 ( .A(a[15]), .B(b[59]), .Z(n19698) );
  XOR U22418 ( .A(n19703), .B(n19332), .Z(n19334) );
  XOR U22419 ( .A(n19704), .B(n19705), .Z(n19332) );
  AND U22420 ( .A(n19706), .B(n19707), .Z(n19704) );
  AND U22421 ( .A(a[16]), .B(b[58]), .Z(n19703) );
  XOR U22422 ( .A(n19708), .B(n19337), .Z(n19339) );
  XOR U22423 ( .A(n19709), .B(n19710), .Z(n19337) );
  AND U22424 ( .A(n19711), .B(n19712), .Z(n19709) );
  AND U22425 ( .A(a[17]), .B(b[57]), .Z(n19708) );
  XOR U22426 ( .A(n19713), .B(n19342), .Z(n19344) );
  XOR U22427 ( .A(n19714), .B(n19715), .Z(n19342) );
  AND U22428 ( .A(n19716), .B(n19717), .Z(n19714) );
  AND U22429 ( .A(a[18]), .B(b[56]), .Z(n19713) );
  XOR U22430 ( .A(n19718), .B(n19347), .Z(n19349) );
  XOR U22431 ( .A(n19719), .B(n19720), .Z(n19347) );
  AND U22432 ( .A(n19721), .B(n19722), .Z(n19719) );
  AND U22433 ( .A(a[19]), .B(b[55]), .Z(n19718) );
  XOR U22434 ( .A(n19723), .B(n19352), .Z(n19354) );
  XOR U22435 ( .A(n19724), .B(n19725), .Z(n19352) );
  AND U22436 ( .A(n19726), .B(n19727), .Z(n19724) );
  AND U22437 ( .A(a[20]), .B(b[54]), .Z(n19723) );
  XOR U22438 ( .A(n19728), .B(n19357), .Z(n19359) );
  XOR U22439 ( .A(n19729), .B(n19730), .Z(n19357) );
  AND U22440 ( .A(n19731), .B(n19732), .Z(n19729) );
  AND U22441 ( .A(a[21]), .B(b[53]), .Z(n19728) );
  XOR U22442 ( .A(n19733), .B(n19362), .Z(n19364) );
  XOR U22443 ( .A(n19734), .B(n19735), .Z(n19362) );
  AND U22444 ( .A(n19736), .B(n19737), .Z(n19734) );
  AND U22445 ( .A(a[22]), .B(b[52]), .Z(n19733) );
  XOR U22446 ( .A(n19738), .B(n19367), .Z(n19369) );
  XOR U22447 ( .A(n19739), .B(n19740), .Z(n19367) );
  AND U22448 ( .A(n19741), .B(n19742), .Z(n19739) );
  AND U22449 ( .A(a[23]), .B(b[51]), .Z(n19738) );
  XOR U22450 ( .A(n19743), .B(n19372), .Z(n19374) );
  XOR U22451 ( .A(n19744), .B(n19745), .Z(n19372) );
  AND U22452 ( .A(n19746), .B(n19747), .Z(n19744) );
  AND U22453 ( .A(a[24]), .B(b[50]), .Z(n19743) );
  XOR U22454 ( .A(n19748), .B(n19377), .Z(n19379) );
  XOR U22455 ( .A(n19749), .B(n19750), .Z(n19377) );
  AND U22456 ( .A(n19751), .B(n19752), .Z(n19749) );
  AND U22457 ( .A(a[25]), .B(b[49]), .Z(n19748) );
  XOR U22458 ( .A(n19753), .B(n19382), .Z(n19384) );
  XOR U22459 ( .A(n19754), .B(n19755), .Z(n19382) );
  AND U22460 ( .A(n19756), .B(n19757), .Z(n19754) );
  AND U22461 ( .A(a[26]), .B(b[48]), .Z(n19753) );
  XOR U22462 ( .A(n19758), .B(n19387), .Z(n19389) );
  XOR U22463 ( .A(n19759), .B(n19760), .Z(n19387) );
  AND U22464 ( .A(n19761), .B(n19762), .Z(n19759) );
  AND U22465 ( .A(a[27]), .B(b[47]), .Z(n19758) );
  XOR U22466 ( .A(n19763), .B(n19392), .Z(n19394) );
  XOR U22467 ( .A(n19764), .B(n19765), .Z(n19392) );
  AND U22468 ( .A(n19766), .B(n19767), .Z(n19764) );
  AND U22469 ( .A(a[28]), .B(b[46]), .Z(n19763) );
  XOR U22470 ( .A(n19768), .B(n19397), .Z(n19399) );
  XOR U22471 ( .A(n19769), .B(n19770), .Z(n19397) );
  AND U22472 ( .A(n19771), .B(n19772), .Z(n19769) );
  AND U22473 ( .A(a[29]), .B(b[45]), .Z(n19768) );
  XOR U22474 ( .A(n19773), .B(n19402), .Z(n19404) );
  XOR U22475 ( .A(n19774), .B(n19775), .Z(n19402) );
  AND U22476 ( .A(n19776), .B(n19777), .Z(n19774) );
  AND U22477 ( .A(a[30]), .B(b[44]), .Z(n19773) );
  XOR U22478 ( .A(n19778), .B(n19407), .Z(n19409) );
  XOR U22479 ( .A(n19779), .B(n19780), .Z(n19407) );
  AND U22480 ( .A(n19781), .B(n19782), .Z(n19779) );
  AND U22481 ( .A(a[31]), .B(b[43]), .Z(n19778) );
  XOR U22482 ( .A(n19783), .B(n19412), .Z(n19414) );
  XOR U22483 ( .A(n19784), .B(n19785), .Z(n19412) );
  AND U22484 ( .A(n19786), .B(n19787), .Z(n19784) );
  AND U22485 ( .A(a[32]), .B(b[42]), .Z(n19783) );
  XOR U22486 ( .A(n19788), .B(n19417), .Z(n19419) );
  XOR U22487 ( .A(n19789), .B(n19790), .Z(n19417) );
  AND U22488 ( .A(n19791), .B(n19792), .Z(n19789) );
  AND U22489 ( .A(a[33]), .B(b[41]), .Z(n19788) );
  XOR U22490 ( .A(n19793), .B(n19422), .Z(n19424) );
  XOR U22491 ( .A(n19794), .B(n19795), .Z(n19422) );
  AND U22492 ( .A(n19796), .B(n19797), .Z(n19794) );
  AND U22493 ( .A(a[34]), .B(b[40]), .Z(n19793) );
  XOR U22494 ( .A(n19798), .B(n19799), .Z(n19426) );
  AND U22495 ( .A(n19800), .B(n19801), .Z(n19798) );
  XOR U22496 ( .A(n19802), .B(n19431), .Z(n19433) );
  XOR U22497 ( .A(n19803), .B(n19804), .Z(n19431) );
  AND U22498 ( .A(n19805), .B(n19806), .Z(n19803) );
  AND U22499 ( .A(a[35]), .B(b[39]), .Z(n19802) );
  XOR U22500 ( .A(n19808), .B(n19809), .Z(n19436) );
  AND U22501 ( .A(n19810), .B(n19811), .Z(n19808) );
  AND U22502 ( .A(a[37]), .B(b[37]), .Z(n19807) );
  XOR U22503 ( .A(n19813), .B(n19814), .Z(n19441) );
  AND U22504 ( .A(n19815), .B(n19816), .Z(n19813) );
  AND U22505 ( .A(b[36]), .B(a[38]), .Z(n19812) );
  XOR U22506 ( .A(n19818), .B(n19819), .Z(n19446) );
  AND U22507 ( .A(n19820), .B(n19821), .Z(n19818) );
  AND U22508 ( .A(b[35]), .B(a[39]), .Z(n19817) );
  XOR U22509 ( .A(n19823), .B(n19824), .Z(n19451) );
  AND U22510 ( .A(n19825), .B(n19826), .Z(n19823) );
  AND U22511 ( .A(b[34]), .B(a[40]), .Z(n19822) );
  XOR U22512 ( .A(n19828), .B(n19829), .Z(n19456) );
  AND U22513 ( .A(n19830), .B(n19831), .Z(n19828) );
  AND U22514 ( .A(b[33]), .B(a[41]), .Z(n19827) );
  XOR U22515 ( .A(n19833), .B(n19834), .Z(n19461) );
  AND U22516 ( .A(n19835), .B(n19836), .Z(n19833) );
  AND U22517 ( .A(b[32]), .B(a[42]), .Z(n19832) );
  XOR U22518 ( .A(n19838), .B(n19839), .Z(n19466) );
  AND U22519 ( .A(n19840), .B(n19841), .Z(n19838) );
  AND U22520 ( .A(b[31]), .B(a[43]), .Z(n19837) );
  XOR U22521 ( .A(n19843), .B(n19844), .Z(n19471) );
  AND U22522 ( .A(n19845), .B(n19846), .Z(n19843) );
  AND U22523 ( .A(b[30]), .B(a[44]), .Z(n19842) );
  XOR U22524 ( .A(n19848), .B(n19849), .Z(n19476) );
  AND U22525 ( .A(n19850), .B(n19851), .Z(n19848) );
  AND U22526 ( .A(b[29]), .B(a[45]), .Z(n19847) );
  XOR U22527 ( .A(n19853), .B(n19854), .Z(n19481) );
  AND U22528 ( .A(n19855), .B(n19856), .Z(n19853) );
  AND U22529 ( .A(b[28]), .B(a[46]), .Z(n19852) );
  XOR U22530 ( .A(n19858), .B(n19859), .Z(n19486) );
  AND U22531 ( .A(n19860), .B(n19861), .Z(n19858) );
  AND U22532 ( .A(b[27]), .B(a[47]), .Z(n19857) );
  XOR U22533 ( .A(n19863), .B(n19864), .Z(n19491) );
  AND U22534 ( .A(n19865), .B(n19866), .Z(n19863) );
  AND U22535 ( .A(b[26]), .B(a[48]), .Z(n19862) );
  XOR U22536 ( .A(n19868), .B(n19869), .Z(n19496) );
  AND U22537 ( .A(n19870), .B(n19871), .Z(n19868) );
  AND U22538 ( .A(b[25]), .B(a[49]), .Z(n19867) );
  XOR U22539 ( .A(n19873), .B(n19874), .Z(n19501) );
  AND U22540 ( .A(n19875), .B(n19876), .Z(n19873) );
  AND U22541 ( .A(b[24]), .B(a[50]), .Z(n19872) );
  XOR U22542 ( .A(n19878), .B(n19879), .Z(n19506) );
  AND U22543 ( .A(n19880), .B(n19881), .Z(n19878) );
  AND U22544 ( .A(b[23]), .B(a[51]), .Z(n19877) );
  XOR U22545 ( .A(n19883), .B(n19884), .Z(n19511) );
  AND U22546 ( .A(n19885), .B(n19886), .Z(n19883) );
  AND U22547 ( .A(b[22]), .B(a[52]), .Z(n19882) );
  XOR U22548 ( .A(n19888), .B(n19889), .Z(n19516) );
  AND U22549 ( .A(n19890), .B(n19891), .Z(n19888) );
  AND U22550 ( .A(b[21]), .B(a[53]), .Z(n19887) );
  XOR U22551 ( .A(n19893), .B(n19894), .Z(n19521) );
  AND U22552 ( .A(n19895), .B(n19896), .Z(n19893) );
  AND U22553 ( .A(b[20]), .B(a[54]), .Z(n19892) );
  XOR U22554 ( .A(n19898), .B(n19899), .Z(n19526) );
  AND U22555 ( .A(n19900), .B(n19901), .Z(n19898) );
  AND U22556 ( .A(b[19]), .B(a[55]), .Z(n19897) );
  XOR U22557 ( .A(n19903), .B(n19904), .Z(n19531) );
  AND U22558 ( .A(n19905), .B(n19906), .Z(n19903) );
  AND U22559 ( .A(b[18]), .B(a[56]), .Z(n19902) );
  XOR U22560 ( .A(n19908), .B(n19909), .Z(n19536) );
  AND U22561 ( .A(n19910), .B(n19911), .Z(n19908) );
  AND U22562 ( .A(b[17]), .B(a[57]), .Z(n19907) );
  XOR U22563 ( .A(n19913), .B(n19914), .Z(n19541) );
  AND U22564 ( .A(n19915), .B(n19916), .Z(n19913) );
  AND U22565 ( .A(b[16]), .B(a[58]), .Z(n19912) );
  XOR U22566 ( .A(n19918), .B(n19919), .Z(n19546) );
  AND U22567 ( .A(n19920), .B(n19921), .Z(n19918) );
  AND U22568 ( .A(b[15]), .B(a[59]), .Z(n19917) );
  XOR U22569 ( .A(n19923), .B(n19924), .Z(n19551) );
  AND U22570 ( .A(n19925), .B(n19926), .Z(n19923) );
  AND U22571 ( .A(b[14]), .B(a[60]), .Z(n19922) );
  XOR U22572 ( .A(n19928), .B(n19929), .Z(n19556) );
  AND U22573 ( .A(n19930), .B(n19931), .Z(n19928) );
  AND U22574 ( .A(b[13]), .B(a[61]), .Z(n19927) );
  XOR U22575 ( .A(n19933), .B(n19934), .Z(n19561) );
  AND U22576 ( .A(n19935), .B(n19936), .Z(n19933) );
  AND U22577 ( .A(b[12]), .B(a[62]), .Z(n19932) );
  XOR U22578 ( .A(n19938), .B(n19939), .Z(n19566) );
  AND U22579 ( .A(n19940), .B(n19941), .Z(n19938) );
  AND U22580 ( .A(b[11]), .B(a[63]), .Z(n19937) );
  XOR U22581 ( .A(n19943), .B(n19944), .Z(n19571) );
  AND U22582 ( .A(n19945), .B(n19946), .Z(n19943) );
  AND U22583 ( .A(b[10]), .B(a[64]), .Z(n19942) );
  XOR U22584 ( .A(n19948), .B(n19949), .Z(n19576) );
  AND U22585 ( .A(n19950), .B(n19951), .Z(n19948) );
  AND U22586 ( .A(b[9]), .B(a[65]), .Z(n19947) );
  XOR U22587 ( .A(n19953), .B(n19954), .Z(n19581) );
  AND U22588 ( .A(n19955), .B(n19956), .Z(n19953) );
  AND U22589 ( .A(b[8]), .B(a[66]), .Z(n19952) );
  XOR U22590 ( .A(n19958), .B(n19959), .Z(n19586) );
  AND U22591 ( .A(n19960), .B(n19961), .Z(n19958) );
  AND U22592 ( .A(b[7]), .B(a[67]), .Z(n19957) );
  XOR U22593 ( .A(n19963), .B(n19964), .Z(n19591) );
  AND U22594 ( .A(n19965), .B(n19966), .Z(n19963) );
  AND U22595 ( .A(b[6]), .B(a[68]), .Z(n19962) );
  XOR U22596 ( .A(n19968), .B(n19969), .Z(n19596) );
  AND U22597 ( .A(n19970), .B(n19971), .Z(n19968) );
  AND U22598 ( .A(b[5]), .B(a[69]), .Z(n19967) );
  XOR U22599 ( .A(n19973), .B(n19974), .Z(n19601) );
  AND U22600 ( .A(n19975), .B(n19976), .Z(n19973) );
  AND U22601 ( .A(b[4]), .B(a[70]), .Z(n19972) );
  XOR U22602 ( .A(n19978), .B(n19979), .Z(n19606) );
  AND U22603 ( .A(n19980), .B(n19981), .Z(n19978) );
  AND U22604 ( .A(b[3]), .B(a[71]), .Z(n19977) );
  XOR U22605 ( .A(n19983), .B(n19984), .Z(n19611) );
  OR U22606 ( .A(n19985), .B(n19986), .Z(n19984) );
  AND U22607 ( .A(b[2]), .B(a[72]), .Z(n19982) );
  XNOR U22608 ( .A(n19621), .B(n19987), .Z(n19617) );
  NAND U22609 ( .A(b[1]), .B(a[73]), .Z(n19987) );
  IV U22610 ( .A(n19615), .Z(n19621) );
  ANDN U22611 ( .B(n10332), .A(n10334), .Z(n19615) );
  NAND U22612 ( .A(a[73]), .B(b[0]), .Z(n10334) );
  XOR U22613 ( .A(n19985), .B(n19986), .Z(n10332) );
  XOR U22614 ( .A(n19989), .B(n19980), .Z(n19988) );
  XOR U22615 ( .A(n19975), .B(n19979), .Z(n19990) );
  XOR U22616 ( .A(n19970), .B(n19974), .Z(n19991) );
  XOR U22617 ( .A(n19965), .B(n19969), .Z(n19992) );
  XOR U22618 ( .A(n19960), .B(n19964), .Z(n19993) );
  XOR U22619 ( .A(n19955), .B(n19959), .Z(n19994) );
  XOR U22620 ( .A(n19950), .B(n19954), .Z(n19995) );
  XOR U22621 ( .A(n19945), .B(n19949), .Z(n19996) );
  XOR U22622 ( .A(n19940), .B(n19944), .Z(n19997) );
  XOR U22623 ( .A(n19935), .B(n19939), .Z(n19998) );
  XOR U22624 ( .A(n19930), .B(n19934), .Z(n19999) );
  XOR U22625 ( .A(n19925), .B(n19929), .Z(n20000) );
  XOR U22626 ( .A(n19920), .B(n19924), .Z(n20001) );
  XOR U22627 ( .A(n19915), .B(n19919), .Z(n20002) );
  XOR U22628 ( .A(n19910), .B(n19914), .Z(n20003) );
  XOR U22629 ( .A(n19905), .B(n19909), .Z(n20004) );
  XOR U22630 ( .A(n19900), .B(n19904), .Z(n20005) );
  XOR U22631 ( .A(n19895), .B(n19899), .Z(n20006) );
  XOR U22632 ( .A(n19890), .B(n19894), .Z(n20007) );
  XOR U22633 ( .A(n19885), .B(n19889), .Z(n20008) );
  XOR U22634 ( .A(n19880), .B(n19884), .Z(n20009) );
  XOR U22635 ( .A(n19875), .B(n19879), .Z(n20010) );
  XOR U22636 ( .A(n19870), .B(n19874), .Z(n20011) );
  XOR U22637 ( .A(n19865), .B(n19869), .Z(n20012) );
  XOR U22638 ( .A(n19860), .B(n19864), .Z(n20013) );
  XOR U22639 ( .A(n19855), .B(n19859), .Z(n20014) );
  XOR U22640 ( .A(n19850), .B(n19854), .Z(n20015) );
  XOR U22641 ( .A(n19845), .B(n19849), .Z(n20016) );
  XOR U22642 ( .A(n19840), .B(n19844), .Z(n20017) );
  XOR U22643 ( .A(n19835), .B(n19839), .Z(n20018) );
  XOR U22644 ( .A(n19830), .B(n19834), .Z(n20019) );
  XOR U22645 ( .A(n19825), .B(n19829), .Z(n20020) );
  XOR U22646 ( .A(n19820), .B(n19824), .Z(n20021) );
  XOR U22647 ( .A(n19815), .B(n19819), .Z(n20022) );
  XOR U22648 ( .A(n19810), .B(n19814), .Z(n20023) );
  XOR U22649 ( .A(n19800), .B(n19809), .Z(n20024) );
  XOR U22650 ( .A(n20025), .B(n19799), .Z(n19800) );
  AND U22651 ( .A(a[36]), .B(b[37]), .Z(n20025) );
  XNOR U22652 ( .A(n19799), .B(n19805), .Z(n20026) );
  XNOR U22653 ( .A(n19804), .B(n19796), .Z(n20027) );
  XNOR U22654 ( .A(n19795), .B(n19791), .Z(n20028) );
  XNOR U22655 ( .A(n19790), .B(n19786), .Z(n20029) );
  XNOR U22656 ( .A(n19785), .B(n19781), .Z(n20030) );
  XNOR U22657 ( .A(n19780), .B(n19776), .Z(n20031) );
  XNOR U22658 ( .A(n19775), .B(n19771), .Z(n20032) );
  XNOR U22659 ( .A(n19770), .B(n19766), .Z(n20033) );
  XNOR U22660 ( .A(n19765), .B(n19761), .Z(n20034) );
  XNOR U22661 ( .A(n19760), .B(n19756), .Z(n20035) );
  XNOR U22662 ( .A(n19755), .B(n19751), .Z(n20036) );
  XNOR U22663 ( .A(n19750), .B(n19746), .Z(n20037) );
  XNOR U22664 ( .A(n19745), .B(n19741), .Z(n20038) );
  XNOR U22665 ( .A(n19740), .B(n19736), .Z(n20039) );
  XNOR U22666 ( .A(n19735), .B(n19731), .Z(n20040) );
  XNOR U22667 ( .A(n19730), .B(n19726), .Z(n20041) );
  XNOR U22668 ( .A(n19725), .B(n19721), .Z(n20042) );
  XNOR U22669 ( .A(n19720), .B(n19716), .Z(n20043) );
  XNOR U22670 ( .A(n19715), .B(n19711), .Z(n20044) );
  XNOR U22671 ( .A(n19710), .B(n19706), .Z(n20045) );
  XNOR U22672 ( .A(n19705), .B(n19701), .Z(n20046) );
  XNOR U22673 ( .A(n19700), .B(n19696), .Z(n20047) );
  XOR U22674 ( .A(n19695), .B(n19692), .Z(n20048) );
  XOR U22675 ( .A(n20049), .B(n20050), .Z(n19692) );
  XOR U22676 ( .A(n19690), .B(n20051), .Z(n20050) );
  XOR U22677 ( .A(n20052), .B(n20053), .Z(n20051) );
  XOR U22678 ( .A(n20054), .B(n20055), .Z(n20053) );
  NAND U22679 ( .A(a[11]), .B(b[62]), .Z(n20055) );
  AND U22680 ( .A(a[10]), .B(b[63]), .Z(n20054) );
  XOR U22681 ( .A(n20056), .B(n20052), .Z(n20049) );
  XOR U22682 ( .A(n20057), .B(n20058), .Z(n20052) );
  ANDN U22683 ( .B(n20059), .A(n20060), .Z(n20057) );
  AND U22684 ( .A(a[12]), .B(b[61]), .Z(n20056) );
  XOR U22685 ( .A(n20061), .B(n19690), .Z(n19691) );
  XOR U22686 ( .A(n20062), .B(n20063), .Z(n19690) );
  AND U22687 ( .A(n20064), .B(n20065), .Z(n20062) );
  AND U22688 ( .A(a[13]), .B(b[60]), .Z(n20061) );
  XOR U22689 ( .A(n20066), .B(n19695), .Z(n19697) );
  XOR U22690 ( .A(n20067), .B(n20068), .Z(n19695) );
  AND U22691 ( .A(n20069), .B(n20070), .Z(n20067) );
  AND U22692 ( .A(a[14]), .B(b[59]), .Z(n20066) );
  XOR U22693 ( .A(n20071), .B(n19700), .Z(n19702) );
  XOR U22694 ( .A(n20072), .B(n20073), .Z(n19700) );
  AND U22695 ( .A(n20074), .B(n20075), .Z(n20072) );
  AND U22696 ( .A(a[15]), .B(b[58]), .Z(n20071) );
  XOR U22697 ( .A(n20076), .B(n19705), .Z(n19707) );
  XOR U22698 ( .A(n20077), .B(n20078), .Z(n19705) );
  AND U22699 ( .A(n20079), .B(n20080), .Z(n20077) );
  AND U22700 ( .A(a[16]), .B(b[57]), .Z(n20076) );
  XOR U22701 ( .A(n20081), .B(n19710), .Z(n19712) );
  XOR U22702 ( .A(n20082), .B(n20083), .Z(n19710) );
  AND U22703 ( .A(n20084), .B(n20085), .Z(n20082) );
  AND U22704 ( .A(a[17]), .B(b[56]), .Z(n20081) );
  XOR U22705 ( .A(n20086), .B(n19715), .Z(n19717) );
  XOR U22706 ( .A(n20087), .B(n20088), .Z(n19715) );
  AND U22707 ( .A(n20089), .B(n20090), .Z(n20087) );
  AND U22708 ( .A(a[18]), .B(b[55]), .Z(n20086) );
  XOR U22709 ( .A(n20091), .B(n19720), .Z(n19722) );
  XOR U22710 ( .A(n20092), .B(n20093), .Z(n19720) );
  AND U22711 ( .A(n20094), .B(n20095), .Z(n20092) );
  AND U22712 ( .A(a[19]), .B(b[54]), .Z(n20091) );
  XOR U22713 ( .A(n20096), .B(n19725), .Z(n19727) );
  XOR U22714 ( .A(n20097), .B(n20098), .Z(n19725) );
  AND U22715 ( .A(n20099), .B(n20100), .Z(n20097) );
  AND U22716 ( .A(a[20]), .B(b[53]), .Z(n20096) );
  XOR U22717 ( .A(n20101), .B(n19730), .Z(n19732) );
  XOR U22718 ( .A(n20102), .B(n20103), .Z(n19730) );
  AND U22719 ( .A(n20104), .B(n20105), .Z(n20102) );
  AND U22720 ( .A(a[21]), .B(b[52]), .Z(n20101) );
  XOR U22721 ( .A(n20106), .B(n19735), .Z(n19737) );
  XOR U22722 ( .A(n20107), .B(n20108), .Z(n19735) );
  AND U22723 ( .A(n20109), .B(n20110), .Z(n20107) );
  AND U22724 ( .A(a[22]), .B(b[51]), .Z(n20106) );
  XOR U22725 ( .A(n20111), .B(n19740), .Z(n19742) );
  XOR U22726 ( .A(n20112), .B(n20113), .Z(n19740) );
  AND U22727 ( .A(n20114), .B(n20115), .Z(n20112) );
  AND U22728 ( .A(a[23]), .B(b[50]), .Z(n20111) );
  XOR U22729 ( .A(n20116), .B(n19745), .Z(n19747) );
  XOR U22730 ( .A(n20117), .B(n20118), .Z(n19745) );
  AND U22731 ( .A(n20119), .B(n20120), .Z(n20117) );
  AND U22732 ( .A(a[24]), .B(b[49]), .Z(n20116) );
  XOR U22733 ( .A(n20121), .B(n19750), .Z(n19752) );
  XOR U22734 ( .A(n20122), .B(n20123), .Z(n19750) );
  AND U22735 ( .A(n20124), .B(n20125), .Z(n20122) );
  AND U22736 ( .A(a[25]), .B(b[48]), .Z(n20121) );
  XOR U22737 ( .A(n20126), .B(n19755), .Z(n19757) );
  XOR U22738 ( .A(n20127), .B(n20128), .Z(n19755) );
  AND U22739 ( .A(n20129), .B(n20130), .Z(n20127) );
  AND U22740 ( .A(a[26]), .B(b[47]), .Z(n20126) );
  XOR U22741 ( .A(n20131), .B(n19760), .Z(n19762) );
  XOR U22742 ( .A(n20132), .B(n20133), .Z(n19760) );
  AND U22743 ( .A(n20134), .B(n20135), .Z(n20132) );
  AND U22744 ( .A(a[27]), .B(b[46]), .Z(n20131) );
  XOR U22745 ( .A(n20136), .B(n19765), .Z(n19767) );
  XOR U22746 ( .A(n20137), .B(n20138), .Z(n19765) );
  AND U22747 ( .A(n20139), .B(n20140), .Z(n20137) );
  AND U22748 ( .A(a[28]), .B(b[45]), .Z(n20136) );
  XOR U22749 ( .A(n20141), .B(n19770), .Z(n19772) );
  XOR U22750 ( .A(n20142), .B(n20143), .Z(n19770) );
  AND U22751 ( .A(n20144), .B(n20145), .Z(n20142) );
  AND U22752 ( .A(a[29]), .B(b[44]), .Z(n20141) );
  XOR U22753 ( .A(n20146), .B(n19775), .Z(n19777) );
  XOR U22754 ( .A(n20147), .B(n20148), .Z(n19775) );
  AND U22755 ( .A(n20149), .B(n20150), .Z(n20147) );
  AND U22756 ( .A(a[30]), .B(b[43]), .Z(n20146) );
  XOR U22757 ( .A(n20151), .B(n19780), .Z(n19782) );
  XOR U22758 ( .A(n20152), .B(n20153), .Z(n19780) );
  AND U22759 ( .A(n20154), .B(n20155), .Z(n20152) );
  AND U22760 ( .A(a[31]), .B(b[42]), .Z(n20151) );
  XOR U22761 ( .A(n20156), .B(n19785), .Z(n19787) );
  XOR U22762 ( .A(n20157), .B(n20158), .Z(n19785) );
  AND U22763 ( .A(n20159), .B(n20160), .Z(n20157) );
  AND U22764 ( .A(a[32]), .B(b[41]), .Z(n20156) );
  XOR U22765 ( .A(n20161), .B(n19790), .Z(n19792) );
  XOR U22766 ( .A(n20162), .B(n20163), .Z(n19790) );
  AND U22767 ( .A(n20164), .B(n20165), .Z(n20162) );
  AND U22768 ( .A(a[33]), .B(b[40]), .Z(n20161) );
  XOR U22769 ( .A(n20166), .B(n19795), .Z(n19797) );
  XOR U22770 ( .A(n20167), .B(n20168), .Z(n19795) );
  AND U22771 ( .A(n20169), .B(n20170), .Z(n20167) );
  AND U22772 ( .A(a[34]), .B(b[39]), .Z(n20166) );
  XOR U22773 ( .A(n20171), .B(n20172), .Z(n19799) );
  AND U22774 ( .A(n20173), .B(n20174), .Z(n20171) );
  XOR U22775 ( .A(n20175), .B(n19804), .Z(n19806) );
  XOR U22776 ( .A(n20176), .B(n20177), .Z(n19804) );
  AND U22777 ( .A(n20178), .B(n20179), .Z(n20176) );
  AND U22778 ( .A(a[35]), .B(b[38]), .Z(n20175) );
  XOR U22779 ( .A(n20181), .B(n20182), .Z(n19809) );
  AND U22780 ( .A(n20183), .B(n20184), .Z(n20181) );
  AND U22781 ( .A(b[36]), .B(a[37]), .Z(n20180) );
  XOR U22782 ( .A(n20186), .B(n20187), .Z(n19814) );
  AND U22783 ( .A(n20188), .B(n20189), .Z(n20186) );
  AND U22784 ( .A(b[35]), .B(a[38]), .Z(n20185) );
  XOR U22785 ( .A(n20191), .B(n20192), .Z(n19819) );
  AND U22786 ( .A(n20193), .B(n20194), .Z(n20191) );
  AND U22787 ( .A(b[34]), .B(a[39]), .Z(n20190) );
  XOR U22788 ( .A(n20196), .B(n20197), .Z(n19824) );
  AND U22789 ( .A(n20198), .B(n20199), .Z(n20196) );
  AND U22790 ( .A(b[33]), .B(a[40]), .Z(n20195) );
  XOR U22791 ( .A(n20201), .B(n20202), .Z(n19829) );
  AND U22792 ( .A(n20203), .B(n20204), .Z(n20201) );
  AND U22793 ( .A(b[32]), .B(a[41]), .Z(n20200) );
  XOR U22794 ( .A(n20206), .B(n20207), .Z(n19834) );
  AND U22795 ( .A(n20208), .B(n20209), .Z(n20206) );
  AND U22796 ( .A(b[31]), .B(a[42]), .Z(n20205) );
  XOR U22797 ( .A(n20211), .B(n20212), .Z(n19839) );
  AND U22798 ( .A(n20213), .B(n20214), .Z(n20211) );
  AND U22799 ( .A(b[30]), .B(a[43]), .Z(n20210) );
  XOR U22800 ( .A(n20216), .B(n20217), .Z(n19844) );
  AND U22801 ( .A(n20218), .B(n20219), .Z(n20216) );
  AND U22802 ( .A(b[29]), .B(a[44]), .Z(n20215) );
  XOR U22803 ( .A(n20221), .B(n20222), .Z(n19849) );
  AND U22804 ( .A(n20223), .B(n20224), .Z(n20221) );
  AND U22805 ( .A(b[28]), .B(a[45]), .Z(n20220) );
  XOR U22806 ( .A(n20226), .B(n20227), .Z(n19854) );
  AND U22807 ( .A(n20228), .B(n20229), .Z(n20226) );
  AND U22808 ( .A(b[27]), .B(a[46]), .Z(n20225) );
  XOR U22809 ( .A(n20231), .B(n20232), .Z(n19859) );
  AND U22810 ( .A(n20233), .B(n20234), .Z(n20231) );
  AND U22811 ( .A(b[26]), .B(a[47]), .Z(n20230) );
  XOR U22812 ( .A(n20236), .B(n20237), .Z(n19864) );
  AND U22813 ( .A(n20238), .B(n20239), .Z(n20236) );
  AND U22814 ( .A(b[25]), .B(a[48]), .Z(n20235) );
  XOR U22815 ( .A(n20241), .B(n20242), .Z(n19869) );
  AND U22816 ( .A(n20243), .B(n20244), .Z(n20241) );
  AND U22817 ( .A(b[24]), .B(a[49]), .Z(n20240) );
  XOR U22818 ( .A(n20246), .B(n20247), .Z(n19874) );
  AND U22819 ( .A(n20248), .B(n20249), .Z(n20246) );
  AND U22820 ( .A(b[23]), .B(a[50]), .Z(n20245) );
  XOR U22821 ( .A(n20251), .B(n20252), .Z(n19879) );
  AND U22822 ( .A(n20253), .B(n20254), .Z(n20251) );
  AND U22823 ( .A(b[22]), .B(a[51]), .Z(n20250) );
  XOR U22824 ( .A(n20256), .B(n20257), .Z(n19884) );
  AND U22825 ( .A(n20258), .B(n20259), .Z(n20256) );
  AND U22826 ( .A(b[21]), .B(a[52]), .Z(n20255) );
  XOR U22827 ( .A(n20261), .B(n20262), .Z(n19889) );
  AND U22828 ( .A(n20263), .B(n20264), .Z(n20261) );
  AND U22829 ( .A(b[20]), .B(a[53]), .Z(n20260) );
  XOR U22830 ( .A(n20266), .B(n20267), .Z(n19894) );
  AND U22831 ( .A(n20268), .B(n20269), .Z(n20266) );
  AND U22832 ( .A(b[19]), .B(a[54]), .Z(n20265) );
  XOR U22833 ( .A(n20271), .B(n20272), .Z(n19899) );
  AND U22834 ( .A(n20273), .B(n20274), .Z(n20271) );
  AND U22835 ( .A(b[18]), .B(a[55]), .Z(n20270) );
  XOR U22836 ( .A(n20276), .B(n20277), .Z(n19904) );
  AND U22837 ( .A(n20278), .B(n20279), .Z(n20276) );
  AND U22838 ( .A(b[17]), .B(a[56]), .Z(n20275) );
  XOR U22839 ( .A(n20281), .B(n20282), .Z(n19909) );
  AND U22840 ( .A(n20283), .B(n20284), .Z(n20281) );
  AND U22841 ( .A(b[16]), .B(a[57]), .Z(n20280) );
  XOR U22842 ( .A(n20286), .B(n20287), .Z(n19914) );
  AND U22843 ( .A(n20288), .B(n20289), .Z(n20286) );
  AND U22844 ( .A(b[15]), .B(a[58]), .Z(n20285) );
  XOR U22845 ( .A(n20291), .B(n20292), .Z(n19919) );
  AND U22846 ( .A(n20293), .B(n20294), .Z(n20291) );
  AND U22847 ( .A(b[14]), .B(a[59]), .Z(n20290) );
  XOR U22848 ( .A(n20296), .B(n20297), .Z(n19924) );
  AND U22849 ( .A(n20298), .B(n20299), .Z(n20296) );
  AND U22850 ( .A(b[13]), .B(a[60]), .Z(n20295) );
  XOR U22851 ( .A(n20301), .B(n20302), .Z(n19929) );
  AND U22852 ( .A(n20303), .B(n20304), .Z(n20301) );
  AND U22853 ( .A(b[12]), .B(a[61]), .Z(n20300) );
  XOR U22854 ( .A(n20306), .B(n20307), .Z(n19934) );
  AND U22855 ( .A(n20308), .B(n20309), .Z(n20306) );
  AND U22856 ( .A(b[11]), .B(a[62]), .Z(n20305) );
  XOR U22857 ( .A(n20311), .B(n20312), .Z(n19939) );
  AND U22858 ( .A(n20313), .B(n20314), .Z(n20311) );
  AND U22859 ( .A(b[10]), .B(a[63]), .Z(n20310) );
  XOR U22860 ( .A(n20316), .B(n20317), .Z(n19944) );
  AND U22861 ( .A(n20318), .B(n20319), .Z(n20316) );
  AND U22862 ( .A(b[9]), .B(a[64]), .Z(n20315) );
  XOR U22863 ( .A(n20321), .B(n20322), .Z(n19949) );
  AND U22864 ( .A(n20323), .B(n20324), .Z(n20321) );
  AND U22865 ( .A(b[8]), .B(a[65]), .Z(n20320) );
  XOR U22866 ( .A(n20326), .B(n20327), .Z(n19954) );
  AND U22867 ( .A(n20328), .B(n20329), .Z(n20326) );
  AND U22868 ( .A(b[7]), .B(a[66]), .Z(n20325) );
  XOR U22869 ( .A(n20331), .B(n20332), .Z(n19959) );
  AND U22870 ( .A(n20333), .B(n20334), .Z(n20331) );
  AND U22871 ( .A(b[6]), .B(a[67]), .Z(n20330) );
  XOR U22872 ( .A(n20336), .B(n20337), .Z(n19964) );
  AND U22873 ( .A(n20338), .B(n20339), .Z(n20336) );
  AND U22874 ( .A(b[5]), .B(a[68]), .Z(n20335) );
  XOR U22875 ( .A(n20341), .B(n20342), .Z(n19969) );
  AND U22876 ( .A(n20343), .B(n20344), .Z(n20341) );
  AND U22877 ( .A(b[4]), .B(a[69]), .Z(n20340) );
  XOR U22878 ( .A(n20346), .B(n20347), .Z(n19974) );
  AND U22879 ( .A(n20348), .B(n20349), .Z(n20346) );
  AND U22880 ( .A(b[3]), .B(a[70]), .Z(n20345) );
  XOR U22881 ( .A(n20351), .B(n20352), .Z(n19979) );
  OR U22882 ( .A(n20353), .B(n20354), .Z(n20352) );
  AND U22883 ( .A(b[2]), .B(a[71]), .Z(n20350) );
  XNOR U22884 ( .A(n19989), .B(n20355), .Z(n19985) );
  NAND U22885 ( .A(b[1]), .B(a[72]), .Z(n20355) );
  IV U22886 ( .A(n19983), .Z(n19989) );
  ANDN U22887 ( .B(n10335), .A(n10337), .Z(n19983) );
  NAND U22888 ( .A(a[72]), .B(b[0]), .Z(n10337) );
  XOR U22889 ( .A(n20353), .B(n20354), .Z(n10335) );
  XOR U22890 ( .A(n20357), .B(n20348), .Z(n20356) );
  XOR U22891 ( .A(n20343), .B(n20347), .Z(n20358) );
  XOR U22892 ( .A(n20338), .B(n20342), .Z(n20359) );
  XOR U22893 ( .A(n20333), .B(n20337), .Z(n20360) );
  XOR U22894 ( .A(n20328), .B(n20332), .Z(n20361) );
  XOR U22895 ( .A(n20323), .B(n20327), .Z(n20362) );
  XOR U22896 ( .A(n20318), .B(n20322), .Z(n20363) );
  XOR U22897 ( .A(n20313), .B(n20317), .Z(n20364) );
  XOR U22898 ( .A(n20308), .B(n20312), .Z(n20365) );
  XOR U22899 ( .A(n20303), .B(n20307), .Z(n20366) );
  XOR U22900 ( .A(n20298), .B(n20302), .Z(n20367) );
  XOR U22901 ( .A(n20293), .B(n20297), .Z(n20368) );
  XOR U22902 ( .A(n20288), .B(n20292), .Z(n20369) );
  XOR U22903 ( .A(n20283), .B(n20287), .Z(n20370) );
  XOR U22904 ( .A(n20278), .B(n20282), .Z(n20371) );
  XOR U22905 ( .A(n20273), .B(n20277), .Z(n20372) );
  XOR U22906 ( .A(n20268), .B(n20272), .Z(n20373) );
  XOR U22907 ( .A(n20263), .B(n20267), .Z(n20374) );
  XOR U22908 ( .A(n20258), .B(n20262), .Z(n20375) );
  XOR U22909 ( .A(n20253), .B(n20257), .Z(n20376) );
  XOR U22910 ( .A(n20248), .B(n20252), .Z(n20377) );
  XOR U22911 ( .A(n20243), .B(n20247), .Z(n20378) );
  XOR U22912 ( .A(n20238), .B(n20242), .Z(n20379) );
  XOR U22913 ( .A(n20233), .B(n20237), .Z(n20380) );
  XOR U22914 ( .A(n20228), .B(n20232), .Z(n20381) );
  XOR U22915 ( .A(n20223), .B(n20227), .Z(n20382) );
  XOR U22916 ( .A(n20218), .B(n20222), .Z(n20383) );
  XOR U22917 ( .A(n20213), .B(n20217), .Z(n20384) );
  XOR U22918 ( .A(n20208), .B(n20212), .Z(n20385) );
  XOR U22919 ( .A(n20203), .B(n20207), .Z(n20386) );
  XOR U22920 ( .A(n20198), .B(n20202), .Z(n20387) );
  XOR U22921 ( .A(n20193), .B(n20197), .Z(n20388) );
  XOR U22922 ( .A(n20188), .B(n20192), .Z(n20389) );
  XOR U22923 ( .A(n20183), .B(n20187), .Z(n20390) );
  XOR U22924 ( .A(n20173), .B(n20182), .Z(n20391) );
  XOR U22925 ( .A(n20392), .B(n20172), .Z(n20173) );
  AND U22926 ( .A(a[36]), .B(b[36]), .Z(n20392) );
  XNOR U22927 ( .A(n20172), .B(n20178), .Z(n20393) );
  XNOR U22928 ( .A(n20177), .B(n20169), .Z(n20394) );
  XNOR U22929 ( .A(n20168), .B(n20164), .Z(n20395) );
  XNOR U22930 ( .A(n20163), .B(n20159), .Z(n20396) );
  XNOR U22931 ( .A(n20158), .B(n20154), .Z(n20397) );
  XNOR U22932 ( .A(n20153), .B(n20149), .Z(n20398) );
  XNOR U22933 ( .A(n20148), .B(n20144), .Z(n20399) );
  XNOR U22934 ( .A(n20143), .B(n20139), .Z(n20400) );
  XNOR U22935 ( .A(n20138), .B(n20134), .Z(n20401) );
  XNOR U22936 ( .A(n20133), .B(n20129), .Z(n20402) );
  XNOR U22937 ( .A(n20128), .B(n20124), .Z(n20403) );
  XNOR U22938 ( .A(n20123), .B(n20119), .Z(n20404) );
  XNOR U22939 ( .A(n20118), .B(n20114), .Z(n20405) );
  XNOR U22940 ( .A(n20113), .B(n20109), .Z(n20406) );
  XNOR U22941 ( .A(n20108), .B(n20104), .Z(n20407) );
  XNOR U22942 ( .A(n20103), .B(n20099), .Z(n20408) );
  XNOR U22943 ( .A(n20098), .B(n20094), .Z(n20409) );
  XNOR U22944 ( .A(n20093), .B(n20089), .Z(n20410) );
  XNOR U22945 ( .A(n20088), .B(n20084), .Z(n20411) );
  XNOR U22946 ( .A(n20083), .B(n20079), .Z(n20412) );
  XNOR U22947 ( .A(n20078), .B(n20074), .Z(n20413) );
  XNOR U22948 ( .A(n20073), .B(n20069), .Z(n20414) );
  XNOR U22949 ( .A(n20068), .B(n20064), .Z(n20415) );
  XOR U22950 ( .A(n20063), .B(n20060), .Z(n20416) );
  XOR U22951 ( .A(n20417), .B(n20418), .Z(n20060) );
  XOR U22952 ( .A(n20058), .B(n20419), .Z(n20418) );
  XOR U22953 ( .A(n20420), .B(n20421), .Z(n20419) );
  XOR U22954 ( .A(n20422), .B(n20423), .Z(n20421) );
  NAND U22955 ( .A(a[10]), .B(b[62]), .Z(n20423) );
  AND U22956 ( .A(a[9]), .B(b[63]), .Z(n20422) );
  XOR U22957 ( .A(n20424), .B(n20420), .Z(n20417) );
  XOR U22958 ( .A(n20425), .B(n20426), .Z(n20420) );
  ANDN U22959 ( .B(n20427), .A(n20428), .Z(n20425) );
  AND U22960 ( .A(a[11]), .B(b[61]), .Z(n20424) );
  XOR U22961 ( .A(n20429), .B(n20058), .Z(n20059) );
  XOR U22962 ( .A(n20430), .B(n20431), .Z(n20058) );
  AND U22963 ( .A(n20432), .B(n20433), .Z(n20430) );
  AND U22964 ( .A(a[12]), .B(b[60]), .Z(n20429) );
  XOR U22965 ( .A(n20434), .B(n20063), .Z(n20065) );
  XOR U22966 ( .A(n20435), .B(n20436), .Z(n20063) );
  AND U22967 ( .A(n20437), .B(n20438), .Z(n20435) );
  AND U22968 ( .A(a[13]), .B(b[59]), .Z(n20434) );
  XOR U22969 ( .A(n20439), .B(n20068), .Z(n20070) );
  XOR U22970 ( .A(n20440), .B(n20441), .Z(n20068) );
  AND U22971 ( .A(n20442), .B(n20443), .Z(n20440) );
  AND U22972 ( .A(a[14]), .B(b[58]), .Z(n20439) );
  XOR U22973 ( .A(n20444), .B(n20073), .Z(n20075) );
  XOR U22974 ( .A(n20445), .B(n20446), .Z(n20073) );
  AND U22975 ( .A(n20447), .B(n20448), .Z(n20445) );
  AND U22976 ( .A(a[15]), .B(b[57]), .Z(n20444) );
  XOR U22977 ( .A(n20449), .B(n20078), .Z(n20080) );
  XOR U22978 ( .A(n20450), .B(n20451), .Z(n20078) );
  AND U22979 ( .A(n20452), .B(n20453), .Z(n20450) );
  AND U22980 ( .A(a[16]), .B(b[56]), .Z(n20449) );
  XOR U22981 ( .A(n20454), .B(n20083), .Z(n20085) );
  XOR U22982 ( .A(n20455), .B(n20456), .Z(n20083) );
  AND U22983 ( .A(n20457), .B(n20458), .Z(n20455) );
  AND U22984 ( .A(a[17]), .B(b[55]), .Z(n20454) );
  XOR U22985 ( .A(n20459), .B(n20088), .Z(n20090) );
  XOR U22986 ( .A(n20460), .B(n20461), .Z(n20088) );
  AND U22987 ( .A(n20462), .B(n20463), .Z(n20460) );
  AND U22988 ( .A(a[18]), .B(b[54]), .Z(n20459) );
  XOR U22989 ( .A(n20464), .B(n20093), .Z(n20095) );
  XOR U22990 ( .A(n20465), .B(n20466), .Z(n20093) );
  AND U22991 ( .A(n20467), .B(n20468), .Z(n20465) );
  AND U22992 ( .A(a[19]), .B(b[53]), .Z(n20464) );
  XOR U22993 ( .A(n20469), .B(n20098), .Z(n20100) );
  XOR U22994 ( .A(n20470), .B(n20471), .Z(n20098) );
  AND U22995 ( .A(n20472), .B(n20473), .Z(n20470) );
  AND U22996 ( .A(a[20]), .B(b[52]), .Z(n20469) );
  XOR U22997 ( .A(n20474), .B(n20103), .Z(n20105) );
  XOR U22998 ( .A(n20475), .B(n20476), .Z(n20103) );
  AND U22999 ( .A(n20477), .B(n20478), .Z(n20475) );
  AND U23000 ( .A(a[21]), .B(b[51]), .Z(n20474) );
  XOR U23001 ( .A(n20479), .B(n20108), .Z(n20110) );
  XOR U23002 ( .A(n20480), .B(n20481), .Z(n20108) );
  AND U23003 ( .A(n20482), .B(n20483), .Z(n20480) );
  AND U23004 ( .A(a[22]), .B(b[50]), .Z(n20479) );
  XOR U23005 ( .A(n20484), .B(n20113), .Z(n20115) );
  XOR U23006 ( .A(n20485), .B(n20486), .Z(n20113) );
  AND U23007 ( .A(n20487), .B(n20488), .Z(n20485) );
  AND U23008 ( .A(a[23]), .B(b[49]), .Z(n20484) );
  XOR U23009 ( .A(n20489), .B(n20118), .Z(n20120) );
  XOR U23010 ( .A(n20490), .B(n20491), .Z(n20118) );
  AND U23011 ( .A(n20492), .B(n20493), .Z(n20490) );
  AND U23012 ( .A(a[24]), .B(b[48]), .Z(n20489) );
  XOR U23013 ( .A(n20494), .B(n20123), .Z(n20125) );
  XOR U23014 ( .A(n20495), .B(n20496), .Z(n20123) );
  AND U23015 ( .A(n20497), .B(n20498), .Z(n20495) );
  AND U23016 ( .A(a[25]), .B(b[47]), .Z(n20494) );
  XOR U23017 ( .A(n20499), .B(n20128), .Z(n20130) );
  XOR U23018 ( .A(n20500), .B(n20501), .Z(n20128) );
  AND U23019 ( .A(n20502), .B(n20503), .Z(n20500) );
  AND U23020 ( .A(a[26]), .B(b[46]), .Z(n20499) );
  XOR U23021 ( .A(n20504), .B(n20133), .Z(n20135) );
  XOR U23022 ( .A(n20505), .B(n20506), .Z(n20133) );
  AND U23023 ( .A(n20507), .B(n20508), .Z(n20505) );
  AND U23024 ( .A(a[27]), .B(b[45]), .Z(n20504) );
  XOR U23025 ( .A(n20509), .B(n20138), .Z(n20140) );
  XOR U23026 ( .A(n20510), .B(n20511), .Z(n20138) );
  AND U23027 ( .A(n20512), .B(n20513), .Z(n20510) );
  AND U23028 ( .A(a[28]), .B(b[44]), .Z(n20509) );
  XOR U23029 ( .A(n20514), .B(n20143), .Z(n20145) );
  XOR U23030 ( .A(n20515), .B(n20516), .Z(n20143) );
  AND U23031 ( .A(n20517), .B(n20518), .Z(n20515) );
  AND U23032 ( .A(a[29]), .B(b[43]), .Z(n20514) );
  XOR U23033 ( .A(n20519), .B(n20148), .Z(n20150) );
  XOR U23034 ( .A(n20520), .B(n20521), .Z(n20148) );
  AND U23035 ( .A(n20522), .B(n20523), .Z(n20520) );
  AND U23036 ( .A(a[30]), .B(b[42]), .Z(n20519) );
  XOR U23037 ( .A(n20524), .B(n20153), .Z(n20155) );
  XOR U23038 ( .A(n20525), .B(n20526), .Z(n20153) );
  AND U23039 ( .A(n20527), .B(n20528), .Z(n20525) );
  AND U23040 ( .A(a[31]), .B(b[41]), .Z(n20524) );
  XOR U23041 ( .A(n20529), .B(n20158), .Z(n20160) );
  XOR U23042 ( .A(n20530), .B(n20531), .Z(n20158) );
  AND U23043 ( .A(n20532), .B(n20533), .Z(n20530) );
  AND U23044 ( .A(a[32]), .B(b[40]), .Z(n20529) );
  XOR U23045 ( .A(n20534), .B(n20163), .Z(n20165) );
  XOR U23046 ( .A(n20535), .B(n20536), .Z(n20163) );
  AND U23047 ( .A(n20537), .B(n20538), .Z(n20535) );
  AND U23048 ( .A(a[33]), .B(b[39]), .Z(n20534) );
  XOR U23049 ( .A(n20539), .B(n20168), .Z(n20170) );
  XOR U23050 ( .A(n20540), .B(n20541), .Z(n20168) );
  AND U23051 ( .A(n20542), .B(n20543), .Z(n20540) );
  AND U23052 ( .A(a[34]), .B(b[38]), .Z(n20539) );
  XOR U23053 ( .A(n20544), .B(n20545), .Z(n20172) );
  AND U23054 ( .A(n20546), .B(n20547), .Z(n20544) );
  XOR U23055 ( .A(n20548), .B(n20177), .Z(n20179) );
  XOR U23056 ( .A(n20549), .B(n20550), .Z(n20177) );
  AND U23057 ( .A(n20551), .B(n20552), .Z(n20549) );
  AND U23058 ( .A(a[35]), .B(b[37]), .Z(n20548) );
  XOR U23059 ( .A(n20554), .B(n20555), .Z(n20182) );
  AND U23060 ( .A(n20556), .B(n20557), .Z(n20554) );
  AND U23061 ( .A(b[35]), .B(a[37]), .Z(n20553) );
  XOR U23062 ( .A(n20559), .B(n20560), .Z(n20187) );
  AND U23063 ( .A(n20561), .B(n20562), .Z(n20559) );
  AND U23064 ( .A(b[34]), .B(a[38]), .Z(n20558) );
  XOR U23065 ( .A(n20564), .B(n20565), .Z(n20192) );
  AND U23066 ( .A(n20566), .B(n20567), .Z(n20564) );
  AND U23067 ( .A(b[33]), .B(a[39]), .Z(n20563) );
  XOR U23068 ( .A(n20569), .B(n20570), .Z(n20197) );
  AND U23069 ( .A(n20571), .B(n20572), .Z(n20569) );
  AND U23070 ( .A(b[32]), .B(a[40]), .Z(n20568) );
  XOR U23071 ( .A(n20574), .B(n20575), .Z(n20202) );
  AND U23072 ( .A(n20576), .B(n20577), .Z(n20574) );
  AND U23073 ( .A(b[31]), .B(a[41]), .Z(n20573) );
  XOR U23074 ( .A(n20579), .B(n20580), .Z(n20207) );
  AND U23075 ( .A(n20581), .B(n20582), .Z(n20579) );
  AND U23076 ( .A(b[30]), .B(a[42]), .Z(n20578) );
  XOR U23077 ( .A(n20584), .B(n20585), .Z(n20212) );
  AND U23078 ( .A(n20586), .B(n20587), .Z(n20584) );
  AND U23079 ( .A(b[29]), .B(a[43]), .Z(n20583) );
  XOR U23080 ( .A(n20589), .B(n20590), .Z(n20217) );
  AND U23081 ( .A(n20591), .B(n20592), .Z(n20589) );
  AND U23082 ( .A(b[28]), .B(a[44]), .Z(n20588) );
  XOR U23083 ( .A(n20594), .B(n20595), .Z(n20222) );
  AND U23084 ( .A(n20596), .B(n20597), .Z(n20594) );
  AND U23085 ( .A(b[27]), .B(a[45]), .Z(n20593) );
  XOR U23086 ( .A(n20599), .B(n20600), .Z(n20227) );
  AND U23087 ( .A(n20601), .B(n20602), .Z(n20599) );
  AND U23088 ( .A(b[26]), .B(a[46]), .Z(n20598) );
  XOR U23089 ( .A(n20604), .B(n20605), .Z(n20232) );
  AND U23090 ( .A(n20606), .B(n20607), .Z(n20604) );
  AND U23091 ( .A(b[25]), .B(a[47]), .Z(n20603) );
  XOR U23092 ( .A(n20609), .B(n20610), .Z(n20237) );
  AND U23093 ( .A(n20611), .B(n20612), .Z(n20609) );
  AND U23094 ( .A(b[24]), .B(a[48]), .Z(n20608) );
  XOR U23095 ( .A(n20614), .B(n20615), .Z(n20242) );
  AND U23096 ( .A(n20616), .B(n20617), .Z(n20614) );
  AND U23097 ( .A(b[23]), .B(a[49]), .Z(n20613) );
  XOR U23098 ( .A(n20619), .B(n20620), .Z(n20247) );
  AND U23099 ( .A(n20621), .B(n20622), .Z(n20619) );
  AND U23100 ( .A(b[22]), .B(a[50]), .Z(n20618) );
  XOR U23101 ( .A(n20624), .B(n20625), .Z(n20252) );
  AND U23102 ( .A(n20626), .B(n20627), .Z(n20624) );
  AND U23103 ( .A(b[21]), .B(a[51]), .Z(n20623) );
  XOR U23104 ( .A(n20629), .B(n20630), .Z(n20257) );
  AND U23105 ( .A(n20631), .B(n20632), .Z(n20629) );
  AND U23106 ( .A(b[20]), .B(a[52]), .Z(n20628) );
  XOR U23107 ( .A(n20634), .B(n20635), .Z(n20262) );
  AND U23108 ( .A(n20636), .B(n20637), .Z(n20634) );
  AND U23109 ( .A(b[19]), .B(a[53]), .Z(n20633) );
  XOR U23110 ( .A(n20639), .B(n20640), .Z(n20267) );
  AND U23111 ( .A(n20641), .B(n20642), .Z(n20639) );
  AND U23112 ( .A(b[18]), .B(a[54]), .Z(n20638) );
  XOR U23113 ( .A(n20644), .B(n20645), .Z(n20272) );
  AND U23114 ( .A(n20646), .B(n20647), .Z(n20644) );
  AND U23115 ( .A(b[17]), .B(a[55]), .Z(n20643) );
  XOR U23116 ( .A(n20649), .B(n20650), .Z(n20277) );
  AND U23117 ( .A(n20651), .B(n20652), .Z(n20649) );
  AND U23118 ( .A(b[16]), .B(a[56]), .Z(n20648) );
  XOR U23119 ( .A(n20654), .B(n20655), .Z(n20282) );
  AND U23120 ( .A(n20656), .B(n20657), .Z(n20654) );
  AND U23121 ( .A(b[15]), .B(a[57]), .Z(n20653) );
  XOR U23122 ( .A(n20659), .B(n20660), .Z(n20287) );
  AND U23123 ( .A(n20661), .B(n20662), .Z(n20659) );
  AND U23124 ( .A(b[14]), .B(a[58]), .Z(n20658) );
  XOR U23125 ( .A(n20664), .B(n20665), .Z(n20292) );
  AND U23126 ( .A(n20666), .B(n20667), .Z(n20664) );
  AND U23127 ( .A(b[13]), .B(a[59]), .Z(n20663) );
  XOR U23128 ( .A(n20669), .B(n20670), .Z(n20297) );
  AND U23129 ( .A(n20671), .B(n20672), .Z(n20669) );
  AND U23130 ( .A(b[12]), .B(a[60]), .Z(n20668) );
  XOR U23131 ( .A(n20674), .B(n20675), .Z(n20302) );
  AND U23132 ( .A(n20676), .B(n20677), .Z(n20674) );
  AND U23133 ( .A(b[11]), .B(a[61]), .Z(n20673) );
  XOR U23134 ( .A(n20679), .B(n20680), .Z(n20307) );
  AND U23135 ( .A(n20681), .B(n20682), .Z(n20679) );
  AND U23136 ( .A(b[10]), .B(a[62]), .Z(n20678) );
  XOR U23137 ( .A(n20684), .B(n20685), .Z(n20312) );
  AND U23138 ( .A(n20686), .B(n20687), .Z(n20684) );
  AND U23139 ( .A(b[9]), .B(a[63]), .Z(n20683) );
  XOR U23140 ( .A(n20689), .B(n20690), .Z(n20317) );
  AND U23141 ( .A(n20691), .B(n20692), .Z(n20689) );
  AND U23142 ( .A(b[8]), .B(a[64]), .Z(n20688) );
  XOR U23143 ( .A(n20694), .B(n20695), .Z(n20322) );
  AND U23144 ( .A(n20696), .B(n20697), .Z(n20694) );
  AND U23145 ( .A(b[7]), .B(a[65]), .Z(n20693) );
  XOR U23146 ( .A(n20699), .B(n20700), .Z(n20327) );
  AND U23147 ( .A(n20701), .B(n20702), .Z(n20699) );
  AND U23148 ( .A(b[6]), .B(a[66]), .Z(n20698) );
  XOR U23149 ( .A(n20704), .B(n20705), .Z(n20332) );
  AND U23150 ( .A(n20706), .B(n20707), .Z(n20704) );
  AND U23151 ( .A(b[5]), .B(a[67]), .Z(n20703) );
  XOR U23152 ( .A(n20709), .B(n20710), .Z(n20337) );
  AND U23153 ( .A(n20711), .B(n20712), .Z(n20709) );
  AND U23154 ( .A(b[4]), .B(a[68]), .Z(n20708) );
  XOR U23155 ( .A(n20714), .B(n20715), .Z(n20342) );
  AND U23156 ( .A(n20716), .B(n20717), .Z(n20714) );
  AND U23157 ( .A(b[3]), .B(a[69]), .Z(n20713) );
  XOR U23158 ( .A(n20719), .B(n20720), .Z(n20347) );
  OR U23159 ( .A(n20721), .B(n20722), .Z(n20720) );
  AND U23160 ( .A(b[2]), .B(a[70]), .Z(n20718) );
  XNOR U23161 ( .A(n20357), .B(n20723), .Z(n20353) );
  NAND U23162 ( .A(b[1]), .B(a[71]), .Z(n20723) );
  IV U23163 ( .A(n20351), .Z(n20357) );
  ANDN U23164 ( .B(n10338), .A(n10340), .Z(n20351) );
  NAND U23165 ( .A(a[71]), .B(b[0]), .Z(n10340) );
  XOR U23166 ( .A(n20721), .B(n20722), .Z(n10338) );
  XOR U23167 ( .A(n20725), .B(n20716), .Z(n20724) );
  XOR U23168 ( .A(n20711), .B(n20715), .Z(n20726) );
  XOR U23169 ( .A(n20706), .B(n20710), .Z(n20727) );
  XOR U23170 ( .A(n20701), .B(n20705), .Z(n20728) );
  XOR U23171 ( .A(n20696), .B(n20700), .Z(n20729) );
  XOR U23172 ( .A(n20691), .B(n20695), .Z(n20730) );
  XOR U23173 ( .A(n20686), .B(n20690), .Z(n20731) );
  XOR U23174 ( .A(n20681), .B(n20685), .Z(n20732) );
  XOR U23175 ( .A(n20676), .B(n20680), .Z(n20733) );
  XOR U23176 ( .A(n20671), .B(n20675), .Z(n20734) );
  XOR U23177 ( .A(n20666), .B(n20670), .Z(n20735) );
  XOR U23178 ( .A(n20661), .B(n20665), .Z(n20736) );
  XOR U23179 ( .A(n20656), .B(n20660), .Z(n20737) );
  XOR U23180 ( .A(n20651), .B(n20655), .Z(n20738) );
  XOR U23181 ( .A(n20646), .B(n20650), .Z(n20739) );
  XOR U23182 ( .A(n20641), .B(n20645), .Z(n20740) );
  XOR U23183 ( .A(n20636), .B(n20640), .Z(n20741) );
  XOR U23184 ( .A(n20631), .B(n20635), .Z(n20742) );
  XOR U23185 ( .A(n20626), .B(n20630), .Z(n20743) );
  XOR U23186 ( .A(n20621), .B(n20625), .Z(n20744) );
  XOR U23187 ( .A(n20616), .B(n20620), .Z(n20745) );
  XOR U23188 ( .A(n20611), .B(n20615), .Z(n20746) );
  XOR U23189 ( .A(n20606), .B(n20610), .Z(n20747) );
  XOR U23190 ( .A(n20601), .B(n20605), .Z(n20748) );
  XOR U23191 ( .A(n20596), .B(n20600), .Z(n20749) );
  XOR U23192 ( .A(n20591), .B(n20595), .Z(n20750) );
  XOR U23193 ( .A(n20586), .B(n20590), .Z(n20751) );
  XOR U23194 ( .A(n20581), .B(n20585), .Z(n20752) );
  XOR U23195 ( .A(n20576), .B(n20580), .Z(n20753) );
  XOR U23196 ( .A(n20571), .B(n20575), .Z(n20754) );
  XOR U23197 ( .A(n20566), .B(n20570), .Z(n20755) );
  XOR U23198 ( .A(n20561), .B(n20565), .Z(n20756) );
  XOR U23199 ( .A(n20556), .B(n20560), .Z(n20757) );
  XOR U23200 ( .A(n20546), .B(n20555), .Z(n20758) );
  XOR U23201 ( .A(n20759), .B(n20545), .Z(n20546) );
  AND U23202 ( .A(b[35]), .B(a[36]), .Z(n20759) );
  XNOR U23203 ( .A(n20545), .B(n20551), .Z(n20760) );
  XNOR U23204 ( .A(n20550), .B(n20542), .Z(n20761) );
  XNOR U23205 ( .A(n20541), .B(n20537), .Z(n20762) );
  XNOR U23206 ( .A(n20536), .B(n20532), .Z(n20763) );
  XNOR U23207 ( .A(n20531), .B(n20527), .Z(n20764) );
  XNOR U23208 ( .A(n20526), .B(n20522), .Z(n20765) );
  XNOR U23209 ( .A(n20521), .B(n20517), .Z(n20766) );
  XNOR U23210 ( .A(n20516), .B(n20512), .Z(n20767) );
  XNOR U23211 ( .A(n20511), .B(n20507), .Z(n20768) );
  XNOR U23212 ( .A(n20506), .B(n20502), .Z(n20769) );
  XNOR U23213 ( .A(n20501), .B(n20497), .Z(n20770) );
  XNOR U23214 ( .A(n20496), .B(n20492), .Z(n20771) );
  XNOR U23215 ( .A(n20491), .B(n20487), .Z(n20772) );
  XNOR U23216 ( .A(n20486), .B(n20482), .Z(n20773) );
  XNOR U23217 ( .A(n20481), .B(n20477), .Z(n20774) );
  XNOR U23218 ( .A(n20476), .B(n20472), .Z(n20775) );
  XNOR U23219 ( .A(n20471), .B(n20467), .Z(n20776) );
  XNOR U23220 ( .A(n20466), .B(n20462), .Z(n20777) );
  XNOR U23221 ( .A(n20461), .B(n20457), .Z(n20778) );
  XNOR U23222 ( .A(n20456), .B(n20452), .Z(n20779) );
  XNOR U23223 ( .A(n20451), .B(n20447), .Z(n20780) );
  XNOR U23224 ( .A(n20446), .B(n20442), .Z(n20781) );
  XNOR U23225 ( .A(n20441), .B(n20437), .Z(n20782) );
  XNOR U23226 ( .A(n20436), .B(n20432), .Z(n20783) );
  XOR U23227 ( .A(n20431), .B(n20428), .Z(n20784) );
  XOR U23228 ( .A(n20785), .B(n20786), .Z(n20428) );
  XOR U23229 ( .A(n20426), .B(n20787), .Z(n20786) );
  XOR U23230 ( .A(n20788), .B(n20789), .Z(n20787) );
  XOR U23231 ( .A(n20790), .B(n20791), .Z(n20789) );
  NAND U23232 ( .A(a[9]), .B(b[62]), .Z(n20791) );
  AND U23233 ( .A(a[8]), .B(b[63]), .Z(n20790) );
  XOR U23234 ( .A(n20792), .B(n20788), .Z(n20785) );
  XOR U23235 ( .A(n20793), .B(n20794), .Z(n20788) );
  ANDN U23236 ( .B(n20795), .A(n20796), .Z(n20793) );
  AND U23237 ( .A(a[10]), .B(b[61]), .Z(n20792) );
  XOR U23238 ( .A(n20797), .B(n20426), .Z(n20427) );
  XOR U23239 ( .A(n20798), .B(n20799), .Z(n20426) );
  AND U23240 ( .A(n20800), .B(n20801), .Z(n20798) );
  AND U23241 ( .A(a[11]), .B(b[60]), .Z(n20797) );
  XOR U23242 ( .A(n20802), .B(n20431), .Z(n20433) );
  XOR U23243 ( .A(n20803), .B(n20804), .Z(n20431) );
  AND U23244 ( .A(n20805), .B(n20806), .Z(n20803) );
  AND U23245 ( .A(a[12]), .B(b[59]), .Z(n20802) );
  XOR U23246 ( .A(n20807), .B(n20436), .Z(n20438) );
  XOR U23247 ( .A(n20808), .B(n20809), .Z(n20436) );
  AND U23248 ( .A(n20810), .B(n20811), .Z(n20808) );
  AND U23249 ( .A(a[13]), .B(b[58]), .Z(n20807) );
  XOR U23250 ( .A(n20812), .B(n20441), .Z(n20443) );
  XOR U23251 ( .A(n20813), .B(n20814), .Z(n20441) );
  AND U23252 ( .A(n20815), .B(n20816), .Z(n20813) );
  AND U23253 ( .A(a[14]), .B(b[57]), .Z(n20812) );
  XOR U23254 ( .A(n20817), .B(n20446), .Z(n20448) );
  XOR U23255 ( .A(n20818), .B(n20819), .Z(n20446) );
  AND U23256 ( .A(n20820), .B(n20821), .Z(n20818) );
  AND U23257 ( .A(a[15]), .B(b[56]), .Z(n20817) );
  XOR U23258 ( .A(n20822), .B(n20451), .Z(n20453) );
  XOR U23259 ( .A(n20823), .B(n20824), .Z(n20451) );
  AND U23260 ( .A(n20825), .B(n20826), .Z(n20823) );
  AND U23261 ( .A(a[16]), .B(b[55]), .Z(n20822) );
  XOR U23262 ( .A(n20827), .B(n20456), .Z(n20458) );
  XOR U23263 ( .A(n20828), .B(n20829), .Z(n20456) );
  AND U23264 ( .A(n20830), .B(n20831), .Z(n20828) );
  AND U23265 ( .A(a[17]), .B(b[54]), .Z(n20827) );
  XOR U23266 ( .A(n20832), .B(n20461), .Z(n20463) );
  XOR U23267 ( .A(n20833), .B(n20834), .Z(n20461) );
  AND U23268 ( .A(n20835), .B(n20836), .Z(n20833) );
  AND U23269 ( .A(a[18]), .B(b[53]), .Z(n20832) );
  XOR U23270 ( .A(n20837), .B(n20466), .Z(n20468) );
  XOR U23271 ( .A(n20838), .B(n20839), .Z(n20466) );
  AND U23272 ( .A(n20840), .B(n20841), .Z(n20838) );
  AND U23273 ( .A(a[19]), .B(b[52]), .Z(n20837) );
  XOR U23274 ( .A(n20842), .B(n20471), .Z(n20473) );
  XOR U23275 ( .A(n20843), .B(n20844), .Z(n20471) );
  AND U23276 ( .A(n20845), .B(n20846), .Z(n20843) );
  AND U23277 ( .A(a[20]), .B(b[51]), .Z(n20842) );
  XOR U23278 ( .A(n20847), .B(n20476), .Z(n20478) );
  XOR U23279 ( .A(n20848), .B(n20849), .Z(n20476) );
  AND U23280 ( .A(n20850), .B(n20851), .Z(n20848) );
  AND U23281 ( .A(a[21]), .B(b[50]), .Z(n20847) );
  XOR U23282 ( .A(n20852), .B(n20481), .Z(n20483) );
  XOR U23283 ( .A(n20853), .B(n20854), .Z(n20481) );
  AND U23284 ( .A(n20855), .B(n20856), .Z(n20853) );
  AND U23285 ( .A(a[22]), .B(b[49]), .Z(n20852) );
  XOR U23286 ( .A(n20857), .B(n20486), .Z(n20488) );
  XOR U23287 ( .A(n20858), .B(n20859), .Z(n20486) );
  AND U23288 ( .A(n20860), .B(n20861), .Z(n20858) );
  AND U23289 ( .A(a[23]), .B(b[48]), .Z(n20857) );
  XOR U23290 ( .A(n20862), .B(n20491), .Z(n20493) );
  XOR U23291 ( .A(n20863), .B(n20864), .Z(n20491) );
  AND U23292 ( .A(n20865), .B(n20866), .Z(n20863) );
  AND U23293 ( .A(a[24]), .B(b[47]), .Z(n20862) );
  XOR U23294 ( .A(n20867), .B(n20496), .Z(n20498) );
  XOR U23295 ( .A(n20868), .B(n20869), .Z(n20496) );
  AND U23296 ( .A(n20870), .B(n20871), .Z(n20868) );
  AND U23297 ( .A(a[25]), .B(b[46]), .Z(n20867) );
  XOR U23298 ( .A(n20872), .B(n20501), .Z(n20503) );
  XOR U23299 ( .A(n20873), .B(n20874), .Z(n20501) );
  AND U23300 ( .A(n20875), .B(n20876), .Z(n20873) );
  AND U23301 ( .A(a[26]), .B(b[45]), .Z(n20872) );
  XOR U23302 ( .A(n20877), .B(n20506), .Z(n20508) );
  XOR U23303 ( .A(n20878), .B(n20879), .Z(n20506) );
  AND U23304 ( .A(n20880), .B(n20881), .Z(n20878) );
  AND U23305 ( .A(a[27]), .B(b[44]), .Z(n20877) );
  XOR U23306 ( .A(n20882), .B(n20511), .Z(n20513) );
  XOR U23307 ( .A(n20883), .B(n20884), .Z(n20511) );
  AND U23308 ( .A(n20885), .B(n20886), .Z(n20883) );
  AND U23309 ( .A(a[28]), .B(b[43]), .Z(n20882) );
  XOR U23310 ( .A(n20887), .B(n20516), .Z(n20518) );
  XOR U23311 ( .A(n20888), .B(n20889), .Z(n20516) );
  AND U23312 ( .A(n20890), .B(n20891), .Z(n20888) );
  AND U23313 ( .A(a[29]), .B(b[42]), .Z(n20887) );
  XOR U23314 ( .A(n20892), .B(n20521), .Z(n20523) );
  XOR U23315 ( .A(n20893), .B(n20894), .Z(n20521) );
  AND U23316 ( .A(n20895), .B(n20896), .Z(n20893) );
  AND U23317 ( .A(a[30]), .B(b[41]), .Z(n20892) );
  XOR U23318 ( .A(n20897), .B(n20526), .Z(n20528) );
  XOR U23319 ( .A(n20898), .B(n20899), .Z(n20526) );
  AND U23320 ( .A(n20900), .B(n20901), .Z(n20898) );
  AND U23321 ( .A(a[31]), .B(b[40]), .Z(n20897) );
  XOR U23322 ( .A(n20902), .B(n20531), .Z(n20533) );
  XOR U23323 ( .A(n20903), .B(n20904), .Z(n20531) );
  AND U23324 ( .A(n20905), .B(n20906), .Z(n20903) );
  AND U23325 ( .A(a[32]), .B(b[39]), .Z(n20902) );
  XOR U23326 ( .A(n20907), .B(n20536), .Z(n20538) );
  XOR U23327 ( .A(n20908), .B(n20909), .Z(n20536) );
  AND U23328 ( .A(n20910), .B(n20911), .Z(n20908) );
  AND U23329 ( .A(a[33]), .B(b[38]), .Z(n20907) );
  XOR U23330 ( .A(n20912), .B(n20541), .Z(n20543) );
  XOR U23331 ( .A(n20913), .B(n20914), .Z(n20541) );
  AND U23332 ( .A(n20915), .B(n20916), .Z(n20913) );
  AND U23333 ( .A(a[34]), .B(b[37]), .Z(n20912) );
  XOR U23334 ( .A(n20917), .B(n20918), .Z(n20545) );
  AND U23335 ( .A(n20919), .B(n20920), .Z(n20917) );
  XOR U23336 ( .A(n20921), .B(n20550), .Z(n20552) );
  XOR U23337 ( .A(n20922), .B(n20923), .Z(n20550) );
  AND U23338 ( .A(n20924), .B(n20925), .Z(n20922) );
  AND U23339 ( .A(a[35]), .B(b[36]), .Z(n20921) );
  XOR U23340 ( .A(n20927), .B(n20928), .Z(n20555) );
  AND U23341 ( .A(n20929), .B(n20930), .Z(n20927) );
  AND U23342 ( .A(b[34]), .B(a[37]), .Z(n20926) );
  XOR U23343 ( .A(n20932), .B(n20933), .Z(n20560) );
  AND U23344 ( .A(n20934), .B(n20935), .Z(n20932) );
  AND U23345 ( .A(b[33]), .B(a[38]), .Z(n20931) );
  XOR U23346 ( .A(n20937), .B(n20938), .Z(n20565) );
  AND U23347 ( .A(n20939), .B(n20940), .Z(n20937) );
  AND U23348 ( .A(b[32]), .B(a[39]), .Z(n20936) );
  XOR U23349 ( .A(n20942), .B(n20943), .Z(n20570) );
  AND U23350 ( .A(n20944), .B(n20945), .Z(n20942) );
  AND U23351 ( .A(b[31]), .B(a[40]), .Z(n20941) );
  XOR U23352 ( .A(n20947), .B(n20948), .Z(n20575) );
  AND U23353 ( .A(n20949), .B(n20950), .Z(n20947) );
  AND U23354 ( .A(b[30]), .B(a[41]), .Z(n20946) );
  XOR U23355 ( .A(n20952), .B(n20953), .Z(n20580) );
  AND U23356 ( .A(n20954), .B(n20955), .Z(n20952) );
  AND U23357 ( .A(b[29]), .B(a[42]), .Z(n20951) );
  XOR U23358 ( .A(n20957), .B(n20958), .Z(n20585) );
  AND U23359 ( .A(n20959), .B(n20960), .Z(n20957) );
  AND U23360 ( .A(b[28]), .B(a[43]), .Z(n20956) );
  XOR U23361 ( .A(n20962), .B(n20963), .Z(n20590) );
  AND U23362 ( .A(n20964), .B(n20965), .Z(n20962) );
  AND U23363 ( .A(b[27]), .B(a[44]), .Z(n20961) );
  XOR U23364 ( .A(n20967), .B(n20968), .Z(n20595) );
  AND U23365 ( .A(n20969), .B(n20970), .Z(n20967) );
  AND U23366 ( .A(b[26]), .B(a[45]), .Z(n20966) );
  XOR U23367 ( .A(n20972), .B(n20973), .Z(n20600) );
  AND U23368 ( .A(n20974), .B(n20975), .Z(n20972) );
  AND U23369 ( .A(b[25]), .B(a[46]), .Z(n20971) );
  XOR U23370 ( .A(n20977), .B(n20978), .Z(n20605) );
  AND U23371 ( .A(n20979), .B(n20980), .Z(n20977) );
  AND U23372 ( .A(b[24]), .B(a[47]), .Z(n20976) );
  XOR U23373 ( .A(n20982), .B(n20983), .Z(n20610) );
  AND U23374 ( .A(n20984), .B(n20985), .Z(n20982) );
  AND U23375 ( .A(b[23]), .B(a[48]), .Z(n20981) );
  XOR U23376 ( .A(n20987), .B(n20988), .Z(n20615) );
  AND U23377 ( .A(n20989), .B(n20990), .Z(n20987) );
  AND U23378 ( .A(b[22]), .B(a[49]), .Z(n20986) );
  XOR U23379 ( .A(n20992), .B(n20993), .Z(n20620) );
  AND U23380 ( .A(n20994), .B(n20995), .Z(n20992) );
  AND U23381 ( .A(b[21]), .B(a[50]), .Z(n20991) );
  XOR U23382 ( .A(n20997), .B(n20998), .Z(n20625) );
  AND U23383 ( .A(n20999), .B(n21000), .Z(n20997) );
  AND U23384 ( .A(b[20]), .B(a[51]), .Z(n20996) );
  XOR U23385 ( .A(n21002), .B(n21003), .Z(n20630) );
  AND U23386 ( .A(n21004), .B(n21005), .Z(n21002) );
  AND U23387 ( .A(b[19]), .B(a[52]), .Z(n21001) );
  XOR U23388 ( .A(n21007), .B(n21008), .Z(n20635) );
  AND U23389 ( .A(n21009), .B(n21010), .Z(n21007) );
  AND U23390 ( .A(b[18]), .B(a[53]), .Z(n21006) );
  XOR U23391 ( .A(n21012), .B(n21013), .Z(n20640) );
  AND U23392 ( .A(n21014), .B(n21015), .Z(n21012) );
  AND U23393 ( .A(b[17]), .B(a[54]), .Z(n21011) );
  XOR U23394 ( .A(n21017), .B(n21018), .Z(n20645) );
  AND U23395 ( .A(n21019), .B(n21020), .Z(n21017) );
  AND U23396 ( .A(b[16]), .B(a[55]), .Z(n21016) );
  XOR U23397 ( .A(n21022), .B(n21023), .Z(n20650) );
  AND U23398 ( .A(n21024), .B(n21025), .Z(n21022) );
  AND U23399 ( .A(b[15]), .B(a[56]), .Z(n21021) );
  XOR U23400 ( .A(n21027), .B(n21028), .Z(n20655) );
  AND U23401 ( .A(n21029), .B(n21030), .Z(n21027) );
  AND U23402 ( .A(b[14]), .B(a[57]), .Z(n21026) );
  XOR U23403 ( .A(n21032), .B(n21033), .Z(n20660) );
  AND U23404 ( .A(n21034), .B(n21035), .Z(n21032) );
  AND U23405 ( .A(b[13]), .B(a[58]), .Z(n21031) );
  XOR U23406 ( .A(n21037), .B(n21038), .Z(n20665) );
  AND U23407 ( .A(n21039), .B(n21040), .Z(n21037) );
  AND U23408 ( .A(b[12]), .B(a[59]), .Z(n21036) );
  XOR U23409 ( .A(n21042), .B(n21043), .Z(n20670) );
  AND U23410 ( .A(n21044), .B(n21045), .Z(n21042) );
  AND U23411 ( .A(b[11]), .B(a[60]), .Z(n21041) );
  XOR U23412 ( .A(n21047), .B(n21048), .Z(n20675) );
  AND U23413 ( .A(n21049), .B(n21050), .Z(n21047) );
  AND U23414 ( .A(b[10]), .B(a[61]), .Z(n21046) );
  XOR U23415 ( .A(n21052), .B(n21053), .Z(n20680) );
  AND U23416 ( .A(n21054), .B(n21055), .Z(n21052) );
  AND U23417 ( .A(b[9]), .B(a[62]), .Z(n21051) );
  XOR U23418 ( .A(n21057), .B(n21058), .Z(n20685) );
  AND U23419 ( .A(n21059), .B(n21060), .Z(n21057) );
  AND U23420 ( .A(b[8]), .B(a[63]), .Z(n21056) );
  XOR U23421 ( .A(n21062), .B(n21063), .Z(n20690) );
  AND U23422 ( .A(n21064), .B(n21065), .Z(n21062) );
  AND U23423 ( .A(b[7]), .B(a[64]), .Z(n21061) );
  XOR U23424 ( .A(n21067), .B(n21068), .Z(n20695) );
  AND U23425 ( .A(n21069), .B(n21070), .Z(n21067) );
  AND U23426 ( .A(b[6]), .B(a[65]), .Z(n21066) );
  XOR U23427 ( .A(n21072), .B(n21073), .Z(n20700) );
  AND U23428 ( .A(n21074), .B(n21075), .Z(n21072) );
  AND U23429 ( .A(b[5]), .B(a[66]), .Z(n21071) );
  XOR U23430 ( .A(n21077), .B(n21078), .Z(n20705) );
  AND U23431 ( .A(n21079), .B(n21080), .Z(n21077) );
  AND U23432 ( .A(b[4]), .B(a[67]), .Z(n21076) );
  XOR U23433 ( .A(n21082), .B(n21083), .Z(n20710) );
  AND U23434 ( .A(n21084), .B(n21085), .Z(n21082) );
  AND U23435 ( .A(b[3]), .B(a[68]), .Z(n21081) );
  XOR U23436 ( .A(n21087), .B(n21088), .Z(n20715) );
  OR U23437 ( .A(n21089), .B(n21090), .Z(n21088) );
  AND U23438 ( .A(b[2]), .B(a[69]), .Z(n21086) );
  XNOR U23439 ( .A(n20725), .B(n21091), .Z(n20721) );
  NAND U23440 ( .A(b[1]), .B(a[70]), .Z(n21091) );
  IV U23441 ( .A(n20719), .Z(n20725) );
  ANDN U23442 ( .B(n10341), .A(n10343), .Z(n20719) );
  NAND U23443 ( .A(a[70]), .B(b[0]), .Z(n10343) );
  XOR U23444 ( .A(n21089), .B(n21090), .Z(n10341) );
  XOR U23445 ( .A(n21093), .B(n21084), .Z(n21092) );
  XOR U23446 ( .A(n21079), .B(n21083), .Z(n21094) );
  XOR U23447 ( .A(n21074), .B(n21078), .Z(n21095) );
  XOR U23448 ( .A(n21069), .B(n21073), .Z(n21096) );
  XOR U23449 ( .A(n21064), .B(n21068), .Z(n21097) );
  XOR U23450 ( .A(n21059), .B(n21063), .Z(n21098) );
  XOR U23451 ( .A(n21054), .B(n21058), .Z(n21099) );
  XOR U23452 ( .A(n21049), .B(n21053), .Z(n21100) );
  XOR U23453 ( .A(n21044), .B(n21048), .Z(n21101) );
  XOR U23454 ( .A(n21039), .B(n21043), .Z(n21102) );
  XOR U23455 ( .A(n21034), .B(n21038), .Z(n21103) );
  XOR U23456 ( .A(n21029), .B(n21033), .Z(n21104) );
  XOR U23457 ( .A(n21024), .B(n21028), .Z(n21105) );
  XOR U23458 ( .A(n21019), .B(n21023), .Z(n21106) );
  XOR U23459 ( .A(n21014), .B(n21018), .Z(n21107) );
  XOR U23460 ( .A(n21009), .B(n21013), .Z(n21108) );
  XOR U23461 ( .A(n21004), .B(n21008), .Z(n21109) );
  XOR U23462 ( .A(n20999), .B(n21003), .Z(n21110) );
  XOR U23463 ( .A(n20994), .B(n20998), .Z(n21111) );
  XOR U23464 ( .A(n20989), .B(n20993), .Z(n21112) );
  XOR U23465 ( .A(n20984), .B(n20988), .Z(n21113) );
  XOR U23466 ( .A(n20979), .B(n20983), .Z(n21114) );
  XOR U23467 ( .A(n20974), .B(n20978), .Z(n21115) );
  XOR U23468 ( .A(n20969), .B(n20973), .Z(n21116) );
  XOR U23469 ( .A(n20964), .B(n20968), .Z(n21117) );
  XOR U23470 ( .A(n20959), .B(n20963), .Z(n21118) );
  XOR U23471 ( .A(n20954), .B(n20958), .Z(n21119) );
  XOR U23472 ( .A(n20949), .B(n20953), .Z(n21120) );
  XOR U23473 ( .A(n20944), .B(n20948), .Z(n21121) );
  XOR U23474 ( .A(n20939), .B(n20943), .Z(n21122) );
  XOR U23475 ( .A(n20934), .B(n20938), .Z(n21123) );
  XOR U23476 ( .A(n20929), .B(n20933), .Z(n21124) );
  XOR U23477 ( .A(n20919), .B(n20928), .Z(n21125) );
  XOR U23478 ( .A(n21126), .B(n20918), .Z(n20919) );
  AND U23479 ( .A(b[34]), .B(a[36]), .Z(n21126) );
  XNOR U23480 ( .A(n20918), .B(n20924), .Z(n21127) );
  XNOR U23481 ( .A(n20923), .B(n20915), .Z(n21128) );
  XNOR U23482 ( .A(n20914), .B(n20910), .Z(n21129) );
  XNOR U23483 ( .A(n20909), .B(n20905), .Z(n21130) );
  XNOR U23484 ( .A(n20904), .B(n20900), .Z(n21131) );
  XNOR U23485 ( .A(n20899), .B(n20895), .Z(n21132) );
  XNOR U23486 ( .A(n20894), .B(n20890), .Z(n21133) );
  XNOR U23487 ( .A(n20889), .B(n20885), .Z(n21134) );
  XNOR U23488 ( .A(n20884), .B(n20880), .Z(n21135) );
  XNOR U23489 ( .A(n20879), .B(n20875), .Z(n21136) );
  XNOR U23490 ( .A(n20874), .B(n20870), .Z(n21137) );
  XNOR U23491 ( .A(n20869), .B(n20865), .Z(n21138) );
  XNOR U23492 ( .A(n20864), .B(n20860), .Z(n21139) );
  XNOR U23493 ( .A(n20859), .B(n20855), .Z(n21140) );
  XNOR U23494 ( .A(n20854), .B(n20850), .Z(n21141) );
  XNOR U23495 ( .A(n20849), .B(n20845), .Z(n21142) );
  XNOR U23496 ( .A(n20844), .B(n20840), .Z(n21143) );
  XNOR U23497 ( .A(n20839), .B(n20835), .Z(n21144) );
  XNOR U23498 ( .A(n20834), .B(n20830), .Z(n21145) );
  XNOR U23499 ( .A(n20829), .B(n20825), .Z(n21146) );
  XNOR U23500 ( .A(n20824), .B(n20820), .Z(n21147) );
  XNOR U23501 ( .A(n20819), .B(n20815), .Z(n21148) );
  XNOR U23502 ( .A(n20814), .B(n20810), .Z(n21149) );
  XNOR U23503 ( .A(n20809), .B(n20805), .Z(n21150) );
  XNOR U23504 ( .A(n20804), .B(n20800), .Z(n21151) );
  XOR U23505 ( .A(n20799), .B(n20796), .Z(n21152) );
  XOR U23506 ( .A(n21153), .B(n21154), .Z(n20796) );
  XOR U23507 ( .A(n20794), .B(n21155), .Z(n21154) );
  XOR U23508 ( .A(n21156), .B(n21157), .Z(n21155) );
  XOR U23509 ( .A(n21158), .B(n21159), .Z(n21157) );
  NAND U23510 ( .A(a[8]), .B(b[62]), .Z(n21159) );
  AND U23511 ( .A(a[7]), .B(b[63]), .Z(n21158) );
  XOR U23512 ( .A(n21160), .B(n21156), .Z(n21153) );
  XOR U23513 ( .A(n21161), .B(n21162), .Z(n21156) );
  ANDN U23514 ( .B(n21163), .A(n21164), .Z(n21161) );
  AND U23515 ( .A(a[9]), .B(b[61]), .Z(n21160) );
  XOR U23516 ( .A(n21165), .B(n20794), .Z(n20795) );
  XOR U23517 ( .A(n21166), .B(n21167), .Z(n20794) );
  AND U23518 ( .A(n21168), .B(n21169), .Z(n21166) );
  AND U23519 ( .A(a[10]), .B(b[60]), .Z(n21165) );
  XOR U23520 ( .A(n21170), .B(n20799), .Z(n20801) );
  XOR U23521 ( .A(n21171), .B(n21172), .Z(n20799) );
  AND U23522 ( .A(n21173), .B(n21174), .Z(n21171) );
  AND U23523 ( .A(a[11]), .B(b[59]), .Z(n21170) );
  XOR U23524 ( .A(n21175), .B(n20804), .Z(n20806) );
  XOR U23525 ( .A(n21176), .B(n21177), .Z(n20804) );
  AND U23526 ( .A(n21178), .B(n21179), .Z(n21176) );
  AND U23527 ( .A(a[12]), .B(b[58]), .Z(n21175) );
  XOR U23528 ( .A(n21180), .B(n20809), .Z(n20811) );
  XOR U23529 ( .A(n21181), .B(n21182), .Z(n20809) );
  AND U23530 ( .A(n21183), .B(n21184), .Z(n21181) );
  AND U23531 ( .A(a[13]), .B(b[57]), .Z(n21180) );
  XOR U23532 ( .A(n21185), .B(n20814), .Z(n20816) );
  XOR U23533 ( .A(n21186), .B(n21187), .Z(n20814) );
  AND U23534 ( .A(n21188), .B(n21189), .Z(n21186) );
  AND U23535 ( .A(a[14]), .B(b[56]), .Z(n21185) );
  XOR U23536 ( .A(n21190), .B(n20819), .Z(n20821) );
  XOR U23537 ( .A(n21191), .B(n21192), .Z(n20819) );
  AND U23538 ( .A(n21193), .B(n21194), .Z(n21191) );
  AND U23539 ( .A(a[15]), .B(b[55]), .Z(n21190) );
  XOR U23540 ( .A(n21195), .B(n20824), .Z(n20826) );
  XOR U23541 ( .A(n21196), .B(n21197), .Z(n20824) );
  AND U23542 ( .A(n21198), .B(n21199), .Z(n21196) );
  AND U23543 ( .A(a[16]), .B(b[54]), .Z(n21195) );
  XOR U23544 ( .A(n21200), .B(n20829), .Z(n20831) );
  XOR U23545 ( .A(n21201), .B(n21202), .Z(n20829) );
  AND U23546 ( .A(n21203), .B(n21204), .Z(n21201) );
  AND U23547 ( .A(a[17]), .B(b[53]), .Z(n21200) );
  XOR U23548 ( .A(n21205), .B(n20834), .Z(n20836) );
  XOR U23549 ( .A(n21206), .B(n21207), .Z(n20834) );
  AND U23550 ( .A(n21208), .B(n21209), .Z(n21206) );
  AND U23551 ( .A(a[18]), .B(b[52]), .Z(n21205) );
  XOR U23552 ( .A(n21210), .B(n20839), .Z(n20841) );
  XOR U23553 ( .A(n21211), .B(n21212), .Z(n20839) );
  AND U23554 ( .A(n21213), .B(n21214), .Z(n21211) );
  AND U23555 ( .A(a[19]), .B(b[51]), .Z(n21210) );
  XOR U23556 ( .A(n21215), .B(n20844), .Z(n20846) );
  XOR U23557 ( .A(n21216), .B(n21217), .Z(n20844) );
  AND U23558 ( .A(n21218), .B(n21219), .Z(n21216) );
  AND U23559 ( .A(a[20]), .B(b[50]), .Z(n21215) );
  XOR U23560 ( .A(n21220), .B(n20849), .Z(n20851) );
  XOR U23561 ( .A(n21221), .B(n21222), .Z(n20849) );
  AND U23562 ( .A(n21223), .B(n21224), .Z(n21221) );
  AND U23563 ( .A(a[21]), .B(b[49]), .Z(n21220) );
  XOR U23564 ( .A(n21225), .B(n20854), .Z(n20856) );
  XOR U23565 ( .A(n21226), .B(n21227), .Z(n20854) );
  AND U23566 ( .A(n21228), .B(n21229), .Z(n21226) );
  AND U23567 ( .A(a[22]), .B(b[48]), .Z(n21225) );
  XOR U23568 ( .A(n21230), .B(n20859), .Z(n20861) );
  XOR U23569 ( .A(n21231), .B(n21232), .Z(n20859) );
  AND U23570 ( .A(n21233), .B(n21234), .Z(n21231) );
  AND U23571 ( .A(a[23]), .B(b[47]), .Z(n21230) );
  XOR U23572 ( .A(n21235), .B(n20864), .Z(n20866) );
  XOR U23573 ( .A(n21236), .B(n21237), .Z(n20864) );
  AND U23574 ( .A(n21238), .B(n21239), .Z(n21236) );
  AND U23575 ( .A(a[24]), .B(b[46]), .Z(n21235) );
  XOR U23576 ( .A(n21240), .B(n20869), .Z(n20871) );
  XOR U23577 ( .A(n21241), .B(n21242), .Z(n20869) );
  AND U23578 ( .A(n21243), .B(n21244), .Z(n21241) );
  AND U23579 ( .A(a[25]), .B(b[45]), .Z(n21240) );
  XOR U23580 ( .A(n21245), .B(n20874), .Z(n20876) );
  XOR U23581 ( .A(n21246), .B(n21247), .Z(n20874) );
  AND U23582 ( .A(n21248), .B(n21249), .Z(n21246) );
  AND U23583 ( .A(a[26]), .B(b[44]), .Z(n21245) );
  XOR U23584 ( .A(n21250), .B(n20879), .Z(n20881) );
  XOR U23585 ( .A(n21251), .B(n21252), .Z(n20879) );
  AND U23586 ( .A(n21253), .B(n21254), .Z(n21251) );
  AND U23587 ( .A(a[27]), .B(b[43]), .Z(n21250) );
  XOR U23588 ( .A(n21255), .B(n20884), .Z(n20886) );
  XOR U23589 ( .A(n21256), .B(n21257), .Z(n20884) );
  AND U23590 ( .A(n21258), .B(n21259), .Z(n21256) );
  AND U23591 ( .A(a[28]), .B(b[42]), .Z(n21255) );
  XOR U23592 ( .A(n21260), .B(n20889), .Z(n20891) );
  XOR U23593 ( .A(n21261), .B(n21262), .Z(n20889) );
  AND U23594 ( .A(n21263), .B(n21264), .Z(n21261) );
  AND U23595 ( .A(a[29]), .B(b[41]), .Z(n21260) );
  XOR U23596 ( .A(n21265), .B(n20894), .Z(n20896) );
  XOR U23597 ( .A(n21266), .B(n21267), .Z(n20894) );
  AND U23598 ( .A(n21268), .B(n21269), .Z(n21266) );
  AND U23599 ( .A(a[30]), .B(b[40]), .Z(n21265) );
  XOR U23600 ( .A(n21270), .B(n20899), .Z(n20901) );
  XOR U23601 ( .A(n21271), .B(n21272), .Z(n20899) );
  AND U23602 ( .A(n21273), .B(n21274), .Z(n21271) );
  AND U23603 ( .A(a[31]), .B(b[39]), .Z(n21270) );
  XOR U23604 ( .A(n21275), .B(n20904), .Z(n20906) );
  XOR U23605 ( .A(n21276), .B(n21277), .Z(n20904) );
  AND U23606 ( .A(n21278), .B(n21279), .Z(n21276) );
  AND U23607 ( .A(a[32]), .B(b[38]), .Z(n21275) );
  XOR U23608 ( .A(n21280), .B(n20909), .Z(n20911) );
  XOR U23609 ( .A(n21281), .B(n21282), .Z(n20909) );
  AND U23610 ( .A(n21283), .B(n21284), .Z(n21281) );
  AND U23611 ( .A(a[33]), .B(b[37]), .Z(n21280) );
  XOR U23612 ( .A(n21285), .B(n20914), .Z(n20916) );
  XOR U23613 ( .A(n21286), .B(n21287), .Z(n20914) );
  AND U23614 ( .A(n21288), .B(n21289), .Z(n21286) );
  AND U23615 ( .A(a[34]), .B(b[36]), .Z(n21285) );
  XOR U23616 ( .A(n21290), .B(n21291), .Z(n20918) );
  AND U23617 ( .A(n21292), .B(n21293), .Z(n21290) );
  XOR U23618 ( .A(n21294), .B(n20923), .Z(n20925) );
  XOR U23619 ( .A(n21295), .B(n21296), .Z(n20923) );
  AND U23620 ( .A(n21297), .B(n21298), .Z(n21295) );
  AND U23621 ( .A(a[35]), .B(b[35]), .Z(n21294) );
  XOR U23622 ( .A(n21300), .B(n21301), .Z(n20928) );
  AND U23623 ( .A(n21302), .B(n21303), .Z(n21300) );
  AND U23624 ( .A(b[33]), .B(a[37]), .Z(n21299) );
  XOR U23625 ( .A(n21305), .B(n21306), .Z(n20933) );
  AND U23626 ( .A(n21307), .B(n21308), .Z(n21305) );
  AND U23627 ( .A(b[32]), .B(a[38]), .Z(n21304) );
  XOR U23628 ( .A(n21310), .B(n21311), .Z(n20938) );
  AND U23629 ( .A(n21312), .B(n21313), .Z(n21310) );
  AND U23630 ( .A(b[31]), .B(a[39]), .Z(n21309) );
  XOR U23631 ( .A(n21315), .B(n21316), .Z(n20943) );
  AND U23632 ( .A(n21317), .B(n21318), .Z(n21315) );
  AND U23633 ( .A(b[30]), .B(a[40]), .Z(n21314) );
  XOR U23634 ( .A(n21320), .B(n21321), .Z(n20948) );
  AND U23635 ( .A(n21322), .B(n21323), .Z(n21320) );
  AND U23636 ( .A(b[29]), .B(a[41]), .Z(n21319) );
  XOR U23637 ( .A(n21325), .B(n21326), .Z(n20953) );
  AND U23638 ( .A(n21327), .B(n21328), .Z(n21325) );
  AND U23639 ( .A(b[28]), .B(a[42]), .Z(n21324) );
  XOR U23640 ( .A(n21330), .B(n21331), .Z(n20958) );
  AND U23641 ( .A(n21332), .B(n21333), .Z(n21330) );
  AND U23642 ( .A(b[27]), .B(a[43]), .Z(n21329) );
  XOR U23643 ( .A(n21335), .B(n21336), .Z(n20963) );
  AND U23644 ( .A(n21337), .B(n21338), .Z(n21335) );
  AND U23645 ( .A(b[26]), .B(a[44]), .Z(n21334) );
  XOR U23646 ( .A(n21340), .B(n21341), .Z(n20968) );
  AND U23647 ( .A(n21342), .B(n21343), .Z(n21340) );
  AND U23648 ( .A(b[25]), .B(a[45]), .Z(n21339) );
  XOR U23649 ( .A(n21345), .B(n21346), .Z(n20973) );
  AND U23650 ( .A(n21347), .B(n21348), .Z(n21345) );
  AND U23651 ( .A(b[24]), .B(a[46]), .Z(n21344) );
  XOR U23652 ( .A(n21350), .B(n21351), .Z(n20978) );
  AND U23653 ( .A(n21352), .B(n21353), .Z(n21350) );
  AND U23654 ( .A(b[23]), .B(a[47]), .Z(n21349) );
  XOR U23655 ( .A(n21355), .B(n21356), .Z(n20983) );
  AND U23656 ( .A(n21357), .B(n21358), .Z(n21355) );
  AND U23657 ( .A(b[22]), .B(a[48]), .Z(n21354) );
  XOR U23658 ( .A(n21360), .B(n21361), .Z(n20988) );
  AND U23659 ( .A(n21362), .B(n21363), .Z(n21360) );
  AND U23660 ( .A(b[21]), .B(a[49]), .Z(n21359) );
  XOR U23661 ( .A(n21365), .B(n21366), .Z(n20993) );
  AND U23662 ( .A(n21367), .B(n21368), .Z(n21365) );
  AND U23663 ( .A(b[20]), .B(a[50]), .Z(n21364) );
  XOR U23664 ( .A(n21370), .B(n21371), .Z(n20998) );
  AND U23665 ( .A(n21372), .B(n21373), .Z(n21370) );
  AND U23666 ( .A(b[19]), .B(a[51]), .Z(n21369) );
  XOR U23667 ( .A(n21375), .B(n21376), .Z(n21003) );
  AND U23668 ( .A(n21377), .B(n21378), .Z(n21375) );
  AND U23669 ( .A(b[18]), .B(a[52]), .Z(n21374) );
  XOR U23670 ( .A(n21380), .B(n21381), .Z(n21008) );
  AND U23671 ( .A(n21382), .B(n21383), .Z(n21380) );
  AND U23672 ( .A(b[17]), .B(a[53]), .Z(n21379) );
  XOR U23673 ( .A(n21385), .B(n21386), .Z(n21013) );
  AND U23674 ( .A(n21387), .B(n21388), .Z(n21385) );
  AND U23675 ( .A(b[16]), .B(a[54]), .Z(n21384) );
  XOR U23676 ( .A(n21390), .B(n21391), .Z(n21018) );
  AND U23677 ( .A(n21392), .B(n21393), .Z(n21390) );
  AND U23678 ( .A(b[15]), .B(a[55]), .Z(n21389) );
  XOR U23679 ( .A(n21395), .B(n21396), .Z(n21023) );
  AND U23680 ( .A(n21397), .B(n21398), .Z(n21395) );
  AND U23681 ( .A(b[14]), .B(a[56]), .Z(n21394) );
  XOR U23682 ( .A(n21400), .B(n21401), .Z(n21028) );
  AND U23683 ( .A(n21402), .B(n21403), .Z(n21400) );
  AND U23684 ( .A(b[13]), .B(a[57]), .Z(n21399) );
  XOR U23685 ( .A(n21405), .B(n21406), .Z(n21033) );
  AND U23686 ( .A(n21407), .B(n21408), .Z(n21405) );
  AND U23687 ( .A(b[12]), .B(a[58]), .Z(n21404) );
  XOR U23688 ( .A(n21410), .B(n21411), .Z(n21038) );
  AND U23689 ( .A(n21412), .B(n21413), .Z(n21410) );
  AND U23690 ( .A(b[11]), .B(a[59]), .Z(n21409) );
  XOR U23691 ( .A(n21415), .B(n21416), .Z(n21043) );
  AND U23692 ( .A(n21417), .B(n21418), .Z(n21415) );
  AND U23693 ( .A(b[10]), .B(a[60]), .Z(n21414) );
  XOR U23694 ( .A(n21420), .B(n21421), .Z(n21048) );
  AND U23695 ( .A(n21422), .B(n21423), .Z(n21420) );
  AND U23696 ( .A(b[9]), .B(a[61]), .Z(n21419) );
  XOR U23697 ( .A(n21425), .B(n21426), .Z(n21053) );
  AND U23698 ( .A(n21427), .B(n21428), .Z(n21425) );
  AND U23699 ( .A(b[8]), .B(a[62]), .Z(n21424) );
  XOR U23700 ( .A(n21430), .B(n21431), .Z(n21058) );
  AND U23701 ( .A(n21432), .B(n21433), .Z(n21430) );
  AND U23702 ( .A(b[7]), .B(a[63]), .Z(n21429) );
  XOR U23703 ( .A(n21435), .B(n21436), .Z(n21063) );
  AND U23704 ( .A(n21437), .B(n21438), .Z(n21435) );
  AND U23705 ( .A(b[6]), .B(a[64]), .Z(n21434) );
  XOR U23706 ( .A(n21440), .B(n21441), .Z(n21068) );
  AND U23707 ( .A(n21442), .B(n21443), .Z(n21440) );
  AND U23708 ( .A(b[5]), .B(a[65]), .Z(n21439) );
  XOR U23709 ( .A(n21445), .B(n21446), .Z(n21073) );
  AND U23710 ( .A(n21447), .B(n21448), .Z(n21445) );
  AND U23711 ( .A(b[4]), .B(a[66]), .Z(n21444) );
  XOR U23712 ( .A(n21450), .B(n21451), .Z(n21078) );
  AND U23713 ( .A(n21452), .B(n21453), .Z(n21450) );
  AND U23714 ( .A(b[3]), .B(a[67]), .Z(n21449) );
  XOR U23715 ( .A(n21455), .B(n21456), .Z(n21083) );
  OR U23716 ( .A(n21457), .B(n21458), .Z(n21456) );
  AND U23717 ( .A(b[2]), .B(a[68]), .Z(n21454) );
  XNOR U23718 ( .A(n21093), .B(n21459), .Z(n21089) );
  NAND U23719 ( .A(b[1]), .B(a[69]), .Z(n21459) );
  IV U23720 ( .A(n21087), .Z(n21093) );
  ANDN U23721 ( .B(n10344), .A(n10346), .Z(n21087) );
  NAND U23722 ( .A(a[69]), .B(b[0]), .Z(n10346) );
  XOR U23723 ( .A(n21457), .B(n21458), .Z(n10344) );
  XOR U23724 ( .A(n21461), .B(n21452), .Z(n21460) );
  XOR U23725 ( .A(n21447), .B(n21451), .Z(n21462) );
  XOR U23726 ( .A(n21442), .B(n21446), .Z(n21463) );
  XOR U23727 ( .A(n21437), .B(n21441), .Z(n21464) );
  XOR U23728 ( .A(n21432), .B(n21436), .Z(n21465) );
  XOR U23729 ( .A(n21427), .B(n21431), .Z(n21466) );
  XOR U23730 ( .A(n21422), .B(n21426), .Z(n21467) );
  XOR U23731 ( .A(n21417), .B(n21421), .Z(n21468) );
  XOR U23732 ( .A(n21412), .B(n21416), .Z(n21469) );
  XOR U23733 ( .A(n21407), .B(n21411), .Z(n21470) );
  XOR U23734 ( .A(n21402), .B(n21406), .Z(n21471) );
  XOR U23735 ( .A(n21397), .B(n21401), .Z(n21472) );
  XOR U23736 ( .A(n21392), .B(n21396), .Z(n21473) );
  XOR U23737 ( .A(n21387), .B(n21391), .Z(n21474) );
  XOR U23738 ( .A(n21382), .B(n21386), .Z(n21475) );
  XOR U23739 ( .A(n21377), .B(n21381), .Z(n21476) );
  XOR U23740 ( .A(n21372), .B(n21376), .Z(n21477) );
  XOR U23741 ( .A(n21367), .B(n21371), .Z(n21478) );
  XOR U23742 ( .A(n21362), .B(n21366), .Z(n21479) );
  XOR U23743 ( .A(n21357), .B(n21361), .Z(n21480) );
  XOR U23744 ( .A(n21352), .B(n21356), .Z(n21481) );
  XOR U23745 ( .A(n21347), .B(n21351), .Z(n21482) );
  XOR U23746 ( .A(n21342), .B(n21346), .Z(n21483) );
  XOR U23747 ( .A(n21337), .B(n21341), .Z(n21484) );
  XOR U23748 ( .A(n21332), .B(n21336), .Z(n21485) );
  XOR U23749 ( .A(n21327), .B(n21331), .Z(n21486) );
  XOR U23750 ( .A(n21322), .B(n21326), .Z(n21487) );
  XOR U23751 ( .A(n21317), .B(n21321), .Z(n21488) );
  XOR U23752 ( .A(n21312), .B(n21316), .Z(n21489) );
  XOR U23753 ( .A(n21307), .B(n21311), .Z(n21490) );
  XOR U23754 ( .A(n21302), .B(n21306), .Z(n21491) );
  XOR U23755 ( .A(n21292), .B(n21301), .Z(n21492) );
  XOR U23756 ( .A(n21493), .B(n21291), .Z(n21292) );
  AND U23757 ( .A(b[33]), .B(a[36]), .Z(n21493) );
  XNOR U23758 ( .A(n21291), .B(n21297), .Z(n21494) );
  XNOR U23759 ( .A(n21296), .B(n21288), .Z(n21495) );
  XNOR U23760 ( .A(n21287), .B(n21283), .Z(n21496) );
  XNOR U23761 ( .A(n21282), .B(n21278), .Z(n21497) );
  XNOR U23762 ( .A(n21277), .B(n21273), .Z(n21498) );
  XNOR U23763 ( .A(n21272), .B(n21268), .Z(n21499) );
  XNOR U23764 ( .A(n21267), .B(n21263), .Z(n21500) );
  XNOR U23765 ( .A(n21262), .B(n21258), .Z(n21501) );
  XNOR U23766 ( .A(n21257), .B(n21253), .Z(n21502) );
  XNOR U23767 ( .A(n21252), .B(n21248), .Z(n21503) );
  XNOR U23768 ( .A(n21247), .B(n21243), .Z(n21504) );
  XNOR U23769 ( .A(n21242), .B(n21238), .Z(n21505) );
  XNOR U23770 ( .A(n21237), .B(n21233), .Z(n21506) );
  XNOR U23771 ( .A(n21232), .B(n21228), .Z(n21507) );
  XNOR U23772 ( .A(n21227), .B(n21223), .Z(n21508) );
  XNOR U23773 ( .A(n21222), .B(n21218), .Z(n21509) );
  XNOR U23774 ( .A(n21217), .B(n21213), .Z(n21510) );
  XNOR U23775 ( .A(n21212), .B(n21208), .Z(n21511) );
  XNOR U23776 ( .A(n21207), .B(n21203), .Z(n21512) );
  XNOR U23777 ( .A(n21202), .B(n21198), .Z(n21513) );
  XNOR U23778 ( .A(n21197), .B(n21193), .Z(n21514) );
  XNOR U23779 ( .A(n21192), .B(n21188), .Z(n21515) );
  XNOR U23780 ( .A(n21187), .B(n21183), .Z(n21516) );
  XNOR U23781 ( .A(n21182), .B(n21178), .Z(n21517) );
  XNOR U23782 ( .A(n21177), .B(n21173), .Z(n21518) );
  XNOR U23783 ( .A(n21172), .B(n21168), .Z(n21519) );
  XOR U23784 ( .A(n21167), .B(n21164), .Z(n21520) );
  XOR U23785 ( .A(n21521), .B(n21522), .Z(n21164) );
  XOR U23786 ( .A(n21162), .B(n21523), .Z(n21522) );
  XOR U23787 ( .A(n21524), .B(n21525), .Z(n21523) );
  XOR U23788 ( .A(n21526), .B(n21527), .Z(n21525) );
  NAND U23789 ( .A(a[7]), .B(b[62]), .Z(n21527) );
  AND U23790 ( .A(a[6]), .B(b[63]), .Z(n21526) );
  XOR U23791 ( .A(n21528), .B(n21524), .Z(n21521) );
  XOR U23792 ( .A(n21529), .B(n21530), .Z(n21524) );
  ANDN U23793 ( .B(n21531), .A(n21532), .Z(n21529) );
  AND U23794 ( .A(a[8]), .B(b[61]), .Z(n21528) );
  XOR U23795 ( .A(n21533), .B(n21162), .Z(n21163) );
  XOR U23796 ( .A(n21534), .B(n21535), .Z(n21162) );
  AND U23797 ( .A(n21536), .B(n21537), .Z(n21534) );
  AND U23798 ( .A(a[9]), .B(b[60]), .Z(n21533) );
  XOR U23799 ( .A(n21538), .B(n21167), .Z(n21169) );
  XOR U23800 ( .A(n21539), .B(n21540), .Z(n21167) );
  AND U23801 ( .A(n21541), .B(n21542), .Z(n21539) );
  AND U23802 ( .A(a[10]), .B(b[59]), .Z(n21538) );
  XOR U23803 ( .A(n21543), .B(n21172), .Z(n21174) );
  XOR U23804 ( .A(n21544), .B(n21545), .Z(n21172) );
  AND U23805 ( .A(n21546), .B(n21547), .Z(n21544) );
  AND U23806 ( .A(a[11]), .B(b[58]), .Z(n21543) );
  XOR U23807 ( .A(n21548), .B(n21177), .Z(n21179) );
  XOR U23808 ( .A(n21549), .B(n21550), .Z(n21177) );
  AND U23809 ( .A(n21551), .B(n21552), .Z(n21549) );
  AND U23810 ( .A(a[12]), .B(b[57]), .Z(n21548) );
  XOR U23811 ( .A(n21553), .B(n21182), .Z(n21184) );
  XOR U23812 ( .A(n21554), .B(n21555), .Z(n21182) );
  AND U23813 ( .A(n21556), .B(n21557), .Z(n21554) );
  AND U23814 ( .A(a[13]), .B(b[56]), .Z(n21553) );
  XOR U23815 ( .A(n21558), .B(n21187), .Z(n21189) );
  XOR U23816 ( .A(n21559), .B(n21560), .Z(n21187) );
  AND U23817 ( .A(n21561), .B(n21562), .Z(n21559) );
  AND U23818 ( .A(a[14]), .B(b[55]), .Z(n21558) );
  XOR U23819 ( .A(n21563), .B(n21192), .Z(n21194) );
  XOR U23820 ( .A(n21564), .B(n21565), .Z(n21192) );
  AND U23821 ( .A(n21566), .B(n21567), .Z(n21564) );
  AND U23822 ( .A(a[15]), .B(b[54]), .Z(n21563) );
  XOR U23823 ( .A(n21568), .B(n21197), .Z(n21199) );
  XOR U23824 ( .A(n21569), .B(n21570), .Z(n21197) );
  AND U23825 ( .A(n21571), .B(n21572), .Z(n21569) );
  AND U23826 ( .A(a[16]), .B(b[53]), .Z(n21568) );
  XOR U23827 ( .A(n21573), .B(n21202), .Z(n21204) );
  XOR U23828 ( .A(n21574), .B(n21575), .Z(n21202) );
  AND U23829 ( .A(n21576), .B(n21577), .Z(n21574) );
  AND U23830 ( .A(a[17]), .B(b[52]), .Z(n21573) );
  XOR U23831 ( .A(n21578), .B(n21207), .Z(n21209) );
  XOR U23832 ( .A(n21579), .B(n21580), .Z(n21207) );
  AND U23833 ( .A(n21581), .B(n21582), .Z(n21579) );
  AND U23834 ( .A(a[18]), .B(b[51]), .Z(n21578) );
  XOR U23835 ( .A(n21583), .B(n21212), .Z(n21214) );
  XOR U23836 ( .A(n21584), .B(n21585), .Z(n21212) );
  AND U23837 ( .A(n21586), .B(n21587), .Z(n21584) );
  AND U23838 ( .A(a[19]), .B(b[50]), .Z(n21583) );
  XOR U23839 ( .A(n21588), .B(n21217), .Z(n21219) );
  XOR U23840 ( .A(n21589), .B(n21590), .Z(n21217) );
  AND U23841 ( .A(n21591), .B(n21592), .Z(n21589) );
  AND U23842 ( .A(a[20]), .B(b[49]), .Z(n21588) );
  XOR U23843 ( .A(n21593), .B(n21222), .Z(n21224) );
  XOR U23844 ( .A(n21594), .B(n21595), .Z(n21222) );
  AND U23845 ( .A(n21596), .B(n21597), .Z(n21594) );
  AND U23846 ( .A(a[21]), .B(b[48]), .Z(n21593) );
  XOR U23847 ( .A(n21598), .B(n21227), .Z(n21229) );
  XOR U23848 ( .A(n21599), .B(n21600), .Z(n21227) );
  AND U23849 ( .A(n21601), .B(n21602), .Z(n21599) );
  AND U23850 ( .A(a[22]), .B(b[47]), .Z(n21598) );
  XOR U23851 ( .A(n21603), .B(n21232), .Z(n21234) );
  XOR U23852 ( .A(n21604), .B(n21605), .Z(n21232) );
  AND U23853 ( .A(n21606), .B(n21607), .Z(n21604) );
  AND U23854 ( .A(a[23]), .B(b[46]), .Z(n21603) );
  XOR U23855 ( .A(n21608), .B(n21237), .Z(n21239) );
  XOR U23856 ( .A(n21609), .B(n21610), .Z(n21237) );
  AND U23857 ( .A(n21611), .B(n21612), .Z(n21609) );
  AND U23858 ( .A(a[24]), .B(b[45]), .Z(n21608) );
  XOR U23859 ( .A(n21613), .B(n21242), .Z(n21244) );
  XOR U23860 ( .A(n21614), .B(n21615), .Z(n21242) );
  AND U23861 ( .A(n21616), .B(n21617), .Z(n21614) );
  AND U23862 ( .A(a[25]), .B(b[44]), .Z(n21613) );
  XOR U23863 ( .A(n21618), .B(n21247), .Z(n21249) );
  XOR U23864 ( .A(n21619), .B(n21620), .Z(n21247) );
  AND U23865 ( .A(n21621), .B(n21622), .Z(n21619) );
  AND U23866 ( .A(a[26]), .B(b[43]), .Z(n21618) );
  XOR U23867 ( .A(n21623), .B(n21252), .Z(n21254) );
  XOR U23868 ( .A(n21624), .B(n21625), .Z(n21252) );
  AND U23869 ( .A(n21626), .B(n21627), .Z(n21624) );
  AND U23870 ( .A(a[27]), .B(b[42]), .Z(n21623) );
  XOR U23871 ( .A(n21628), .B(n21257), .Z(n21259) );
  XOR U23872 ( .A(n21629), .B(n21630), .Z(n21257) );
  AND U23873 ( .A(n21631), .B(n21632), .Z(n21629) );
  AND U23874 ( .A(a[28]), .B(b[41]), .Z(n21628) );
  XOR U23875 ( .A(n21633), .B(n21262), .Z(n21264) );
  XOR U23876 ( .A(n21634), .B(n21635), .Z(n21262) );
  AND U23877 ( .A(n21636), .B(n21637), .Z(n21634) );
  AND U23878 ( .A(a[29]), .B(b[40]), .Z(n21633) );
  XOR U23879 ( .A(n21638), .B(n21267), .Z(n21269) );
  XOR U23880 ( .A(n21639), .B(n21640), .Z(n21267) );
  AND U23881 ( .A(n21641), .B(n21642), .Z(n21639) );
  AND U23882 ( .A(a[30]), .B(b[39]), .Z(n21638) );
  XOR U23883 ( .A(n21643), .B(n21272), .Z(n21274) );
  XOR U23884 ( .A(n21644), .B(n21645), .Z(n21272) );
  AND U23885 ( .A(n21646), .B(n21647), .Z(n21644) );
  AND U23886 ( .A(a[31]), .B(b[38]), .Z(n21643) );
  XOR U23887 ( .A(n21648), .B(n21277), .Z(n21279) );
  XOR U23888 ( .A(n21649), .B(n21650), .Z(n21277) );
  AND U23889 ( .A(n21651), .B(n21652), .Z(n21649) );
  AND U23890 ( .A(a[32]), .B(b[37]), .Z(n21648) );
  XOR U23891 ( .A(n21653), .B(n21282), .Z(n21284) );
  XOR U23892 ( .A(n21654), .B(n21655), .Z(n21282) );
  AND U23893 ( .A(n21656), .B(n21657), .Z(n21654) );
  AND U23894 ( .A(a[33]), .B(b[36]), .Z(n21653) );
  XOR U23895 ( .A(n21658), .B(n21287), .Z(n21289) );
  XOR U23896 ( .A(n21659), .B(n21660), .Z(n21287) );
  AND U23897 ( .A(n21661), .B(n21662), .Z(n21659) );
  AND U23898 ( .A(a[34]), .B(b[35]), .Z(n21658) );
  XOR U23899 ( .A(n21663), .B(n21664), .Z(n21291) );
  AND U23900 ( .A(n21665), .B(n21666), .Z(n21663) );
  XOR U23901 ( .A(n21667), .B(n21296), .Z(n21298) );
  XOR U23902 ( .A(n21668), .B(n21669), .Z(n21296) );
  AND U23903 ( .A(n21670), .B(n21671), .Z(n21668) );
  AND U23904 ( .A(b[34]), .B(a[35]), .Z(n21667) );
  XOR U23905 ( .A(n21673), .B(n21674), .Z(n21301) );
  AND U23906 ( .A(n21675), .B(n21676), .Z(n21673) );
  AND U23907 ( .A(b[32]), .B(a[37]), .Z(n21672) );
  XOR U23908 ( .A(n21678), .B(n21679), .Z(n21306) );
  AND U23909 ( .A(n21680), .B(n21681), .Z(n21678) );
  AND U23910 ( .A(b[31]), .B(a[38]), .Z(n21677) );
  XOR U23911 ( .A(n21683), .B(n21684), .Z(n21311) );
  AND U23912 ( .A(n21685), .B(n21686), .Z(n21683) );
  AND U23913 ( .A(b[30]), .B(a[39]), .Z(n21682) );
  XOR U23914 ( .A(n21688), .B(n21689), .Z(n21316) );
  AND U23915 ( .A(n21690), .B(n21691), .Z(n21688) );
  AND U23916 ( .A(b[29]), .B(a[40]), .Z(n21687) );
  XOR U23917 ( .A(n21693), .B(n21694), .Z(n21321) );
  AND U23918 ( .A(n21695), .B(n21696), .Z(n21693) );
  AND U23919 ( .A(b[28]), .B(a[41]), .Z(n21692) );
  XOR U23920 ( .A(n21698), .B(n21699), .Z(n21326) );
  AND U23921 ( .A(n21700), .B(n21701), .Z(n21698) );
  AND U23922 ( .A(b[27]), .B(a[42]), .Z(n21697) );
  XOR U23923 ( .A(n21703), .B(n21704), .Z(n21331) );
  AND U23924 ( .A(n21705), .B(n21706), .Z(n21703) );
  AND U23925 ( .A(b[26]), .B(a[43]), .Z(n21702) );
  XOR U23926 ( .A(n21708), .B(n21709), .Z(n21336) );
  AND U23927 ( .A(n21710), .B(n21711), .Z(n21708) );
  AND U23928 ( .A(b[25]), .B(a[44]), .Z(n21707) );
  XOR U23929 ( .A(n21713), .B(n21714), .Z(n21341) );
  AND U23930 ( .A(n21715), .B(n21716), .Z(n21713) );
  AND U23931 ( .A(b[24]), .B(a[45]), .Z(n21712) );
  XOR U23932 ( .A(n21718), .B(n21719), .Z(n21346) );
  AND U23933 ( .A(n21720), .B(n21721), .Z(n21718) );
  AND U23934 ( .A(b[23]), .B(a[46]), .Z(n21717) );
  XOR U23935 ( .A(n21723), .B(n21724), .Z(n21351) );
  AND U23936 ( .A(n21725), .B(n21726), .Z(n21723) );
  AND U23937 ( .A(b[22]), .B(a[47]), .Z(n21722) );
  XOR U23938 ( .A(n21728), .B(n21729), .Z(n21356) );
  AND U23939 ( .A(n21730), .B(n21731), .Z(n21728) );
  AND U23940 ( .A(b[21]), .B(a[48]), .Z(n21727) );
  XOR U23941 ( .A(n21733), .B(n21734), .Z(n21361) );
  AND U23942 ( .A(n21735), .B(n21736), .Z(n21733) );
  AND U23943 ( .A(b[20]), .B(a[49]), .Z(n21732) );
  XOR U23944 ( .A(n21738), .B(n21739), .Z(n21366) );
  AND U23945 ( .A(n21740), .B(n21741), .Z(n21738) );
  AND U23946 ( .A(b[19]), .B(a[50]), .Z(n21737) );
  XOR U23947 ( .A(n21743), .B(n21744), .Z(n21371) );
  AND U23948 ( .A(n21745), .B(n21746), .Z(n21743) );
  AND U23949 ( .A(b[18]), .B(a[51]), .Z(n21742) );
  XOR U23950 ( .A(n21748), .B(n21749), .Z(n21376) );
  AND U23951 ( .A(n21750), .B(n21751), .Z(n21748) );
  AND U23952 ( .A(b[17]), .B(a[52]), .Z(n21747) );
  XOR U23953 ( .A(n21753), .B(n21754), .Z(n21381) );
  AND U23954 ( .A(n21755), .B(n21756), .Z(n21753) );
  AND U23955 ( .A(b[16]), .B(a[53]), .Z(n21752) );
  XOR U23956 ( .A(n21758), .B(n21759), .Z(n21386) );
  AND U23957 ( .A(n21760), .B(n21761), .Z(n21758) );
  AND U23958 ( .A(b[15]), .B(a[54]), .Z(n21757) );
  XOR U23959 ( .A(n21763), .B(n21764), .Z(n21391) );
  AND U23960 ( .A(n21765), .B(n21766), .Z(n21763) );
  AND U23961 ( .A(b[14]), .B(a[55]), .Z(n21762) );
  XOR U23962 ( .A(n21768), .B(n21769), .Z(n21396) );
  AND U23963 ( .A(n21770), .B(n21771), .Z(n21768) );
  AND U23964 ( .A(b[13]), .B(a[56]), .Z(n21767) );
  XOR U23965 ( .A(n21773), .B(n21774), .Z(n21401) );
  AND U23966 ( .A(n21775), .B(n21776), .Z(n21773) );
  AND U23967 ( .A(b[12]), .B(a[57]), .Z(n21772) );
  XOR U23968 ( .A(n21778), .B(n21779), .Z(n21406) );
  AND U23969 ( .A(n21780), .B(n21781), .Z(n21778) );
  AND U23970 ( .A(b[11]), .B(a[58]), .Z(n21777) );
  XOR U23971 ( .A(n21783), .B(n21784), .Z(n21411) );
  AND U23972 ( .A(n21785), .B(n21786), .Z(n21783) );
  AND U23973 ( .A(b[10]), .B(a[59]), .Z(n21782) );
  XOR U23974 ( .A(n21788), .B(n21789), .Z(n21416) );
  AND U23975 ( .A(n21790), .B(n21791), .Z(n21788) );
  AND U23976 ( .A(b[9]), .B(a[60]), .Z(n21787) );
  XOR U23977 ( .A(n21793), .B(n21794), .Z(n21421) );
  AND U23978 ( .A(n21795), .B(n21796), .Z(n21793) );
  AND U23979 ( .A(b[8]), .B(a[61]), .Z(n21792) );
  XOR U23980 ( .A(n21798), .B(n21799), .Z(n21426) );
  AND U23981 ( .A(n21800), .B(n21801), .Z(n21798) );
  AND U23982 ( .A(b[7]), .B(a[62]), .Z(n21797) );
  XOR U23983 ( .A(n21803), .B(n21804), .Z(n21431) );
  AND U23984 ( .A(n21805), .B(n21806), .Z(n21803) );
  AND U23985 ( .A(b[6]), .B(a[63]), .Z(n21802) );
  XOR U23986 ( .A(n21808), .B(n21809), .Z(n21436) );
  AND U23987 ( .A(n21810), .B(n21811), .Z(n21808) );
  AND U23988 ( .A(b[5]), .B(a[64]), .Z(n21807) );
  XOR U23989 ( .A(n21813), .B(n21814), .Z(n21441) );
  AND U23990 ( .A(n21815), .B(n21816), .Z(n21813) );
  AND U23991 ( .A(b[4]), .B(a[65]), .Z(n21812) );
  XOR U23992 ( .A(n21818), .B(n21819), .Z(n21446) );
  AND U23993 ( .A(n21820), .B(n21821), .Z(n21818) );
  AND U23994 ( .A(b[3]), .B(a[66]), .Z(n21817) );
  XOR U23995 ( .A(n21823), .B(n21824), .Z(n21451) );
  OR U23996 ( .A(n21825), .B(n21826), .Z(n21824) );
  AND U23997 ( .A(b[2]), .B(a[67]), .Z(n21822) );
  XNOR U23998 ( .A(n21461), .B(n21827), .Z(n21457) );
  NAND U23999 ( .A(b[1]), .B(a[68]), .Z(n21827) );
  IV U24000 ( .A(n21455), .Z(n21461) );
  ANDN U24001 ( .B(n10347), .A(n10349), .Z(n21455) );
  NAND U24002 ( .A(a[68]), .B(b[0]), .Z(n10349) );
  XOR U24003 ( .A(n21825), .B(n21826), .Z(n10347) );
  XOR U24004 ( .A(n21829), .B(n21820), .Z(n21828) );
  XOR U24005 ( .A(n21815), .B(n21819), .Z(n21830) );
  XOR U24006 ( .A(n21810), .B(n21814), .Z(n21831) );
  XOR U24007 ( .A(n21805), .B(n21809), .Z(n21832) );
  XOR U24008 ( .A(n21800), .B(n21804), .Z(n21833) );
  XOR U24009 ( .A(n21795), .B(n21799), .Z(n21834) );
  XOR U24010 ( .A(n21790), .B(n21794), .Z(n21835) );
  XOR U24011 ( .A(n21785), .B(n21789), .Z(n21836) );
  XOR U24012 ( .A(n21780), .B(n21784), .Z(n21837) );
  XOR U24013 ( .A(n21775), .B(n21779), .Z(n21838) );
  XOR U24014 ( .A(n21770), .B(n21774), .Z(n21839) );
  XOR U24015 ( .A(n21765), .B(n21769), .Z(n21840) );
  XOR U24016 ( .A(n21760), .B(n21764), .Z(n21841) );
  XOR U24017 ( .A(n21755), .B(n21759), .Z(n21842) );
  XOR U24018 ( .A(n21750), .B(n21754), .Z(n21843) );
  XOR U24019 ( .A(n21745), .B(n21749), .Z(n21844) );
  XOR U24020 ( .A(n21740), .B(n21744), .Z(n21845) );
  XOR U24021 ( .A(n21735), .B(n21739), .Z(n21846) );
  XOR U24022 ( .A(n21730), .B(n21734), .Z(n21847) );
  XOR U24023 ( .A(n21725), .B(n21729), .Z(n21848) );
  XOR U24024 ( .A(n21720), .B(n21724), .Z(n21849) );
  XOR U24025 ( .A(n21715), .B(n21719), .Z(n21850) );
  XOR U24026 ( .A(n21710), .B(n21714), .Z(n21851) );
  XOR U24027 ( .A(n21705), .B(n21709), .Z(n21852) );
  XOR U24028 ( .A(n21700), .B(n21704), .Z(n21853) );
  XOR U24029 ( .A(n21695), .B(n21699), .Z(n21854) );
  XOR U24030 ( .A(n21690), .B(n21694), .Z(n21855) );
  XOR U24031 ( .A(n21685), .B(n21689), .Z(n21856) );
  XOR U24032 ( .A(n21680), .B(n21684), .Z(n21857) );
  XOR U24033 ( .A(n21675), .B(n21679), .Z(n21858) );
  XOR U24034 ( .A(n21665), .B(n21674), .Z(n21859) );
  XOR U24035 ( .A(n21860), .B(n21664), .Z(n21665) );
  AND U24036 ( .A(b[32]), .B(a[36]), .Z(n21860) );
  XNOR U24037 ( .A(n21664), .B(n21670), .Z(n21861) );
  XNOR U24038 ( .A(n21669), .B(n21661), .Z(n21862) );
  XNOR U24039 ( .A(n21660), .B(n21656), .Z(n21863) );
  XNOR U24040 ( .A(n21655), .B(n21651), .Z(n21864) );
  XNOR U24041 ( .A(n21650), .B(n21646), .Z(n21865) );
  XNOR U24042 ( .A(n21645), .B(n21641), .Z(n21866) );
  XNOR U24043 ( .A(n21640), .B(n21636), .Z(n21867) );
  XNOR U24044 ( .A(n21635), .B(n21631), .Z(n21868) );
  XNOR U24045 ( .A(n21630), .B(n21626), .Z(n21869) );
  XNOR U24046 ( .A(n21625), .B(n21621), .Z(n21870) );
  XNOR U24047 ( .A(n21620), .B(n21616), .Z(n21871) );
  XNOR U24048 ( .A(n21615), .B(n21611), .Z(n21872) );
  XNOR U24049 ( .A(n21610), .B(n21606), .Z(n21873) );
  XNOR U24050 ( .A(n21605), .B(n21601), .Z(n21874) );
  XNOR U24051 ( .A(n21600), .B(n21596), .Z(n21875) );
  XNOR U24052 ( .A(n21595), .B(n21591), .Z(n21876) );
  XNOR U24053 ( .A(n21590), .B(n21586), .Z(n21877) );
  XNOR U24054 ( .A(n21585), .B(n21581), .Z(n21878) );
  XNOR U24055 ( .A(n21580), .B(n21576), .Z(n21879) );
  XNOR U24056 ( .A(n21575), .B(n21571), .Z(n21880) );
  XNOR U24057 ( .A(n21570), .B(n21566), .Z(n21881) );
  XNOR U24058 ( .A(n21565), .B(n21561), .Z(n21882) );
  XNOR U24059 ( .A(n21560), .B(n21556), .Z(n21883) );
  XNOR U24060 ( .A(n21555), .B(n21551), .Z(n21884) );
  XNOR U24061 ( .A(n21550), .B(n21546), .Z(n21885) );
  XNOR U24062 ( .A(n21545), .B(n21541), .Z(n21886) );
  XNOR U24063 ( .A(n21540), .B(n21536), .Z(n21887) );
  XOR U24064 ( .A(n21535), .B(n21532), .Z(n21888) );
  XOR U24065 ( .A(n21889), .B(n21890), .Z(n21532) );
  XOR U24066 ( .A(n21530), .B(n21891), .Z(n21890) );
  XOR U24067 ( .A(n21892), .B(n21893), .Z(n21891) );
  XOR U24068 ( .A(n21894), .B(n21895), .Z(n21893) );
  NAND U24069 ( .A(a[6]), .B(b[62]), .Z(n21895) );
  AND U24070 ( .A(a[5]), .B(b[63]), .Z(n21894) );
  XOR U24071 ( .A(n21896), .B(n21892), .Z(n21889) );
  XOR U24072 ( .A(n21897), .B(n21898), .Z(n21892) );
  ANDN U24073 ( .B(n21899), .A(n21900), .Z(n21897) );
  AND U24074 ( .A(a[7]), .B(b[61]), .Z(n21896) );
  XOR U24075 ( .A(n21901), .B(n21530), .Z(n21531) );
  XOR U24076 ( .A(n21902), .B(n21903), .Z(n21530) );
  AND U24077 ( .A(n21904), .B(n21905), .Z(n21902) );
  AND U24078 ( .A(a[8]), .B(b[60]), .Z(n21901) );
  XOR U24079 ( .A(n21906), .B(n21535), .Z(n21537) );
  XOR U24080 ( .A(n21907), .B(n21908), .Z(n21535) );
  AND U24081 ( .A(n21909), .B(n21910), .Z(n21907) );
  AND U24082 ( .A(a[9]), .B(b[59]), .Z(n21906) );
  XOR U24083 ( .A(n21911), .B(n21540), .Z(n21542) );
  XOR U24084 ( .A(n21912), .B(n21913), .Z(n21540) );
  AND U24085 ( .A(n21914), .B(n21915), .Z(n21912) );
  AND U24086 ( .A(a[10]), .B(b[58]), .Z(n21911) );
  XOR U24087 ( .A(n21916), .B(n21545), .Z(n21547) );
  XOR U24088 ( .A(n21917), .B(n21918), .Z(n21545) );
  AND U24089 ( .A(n21919), .B(n21920), .Z(n21917) );
  AND U24090 ( .A(a[11]), .B(b[57]), .Z(n21916) );
  XOR U24091 ( .A(n21921), .B(n21550), .Z(n21552) );
  XOR U24092 ( .A(n21922), .B(n21923), .Z(n21550) );
  AND U24093 ( .A(n21924), .B(n21925), .Z(n21922) );
  AND U24094 ( .A(a[12]), .B(b[56]), .Z(n21921) );
  XOR U24095 ( .A(n21926), .B(n21555), .Z(n21557) );
  XOR U24096 ( .A(n21927), .B(n21928), .Z(n21555) );
  AND U24097 ( .A(n21929), .B(n21930), .Z(n21927) );
  AND U24098 ( .A(a[13]), .B(b[55]), .Z(n21926) );
  XOR U24099 ( .A(n21931), .B(n21560), .Z(n21562) );
  XOR U24100 ( .A(n21932), .B(n21933), .Z(n21560) );
  AND U24101 ( .A(n21934), .B(n21935), .Z(n21932) );
  AND U24102 ( .A(a[14]), .B(b[54]), .Z(n21931) );
  XOR U24103 ( .A(n21936), .B(n21565), .Z(n21567) );
  XOR U24104 ( .A(n21937), .B(n21938), .Z(n21565) );
  AND U24105 ( .A(n21939), .B(n21940), .Z(n21937) );
  AND U24106 ( .A(a[15]), .B(b[53]), .Z(n21936) );
  XOR U24107 ( .A(n21941), .B(n21570), .Z(n21572) );
  XOR U24108 ( .A(n21942), .B(n21943), .Z(n21570) );
  AND U24109 ( .A(n21944), .B(n21945), .Z(n21942) );
  AND U24110 ( .A(a[16]), .B(b[52]), .Z(n21941) );
  XOR U24111 ( .A(n21946), .B(n21575), .Z(n21577) );
  XOR U24112 ( .A(n21947), .B(n21948), .Z(n21575) );
  AND U24113 ( .A(n21949), .B(n21950), .Z(n21947) );
  AND U24114 ( .A(a[17]), .B(b[51]), .Z(n21946) );
  XOR U24115 ( .A(n21951), .B(n21580), .Z(n21582) );
  XOR U24116 ( .A(n21952), .B(n21953), .Z(n21580) );
  AND U24117 ( .A(n21954), .B(n21955), .Z(n21952) );
  AND U24118 ( .A(a[18]), .B(b[50]), .Z(n21951) );
  XOR U24119 ( .A(n21956), .B(n21585), .Z(n21587) );
  XOR U24120 ( .A(n21957), .B(n21958), .Z(n21585) );
  AND U24121 ( .A(n21959), .B(n21960), .Z(n21957) );
  AND U24122 ( .A(a[19]), .B(b[49]), .Z(n21956) );
  XOR U24123 ( .A(n21961), .B(n21590), .Z(n21592) );
  XOR U24124 ( .A(n21962), .B(n21963), .Z(n21590) );
  AND U24125 ( .A(n21964), .B(n21965), .Z(n21962) );
  AND U24126 ( .A(a[20]), .B(b[48]), .Z(n21961) );
  XOR U24127 ( .A(n21966), .B(n21595), .Z(n21597) );
  XOR U24128 ( .A(n21967), .B(n21968), .Z(n21595) );
  AND U24129 ( .A(n21969), .B(n21970), .Z(n21967) );
  AND U24130 ( .A(a[21]), .B(b[47]), .Z(n21966) );
  XOR U24131 ( .A(n21971), .B(n21600), .Z(n21602) );
  XOR U24132 ( .A(n21972), .B(n21973), .Z(n21600) );
  AND U24133 ( .A(n21974), .B(n21975), .Z(n21972) );
  AND U24134 ( .A(a[22]), .B(b[46]), .Z(n21971) );
  XOR U24135 ( .A(n21976), .B(n21605), .Z(n21607) );
  XOR U24136 ( .A(n21977), .B(n21978), .Z(n21605) );
  AND U24137 ( .A(n21979), .B(n21980), .Z(n21977) );
  AND U24138 ( .A(a[23]), .B(b[45]), .Z(n21976) );
  XOR U24139 ( .A(n21981), .B(n21610), .Z(n21612) );
  XOR U24140 ( .A(n21982), .B(n21983), .Z(n21610) );
  AND U24141 ( .A(n21984), .B(n21985), .Z(n21982) );
  AND U24142 ( .A(a[24]), .B(b[44]), .Z(n21981) );
  XOR U24143 ( .A(n21986), .B(n21615), .Z(n21617) );
  XOR U24144 ( .A(n21987), .B(n21988), .Z(n21615) );
  AND U24145 ( .A(n21989), .B(n21990), .Z(n21987) );
  AND U24146 ( .A(a[25]), .B(b[43]), .Z(n21986) );
  XOR U24147 ( .A(n21991), .B(n21620), .Z(n21622) );
  XOR U24148 ( .A(n21992), .B(n21993), .Z(n21620) );
  AND U24149 ( .A(n21994), .B(n21995), .Z(n21992) );
  AND U24150 ( .A(a[26]), .B(b[42]), .Z(n21991) );
  XOR U24151 ( .A(n21996), .B(n21625), .Z(n21627) );
  XOR U24152 ( .A(n21997), .B(n21998), .Z(n21625) );
  AND U24153 ( .A(n21999), .B(n22000), .Z(n21997) );
  AND U24154 ( .A(a[27]), .B(b[41]), .Z(n21996) );
  XOR U24155 ( .A(n22001), .B(n21630), .Z(n21632) );
  XOR U24156 ( .A(n22002), .B(n22003), .Z(n21630) );
  AND U24157 ( .A(n22004), .B(n22005), .Z(n22002) );
  AND U24158 ( .A(a[28]), .B(b[40]), .Z(n22001) );
  XOR U24159 ( .A(n22006), .B(n21635), .Z(n21637) );
  XOR U24160 ( .A(n22007), .B(n22008), .Z(n21635) );
  AND U24161 ( .A(n22009), .B(n22010), .Z(n22007) );
  AND U24162 ( .A(a[29]), .B(b[39]), .Z(n22006) );
  XOR U24163 ( .A(n22011), .B(n21640), .Z(n21642) );
  XOR U24164 ( .A(n22012), .B(n22013), .Z(n21640) );
  AND U24165 ( .A(n22014), .B(n22015), .Z(n22012) );
  AND U24166 ( .A(a[30]), .B(b[38]), .Z(n22011) );
  XOR U24167 ( .A(n22016), .B(n21645), .Z(n21647) );
  XOR U24168 ( .A(n22017), .B(n22018), .Z(n21645) );
  AND U24169 ( .A(n22019), .B(n22020), .Z(n22017) );
  AND U24170 ( .A(a[31]), .B(b[37]), .Z(n22016) );
  XOR U24171 ( .A(n22021), .B(n21650), .Z(n21652) );
  XOR U24172 ( .A(n22022), .B(n22023), .Z(n21650) );
  AND U24173 ( .A(n22024), .B(n22025), .Z(n22022) );
  AND U24174 ( .A(a[32]), .B(b[36]), .Z(n22021) );
  XOR U24175 ( .A(n22026), .B(n21655), .Z(n21657) );
  XOR U24176 ( .A(n22027), .B(n22028), .Z(n21655) );
  AND U24177 ( .A(n22029), .B(n22030), .Z(n22027) );
  AND U24178 ( .A(a[33]), .B(b[35]), .Z(n22026) );
  XOR U24179 ( .A(n22031), .B(n21660), .Z(n21662) );
  XOR U24180 ( .A(n22032), .B(n22033), .Z(n21660) );
  AND U24181 ( .A(n22034), .B(n22035), .Z(n22032) );
  AND U24182 ( .A(a[34]), .B(b[34]), .Z(n22031) );
  XOR U24183 ( .A(n22036), .B(n22037), .Z(n21664) );
  AND U24184 ( .A(n22038), .B(n22039), .Z(n22036) );
  XOR U24185 ( .A(n22040), .B(n21669), .Z(n21671) );
  XOR U24186 ( .A(n22041), .B(n22042), .Z(n21669) );
  AND U24187 ( .A(n22043), .B(n22044), .Z(n22041) );
  AND U24188 ( .A(b[33]), .B(a[35]), .Z(n22040) );
  XOR U24189 ( .A(n22046), .B(n22047), .Z(n21674) );
  AND U24190 ( .A(n22048), .B(n22049), .Z(n22046) );
  AND U24191 ( .A(b[31]), .B(a[37]), .Z(n22045) );
  XOR U24192 ( .A(n22051), .B(n22052), .Z(n21679) );
  AND U24193 ( .A(n22053), .B(n22054), .Z(n22051) );
  AND U24194 ( .A(b[30]), .B(a[38]), .Z(n22050) );
  XOR U24195 ( .A(n22056), .B(n22057), .Z(n21684) );
  AND U24196 ( .A(n22058), .B(n22059), .Z(n22056) );
  AND U24197 ( .A(b[29]), .B(a[39]), .Z(n22055) );
  XOR U24198 ( .A(n22061), .B(n22062), .Z(n21689) );
  AND U24199 ( .A(n22063), .B(n22064), .Z(n22061) );
  AND U24200 ( .A(b[28]), .B(a[40]), .Z(n22060) );
  XOR U24201 ( .A(n22066), .B(n22067), .Z(n21694) );
  AND U24202 ( .A(n22068), .B(n22069), .Z(n22066) );
  AND U24203 ( .A(b[27]), .B(a[41]), .Z(n22065) );
  XOR U24204 ( .A(n22071), .B(n22072), .Z(n21699) );
  AND U24205 ( .A(n22073), .B(n22074), .Z(n22071) );
  AND U24206 ( .A(b[26]), .B(a[42]), .Z(n22070) );
  XOR U24207 ( .A(n22076), .B(n22077), .Z(n21704) );
  AND U24208 ( .A(n22078), .B(n22079), .Z(n22076) );
  AND U24209 ( .A(b[25]), .B(a[43]), .Z(n22075) );
  XOR U24210 ( .A(n22081), .B(n22082), .Z(n21709) );
  AND U24211 ( .A(n22083), .B(n22084), .Z(n22081) );
  AND U24212 ( .A(b[24]), .B(a[44]), .Z(n22080) );
  XOR U24213 ( .A(n22086), .B(n22087), .Z(n21714) );
  AND U24214 ( .A(n22088), .B(n22089), .Z(n22086) );
  AND U24215 ( .A(b[23]), .B(a[45]), .Z(n22085) );
  XOR U24216 ( .A(n22091), .B(n22092), .Z(n21719) );
  AND U24217 ( .A(n22093), .B(n22094), .Z(n22091) );
  AND U24218 ( .A(b[22]), .B(a[46]), .Z(n22090) );
  XOR U24219 ( .A(n22096), .B(n22097), .Z(n21724) );
  AND U24220 ( .A(n22098), .B(n22099), .Z(n22096) );
  AND U24221 ( .A(b[21]), .B(a[47]), .Z(n22095) );
  XOR U24222 ( .A(n22101), .B(n22102), .Z(n21729) );
  AND U24223 ( .A(n22103), .B(n22104), .Z(n22101) );
  AND U24224 ( .A(b[20]), .B(a[48]), .Z(n22100) );
  XOR U24225 ( .A(n22106), .B(n22107), .Z(n21734) );
  AND U24226 ( .A(n22108), .B(n22109), .Z(n22106) );
  AND U24227 ( .A(b[19]), .B(a[49]), .Z(n22105) );
  XOR U24228 ( .A(n22111), .B(n22112), .Z(n21739) );
  AND U24229 ( .A(n22113), .B(n22114), .Z(n22111) );
  AND U24230 ( .A(b[18]), .B(a[50]), .Z(n22110) );
  XOR U24231 ( .A(n22116), .B(n22117), .Z(n21744) );
  AND U24232 ( .A(n22118), .B(n22119), .Z(n22116) );
  AND U24233 ( .A(b[17]), .B(a[51]), .Z(n22115) );
  XOR U24234 ( .A(n22121), .B(n22122), .Z(n21749) );
  AND U24235 ( .A(n22123), .B(n22124), .Z(n22121) );
  AND U24236 ( .A(b[16]), .B(a[52]), .Z(n22120) );
  XOR U24237 ( .A(n22126), .B(n22127), .Z(n21754) );
  AND U24238 ( .A(n22128), .B(n22129), .Z(n22126) );
  AND U24239 ( .A(b[15]), .B(a[53]), .Z(n22125) );
  XOR U24240 ( .A(n22131), .B(n22132), .Z(n21759) );
  AND U24241 ( .A(n22133), .B(n22134), .Z(n22131) );
  AND U24242 ( .A(b[14]), .B(a[54]), .Z(n22130) );
  XOR U24243 ( .A(n22136), .B(n22137), .Z(n21764) );
  AND U24244 ( .A(n22138), .B(n22139), .Z(n22136) );
  AND U24245 ( .A(b[13]), .B(a[55]), .Z(n22135) );
  XOR U24246 ( .A(n22141), .B(n22142), .Z(n21769) );
  AND U24247 ( .A(n22143), .B(n22144), .Z(n22141) );
  AND U24248 ( .A(b[12]), .B(a[56]), .Z(n22140) );
  XOR U24249 ( .A(n22146), .B(n22147), .Z(n21774) );
  AND U24250 ( .A(n22148), .B(n22149), .Z(n22146) );
  AND U24251 ( .A(b[11]), .B(a[57]), .Z(n22145) );
  XOR U24252 ( .A(n22151), .B(n22152), .Z(n21779) );
  AND U24253 ( .A(n22153), .B(n22154), .Z(n22151) );
  AND U24254 ( .A(b[10]), .B(a[58]), .Z(n22150) );
  XOR U24255 ( .A(n22156), .B(n22157), .Z(n21784) );
  AND U24256 ( .A(n22158), .B(n22159), .Z(n22156) );
  AND U24257 ( .A(b[9]), .B(a[59]), .Z(n22155) );
  XOR U24258 ( .A(n22161), .B(n22162), .Z(n21789) );
  AND U24259 ( .A(n22163), .B(n22164), .Z(n22161) );
  AND U24260 ( .A(b[8]), .B(a[60]), .Z(n22160) );
  XOR U24261 ( .A(n22166), .B(n22167), .Z(n21794) );
  AND U24262 ( .A(n22168), .B(n22169), .Z(n22166) );
  AND U24263 ( .A(b[7]), .B(a[61]), .Z(n22165) );
  XOR U24264 ( .A(n22171), .B(n22172), .Z(n21799) );
  AND U24265 ( .A(n22173), .B(n22174), .Z(n22171) );
  AND U24266 ( .A(b[6]), .B(a[62]), .Z(n22170) );
  XOR U24267 ( .A(n22176), .B(n22177), .Z(n21804) );
  AND U24268 ( .A(n22178), .B(n22179), .Z(n22176) );
  AND U24269 ( .A(b[5]), .B(a[63]), .Z(n22175) );
  XOR U24270 ( .A(n22181), .B(n22182), .Z(n21809) );
  AND U24271 ( .A(n22183), .B(n22184), .Z(n22181) );
  AND U24272 ( .A(b[4]), .B(a[64]), .Z(n22180) );
  XOR U24273 ( .A(n22186), .B(n22187), .Z(n21814) );
  AND U24274 ( .A(n22188), .B(n22189), .Z(n22186) );
  AND U24275 ( .A(b[3]), .B(a[65]), .Z(n22185) );
  XOR U24276 ( .A(n22191), .B(n22192), .Z(n21819) );
  OR U24277 ( .A(n22193), .B(n22194), .Z(n22192) );
  AND U24278 ( .A(b[2]), .B(a[66]), .Z(n22190) );
  XNOR U24279 ( .A(n21829), .B(n22195), .Z(n21825) );
  NAND U24280 ( .A(b[1]), .B(a[67]), .Z(n22195) );
  IV U24281 ( .A(n21823), .Z(n21829) );
  ANDN U24282 ( .B(n10350), .A(n10352), .Z(n21823) );
  NAND U24283 ( .A(a[67]), .B(b[0]), .Z(n10352) );
  XOR U24284 ( .A(n22193), .B(n22194), .Z(n10350) );
  XOR U24285 ( .A(n22197), .B(n22188), .Z(n22196) );
  XOR U24286 ( .A(n22183), .B(n22187), .Z(n22198) );
  XOR U24287 ( .A(n22178), .B(n22182), .Z(n22199) );
  XOR U24288 ( .A(n22173), .B(n22177), .Z(n22200) );
  XOR U24289 ( .A(n22168), .B(n22172), .Z(n22201) );
  XOR U24290 ( .A(n22163), .B(n22167), .Z(n22202) );
  XOR U24291 ( .A(n22158), .B(n22162), .Z(n22203) );
  XOR U24292 ( .A(n22153), .B(n22157), .Z(n22204) );
  XOR U24293 ( .A(n22148), .B(n22152), .Z(n22205) );
  XOR U24294 ( .A(n22143), .B(n22147), .Z(n22206) );
  XOR U24295 ( .A(n22138), .B(n22142), .Z(n22207) );
  XOR U24296 ( .A(n22133), .B(n22137), .Z(n22208) );
  XOR U24297 ( .A(n22128), .B(n22132), .Z(n22209) );
  XOR U24298 ( .A(n22123), .B(n22127), .Z(n22210) );
  XOR U24299 ( .A(n22118), .B(n22122), .Z(n22211) );
  XOR U24300 ( .A(n22113), .B(n22117), .Z(n22212) );
  XOR U24301 ( .A(n22108), .B(n22112), .Z(n22213) );
  XOR U24302 ( .A(n22103), .B(n22107), .Z(n22214) );
  XOR U24303 ( .A(n22098), .B(n22102), .Z(n22215) );
  XOR U24304 ( .A(n22093), .B(n22097), .Z(n22216) );
  XOR U24305 ( .A(n22088), .B(n22092), .Z(n22217) );
  XOR U24306 ( .A(n22083), .B(n22087), .Z(n22218) );
  XOR U24307 ( .A(n22078), .B(n22082), .Z(n22219) );
  XOR U24308 ( .A(n22073), .B(n22077), .Z(n22220) );
  XOR U24309 ( .A(n22068), .B(n22072), .Z(n22221) );
  XOR U24310 ( .A(n22063), .B(n22067), .Z(n22222) );
  XOR U24311 ( .A(n22058), .B(n22062), .Z(n22223) );
  XOR U24312 ( .A(n22053), .B(n22057), .Z(n22224) );
  XOR U24313 ( .A(n22048), .B(n22052), .Z(n22225) );
  XOR U24314 ( .A(n22038), .B(n22047), .Z(n22226) );
  XOR U24315 ( .A(n22227), .B(n22037), .Z(n22038) );
  AND U24316 ( .A(b[31]), .B(a[36]), .Z(n22227) );
  XNOR U24317 ( .A(n22037), .B(n22043), .Z(n22228) );
  XNOR U24318 ( .A(n22042), .B(n22034), .Z(n22229) );
  XNOR U24319 ( .A(n22033), .B(n22029), .Z(n22230) );
  XNOR U24320 ( .A(n22028), .B(n22024), .Z(n22231) );
  XNOR U24321 ( .A(n22023), .B(n22019), .Z(n22232) );
  XNOR U24322 ( .A(n22018), .B(n22014), .Z(n22233) );
  XNOR U24323 ( .A(n22013), .B(n22009), .Z(n22234) );
  XNOR U24324 ( .A(n22008), .B(n22004), .Z(n22235) );
  XNOR U24325 ( .A(n22003), .B(n21999), .Z(n22236) );
  XNOR U24326 ( .A(n21998), .B(n21994), .Z(n22237) );
  XNOR U24327 ( .A(n21993), .B(n21989), .Z(n22238) );
  XNOR U24328 ( .A(n21988), .B(n21984), .Z(n22239) );
  XNOR U24329 ( .A(n21983), .B(n21979), .Z(n22240) );
  XNOR U24330 ( .A(n21978), .B(n21974), .Z(n22241) );
  XNOR U24331 ( .A(n21973), .B(n21969), .Z(n22242) );
  XNOR U24332 ( .A(n21968), .B(n21964), .Z(n22243) );
  XNOR U24333 ( .A(n21963), .B(n21959), .Z(n22244) );
  XNOR U24334 ( .A(n21958), .B(n21954), .Z(n22245) );
  XNOR U24335 ( .A(n21953), .B(n21949), .Z(n22246) );
  XNOR U24336 ( .A(n21948), .B(n21944), .Z(n22247) );
  XNOR U24337 ( .A(n21943), .B(n21939), .Z(n22248) );
  XNOR U24338 ( .A(n21938), .B(n21934), .Z(n22249) );
  XNOR U24339 ( .A(n21933), .B(n21929), .Z(n22250) );
  XNOR U24340 ( .A(n21928), .B(n21924), .Z(n22251) );
  XNOR U24341 ( .A(n21923), .B(n21919), .Z(n22252) );
  XNOR U24342 ( .A(n21918), .B(n21914), .Z(n22253) );
  XNOR U24343 ( .A(n21913), .B(n21909), .Z(n22254) );
  XNOR U24344 ( .A(n21908), .B(n21904), .Z(n22255) );
  XOR U24345 ( .A(n21903), .B(n21900), .Z(n22256) );
  XOR U24346 ( .A(n22257), .B(n22258), .Z(n21900) );
  XOR U24347 ( .A(n21898), .B(n22259), .Z(n22258) );
  XOR U24348 ( .A(n22260), .B(n22261), .Z(n22259) );
  XOR U24349 ( .A(n22262), .B(n22263), .Z(n22261) );
  NAND U24350 ( .A(a[5]), .B(b[62]), .Z(n22263) );
  AND U24351 ( .A(a[4]), .B(b[63]), .Z(n22262) );
  XOR U24352 ( .A(n22264), .B(n22260), .Z(n22257) );
  XOR U24353 ( .A(n22265), .B(n22266), .Z(n22260) );
  ANDN U24354 ( .B(n22267), .A(n22268), .Z(n22265) );
  AND U24355 ( .A(a[6]), .B(b[61]), .Z(n22264) );
  XOR U24356 ( .A(n22269), .B(n21898), .Z(n21899) );
  XOR U24357 ( .A(n22270), .B(n22271), .Z(n21898) );
  AND U24358 ( .A(n22272), .B(n22273), .Z(n22270) );
  AND U24359 ( .A(a[7]), .B(b[60]), .Z(n22269) );
  XOR U24360 ( .A(n22274), .B(n21903), .Z(n21905) );
  XOR U24361 ( .A(n22275), .B(n22276), .Z(n21903) );
  AND U24362 ( .A(n22277), .B(n22278), .Z(n22275) );
  AND U24363 ( .A(a[8]), .B(b[59]), .Z(n22274) );
  XOR U24364 ( .A(n22279), .B(n21908), .Z(n21910) );
  XOR U24365 ( .A(n22280), .B(n22281), .Z(n21908) );
  AND U24366 ( .A(n22282), .B(n22283), .Z(n22280) );
  AND U24367 ( .A(a[9]), .B(b[58]), .Z(n22279) );
  XOR U24368 ( .A(n22284), .B(n21913), .Z(n21915) );
  XOR U24369 ( .A(n22285), .B(n22286), .Z(n21913) );
  AND U24370 ( .A(n22287), .B(n22288), .Z(n22285) );
  AND U24371 ( .A(a[10]), .B(b[57]), .Z(n22284) );
  XOR U24372 ( .A(n22289), .B(n21918), .Z(n21920) );
  XOR U24373 ( .A(n22290), .B(n22291), .Z(n21918) );
  AND U24374 ( .A(n22292), .B(n22293), .Z(n22290) );
  AND U24375 ( .A(a[11]), .B(b[56]), .Z(n22289) );
  XOR U24376 ( .A(n22294), .B(n21923), .Z(n21925) );
  XOR U24377 ( .A(n22295), .B(n22296), .Z(n21923) );
  AND U24378 ( .A(n22297), .B(n22298), .Z(n22295) );
  AND U24379 ( .A(a[12]), .B(b[55]), .Z(n22294) );
  XOR U24380 ( .A(n22299), .B(n21928), .Z(n21930) );
  XOR U24381 ( .A(n22300), .B(n22301), .Z(n21928) );
  AND U24382 ( .A(n22302), .B(n22303), .Z(n22300) );
  AND U24383 ( .A(a[13]), .B(b[54]), .Z(n22299) );
  XOR U24384 ( .A(n22304), .B(n21933), .Z(n21935) );
  XOR U24385 ( .A(n22305), .B(n22306), .Z(n21933) );
  AND U24386 ( .A(n22307), .B(n22308), .Z(n22305) );
  AND U24387 ( .A(a[14]), .B(b[53]), .Z(n22304) );
  XOR U24388 ( .A(n22309), .B(n21938), .Z(n21940) );
  XOR U24389 ( .A(n22310), .B(n22311), .Z(n21938) );
  AND U24390 ( .A(n22312), .B(n22313), .Z(n22310) );
  AND U24391 ( .A(a[15]), .B(b[52]), .Z(n22309) );
  XOR U24392 ( .A(n22314), .B(n21943), .Z(n21945) );
  XOR U24393 ( .A(n22315), .B(n22316), .Z(n21943) );
  AND U24394 ( .A(n22317), .B(n22318), .Z(n22315) );
  AND U24395 ( .A(a[16]), .B(b[51]), .Z(n22314) );
  XOR U24396 ( .A(n22319), .B(n21948), .Z(n21950) );
  XOR U24397 ( .A(n22320), .B(n22321), .Z(n21948) );
  AND U24398 ( .A(n22322), .B(n22323), .Z(n22320) );
  AND U24399 ( .A(a[17]), .B(b[50]), .Z(n22319) );
  XOR U24400 ( .A(n22324), .B(n21953), .Z(n21955) );
  XOR U24401 ( .A(n22325), .B(n22326), .Z(n21953) );
  AND U24402 ( .A(n22327), .B(n22328), .Z(n22325) );
  AND U24403 ( .A(a[18]), .B(b[49]), .Z(n22324) );
  XOR U24404 ( .A(n22329), .B(n21958), .Z(n21960) );
  XOR U24405 ( .A(n22330), .B(n22331), .Z(n21958) );
  AND U24406 ( .A(n22332), .B(n22333), .Z(n22330) );
  AND U24407 ( .A(a[19]), .B(b[48]), .Z(n22329) );
  XOR U24408 ( .A(n22334), .B(n21963), .Z(n21965) );
  XOR U24409 ( .A(n22335), .B(n22336), .Z(n21963) );
  AND U24410 ( .A(n22337), .B(n22338), .Z(n22335) );
  AND U24411 ( .A(a[20]), .B(b[47]), .Z(n22334) );
  XOR U24412 ( .A(n22339), .B(n21968), .Z(n21970) );
  XOR U24413 ( .A(n22340), .B(n22341), .Z(n21968) );
  AND U24414 ( .A(n22342), .B(n22343), .Z(n22340) );
  AND U24415 ( .A(a[21]), .B(b[46]), .Z(n22339) );
  XOR U24416 ( .A(n22344), .B(n21973), .Z(n21975) );
  XOR U24417 ( .A(n22345), .B(n22346), .Z(n21973) );
  AND U24418 ( .A(n22347), .B(n22348), .Z(n22345) );
  AND U24419 ( .A(a[22]), .B(b[45]), .Z(n22344) );
  XOR U24420 ( .A(n22349), .B(n21978), .Z(n21980) );
  XOR U24421 ( .A(n22350), .B(n22351), .Z(n21978) );
  AND U24422 ( .A(n22352), .B(n22353), .Z(n22350) );
  AND U24423 ( .A(a[23]), .B(b[44]), .Z(n22349) );
  XOR U24424 ( .A(n22354), .B(n21983), .Z(n21985) );
  XOR U24425 ( .A(n22355), .B(n22356), .Z(n21983) );
  AND U24426 ( .A(n22357), .B(n22358), .Z(n22355) );
  AND U24427 ( .A(a[24]), .B(b[43]), .Z(n22354) );
  XOR U24428 ( .A(n22359), .B(n21988), .Z(n21990) );
  XOR U24429 ( .A(n22360), .B(n22361), .Z(n21988) );
  AND U24430 ( .A(n22362), .B(n22363), .Z(n22360) );
  AND U24431 ( .A(a[25]), .B(b[42]), .Z(n22359) );
  XOR U24432 ( .A(n22364), .B(n21993), .Z(n21995) );
  XOR U24433 ( .A(n22365), .B(n22366), .Z(n21993) );
  AND U24434 ( .A(n22367), .B(n22368), .Z(n22365) );
  AND U24435 ( .A(a[26]), .B(b[41]), .Z(n22364) );
  XOR U24436 ( .A(n22369), .B(n21998), .Z(n22000) );
  XOR U24437 ( .A(n22370), .B(n22371), .Z(n21998) );
  AND U24438 ( .A(n22372), .B(n22373), .Z(n22370) );
  AND U24439 ( .A(a[27]), .B(b[40]), .Z(n22369) );
  XOR U24440 ( .A(n22374), .B(n22003), .Z(n22005) );
  XOR U24441 ( .A(n22375), .B(n22376), .Z(n22003) );
  AND U24442 ( .A(n22377), .B(n22378), .Z(n22375) );
  AND U24443 ( .A(a[28]), .B(b[39]), .Z(n22374) );
  XOR U24444 ( .A(n22379), .B(n22008), .Z(n22010) );
  XOR U24445 ( .A(n22380), .B(n22381), .Z(n22008) );
  AND U24446 ( .A(n22382), .B(n22383), .Z(n22380) );
  AND U24447 ( .A(a[29]), .B(b[38]), .Z(n22379) );
  XOR U24448 ( .A(n22384), .B(n22013), .Z(n22015) );
  XOR U24449 ( .A(n22385), .B(n22386), .Z(n22013) );
  AND U24450 ( .A(n22387), .B(n22388), .Z(n22385) );
  AND U24451 ( .A(a[30]), .B(b[37]), .Z(n22384) );
  XOR U24452 ( .A(n22389), .B(n22018), .Z(n22020) );
  XOR U24453 ( .A(n22390), .B(n22391), .Z(n22018) );
  AND U24454 ( .A(n22392), .B(n22393), .Z(n22390) );
  AND U24455 ( .A(a[31]), .B(b[36]), .Z(n22389) );
  XOR U24456 ( .A(n22394), .B(n22023), .Z(n22025) );
  XOR U24457 ( .A(n22395), .B(n22396), .Z(n22023) );
  AND U24458 ( .A(n22397), .B(n22398), .Z(n22395) );
  AND U24459 ( .A(a[32]), .B(b[35]), .Z(n22394) );
  XOR U24460 ( .A(n22399), .B(n22028), .Z(n22030) );
  XOR U24461 ( .A(n22400), .B(n22401), .Z(n22028) );
  AND U24462 ( .A(n22402), .B(n22403), .Z(n22400) );
  AND U24463 ( .A(a[33]), .B(b[34]), .Z(n22399) );
  XOR U24464 ( .A(n22404), .B(n22033), .Z(n22035) );
  XOR U24465 ( .A(n22405), .B(n22406), .Z(n22033) );
  AND U24466 ( .A(n22407), .B(n22408), .Z(n22405) );
  AND U24467 ( .A(b[33]), .B(a[34]), .Z(n22404) );
  XOR U24468 ( .A(n22409), .B(n22410), .Z(n22037) );
  AND U24469 ( .A(n22411), .B(n22412), .Z(n22409) );
  XOR U24470 ( .A(n22413), .B(n22042), .Z(n22044) );
  XOR U24471 ( .A(n22414), .B(n22415), .Z(n22042) );
  AND U24472 ( .A(n22416), .B(n22417), .Z(n22414) );
  AND U24473 ( .A(b[32]), .B(a[35]), .Z(n22413) );
  XOR U24474 ( .A(n22419), .B(n22420), .Z(n22047) );
  AND U24475 ( .A(n22421), .B(n22422), .Z(n22419) );
  AND U24476 ( .A(b[30]), .B(a[37]), .Z(n22418) );
  XOR U24477 ( .A(n22424), .B(n22425), .Z(n22052) );
  AND U24478 ( .A(n22426), .B(n22427), .Z(n22424) );
  AND U24479 ( .A(b[29]), .B(a[38]), .Z(n22423) );
  XOR U24480 ( .A(n22429), .B(n22430), .Z(n22057) );
  AND U24481 ( .A(n22431), .B(n22432), .Z(n22429) );
  AND U24482 ( .A(b[28]), .B(a[39]), .Z(n22428) );
  XOR U24483 ( .A(n22434), .B(n22435), .Z(n22062) );
  AND U24484 ( .A(n22436), .B(n22437), .Z(n22434) );
  AND U24485 ( .A(b[27]), .B(a[40]), .Z(n22433) );
  XOR U24486 ( .A(n22439), .B(n22440), .Z(n22067) );
  AND U24487 ( .A(n22441), .B(n22442), .Z(n22439) );
  AND U24488 ( .A(b[26]), .B(a[41]), .Z(n22438) );
  XOR U24489 ( .A(n22444), .B(n22445), .Z(n22072) );
  AND U24490 ( .A(n22446), .B(n22447), .Z(n22444) );
  AND U24491 ( .A(b[25]), .B(a[42]), .Z(n22443) );
  XOR U24492 ( .A(n22449), .B(n22450), .Z(n22077) );
  AND U24493 ( .A(n22451), .B(n22452), .Z(n22449) );
  AND U24494 ( .A(b[24]), .B(a[43]), .Z(n22448) );
  XOR U24495 ( .A(n22454), .B(n22455), .Z(n22082) );
  AND U24496 ( .A(n22456), .B(n22457), .Z(n22454) );
  AND U24497 ( .A(b[23]), .B(a[44]), .Z(n22453) );
  XOR U24498 ( .A(n22459), .B(n22460), .Z(n22087) );
  AND U24499 ( .A(n22461), .B(n22462), .Z(n22459) );
  AND U24500 ( .A(b[22]), .B(a[45]), .Z(n22458) );
  XOR U24501 ( .A(n22464), .B(n22465), .Z(n22092) );
  AND U24502 ( .A(n22466), .B(n22467), .Z(n22464) );
  AND U24503 ( .A(b[21]), .B(a[46]), .Z(n22463) );
  XOR U24504 ( .A(n22469), .B(n22470), .Z(n22097) );
  AND U24505 ( .A(n22471), .B(n22472), .Z(n22469) );
  AND U24506 ( .A(b[20]), .B(a[47]), .Z(n22468) );
  XOR U24507 ( .A(n22474), .B(n22475), .Z(n22102) );
  AND U24508 ( .A(n22476), .B(n22477), .Z(n22474) );
  AND U24509 ( .A(b[19]), .B(a[48]), .Z(n22473) );
  XOR U24510 ( .A(n22479), .B(n22480), .Z(n22107) );
  AND U24511 ( .A(n22481), .B(n22482), .Z(n22479) );
  AND U24512 ( .A(b[18]), .B(a[49]), .Z(n22478) );
  XOR U24513 ( .A(n22484), .B(n22485), .Z(n22112) );
  AND U24514 ( .A(n22486), .B(n22487), .Z(n22484) );
  AND U24515 ( .A(b[17]), .B(a[50]), .Z(n22483) );
  XOR U24516 ( .A(n22489), .B(n22490), .Z(n22117) );
  AND U24517 ( .A(n22491), .B(n22492), .Z(n22489) );
  AND U24518 ( .A(b[16]), .B(a[51]), .Z(n22488) );
  XOR U24519 ( .A(n22494), .B(n22495), .Z(n22122) );
  AND U24520 ( .A(n22496), .B(n22497), .Z(n22494) );
  AND U24521 ( .A(b[15]), .B(a[52]), .Z(n22493) );
  XOR U24522 ( .A(n22499), .B(n22500), .Z(n22127) );
  AND U24523 ( .A(n22501), .B(n22502), .Z(n22499) );
  AND U24524 ( .A(b[14]), .B(a[53]), .Z(n22498) );
  XOR U24525 ( .A(n22504), .B(n22505), .Z(n22132) );
  AND U24526 ( .A(n22506), .B(n22507), .Z(n22504) );
  AND U24527 ( .A(b[13]), .B(a[54]), .Z(n22503) );
  XOR U24528 ( .A(n22509), .B(n22510), .Z(n22137) );
  AND U24529 ( .A(n22511), .B(n22512), .Z(n22509) );
  AND U24530 ( .A(b[12]), .B(a[55]), .Z(n22508) );
  XOR U24531 ( .A(n22514), .B(n22515), .Z(n22142) );
  AND U24532 ( .A(n22516), .B(n22517), .Z(n22514) );
  AND U24533 ( .A(b[11]), .B(a[56]), .Z(n22513) );
  XOR U24534 ( .A(n22519), .B(n22520), .Z(n22147) );
  AND U24535 ( .A(n22521), .B(n22522), .Z(n22519) );
  AND U24536 ( .A(b[10]), .B(a[57]), .Z(n22518) );
  XOR U24537 ( .A(n22524), .B(n22525), .Z(n22152) );
  AND U24538 ( .A(n22526), .B(n22527), .Z(n22524) );
  AND U24539 ( .A(b[9]), .B(a[58]), .Z(n22523) );
  XOR U24540 ( .A(n22529), .B(n22530), .Z(n22157) );
  AND U24541 ( .A(n22531), .B(n22532), .Z(n22529) );
  AND U24542 ( .A(b[8]), .B(a[59]), .Z(n22528) );
  XOR U24543 ( .A(n22534), .B(n22535), .Z(n22162) );
  AND U24544 ( .A(n22536), .B(n22537), .Z(n22534) );
  AND U24545 ( .A(b[7]), .B(a[60]), .Z(n22533) );
  XOR U24546 ( .A(n22539), .B(n22540), .Z(n22167) );
  AND U24547 ( .A(n22541), .B(n22542), .Z(n22539) );
  AND U24548 ( .A(b[6]), .B(a[61]), .Z(n22538) );
  XOR U24549 ( .A(n22544), .B(n22545), .Z(n22172) );
  AND U24550 ( .A(n22546), .B(n22547), .Z(n22544) );
  AND U24551 ( .A(b[5]), .B(a[62]), .Z(n22543) );
  XOR U24552 ( .A(n22549), .B(n22550), .Z(n22177) );
  AND U24553 ( .A(n22551), .B(n22552), .Z(n22549) );
  AND U24554 ( .A(b[4]), .B(a[63]), .Z(n22548) );
  XOR U24555 ( .A(n22554), .B(n22555), .Z(n22182) );
  AND U24556 ( .A(n22556), .B(n22557), .Z(n22554) );
  AND U24557 ( .A(b[3]), .B(a[64]), .Z(n22553) );
  XOR U24558 ( .A(n22559), .B(n22560), .Z(n22187) );
  OR U24559 ( .A(n22561), .B(n22562), .Z(n22560) );
  AND U24560 ( .A(b[2]), .B(a[65]), .Z(n22558) );
  XNOR U24561 ( .A(n22197), .B(n22563), .Z(n22193) );
  NAND U24562 ( .A(b[1]), .B(a[66]), .Z(n22563) );
  IV U24563 ( .A(n22191), .Z(n22197) );
  ANDN U24564 ( .B(n10353), .A(n10355), .Z(n22191) );
  NAND U24565 ( .A(a[66]), .B(b[0]), .Z(n10355) );
  XOR U24566 ( .A(n22561), .B(n22562), .Z(n10353) );
  XOR U24567 ( .A(n22565), .B(n22556), .Z(n22564) );
  XOR U24568 ( .A(n22551), .B(n22555), .Z(n22566) );
  XOR U24569 ( .A(n22546), .B(n22550), .Z(n22567) );
  XOR U24570 ( .A(n22541), .B(n22545), .Z(n22568) );
  XOR U24571 ( .A(n22536), .B(n22540), .Z(n22569) );
  XOR U24572 ( .A(n22531), .B(n22535), .Z(n22570) );
  XOR U24573 ( .A(n22526), .B(n22530), .Z(n22571) );
  XOR U24574 ( .A(n22521), .B(n22525), .Z(n22572) );
  XOR U24575 ( .A(n22516), .B(n22520), .Z(n22573) );
  XOR U24576 ( .A(n22511), .B(n22515), .Z(n22574) );
  XOR U24577 ( .A(n22506), .B(n22510), .Z(n22575) );
  XOR U24578 ( .A(n22501), .B(n22505), .Z(n22576) );
  XOR U24579 ( .A(n22496), .B(n22500), .Z(n22577) );
  XOR U24580 ( .A(n22491), .B(n22495), .Z(n22578) );
  XOR U24581 ( .A(n22486), .B(n22490), .Z(n22579) );
  XOR U24582 ( .A(n22481), .B(n22485), .Z(n22580) );
  XOR U24583 ( .A(n22476), .B(n22480), .Z(n22581) );
  XOR U24584 ( .A(n22471), .B(n22475), .Z(n22582) );
  XOR U24585 ( .A(n22466), .B(n22470), .Z(n22583) );
  XOR U24586 ( .A(n22461), .B(n22465), .Z(n22584) );
  XOR U24587 ( .A(n22456), .B(n22460), .Z(n22585) );
  XOR U24588 ( .A(n22451), .B(n22455), .Z(n22586) );
  XOR U24589 ( .A(n22446), .B(n22450), .Z(n22587) );
  XOR U24590 ( .A(n22441), .B(n22445), .Z(n22588) );
  XOR U24591 ( .A(n22436), .B(n22440), .Z(n22589) );
  XOR U24592 ( .A(n22431), .B(n22435), .Z(n22590) );
  XOR U24593 ( .A(n22426), .B(n22430), .Z(n22591) );
  XOR U24594 ( .A(n22421), .B(n22425), .Z(n22592) );
  XOR U24595 ( .A(n22411), .B(n22420), .Z(n22593) );
  XOR U24596 ( .A(n22594), .B(n22410), .Z(n22411) );
  AND U24597 ( .A(b[30]), .B(a[36]), .Z(n22594) );
  XNOR U24598 ( .A(n22410), .B(n22416), .Z(n22595) );
  XNOR U24599 ( .A(n22415), .B(n22407), .Z(n22596) );
  XNOR U24600 ( .A(n22406), .B(n22402), .Z(n22597) );
  XNOR U24601 ( .A(n22401), .B(n22397), .Z(n22598) );
  XNOR U24602 ( .A(n22396), .B(n22392), .Z(n22599) );
  XNOR U24603 ( .A(n22391), .B(n22387), .Z(n22600) );
  XNOR U24604 ( .A(n22386), .B(n22382), .Z(n22601) );
  XNOR U24605 ( .A(n22381), .B(n22377), .Z(n22602) );
  XNOR U24606 ( .A(n22376), .B(n22372), .Z(n22603) );
  XNOR U24607 ( .A(n22371), .B(n22367), .Z(n22604) );
  XNOR U24608 ( .A(n22366), .B(n22362), .Z(n22605) );
  XNOR U24609 ( .A(n22361), .B(n22357), .Z(n22606) );
  XNOR U24610 ( .A(n22356), .B(n22352), .Z(n22607) );
  XNOR U24611 ( .A(n22351), .B(n22347), .Z(n22608) );
  XNOR U24612 ( .A(n22346), .B(n22342), .Z(n22609) );
  XNOR U24613 ( .A(n22341), .B(n22337), .Z(n22610) );
  XNOR U24614 ( .A(n22336), .B(n22332), .Z(n22611) );
  XNOR U24615 ( .A(n22331), .B(n22327), .Z(n22612) );
  XNOR U24616 ( .A(n22326), .B(n22322), .Z(n22613) );
  XNOR U24617 ( .A(n22321), .B(n22317), .Z(n22614) );
  XNOR U24618 ( .A(n22316), .B(n22312), .Z(n22615) );
  XNOR U24619 ( .A(n22311), .B(n22307), .Z(n22616) );
  XNOR U24620 ( .A(n22306), .B(n22302), .Z(n22617) );
  XNOR U24621 ( .A(n22301), .B(n22297), .Z(n22618) );
  XNOR U24622 ( .A(n22296), .B(n22292), .Z(n22619) );
  XNOR U24623 ( .A(n22291), .B(n22287), .Z(n22620) );
  XNOR U24624 ( .A(n22286), .B(n22282), .Z(n22621) );
  XNOR U24625 ( .A(n22281), .B(n22277), .Z(n22622) );
  XNOR U24626 ( .A(n22276), .B(n22272), .Z(n22623) );
  XOR U24627 ( .A(n22271), .B(n22268), .Z(n22624) );
  XOR U24628 ( .A(n22625), .B(n22626), .Z(n22268) );
  XOR U24629 ( .A(n22266), .B(n22627), .Z(n22626) );
  XOR U24630 ( .A(n22628), .B(n22629), .Z(n22627) );
  XOR U24631 ( .A(n22630), .B(n22631), .Z(n22629) );
  NAND U24632 ( .A(a[4]), .B(b[62]), .Z(n22631) );
  AND U24633 ( .A(a[3]), .B(b[63]), .Z(n22630) );
  XOR U24634 ( .A(n22632), .B(n22628), .Z(n22625) );
  XOR U24635 ( .A(n22633), .B(n22634), .Z(n22628) );
  ANDN U24636 ( .B(n22635), .A(n22636), .Z(n22633) );
  AND U24637 ( .A(a[5]), .B(b[61]), .Z(n22632) );
  XOR U24638 ( .A(n22637), .B(n22266), .Z(n22267) );
  XOR U24639 ( .A(n22638), .B(n22639), .Z(n22266) );
  AND U24640 ( .A(n22640), .B(n22641), .Z(n22638) );
  AND U24641 ( .A(a[6]), .B(b[60]), .Z(n22637) );
  XOR U24642 ( .A(n22642), .B(n22271), .Z(n22273) );
  XOR U24643 ( .A(n22643), .B(n22644), .Z(n22271) );
  AND U24644 ( .A(n22645), .B(n22646), .Z(n22643) );
  AND U24645 ( .A(a[7]), .B(b[59]), .Z(n22642) );
  XOR U24646 ( .A(n22647), .B(n22276), .Z(n22278) );
  XOR U24647 ( .A(n22648), .B(n22649), .Z(n22276) );
  AND U24648 ( .A(n22650), .B(n22651), .Z(n22648) );
  AND U24649 ( .A(a[8]), .B(b[58]), .Z(n22647) );
  XOR U24650 ( .A(n22652), .B(n22281), .Z(n22283) );
  XOR U24651 ( .A(n22653), .B(n22654), .Z(n22281) );
  AND U24652 ( .A(n22655), .B(n22656), .Z(n22653) );
  AND U24653 ( .A(a[9]), .B(b[57]), .Z(n22652) );
  XOR U24654 ( .A(n22657), .B(n22286), .Z(n22288) );
  XOR U24655 ( .A(n22658), .B(n22659), .Z(n22286) );
  AND U24656 ( .A(n22660), .B(n22661), .Z(n22658) );
  AND U24657 ( .A(a[10]), .B(b[56]), .Z(n22657) );
  XOR U24658 ( .A(n22662), .B(n22291), .Z(n22293) );
  XOR U24659 ( .A(n22663), .B(n22664), .Z(n22291) );
  AND U24660 ( .A(n22665), .B(n22666), .Z(n22663) );
  AND U24661 ( .A(a[11]), .B(b[55]), .Z(n22662) );
  XOR U24662 ( .A(n22667), .B(n22296), .Z(n22298) );
  XOR U24663 ( .A(n22668), .B(n22669), .Z(n22296) );
  AND U24664 ( .A(n22670), .B(n22671), .Z(n22668) );
  AND U24665 ( .A(a[12]), .B(b[54]), .Z(n22667) );
  XOR U24666 ( .A(n22672), .B(n22301), .Z(n22303) );
  XOR U24667 ( .A(n22673), .B(n22674), .Z(n22301) );
  AND U24668 ( .A(n22675), .B(n22676), .Z(n22673) );
  AND U24669 ( .A(a[13]), .B(b[53]), .Z(n22672) );
  XOR U24670 ( .A(n22677), .B(n22306), .Z(n22308) );
  XOR U24671 ( .A(n22678), .B(n22679), .Z(n22306) );
  AND U24672 ( .A(n22680), .B(n22681), .Z(n22678) );
  AND U24673 ( .A(a[14]), .B(b[52]), .Z(n22677) );
  XOR U24674 ( .A(n22682), .B(n22311), .Z(n22313) );
  XOR U24675 ( .A(n22683), .B(n22684), .Z(n22311) );
  AND U24676 ( .A(n22685), .B(n22686), .Z(n22683) );
  AND U24677 ( .A(a[15]), .B(b[51]), .Z(n22682) );
  XOR U24678 ( .A(n22687), .B(n22316), .Z(n22318) );
  XOR U24679 ( .A(n22688), .B(n22689), .Z(n22316) );
  AND U24680 ( .A(n22690), .B(n22691), .Z(n22688) );
  AND U24681 ( .A(a[16]), .B(b[50]), .Z(n22687) );
  XOR U24682 ( .A(n22692), .B(n22321), .Z(n22323) );
  XOR U24683 ( .A(n22693), .B(n22694), .Z(n22321) );
  AND U24684 ( .A(n22695), .B(n22696), .Z(n22693) );
  AND U24685 ( .A(a[17]), .B(b[49]), .Z(n22692) );
  XOR U24686 ( .A(n22697), .B(n22326), .Z(n22328) );
  XOR U24687 ( .A(n22698), .B(n22699), .Z(n22326) );
  AND U24688 ( .A(n22700), .B(n22701), .Z(n22698) );
  AND U24689 ( .A(a[18]), .B(b[48]), .Z(n22697) );
  XOR U24690 ( .A(n22702), .B(n22331), .Z(n22333) );
  XOR U24691 ( .A(n22703), .B(n22704), .Z(n22331) );
  AND U24692 ( .A(n22705), .B(n22706), .Z(n22703) );
  AND U24693 ( .A(a[19]), .B(b[47]), .Z(n22702) );
  XOR U24694 ( .A(n22707), .B(n22336), .Z(n22338) );
  XOR U24695 ( .A(n22708), .B(n22709), .Z(n22336) );
  AND U24696 ( .A(n22710), .B(n22711), .Z(n22708) );
  AND U24697 ( .A(a[20]), .B(b[46]), .Z(n22707) );
  XOR U24698 ( .A(n22712), .B(n22341), .Z(n22343) );
  XOR U24699 ( .A(n22713), .B(n22714), .Z(n22341) );
  AND U24700 ( .A(n22715), .B(n22716), .Z(n22713) );
  AND U24701 ( .A(a[21]), .B(b[45]), .Z(n22712) );
  XOR U24702 ( .A(n22717), .B(n22346), .Z(n22348) );
  XOR U24703 ( .A(n22718), .B(n22719), .Z(n22346) );
  AND U24704 ( .A(n22720), .B(n22721), .Z(n22718) );
  AND U24705 ( .A(a[22]), .B(b[44]), .Z(n22717) );
  XOR U24706 ( .A(n22722), .B(n22351), .Z(n22353) );
  XOR U24707 ( .A(n22723), .B(n22724), .Z(n22351) );
  AND U24708 ( .A(n22725), .B(n22726), .Z(n22723) );
  AND U24709 ( .A(a[23]), .B(b[43]), .Z(n22722) );
  XOR U24710 ( .A(n22727), .B(n22356), .Z(n22358) );
  XOR U24711 ( .A(n22728), .B(n22729), .Z(n22356) );
  AND U24712 ( .A(n22730), .B(n22731), .Z(n22728) );
  AND U24713 ( .A(a[24]), .B(b[42]), .Z(n22727) );
  XOR U24714 ( .A(n22732), .B(n22361), .Z(n22363) );
  XOR U24715 ( .A(n22733), .B(n22734), .Z(n22361) );
  AND U24716 ( .A(n22735), .B(n22736), .Z(n22733) );
  AND U24717 ( .A(a[25]), .B(b[41]), .Z(n22732) );
  XOR U24718 ( .A(n22737), .B(n22366), .Z(n22368) );
  XOR U24719 ( .A(n22738), .B(n22739), .Z(n22366) );
  AND U24720 ( .A(n22740), .B(n22741), .Z(n22738) );
  AND U24721 ( .A(a[26]), .B(b[40]), .Z(n22737) );
  XOR U24722 ( .A(n22742), .B(n22371), .Z(n22373) );
  XOR U24723 ( .A(n22743), .B(n22744), .Z(n22371) );
  AND U24724 ( .A(n22745), .B(n22746), .Z(n22743) );
  AND U24725 ( .A(a[27]), .B(b[39]), .Z(n22742) );
  XOR U24726 ( .A(n22747), .B(n22376), .Z(n22378) );
  XOR U24727 ( .A(n22748), .B(n22749), .Z(n22376) );
  AND U24728 ( .A(n22750), .B(n22751), .Z(n22748) );
  AND U24729 ( .A(a[28]), .B(b[38]), .Z(n22747) );
  XOR U24730 ( .A(n22752), .B(n22381), .Z(n22383) );
  XOR U24731 ( .A(n22753), .B(n22754), .Z(n22381) );
  AND U24732 ( .A(n22755), .B(n22756), .Z(n22753) );
  AND U24733 ( .A(a[29]), .B(b[37]), .Z(n22752) );
  XOR U24734 ( .A(n22757), .B(n22386), .Z(n22388) );
  XOR U24735 ( .A(n22758), .B(n22759), .Z(n22386) );
  AND U24736 ( .A(n22760), .B(n22761), .Z(n22758) );
  AND U24737 ( .A(a[30]), .B(b[36]), .Z(n22757) );
  XOR U24738 ( .A(n22762), .B(n22391), .Z(n22393) );
  XOR U24739 ( .A(n22763), .B(n22764), .Z(n22391) );
  AND U24740 ( .A(n22765), .B(n22766), .Z(n22763) );
  AND U24741 ( .A(a[31]), .B(b[35]), .Z(n22762) );
  XOR U24742 ( .A(n22767), .B(n22396), .Z(n22398) );
  XOR U24743 ( .A(n22768), .B(n22769), .Z(n22396) );
  AND U24744 ( .A(n22770), .B(n22771), .Z(n22768) );
  AND U24745 ( .A(a[32]), .B(b[34]), .Z(n22767) );
  XOR U24746 ( .A(n22772), .B(n22401), .Z(n22403) );
  XOR U24747 ( .A(n22773), .B(n22774), .Z(n22401) );
  AND U24748 ( .A(n22775), .B(n22776), .Z(n22773) );
  AND U24749 ( .A(a[33]), .B(b[33]), .Z(n22772) );
  XOR U24750 ( .A(n22777), .B(n22406), .Z(n22408) );
  XOR U24751 ( .A(n22778), .B(n22779), .Z(n22406) );
  AND U24752 ( .A(n22780), .B(n22781), .Z(n22778) );
  AND U24753 ( .A(b[32]), .B(a[34]), .Z(n22777) );
  XOR U24754 ( .A(n22782), .B(n22783), .Z(n22410) );
  AND U24755 ( .A(n22784), .B(n22785), .Z(n22782) );
  XOR U24756 ( .A(n22786), .B(n22415), .Z(n22417) );
  XOR U24757 ( .A(n22787), .B(n22788), .Z(n22415) );
  AND U24758 ( .A(n22789), .B(n22790), .Z(n22787) );
  AND U24759 ( .A(b[31]), .B(a[35]), .Z(n22786) );
  XOR U24760 ( .A(n22792), .B(n22793), .Z(n22420) );
  AND U24761 ( .A(n22794), .B(n22795), .Z(n22792) );
  AND U24762 ( .A(b[29]), .B(a[37]), .Z(n22791) );
  XOR U24763 ( .A(n22797), .B(n22798), .Z(n22425) );
  AND U24764 ( .A(n22799), .B(n22800), .Z(n22797) );
  AND U24765 ( .A(b[28]), .B(a[38]), .Z(n22796) );
  XOR U24766 ( .A(n22802), .B(n22803), .Z(n22430) );
  AND U24767 ( .A(n22804), .B(n22805), .Z(n22802) );
  AND U24768 ( .A(b[27]), .B(a[39]), .Z(n22801) );
  XOR U24769 ( .A(n22807), .B(n22808), .Z(n22435) );
  AND U24770 ( .A(n22809), .B(n22810), .Z(n22807) );
  AND U24771 ( .A(b[26]), .B(a[40]), .Z(n22806) );
  XOR U24772 ( .A(n22812), .B(n22813), .Z(n22440) );
  AND U24773 ( .A(n22814), .B(n22815), .Z(n22812) );
  AND U24774 ( .A(b[25]), .B(a[41]), .Z(n22811) );
  XOR U24775 ( .A(n22817), .B(n22818), .Z(n22445) );
  AND U24776 ( .A(n22819), .B(n22820), .Z(n22817) );
  AND U24777 ( .A(b[24]), .B(a[42]), .Z(n22816) );
  XOR U24778 ( .A(n22822), .B(n22823), .Z(n22450) );
  AND U24779 ( .A(n22824), .B(n22825), .Z(n22822) );
  AND U24780 ( .A(b[23]), .B(a[43]), .Z(n22821) );
  XOR U24781 ( .A(n22827), .B(n22828), .Z(n22455) );
  AND U24782 ( .A(n22829), .B(n22830), .Z(n22827) );
  AND U24783 ( .A(b[22]), .B(a[44]), .Z(n22826) );
  XOR U24784 ( .A(n22832), .B(n22833), .Z(n22460) );
  AND U24785 ( .A(n22834), .B(n22835), .Z(n22832) );
  AND U24786 ( .A(b[21]), .B(a[45]), .Z(n22831) );
  XOR U24787 ( .A(n22837), .B(n22838), .Z(n22465) );
  AND U24788 ( .A(n22839), .B(n22840), .Z(n22837) );
  AND U24789 ( .A(b[20]), .B(a[46]), .Z(n22836) );
  XOR U24790 ( .A(n22842), .B(n22843), .Z(n22470) );
  AND U24791 ( .A(n22844), .B(n22845), .Z(n22842) );
  AND U24792 ( .A(b[19]), .B(a[47]), .Z(n22841) );
  XOR U24793 ( .A(n22847), .B(n22848), .Z(n22475) );
  AND U24794 ( .A(n22849), .B(n22850), .Z(n22847) );
  AND U24795 ( .A(b[18]), .B(a[48]), .Z(n22846) );
  XOR U24796 ( .A(n22852), .B(n22853), .Z(n22480) );
  AND U24797 ( .A(n22854), .B(n22855), .Z(n22852) );
  AND U24798 ( .A(b[17]), .B(a[49]), .Z(n22851) );
  XOR U24799 ( .A(n22857), .B(n22858), .Z(n22485) );
  AND U24800 ( .A(n22859), .B(n22860), .Z(n22857) );
  AND U24801 ( .A(b[16]), .B(a[50]), .Z(n22856) );
  XOR U24802 ( .A(n22862), .B(n22863), .Z(n22490) );
  AND U24803 ( .A(n22864), .B(n22865), .Z(n22862) );
  AND U24804 ( .A(b[15]), .B(a[51]), .Z(n22861) );
  XOR U24805 ( .A(n22867), .B(n22868), .Z(n22495) );
  AND U24806 ( .A(n22869), .B(n22870), .Z(n22867) );
  AND U24807 ( .A(b[14]), .B(a[52]), .Z(n22866) );
  XOR U24808 ( .A(n22872), .B(n22873), .Z(n22500) );
  AND U24809 ( .A(n22874), .B(n22875), .Z(n22872) );
  AND U24810 ( .A(b[13]), .B(a[53]), .Z(n22871) );
  XOR U24811 ( .A(n22877), .B(n22878), .Z(n22505) );
  AND U24812 ( .A(n22879), .B(n22880), .Z(n22877) );
  AND U24813 ( .A(b[12]), .B(a[54]), .Z(n22876) );
  XOR U24814 ( .A(n22882), .B(n22883), .Z(n22510) );
  AND U24815 ( .A(n22884), .B(n22885), .Z(n22882) );
  AND U24816 ( .A(b[11]), .B(a[55]), .Z(n22881) );
  XOR U24817 ( .A(n22887), .B(n22888), .Z(n22515) );
  AND U24818 ( .A(n22889), .B(n22890), .Z(n22887) );
  AND U24819 ( .A(b[10]), .B(a[56]), .Z(n22886) );
  XOR U24820 ( .A(n22892), .B(n22893), .Z(n22520) );
  AND U24821 ( .A(n22894), .B(n22895), .Z(n22892) );
  AND U24822 ( .A(b[9]), .B(a[57]), .Z(n22891) );
  XOR U24823 ( .A(n22897), .B(n22898), .Z(n22525) );
  AND U24824 ( .A(n22899), .B(n22900), .Z(n22897) );
  AND U24825 ( .A(b[8]), .B(a[58]), .Z(n22896) );
  XOR U24826 ( .A(n22902), .B(n22903), .Z(n22530) );
  AND U24827 ( .A(n22904), .B(n22905), .Z(n22902) );
  AND U24828 ( .A(b[7]), .B(a[59]), .Z(n22901) );
  XOR U24829 ( .A(n22907), .B(n22908), .Z(n22535) );
  AND U24830 ( .A(n22909), .B(n22910), .Z(n22907) );
  AND U24831 ( .A(b[6]), .B(a[60]), .Z(n22906) );
  XOR U24832 ( .A(n22912), .B(n22913), .Z(n22540) );
  AND U24833 ( .A(n22914), .B(n22915), .Z(n22912) );
  AND U24834 ( .A(b[5]), .B(a[61]), .Z(n22911) );
  XOR U24835 ( .A(n22917), .B(n22918), .Z(n22545) );
  AND U24836 ( .A(n22919), .B(n22920), .Z(n22917) );
  AND U24837 ( .A(b[4]), .B(a[62]), .Z(n22916) );
  XOR U24838 ( .A(n22922), .B(n22923), .Z(n22550) );
  AND U24839 ( .A(n22924), .B(n22925), .Z(n22922) );
  AND U24840 ( .A(b[3]), .B(a[63]), .Z(n22921) );
  XOR U24841 ( .A(n22927), .B(n22928), .Z(n22555) );
  OR U24842 ( .A(n22929), .B(n22930), .Z(n22928) );
  AND U24843 ( .A(b[2]), .B(a[64]), .Z(n22926) );
  XNOR U24844 ( .A(n22565), .B(n22931), .Z(n22561) );
  NAND U24845 ( .A(b[1]), .B(a[65]), .Z(n22931) );
  IV U24846 ( .A(n22559), .Z(n22565) );
  ANDN U24847 ( .B(n10356), .A(n10358), .Z(n22559) );
  NAND U24848 ( .A(a[65]), .B(b[0]), .Z(n10358) );
  XOR U24849 ( .A(n22929), .B(n22930), .Z(n10356) );
  XOR U24850 ( .A(n22933), .B(n22924), .Z(n22932) );
  XOR U24851 ( .A(n22919), .B(n22923), .Z(n22934) );
  XOR U24852 ( .A(n22914), .B(n22918), .Z(n22935) );
  XOR U24853 ( .A(n22909), .B(n22913), .Z(n22936) );
  XOR U24854 ( .A(n22904), .B(n22908), .Z(n22937) );
  XOR U24855 ( .A(n22899), .B(n22903), .Z(n22938) );
  XOR U24856 ( .A(n22894), .B(n22898), .Z(n22939) );
  XOR U24857 ( .A(n22889), .B(n22893), .Z(n22940) );
  XOR U24858 ( .A(n22884), .B(n22888), .Z(n22941) );
  XOR U24859 ( .A(n22879), .B(n22883), .Z(n22942) );
  XOR U24860 ( .A(n22874), .B(n22878), .Z(n22943) );
  XOR U24861 ( .A(n22869), .B(n22873), .Z(n22944) );
  XOR U24862 ( .A(n22864), .B(n22868), .Z(n22945) );
  XOR U24863 ( .A(n22859), .B(n22863), .Z(n22946) );
  XOR U24864 ( .A(n22854), .B(n22858), .Z(n22947) );
  XOR U24865 ( .A(n22849), .B(n22853), .Z(n22948) );
  XOR U24866 ( .A(n22844), .B(n22848), .Z(n22949) );
  XOR U24867 ( .A(n22839), .B(n22843), .Z(n22950) );
  XOR U24868 ( .A(n22834), .B(n22838), .Z(n22951) );
  XOR U24869 ( .A(n22829), .B(n22833), .Z(n22952) );
  XOR U24870 ( .A(n22824), .B(n22828), .Z(n22953) );
  XOR U24871 ( .A(n22819), .B(n22823), .Z(n22954) );
  XOR U24872 ( .A(n22814), .B(n22818), .Z(n22955) );
  XOR U24873 ( .A(n22809), .B(n22813), .Z(n22956) );
  XOR U24874 ( .A(n22804), .B(n22808), .Z(n22957) );
  XOR U24875 ( .A(n22799), .B(n22803), .Z(n22958) );
  XOR U24876 ( .A(n22794), .B(n22798), .Z(n22959) );
  XOR U24877 ( .A(n22784), .B(n22793), .Z(n22960) );
  XOR U24878 ( .A(n22961), .B(n22783), .Z(n22784) );
  AND U24879 ( .A(b[29]), .B(a[36]), .Z(n22961) );
  XNOR U24880 ( .A(n22783), .B(n22789), .Z(n22962) );
  XNOR U24881 ( .A(n22788), .B(n22780), .Z(n22963) );
  XNOR U24882 ( .A(n22779), .B(n22775), .Z(n22964) );
  XNOR U24883 ( .A(n22774), .B(n22770), .Z(n22965) );
  XNOR U24884 ( .A(n22769), .B(n22765), .Z(n22966) );
  XNOR U24885 ( .A(n22764), .B(n22760), .Z(n22967) );
  XNOR U24886 ( .A(n22759), .B(n22755), .Z(n22968) );
  XNOR U24887 ( .A(n22754), .B(n22750), .Z(n22969) );
  XNOR U24888 ( .A(n22749), .B(n22745), .Z(n22970) );
  XNOR U24889 ( .A(n22744), .B(n22740), .Z(n22971) );
  XNOR U24890 ( .A(n22739), .B(n22735), .Z(n22972) );
  XNOR U24891 ( .A(n22734), .B(n22730), .Z(n22973) );
  XNOR U24892 ( .A(n22729), .B(n22725), .Z(n22974) );
  XNOR U24893 ( .A(n22724), .B(n22720), .Z(n22975) );
  XNOR U24894 ( .A(n22719), .B(n22715), .Z(n22976) );
  XNOR U24895 ( .A(n22714), .B(n22710), .Z(n22977) );
  XNOR U24896 ( .A(n22709), .B(n22705), .Z(n22978) );
  XNOR U24897 ( .A(n22704), .B(n22700), .Z(n22979) );
  XNOR U24898 ( .A(n22699), .B(n22695), .Z(n22980) );
  XNOR U24899 ( .A(n22694), .B(n22690), .Z(n22981) );
  XNOR U24900 ( .A(n22689), .B(n22685), .Z(n22982) );
  XNOR U24901 ( .A(n22684), .B(n22680), .Z(n22983) );
  XNOR U24902 ( .A(n22679), .B(n22675), .Z(n22984) );
  XNOR U24903 ( .A(n22674), .B(n22670), .Z(n22985) );
  XNOR U24904 ( .A(n22669), .B(n22665), .Z(n22986) );
  XNOR U24905 ( .A(n22664), .B(n22660), .Z(n22987) );
  XNOR U24906 ( .A(n22659), .B(n22655), .Z(n22988) );
  XNOR U24907 ( .A(n22654), .B(n22650), .Z(n22989) );
  XNOR U24908 ( .A(n22649), .B(n22645), .Z(n22990) );
  XNOR U24909 ( .A(n22644), .B(n22640), .Z(n22991) );
  XOR U24910 ( .A(n22639), .B(n22636), .Z(n22992) );
  XOR U24911 ( .A(n22993), .B(n22994), .Z(n22636) );
  XOR U24912 ( .A(n22634), .B(n22995), .Z(n22994) );
  XOR U24913 ( .A(n22996), .B(n22997), .Z(n22995) );
  XOR U24914 ( .A(n22998), .B(n22999), .Z(n22997) );
  NAND U24915 ( .A(a[3]), .B(b[62]), .Z(n22999) );
  AND U24916 ( .A(a[2]), .B(b[63]), .Z(n22998) );
  XOR U24917 ( .A(n23000), .B(n22996), .Z(n22993) );
  XOR U24918 ( .A(n23001), .B(n23002), .Z(n22996) );
  ANDN U24919 ( .B(n23003), .A(n23004), .Z(n23001) );
  AND U24920 ( .A(a[4]), .B(b[61]), .Z(n23000) );
  XOR U24921 ( .A(n23005), .B(n22634), .Z(n22635) );
  XOR U24922 ( .A(n23006), .B(n23007), .Z(n22634) );
  AND U24923 ( .A(n23008), .B(n23009), .Z(n23006) );
  AND U24924 ( .A(a[5]), .B(b[60]), .Z(n23005) );
  XOR U24925 ( .A(n23010), .B(n22639), .Z(n22641) );
  XOR U24926 ( .A(n23011), .B(n23012), .Z(n22639) );
  AND U24927 ( .A(n23013), .B(n23014), .Z(n23011) );
  AND U24928 ( .A(a[6]), .B(b[59]), .Z(n23010) );
  XOR U24929 ( .A(n23015), .B(n22644), .Z(n22646) );
  XOR U24930 ( .A(n23016), .B(n23017), .Z(n22644) );
  AND U24931 ( .A(n23018), .B(n23019), .Z(n23016) );
  AND U24932 ( .A(a[7]), .B(b[58]), .Z(n23015) );
  XOR U24933 ( .A(n23020), .B(n22649), .Z(n22651) );
  XOR U24934 ( .A(n23021), .B(n23022), .Z(n22649) );
  AND U24935 ( .A(n23023), .B(n23024), .Z(n23021) );
  AND U24936 ( .A(a[8]), .B(b[57]), .Z(n23020) );
  XOR U24937 ( .A(n23025), .B(n22654), .Z(n22656) );
  XOR U24938 ( .A(n23026), .B(n23027), .Z(n22654) );
  AND U24939 ( .A(n23028), .B(n23029), .Z(n23026) );
  AND U24940 ( .A(a[9]), .B(b[56]), .Z(n23025) );
  XOR U24941 ( .A(n23030), .B(n22659), .Z(n22661) );
  XOR U24942 ( .A(n23031), .B(n23032), .Z(n22659) );
  AND U24943 ( .A(n23033), .B(n23034), .Z(n23031) );
  AND U24944 ( .A(a[10]), .B(b[55]), .Z(n23030) );
  XOR U24945 ( .A(n23035), .B(n22664), .Z(n22666) );
  XOR U24946 ( .A(n23036), .B(n23037), .Z(n22664) );
  AND U24947 ( .A(n23038), .B(n23039), .Z(n23036) );
  AND U24948 ( .A(a[11]), .B(b[54]), .Z(n23035) );
  XOR U24949 ( .A(n23040), .B(n22669), .Z(n22671) );
  XOR U24950 ( .A(n23041), .B(n23042), .Z(n22669) );
  AND U24951 ( .A(n23043), .B(n23044), .Z(n23041) );
  AND U24952 ( .A(a[12]), .B(b[53]), .Z(n23040) );
  XOR U24953 ( .A(n23045), .B(n22674), .Z(n22676) );
  XOR U24954 ( .A(n23046), .B(n23047), .Z(n22674) );
  AND U24955 ( .A(n23048), .B(n23049), .Z(n23046) );
  AND U24956 ( .A(a[13]), .B(b[52]), .Z(n23045) );
  XOR U24957 ( .A(n23050), .B(n22679), .Z(n22681) );
  XOR U24958 ( .A(n23051), .B(n23052), .Z(n22679) );
  AND U24959 ( .A(n23053), .B(n23054), .Z(n23051) );
  AND U24960 ( .A(a[14]), .B(b[51]), .Z(n23050) );
  XOR U24961 ( .A(n23055), .B(n22684), .Z(n22686) );
  XOR U24962 ( .A(n23056), .B(n23057), .Z(n22684) );
  AND U24963 ( .A(n23058), .B(n23059), .Z(n23056) );
  AND U24964 ( .A(a[15]), .B(b[50]), .Z(n23055) );
  XOR U24965 ( .A(n23060), .B(n22689), .Z(n22691) );
  XOR U24966 ( .A(n23061), .B(n23062), .Z(n22689) );
  AND U24967 ( .A(n23063), .B(n23064), .Z(n23061) );
  AND U24968 ( .A(a[16]), .B(b[49]), .Z(n23060) );
  XOR U24969 ( .A(n23065), .B(n22694), .Z(n22696) );
  XOR U24970 ( .A(n23066), .B(n23067), .Z(n22694) );
  AND U24971 ( .A(n23068), .B(n23069), .Z(n23066) );
  AND U24972 ( .A(a[17]), .B(b[48]), .Z(n23065) );
  XOR U24973 ( .A(n23070), .B(n22699), .Z(n22701) );
  XOR U24974 ( .A(n23071), .B(n23072), .Z(n22699) );
  AND U24975 ( .A(n23073), .B(n23074), .Z(n23071) );
  AND U24976 ( .A(a[18]), .B(b[47]), .Z(n23070) );
  XOR U24977 ( .A(n23075), .B(n22704), .Z(n22706) );
  XOR U24978 ( .A(n23076), .B(n23077), .Z(n22704) );
  AND U24979 ( .A(n23078), .B(n23079), .Z(n23076) );
  AND U24980 ( .A(a[19]), .B(b[46]), .Z(n23075) );
  XOR U24981 ( .A(n23080), .B(n22709), .Z(n22711) );
  XOR U24982 ( .A(n23081), .B(n23082), .Z(n22709) );
  AND U24983 ( .A(n23083), .B(n23084), .Z(n23081) );
  AND U24984 ( .A(a[20]), .B(b[45]), .Z(n23080) );
  XOR U24985 ( .A(n23085), .B(n22714), .Z(n22716) );
  XOR U24986 ( .A(n23086), .B(n23087), .Z(n22714) );
  AND U24987 ( .A(n23088), .B(n23089), .Z(n23086) );
  AND U24988 ( .A(a[21]), .B(b[44]), .Z(n23085) );
  XOR U24989 ( .A(n23090), .B(n22719), .Z(n22721) );
  XOR U24990 ( .A(n23091), .B(n23092), .Z(n22719) );
  AND U24991 ( .A(n23093), .B(n23094), .Z(n23091) );
  AND U24992 ( .A(a[22]), .B(b[43]), .Z(n23090) );
  XOR U24993 ( .A(n23095), .B(n22724), .Z(n22726) );
  XOR U24994 ( .A(n23096), .B(n23097), .Z(n22724) );
  AND U24995 ( .A(n23098), .B(n23099), .Z(n23096) );
  AND U24996 ( .A(a[23]), .B(b[42]), .Z(n23095) );
  XOR U24997 ( .A(n23100), .B(n22729), .Z(n22731) );
  XOR U24998 ( .A(n23101), .B(n23102), .Z(n22729) );
  AND U24999 ( .A(n23103), .B(n23104), .Z(n23101) );
  AND U25000 ( .A(a[24]), .B(b[41]), .Z(n23100) );
  XOR U25001 ( .A(n23105), .B(n22734), .Z(n22736) );
  XOR U25002 ( .A(n23106), .B(n23107), .Z(n22734) );
  AND U25003 ( .A(n23108), .B(n23109), .Z(n23106) );
  AND U25004 ( .A(a[25]), .B(b[40]), .Z(n23105) );
  XOR U25005 ( .A(n23110), .B(n22739), .Z(n22741) );
  XOR U25006 ( .A(n23111), .B(n23112), .Z(n22739) );
  AND U25007 ( .A(n23113), .B(n23114), .Z(n23111) );
  AND U25008 ( .A(a[26]), .B(b[39]), .Z(n23110) );
  XOR U25009 ( .A(n23115), .B(n22744), .Z(n22746) );
  XOR U25010 ( .A(n23116), .B(n23117), .Z(n22744) );
  AND U25011 ( .A(n23118), .B(n23119), .Z(n23116) );
  AND U25012 ( .A(a[27]), .B(b[38]), .Z(n23115) );
  XOR U25013 ( .A(n23120), .B(n22749), .Z(n22751) );
  XOR U25014 ( .A(n23121), .B(n23122), .Z(n22749) );
  AND U25015 ( .A(n23123), .B(n23124), .Z(n23121) );
  AND U25016 ( .A(a[28]), .B(b[37]), .Z(n23120) );
  XOR U25017 ( .A(n23125), .B(n22754), .Z(n22756) );
  XOR U25018 ( .A(n23126), .B(n23127), .Z(n22754) );
  AND U25019 ( .A(n23128), .B(n23129), .Z(n23126) );
  AND U25020 ( .A(a[29]), .B(b[36]), .Z(n23125) );
  XOR U25021 ( .A(n23130), .B(n22759), .Z(n22761) );
  XOR U25022 ( .A(n23131), .B(n23132), .Z(n22759) );
  AND U25023 ( .A(n23133), .B(n23134), .Z(n23131) );
  AND U25024 ( .A(a[30]), .B(b[35]), .Z(n23130) );
  XOR U25025 ( .A(n23135), .B(n22764), .Z(n22766) );
  XOR U25026 ( .A(n23136), .B(n23137), .Z(n22764) );
  AND U25027 ( .A(n23138), .B(n23139), .Z(n23136) );
  AND U25028 ( .A(a[31]), .B(b[34]), .Z(n23135) );
  XOR U25029 ( .A(n23140), .B(n22769), .Z(n22771) );
  XOR U25030 ( .A(n23141), .B(n23142), .Z(n22769) );
  AND U25031 ( .A(n23143), .B(n23144), .Z(n23141) );
  AND U25032 ( .A(a[32]), .B(b[33]), .Z(n23140) );
  XOR U25033 ( .A(n23145), .B(n22774), .Z(n22776) );
  XOR U25034 ( .A(n23146), .B(n23147), .Z(n22774) );
  AND U25035 ( .A(n23148), .B(n23149), .Z(n23146) );
  AND U25036 ( .A(b[32]), .B(a[33]), .Z(n23145) );
  XOR U25037 ( .A(n23150), .B(n22779), .Z(n22781) );
  XOR U25038 ( .A(n23151), .B(n23152), .Z(n22779) );
  AND U25039 ( .A(n23153), .B(n23154), .Z(n23151) );
  AND U25040 ( .A(b[31]), .B(a[34]), .Z(n23150) );
  XOR U25041 ( .A(n23155), .B(n23156), .Z(n22783) );
  AND U25042 ( .A(n23157), .B(n23158), .Z(n23155) );
  XOR U25043 ( .A(n23159), .B(n22788), .Z(n22790) );
  XOR U25044 ( .A(n23160), .B(n23161), .Z(n22788) );
  AND U25045 ( .A(n23162), .B(n23163), .Z(n23160) );
  AND U25046 ( .A(b[30]), .B(a[35]), .Z(n23159) );
  XNOR U25047 ( .A(n23165), .B(n23166), .Z(n22793) );
  AND U25048 ( .A(n23167), .B(n23168), .Z(n23165) );
  AND U25049 ( .A(b[28]), .B(a[37]), .Z(n23164) );
  XNOR U25050 ( .A(n23170), .B(n23171), .Z(n22798) );
  AND U25051 ( .A(n23172), .B(n23173), .Z(n23170) );
  AND U25052 ( .A(b[27]), .B(a[38]), .Z(n23169) );
  XNOR U25053 ( .A(n23175), .B(n23176), .Z(n22803) );
  AND U25054 ( .A(n23177), .B(n23178), .Z(n23175) );
  AND U25055 ( .A(b[26]), .B(a[39]), .Z(n23174) );
  XNOR U25056 ( .A(n23180), .B(n23181), .Z(n22808) );
  AND U25057 ( .A(n23182), .B(n23183), .Z(n23180) );
  AND U25058 ( .A(b[25]), .B(a[40]), .Z(n23179) );
  XNOR U25059 ( .A(n23185), .B(n23186), .Z(n22813) );
  AND U25060 ( .A(n23187), .B(n23188), .Z(n23185) );
  AND U25061 ( .A(b[24]), .B(a[41]), .Z(n23184) );
  XNOR U25062 ( .A(n23190), .B(n23191), .Z(n22818) );
  AND U25063 ( .A(n23192), .B(n23193), .Z(n23190) );
  AND U25064 ( .A(b[23]), .B(a[42]), .Z(n23189) );
  XNOR U25065 ( .A(n23195), .B(n23196), .Z(n22823) );
  AND U25066 ( .A(n23197), .B(n23198), .Z(n23195) );
  AND U25067 ( .A(b[22]), .B(a[43]), .Z(n23194) );
  XNOR U25068 ( .A(n23200), .B(n23201), .Z(n22828) );
  AND U25069 ( .A(n23202), .B(n23203), .Z(n23200) );
  AND U25070 ( .A(b[21]), .B(a[44]), .Z(n23199) );
  XNOR U25071 ( .A(n23205), .B(n23206), .Z(n22833) );
  AND U25072 ( .A(n23207), .B(n23208), .Z(n23205) );
  AND U25073 ( .A(b[20]), .B(a[45]), .Z(n23204) );
  XNOR U25074 ( .A(n23210), .B(n23211), .Z(n22838) );
  AND U25075 ( .A(n23212), .B(n23213), .Z(n23210) );
  AND U25076 ( .A(b[19]), .B(a[46]), .Z(n23209) );
  XNOR U25077 ( .A(n23215), .B(n23216), .Z(n22843) );
  AND U25078 ( .A(n23217), .B(n23218), .Z(n23215) );
  AND U25079 ( .A(b[18]), .B(a[47]), .Z(n23214) );
  XNOR U25080 ( .A(n23220), .B(n23221), .Z(n22848) );
  AND U25081 ( .A(n23222), .B(n23223), .Z(n23220) );
  AND U25082 ( .A(b[17]), .B(a[48]), .Z(n23219) );
  XNOR U25083 ( .A(n23225), .B(n23226), .Z(n22853) );
  AND U25084 ( .A(n23227), .B(n23228), .Z(n23225) );
  AND U25085 ( .A(b[16]), .B(a[49]), .Z(n23224) );
  XNOR U25086 ( .A(n23230), .B(n23231), .Z(n22858) );
  AND U25087 ( .A(n23232), .B(n23233), .Z(n23230) );
  AND U25088 ( .A(b[15]), .B(a[50]), .Z(n23229) );
  XNOR U25089 ( .A(n23235), .B(n23236), .Z(n22863) );
  AND U25090 ( .A(n23237), .B(n23238), .Z(n23235) );
  AND U25091 ( .A(b[14]), .B(a[51]), .Z(n23234) );
  XNOR U25092 ( .A(n23240), .B(n23241), .Z(n22868) );
  AND U25093 ( .A(n23242), .B(n23243), .Z(n23240) );
  AND U25094 ( .A(b[13]), .B(a[52]), .Z(n23239) );
  XNOR U25095 ( .A(n23245), .B(n23246), .Z(n22873) );
  AND U25096 ( .A(n23247), .B(n23248), .Z(n23245) );
  AND U25097 ( .A(b[12]), .B(a[53]), .Z(n23244) );
  XNOR U25098 ( .A(n23250), .B(n23251), .Z(n22878) );
  AND U25099 ( .A(n23252), .B(n23253), .Z(n23250) );
  AND U25100 ( .A(b[11]), .B(a[54]), .Z(n23249) );
  XNOR U25101 ( .A(n23255), .B(n23256), .Z(n22883) );
  AND U25102 ( .A(n23257), .B(n23258), .Z(n23255) );
  AND U25103 ( .A(b[10]), .B(a[55]), .Z(n23254) );
  XNOR U25104 ( .A(n23260), .B(n23261), .Z(n22888) );
  AND U25105 ( .A(n23262), .B(n23263), .Z(n23260) );
  AND U25106 ( .A(b[9]), .B(a[56]), .Z(n23259) );
  XNOR U25107 ( .A(n23265), .B(n23266), .Z(n22893) );
  AND U25108 ( .A(n23267), .B(n23268), .Z(n23265) );
  AND U25109 ( .A(b[8]), .B(a[57]), .Z(n23264) );
  XNOR U25110 ( .A(n23270), .B(n23271), .Z(n22898) );
  AND U25111 ( .A(n23272), .B(n23273), .Z(n23270) );
  AND U25112 ( .A(b[7]), .B(a[58]), .Z(n23269) );
  XNOR U25113 ( .A(n23275), .B(n23276), .Z(n22903) );
  AND U25114 ( .A(n23277), .B(n23278), .Z(n23275) );
  AND U25115 ( .A(b[6]), .B(a[59]), .Z(n23274) );
  XNOR U25116 ( .A(n23280), .B(n23281), .Z(n22908) );
  AND U25117 ( .A(n23282), .B(n23283), .Z(n23280) );
  AND U25118 ( .A(b[5]), .B(a[60]), .Z(n23279) );
  XNOR U25119 ( .A(n23285), .B(n23286), .Z(n22913) );
  AND U25120 ( .A(n23287), .B(n23288), .Z(n23285) );
  AND U25121 ( .A(b[4]), .B(a[61]), .Z(n23284) );
  XOR U25122 ( .A(n23290), .B(n23291), .Z(n22918) );
  AND U25123 ( .A(n23292), .B(n23293), .Z(n23290) );
  AND U25124 ( .A(b[3]), .B(a[62]), .Z(n23289) );
  XOR U25125 ( .A(n23295), .B(n23296), .Z(n22923) );
  OR U25126 ( .A(n23297), .B(n23298), .Z(n23296) );
  AND U25127 ( .A(b[2]), .B(a[63]), .Z(n23294) );
  XNOR U25128 ( .A(n22933), .B(n23299), .Z(n22929) );
  NAND U25129 ( .A(b[1]), .B(a[64]), .Z(n23299) );
  IV U25130 ( .A(n22927), .Z(n22933) );
  ANDN U25131 ( .B(n10359), .A(n10361), .Z(n22927) );
  NAND U25132 ( .A(a[64]), .B(b[0]), .Z(n10361) );
  XOR U25133 ( .A(n23297), .B(n23298), .Z(n10359) );
  XOR U25134 ( .A(n23301), .B(n23292), .Z(n23300) );
  XOR U25135 ( .A(n23287), .B(n23291), .Z(n23302) );
  XNOR U25136 ( .A(n23282), .B(n23286), .Z(n23303) );
  XNOR U25137 ( .A(n23277), .B(n23281), .Z(n23304) );
  XNOR U25138 ( .A(n23272), .B(n23276), .Z(n23305) );
  XNOR U25139 ( .A(n23267), .B(n23271), .Z(n23306) );
  XNOR U25140 ( .A(n23262), .B(n23266), .Z(n23307) );
  XNOR U25141 ( .A(n23257), .B(n23261), .Z(n23308) );
  XNOR U25142 ( .A(n23252), .B(n23256), .Z(n23309) );
  XNOR U25143 ( .A(n23247), .B(n23251), .Z(n23310) );
  XNOR U25144 ( .A(n23242), .B(n23246), .Z(n23311) );
  XNOR U25145 ( .A(n23237), .B(n23241), .Z(n23312) );
  XNOR U25146 ( .A(n23232), .B(n23236), .Z(n23313) );
  XNOR U25147 ( .A(n23227), .B(n23231), .Z(n23314) );
  XNOR U25148 ( .A(n23222), .B(n23226), .Z(n23315) );
  XNOR U25149 ( .A(n23217), .B(n23221), .Z(n23316) );
  XNOR U25150 ( .A(n23212), .B(n23216), .Z(n23317) );
  XNOR U25151 ( .A(n23207), .B(n23211), .Z(n23318) );
  XNOR U25152 ( .A(n23202), .B(n23206), .Z(n23319) );
  XNOR U25153 ( .A(n23197), .B(n23201), .Z(n23320) );
  XNOR U25154 ( .A(n23192), .B(n23196), .Z(n23321) );
  XNOR U25155 ( .A(n23187), .B(n23191), .Z(n23322) );
  XNOR U25156 ( .A(n23182), .B(n23186), .Z(n23323) );
  XNOR U25157 ( .A(n23177), .B(n23181), .Z(n23324) );
  XNOR U25158 ( .A(n23172), .B(n23176), .Z(n23325) );
  XNOR U25159 ( .A(n23167), .B(n23171), .Z(n23326) );
  XNOR U25160 ( .A(n23157), .B(n23166), .Z(n23327) );
  XOR U25161 ( .A(n23328), .B(n23156), .Z(n23157) );
  AND U25162 ( .A(b[28]), .B(a[36]), .Z(n23328) );
  XNOR U25163 ( .A(n23156), .B(n23162), .Z(n23329) );
  XNOR U25164 ( .A(n23161), .B(n23153), .Z(n23330) );
  XNOR U25165 ( .A(n23152), .B(n23148), .Z(n23331) );
  XNOR U25166 ( .A(n23147), .B(n23143), .Z(n23332) );
  XNOR U25167 ( .A(n23142), .B(n23138), .Z(n23333) );
  XNOR U25168 ( .A(n23137), .B(n23133), .Z(n23334) );
  XNOR U25169 ( .A(n23132), .B(n23128), .Z(n23335) );
  XNOR U25170 ( .A(n23127), .B(n23123), .Z(n23336) );
  XNOR U25171 ( .A(n23122), .B(n23118), .Z(n23337) );
  XNOR U25172 ( .A(n23117), .B(n23113), .Z(n23338) );
  XNOR U25173 ( .A(n23112), .B(n23108), .Z(n23339) );
  XNOR U25174 ( .A(n23107), .B(n23103), .Z(n23340) );
  XNOR U25175 ( .A(n23102), .B(n23098), .Z(n23341) );
  XNOR U25176 ( .A(n23097), .B(n23093), .Z(n23342) );
  XNOR U25177 ( .A(n23092), .B(n23088), .Z(n23343) );
  XNOR U25178 ( .A(n23087), .B(n23083), .Z(n23344) );
  XNOR U25179 ( .A(n23082), .B(n23078), .Z(n23345) );
  XNOR U25180 ( .A(n23077), .B(n23073), .Z(n23346) );
  XNOR U25181 ( .A(n23072), .B(n23068), .Z(n23347) );
  XNOR U25182 ( .A(n23067), .B(n23063), .Z(n23348) );
  XNOR U25183 ( .A(n23062), .B(n23058), .Z(n23349) );
  XNOR U25184 ( .A(n23057), .B(n23053), .Z(n23350) );
  XNOR U25185 ( .A(n23052), .B(n23048), .Z(n23351) );
  XNOR U25186 ( .A(n23047), .B(n23043), .Z(n23352) );
  XNOR U25187 ( .A(n23042), .B(n23038), .Z(n23353) );
  XNOR U25188 ( .A(n23037), .B(n23033), .Z(n23354) );
  XNOR U25189 ( .A(n23032), .B(n23028), .Z(n23355) );
  XNOR U25190 ( .A(n23027), .B(n23023), .Z(n23356) );
  XNOR U25191 ( .A(n23022), .B(n23018), .Z(n23357) );
  XNOR U25192 ( .A(n23017), .B(n23013), .Z(n23358) );
  XNOR U25193 ( .A(n23012), .B(n23008), .Z(n23359) );
  XOR U25194 ( .A(n23007), .B(n23004), .Z(n23360) );
  XOR U25195 ( .A(n23361), .B(n23362), .Z(n23004) );
  XOR U25196 ( .A(n23002), .B(n23363), .Z(n23362) );
  XOR U25197 ( .A(n23364), .B(n23365), .Z(n23363) );
  XOR U25198 ( .A(n23366), .B(n23367), .Z(n23365) );
  NAND U25199 ( .A(a[2]), .B(b[62]), .Z(n23367) );
  AND U25200 ( .A(a[1]), .B(b[63]), .Z(n23366) );
  XOR U25201 ( .A(n23368), .B(n23364), .Z(n23361) );
  XOR U25202 ( .A(n23369), .B(n23370), .Z(n23364) );
  ANDN U25203 ( .B(n23371), .A(n23372), .Z(n23369) );
  AND U25204 ( .A(a[3]), .B(b[61]), .Z(n23368) );
  XOR U25205 ( .A(n23373), .B(n23002), .Z(n23003) );
  XOR U25206 ( .A(n23374), .B(n23375), .Z(n23002) );
  AND U25207 ( .A(n23376), .B(n23377), .Z(n23374) );
  AND U25208 ( .A(a[4]), .B(b[60]), .Z(n23373) );
  XOR U25209 ( .A(n23378), .B(n23007), .Z(n23009) );
  XOR U25210 ( .A(n23379), .B(n23380), .Z(n23007) );
  AND U25211 ( .A(n23381), .B(n23382), .Z(n23379) );
  AND U25212 ( .A(a[5]), .B(b[59]), .Z(n23378) );
  XOR U25213 ( .A(n23383), .B(n23012), .Z(n23014) );
  XOR U25214 ( .A(n23384), .B(n23385), .Z(n23012) );
  AND U25215 ( .A(n23386), .B(n23387), .Z(n23384) );
  AND U25216 ( .A(a[6]), .B(b[58]), .Z(n23383) );
  XOR U25217 ( .A(n23388), .B(n23017), .Z(n23019) );
  XOR U25218 ( .A(n23389), .B(n23390), .Z(n23017) );
  AND U25219 ( .A(n23391), .B(n23392), .Z(n23389) );
  AND U25220 ( .A(a[7]), .B(b[57]), .Z(n23388) );
  XOR U25221 ( .A(n23393), .B(n23022), .Z(n23024) );
  XOR U25222 ( .A(n23394), .B(n23395), .Z(n23022) );
  AND U25223 ( .A(n23396), .B(n23397), .Z(n23394) );
  AND U25224 ( .A(a[8]), .B(b[56]), .Z(n23393) );
  XOR U25225 ( .A(n23398), .B(n23027), .Z(n23029) );
  XOR U25226 ( .A(n23399), .B(n23400), .Z(n23027) );
  AND U25227 ( .A(n23401), .B(n23402), .Z(n23399) );
  AND U25228 ( .A(a[9]), .B(b[55]), .Z(n23398) );
  XOR U25229 ( .A(n23403), .B(n23032), .Z(n23034) );
  XOR U25230 ( .A(n23404), .B(n23405), .Z(n23032) );
  AND U25231 ( .A(n23406), .B(n23407), .Z(n23404) );
  AND U25232 ( .A(a[10]), .B(b[54]), .Z(n23403) );
  XOR U25233 ( .A(n23408), .B(n23037), .Z(n23039) );
  XOR U25234 ( .A(n23409), .B(n23410), .Z(n23037) );
  AND U25235 ( .A(n23411), .B(n23412), .Z(n23409) );
  AND U25236 ( .A(a[11]), .B(b[53]), .Z(n23408) );
  XOR U25237 ( .A(n23413), .B(n23042), .Z(n23044) );
  XOR U25238 ( .A(n23414), .B(n23415), .Z(n23042) );
  AND U25239 ( .A(n23416), .B(n23417), .Z(n23414) );
  AND U25240 ( .A(a[12]), .B(b[52]), .Z(n23413) );
  XOR U25241 ( .A(n23418), .B(n23047), .Z(n23049) );
  XOR U25242 ( .A(n23419), .B(n23420), .Z(n23047) );
  AND U25243 ( .A(n23421), .B(n23422), .Z(n23419) );
  AND U25244 ( .A(a[13]), .B(b[51]), .Z(n23418) );
  XOR U25245 ( .A(n23423), .B(n23052), .Z(n23054) );
  XOR U25246 ( .A(n23424), .B(n23425), .Z(n23052) );
  AND U25247 ( .A(n23426), .B(n23427), .Z(n23424) );
  AND U25248 ( .A(a[14]), .B(b[50]), .Z(n23423) );
  XOR U25249 ( .A(n23428), .B(n23057), .Z(n23059) );
  XOR U25250 ( .A(n23429), .B(n23430), .Z(n23057) );
  AND U25251 ( .A(n23431), .B(n23432), .Z(n23429) );
  AND U25252 ( .A(a[15]), .B(b[49]), .Z(n23428) );
  XOR U25253 ( .A(n23433), .B(n23062), .Z(n23064) );
  XOR U25254 ( .A(n23434), .B(n23435), .Z(n23062) );
  AND U25255 ( .A(n23436), .B(n23437), .Z(n23434) );
  AND U25256 ( .A(a[16]), .B(b[48]), .Z(n23433) );
  XOR U25257 ( .A(n23438), .B(n23067), .Z(n23069) );
  XOR U25258 ( .A(n23439), .B(n23440), .Z(n23067) );
  AND U25259 ( .A(n23441), .B(n23442), .Z(n23439) );
  AND U25260 ( .A(a[17]), .B(b[47]), .Z(n23438) );
  XOR U25261 ( .A(n23443), .B(n23072), .Z(n23074) );
  XOR U25262 ( .A(n23444), .B(n23445), .Z(n23072) );
  AND U25263 ( .A(n23446), .B(n23447), .Z(n23444) );
  AND U25264 ( .A(a[18]), .B(b[46]), .Z(n23443) );
  XOR U25265 ( .A(n23448), .B(n23077), .Z(n23079) );
  XOR U25266 ( .A(n23449), .B(n23450), .Z(n23077) );
  AND U25267 ( .A(n23451), .B(n23452), .Z(n23449) );
  AND U25268 ( .A(a[19]), .B(b[45]), .Z(n23448) );
  XOR U25269 ( .A(n23453), .B(n23082), .Z(n23084) );
  XOR U25270 ( .A(n23454), .B(n23455), .Z(n23082) );
  AND U25271 ( .A(n23456), .B(n23457), .Z(n23454) );
  AND U25272 ( .A(a[20]), .B(b[44]), .Z(n23453) );
  XOR U25273 ( .A(n23458), .B(n23087), .Z(n23089) );
  XOR U25274 ( .A(n23459), .B(n23460), .Z(n23087) );
  AND U25275 ( .A(n23461), .B(n23462), .Z(n23459) );
  AND U25276 ( .A(a[21]), .B(b[43]), .Z(n23458) );
  XOR U25277 ( .A(n23463), .B(n23092), .Z(n23094) );
  XOR U25278 ( .A(n23464), .B(n23465), .Z(n23092) );
  AND U25279 ( .A(n23466), .B(n23467), .Z(n23464) );
  AND U25280 ( .A(a[22]), .B(b[42]), .Z(n23463) );
  XOR U25281 ( .A(n23468), .B(n23097), .Z(n23099) );
  XOR U25282 ( .A(n23469), .B(n23470), .Z(n23097) );
  AND U25283 ( .A(n23471), .B(n23472), .Z(n23469) );
  AND U25284 ( .A(a[23]), .B(b[41]), .Z(n23468) );
  XOR U25285 ( .A(n23473), .B(n23102), .Z(n23104) );
  XOR U25286 ( .A(n23474), .B(n23475), .Z(n23102) );
  AND U25287 ( .A(n23476), .B(n23477), .Z(n23474) );
  AND U25288 ( .A(a[24]), .B(b[40]), .Z(n23473) );
  XOR U25289 ( .A(n23478), .B(n23107), .Z(n23109) );
  XOR U25290 ( .A(n23479), .B(n23480), .Z(n23107) );
  AND U25291 ( .A(n23481), .B(n23482), .Z(n23479) );
  AND U25292 ( .A(a[25]), .B(b[39]), .Z(n23478) );
  XOR U25293 ( .A(n23483), .B(n23112), .Z(n23114) );
  XOR U25294 ( .A(n23484), .B(n23485), .Z(n23112) );
  AND U25295 ( .A(n23486), .B(n23487), .Z(n23484) );
  AND U25296 ( .A(a[26]), .B(b[38]), .Z(n23483) );
  XOR U25297 ( .A(n23488), .B(n23117), .Z(n23119) );
  XOR U25298 ( .A(n23489), .B(n23490), .Z(n23117) );
  AND U25299 ( .A(n23491), .B(n23492), .Z(n23489) );
  AND U25300 ( .A(a[27]), .B(b[37]), .Z(n23488) );
  XOR U25301 ( .A(n23493), .B(n23122), .Z(n23124) );
  XOR U25302 ( .A(n23494), .B(n23495), .Z(n23122) );
  AND U25303 ( .A(n23496), .B(n23497), .Z(n23494) );
  AND U25304 ( .A(a[28]), .B(b[36]), .Z(n23493) );
  XOR U25305 ( .A(n23498), .B(n23127), .Z(n23129) );
  XOR U25306 ( .A(n23499), .B(n23500), .Z(n23127) );
  AND U25307 ( .A(n23501), .B(n23502), .Z(n23499) );
  AND U25308 ( .A(a[29]), .B(b[35]), .Z(n23498) );
  XOR U25309 ( .A(n23503), .B(n23132), .Z(n23134) );
  XOR U25310 ( .A(n23504), .B(n23505), .Z(n23132) );
  AND U25311 ( .A(n23506), .B(n23507), .Z(n23504) );
  AND U25312 ( .A(a[30]), .B(b[34]), .Z(n23503) );
  XOR U25313 ( .A(n23508), .B(n23137), .Z(n23139) );
  XOR U25314 ( .A(n23509), .B(n23510), .Z(n23137) );
  AND U25315 ( .A(n23511), .B(n23512), .Z(n23509) );
  AND U25316 ( .A(a[31]), .B(b[33]), .Z(n23508) );
  XOR U25317 ( .A(n23513), .B(n23142), .Z(n23144) );
  XOR U25318 ( .A(n23514), .B(n23515), .Z(n23142) );
  AND U25319 ( .A(n23516), .B(n23517), .Z(n23514) );
  AND U25320 ( .A(a[32]), .B(b[32]), .Z(n23513) );
  XOR U25321 ( .A(n23518), .B(n23147), .Z(n23149) );
  XOR U25322 ( .A(n23519), .B(n23520), .Z(n23147) );
  AND U25323 ( .A(n23521), .B(n23522), .Z(n23519) );
  AND U25324 ( .A(b[31]), .B(a[33]), .Z(n23518) );
  XOR U25325 ( .A(n23523), .B(n23152), .Z(n23154) );
  XOR U25326 ( .A(n23524), .B(n23525), .Z(n23152) );
  AND U25327 ( .A(n23526), .B(n23527), .Z(n23524) );
  AND U25328 ( .A(b[30]), .B(a[34]), .Z(n23523) );
  XOR U25329 ( .A(n23528), .B(n23529), .Z(n23156) );
  AND U25330 ( .A(n23530), .B(n23531), .Z(n23528) );
  XOR U25331 ( .A(n23532), .B(n23161), .Z(n23163) );
  XOR U25332 ( .A(n23533), .B(n23534), .Z(n23161) );
  AND U25333 ( .A(n23535), .B(n23536), .Z(n23533) );
  AND U25334 ( .A(b[29]), .B(a[35]), .Z(n23532) );
  XOR U25335 ( .A(n23537), .B(n23166), .Z(n23168) );
  XOR U25336 ( .A(n23538), .B(n23539), .Z(n23166) );
  AND U25337 ( .A(n23540), .B(n23541), .Z(n23538) );
  AND U25338 ( .A(b[27]), .B(a[37]), .Z(n23537) );
  XOR U25339 ( .A(n23542), .B(n23171), .Z(n23173) );
  XOR U25340 ( .A(n23543), .B(n23544), .Z(n23171) );
  AND U25341 ( .A(n23545), .B(n23546), .Z(n23543) );
  AND U25342 ( .A(b[26]), .B(a[38]), .Z(n23542) );
  XOR U25343 ( .A(n23547), .B(n23176), .Z(n23178) );
  XOR U25344 ( .A(n23548), .B(n23549), .Z(n23176) );
  AND U25345 ( .A(n23550), .B(n23551), .Z(n23548) );
  AND U25346 ( .A(b[25]), .B(a[39]), .Z(n23547) );
  XOR U25347 ( .A(n23552), .B(n23181), .Z(n23183) );
  XOR U25348 ( .A(n23553), .B(n23554), .Z(n23181) );
  AND U25349 ( .A(n23555), .B(n23556), .Z(n23553) );
  AND U25350 ( .A(b[24]), .B(a[40]), .Z(n23552) );
  XOR U25351 ( .A(n23557), .B(n23186), .Z(n23188) );
  XOR U25352 ( .A(n23558), .B(n23559), .Z(n23186) );
  AND U25353 ( .A(n23560), .B(n23561), .Z(n23558) );
  AND U25354 ( .A(b[23]), .B(a[41]), .Z(n23557) );
  XOR U25355 ( .A(n23562), .B(n23191), .Z(n23193) );
  XOR U25356 ( .A(n23563), .B(n23564), .Z(n23191) );
  AND U25357 ( .A(n23565), .B(n23566), .Z(n23563) );
  AND U25358 ( .A(b[22]), .B(a[42]), .Z(n23562) );
  XOR U25359 ( .A(n23567), .B(n23196), .Z(n23198) );
  XOR U25360 ( .A(n23568), .B(n23569), .Z(n23196) );
  AND U25361 ( .A(n23570), .B(n23571), .Z(n23568) );
  AND U25362 ( .A(b[21]), .B(a[43]), .Z(n23567) );
  XOR U25363 ( .A(n23572), .B(n23201), .Z(n23203) );
  XOR U25364 ( .A(n23573), .B(n23574), .Z(n23201) );
  AND U25365 ( .A(n23575), .B(n23576), .Z(n23573) );
  AND U25366 ( .A(b[20]), .B(a[44]), .Z(n23572) );
  XOR U25367 ( .A(n23577), .B(n23206), .Z(n23208) );
  XOR U25368 ( .A(n23578), .B(n23579), .Z(n23206) );
  AND U25369 ( .A(n23580), .B(n23581), .Z(n23578) );
  AND U25370 ( .A(b[19]), .B(a[45]), .Z(n23577) );
  XOR U25371 ( .A(n23582), .B(n23211), .Z(n23213) );
  XOR U25372 ( .A(n23583), .B(n23584), .Z(n23211) );
  AND U25373 ( .A(n23585), .B(n23586), .Z(n23583) );
  AND U25374 ( .A(b[18]), .B(a[46]), .Z(n23582) );
  XOR U25375 ( .A(n23587), .B(n23216), .Z(n23218) );
  XOR U25376 ( .A(n23588), .B(n23589), .Z(n23216) );
  AND U25377 ( .A(n23590), .B(n23591), .Z(n23588) );
  AND U25378 ( .A(b[17]), .B(a[47]), .Z(n23587) );
  XOR U25379 ( .A(n23592), .B(n23221), .Z(n23223) );
  XOR U25380 ( .A(n23593), .B(n23594), .Z(n23221) );
  AND U25381 ( .A(n23595), .B(n23596), .Z(n23593) );
  AND U25382 ( .A(b[16]), .B(a[48]), .Z(n23592) );
  XOR U25383 ( .A(n23597), .B(n23226), .Z(n23228) );
  XOR U25384 ( .A(n23598), .B(n23599), .Z(n23226) );
  AND U25385 ( .A(n23600), .B(n23601), .Z(n23598) );
  AND U25386 ( .A(b[15]), .B(a[49]), .Z(n23597) );
  XOR U25387 ( .A(n23602), .B(n23231), .Z(n23233) );
  XOR U25388 ( .A(n23603), .B(n23604), .Z(n23231) );
  AND U25389 ( .A(n23605), .B(n23606), .Z(n23603) );
  AND U25390 ( .A(b[14]), .B(a[50]), .Z(n23602) );
  XOR U25391 ( .A(n23607), .B(n23236), .Z(n23238) );
  XOR U25392 ( .A(n23608), .B(n23609), .Z(n23236) );
  AND U25393 ( .A(n23610), .B(n23611), .Z(n23608) );
  AND U25394 ( .A(b[13]), .B(a[51]), .Z(n23607) );
  XOR U25395 ( .A(n23612), .B(n23241), .Z(n23243) );
  XOR U25396 ( .A(n23613), .B(n23614), .Z(n23241) );
  AND U25397 ( .A(n23615), .B(n23616), .Z(n23613) );
  AND U25398 ( .A(b[12]), .B(a[52]), .Z(n23612) );
  XOR U25399 ( .A(n23617), .B(n23246), .Z(n23248) );
  XOR U25400 ( .A(n23618), .B(n23619), .Z(n23246) );
  AND U25401 ( .A(n23620), .B(n23621), .Z(n23618) );
  AND U25402 ( .A(b[11]), .B(a[53]), .Z(n23617) );
  XOR U25403 ( .A(n23622), .B(n23251), .Z(n23253) );
  XOR U25404 ( .A(n23623), .B(n23624), .Z(n23251) );
  AND U25405 ( .A(n23625), .B(n23626), .Z(n23623) );
  AND U25406 ( .A(b[10]), .B(a[54]), .Z(n23622) );
  XOR U25407 ( .A(n23627), .B(n23256), .Z(n23258) );
  XOR U25408 ( .A(n23628), .B(n23629), .Z(n23256) );
  AND U25409 ( .A(n23630), .B(n23631), .Z(n23628) );
  AND U25410 ( .A(b[9]), .B(a[55]), .Z(n23627) );
  XOR U25411 ( .A(n23632), .B(n23261), .Z(n23263) );
  XOR U25412 ( .A(n23633), .B(n23634), .Z(n23261) );
  AND U25413 ( .A(n23635), .B(n23636), .Z(n23633) );
  AND U25414 ( .A(b[8]), .B(a[56]), .Z(n23632) );
  XOR U25415 ( .A(n23637), .B(n23266), .Z(n23268) );
  XOR U25416 ( .A(n23638), .B(n23639), .Z(n23266) );
  AND U25417 ( .A(n23640), .B(n23641), .Z(n23638) );
  AND U25418 ( .A(b[7]), .B(a[57]), .Z(n23637) );
  XOR U25419 ( .A(n23642), .B(n23271), .Z(n23273) );
  XOR U25420 ( .A(n23643), .B(n23644), .Z(n23271) );
  AND U25421 ( .A(n23645), .B(n23646), .Z(n23643) );
  AND U25422 ( .A(b[6]), .B(a[58]), .Z(n23642) );
  XOR U25423 ( .A(n23647), .B(n23276), .Z(n23278) );
  XOR U25424 ( .A(n23648), .B(n23649), .Z(n23276) );
  AND U25425 ( .A(n23650), .B(n23651), .Z(n23648) );
  AND U25426 ( .A(b[5]), .B(a[59]), .Z(n23647) );
  XOR U25427 ( .A(n23652), .B(n23281), .Z(n23283) );
  XOR U25428 ( .A(n23653), .B(n23654), .Z(n23281) );
  AND U25429 ( .A(n23655), .B(n23656), .Z(n23653) );
  AND U25430 ( .A(b[4]), .B(a[60]), .Z(n23652) );
  XOR U25431 ( .A(n23657), .B(n23286), .Z(n23288) );
  XNOR U25432 ( .A(n23658), .B(n23659), .Z(n23286) );
  ANDN U25433 ( .B(n23660), .A(n23661), .Z(n23658) );
  AND U25434 ( .A(b[3]), .B(a[61]), .Z(n23657) );
  XOR U25435 ( .A(n23663), .B(n23664), .Z(n23291) );
  OR U25436 ( .A(n23665), .B(n23666), .Z(n23664) );
  AND U25437 ( .A(b[2]), .B(a[62]), .Z(n23662) );
  XNOR U25438 ( .A(n23301), .B(n23667), .Z(n23297) );
  NAND U25439 ( .A(b[1]), .B(a[63]), .Z(n23667) );
  IV U25440 ( .A(n23295), .Z(n23301) );
  ANDN U25441 ( .B(n23668), .A(n23669), .Z(n23295) );
  NAND U25442 ( .A(a[97]), .B(b[0]), .Z(n10262) );
  NAND U25443 ( .A(a[98]), .B(b[0]), .Z(n10259) );
  XOR U25444 ( .A(n23670), .B(n23671), .Z(c[99]) );
  XOR U25445 ( .A(n23672), .B(n23673), .Z(c[98]) );
  XOR U25446 ( .A(n23674), .B(n23675), .Z(c[97]) );
  XOR U25447 ( .A(n23676), .B(n23677), .Z(c[96]) );
  XOR U25448 ( .A(n23678), .B(n23679), .Z(c[95]) );
  XOR U25449 ( .A(n23680), .B(n23681), .Z(c[94]) );
  XOR U25450 ( .A(n23682), .B(n23683), .Z(c[93]) );
  XOR U25451 ( .A(n23684), .B(n23685), .Z(c[92]) );
  XOR U25452 ( .A(n23686), .B(n23687), .Z(c[91]) );
  XOR U25453 ( .A(n23688), .B(n23689), .Z(c[90]) );
  XOR U25454 ( .A(n23690), .B(n23691), .Z(c[89]) );
  XOR U25455 ( .A(n23692), .B(n23693), .Z(c[88]) );
  XOR U25456 ( .A(n23694), .B(n23695), .Z(c[87]) );
  XOR U25457 ( .A(n23696), .B(n23697), .Z(c[86]) );
  XOR U25458 ( .A(n23698), .B(n23699), .Z(c[85]) );
  XOR U25459 ( .A(n23700), .B(n23701), .Z(c[84]) );
  XOR U25460 ( .A(n23702), .B(n23703), .Z(c[83]) );
  XOR U25461 ( .A(n23704), .B(n23705), .Z(c[82]) );
  XOR U25462 ( .A(n23706), .B(n23707), .Z(c[81]) );
  XOR U25463 ( .A(n23708), .B(n23709), .Z(c[80]) );
  XOR U25464 ( .A(n23710), .B(n23711), .Z(c[79]) );
  XOR U25465 ( .A(n23712), .B(n23713), .Z(c[78]) );
  XOR U25466 ( .A(n23714), .B(n23715), .Z(c[77]) );
  XOR U25467 ( .A(n23716), .B(n23717), .Z(c[76]) );
  XOR U25468 ( .A(n23718), .B(n23719), .Z(c[75]) );
  XOR U25469 ( .A(n23720), .B(n23721), .Z(c[74]) );
  XOR U25470 ( .A(n23722), .B(n23723), .Z(c[73]) );
  XOR U25471 ( .A(n23724), .B(n23725), .Z(c[72]) );
  XOR U25472 ( .A(n23726), .B(n23727), .Z(c[71]) );
  XOR U25473 ( .A(n23728), .B(n23729), .Z(c[70]) );
  XOR U25474 ( .A(n23730), .B(n23731), .Z(c[69]) );
  XOR U25475 ( .A(n23732), .B(n23733), .Z(c[68]) );
  XOR U25476 ( .A(n23734), .B(n23735), .Z(c[67]) );
  XOR U25477 ( .A(n23736), .B(n23737), .Z(c[66]) );
  XOR U25478 ( .A(n23738), .B(n23739), .Z(c[65]) );
  XNOR U25479 ( .A(sreg[128]), .B(n23740), .Z(c[64]) );
  XOR U25480 ( .A(n10365), .B(n10364), .Z(c[127]) );
  XOR U25481 ( .A(sreg[191]), .B(n10363), .Z(n10364) );
  XOR U25482 ( .A(n23668), .B(n23741), .Z(n10365) );
  XNOR U25483 ( .A(n23669), .B(n10363), .Z(n23741) );
  XOR U25484 ( .A(n23742), .B(n23743), .Z(n10363) );
  NOR U25485 ( .A(n23744), .B(n23745), .Z(n23742) );
  NAND U25486 ( .A(a[63]), .B(b[0]), .Z(n23669) );
  XOR U25487 ( .A(n23666), .B(n23665), .Z(n23668) );
  XOR U25488 ( .A(n23663), .B(n23746), .Z(n23665) );
  NAND U25489 ( .A(b[1]), .B(a[62]), .Z(n23746) );
  XOR U25490 ( .A(n23663), .B(n23661), .Z(n23747) );
  XOR U25491 ( .A(n23748), .B(n23659), .Z(n23661) );
  AND U25492 ( .A(b[2]), .B(a[61]), .Z(n23748) );
  ANDN U25493 ( .B(n23749), .A(n23750), .Z(n23663) );
  XOR U25494 ( .A(n23659), .B(n23655), .Z(n23751) );
  XNOR U25495 ( .A(n23654), .B(n23650), .Z(n23752) );
  XNOR U25496 ( .A(n23649), .B(n23645), .Z(n23753) );
  XNOR U25497 ( .A(n23644), .B(n23640), .Z(n23754) );
  XNOR U25498 ( .A(n23639), .B(n23635), .Z(n23755) );
  XNOR U25499 ( .A(n23634), .B(n23630), .Z(n23756) );
  XNOR U25500 ( .A(n23629), .B(n23625), .Z(n23757) );
  XNOR U25501 ( .A(n23624), .B(n23620), .Z(n23758) );
  XNOR U25502 ( .A(n23619), .B(n23615), .Z(n23759) );
  XNOR U25503 ( .A(n23614), .B(n23610), .Z(n23760) );
  XNOR U25504 ( .A(n23609), .B(n23605), .Z(n23761) );
  XNOR U25505 ( .A(n23604), .B(n23600), .Z(n23762) );
  XNOR U25506 ( .A(n23599), .B(n23595), .Z(n23763) );
  XNOR U25507 ( .A(n23594), .B(n23590), .Z(n23764) );
  XNOR U25508 ( .A(n23589), .B(n23585), .Z(n23765) );
  XNOR U25509 ( .A(n23584), .B(n23580), .Z(n23766) );
  XNOR U25510 ( .A(n23579), .B(n23575), .Z(n23767) );
  XNOR U25511 ( .A(n23574), .B(n23570), .Z(n23768) );
  XNOR U25512 ( .A(n23569), .B(n23565), .Z(n23769) );
  XNOR U25513 ( .A(n23564), .B(n23560), .Z(n23770) );
  XNOR U25514 ( .A(n23559), .B(n23555), .Z(n23771) );
  XNOR U25515 ( .A(n23554), .B(n23550), .Z(n23772) );
  XNOR U25516 ( .A(n23549), .B(n23545), .Z(n23773) );
  XNOR U25517 ( .A(n23544), .B(n23540), .Z(n23774) );
  XNOR U25518 ( .A(n23539), .B(n23530), .Z(n23775) );
  XNOR U25519 ( .A(n23529), .B(n23535), .Z(n23776) );
  XNOR U25520 ( .A(n23534), .B(n23526), .Z(n23777) );
  XNOR U25521 ( .A(n23525), .B(n23521), .Z(n23778) );
  XNOR U25522 ( .A(n23520), .B(n23516), .Z(n23779) );
  XNOR U25523 ( .A(n23515), .B(n23511), .Z(n23780) );
  XNOR U25524 ( .A(n23510), .B(n23506), .Z(n23781) );
  XNOR U25525 ( .A(n23505), .B(n23501), .Z(n23782) );
  XNOR U25526 ( .A(n23500), .B(n23496), .Z(n23783) );
  XNOR U25527 ( .A(n23495), .B(n23491), .Z(n23784) );
  XNOR U25528 ( .A(n23490), .B(n23486), .Z(n23785) );
  XNOR U25529 ( .A(n23485), .B(n23481), .Z(n23786) );
  XNOR U25530 ( .A(n23480), .B(n23476), .Z(n23787) );
  XNOR U25531 ( .A(n23475), .B(n23471), .Z(n23788) );
  XNOR U25532 ( .A(n23470), .B(n23466), .Z(n23789) );
  XNOR U25533 ( .A(n23465), .B(n23461), .Z(n23790) );
  XNOR U25534 ( .A(n23460), .B(n23456), .Z(n23791) );
  XNOR U25535 ( .A(n23455), .B(n23451), .Z(n23792) );
  XNOR U25536 ( .A(n23450), .B(n23446), .Z(n23793) );
  XNOR U25537 ( .A(n23445), .B(n23441), .Z(n23794) );
  XNOR U25538 ( .A(n23440), .B(n23436), .Z(n23795) );
  XNOR U25539 ( .A(n23435), .B(n23431), .Z(n23796) );
  XNOR U25540 ( .A(n23430), .B(n23426), .Z(n23797) );
  XNOR U25541 ( .A(n23425), .B(n23421), .Z(n23798) );
  XNOR U25542 ( .A(n23420), .B(n23416), .Z(n23799) );
  XNOR U25543 ( .A(n23415), .B(n23411), .Z(n23800) );
  XNOR U25544 ( .A(n23410), .B(n23406), .Z(n23801) );
  XNOR U25545 ( .A(n23405), .B(n23401), .Z(n23802) );
  XNOR U25546 ( .A(n23400), .B(n23396), .Z(n23803) );
  XNOR U25547 ( .A(n23395), .B(n23391), .Z(n23804) );
  XNOR U25548 ( .A(n23390), .B(n23386), .Z(n23805) );
  XNOR U25549 ( .A(n23385), .B(n23381), .Z(n23806) );
  XNOR U25550 ( .A(n23380), .B(n23376), .Z(n23807) );
  XOR U25551 ( .A(n23375), .B(n23372), .Z(n23808) );
  XOR U25552 ( .A(n23809), .B(n23810), .Z(n23372) );
  XOR U25553 ( .A(n23370), .B(n23811), .Z(n23810) );
  XOR U25554 ( .A(n23812), .B(n23813), .Z(n23811) );
  XOR U25555 ( .A(n23814), .B(n23815), .Z(n23813) );
  NAND U25556 ( .A(a[1]), .B(b[62]), .Z(n23815) );
  AND U25557 ( .A(a[0]), .B(b[63]), .Z(n23814) );
  XOR U25558 ( .A(n23816), .B(n23812), .Z(n23809) );
  XOR U25559 ( .A(n23817), .B(n23818), .Z(n23812) );
  ANDN U25560 ( .B(n23819), .A(n23820), .Z(n23817) );
  AND U25561 ( .A(a[2]), .B(b[61]), .Z(n23816) );
  XOR U25562 ( .A(n23821), .B(n23370), .Z(n23371) );
  XOR U25563 ( .A(n23822), .B(n23823), .Z(n23370) );
  AND U25564 ( .A(n23824), .B(n23825), .Z(n23822) );
  AND U25565 ( .A(a[3]), .B(b[60]), .Z(n23821) );
  XOR U25566 ( .A(n23826), .B(n23375), .Z(n23377) );
  XOR U25567 ( .A(n23827), .B(n23828), .Z(n23375) );
  AND U25568 ( .A(n23829), .B(n23830), .Z(n23827) );
  AND U25569 ( .A(a[4]), .B(b[59]), .Z(n23826) );
  XOR U25570 ( .A(n23831), .B(n23380), .Z(n23382) );
  XOR U25571 ( .A(n23832), .B(n23833), .Z(n23380) );
  AND U25572 ( .A(n23834), .B(n23835), .Z(n23832) );
  AND U25573 ( .A(a[5]), .B(b[58]), .Z(n23831) );
  XOR U25574 ( .A(n23836), .B(n23385), .Z(n23387) );
  XOR U25575 ( .A(n23837), .B(n23838), .Z(n23385) );
  AND U25576 ( .A(n23839), .B(n23840), .Z(n23837) );
  AND U25577 ( .A(a[6]), .B(b[57]), .Z(n23836) );
  XOR U25578 ( .A(n23841), .B(n23390), .Z(n23392) );
  XOR U25579 ( .A(n23842), .B(n23843), .Z(n23390) );
  AND U25580 ( .A(n23844), .B(n23845), .Z(n23842) );
  AND U25581 ( .A(a[7]), .B(b[56]), .Z(n23841) );
  XOR U25582 ( .A(n23846), .B(n23395), .Z(n23397) );
  XOR U25583 ( .A(n23847), .B(n23848), .Z(n23395) );
  AND U25584 ( .A(n23849), .B(n23850), .Z(n23847) );
  AND U25585 ( .A(a[8]), .B(b[55]), .Z(n23846) );
  XOR U25586 ( .A(n23851), .B(n23400), .Z(n23402) );
  XOR U25587 ( .A(n23852), .B(n23853), .Z(n23400) );
  AND U25588 ( .A(n23854), .B(n23855), .Z(n23852) );
  AND U25589 ( .A(a[9]), .B(b[54]), .Z(n23851) );
  XOR U25590 ( .A(n23856), .B(n23405), .Z(n23407) );
  XOR U25591 ( .A(n23857), .B(n23858), .Z(n23405) );
  AND U25592 ( .A(n23859), .B(n23860), .Z(n23857) );
  AND U25593 ( .A(a[10]), .B(b[53]), .Z(n23856) );
  XOR U25594 ( .A(n23861), .B(n23410), .Z(n23412) );
  XOR U25595 ( .A(n23862), .B(n23863), .Z(n23410) );
  AND U25596 ( .A(n23864), .B(n23865), .Z(n23862) );
  AND U25597 ( .A(a[11]), .B(b[52]), .Z(n23861) );
  XOR U25598 ( .A(n23866), .B(n23415), .Z(n23417) );
  XOR U25599 ( .A(n23867), .B(n23868), .Z(n23415) );
  AND U25600 ( .A(n23869), .B(n23870), .Z(n23867) );
  AND U25601 ( .A(a[12]), .B(b[51]), .Z(n23866) );
  XOR U25602 ( .A(n23871), .B(n23420), .Z(n23422) );
  XOR U25603 ( .A(n23872), .B(n23873), .Z(n23420) );
  AND U25604 ( .A(n23874), .B(n23875), .Z(n23872) );
  AND U25605 ( .A(a[13]), .B(b[50]), .Z(n23871) );
  XOR U25606 ( .A(n23876), .B(n23425), .Z(n23427) );
  XOR U25607 ( .A(n23877), .B(n23878), .Z(n23425) );
  AND U25608 ( .A(n23879), .B(n23880), .Z(n23877) );
  AND U25609 ( .A(a[14]), .B(b[49]), .Z(n23876) );
  XOR U25610 ( .A(n23881), .B(n23430), .Z(n23432) );
  XOR U25611 ( .A(n23882), .B(n23883), .Z(n23430) );
  AND U25612 ( .A(n23884), .B(n23885), .Z(n23882) );
  AND U25613 ( .A(a[15]), .B(b[48]), .Z(n23881) );
  XOR U25614 ( .A(n23886), .B(n23435), .Z(n23437) );
  XOR U25615 ( .A(n23887), .B(n23888), .Z(n23435) );
  AND U25616 ( .A(n23889), .B(n23890), .Z(n23887) );
  AND U25617 ( .A(a[16]), .B(b[47]), .Z(n23886) );
  XOR U25618 ( .A(n23891), .B(n23440), .Z(n23442) );
  XOR U25619 ( .A(n23892), .B(n23893), .Z(n23440) );
  AND U25620 ( .A(n23894), .B(n23895), .Z(n23892) );
  AND U25621 ( .A(a[17]), .B(b[46]), .Z(n23891) );
  XOR U25622 ( .A(n23896), .B(n23445), .Z(n23447) );
  XOR U25623 ( .A(n23897), .B(n23898), .Z(n23445) );
  AND U25624 ( .A(n23899), .B(n23900), .Z(n23897) );
  AND U25625 ( .A(a[18]), .B(b[45]), .Z(n23896) );
  XOR U25626 ( .A(n23901), .B(n23450), .Z(n23452) );
  XOR U25627 ( .A(n23902), .B(n23903), .Z(n23450) );
  AND U25628 ( .A(n23904), .B(n23905), .Z(n23902) );
  AND U25629 ( .A(a[19]), .B(b[44]), .Z(n23901) );
  XOR U25630 ( .A(n23906), .B(n23455), .Z(n23457) );
  XOR U25631 ( .A(n23907), .B(n23908), .Z(n23455) );
  AND U25632 ( .A(n23909), .B(n23910), .Z(n23907) );
  AND U25633 ( .A(a[20]), .B(b[43]), .Z(n23906) );
  XOR U25634 ( .A(n23911), .B(n23460), .Z(n23462) );
  XOR U25635 ( .A(n23912), .B(n23913), .Z(n23460) );
  AND U25636 ( .A(n23914), .B(n23915), .Z(n23912) );
  AND U25637 ( .A(a[21]), .B(b[42]), .Z(n23911) );
  XOR U25638 ( .A(n23916), .B(n23465), .Z(n23467) );
  XOR U25639 ( .A(n23917), .B(n23918), .Z(n23465) );
  AND U25640 ( .A(n23919), .B(n23920), .Z(n23917) );
  AND U25641 ( .A(a[22]), .B(b[41]), .Z(n23916) );
  XOR U25642 ( .A(n23921), .B(n23470), .Z(n23472) );
  XOR U25643 ( .A(n23922), .B(n23923), .Z(n23470) );
  AND U25644 ( .A(n23924), .B(n23925), .Z(n23922) );
  AND U25645 ( .A(a[23]), .B(b[40]), .Z(n23921) );
  XOR U25646 ( .A(n23926), .B(n23475), .Z(n23477) );
  XOR U25647 ( .A(n23927), .B(n23928), .Z(n23475) );
  AND U25648 ( .A(n23929), .B(n23930), .Z(n23927) );
  AND U25649 ( .A(a[24]), .B(b[39]), .Z(n23926) );
  XOR U25650 ( .A(n23931), .B(n23480), .Z(n23482) );
  XOR U25651 ( .A(n23932), .B(n23933), .Z(n23480) );
  AND U25652 ( .A(n23934), .B(n23935), .Z(n23932) );
  AND U25653 ( .A(a[25]), .B(b[38]), .Z(n23931) );
  XOR U25654 ( .A(n23936), .B(n23485), .Z(n23487) );
  XOR U25655 ( .A(n23937), .B(n23938), .Z(n23485) );
  AND U25656 ( .A(n23939), .B(n23940), .Z(n23937) );
  AND U25657 ( .A(a[26]), .B(b[37]), .Z(n23936) );
  XOR U25658 ( .A(n23941), .B(n23490), .Z(n23492) );
  XOR U25659 ( .A(n23942), .B(n23943), .Z(n23490) );
  AND U25660 ( .A(n23944), .B(n23945), .Z(n23942) );
  AND U25661 ( .A(a[27]), .B(b[36]), .Z(n23941) );
  XOR U25662 ( .A(n23946), .B(n23495), .Z(n23497) );
  XOR U25663 ( .A(n23947), .B(n23948), .Z(n23495) );
  AND U25664 ( .A(n23949), .B(n23950), .Z(n23947) );
  AND U25665 ( .A(a[28]), .B(b[35]), .Z(n23946) );
  XOR U25666 ( .A(n23951), .B(n23500), .Z(n23502) );
  XOR U25667 ( .A(n23952), .B(n23953), .Z(n23500) );
  AND U25668 ( .A(n23954), .B(n23955), .Z(n23952) );
  AND U25669 ( .A(a[29]), .B(b[34]), .Z(n23951) );
  XOR U25670 ( .A(n23956), .B(n23505), .Z(n23507) );
  XOR U25671 ( .A(n23957), .B(n23958), .Z(n23505) );
  AND U25672 ( .A(n23959), .B(n23960), .Z(n23957) );
  AND U25673 ( .A(a[30]), .B(b[33]), .Z(n23956) );
  XOR U25674 ( .A(n23961), .B(n23510), .Z(n23512) );
  XOR U25675 ( .A(n23962), .B(n23963), .Z(n23510) );
  AND U25676 ( .A(n23964), .B(n23965), .Z(n23962) );
  AND U25677 ( .A(a[31]), .B(b[32]), .Z(n23961) );
  XOR U25678 ( .A(n23966), .B(n23515), .Z(n23517) );
  XOR U25679 ( .A(n23967), .B(n23968), .Z(n23515) );
  AND U25680 ( .A(n23969), .B(n23970), .Z(n23967) );
  AND U25681 ( .A(b[31]), .B(a[32]), .Z(n23966) );
  XOR U25682 ( .A(n23971), .B(n23520), .Z(n23522) );
  XOR U25683 ( .A(n23972), .B(n23973), .Z(n23520) );
  AND U25684 ( .A(n23974), .B(n23975), .Z(n23972) );
  AND U25685 ( .A(b[30]), .B(a[33]), .Z(n23971) );
  XOR U25686 ( .A(n23976), .B(n23525), .Z(n23527) );
  XOR U25687 ( .A(n23977), .B(n23978), .Z(n23525) );
  AND U25688 ( .A(n23979), .B(n23980), .Z(n23977) );
  AND U25689 ( .A(b[29]), .B(a[34]), .Z(n23976) );
  XOR U25690 ( .A(n23981), .B(n23534), .Z(n23536) );
  XOR U25691 ( .A(n23982), .B(n23983), .Z(n23534) );
  AND U25692 ( .A(n23984), .B(n23985), .Z(n23982) );
  AND U25693 ( .A(b[28]), .B(a[35]), .Z(n23981) );
  XOR U25694 ( .A(n23986), .B(n23529), .Z(n23531) );
  XOR U25695 ( .A(n23987), .B(n23988), .Z(n23529) );
  AND U25696 ( .A(n23989), .B(n23990), .Z(n23987) );
  AND U25697 ( .A(b[27]), .B(a[36]), .Z(n23986) );
  XOR U25698 ( .A(n23991), .B(n23539), .Z(n23541) );
  XOR U25699 ( .A(n23992), .B(n23993), .Z(n23539) );
  AND U25700 ( .A(n23994), .B(n23995), .Z(n23992) );
  AND U25701 ( .A(b[26]), .B(a[37]), .Z(n23991) );
  XOR U25702 ( .A(n23996), .B(n23544), .Z(n23546) );
  XOR U25703 ( .A(n23997), .B(n23998), .Z(n23544) );
  AND U25704 ( .A(n23999), .B(n24000), .Z(n23997) );
  AND U25705 ( .A(b[25]), .B(a[38]), .Z(n23996) );
  XOR U25706 ( .A(n24001), .B(n23549), .Z(n23551) );
  XOR U25707 ( .A(n24002), .B(n24003), .Z(n23549) );
  AND U25708 ( .A(n24004), .B(n24005), .Z(n24002) );
  AND U25709 ( .A(b[24]), .B(a[39]), .Z(n24001) );
  XOR U25710 ( .A(n24006), .B(n23554), .Z(n23556) );
  XOR U25711 ( .A(n24007), .B(n24008), .Z(n23554) );
  AND U25712 ( .A(n24009), .B(n24010), .Z(n24007) );
  AND U25713 ( .A(b[23]), .B(a[40]), .Z(n24006) );
  XOR U25714 ( .A(n24011), .B(n23559), .Z(n23561) );
  XOR U25715 ( .A(n24012), .B(n24013), .Z(n23559) );
  AND U25716 ( .A(n24014), .B(n24015), .Z(n24012) );
  AND U25717 ( .A(b[22]), .B(a[41]), .Z(n24011) );
  XOR U25718 ( .A(n24016), .B(n23564), .Z(n23566) );
  XOR U25719 ( .A(n24017), .B(n24018), .Z(n23564) );
  AND U25720 ( .A(n24019), .B(n24020), .Z(n24017) );
  AND U25721 ( .A(b[21]), .B(a[42]), .Z(n24016) );
  XOR U25722 ( .A(n24021), .B(n23569), .Z(n23571) );
  XOR U25723 ( .A(n24022), .B(n24023), .Z(n23569) );
  AND U25724 ( .A(n24024), .B(n24025), .Z(n24022) );
  AND U25725 ( .A(b[20]), .B(a[43]), .Z(n24021) );
  XOR U25726 ( .A(n24026), .B(n23574), .Z(n23576) );
  XOR U25727 ( .A(n24027), .B(n24028), .Z(n23574) );
  AND U25728 ( .A(n24029), .B(n24030), .Z(n24027) );
  AND U25729 ( .A(b[19]), .B(a[44]), .Z(n24026) );
  XOR U25730 ( .A(n24031), .B(n23579), .Z(n23581) );
  XOR U25731 ( .A(n24032), .B(n24033), .Z(n23579) );
  AND U25732 ( .A(n24034), .B(n24035), .Z(n24032) );
  AND U25733 ( .A(b[18]), .B(a[45]), .Z(n24031) );
  XOR U25734 ( .A(n24036), .B(n23584), .Z(n23586) );
  XOR U25735 ( .A(n24037), .B(n24038), .Z(n23584) );
  AND U25736 ( .A(n24039), .B(n24040), .Z(n24037) );
  AND U25737 ( .A(b[17]), .B(a[46]), .Z(n24036) );
  XOR U25738 ( .A(n24041), .B(n23589), .Z(n23591) );
  XOR U25739 ( .A(n24042), .B(n24043), .Z(n23589) );
  AND U25740 ( .A(n24044), .B(n24045), .Z(n24042) );
  AND U25741 ( .A(b[16]), .B(a[47]), .Z(n24041) );
  XOR U25742 ( .A(n24046), .B(n23594), .Z(n23596) );
  XOR U25743 ( .A(n24047), .B(n24048), .Z(n23594) );
  AND U25744 ( .A(n24049), .B(n24050), .Z(n24047) );
  AND U25745 ( .A(b[15]), .B(a[48]), .Z(n24046) );
  XOR U25746 ( .A(n24051), .B(n23599), .Z(n23601) );
  XOR U25747 ( .A(n24052), .B(n24053), .Z(n23599) );
  AND U25748 ( .A(n24054), .B(n24055), .Z(n24052) );
  AND U25749 ( .A(b[14]), .B(a[49]), .Z(n24051) );
  XOR U25750 ( .A(n24056), .B(n23604), .Z(n23606) );
  XOR U25751 ( .A(n24057), .B(n24058), .Z(n23604) );
  AND U25752 ( .A(n24059), .B(n24060), .Z(n24057) );
  AND U25753 ( .A(b[13]), .B(a[50]), .Z(n24056) );
  XOR U25754 ( .A(n24061), .B(n23609), .Z(n23611) );
  XOR U25755 ( .A(n24062), .B(n24063), .Z(n23609) );
  AND U25756 ( .A(n24064), .B(n24065), .Z(n24062) );
  AND U25757 ( .A(b[12]), .B(a[51]), .Z(n24061) );
  XOR U25758 ( .A(n24066), .B(n23614), .Z(n23616) );
  XOR U25759 ( .A(n24067), .B(n24068), .Z(n23614) );
  AND U25760 ( .A(n24069), .B(n24070), .Z(n24067) );
  AND U25761 ( .A(b[11]), .B(a[52]), .Z(n24066) );
  XOR U25762 ( .A(n24071), .B(n23619), .Z(n23621) );
  XOR U25763 ( .A(n24072), .B(n24073), .Z(n23619) );
  AND U25764 ( .A(n24074), .B(n24075), .Z(n24072) );
  AND U25765 ( .A(b[10]), .B(a[53]), .Z(n24071) );
  XOR U25766 ( .A(n24076), .B(n23624), .Z(n23626) );
  XOR U25767 ( .A(n24077), .B(n24078), .Z(n23624) );
  AND U25768 ( .A(n24079), .B(n24080), .Z(n24077) );
  AND U25769 ( .A(b[9]), .B(a[54]), .Z(n24076) );
  XOR U25770 ( .A(n24081), .B(n23629), .Z(n23631) );
  XOR U25771 ( .A(n24082), .B(n24083), .Z(n23629) );
  AND U25772 ( .A(n24084), .B(n24085), .Z(n24082) );
  AND U25773 ( .A(b[8]), .B(a[55]), .Z(n24081) );
  XOR U25774 ( .A(n24086), .B(n23634), .Z(n23636) );
  XOR U25775 ( .A(n24087), .B(n24088), .Z(n23634) );
  AND U25776 ( .A(n24089), .B(n24090), .Z(n24087) );
  AND U25777 ( .A(b[7]), .B(a[56]), .Z(n24086) );
  XOR U25778 ( .A(n24091), .B(n23639), .Z(n23641) );
  XOR U25779 ( .A(n24092), .B(n24093), .Z(n23639) );
  AND U25780 ( .A(n24094), .B(n24095), .Z(n24092) );
  AND U25781 ( .A(b[6]), .B(a[57]), .Z(n24091) );
  XOR U25782 ( .A(n24096), .B(n23644), .Z(n23646) );
  XOR U25783 ( .A(n24097), .B(n24098), .Z(n23644) );
  AND U25784 ( .A(n24099), .B(n24100), .Z(n24097) );
  AND U25785 ( .A(b[5]), .B(a[58]), .Z(n24096) );
  XOR U25786 ( .A(n24101), .B(n23649), .Z(n23651) );
  XOR U25787 ( .A(n24102), .B(n24103), .Z(n23649) );
  AND U25788 ( .A(n24104), .B(n24105), .Z(n24102) );
  AND U25789 ( .A(b[4]), .B(a[59]), .Z(n24101) );
  XNOR U25790 ( .A(n24106), .B(n24107), .Z(n23659) );
  NANDN U25791 ( .A(n24108), .B(n24109), .Z(n24107) );
  XOR U25792 ( .A(n24110), .B(n23654), .Z(n23656) );
  XNOR U25793 ( .A(n24111), .B(n24112), .Z(n23654) );
  AND U25794 ( .A(n24113), .B(n24114), .Z(n24111) );
  AND U25795 ( .A(b[3]), .B(a[60]), .Z(n24110) );
  XOR U25796 ( .A(n23745), .B(n23744), .Z(c[126]) );
  XOR U25797 ( .A(sreg[190]), .B(n23743), .Z(n23744) );
  XOR U25798 ( .A(n23749), .B(n24115), .Z(n23745) );
  XNOR U25799 ( .A(n23750), .B(n23743), .Z(n24115) );
  XOR U25800 ( .A(n24116), .B(n24117), .Z(n23743) );
  NOR U25801 ( .A(n24118), .B(n24119), .Z(n24116) );
  NAND U25802 ( .A(a[62]), .B(b[0]), .Z(n23750) );
  XNOR U25803 ( .A(n24108), .B(n24109), .Z(n23749) );
  XOR U25804 ( .A(n24106), .B(n24120), .Z(n24109) );
  NAND U25805 ( .A(b[1]), .B(a[61]), .Z(n24120) );
  XOR U25806 ( .A(n24114), .B(n24121), .Z(n24108) );
  XOR U25807 ( .A(n24106), .B(n24113), .Z(n24121) );
  XNOR U25808 ( .A(n24122), .B(n24112), .Z(n24113) );
  AND U25809 ( .A(b[2]), .B(a[60]), .Z(n24122) );
  NANDN U25810 ( .A(n24123), .B(n24124), .Z(n24106) );
  XOR U25811 ( .A(n24112), .B(n24104), .Z(n24125) );
  XNOR U25812 ( .A(n24103), .B(n24099), .Z(n24126) );
  XNOR U25813 ( .A(n24098), .B(n24094), .Z(n24127) );
  XNOR U25814 ( .A(n24093), .B(n24089), .Z(n24128) );
  XNOR U25815 ( .A(n24088), .B(n24084), .Z(n24129) );
  XNOR U25816 ( .A(n24083), .B(n24079), .Z(n24130) );
  XNOR U25817 ( .A(n24078), .B(n24074), .Z(n24131) );
  XNOR U25818 ( .A(n24073), .B(n24069), .Z(n24132) );
  XNOR U25819 ( .A(n24068), .B(n24064), .Z(n24133) );
  XNOR U25820 ( .A(n24063), .B(n24059), .Z(n24134) );
  XNOR U25821 ( .A(n24058), .B(n24054), .Z(n24135) );
  XNOR U25822 ( .A(n24053), .B(n24049), .Z(n24136) );
  XNOR U25823 ( .A(n24048), .B(n24044), .Z(n24137) );
  XNOR U25824 ( .A(n24043), .B(n24039), .Z(n24138) );
  XNOR U25825 ( .A(n24038), .B(n24034), .Z(n24139) );
  XNOR U25826 ( .A(n24033), .B(n24029), .Z(n24140) );
  XNOR U25827 ( .A(n24028), .B(n24024), .Z(n24141) );
  XNOR U25828 ( .A(n24023), .B(n24019), .Z(n24142) );
  XNOR U25829 ( .A(n24018), .B(n24014), .Z(n24143) );
  XNOR U25830 ( .A(n24013), .B(n24009), .Z(n24144) );
  XNOR U25831 ( .A(n24008), .B(n24004), .Z(n24145) );
  XNOR U25832 ( .A(n24003), .B(n23999), .Z(n24146) );
  XNOR U25833 ( .A(n23998), .B(n23994), .Z(n24147) );
  XNOR U25834 ( .A(n23993), .B(n23989), .Z(n24148) );
  XNOR U25835 ( .A(n23988), .B(n23984), .Z(n24149) );
  XNOR U25836 ( .A(n23983), .B(n23979), .Z(n24150) );
  XNOR U25837 ( .A(n23978), .B(n23974), .Z(n24151) );
  XNOR U25838 ( .A(n23973), .B(n23969), .Z(n24152) );
  XNOR U25839 ( .A(n23968), .B(n23964), .Z(n24153) );
  XNOR U25840 ( .A(n23963), .B(n23959), .Z(n24154) );
  XNOR U25841 ( .A(n23958), .B(n23954), .Z(n24155) );
  XNOR U25842 ( .A(n23953), .B(n23949), .Z(n24156) );
  XNOR U25843 ( .A(n23948), .B(n23944), .Z(n24157) );
  XNOR U25844 ( .A(n23943), .B(n23939), .Z(n24158) );
  XNOR U25845 ( .A(n23938), .B(n23934), .Z(n24159) );
  XNOR U25846 ( .A(n23933), .B(n23929), .Z(n24160) );
  XNOR U25847 ( .A(n23928), .B(n23924), .Z(n24161) );
  XNOR U25848 ( .A(n23923), .B(n23919), .Z(n24162) );
  XNOR U25849 ( .A(n23918), .B(n23914), .Z(n24163) );
  XNOR U25850 ( .A(n23913), .B(n23909), .Z(n24164) );
  XNOR U25851 ( .A(n23908), .B(n23904), .Z(n24165) );
  XNOR U25852 ( .A(n23903), .B(n23899), .Z(n24166) );
  XNOR U25853 ( .A(n23898), .B(n23894), .Z(n24167) );
  XNOR U25854 ( .A(n23893), .B(n23889), .Z(n24168) );
  XNOR U25855 ( .A(n23888), .B(n23884), .Z(n24169) );
  XNOR U25856 ( .A(n23883), .B(n23879), .Z(n24170) );
  XNOR U25857 ( .A(n23878), .B(n23874), .Z(n24171) );
  XNOR U25858 ( .A(n23873), .B(n23869), .Z(n24172) );
  XNOR U25859 ( .A(n23868), .B(n23864), .Z(n24173) );
  XNOR U25860 ( .A(n23863), .B(n23859), .Z(n24174) );
  XNOR U25861 ( .A(n23858), .B(n23854), .Z(n24175) );
  XNOR U25862 ( .A(n23853), .B(n23849), .Z(n24176) );
  XNOR U25863 ( .A(n23848), .B(n23844), .Z(n24177) );
  XNOR U25864 ( .A(n23843), .B(n23839), .Z(n24178) );
  XNOR U25865 ( .A(n23838), .B(n23834), .Z(n24179) );
  XNOR U25866 ( .A(n23833), .B(n23829), .Z(n24180) );
  XNOR U25867 ( .A(n23828), .B(n23824), .Z(n24181) );
  XOR U25868 ( .A(n23823), .B(n23820), .Z(n24182) );
  XOR U25869 ( .A(n24183), .B(n24184), .Z(n23820) );
  XOR U25870 ( .A(n23818), .B(n24185), .Z(n24184) );
  XOR U25871 ( .A(n24186), .B(n24187), .Z(n24185) );
  AND U25872 ( .A(a[0]), .B(b[62]), .Z(n24186) );
  XNOR U25873 ( .A(n24188), .B(n24187), .Z(n24183) );
  XNOR U25874 ( .A(n24189), .B(n24190), .Z(n24187) );
  AND U25875 ( .A(n24191), .B(n24192), .Z(n24189) );
  AND U25876 ( .A(a[1]), .B(b[61]), .Z(n24188) );
  XOR U25877 ( .A(n24193), .B(n23818), .Z(n23819) );
  XOR U25878 ( .A(n24194), .B(n24195), .Z(n23818) );
  AND U25879 ( .A(n24196), .B(n24197), .Z(n24194) );
  AND U25880 ( .A(a[2]), .B(b[60]), .Z(n24193) );
  XOR U25881 ( .A(n24198), .B(n23823), .Z(n23825) );
  XOR U25882 ( .A(n24199), .B(n24200), .Z(n23823) );
  AND U25883 ( .A(n24201), .B(n24202), .Z(n24199) );
  AND U25884 ( .A(a[3]), .B(b[59]), .Z(n24198) );
  XOR U25885 ( .A(n24203), .B(n23828), .Z(n23830) );
  XOR U25886 ( .A(n24204), .B(n24205), .Z(n23828) );
  AND U25887 ( .A(n24206), .B(n24207), .Z(n24204) );
  AND U25888 ( .A(a[4]), .B(b[58]), .Z(n24203) );
  XOR U25889 ( .A(n24208), .B(n23833), .Z(n23835) );
  XOR U25890 ( .A(n24209), .B(n24210), .Z(n23833) );
  AND U25891 ( .A(n24211), .B(n24212), .Z(n24209) );
  AND U25892 ( .A(a[5]), .B(b[57]), .Z(n24208) );
  XOR U25893 ( .A(n24213), .B(n23838), .Z(n23840) );
  XOR U25894 ( .A(n24214), .B(n24215), .Z(n23838) );
  AND U25895 ( .A(n24216), .B(n24217), .Z(n24214) );
  AND U25896 ( .A(a[6]), .B(b[56]), .Z(n24213) );
  XOR U25897 ( .A(n24218), .B(n23843), .Z(n23845) );
  XOR U25898 ( .A(n24219), .B(n24220), .Z(n23843) );
  AND U25899 ( .A(n24221), .B(n24222), .Z(n24219) );
  AND U25900 ( .A(a[7]), .B(b[55]), .Z(n24218) );
  XOR U25901 ( .A(n24223), .B(n23848), .Z(n23850) );
  XOR U25902 ( .A(n24224), .B(n24225), .Z(n23848) );
  AND U25903 ( .A(n24226), .B(n24227), .Z(n24224) );
  AND U25904 ( .A(a[8]), .B(b[54]), .Z(n24223) );
  XOR U25905 ( .A(n24228), .B(n23853), .Z(n23855) );
  XOR U25906 ( .A(n24229), .B(n24230), .Z(n23853) );
  AND U25907 ( .A(n24231), .B(n24232), .Z(n24229) );
  AND U25908 ( .A(a[9]), .B(b[53]), .Z(n24228) );
  XOR U25909 ( .A(n24233), .B(n23858), .Z(n23860) );
  XOR U25910 ( .A(n24234), .B(n24235), .Z(n23858) );
  AND U25911 ( .A(n24236), .B(n24237), .Z(n24234) );
  AND U25912 ( .A(a[10]), .B(b[52]), .Z(n24233) );
  XOR U25913 ( .A(n24238), .B(n23863), .Z(n23865) );
  XOR U25914 ( .A(n24239), .B(n24240), .Z(n23863) );
  AND U25915 ( .A(n24241), .B(n24242), .Z(n24239) );
  AND U25916 ( .A(a[11]), .B(b[51]), .Z(n24238) );
  XOR U25917 ( .A(n24243), .B(n23868), .Z(n23870) );
  XOR U25918 ( .A(n24244), .B(n24245), .Z(n23868) );
  AND U25919 ( .A(n24246), .B(n24247), .Z(n24244) );
  AND U25920 ( .A(a[12]), .B(b[50]), .Z(n24243) );
  XOR U25921 ( .A(n24248), .B(n23873), .Z(n23875) );
  XOR U25922 ( .A(n24249), .B(n24250), .Z(n23873) );
  AND U25923 ( .A(n24251), .B(n24252), .Z(n24249) );
  AND U25924 ( .A(a[13]), .B(b[49]), .Z(n24248) );
  XOR U25925 ( .A(n24253), .B(n23878), .Z(n23880) );
  XOR U25926 ( .A(n24254), .B(n24255), .Z(n23878) );
  AND U25927 ( .A(n24256), .B(n24257), .Z(n24254) );
  AND U25928 ( .A(a[14]), .B(b[48]), .Z(n24253) );
  XOR U25929 ( .A(n24258), .B(n23883), .Z(n23885) );
  XOR U25930 ( .A(n24259), .B(n24260), .Z(n23883) );
  AND U25931 ( .A(n24261), .B(n24262), .Z(n24259) );
  AND U25932 ( .A(a[15]), .B(b[47]), .Z(n24258) );
  XOR U25933 ( .A(n24263), .B(n23888), .Z(n23890) );
  XOR U25934 ( .A(n24264), .B(n24265), .Z(n23888) );
  AND U25935 ( .A(n24266), .B(n24267), .Z(n24264) );
  AND U25936 ( .A(a[16]), .B(b[46]), .Z(n24263) );
  XOR U25937 ( .A(n24268), .B(n23893), .Z(n23895) );
  XOR U25938 ( .A(n24269), .B(n24270), .Z(n23893) );
  AND U25939 ( .A(n24271), .B(n24272), .Z(n24269) );
  AND U25940 ( .A(a[17]), .B(b[45]), .Z(n24268) );
  XOR U25941 ( .A(n24273), .B(n23898), .Z(n23900) );
  XOR U25942 ( .A(n24274), .B(n24275), .Z(n23898) );
  AND U25943 ( .A(n24276), .B(n24277), .Z(n24274) );
  AND U25944 ( .A(a[18]), .B(b[44]), .Z(n24273) );
  XOR U25945 ( .A(n24278), .B(n23903), .Z(n23905) );
  XOR U25946 ( .A(n24279), .B(n24280), .Z(n23903) );
  AND U25947 ( .A(n24281), .B(n24282), .Z(n24279) );
  AND U25948 ( .A(a[19]), .B(b[43]), .Z(n24278) );
  XOR U25949 ( .A(n24283), .B(n23908), .Z(n23910) );
  XOR U25950 ( .A(n24284), .B(n24285), .Z(n23908) );
  AND U25951 ( .A(n24286), .B(n24287), .Z(n24284) );
  AND U25952 ( .A(a[20]), .B(b[42]), .Z(n24283) );
  XOR U25953 ( .A(n24288), .B(n23913), .Z(n23915) );
  XOR U25954 ( .A(n24289), .B(n24290), .Z(n23913) );
  AND U25955 ( .A(n24291), .B(n24292), .Z(n24289) );
  AND U25956 ( .A(a[21]), .B(b[41]), .Z(n24288) );
  XOR U25957 ( .A(n24293), .B(n23918), .Z(n23920) );
  XOR U25958 ( .A(n24294), .B(n24295), .Z(n23918) );
  AND U25959 ( .A(n24296), .B(n24297), .Z(n24294) );
  AND U25960 ( .A(a[22]), .B(b[40]), .Z(n24293) );
  XOR U25961 ( .A(n24298), .B(n23923), .Z(n23925) );
  XOR U25962 ( .A(n24299), .B(n24300), .Z(n23923) );
  AND U25963 ( .A(n24301), .B(n24302), .Z(n24299) );
  AND U25964 ( .A(a[23]), .B(b[39]), .Z(n24298) );
  XOR U25965 ( .A(n24303), .B(n23928), .Z(n23930) );
  XOR U25966 ( .A(n24304), .B(n24305), .Z(n23928) );
  AND U25967 ( .A(n24306), .B(n24307), .Z(n24304) );
  AND U25968 ( .A(a[24]), .B(b[38]), .Z(n24303) );
  XOR U25969 ( .A(n24308), .B(n23933), .Z(n23935) );
  XOR U25970 ( .A(n24309), .B(n24310), .Z(n23933) );
  AND U25971 ( .A(n24311), .B(n24312), .Z(n24309) );
  AND U25972 ( .A(a[25]), .B(b[37]), .Z(n24308) );
  XOR U25973 ( .A(n24313), .B(n23938), .Z(n23940) );
  XOR U25974 ( .A(n24314), .B(n24315), .Z(n23938) );
  AND U25975 ( .A(n24316), .B(n24317), .Z(n24314) );
  AND U25976 ( .A(a[26]), .B(b[36]), .Z(n24313) );
  XOR U25977 ( .A(n24318), .B(n23943), .Z(n23945) );
  XOR U25978 ( .A(n24319), .B(n24320), .Z(n23943) );
  AND U25979 ( .A(n24321), .B(n24322), .Z(n24319) );
  AND U25980 ( .A(a[27]), .B(b[35]), .Z(n24318) );
  XOR U25981 ( .A(n24323), .B(n23948), .Z(n23950) );
  XOR U25982 ( .A(n24324), .B(n24325), .Z(n23948) );
  AND U25983 ( .A(n24326), .B(n24327), .Z(n24324) );
  AND U25984 ( .A(a[28]), .B(b[34]), .Z(n24323) );
  XOR U25985 ( .A(n24328), .B(n23953), .Z(n23955) );
  XOR U25986 ( .A(n24329), .B(n24330), .Z(n23953) );
  AND U25987 ( .A(n24331), .B(n24332), .Z(n24329) );
  AND U25988 ( .A(a[29]), .B(b[33]), .Z(n24328) );
  XOR U25989 ( .A(n24333), .B(n23958), .Z(n23960) );
  XOR U25990 ( .A(n24334), .B(n24335), .Z(n23958) );
  AND U25991 ( .A(n24336), .B(n24337), .Z(n24334) );
  AND U25992 ( .A(a[30]), .B(b[32]), .Z(n24333) );
  XOR U25993 ( .A(n24338), .B(n23963), .Z(n23965) );
  XOR U25994 ( .A(n24339), .B(n24340), .Z(n23963) );
  AND U25995 ( .A(n24341), .B(n24342), .Z(n24339) );
  AND U25996 ( .A(a[31]), .B(b[31]), .Z(n24338) );
  XOR U25997 ( .A(n24343), .B(n23968), .Z(n23970) );
  XOR U25998 ( .A(n24344), .B(n24345), .Z(n23968) );
  AND U25999 ( .A(n24346), .B(n24347), .Z(n24344) );
  AND U26000 ( .A(b[30]), .B(a[32]), .Z(n24343) );
  XOR U26001 ( .A(n24348), .B(n23973), .Z(n23975) );
  XOR U26002 ( .A(n24349), .B(n24350), .Z(n23973) );
  AND U26003 ( .A(n24351), .B(n24352), .Z(n24349) );
  AND U26004 ( .A(b[29]), .B(a[33]), .Z(n24348) );
  XOR U26005 ( .A(n24353), .B(n23978), .Z(n23980) );
  XOR U26006 ( .A(n24354), .B(n24355), .Z(n23978) );
  AND U26007 ( .A(n24356), .B(n24357), .Z(n24354) );
  AND U26008 ( .A(b[28]), .B(a[34]), .Z(n24353) );
  XOR U26009 ( .A(n24358), .B(n23983), .Z(n23985) );
  XOR U26010 ( .A(n24359), .B(n24360), .Z(n23983) );
  AND U26011 ( .A(n24361), .B(n24362), .Z(n24359) );
  AND U26012 ( .A(b[27]), .B(a[35]), .Z(n24358) );
  XOR U26013 ( .A(n24363), .B(n23988), .Z(n23990) );
  XOR U26014 ( .A(n24364), .B(n24365), .Z(n23988) );
  AND U26015 ( .A(n24366), .B(n24367), .Z(n24364) );
  AND U26016 ( .A(b[26]), .B(a[36]), .Z(n24363) );
  XOR U26017 ( .A(n24368), .B(n23993), .Z(n23995) );
  XOR U26018 ( .A(n24369), .B(n24370), .Z(n23993) );
  AND U26019 ( .A(n24371), .B(n24372), .Z(n24369) );
  AND U26020 ( .A(b[25]), .B(a[37]), .Z(n24368) );
  XOR U26021 ( .A(n24373), .B(n23998), .Z(n24000) );
  XOR U26022 ( .A(n24374), .B(n24375), .Z(n23998) );
  AND U26023 ( .A(n24376), .B(n24377), .Z(n24374) );
  AND U26024 ( .A(b[24]), .B(a[38]), .Z(n24373) );
  XOR U26025 ( .A(n24378), .B(n24003), .Z(n24005) );
  XOR U26026 ( .A(n24379), .B(n24380), .Z(n24003) );
  AND U26027 ( .A(n24381), .B(n24382), .Z(n24379) );
  AND U26028 ( .A(b[23]), .B(a[39]), .Z(n24378) );
  XOR U26029 ( .A(n24383), .B(n24008), .Z(n24010) );
  XOR U26030 ( .A(n24384), .B(n24385), .Z(n24008) );
  AND U26031 ( .A(n24386), .B(n24387), .Z(n24384) );
  AND U26032 ( .A(b[22]), .B(a[40]), .Z(n24383) );
  XOR U26033 ( .A(n24388), .B(n24013), .Z(n24015) );
  XOR U26034 ( .A(n24389), .B(n24390), .Z(n24013) );
  AND U26035 ( .A(n24391), .B(n24392), .Z(n24389) );
  AND U26036 ( .A(b[21]), .B(a[41]), .Z(n24388) );
  XOR U26037 ( .A(n24393), .B(n24018), .Z(n24020) );
  XOR U26038 ( .A(n24394), .B(n24395), .Z(n24018) );
  AND U26039 ( .A(n24396), .B(n24397), .Z(n24394) );
  AND U26040 ( .A(b[20]), .B(a[42]), .Z(n24393) );
  XOR U26041 ( .A(n24398), .B(n24023), .Z(n24025) );
  XOR U26042 ( .A(n24399), .B(n24400), .Z(n24023) );
  AND U26043 ( .A(n24401), .B(n24402), .Z(n24399) );
  AND U26044 ( .A(b[19]), .B(a[43]), .Z(n24398) );
  XOR U26045 ( .A(n24403), .B(n24028), .Z(n24030) );
  XOR U26046 ( .A(n24404), .B(n24405), .Z(n24028) );
  AND U26047 ( .A(n24406), .B(n24407), .Z(n24404) );
  AND U26048 ( .A(b[18]), .B(a[44]), .Z(n24403) );
  XOR U26049 ( .A(n24408), .B(n24033), .Z(n24035) );
  XOR U26050 ( .A(n24409), .B(n24410), .Z(n24033) );
  AND U26051 ( .A(n24411), .B(n24412), .Z(n24409) );
  AND U26052 ( .A(b[17]), .B(a[45]), .Z(n24408) );
  XOR U26053 ( .A(n24413), .B(n24038), .Z(n24040) );
  XOR U26054 ( .A(n24414), .B(n24415), .Z(n24038) );
  AND U26055 ( .A(n24416), .B(n24417), .Z(n24414) );
  AND U26056 ( .A(b[16]), .B(a[46]), .Z(n24413) );
  XOR U26057 ( .A(n24418), .B(n24043), .Z(n24045) );
  XOR U26058 ( .A(n24419), .B(n24420), .Z(n24043) );
  AND U26059 ( .A(n24421), .B(n24422), .Z(n24419) );
  AND U26060 ( .A(b[15]), .B(a[47]), .Z(n24418) );
  XOR U26061 ( .A(n24423), .B(n24048), .Z(n24050) );
  XOR U26062 ( .A(n24424), .B(n24425), .Z(n24048) );
  AND U26063 ( .A(n24426), .B(n24427), .Z(n24424) );
  AND U26064 ( .A(b[14]), .B(a[48]), .Z(n24423) );
  XOR U26065 ( .A(n24428), .B(n24053), .Z(n24055) );
  XOR U26066 ( .A(n24429), .B(n24430), .Z(n24053) );
  AND U26067 ( .A(n24431), .B(n24432), .Z(n24429) );
  AND U26068 ( .A(b[13]), .B(a[49]), .Z(n24428) );
  XOR U26069 ( .A(n24433), .B(n24058), .Z(n24060) );
  XOR U26070 ( .A(n24434), .B(n24435), .Z(n24058) );
  AND U26071 ( .A(n24436), .B(n24437), .Z(n24434) );
  AND U26072 ( .A(b[12]), .B(a[50]), .Z(n24433) );
  XOR U26073 ( .A(n24438), .B(n24063), .Z(n24065) );
  XOR U26074 ( .A(n24439), .B(n24440), .Z(n24063) );
  AND U26075 ( .A(n24441), .B(n24442), .Z(n24439) );
  AND U26076 ( .A(b[11]), .B(a[51]), .Z(n24438) );
  XOR U26077 ( .A(n24443), .B(n24068), .Z(n24070) );
  XOR U26078 ( .A(n24444), .B(n24445), .Z(n24068) );
  AND U26079 ( .A(n24446), .B(n24447), .Z(n24444) );
  AND U26080 ( .A(b[10]), .B(a[52]), .Z(n24443) );
  XOR U26081 ( .A(n24448), .B(n24073), .Z(n24075) );
  XOR U26082 ( .A(n24449), .B(n24450), .Z(n24073) );
  AND U26083 ( .A(n24451), .B(n24452), .Z(n24449) );
  AND U26084 ( .A(b[9]), .B(a[53]), .Z(n24448) );
  XOR U26085 ( .A(n24453), .B(n24078), .Z(n24080) );
  XOR U26086 ( .A(n24454), .B(n24455), .Z(n24078) );
  AND U26087 ( .A(n24456), .B(n24457), .Z(n24454) );
  AND U26088 ( .A(b[8]), .B(a[54]), .Z(n24453) );
  XOR U26089 ( .A(n24458), .B(n24083), .Z(n24085) );
  XOR U26090 ( .A(n24459), .B(n24460), .Z(n24083) );
  AND U26091 ( .A(n24461), .B(n24462), .Z(n24459) );
  AND U26092 ( .A(b[7]), .B(a[55]), .Z(n24458) );
  XOR U26093 ( .A(n24463), .B(n24088), .Z(n24090) );
  XOR U26094 ( .A(n24464), .B(n24465), .Z(n24088) );
  AND U26095 ( .A(n24466), .B(n24467), .Z(n24464) );
  AND U26096 ( .A(b[6]), .B(a[56]), .Z(n24463) );
  XOR U26097 ( .A(n24468), .B(n24093), .Z(n24095) );
  XOR U26098 ( .A(n24469), .B(n24470), .Z(n24093) );
  AND U26099 ( .A(n24471), .B(n24472), .Z(n24469) );
  AND U26100 ( .A(b[5]), .B(a[57]), .Z(n24468) );
  XOR U26101 ( .A(n24473), .B(n24098), .Z(n24100) );
  XOR U26102 ( .A(n24474), .B(n24475), .Z(n24098) );
  AND U26103 ( .A(n24476), .B(n24477), .Z(n24474) );
  AND U26104 ( .A(b[4]), .B(a[58]), .Z(n24473) );
  XNOR U26105 ( .A(n24478), .B(n24479), .Z(n24112) );
  NANDN U26106 ( .A(n24480), .B(n24481), .Z(n24479) );
  XOR U26107 ( .A(n24482), .B(n24103), .Z(n24105) );
  XNOR U26108 ( .A(n24483), .B(n24484), .Z(n24103) );
  AND U26109 ( .A(n24485), .B(n24486), .Z(n24483) );
  AND U26110 ( .A(b[3]), .B(a[59]), .Z(n24482) );
  XOR U26111 ( .A(n24119), .B(n24118), .Z(c[125]) );
  XOR U26112 ( .A(sreg[189]), .B(n24117), .Z(n24118) );
  XOR U26113 ( .A(n24124), .B(n24487), .Z(n24119) );
  XNOR U26114 ( .A(n24123), .B(n24117), .Z(n24487) );
  XOR U26115 ( .A(n24488), .B(n24489), .Z(n24117) );
  NOR U26116 ( .A(n24490), .B(n24491), .Z(n24488) );
  NAND U26117 ( .A(a[61]), .B(b[0]), .Z(n24123) );
  XNOR U26118 ( .A(n24480), .B(n24481), .Z(n24124) );
  XOR U26119 ( .A(n24478), .B(n24492), .Z(n24481) );
  NAND U26120 ( .A(b[1]), .B(a[60]), .Z(n24492) );
  XOR U26121 ( .A(n24486), .B(n24493), .Z(n24480) );
  XOR U26122 ( .A(n24478), .B(n24485), .Z(n24493) );
  XNOR U26123 ( .A(n24494), .B(n24484), .Z(n24485) );
  AND U26124 ( .A(b[2]), .B(a[59]), .Z(n24494) );
  NANDN U26125 ( .A(n24495), .B(n24496), .Z(n24478) );
  XOR U26126 ( .A(n24484), .B(n24476), .Z(n24497) );
  XNOR U26127 ( .A(n24475), .B(n24471), .Z(n24498) );
  XNOR U26128 ( .A(n24470), .B(n24466), .Z(n24499) );
  XNOR U26129 ( .A(n24465), .B(n24461), .Z(n24500) );
  XNOR U26130 ( .A(n24460), .B(n24456), .Z(n24501) );
  XNOR U26131 ( .A(n24455), .B(n24451), .Z(n24502) );
  XNOR U26132 ( .A(n24450), .B(n24446), .Z(n24503) );
  XNOR U26133 ( .A(n24445), .B(n24441), .Z(n24504) );
  XNOR U26134 ( .A(n24440), .B(n24436), .Z(n24505) );
  XNOR U26135 ( .A(n24435), .B(n24431), .Z(n24506) );
  XNOR U26136 ( .A(n24430), .B(n24426), .Z(n24507) );
  XNOR U26137 ( .A(n24425), .B(n24421), .Z(n24508) );
  XNOR U26138 ( .A(n24420), .B(n24416), .Z(n24509) );
  XNOR U26139 ( .A(n24415), .B(n24411), .Z(n24510) );
  XNOR U26140 ( .A(n24410), .B(n24406), .Z(n24511) );
  XNOR U26141 ( .A(n24405), .B(n24401), .Z(n24512) );
  XNOR U26142 ( .A(n24400), .B(n24396), .Z(n24513) );
  XNOR U26143 ( .A(n24395), .B(n24391), .Z(n24514) );
  XNOR U26144 ( .A(n24390), .B(n24386), .Z(n24515) );
  XNOR U26145 ( .A(n24385), .B(n24381), .Z(n24516) );
  XNOR U26146 ( .A(n24380), .B(n24376), .Z(n24517) );
  XNOR U26147 ( .A(n24375), .B(n24371), .Z(n24518) );
  XNOR U26148 ( .A(n24370), .B(n24366), .Z(n24519) );
  XNOR U26149 ( .A(n24365), .B(n24361), .Z(n24520) );
  XNOR U26150 ( .A(n24360), .B(n24356), .Z(n24521) );
  XNOR U26151 ( .A(n24355), .B(n24351), .Z(n24522) );
  XNOR U26152 ( .A(n24350), .B(n24346), .Z(n24523) );
  XNOR U26153 ( .A(n24345), .B(n24341), .Z(n24524) );
  XNOR U26154 ( .A(n24340), .B(n24336), .Z(n24525) );
  XNOR U26155 ( .A(n24335), .B(n24331), .Z(n24526) );
  XNOR U26156 ( .A(n24330), .B(n24326), .Z(n24527) );
  XNOR U26157 ( .A(n24325), .B(n24321), .Z(n24528) );
  XNOR U26158 ( .A(n24320), .B(n24316), .Z(n24529) );
  XNOR U26159 ( .A(n24315), .B(n24311), .Z(n24530) );
  XNOR U26160 ( .A(n24310), .B(n24306), .Z(n24531) );
  XNOR U26161 ( .A(n24305), .B(n24301), .Z(n24532) );
  XNOR U26162 ( .A(n24300), .B(n24296), .Z(n24533) );
  XNOR U26163 ( .A(n24295), .B(n24291), .Z(n24534) );
  XNOR U26164 ( .A(n24290), .B(n24286), .Z(n24535) );
  XNOR U26165 ( .A(n24285), .B(n24281), .Z(n24536) );
  XNOR U26166 ( .A(n24280), .B(n24276), .Z(n24537) );
  XNOR U26167 ( .A(n24275), .B(n24271), .Z(n24538) );
  XNOR U26168 ( .A(n24270), .B(n24266), .Z(n24539) );
  XNOR U26169 ( .A(n24265), .B(n24261), .Z(n24540) );
  XNOR U26170 ( .A(n24260), .B(n24256), .Z(n24541) );
  XNOR U26171 ( .A(n24255), .B(n24251), .Z(n24542) );
  XNOR U26172 ( .A(n24250), .B(n24246), .Z(n24543) );
  XNOR U26173 ( .A(n24245), .B(n24241), .Z(n24544) );
  XNOR U26174 ( .A(n24240), .B(n24236), .Z(n24545) );
  XNOR U26175 ( .A(n24235), .B(n24231), .Z(n24546) );
  XNOR U26176 ( .A(n24230), .B(n24226), .Z(n24547) );
  XNOR U26177 ( .A(n24225), .B(n24221), .Z(n24548) );
  XNOR U26178 ( .A(n24220), .B(n24216), .Z(n24549) );
  XNOR U26179 ( .A(n24215), .B(n24211), .Z(n24550) );
  XNOR U26180 ( .A(n24210), .B(n24206), .Z(n24551) );
  XNOR U26181 ( .A(n24205), .B(n24201), .Z(n24552) );
  XNOR U26182 ( .A(n24200), .B(n24196), .Z(n24553) );
  XNOR U26183 ( .A(n24195), .B(n24191), .Z(n24554) );
  XOR U26184 ( .A(n24555), .B(n24190), .Z(n24191) );
  AND U26185 ( .A(a[0]), .B(b[61]), .Z(n24555) );
  XOR U26186 ( .A(n24556), .B(n24190), .Z(n24192) );
  XNOR U26187 ( .A(n24557), .B(n24558), .Z(n24190) );
  AND U26188 ( .A(n24559), .B(n24560), .Z(n24557) );
  AND U26189 ( .A(a[1]), .B(b[60]), .Z(n24556) );
  XOR U26190 ( .A(n24561), .B(n24195), .Z(n24197) );
  XOR U26191 ( .A(n24562), .B(n24563), .Z(n24195) );
  AND U26192 ( .A(n24564), .B(n24565), .Z(n24562) );
  AND U26193 ( .A(a[2]), .B(b[59]), .Z(n24561) );
  XOR U26194 ( .A(n24566), .B(n24200), .Z(n24202) );
  XOR U26195 ( .A(n24567), .B(n24568), .Z(n24200) );
  AND U26196 ( .A(n24569), .B(n24570), .Z(n24567) );
  AND U26197 ( .A(a[3]), .B(b[58]), .Z(n24566) );
  XOR U26198 ( .A(n24571), .B(n24205), .Z(n24207) );
  XOR U26199 ( .A(n24572), .B(n24573), .Z(n24205) );
  AND U26200 ( .A(n24574), .B(n24575), .Z(n24572) );
  AND U26201 ( .A(a[4]), .B(b[57]), .Z(n24571) );
  XOR U26202 ( .A(n24576), .B(n24210), .Z(n24212) );
  XOR U26203 ( .A(n24577), .B(n24578), .Z(n24210) );
  AND U26204 ( .A(n24579), .B(n24580), .Z(n24577) );
  AND U26205 ( .A(a[5]), .B(b[56]), .Z(n24576) );
  XOR U26206 ( .A(n24581), .B(n24215), .Z(n24217) );
  XOR U26207 ( .A(n24582), .B(n24583), .Z(n24215) );
  AND U26208 ( .A(n24584), .B(n24585), .Z(n24582) );
  AND U26209 ( .A(a[6]), .B(b[55]), .Z(n24581) );
  XOR U26210 ( .A(n24586), .B(n24220), .Z(n24222) );
  XOR U26211 ( .A(n24587), .B(n24588), .Z(n24220) );
  AND U26212 ( .A(n24589), .B(n24590), .Z(n24587) );
  AND U26213 ( .A(a[7]), .B(b[54]), .Z(n24586) );
  XOR U26214 ( .A(n24591), .B(n24225), .Z(n24227) );
  XOR U26215 ( .A(n24592), .B(n24593), .Z(n24225) );
  AND U26216 ( .A(n24594), .B(n24595), .Z(n24592) );
  AND U26217 ( .A(a[8]), .B(b[53]), .Z(n24591) );
  XOR U26218 ( .A(n24596), .B(n24230), .Z(n24232) );
  XOR U26219 ( .A(n24597), .B(n24598), .Z(n24230) );
  AND U26220 ( .A(n24599), .B(n24600), .Z(n24597) );
  AND U26221 ( .A(a[9]), .B(b[52]), .Z(n24596) );
  XOR U26222 ( .A(n24601), .B(n24235), .Z(n24237) );
  XOR U26223 ( .A(n24602), .B(n24603), .Z(n24235) );
  AND U26224 ( .A(n24604), .B(n24605), .Z(n24602) );
  AND U26225 ( .A(a[10]), .B(b[51]), .Z(n24601) );
  XOR U26226 ( .A(n24606), .B(n24240), .Z(n24242) );
  XOR U26227 ( .A(n24607), .B(n24608), .Z(n24240) );
  AND U26228 ( .A(n24609), .B(n24610), .Z(n24607) );
  AND U26229 ( .A(a[11]), .B(b[50]), .Z(n24606) );
  XOR U26230 ( .A(n24611), .B(n24245), .Z(n24247) );
  XOR U26231 ( .A(n24612), .B(n24613), .Z(n24245) );
  AND U26232 ( .A(n24614), .B(n24615), .Z(n24612) );
  AND U26233 ( .A(a[12]), .B(b[49]), .Z(n24611) );
  XOR U26234 ( .A(n24616), .B(n24250), .Z(n24252) );
  XOR U26235 ( .A(n24617), .B(n24618), .Z(n24250) );
  AND U26236 ( .A(n24619), .B(n24620), .Z(n24617) );
  AND U26237 ( .A(a[13]), .B(b[48]), .Z(n24616) );
  XOR U26238 ( .A(n24621), .B(n24255), .Z(n24257) );
  XOR U26239 ( .A(n24622), .B(n24623), .Z(n24255) );
  AND U26240 ( .A(n24624), .B(n24625), .Z(n24622) );
  AND U26241 ( .A(a[14]), .B(b[47]), .Z(n24621) );
  XOR U26242 ( .A(n24626), .B(n24260), .Z(n24262) );
  XOR U26243 ( .A(n24627), .B(n24628), .Z(n24260) );
  AND U26244 ( .A(n24629), .B(n24630), .Z(n24627) );
  AND U26245 ( .A(a[15]), .B(b[46]), .Z(n24626) );
  XOR U26246 ( .A(n24631), .B(n24265), .Z(n24267) );
  XOR U26247 ( .A(n24632), .B(n24633), .Z(n24265) );
  AND U26248 ( .A(n24634), .B(n24635), .Z(n24632) );
  AND U26249 ( .A(a[16]), .B(b[45]), .Z(n24631) );
  XOR U26250 ( .A(n24636), .B(n24270), .Z(n24272) );
  XOR U26251 ( .A(n24637), .B(n24638), .Z(n24270) );
  AND U26252 ( .A(n24639), .B(n24640), .Z(n24637) );
  AND U26253 ( .A(a[17]), .B(b[44]), .Z(n24636) );
  XOR U26254 ( .A(n24641), .B(n24275), .Z(n24277) );
  XOR U26255 ( .A(n24642), .B(n24643), .Z(n24275) );
  AND U26256 ( .A(n24644), .B(n24645), .Z(n24642) );
  AND U26257 ( .A(a[18]), .B(b[43]), .Z(n24641) );
  XOR U26258 ( .A(n24646), .B(n24280), .Z(n24282) );
  XOR U26259 ( .A(n24647), .B(n24648), .Z(n24280) );
  AND U26260 ( .A(n24649), .B(n24650), .Z(n24647) );
  AND U26261 ( .A(a[19]), .B(b[42]), .Z(n24646) );
  XOR U26262 ( .A(n24651), .B(n24285), .Z(n24287) );
  XOR U26263 ( .A(n24652), .B(n24653), .Z(n24285) );
  AND U26264 ( .A(n24654), .B(n24655), .Z(n24652) );
  AND U26265 ( .A(a[20]), .B(b[41]), .Z(n24651) );
  XOR U26266 ( .A(n24656), .B(n24290), .Z(n24292) );
  XOR U26267 ( .A(n24657), .B(n24658), .Z(n24290) );
  AND U26268 ( .A(n24659), .B(n24660), .Z(n24657) );
  AND U26269 ( .A(a[21]), .B(b[40]), .Z(n24656) );
  XOR U26270 ( .A(n24661), .B(n24295), .Z(n24297) );
  XOR U26271 ( .A(n24662), .B(n24663), .Z(n24295) );
  AND U26272 ( .A(n24664), .B(n24665), .Z(n24662) );
  AND U26273 ( .A(a[22]), .B(b[39]), .Z(n24661) );
  XOR U26274 ( .A(n24666), .B(n24300), .Z(n24302) );
  XOR U26275 ( .A(n24667), .B(n24668), .Z(n24300) );
  AND U26276 ( .A(n24669), .B(n24670), .Z(n24667) );
  AND U26277 ( .A(a[23]), .B(b[38]), .Z(n24666) );
  XOR U26278 ( .A(n24671), .B(n24305), .Z(n24307) );
  XOR U26279 ( .A(n24672), .B(n24673), .Z(n24305) );
  AND U26280 ( .A(n24674), .B(n24675), .Z(n24672) );
  AND U26281 ( .A(a[24]), .B(b[37]), .Z(n24671) );
  XOR U26282 ( .A(n24676), .B(n24310), .Z(n24312) );
  XOR U26283 ( .A(n24677), .B(n24678), .Z(n24310) );
  AND U26284 ( .A(n24679), .B(n24680), .Z(n24677) );
  AND U26285 ( .A(a[25]), .B(b[36]), .Z(n24676) );
  XOR U26286 ( .A(n24681), .B(n24315), .Z(n24317) );
  XOR U26287 ( .A(n24682), .B(n24683), .Z(n24315) );
  AND U26288 ( .A(n24684), .B(n24685), .Z(n24682) );
  AND U26289 ( .A(a[26]), .B(b[35]), .Z(n24681) );
  XOR U26290 ( .A(n24686), .B(n24320), .Z(n24322) );
  XOR U26291 ( .A(n24687), .B(n24688), .Z(n24320) );
  AND U26292 ( .A(n24689), .B(n24690), .Z(n24687) );
  AND U26293 ( .A(a[27]), .B(b[34]), .Z(n24686) );
  XOR U26294 ( .A(n24691), .B(n24325), .Z(n24327) );
  XOR U26295 ( .A(n24692), .B(n24693), .Z(n24325) );
  AND U26296 ( .A(n24694), .B(n24695), .Z(n24692) );
  AND U26297 ( .A(a[28]), .B(b[33]), .Z(n24691) );
  XOR U26298 ( .A(n24696), .B(n24330), .Z(n24332) );
  XOR U26299 ( .A(n24697), .B(n24698), .Z(n24330) );
  AND U26300 ( .A(n24699), .B(n24700), .Z(n24697) );
  AND U26301 ( .A(a[29]), .B(b[32]), .Z(n24696) );
  XOR U26302 ( .A(n24701), .B(n24335), .Z(n24337) );
  XOR U26303 ( .A(n24702), .B(n24703), .Z(n24335) );
  AND U26304 ( .A(n24704), .B(n24705), .Z(n24702) );
  AND U26305 ( .A(a[30]), .B(b[31]), .Z(n24701) );
  XOR U26306 ( .A(n24706), .B(n24340), .Z(n24342) );
  XOR U26307 ( .A(n24707), .B(n24708), .Z(n24340) );
  AND U26308 ( .A(n24709), .B(n24710), .Z(n24707) );
  AND U26309 ( .A(b[30]), .B(a[31]), .Z(n24706) );
  XOR U26310 ( .A(n24711), .B(n24345), .Z(n24347) );
  XOR U26311 ( .A(n24712), .B(n24713), .Z(n24345) );
  AND U26312 ( .A(n24714), .B(n24715), .Z(n24712) );
  AND U26313 ( .A(b[29]), .B(a[32]), .Z(n24711) );
  XOR U26314 ( .A(n24716), .B(n24350), .Z(n24352) );
  XOR U26315 ( .A(n24717), .B(n24718), .Z(n24350) );
  AND U26316 ( .A(n24719), .B(n24720), .Z(n24717) );
  AND U26317 ( .A(b[28]), .B(a[33]), .Z(n24716) );
  XOR U26318 ( .A(n24721), .B(n24355), .Z(n24357) );
  XOR U26319 ( .A(n24722), .B(n24723), .Z(n24355) );
  AND U26320 ( .A(n24724), .B(n24725), .Z(n24722) );
  AND U26321 ( .A(b[27]), .B(a[34]), .Z(n24721) );
  XOR U26322 ( .A(n24726), .B(n24360), .Z(n24362) );
  XOR U26323 ( .A(n24727), .B(n24728), .Z(n24360) );
  AND U26324 ( .A(n24729), .B(n24730), .Z(n24727) );
  AND U26325 ( .A(b[26]), .B(a[35]), .Z(n24726) );
  XOR U26326 ( .A(n24731), .B(n24365), .Z(n24367) );
  XOR U26327 ( .A(n24732), .B(n24733), .Z(n24365) );
  AND U26328 ( .A(n24734), .B(n24735), .Z(n24732) );
  AND U26329 ( .A(b[25]), .B(a[36]), .Z(n24731) );
  XOR U26330 ( .A(n24736), .B(n24370), .Z(n24372) );
  XOR U26331 ( .A(n24737), .B(n24738), .Z(n24370) );
  AND U26332 ( .A(n24739), .B(n24740), .Z(n24737) );
  AND U26333 ( .A(b[24]), .B(a[37]), .Z(n24736) );
  XOR U26334 ( .A(n24741), .B(n24375), .Z(n24377) );
  XOR U26335 ( .A(n24742), .B(n24743), .Z(n24375) );
  AND U26336 ( .A(n24744), .B(n24745), .Z(n24742) );
  AND U26337 ( .A(b[23]), .B(a[38]), .Z(n24741) );
  XOR U26338 ( .A(n24746), .B(n24380), .Z(n24382) );
  XOR U26339 ( .A(n24747), .B(n24748), .Z(n24380) );
  AND U26340 ( .A(n24749), .B(n24750), .Z(n24747) );
  AND U26341 ( .A(b[22]), .B(a[39]), .Z(n24746) );
  XOR U26342 ( .A(n24751), .B(n24385), .Z(n24387) );
  XOR U26343 ( .A(n24752), .B(n24753), .Z(n24385) );
  AND U26344 ( .A(n24754), .B(n24755), .Z(n24752) );
  AND U26345 ( .A(b[21]), .B(a[40]), .Z(n24751) );
  XOR U26346 ( .A(n24756), .B(n24390), .Z(n24392) );
  XOR U26347 ( .A(n24757), .B(n24758), .Z(n24390) );
  AND U26348 ( .A(n24759), .B(n24760), .Z(n24757) );
  AND U26349 ( .A(b[20]), .B(a[41]), .Z(n24756) );
  XOR U26350 ( .A(n24761), .B(n24395), .Z(n24397) );
  XOR U26351 ( .A(n24762), .B(n24763), .Z(n24395) );
  AND U26352 ( .A(n24764), .B(n24765), .Z(n24762) );
  AND U26353 ( .A(b[19]), .B(a[42]), .Z(n24761) );
  XOR U26354 ( .A(n24766), .B(n24400), .Z(n24402) );
  XOR U26355 ( .A(n24767), .B(n24768), .Z(n24400) );
  AND U26356 ( .A(n24769), .B(n24770), .Z(n24767) );
  AND U26357 ( .A(b[18]), .B(a[43]), .Z(n24766) );
  XOR U26358 ( .A(n24771), .B(n24405), .Z(n24407) );
  XOR U26359 ( .A(n24772), .B(n24773), .Z(n24405) );
  AND U26360 ( .A(n24774), .B(n24775), .Z(n24772) );
  AND U26361 ( .A(b[17]), .B(a[44]), .Z(n24771) );
  XOR U26362 ( .A(n24776), .B(n24410), .Z(n24412) );
  XOR U26363 ( .A(n24777), .B(n24778), .Z(n24410) );
  AND U26364 ( .A(n24779), .B(n24780), .Z(n24777) );
  AND U26365 ( .A(b[16]), .B(a[45]), .Z(n24776) );
  XOR U26366 ( .A(n24781), .B(n24415), .Z(n24417) );
  XOR U26367 ( .A(n24782), .B(n24783), .Z(n24415) );
  AND U26368 ( .A(n24784), .B(n24785), .Z(n24782) );
  AND U26369 ( .A(b[15]), .B(a[46]), .Z(n24781) );
  XOR U26370 ( .A(n24786), .B(n24420), .Z(n24422) );
  XOR U26371 ( .A(n24787), .B(n24788), .Z(n24420) );
  AND U26372 ( .A(n24789), .B(n24790), .Z(n24787) );
  AND U26373 ( .A(b[14]), .B(a[47]), .Z(n24786) );
  XOR U26374 ( .A(n24791), .B(n24425), .Z(n24427) );
  XOR U26375 ( .A(n24792), .B(n24793), .Z(n24425) );
  AND U26376 ( .A(n24794), .B(n24795), .Z(n24792) );
  AND U26377 ( .A(b[13]), .B(a[48]), .Z(n24791) );
  XOR U26378 ( .A(n24796), .B(n24430), .Z(n24432) );
  XOR U26379 ( .A(n24797), .B(n24798), .Z(n24430) );
  AND U26380 ( .A(n24799), .B(n24800), .Z(n24797) );
  AND U26381 ( .A(b[12]), .B(a[49]), .Z(n24796) );
  XOR U26382 ( .A(n24801), .B(n24435), .Z(n24437) );
  XOR U26383 ( .A(n24802), .B(n24803), .Z(n24435) );
  AND U26384 ( .A(n24804), .B(n24805), .Z(n24802) );
  AND U26385 ( .A(b[11]), .B(a[50]), .Z(n24801) );
  XOR U26386 ( .A(n24806), .B(n24440), .Z(n24442) );
  XOR U26387 ( .A(n24807), .B(n24808), .Z(n24440) );
  AND U26388 ( .A(n24809), .B(n24810), .Z(n24807) );
  AND U26389 ( .A(b[10]), .B(a[51]), .Z(n24806) );
  XOR U26390 ( .A(n24811), .B(n24445), .Z(n24447) );
  XOR U26391 ( .A(n24812), .B(n24813), .Z(n24445) );
  AND U26392 ( .A(n24814), .B(n24815), .Z(n24812) );
  AND U26393 ( .A(b[9]), .B(a[52]), .Z(n24811) );
  XOR U26394 ( .A(n24816), .B(n24450), .Z(n24452) );
  XOR U26395 ( .A(n24817), .B(n24818), .Z(n24450) );
  AND U26396 ( .A(n24819), .B(n24820), .Z(n24817) );
  AND U26397 ( .A(b[8]), .B(a[53]), .Z(n24816) );
  XOR U26398 ( .A(n24821), .B(n24455), .Z(n24457) );
  XOR U26399 ( .A(n24822), .B(n24823), .Z(n24455) );
  AND U26400 ( .A(n24824), .B(n24825), .Z(n24822) );
  AND U26401 ( .A(b[7]), .B(a[54]), .Z(n24821) );
  XOR U26402 ( .A(n24826), .B(n24460), .Z(n24462) );
  XOR U26403 ( .A(n24827), .B(n24828), .Z(n24460) );
  AND U26404 ( .A(n24829), .B(n24830), .Z(n24827) );
  AND U26405 ( .A(b[6]), .B(a[55]), .Z(n24826) );
  XOR U26406 ( .A(n24831), .B(n24465), .Z(n24467) );
  XOR U26407 ( .A(n24832), .B(n24833), .Z(n24465) );
  AND U26408 ( .A(n24834), .B(n24835), .Z(n24832) );
  AND U26409 ( .A(b[5]), .B(a[56]), .Z(n24831) );
  XOR U26410 ( .A(n24836), .B(n24470), .Z(n24472) );
  XOR U26411 ( .A(n24837), .B(n24838), .Z(n24470) );
  AND U26412 ( .A(n24839), .B(n24840), .Z(n24837) );
  AND U26413 ( .A(b[4]), .B(a[57]), .Z(n24836) );
  XNOR U26414 ( .A(n24841), .B(n24842), .Z(n24484) );
  NANDN U26415 ( .A(n24843), .B(n24844), .Z(n24842) );
  XOR U26416 ( .A(n24845), .B(n24475), .Z(n24477) );
  XNOR U26417 ( .A(n24846), .B(n24847), .Z(n24475) );
  AND U26418 ( .A(n24848), .B(n24849), .Z(n24846) );
  AND U26419 ( .A(b[3]), .B(a[58]), .Z(n24845) );
  XOR U26420 ( .A(n24491), .B(n24490), .Z(c[124]) );
  XOR U26421 ( .A(sreg[188]), .B(n24489), .Z(n24490) );
  XOR U26422 ( .A(n24496), .B(n24850), .Z(n24491) );
  XNOR U26423 ( .A(n24495), .B(n24489), .Z(n24850) );
  XOR U26424 ( .A(n24851), .B(n24852), .Z(n24489) );
  NOR U26425 ( .A(n24853), .B(n24854), .Z(n24851) );
  NAND U26426 ( .A(a[60]), .B(b[0]), .Z(n24495) );
  XNOR U26427 ( .A(n24843), .B(n24844), .Z(n24496) );
  XOR U26428 ( .A(n24841), .B(n24855), .Z(n24844) );
  NAND U26429 ( .A(b[1]), .B(a[59]), .Z(n24855) );
  XOR U26430 ( .A(n24849), .B(n24856), .Z(n24843) );
  XOR U26431 ( .A(n24841), .B(n24848), .Z(n24856) );
  XNOR U26432 ( .A(n24857), .B(n24847), .Z(n24848) );
  AND U26433 ( .A(b[2]), .B(a[58]), .Z(n24857) );
  NANDN U26434 ( .A(n24858), .B(n24859), .Z(n24841) );
  XOR U26435 ( .A(n24847), .B(n24839), .Z(n24860) );
  XNOR U26436 ( .A(n24838), .B(n24834), .Z(n24861) );
  XNOR U26437 ( .A(n24833), .B(n24829), .Z(n24862) );
  XNOR U26438 ( .A(n24828), .B(n24824), .Z(n24863) );
  XNOR U26439 ( .A(n24823), .B(n24819), .Z(n24864) );
  XNOR U26440 ( .A(n24818), .B(n24814), .Z(n24865) );
  XNOR U26441 ( .A(n24813), .B(n24809), .Z(n24866) );
  XNOR U26442 ( .A(n24808), .B(n24804), .Z(n24867) );
  XNOR U26443 ( .A(n24803), .B(n24799), .Z(n24868) );
  XNOR U26444 ( .A(n24798), .B(n24794), .Z(n24869) );
  XNOR U26445 ( .A(n24793), .B(n24789), .Z(n24870) );
  XNOR U26446 ( .A(n24788), .B(n24784), .Z(n24871) );
  XNOR U26447 ( .A(n24783), .B(n24779), .Z(n24872) );
  XNOR U26448 ( .A(n24778), .B(n24774), .Z(n24873) );
  XNOR U26449 ( .A(n24773), .B(n24769), .Z(n24874) );
  XNOR U26450 ( .A(n24768), .B(n24764), .Z(n24875) );
  XNOR U26451 ( .A(n24763), .B(n24759), .Z(n24876) );
  XNOR U26452 ( .A(n24758), .B(n24754), .Z(n24877) );
  XNOR U26453 ( .A(n24753), .B(n24749), .Z(n24878) );
  XNOR U26454 ( .A(n24748), .B(n24744), .Z(n24879) );
  XNOR U26455 ( .A(n24743), .B(n24739), .Z(n24880) );
  XNOR U26456 ( .A(n24738), .B(n24734), .Z(n24881) );
  XNOR U26457 ( .A(n24733), .B(n24729), .Z(n24882) );
  XNOR U26458 ( .A(n24728), .B(n24724), .Z(n24883) );
  XNOR U26459 ( .A(n24723), .B(n24719), .Z(n24884) );
  XNOR U26460 ( .A(n24718), .B(n24714), .Z(n24885) );
  XNOR U26461 ( .A(n24713), .B(n24709), .Z(n24886) );
  XNOR U26462 ( .A(n24708), .B(n24704), .Z(n24887) );
  XNOR U26463 ( .A(n24703), .B(n24699), .Z(n24888) );
  XNOR U26464 ( .A(n24698), .B(n24694), .Z(n24889) );
  XNOR U26465 ( .A(n24693), .B(n24689), .Z(n24890) );
  XNOR U26466 ( .A(n24688), .B(n24684), .Z(n24891) );
  XNOR U26467 ( .A(n24683), .B(n24679), .Z(n24892) );
  XNOR U26468 ( .A(n24678), .B(n24674), .Z(n24893) );
  XNOR U26469 ( .A(n24673), .B(n24669), .Z(n24894) );
  XNOR U26470 ( .A(n24668), .B(n24664), .Z(n24895) );
  XNOR U26471 ( .A(n24663), .B(n24659), .Z(n24896) );
  XNOR U26472 ( .A(n24658), .B(n24654), .Z(n24897) );
  XNOR U26473 ( .A(n24653), .B(n24649), .Z(n24898) );
  XNOR U26474 ( .A(n24648), .B(n24644), .Z(n24899) );
  XNOR U26475 ( .A(n24643), .B(n24639), .Z(n24900) );
  XNOR U26476 ( .A(n24638), .B(n24634), .Z(n24901) );
  XNOR U26477 ( .A(n24633), .B(n24629), .Z(n24902) );
  XNOR U26478 ( .A(n24628), .B(n24624), .Z(n24903) );
  XNOR U26479 ( .A(n24623), .B(n24619), .Z(n24904) );
  XNOR U26480 ( .A(n24618), .B(n24614), .Z(n24905) );
  XNOR U26481 ( .A(n24613), .B(n24609), .Z(n24906) );
  XNOR U26482 ( .A(n24608), .B(n24604), .Z(n24907) );
  XNOR U26483 ( .A(n24603), .B(n24599), .Z(n24908) );
  XNOR U26484 ( .A(n24598), .B(n24594), .Z(n24909) );
  XNOR U26485 ( .A(n24593), .B(n24589), .Z(n24910) );
  XNOR U26486 ( .A(n24588), .B(n24584), .Z(n24911) );
  XNOR U26487 ( .A(n24583), .B(n24579), .Z(n24912) );
  XNOR U26488 ( .A(n24578), .B(n24574), .Z(n24913) );
  XNOR U26489 ( .A(n24573), .B(n24569), .Z(n24914) );
  XNOR U26490 ( .A(n24568), .B(n24564), .Z(n24915) );
  XNOR U26491 ( .A(n24563), .B(n24559), .Z(n24916) );
  XNOR U26492 ( .A(n24917), .B(n24558), .Z(n24559) );
  AND U26493 ( .A(a[0]), .B(b[60]), .Z(n24917) );
  XNOR U26494 ( .A(n24918), .B(n24558), .Z(n24560) );
  XNOR U26495 ( .A(n24919), .B(n24920), .Z(n24558) );
  AND U26496 ( .A(n24921), .B(n24922), .Z(n24919) );
  AND U26497 ( .A(a[1]), .B(b[59]), .Z(n24918) );
  XOR U26498 ( .A(n24923), .B(n24563), .Z(n24565) );
  XOR U26499 ( .A(n24924), .B(n24925), .Z(n24563) );
  AND U26500 ( .A(n24926), .B(n24927), .Z(n24924) );
  AND U26501 ( .A(a[2]), .B(b[58]), .Z(n24923) );
  XOR U26502 ( .A(n24928), .B(n24568), .Z(n24570) );
  XOR U26503 ( .A(n24929), .B(n24930), .Z(n24568) );
  AND U26504 ( .A(n24931), .B(n24932), .Z(n24929) );
  AND U26505 ( .A(a[3]), .B(b[57]), .Z(n24928) );
  XOR U26506 ( .A(n24933), .B(n24573), .Z(n24575) );
  XOR U26507 ( .A(n24934), .B(n24935), .Z(n24573) );
  AND U26508 ( .A(n24936), .B(n24937), .Z(n24934) );
  AND U26509 ( .A(a[4]), .B(b[56]), .Z(n24933) );
  XOR U26510 ( .A(n24938), .B(n24578), .Z(n24580) );
  XOR U26511 ( .A(n24939), .B(n24940), .Z(n24578) );
  AND U26512 ( .A(n24941), .B(n24942), .Z(n24939) );
  AND U26513 ( .A(a[5]), .B(b[55]), .Z(n24938) );
  XOR U26514 ( .A(n24943), .B(n24583), .Z(n24585) );
  XOR U26515 ( .A(n24944), .B(n24945), .Z(n24583) );
  AND U26516 ( .A(n24946), .B(n24947), .Z(n24944) );
  AND U26517 ( .A(a[6]), .B(b[54]), .Z(n24943) );
  XOR U26518 ( .A(n24948), .B(n24588), .Z(n24590) );
  XOR U26519 ( .A(n24949), .B(n24950), .Z(n24588) );
  AND U26520 ( .A(n24951), .B(n24952), .Z(n24949) );
  AND U26521 ( .A(a[7]), .B(b[53]), .Z(n24948) );
  XOR U26522 ( .A(n24953), .B(n24593), .Z(n24595) );
  XOR U26523 ( .A(n24954), .B(n24955), .Z(n24593) );
  AND U26524 ( .A(n24956), .B(n24957), .Z(n24954) );
  AND U26525 ( .A(a[8]), .B(b[52]), .Z(n24953) );
  XOR U26526 ( .A(n24958), .B(n24598), .Z(n24600) );
  XOR U26527 ( .A(n24959), .B(n24960), .Z(n24598) );
  AND U26528 ( .A(n24961), .B(n24962), .Z(n24959) );
  AND U26529 ( .A(a[9]), .B(b[51]), .Z(n24958) );
  XOR U26530 ( .A(n24963), .B(n24603), .Z(n24605) );
  XOR U26531 ( .A(n24964), .B(n24965), .Z(n24603) );
  AND U26532 ( .A(n24966), .B(n24967), .Z(n24964) );
  AND U26533 ( .A(a[10]), .B(b[50]), .Z(n24963) );
  XOR U26534 ( .A(n24968), .B(n24608), .Z(n24610) );
  XOR U26535 ( .A(n24969), .B(n24970), .Z(n24608) );
  AND U26536 ( .A(n24971), .B(n24972), .Z(n24969) );
  AND U26537 ( .A(a[11]), .B(b[49]), .Z(n24968) );
  XOR U26538 ( .A(n24973), .B(n24613), .Z(n24615) );
  XOR U26539 ( .A(n24974), .B(n24975), .Z(n24613) );
  AND U26540 ( .A(n24976), .B(n24977), .Z(n24974) );
  AND U26541 ( .A(a[12]), .B(b[48]), .Z(n24973) );
  XOR U26542 ( .A(n24978), .B(n24618), .Z(n24620) );
  XOR U26543 ( .A(n24979), .B(n24980), .Z(n24618) );
  AND U26544 ( .A(n24981), .B(n24982), .Z(n24979) );
  AND U26545 ( .A(a[13]), .B(b[47]), .Z(n24978) );
  XOR U26546 ( .A(n24983), .B(n24623), .Z(n24625) );
  XOR U26547 ( .A(n24984), .B(n24985), .Z(n24623) );
  AND U26548 ( .A(n24986), .B(n24987), .Z(n24984) );
  AND U26549 ( .A(a[14]), .B(b[46]), .Z(n24983) );
  XOR U26550 ( .A(n24988), .B(n24628), .Z(n24630) );
  XOR U26551 ( .A(n24989), .B(n24990), .Z(n24628) );
  AND U26552 ( .A(n24991), .B(n24992), .Z(n24989) );
  AND U26553 ( .A(a[15]), .B(b[45]), .Z(n24988) );
  XOR U26554 ( .A(n24993), .B(n24633), .Z(n24635) );
  XOR U26555 ( .A(n24994), .B(n24995), .Z(n24633) );
  AND U26556 ( .A(n24996), .B(n24997), .Z(n24994) );
  AND U26557 ( .A(a[16]), .B(b[44]), .Z(n24993) );
  XOR U26558 ( .A(n24998), .B(n24638), .Z(n24640) );
  XOR U26559 ( .A(n24999), .B(n25000), .Z(n24638) );
  AND U26560 ( .A(n25001), .B(n25002), .Z(n24999) );
  AND U26561 ( .A(a[17]), .B(b[43]), .Z(n24998) );
  XOR U26562 ( .A(n25003), .B(n24643), .Z(n24645) );
  XOR U26563 ( .A(n25004), .B(n25005), .Z(n24643) );
  AND U26564 ( .A(n25006), .B(n25007), .Z(n25004) );
  AND U26565 ( .A(a[18]), .B(b[42]), .Z(n25003) );
  XOR U26566 ( .A(n25008), .B(n24648), .Z(n24650) );
  XOR U26567 ( .A(n25009), .B(n25010), .Z(n24648) );
  AND U26568 ( .A(n25011), .B(n25012), .Z(n25009) );
  AND U26569 ( .A(a[19]), .B(b[41]), .Z(n25008) );
  XOR U26570 ( .A(n25013), .B(n24653), .Z(n24655) );
  XOR U26571 ( .A(n25014), .B(n25015), .Z(n24653) );
  AND U26572 ( .A(n25016), .B(n25017), .Z(n25014) );
  AND U26573 ( .A(a[20]), .B(b[40]), .Z(n25013) );
  XOR U26574 ( .A(n25018), .B(n24658), .Z(n24660) );
  XOR U26575 ( .A(n25019), .B(n25020), .Z(n24658) );
  AND U26576 ( .A(n25021), .B(n25022), .Z(n25019) );
  AND U26577 ( .A(a[21]), .B(b[39]), .Z(n25018) );
  XOR U26578 ( .A(n25023), .B(n24663), .Z(n24665) );
  XOR U26579 ( .A(n25024), .B(n25025), .Z(n24663) );
  AND U26580 ( .A(n25026), .B(n25027), .Z(n25024) );
  AND U26581 ( .A(a[22]), .B(b[38]), .Z(n25023) );
  XOR U26582 ( .A(n25028), .B(n24668), .Z(n24670) );
  XOR U26583 ( .A(n25029), .B(n25030), .Z(n24668) );
  AND U26584 ( .A(n25031), .B(n25032), .Z(n25029) );
  AND U26585 ( .A(a[23]), .B(b[37]), .Z(n25028) );
  XOR U26586 ( .A(n25033), .B(n24673), .Z(n24675) );
  XOR U26587 ( .A(n25034), .B(n25035), .Z(n24673) );
  AND U26588 ( .A(n25036), .B(n25037), .Z(n25034) );
  AND U26589 ( .A(a[24]), .B(b[36]), .Z(n25033) );
  XOR U26590 ( .A(n25038), .B(n24678), .Z(n24680) );
  XOR U26591 ( .A(n25039), .B(n25040), .Z(n24678) );
  AND U26592 ( .A(n25041), .B(n25042), .Z(n25039) );
  AND U26593 ( .A(a[25]), .B(b[35]), .Z(n25038) );
  XOR U26594 ( .A(n25043), .B(n24683), .Z(n24685) );
  XOR U26595 ( .A(n25044), .B(n25045), .Z(n24683) );
  AND U26596 ( .A(n25046), .B(n25047), .Z(n25044) );
  AND U26597 ( .A(a[26]), .B(b[34]), .Z(n25043) );
  XOR U26598 ( .A(n25048), .B(n24688), .Z(n24690) );
  XOR U26599 ( .A(n25049), .B(n25050), .Z(n24688) );
  AND U26600 ( .A(n25051), .B(n25052), .Z(n25049) );
  AND U26601 ( .A(a[27]), .B(b[33]), .Z(n25048) );
  XOR U26602 ( .A(n25053), .B(n24693), .Z(n24695) );
  XOR U26603 ( .A(n25054), .B(n25055), .Z(n24693) );
  AND U26604 ( .A(n25056), .B(n25057), .Z(n25054) );
  AND U26605 ( .A(a[28]), .B(b[32]), .Z(n25053) );
  XOR U26606 ( .A(n25058), .B(n24698), .Z(n24700) );
  XOR U26607 ( .A(n25059), .B(n25060), .Z(n24698) );
  AND U26608 ( .A(n25061), .B(n25062), .Z(n25059) );
  AND U26609 ( .A(a[29]), .B(b[31]), .Z(n25058) );
  XOR U26610 ( .A(n25063), .B(n24703), .Z(n24705) );
  XOR U26611 ( .A(n25064), .B(n25065), .Z(n24703) );
  AND U26612 ( .A(n25066), .B(n25067), .Z(n25064) );
  AND U26613 ( .A(a[30]), .B(b[30]), .Z(n25063) );
  XOR U26614 ( .A(n25068), .B(n24708), .Z(n24710) );
  XOR U26615 ( .A(n25069), .B(n25070), .Z(n24708) );
  AND U26616 ( .A(n25071), .B(n25072), .Z(n25069) );
  AND U26617 ( .A(b[29]), .B(a[31]), .Z(n25068) );
  XOR U26618 ( .A(n25073), .B(n24713), .Z(n24715) );
  XOR U26619 ( .A(n25074), .B(n25075), .Z(n24713) );
  AND U26620 ( .A(n25076), .B(n25077), .Z(n25074) );
  AND U26621 ( .A(b[28]), .B(a[32]), .Z(n25073) );
  XOR U26622 ( .A(n25078), .B(n24718), .Z(n24720) );
  XOR U26623 ( .A(n25079), .B(n25080), .Z(n24718) );
  AND U26624 ( .A(n25081), .B(n25082), .Z(n25079) );
  AND U26625 ( .A(b[27]), .B(a[33]), .Z(n25078) );
  XOR U26626 ( .A(n25083), .B(n24723), .Z(n24725) );
  XOR U26627 ( .A(n25084), .B(n25085), .Z(n24723) );
  AND U26628 ( .A(n25086), .B(n25087), .Z(n25084) );
  AND U26629 ( .A(b[26]), .B(a[34]), .Z(n25083) );
  XOR U26630 ( .A(n25088), .B(n24728), .Z(n24730) );
  XOR U26631 ( .A(n25089), .B(n25090), .Z(n24728) );
  AND U26632 ( .A(n25091), .B(n25092), .Z(n25089) );
  AND U26633 ( .A(b[25]), .B(a[35]), .Z(n25088) );
  XOR U26634 ( .A(n25093), .B(n24733), .Z(n24735) );
  XOR U26635 ( .A(n25094), .B(n25095), .Z(n24733) );
  AND U26636 ( .A(n25096), .B(n25097), .Z(n25094) );
  AND U26637 ( .A(b[24]), .B(a[36]), .Z(n25093) );
  XOR U26638 ( .A(n25098), .B(n24738), .Z(n24740) );
  XOR U26639 ( .A(n25099), .B(n25100), .Z(n24738) );
  AND U26640 ( .A(n25101), .B(n25102), .Z(n25099) );
  AND U26641 ( .A(b[23]), .B(a[37]), .Z(n25098) );
  XOR U26642 ( .A(n25103), .B(n24743), .Z(n24745) );
  XOR U26643 ( .A(n25104), .B(n25105), .Z(n24743) );
  AND U26644 ( .A(n25106), .B(n25107), .Z(n25104) );
  AND U26645 ( .A(b[22]), .B(a[38]), .Z(n25103) );
  XOR U26646 ( .A(n25108), .B(n24748), .Z(n24750) );
  XOR U26647 ( .A(n25109), .B(n25110), .Z(n24748) );
  AND U26648 ( .A(n25111), .B(n25112), .Z(n25109) );
  AND U26649 ( .A(b[21]), .B(a[39]), .Z(n25108) );
  XOR U26650 ( .A(n25113), .B(n24753), .Z(n24755) );
  XOR U26651 ( .A(n25114), .B(n25115), .Z(n24753) );
  AND U26652 ( .A(n25116), .B(n25117), .Z(n25114) );
  AND U26653 ( .A(b[20]), .B(a[40]), .Z(n25113) );
  XOR U26654 ( .A(n25118), .B(n24758), .Z(n24760) );
  XOR U26655 ( .A(n25119), .B(n25120), .Z(n24758) );
  AND U26656 ( .A(n25121), .B(n25122), .Z(n25119) );
  AND U26657 ( .A(b[19]), .B(a[41]), .Z(n25118) );
  XOR U26658 ( .A(n25123), .B(n24763), .Z(n24765) );
  XOR U26659 ( .A(n25124), .B(n25125), .Z(n24763) );
  AND U26660 ( .A(n25126), .B(n25127), .Z(n25124) );
  AND U26661 ( .A(b[18]), .B(a[42]), .Z(n25123) );
  XOR U26662 ( .A(n25128), .B(n24768), .Z(n24770) );
  XOR U26663 ( .A(n25129), .B(n25130), .Z(n24768) );
  AND U26664 ( .A(n25131), .B(n25132), .Z(n25129) );
  AND U26665 ( .A(b[17]), .B(a[43]), .Z(n25128) );
  XOR U26666 ( .A(n25133), .B(n24773), .Z(n24775) );
  XOR U26667 ( .A(n25134), .B(n25135), .Z(n24773) );
  AND U26668 ( .A(n25136), .B(n25137), .Z(n25134) );
  AND U26669 ( .A(b[16]), .B(a[44]), .Z(n25133) );
  XOR U26670 ( .A(n25138), .B(n24778), .Z(n24780) );
  XOR U26671 ( .A(n25139), .B(n25140), .Z(n24778) );
  AND U26672 ( .A(n25141), .B(n25142), .Z(n25139) );
  AND U26673 ( .A(b[15]), .B(a[45]), .Z(n25138) );
  XOR U26674 ( .A(n25143), .B(n24783), .Z(n24785) );
  XOR U26675 ( .A(n25144), .B(n25145), .Z(n24783) );
  AND U26676 ( .A(n25146), .B(n25147), .Z(n25144) );
  AND U26677 ( .A(b[14]), .B(a[46]), .Z(n25143) );
  XOR U26678 ( .A(n25148), .B(n24788), .Z(n24790) );
  XOR U26679 ( .A(n25149), .B(n25150), .Z(n24788) );
  AND U26680 ( .A(n25151), .B(n25152), .Z(n25149) );
  AND U26681 ( .A(b[13]), .B(a[47]), .Z(n25148) );
  XOR U26682 ( .A(n25153), .B(n24793), .Z(n24795) );
  XOR U26683 ( .A(n25154), .B(n25155), .Z(n24793) );
  AND U26684 ( .A(n25156), .B(n25157), .Z(n25154) );
  AND U26685 ( .A(b[12]), .B(a[48]), .Z(n25153) );
  XOR U26686 ( .A(n25158), .B(n24798), .Z(n24800) );
  XOR U26687 ( .A(n25159), .B(n25160), .Z(n24798) );
  AND U26688 ( .A(n25161), .B(n25162), .Z(n25159) );
  AND U26689 ( .A(b[11]), .B(a[49]), .Z(n25158) );
  XOR U26690 ( .A(n25163), .B(n24803), .Z(n24805) );
  XOR U26691 ( .A(n25164), .B(n25165), .Z(n24803) );
  AND U26692 ( .A(n25166), .B(n25167), .Z(n25164) );
  AND U26693 ( .A(b[10]), .B(a[50]), .Z(n25163) );
  XOR U26694 ( .A(n25168), .B(n24808), .Z(n24810) );
  XOR U26695 ( .A(n25169), .B(n25170), .Z(n24808) );
  AND U26696 ( .A(n25171), .B(n25172), .Z(n25169) );
  AND U26697 ( .A(b[9]), .B(a[51]), .Z(n25168) );
  XOR U26698 ( .A(n25173), .B(n24813), .Z(n24815) );
  XOR U26699 ( .A(n25174), .B(n25175), .Z(n24813) );
  AND U26700 ( .A(n25176), .B(n25177), .Z(n25174) );
  AND U26701 ( .A(b[8]), .B(a[52]), .Z(n25173) );
  XOR U26702 ( .A(n25178), .B(n24818), .Z(n24820) );
  XOR U26703 ( .A(n25179), .B(n25180), .Z(n24818) );
  AND U26704 ( .A(n25181), .B(n25182), .Z(n25179) );
  AND U26705 ( .A(b[7]), .B(a[53]), .Z(n25178) );
  XOR U26706 ( .A(n25183), .B(n24823), .Z(n24825) );
  XOR U26707 ( .A(n25184), .B(n25185), .Z(n24823) );
  AND U26708 ( .A(n25186), .B(n25187), .Z(n25184) );
  AND U26709 ( .A(b[6]), .B(a[54]), .Z(n25183) );
  XOR U26710 ( .A(n25188), .B(n24828), .Z(n24830) );
  XOR U26711 ( .A(n25189), .B(n25190), .Z(n24828) );
  AND U26712 ( .A(n25191), .B(n25192), .Z(n25189) );
  AND U26713 ( .A(b[5]), .B(a[55]), .Z(n25188) );
  XOR U26714 ( .A(n25193), .B(n24833), .Z(n24835) );
  XOR U26715 ( .A(n25194), .B(n25195), .Z(n24833) );
  AND U26716 ( .A(n25196), .B(n25197), .Z(n25194) );
  AND U26717 ( .A(b[4]), .B(a[56]), .Z(n25193) );
  XNOR U26718 ( .A(n25198), .B(n25199), .Z(n24847) );
  NANDN U26719 ( .A(n25200), .B(n25201), .Z(n25199) );
  XOR U26720 ( .A(n25202), .B(n24838), .Z(n24840) );
  XNOR U26721 ( .A(n25203), .B(n25204), .Z(n24838) );
  AND U26722 ( .A(n25205), .B(n25206), .Z(n25203) );
  AND U26723 ( .A(b[3]), .B(a[57]), .Z(n25202) );
  XOR U26724 ( .A(n24854), .B(n24853), .Z(c[123]) );
  XOR U26725 ( .A(sreg[187]), .B(n24852), .Z(n24853) );
  XOR U26726 ( .A(n24859), .B(n25207), .Z(n24854) );
  XNOR U26727 ( .A(n24858), .B(n24852), .Z(n25207) );
  XOR U26728 ( .A(n25208), .B(n25209), .Z(n24852) );
  NOR U26729 ( .A(n25210), .B(n25211), .Z(n25208) );
  NAND U26730 ( .A(a[59]), .B(b[0]), .Z(n24858) );
  XNOR U26731 ( .A(n25200), .B(n25201), .Z(n24859) );
  XOR U26732 ( .A(n25198), .B(n25212), .Z(n25201) );
  NAND U26733 ( .A(b[1]), .B(a[58]), .Z(n25212) );
  XOR U26734 ( .A(n25206), .B(n25213), .Z(n25200) );
  XOR U26735 ( .A(n25198), .B(n25205), .Z(n25213) );
  XNOR U26736 ( .A(n25214), .B(n25204), .Z(n25205) );
  AND U26737 ( .A(b[2]), .B(a[57]), .Z(n25214) );
  NANDN U26738 ( .A(n25215), .B(n25216), .Z(n25198) );
  XOR U26739 ( .A(n25204), .B(n25196), .Z(n25217) );
  XNOR U26740 ( .A(n25195), .B(n25191), .Z(n25218) );
  XNOR U26741 ( .A(n25190), .B(n25186), .Z(n25219) );
  XNOR U26742 ( .A(n25185), .B(n25181), .Z(n25220) );
  XNOR U26743 ( .A(n25180), .B(n25176), .Z(n25221) );
  XNOR U26744 ( .A(n25175), .B(n25171), .Z(n25222) );
  XNOR U26745 ( .A(n25170), .B(n25166), .Z(n25223) );
  XNOR U26746 ( .A(n25165), .B(n25161), .Z(n25224) );
  XNOR U26747 ( .A(n25160), .B(n25156), .Z(n25225) );
  XNOR U26748 ( .A(n25155), .B(n25151), .Z(n25226) );
  XNOR U26749 ( .A(n25150), .B(n25146), .Z(n25227) );
  XNOR U26750 ( .A(n25145), .B(n25141), .Z(n25228) );
  XNOR U26751 ( .A(n25140), .B(n25136), .Z(n25229) );
  XNOR U26752 ( .A(n25135), .B(n25131), .Z(n25230) );
  XNOR U26753 ( .A(n25130), .B(n25126), .Z(n25231) );
  XNOR U26754 ( .A(n25125), .B(n25121), .Z(n25232) );
  XNOR U26755 ( .A(n25120), .B(n25116), .Z(n25233) );
  XNOR U26756 ( .A(n25115), .B(n25111), .Z(n25234) );
  XNOR U26757 ( .A(n25110), .B(n25106), .Z(n25235) );
  XNOR U26758 ( .A(n25105), .B(n25101), .Z(n25236) );
  XNOR U26759 ( .A(n25100), .B(n25096), .Z(n25237) );
  XNOR U26760 ( .A(n25095), .B(n25091), .Z(n25238) );
  XNOR U26761 ( .A(n25090), .B(n25086), .Z(n25239) );
  XNOR U26762 ( .A(n25085), .B(n25081), .Z(n25240) );
  XNOR U26763 ( .A(n25080), .B(n25076), .Z(n25241) );
  XNOR U26764 ( .A(n25075), .B(n25071), .Z(n25242) );
  XNOR U26765 ( .A(n25070), .B(n25066), .Z(n25243) );
  XNOR U26766 ( .A(n25065), .B(n25061), .Z(n25244) );
  XNOR U26767 ( .A(n25060), .B(n25056), .Z(n25245) );
  XNOR U26768 ( .A(n25055), .B(n25051), .Z(n25246) );
  XNOR U26769 ( .A(n25050), .B(n25046), .Z(n25247) );
  XNOR U26770 ( .A(n25045), .B(n25041), .Z(n25248) );
  XNOR U26771 ( .A(n25040), .B(n25036), .Z(n25249) );
  XNOR U26772 ( .A(n25035), .B(n25031), .Z(n25250) );
  XNOR U26773 ( .A(n25030), .B(n25026), .Z(n25251) );
  XNOR U26774 ( .A(n25025), .B(n25021), .Z(n25252) );
  XNOR U26775 ( .A(n25020), .B(n25016), .Z(n25253) );
  XNOR U26776 ( .A(n25015), .B(n25011), .Z(n25254) );
  XNOR U26777 ( .A(n25010), .B(n25006), .Z(n25255) );
  XNOR U26778 ( .A(n25005), .B(n25001), .Z(n25256) );
  XNOR U26779 ( .A(n25000), .B(n24996), .Z(n25257) );
  XNOR U26780 ( .A(n24995), .B(n24991), .Z(n25258) );
  XNOR U26781 ( .A(n24990), .B(n24986), .Z(n25259) );
  XNOR U26782 ( .A(n24985), .B(n24981), .Z(n25260) );
  XNOR U26783 ( .A(n24980), .B(n24976), .Z(n25261) );
  XNOR U26784 ( .A(n24975), .B(n24971), .Z(n25262) );
  XNOR U26785 ( .A(n24970), .B(n24966), .Z(n25263) );
  XNOR U26786 ( .A(n24965), .B(n24961), .Z(n25264) );
  XNOR U26787 ( .A(n24960), .B(n24956), .Z(n25265) );
  XNOR U26788 ( .A(n24955), .B(n24951), .Z(n25266) );
  XNOR U26789 ( .A(n24950), .B(n24946), .Z(n25267) );
  XNOR U26790 ( .A(n24945), .B(n24941), .Z(n25268) );
  XNOR U26791 ( .A(n24940), .B(n24936), .Z(n25269) );
  XNOR U26792 ( .A(n24935), .B(n24931), .Z(n25270) );
  XNOR U26793 ( .A(n24930), .B(n24926), .Z(n25271) );
  XNOR U26794 ( .A(n24925), .B(n24921), .Z(n25272) );
  XOR U26795 ( .A(n25273), .B(n24920), .Z(n24921) );
  AND U26796 ( .A(a[0]), .B(b[59]), .Z(n25273) );
  XOR U26797 ( .A(n25274), .B(n24920), .Z(n24922) );
  XNOR U26798 ( .A(n25275), .B(n25276), .Z(n24920) );
  AND U26799 ( .A(n25277), .B(n25278), .Z(n25275) );
  AND U26800 ( .A(a[1]), .B(b[58]), .Z(n25274) );
  XOR U26801 ( .A(n25279), .B(n24925), .Z(n24927) );
  XOR U26802 ( .A(n25280), .B(n25281), .Z(n24925) );
  AND U26803 ( .A(n25282), .B(n25283), .Z(n25280) );
  AND U26804 ( .A(a[2]), .B(b[57]), .Z(n25279) );
  XOR U26805 ( .A(n25284), .B(n24930), .Z(n24932) );
  XOR U26806 ( .A(n25285), .B(n25286), .Z(n24930) );
  AND U26807 ( .A(n25287), .B(n25288), .Z(n25285) );
  AND U26808 ( .A(a[3]), .B(b[56]), .Z(n25284) );
  XOR U26809 ( .A(n25289), .B(n24935), .Z(n24937) );
  XOR U26810 ( .A(n25290), .B(n25291), .Z(n24935) );
  AND U26811 ( .A(n25292), .B(n25293), .Z(n25290) );
  AND U26812 ( .A(a[4]), .B(b[55]), .Z(n25289) );
  XOR U26813 ( .A(n25294), .B(n24940), .Z(n24942) );
  XOR U26814 ( .A(n25295), .B(n25296), .Z(n24940) );
  AND U26815 ( .A(n25297), .B(n25298), .Z(n25295) );
  AND U26816 ( .A(a[5]), .B(b[54]), .Z(n25294) );
  XOR U26817 ( .A(n25299), .B(n24945), .Z(n24947) );
  XOR U26818 ( .A(n25300), .B(n25301), .Z(n24945) );
  AND U26819 ( .A(n25302), .B(n25303), .Z(n25300) );
  AND U26820 ( .A(a[6]), .B(b[53]), .Z(n25299) );
  XOR U26821 ( .A(n25304), .B(n24950), .Z(n24952) );
  XOR U26822 ( .A(n25305), .B(n25306), .Z(n24950) );
  AND U26823 ( .A(n25307), .B(n25308), .Z(n25305) );
  AND U26824 ( .A(a[7]), .B(b[52]), .Z(n25304) );
  XOR U26825 ( .A(n25309), .B(n24955), .Z(n24957) );
  XOR U26826 ( .A(n25310), .B(n25311), .Z(n24955) );
  AND U26827 ( .A(n25312), .B(n25313), .Z(n25310) );
  AND U26828 ( .A(a[8]), .B(b[51]), .Z(n25309) );
  XOR U26829 ( .A(n25314), .B(n24960), .Z(n24962) );
  XOR U26830 ( .A(n25315), .B(n25316), .Z(n24960) );
  AND U26831 ( .A(n25317), .B(n25318), .Z(n25315) );
  AND U26832 ( .A(a[9]), .B(b[50]), .Z(n25314) );
  XOR U26833 ( .A(n25319), .B(n24965), .Z(n24967) );
  XOR U26834 ( .A(n25320), .B(n25321), .Z(n24965) );
  AND U26835 ( .A(n25322), .B(n25323), .Z(n25320) );
  AND U26836 ( .A(a[10]), .B(b[49]), .Z(n25319) );
  XOR U26837 ( .A(n25324), .B(n24970), .Z(n24972) );
  XOR U26838 ( .A(n25325), .B(n25326), .Z(n24970) );
  AND U26839 ( .A(n25327), .B(n25328), .Z(n25325) );
  AND U26840 ( .A(a[11]), .B(b[48]), .Z(n25324) );
  XOR U26841 ( .A(n25329), .B(n24975), .Z(n24977) );
  XOR U26842 ( .A(n25330), .B(n25331), .Z(n24975) );
  AND U26843 ( .A(n25332), .B(n25333), .Z(n25330) );
  AND U26844 ( .A(a[12]), .B(b[47]), .Z(n25329) );
  XOR U26845 ( .A(n25334), .B(n24980), .Z(n24982) );
  XOR U26846 ( .A(n25335), .B(n25336), .Z(n24980) );
  AND U26847 ( .A(n25337), .B(n25338), .Z(n25335) );
  AND U26848 ( .A(a[13]), .B(b[46]), .Z(n25334) );
  XOR U26849 ( .A(n25339), .B(n24985), .Z(n24987) );
  XOR U26850 ( .A(n25340), .B(n25341), .Z(n24985) );
  AND U26851 ( .A(n25342), .B(n25343), .Z(n25340) );
  AND U26852 ( .A(a[14]), .B(b[45]), .Z(n25339) );
  XOR U26853 ( .A(n25344), .B(n24990), .Z(n24992) );
  XOR U26854 ( .A(n25345), .B(n25346), .Z(n24990) );
  AND U26855 ( .A(n25347), .B(n25348), .Z(n25345) );
  AND U26856 ( .A(a[15]), .B(b[44]), .Z(n25344) );
  XOR U26857 ( .A(n25349), .B(n24995), .Z(n24997) );
  XOR U26858 ( .A(n25350), .B(n25351), .Z(n24995) );
  AND U26859 ( .A(n25352), .B(n25353), .Z(n25350) );
  AND U26860 ( .A(a[16]), .B(b[43]), .Z(n25349) );
  XOR U26861 ( .A(n25354), .B(n25000), .Z(n25002) );
  XOR U26862 ( .A(n25355), .B(n25356), .Z(n25000) );
  AND U26863 ( .A(n25357), .B(n25358), .Z(n25355) );
  AND U26864 ( .A(a[17]), .B(b[42]), .Z(n25354) );
  XOR U26865 ( .A(n25359), .B(n25005), .Z(n25007) );
  XOR U26866 ( .A(n25360), .B(n25361), .Z(n25005) );
  AND U26867 ( .A(n25362), .B(n25363), .Z(n25360) );
  AND U26868 ( .A(a[18]), .B(b[41]), .Z(n25359) );
  XOR U26869 ( .A(n25364), .B(n25010), .Z(n25012) );
  XOR U26870 ( .A(n25365), .B(n25366), .Z(n25010) );
  AND U26871 ( .A(n25367), .B(n25368), .Z(n25365) );
  AND U26872 ( .A(a[19]), .B(b[40]), .Z(n25364) );
  XOR U26873 ( .A(n25369), .B(n25015), .Z(n25017) );
  XOR U26874 ( .A(n25370), .B(n25371), .Z(n25015) );
  AND U26875 ( .A(n25372), .B(n25373), .Z(n25370) );
  AND U26876 ( .A(a[20]), .B(b[39]), .Z(n25369) );
  XOR U26877 ( .A(n25374), .B(n25020), .Z(n25022) );
  XOR U26878 ( .A(n25375), .B(n25376), .Z(n25020) );
  AND U26879 ( .A(n25377), .B(n25378), .Z(n25375) );
  AND U26880 ( .A(a[21]), .B(b[38]), .Z(n25374) );
  XOR U26881 ( .A(n25379), .B(n25025), .Z(n25027) );
  XOR U26882 ( .A(n25380), .B(n25381), .Z(n25025) );
  AND U26883 ( .A(n25382), .B(n25383), .Z(n25380) );
  AND U26884 ( .A(a[22]), .B(b[37]), .Z(n25379) );
  XOR U26885 ( .A(n25384), .B(n25030), .Z(n25032) );
  XOR U26886 ( .A(n25385), .B(n25386), .Z(n25030) );
  AND U26887 ( .A(n25387), .B(n25388), .Z(n25385) );
  AND U26888 ( .A(a[23]), .B(b[36]), .Z(n25384) );
  XOR U26889 ( .A(n25389), .B(n25035), .Z(n25037) );
  XOR U26890 ( .A(n25390), .B(n25391), .Z(n25035) );
  AND U26891 ( .A(n25392), .B(n25393), .Z(n25390) );
  AND U26892 ( .A(a[24]), .B(b[35]), .Z(n25389) );
  XOR U26893 ( .A(n25394), .B(n25040), .Z(n25042) );
  XOR U26894 ( .A(n25395), .B(n25396), .Z(n25040) );
  AND U26895 ( .A(n25397), .B(n25398), .Z(n25395) );
  AND U26896 ( .A(a[25]), .B(b[34]), .Z(n25394) );
  XOR U26897 ( .A(n25399), .B(n25045), .Z(n25047) );
  XOR U26898 ( .A(n25400), .B(n25401), .Z(n25045) );
  AND U26899 ( .A(n25402), .B(n25403), .Z(n25400) );
  AND U26900 ( .A(a[26]), .B(b[33]), .Z(n25399) );
  XOR U26901 ( .A(n25404), .B(n25050), .Z(n25052) );
  XOR U26902 ( .A(n25405), .B(n25406), .Z(n25050) );
  AND U26903 ( .A(n25407), .B(n25408), .Z(n25405) );
  AND U26904 ( .A(a[27]), .B(b[32]), .Z(n25404) );
  XOR U26905 ( .A(n25409), .B(n25055), .Z(n25057) );
  XOR U26906 ( .A(n25410), .B(n25411), .Z(n25055) );
  AND U26907 ( .A(n25412), .B(n25413), .Z(n25410) );
  AND U26908 ( .A(a[28]), .B(b[31]), .Z(n25409) );
  XOR U26909 ( .A(n25414), .B(n25060), .Z(n25062) );
  XOR U26910 ( .A(n25415), .B(n25416), .Z(n25060) );
  AND U26911 ( .A(n25417), .B(n25418), .Z(n25415) );
  AND U26912 ( .A(a[29]), .B(b[30]), .Z(n25414) );
  XOR U26913 ( .A(n25419), .B(n25065), .Z(n25067) );
  XOR U26914 ( .A(n25420), .B(n25421), .Z(n25065) );
  AND U26915 ( .A(n25422), .B(n25423), .Z(n25420) );
  AND U26916 ( .A(b[29]), .B(a[30]), .Z(n25419) );
  XOR U26917 ( .A(n25424), .B(n25070), .Z(n25072) );
  XOR U26918 ( .A(n25425), .B(n25426), .Z(n25070) );
  AND U26919 ( .A(n25427), .B(n25428), .Z(n25425) );
  AND U26920 ( .A(b[28]), .B(a[31]), .Z(n25424) );
  XOR U26921 ( .A(n25429), .B(n25075), .Z(n25077) );
  XOR U26922 ( .A(n25430), .B(n25431), .Z(n25075) );
  AND U26923 ( .A(n25432), .B(n25433), .Z(n25430) );
  AND U26924 ( .A(b[27]), .B(a[32]), .Z(n25429) );
  XOR U26925 ( .A(n25434), .B(n25080), .Z(n25082) );
  XOR U26926 ( .A(n25435), .B(n25436), .Z(n25080) );
  AND U26927 ( .A(n25437), .B(n25438), .Z(n25435) );
  AND U26928 ( .A(b[26]), .B(a[33]), .Z(n25434) );
  XOR U26929 ( .A(n25439), .B(n25085), .Z(n25087) );
  XOR U26930 ( .A(n25440), .B(n25441), .Z(n25085) );
  AND U26931 ( .A(n25442), .B(n25443), .Z(n25440) );
  AND U26932 ( .A(b[25]), .B(a[34]), .Z(n25439) );
  XOR U26933 ( .A(n25444), .B(n25090), .Z(n25092) );
  XOR U26934 ( .A(n25445), .B(n25446), .Z(n25090) );
  AND U26935 ( .A(n25447), .B(n25448), .Z(n25445) );
  AND U26936 ( .A(b[24]), .B(a[35]), .Z(n25444) );
  XOR U26937 ( .A(n25449), .B(n25095), .Z(n25097) );
  XOR U26938 ( .A(n25450), .B(n25451), .Z(n25095) );
  AND U26939 ( .A(n25452), .B(n25453), .Z(n25450) );
  AND U26940 ( .A(b[23]), .B(a[36]), .Z(n25449) );
  XOR U26941 ( .A(n25454), .B(n25100), .Z(n25102) );
  XOR U26942 ( .A(n25455), .B(n25456), .Z(n25100) );
  AND U26943 ( .A(n25457), .B(n25458), .Z(n25455) );
  AND U26944 ( .A(b[22]), .B(a[37]), .Z(n25454) );
  XOR U26945 ( .A(n25459), .B(n25105), .Z(n25107) );
  XOR U26946 ( .A(n25460), .B(n25461), .Z(n25105) );
  AND U26947 ( .A(n25462), .B(n25463), .Z(n25460) );
  AND U26948 ( .A(b[21]), .B(a[38]), .Z(n25459) );
  XOR U26949 ( .A(n25464), .B(n25110), .Z(n25112) );
  XOR U26950 ( .A(n25465), .B(n25466), .Z(n25110) );
  AND U26951 ( .A(n25467), .B(n25468), .Z(n25465) );
  AND U26952 ( .A(b[20]), .B(a[39]), .Z(n25464) );
  XOR U26953 ( .A(n25469), .B(n25115), .Z(n25117) );
  XOR U26954 ( .A(n25470), .B(n25471), .Z(n25115) );
  AND U26955 ( .A(n25472), .B(n25473), .Z(n25470) );
  AND U26956 ( .A(b[19]), .B(a[40]), .Z(n25469) );
  XOR U26957 ( .A(n25474), .B(n25120), .Z(n25122) );
  XOR U26958 ( .A(n25475), .B(n25476), .Z(n25120) );
  AND U26959 ( .A(n25477), .B(n25478), .Z(n25475) );
  AND U26960 ( .A(b[18]), .B(a[41]), .Z(n25474) );
  XOR U26961 ( .A(n25479), .B(n25125), .Z(n25127) );
  XOR U26962 ( .A(n25480), .B(n25481), .Z(n25125) );
  AND U26963 ( .A(n25482), .B(n25483), .Z(n25480) );
  AND U26964 ( .A(b[17]), .B(a[42]), .Z(n25479) );
  XOR U26965 ( .A(n25484), .B(n25130), .Z(n25132) );
  XOR U26966 ( .A(n25485), .B(n25486), .Z(n25130) );
  AND U26967 ( .A(n25487), .B(n25488), .Z(n25485) );
  AND U26968 ( .A(b[16]), .B(a[43]), .Z(n25484) );
  XOR U26969 ( .A(n25489), .B(n25135), .Z(n25137) );
  XOR U26970 ( .A(n25490), .B(n25491), .Z(n25135) );
  AND U26971 ( .A(n25492), .B(n25493), .Z(n25490) );
  AND U26972 ( .A(b[15]), .B(a[44]), .Z(n25489) );
  XOR U26973 ( .A(n25494), .B(n25140), .Z(n25142) );
  XOR U26974 ( .A(n25495), .B(n25496), .Z(n25140) );
  AND U26975 ( .A(n25497), .B(n25498), .Z(n25495) );
  AND U26976 ( .A(b[14]), .B(a[45]), .Z(n25494) );
  XOR U26977 ( .A(n25499), .B(n25145), .Z(n25147) );
  XOR U26978 ( .A(n25500), .B(n25501), .Z(n25145) );
  AND U26979 ( .A(n25502), .B(n25503), .Z(n25500) );
  AND U26980 ( .A(b[13]), .B(a[46]), .Z(n25499) );
  XOR U26981 ( .A(n25504), .B(n25150), .Z(n25152) );
  XOR U26982 ( .A(n25505), .B(n25506), .Z(n25150) );
  AND U26983 ( .A(n25507), .B(n25508), .Z(n25505) );
  AND U26984 ( .A(b[12]), .B(a[47]), .Z(n25504) );
  XOR U26985 ( .A(n25509), .B(n25155), .Z(n25157) );
  XOR U26986 ( .A(n25510), .B(n25511), .Z(n25155) );
  AND U26987 ( .A(n25512), .B(n25513), .Z(n25510) );
  AND U26988 ( .A(b[11]), .B(a[48]), .Z(n25509) );
  XOR U26989 ( .A(n25514), .B(n25160), .Z(n25162) );
  XOR U26990 ( .A(n25515), .B(n25516), .Z(n25160) );
  AND U26991 ( .A(n25517), .B(n25518), .Z(n25515) );
  AND U26992 ( .A(b[10]), .B(a[49]), .Z(n25514) );
  XOR U26993 ( .A(n25519), .B(n25165), .Z(n25167) );
  XOR U26994 ( .A(n25520), .B(n25521), .Z(n25165) );
  AND U26995 ( .A(n25522), .B(n25523), .Z(n25520) );
  AND U26996 ( .A(b[9]), .B(a[50]), .Z(n25519) );
  XOR U26997 ( .A(n25524), .B(n25170), .Z(n25172) );
  XOR U26998 ( .A(n25525), .B(n25526), .Z(n25170) );
  AND U26999 ( .A(n25527), .B(n25528), .Z(n25525) );
  AND U27000 ( .A(b[8]), .B(a[51]), .Z(n25524) );
  XOR U27001 ( .A(n25529), .B(n25175), .Z(n25177) );
  XOR U27002 ( .A(n25530), .B(n25531), .Z(n25175) );
  AND U27003 ( .A(n25532), .B(n25533), .Z(n25530) );
  AND U27004 ( .A(b[7]), .B(a[52]), .Z(n25529) );
  XOR U27005 ( .A(n25534), .B(n25180), .Z(n25182) );
  XOR U27006 ( .A(n25535), .B(n25536), .Z(n25180) );
  AND U27007 ( .A(n25537), .B(n25538), .Z(n25535) );
  AND U27008 ( .A(b[6]), .B(a[53]), .Z(n25534) );
  XOR U27009 ( .A(n25539), .B(n25185), .Z(n25187) );
  XOR U27010 ( .A(n25540), .B(n25541), .Z(n25185) );
  AND U27011 ( .A(n25542), .B(n25543), .Z(n25540) );
  AND U27012 ( .A(b[5]), .B(a[54]), .Z(n25539) );
  XOR U27013 ( .A(n25544), .B(n25190), .Z(n25192) );
  XOR U27014 ( .A(n25545), .B(n25546), .Z(n25190) );
  AND U27015 ( .A(n25547), .B(n25548), .Z(n25545) );
  AND U27016 ( .A(b[4]), .B(a[55]), .Z(n25544) );
  XNOR U27017 ( .A(n25549), .B(n25550), .Z(n25204) );
  NANDN U27018 ( .A(n25551), .B(n25552), .Z(n25550) );
  XOR U27019 ( .A(n25553), .B(n25195), .Z(n25197) );
  XNOR U27020 ( .A(n25554), .B(n25555), .Z(n25195) );
  AND U27021 ( .A(n25556), .B(n25557), .Z(n25554) );
  AND U27022 ( .A(b[3]), .B(a[56]), .Z(n25553) );
  XOR U27023 ( .A(n25211), .B(n25210), .Z(c[122]) );
  XOR U27024 ( .A(sreg[186]), .B(n25209), .Z(n25210) );
  XOR U27025 ( .A(n25216), .B(n25558), .Z(n25211) );
  XNOR U27026 ( .A(n25215), .B(n25209), .Z(n25558) );
  XOR U27027 ( .A(n25559), .B(n25560), .Z(n25209) );
  NOR U27028 ( .A(n25561), .B(n25562), .Z(n25559) );
  NAND U27029 ( .A(a[58]), .B(b[0]), .Z(n25215) );
  XNOR U27030 ( .A(n25551), .B(n25552), .Z(n25216) );
  XOR U27031 ( .A(n25549), .B(n25563), .Z(n25552) );
  NAND U27032 ( .A(b[1]), .B(a[57]), .Z(n25563) );
  XOR U27033 ( .A(n25557), .B(n25564), .Z(n25551) );
  XOR U27034 ( .A(n25549), .B(n25556), .Z(n25564) );
  XNOR U27035 ( .A(n25565), .B(n25555), .Z(n25556) );
  AND U27036 ( .A(b[2]), .B(a[56]), .Z(n25565) );
  NANDN U27037 ( .A(n25566), .B(n25567), .Z(n25549) );
  XOR U27038 ( .A(n25555), .B(n25547), .Z(n25568) );
  XNOR U27039 ( .A(n25546), .B(n25542), .Z(n25569) );
  XNOR U27040 ( .A(n25541), .B(n25537), .Z(n25570) );
  XNOR U27041 ( .A(n25536), .B(n25532), .Z(n25571) );
  XNOR U27042 ( .A(n25531), .B(n25527), .Z(n25572) );
  XNOR U27043 ( .A(n25526), .B(n25522), .Z(n25573) );
  XNOR U27044 ( .A(n25521), .B(n25517), .Z(n25574) );
  XNOR U27045 ( .A(n25516), .B(n25512), .Z(n25575) );
  XNOR U27046 ( .A(n25511), .B(n25507), .Z(n25576) );
  XNOR U27047 ( .A(n25506), .B(n25502), .Z(n25577) );
  XNOR U27048 ( .A(n25501), .B(n25497), .Z(n25578) );
  XNOR U27049 ( .A(n25496), .B(n25492), .Z(n25579) );
  XNOR U27050 ( .A(n25491), .B(n25487), .Z(n25580) );
  XNOR U27051 ( .A(n25486), .B(n25482), .Z(n25581) );
  XNOR U27052 ( .A(n25481), .B(n25477), .Z(n25582) );
  XNOR U27053 ( .A(n25476), .B(n25472), .Z(n25583) );
  XNOR U27054 ( .A(n25471), .B(n25467), .Z(n25584) );
  XNOR U27055 ( .A(n25466), .B(n25462), .Z(n25585) );
  XNOR U27056 ( .A(n25461), .B(n25457), .Z(n25586) );
  XNOR U27057 ( .A(n25456), .B(n25452), .Z(n25587) );
  XNOR U27058 ( .A(n25451), .B(n25447), .Z(n25588) );
  XNOR U27059 ( .A(n25446), .B(n25442), .Z(n25589) );
  XNOR U27060 ( .A(n25441), .B(n25437), .Z(n25590) );
  XNOR U27061 ( .A(n25436), .B(n25432), .Z(n25591) );
  XNOR U27062 ( .A(n25431), .B(n25427), .Z(n25592) );
  XNOR U27063 ( .A(n25426), .B(n25422), .Z(n25593) );
  XNOR U27064 ( .A(n25421), .B(n25417), .Z(n25594) );
  XNOR U27065 ( .A(n25416), .B(n25412), .Z(n25595) );
  XNOR U27066 ( .A(n25411), .B(n25407), .Z(n25596) );
  XNOR U27067 ( .A(n25406), .B(n25402), .Z(n25597) );
  XNOR U27068 ( .A(n25401), .B(n25397), .Z(n25598) );
  XNOR U27069 ( .A(n25396), .B(n25392), .Z(n25599) );
  XNOR U27070 ( .A(n25391), .B(n25387), .Z(n25600) );
  XNOR U27071 ( .A(n25386), .B(n25382), .Z(n25601) );
  XNOR U27072 ( .A(n25381), .B(n25377), .Z(n25602) );
  XNOR U27073 ( .A(n25376), .B(n25372), .Z(n25603) );
  XNOR U27074 ( .A(n25371), .B(n25367), .Z(n25604) );
  XNOR U27075 ( .A(n25366), .B(n25362), .Z(n25605) );
  XNOR U27076 ( .A(n25361), .B(n25357), .Z(n25606) );
  XNOR U27077 ( .A(n25356), .B(n25352), .Z(n25607) );
  XNOR U27078 ( .A(n25351), .B(n25347), .Z(n25608) );
  XNOR U27079 ( .A(n25346), .B(n25342), .Z(n25609) );
  XNOR U27080 ( .A(n25341), .B(n25337), .Z(n25610) );
  XNOR U27081 ( .A(n25336), .B(n25332), .Z(n25611) );
  XNOR U27082 ( .A(n25331), .B(n25327), .Z(n25612) );
  XNOR U27083 ( .A(n25326), .B(n25322), .Z(n25613) );
  XNOR U27084 ( .A(n25321), .B(n25317), .Z(n25614) );
  XNOR U27085 ( .A(n25316), .B(n25312), .Z(n25615) );
  XNOR U27086 ( .A(n25311), .B(n25307), .Z(n25616) );
  XNOR U27087 ( .A(n25306), .B(n25302), .Z(n25617) );
  XNOR U27088 ( .A(n25301), .B(n25297), .Z(n25618) );
  XNOR U27089 ( .A(n25296), .B(n25292), .Z(n25619) );
  XNOR U27090 ( .A(n25291), .B(n25287), .Z(n25620) );
  XNOR U27091 ( .A(n25286), .B(n25282), .Z(n25621) );
  XNOR U27092 ( .A(n25281), .B(n25277), .Z(n25622) );
  XNOR U27093 ( .A(n25623), .B(n25276), .Z(n25277) );
  AND U27094 ( .A(a[0]), .B(b[58]), .Z(n25623) );
  XNOR U27095 ( .A(n25624), .B(n25276), .Z(n25278) );
  XNOR U27096 ( .A(n25625), .B(n25626), .Z(n25276) );
  AND U27097 ( .A(n25627), .B(n25628), .Z(n25625) );
  AND U27098 ( .A(a[1]), .B(b[57]), .Z(n25624) );
  XOR U27099 ( .A(n25629), .B(n25281), .Z(n25283) );
  XOR U27100 ( .A(n25630), .B(n25631), .Z(n25281) );
  AND U27101 ( .A(n25632), .B(n25633), .Z(n25630) );
  AND U27102 ( .A(a[2]), .B(b[56]), .Z(n25629) );
  XOR U27103 ( .A(n25634), .B(n25286), .Z(n25288) );
  XOR U27104 ( .A(n25635), .B(n25636), .Z(n25286) );
  AND U27105 ( .A(n25637), .B(n25638), .Z(n25635) );
  AND U27106 ( .A(a[3]), .B(b[55]), .Z(n25634) );
  XOR U27107 ( .A(n25639), .B(n25291), .Z(n25293) );
  XOR U27108 ( .A(n25640), .B(n25641), .Z(n25291) );
  AND U27109 ( .A(n25642), .B(n25643), .Z(n25640) );
  AND U27110 ( .A(a[4]), .B(b[54]), .Z(n25639) );
  XOR U27111 ( .A(n25644), .B(n25296), .Z(n25298) );
  XOR U27112 ( .A(n25645), .B(n25646), .Z(n25296) );
  AND U27113 ( .A(n25647), .B(n25648), .Z(n25645) );
  AND U27114 ( .A(a[5]), .B(b[53]), .Z(n25644) );
  XOR U27115 ( .A(n25649), .B(n25301), .Z(n25303) );
  XOR U27116 ( .A(n25650), .B(n25651), .Z(n25301) );
  AND U27117 ( .A(n25652), .B(n25653), .Z(n25650) );
  AND U27118 ( .A(a[6]), .B(b[52]), .Z(n25649) );
  XOR U27119 ( .A(n25654), .B(n25306), .Z(n25308) );
  XOR U27120 ( .A(n25655), .B(n25656), .Z(n25306) );
  AND U27121 ( .A(n25657), .B(n25658), .Z(n25655) );
  AND U27122 ( .A(a[7]), .B(b[51]), .Z(n25654) );
  XOR U27123 ( .A(n25659), .B(n25311), .Z(n25313) );
  XOR U27124 ( .A(n25660), .B(n25661), .Z(n25311) );
  AND U27125 ( .A(n25662), .B(n25663), .Z(n25660) );
  AND U27126 ( .A(a[8]), .B(b[50]), .Z(n25659) );
  XOR U27127 ( .A(n25664), .B(n25316), .Z(n25318) );
  XOR U27128 ( .A(n25665), .B(n25666), .Z(n25316) );
  AND U27129 ( .A(n25667), .B(n25668), .Z(n25665) );
  AND U27130 ( .A(a[9]), .B(b[49]), .Z(n25664) );
  XOR U27131 ( .A(n25669), .B(n25321), .Z(n25323) );
  XOR U27132 ( .A(n25670), .B(n25671), .Z(n25321) );
  AND U27133 ( .A(n25672), .B(n25673), .Z(n25670) );
  AND U27134 ( .A(a[10]), .B(b[48]), .Z(n25669) );
  XOR U27135 ( .A(n25674), .B(n25326), .Z(n25328) );
  XOR U27136 ( .A(n25675), .B(n25676), .Z(n25326) );
  AND U27137 ( .A(n25677), .B(n25678), .Z(n25675) );
  AND U27138 ( .A(a[11]), .B(b[47]), .Z(n25674) );
  XOR U27139 ( .A(n25679), .B(n25331), .Z(n25333) );
  XOR U27140 ( .A(n25680), .B(n25681), .Z(n25331) );
  AND U27141 ( .A(n25682), .B(n25683), .Z(n25680) );
  AND U27142 ( .A(a[12]), .B(b[46]), .Z(n25679) );
  XOR U27143 ( .A(n25684), .B(n25336), .Z(n25338) );
  XOR U27144 ( .A(n25685), .B(n25686), .Z(n25336) );
  AND U27145 ( .A(n25687), .B(n25688), .Z(n25685) );
  AND U27146 ( .A(a[13]), .B(b[45]), .Z(n25684) );
  XOR U27147 ( .A(n25689), .B(n25341), .Z(n25343) );
  XOR U27148 ( .A(n25690), .B(n25691), .Z(n25341) );
  AND U27149 ( .A(n25692), .B(n25693), .Z(n25690) );
  AND U27150 ( .A(a[14]), .B(b[44]), .Z(n25689) );
  XOR U27151 ( .A(n25694), .B(n25346), .Z(n25348) );
  XOR U27152 ( .A(n25695), .B(n25696), .Z(n25346) );
  AND U27153 ( .A(n25697), .B(n25698), .Z(n25695) );
  AND U27154 ( .A(a[15]), .B(b[43]), .Z(n25694) );
  XOR U27155 ( .A(n25699), .B(n25351), .Z(n25353) );
  XOR U27156 ( .A(n25700), .B(n25701), .Z(n25351) );
  AND U27157 ( .A(n25702), .B(n25703), .Z(n25700) );
  AND U27158 ( .A(a[16]), .B(b[42]), .Z(n25699) );
  XOR U27159 ( .A(n25704), .B(n25356), .Z(n25358) );
  XOR U27160 ( .A(n25705), .B(n25706), .Z(n25356) );
  AND U27161 ( .A(n25707), .B(n25708), .Z(n25705) );
  AND U27162 ( .A(a[17]), .B(b[41]), .Z(n25704) );
  XOR U27163 ( .A(n25709), .B(n25361), .Z(n25363) );
  XOR U27164 ( .A(n25710), .B(n25711), .Z(n25361) );
  AND U27165 ( .A(n25712), .B(n25713), .Z(n25710) );
  AND U27166 ( .A(a[18]), .B(b[40]), .Z(n25709) );
  XOR U27167 ( .A(n25714), .B(n25366), .Z(n25368) );
  XOR U27168 ( .A(n25715), .B(n25716), .Z(n25366) );
  AND U27169 ( .A(n25717), .B(n25718), .Z(n25715) );
  AND U27170 ( .A(a[19]), .B(b[39]), .Z(n25714) );
  XOR U27171 ( .A(n25719), .B(n25371), .Z(n25373) );
  XOR U27172 ( .A(n25720), .B(n25721), .Z(n25371) );
  AND U27173 ( .A(n25722), .B(n25723), .Z(n25720) );
  AND U27174 ( .A(a[20]), .B(b[38]), .Z(n25719) );
  XOR U27175 ( .A(n25724), .B(n25376), .Z(n25378) );
  XOR U27176 ( .A(n25725), .B(n25726), .Z(n25376) );
  AND U27177 ( .A(n25727), .B(n25728), .Z(n25725) );
  AND U27178 ( .A(a[21]), .B(b[37]), .Z(n25724) );
  XOR U27179 ( .A(n25729), .B(n25381), .Z(n25383) );
  XOR U27180 ( .A(n25730), .B(n25731), .Z(n25381) );
  AND U27181 ( .A(n25732), .B(n25733), .Z(n25730) );
  AND U27182 ( .A(a[22]), .B(b[36]), .Z(n25729) );
  XOR U27183 ( .A(n25734), .B(n25386), .Z(n25388) );
  XOR U27184 ( .A(n25735), .B(n25736), .Z(n25386) );
  AND U27185 ( .A(n25737), .B(n25738), .Z(n25735) );
  AND U27186 ( .A(a[23]), .B(b[35]), .Z(n25734) );
  XOR U27187 ( .A(n25739), .B(n25391), .Z(n25393) );
  XOR U27188 ( .A(n25740), .B(n25741), .Z(n25391) );
  AND U27189 ( .A(n25742), .B(n25743), .Z(n25740) );
  AND U27190 ( .A(a[24]), .B(b[34]), .Z(n25739) );
  XOR U27191 ( .A(n25744), .B(n25396), .Z(n25398) );
  XOR U27192 ( .A(n25745), .B(n25746), .Z(n25396) );
  AND U27193 ( .A(n25747), .B(n25748), .Z(n25745) );
  AND U27194 ( .A(a[25]), .B(b[33]), .Z(n25744) );
  XOR U27195 ( .A(n25749), .B(n25401), .Z(n25403) );
  XOR U27196 ( .A(n25750), .B(n25751), .Z(n25401) );
  AND U27197 ( .A(n25752), .B(n25753), .Z(n25750) );
  AND U27198 ( .A(a[26]), .B(b[32]), .Z(n25749) );
  XOR U27199 ( .A(n25754), .B(n25406), .Z(n25408) );
  XOR U27200 ( .A(n25755), .B(n25756), .Z(n25406) );
  AND U27201 ( .A(n25757), .B(n25758), .Z(n25755) );
  AND U27202 ( .A(a[27]), .B(b[31]), .Z(n25754) );
  XOR U27203 ( .A(n25759), .B(n25411), .Z(n25413) );
  XOR U27204 ( .A(n25760), .B(n25761), .Z(n25411) );
  AND U27205 ( .A(n25762), .B(n25763), .Z(n25760) );
  AND U27206 ( .A(a[28]), .B(b[30]), .Z(n25759) );
  XOR U27207 ( .A(n25764), .B(n25416), .Z(n25418) );
  XOR U27208 ( .A(n25765), .B(n25766), .Z(n25416) );
  AND U27209 ( .A(n25767), .B(n25768), .Z(n25765) );
  AND U27210 ( .A(a[29]), .B(b[29]), .Z(n25764) );
  XOR U27211 ( .A(n25769), .B(n25421), .Z(n25423) );
  XOR U27212 ( .A(n25770), .B(n25771), .Z(n25421) );
  AND U27213 ( .A(n25772), .B(n25773), .Z(n25770) );
  AND U27214 ( .A(b[28]), .B(a[30]), .Z(n25769) );
  XOR U27215 ( .A(n25774), .B(n25426), .Z(n25428) );
  XOR U27216 ( .A(n25775), .B(n25776), .Z(n25426) );
  AND U27217 ( .A(n25777), .B(n25778), .Z(n25775) );
  AND U27218 ( .A(b[27]), .B(a[31]), .Z(n25774) );
  XOR U27219 ( .A(n25779), .B(n25431), .Z(n25433) );
  XOR U27220 ( .A(n25780), .B(n25781), .Z(n25431) );
  AND U27221 ( .A(n25782), .B(n25783), .Z(n25780) );
  AND U27222 ( .A(b[26]), .B(a[32]), .Z(n25779) );
  XOR U27223 ( .A(n25784), .B(n25436), .Z(n25438) );
  XOR U27224 ( .A(n25785), .B(n25786), .Z(n25436) );
  AND U27225 ( .A(n25787), .B(n25788), .Z(n25785) );
  AND U27226 ( .A(b[25]), .B(a[33]), .Z(n25784) );
  XOR U27227 ( .A(n25789), .B(n25441), .Z(n25443) );
  XOR U27228 ( .A(n25790), .B(n25791), .Z(n25441) );
  AND U27229 ( .A(n25792), .B(n25793), .Z(n25790) );
  AND U27230 ( .A(b[24]), .B(a[34]), .Z(n25789) );
  XOR U27231 ( .A(n25794), .B(n25446), .Z(n25448) );
  XOR U27232 ( .A(n25795), .B(n25796), .Z(n25446) );
  AND U27233 ( .A(n25797), .B(n25798), .Z(n25795) );
  AND U27234 ( .A(b[23]), .B(a[35]), .Z(n25794) );
  XOR U27235 ( .A(n25799), .B(n25451), .Z(n25453) );
  XOR U27236 ( .A(n25800), .B(n25801), .Z(n25451) );
  AND U27237 ( .A(n25802), .B(n25803), .Z(n25800) );
  AND U27238 ( .A(b[22]), .B(a[36]), .Z(n25799) );
  XOR U27239 ( .A(n25804), .B(n25456), .Z(n25458) );
  XOR U27240 ( .A(n25805), .B(n25806), .Z(n25456) );
  AND U27241 ( .A(n25807), .B(n25808), .Z(n25805) );
  AND U27242 ( .A(b[21]), .B(a[37]), .Z(n25804) );
  XOR U27243 ( .A(n25809), .B(n25461), .Z(n25463) );
  XOR U27244 ( .A(n25810), .B(n25811), .Z(n25461) );
  AND U27245 ( .A(n25812), .B(n25813), .Z(n25810) );
  AND U27246 ( .A(b[20]), .B(a[38]), .Z(n25809) );
  XOR U27247 ( .A(n25814), .B(n25466), .Z(n25468) );
  XOR U27248 ( .A(n25815), .B(n25816), .Z(n25466) );
  AND U27249 ( .A(n25817), .B(n25818), .Z(n25815) );
  AND U27250 ( .A(b[19]), .B(a[39]), .Z(n25814) );
  XOR U27251 ( .A(n25819), .B(n25471), .Z(n25473) );
  XOR U27252 ( .A(n25820), .B(n25821), .Z(n25471) );
  AND U27253 ( .A(n25822), .B(n25823), .Z(n25820) );
  AND U27254 ( .A(b[18]), .B(a[40]), .Z(n25819) );
  XOR U27255 ( .A(n25824), .B(n25476), .Z(n25478) );
  XOR U27256 ( .A(n25825), .B(n25826), .Z(n25476) );
  AND U27257 ( .A(n25827), .B(n25828), .Z(n25825) );
  AND U27258 ( .A(b[17]), .B(a[41]), .Z(n25824) );
  XOR U27259 ( .A(n25829), .B(n25481), .Z(n25483) );
  XOR U27260 ( .A(n25830), .B(n25831), .Z(n25481) );
  AND U27261 ( .A(n25832), .B(n25833), .Z(n25830) );
  AND U27262 ( .A(b[16]), .B(a[42]), .Z(n25829) );
  XOR U27263 ( .A(n25834), .B(n25486), .Z(n25488) );
  XOR U27264 ( .A(n25835), .B(n25836), .Z(n25486) );
  AND U27265 ( .A(n25837), .B(n25838), .Z(n25835) );
  AND U27266 ( .A(b[15]), .B(a[43]), .Z(n25834) );
  XOR U27267 ( .A(n25839), .B(n25491), .Z(n25493) );
  XOR U27268 ( .A(n25840), .B(n25841), .Z(n25491) );
  AND U27269 ( .A(n25842), .B(n25843), .Z(n25840) );
  AND U27270 ( .A(b[14]), .B(a[44]), .Z(n25839) );
  XOR U27271 ( .A(n25844), .B(n25496), .Z(n25498) );
  XOR U27272 ( .A(n25845), .B(n25846), .Z(n25496) );
  AND U27273 ( .A(n25847), .B(n25848), .Z(n25845) );
  AND U27274 ( .A(b[13]), .B(a[45]), .Z(n25844) );
  XOR U27275 ( .A(n25849), .B(n25501), .Z(n25503) );
  XOR U27276 ( .A(n25850), .B(n25851), .Z(n25501) );
  AND U27277 ( .A(n25852), .B(n25853), .Z(n25850) );
  AND U27278 ( .A(b[12]), .B(a[46]), .Z(n25849) );
  XOR U27279 ( .A(n25854), .B(n25506), .Z(n25508) );
  XOR U27280 ( .A(n25855), .B(n25856), .Z(n25506) );
  AND U27281 ( .A(n25857), .B(n25858), .Z(n25855) );
  AND U27282 ( .A(b[11]), .B(a[47]), .Z(n25854) );
  XOR U27283 ( .A(n25859), .B(n25511), .Z(n25513) );
  XOR U27284 ( .A(n25860), .B(n25861), .Z(n25511) );
  AND U27285 ( .A(n25862), .B(n25863), .Z(n25860) );
  AND U27286 ( .A(b[10]), .B(a[48]), .Z(n25859) );
  XOR U27287 ( .A(n25864), .B(n25516), .Z(n25518) );
  XOR U27288 ( .A(n25865), .B(n25866), .Z(n25516) );
  AND U27289 ( .A(n25867), .B(n25868), .Z(n25865) );
  AND U27290 ( .A(b[9]), .B(a[49]), .Z(n25864) );
  XOR U27291 ( .A(n25869), .B(n25521), .Z(n25523) );
  XOR U27292 ( .A(n25870), .B(n25871), .Z(n25521) );
  AND U27293 ( .A(n25872), .B(n25873), .Z(n25870) );
  AND U27294 ( .A(b[8]), .B(a[50]), .Z(n25869) );
  XOR U27295 ( .A(n25874), .B(n25526), .Z(n25528) );
  XOR U27296 ( .A(n25875), .B(n25876), .Z(n25526) );
  AND U27297 ( .A(n25877), .B(n25878), .Z(n25875) );
  AND U27298 ( .A(b[7]), .B(a[51]), .Z(n25874) );
  XOR U27299 ( .A(n25879), .B(n25531), .Z(n25533) );
  XOR U27300 ( .A(n25880), .B(n25881), .Z(n25531) );
  AND U27301 ( .A(n25882), .B(n25883), .Z(n25880) );
  AND U27302 ( .A(b[6]), .B(a[52]), .Z(n25879) );
  XOR U27303 ( .A(n25884), .B(n25536), .Z(n25538) );
  XOR U27304 ( .A(n25885), .B(n25886), .Z(n25536) );
  AND U27305 ( .A(n25887), .B(n25888), .Z(n25885) );
  AND U27306 ( .A(b[5]), .B(a[53]), .Z(n25884) );
  XOR U27307 ( .A(n25889), .B(n25541), .Z(n25543) );
  XOR U27308 ( .A(n25890), .B(n25891), .Z(n25541) );
  AND U27309 ( .A(n25892), .B(n25893), .Z(n25890) );
  AND U27310 ( .A(b[4]), .B(a[54]), .Z(n25889) );
  XNOR U27311 ( .A(n25894), .B(n25895), .Z(n25555) );
  NANDN U27312 ( .A(n25896), .B(n25897), .Z(n25895) );
  XOR U27313 ( .A(n25898), .B(n25546), .Z(n25548) );
  XNOR U27314 ( .A(n25899), .B(n25900), .Z(n25546) );
  AND U27315 ( .A(n25901), .B(n25902), .Z(n25899) );
  AND U27316 ( .A(b[3]), .B(a[55]), .Z(n25898) );
  XOR U27317 ( .A(n25562), .B(n25561), .Z(c[121]) );
  XOR U27318 ( .A(sreg[185]), .B(n25560), .Z(n25561) );
  XOR U27319 ( .A(n25567), .B(n25903), .Z(n25562) );
  XNOR U27320 ( .A(n25566), .B(n25560), .Z(n25903) );
  XOR U27321 ( .A(n25904), .B(n25905), .Z(n25560) );
  NOR U27322 ( .A(n25906), .B(n25907), .Z(n25904) );
  NAND U27323 ( .A(a[57]), .B(b[0]), .Z(n25566) );
  XNOR U27324 ( .A(n25896), .B(n25897), .Z(n25567) );
  XOR U27325 ( .A(n25894), .B(n25908), .Z(n25897) );
  NAND U27326 ( .A(b[1]), .B(a[56]), .Z(n25908) );
  XOR U27327 ( .A(n25902), .B(n25909), .Z(n25896) );
  XOR U27328 ( .A(n25894), .B(n25901), .Z(n25909) );
  XNOR U27329 ( .A(n25910), .B(n25900), .Z(n25901) );
  AND U27330 ( .A(b[2]), .B(a[55]), .Z(n25910) );
  NANDN U27331 ( .A(n25911), .B(n25912), .Z(n25894) );
  XOR U27332 ( .A(n25900), .B(n25892), .Z(n25913) );
  XNOR U27333 ( .A(n25891), .B(n25887), .Z(n25914) );
  XNOR U27334 ( .A(n25886), .B(n25882), .Z(n25915) );
  XNOR U27335 ( .A(n25881), .B(n25877), .Z(n25916) );
  XNOR U27336 ( .A(n25876), .B(n25872), .Z(n25917) );
  XNOR U27337 ( .A(n25871), .B(n25867), .Z(n25918) );
  XNOR U27338 ( .A(n25866), .B(n25862), .Z(n25919) );
  XNOR U27339 ( .A(n25861), .B(n25857), .Z(n25920) );
  XNOR U27340 ( .A(n25856), .B(n25852), .Z(n25921) );
  XNOR U27341 ( .A(n25851), .B(n25847), .Z(n25922) );
  XNOR U27342 ( .A(n25846), .B(n25842), .Z(n25923) );
  XNOR U27343 ( .A(n25841), .B(n25837), .Z(n25924) );
  XNOR U27344 ( .A(n25836), .B(n25832), .Z(n25925) );
  XNOR U27345 ( .A(n25831), .B(n25827), .Z(n25926) );
  XNOR U27346 ( .A(n25826), .B(n25822), .Z(n25927) );
  XNOR U27347 ( .A(n25821), .B(n25817), .Z(n25928) );
  XNOR U27348 ( .A(n25816), .B(n25812), .Z(n25929) );
  XNOR U27349 ( .A(n25811), .B(n25807), .Z(n25930) );
  XNOR U27350 ( .A(n25806), .B(n25802), .Z(n25931) );
  XNOR U27351 ( .A(n25801), .B(n25797), .Z(n25932) );
  XNOR U27352 ( .A(n25796), .B(n25792), .Z(n25933) );
  XNOR U27353 ( .A(n25791), .B(n25787), .Z(n25934) );
  XNOR U27354 ( .A(n25786), .B(n25782), .Z(n25935) );
  XNOR U27355 ( .A(n25781), .B(n25777), .Z(n25936) );
  XNOR U27356 ( .A(n25776), .B(n25772), .Z(n25937) );
  XNOR U27357 ( .A(n25771), .B(n25767), .Z(n25938) );
  XNOR U27358 ( .A(n25766), .B(n25762), .Z(n25939) );
  XNOR U27359 ( .A(n25761), .B(n25757), .Z(n25940) );
  XNOR U27360 ( .A(n25756), .B(n25752), .Z(n25941) );
  XNOR U27361 ( .A(n25751), .B(n25747), .Z(n25942) );
  XNOR U27362 ( .A(n25746), .B(n25742), .Z(n25943) );
  XNOR U27363 ( .A(n25741), .B(n25737), .Z(n25944) );
  XNOR U27364 ( .A(n25736), .B(n25732), .Z(n25945) );
  XNOR U27365 ( .A(n25731), .B(n25727), .Z(n25946) );
  XNOR U27366 ( .A(n25726), .B(n25722), .Z(n25947) );
  XNOR U27367 ( .A(n25721), .B(n25717), .Z(n25948) );
  XNOR U27368 ( .A(n25716), .B(n25712), .Z(n25949) );
  XNOR U27369 ( .A(n25711), .B(n25707), .Z(n25950) );
  XNOR U27370 ( .A(n25706), .B(n25702), .Z(n25951) );
  XNOR U27371 ( .A(n25701), .B(n25697), .Z(n25952) );
  XNOR U27372 ( .A(n25696), .B(n25692), .Z(n25953) );
  XNOR U27373 ( .A(n25691), .B(n25687), .Z(n25954) );
  XNOR U27374 ( .A(n25686), .B(n25682), .Z(n25955) );
  XNOR U27375 ( .A(n25681), .B(n25677), .Z(n25956) );
  XNOR U27376 ( .A(n25676), .B(n25672), .Z(n25957) );
  XNOR U27377 ( .A(n25671), .B(n25667), .Z(n25958) );
  XNOR U27378 ( .A(n25666), .B(n25662), .Z(n25959) );
  XNOR U27379 ( .A(n25661), .B(n25657), .Z(n25960) );
  XNOR U27380 ( .A(n25656), .B(n25652), .Z(n25961) );
  XNOR U27381 ( .A(n25651), .B(n25647), .Z(n25962) );
  XNOR U27382 ( .A(n25646), .B(n25642), .Z(n25963) );
  XNOR U27383 ( .A(n25641), .B(n25637), .Z(n25964) );
  XNOR U27384 ( .A(n25636), .B(n25632), .Z(n25965) );
  XNOR U27385 ( .A(n25631), .B(n25627), .Z(n25966) );
  XOR U27386 ( .A(n25967), .B(n25626), .Z(n25627) );
  AND U27387 ( .A(a[0]), .B(b[57]), .Z(n25967) );
  XOR U27388 ( .A(n25968), .B(n25626), .Z(n25628) );
  XNOR U27389 ( .A(n25969), .B(n25970), .Z(n25626) );
  AND U27390 ( .A(n25971), .B(n25972), .Z(n25969) );
  AND U27391 ( .A(a[1]), .B(b[56]), .Z(n25968) );
  XOR U27392 ( .A(n25973), .B(n25631), .Z(n25633) );
  XOR U27393 ( .A(n25974), .B(n25975), .Z(n25631) );
  AND U27394 ( .A(n25976), .B(n25977), .Z(n25974) );
  AND U27395 ( .A(a[2]), .B(b[55]), .Z(n25973) );
  XOR U27396 ( .A(n25978), .B(n25636), .Z(n25638) );
  XOR U27397 ( .A(n25979), .B(n25980), .Z(n25636) );
  AND U27398 ( .A(n25981), .B(n25982), .Z(n25979) );
  AND U27399 ( .A(a[3]), .B(b[54]), .Z(n25978) );
  XOR U27400 ( .A(n25983), .B(n25641), .Z(n25643) );
  XOR U27401 ( .A(n25984), .B(n25985), .Z(n25641) );
  AND U27402 ( .A(n25986), .B(n25987), .Z(n25984) );
  AND U27403 ( .A(a[4]), .B(b[53]), .Z(n25983) );
  XOR U27404 ( .A(n25988), .B(n25646), .Z(n25648) );
  XOR U27405 ( .A(n25989), .B(n25990), .Z(n25646) );
  AND U27406 ( .A(n25991), .B(n25992), .Z(n25989) );
  AND U27407 ( .A(a[5]), .B(b[52]), .Z(n25988) );
  XOR U27408 ( .A(n25993), .B(n25651), .Z(n25653) );
  XOR U27409 ( .A(n25994), .B(n25995), .Z(n25651) );
  AND U27410 ( .A(n25996), .B(n25997), .Z(n25994) );
  AND U27411 ( .A(a[6]), .B(b[51]), .Z(n25993) );
  XOR U27412 ( .A(n25998), .B(n25656), .Z(n25658) );
  XOR U27413 ( .A(n25999), .B(n26000), .Z(n25656) );
  AND U27414 ( .A(n26001), .B(n26002), .Z(n25999) );
  AND U27415 ( .A(a[7]), .B(b[50]), .Z(n25998) );
  XOR U27416 ( .A(n26003), .B(n25661), .Z(n25663) );
  XOR U27417 ( .A(n26004), .B(n26005), .Z(n25661) );
  AND U27418 ( .A(n26006), .B(n26007), .Z(n26004) );
  AND U27419 ( .A(a[8]), .B(b[49]), .Z(n26003) );
  XOR U27420 ( .A(n26008), .B(n25666), .Z(n25668) );
  XOR U27421 ( .A(n26009), .B(n26010), .Z(n25666) );
  AND U27422 ( .A(n26011), .B(n26012), .Z(n26009) );
  AND U27423 ( .A(a[9]), .B(b[48]), .Z(n26008) );
  XOR U27424 ( .A(n26013), .B(n25671), .Z(n25673) );
  XOR U27425 ( .A(n26014), .B(n26015), .Z(n25671) );
  AND U27426 ( .A(n26016), .B(n26017), .Z(n26014) );
  AND U27427 ( .A(a[10]), .B(b[47]), .Z(n26013) );
  XOR U27428 ( .A(n26018), .B(n25676), .Z(n25678) );
  XOR U27429 ( .A(n26019), .B(n26020), .Z(n25676) );
  AND U27430 ( .A(n26021), .B(n26022), .Z(n26019) );
  AND U27431 ( .A(a[11]), .B(b[46]), .Z(n26018) );
  XOR U27432 ( .A(n26023), .B(n25681), .Z(n25683) );
  XOR U27433 ( .A(n26024), .B(n26025), .Z(n25681) );
  AND U27434 ( .A(n26026), .B(n26027), .Z(n26024) );
  AND U27435 ( .A(a[12]), .B(b[45]), .Z(n26023) );
  XOR U27436 ( .A(n26028), .B(n25686), .Z(n25688) );
  XOR U27437 ( .A(n26029), .B(n26030), .Z(n25686) );
  AND U27438 ( .A(n26031), .B(n26032), .Z(n26029) );
  AND U27439 ( .A(a[13]), .B(b[44]), .Z(n26028) );
  XOR U27440 ( .A(n26033), .B(n25691), .Z(n25693) );
  XOR U27441 ( .A(n26034), .B(n26035), .Z(n25691) );
  AND U27442 ( .A(n26036), .B(n26037), .Z(n26034) );
  AND U27443 ( .A(a[14]), .B(b[43]), .Z(n26033) );
  XOR U27444 ( .A(n26038), .B(n25696), .Z(n25698) );
  XOR U27445 ( .A(n26039), .B(n26040), .Z(n25696) );
  AND U27446 ( .A(n26041), .B(n26042), .Z(n26039) );
  AND U27447 ( .A(a[15]), .B(b[42]), .Z(n26038) );
  XOR U27448 ( .A(n26043), .B(n25701), .Z(n25703) );
  XOR U27449 ( .A(n26044), .B(n26045), .Z(n25701) );
  AND U27450 ( .A(n26046), .B(n26047), .Z(n26044) );
  AND U27451 ( .A(a[16]), .B(b[41]), .Z(n26043) );
  XOR U27452 ( .A(n26048), .B(n25706), .Z(n25708) );
  XOR U27453 ( .A(n26049), .B(n26050), .Z(n25706) );
  AND U27454 ( .A(n26051), .B(n26052), .Z(n26049) );
  AND U27455 ( .A(a[17]), .B(b[40]), .Z(n26048) );
  XOR U27456 ( .A(n26053), .B(n25711), .Z(n25713) );
  XOR U27457 ( .A(n26054), .B(n26055), .Z(n25711) );
  AND U27458 ( .A(n26056), .B(n26057), .Z(n26054) );
  AND U27459 ( .A(a[18]), .B(b[39]), .Z(n26053) );
  XOR U27460 ( .A(n26058), .B(n25716), .Z(n25718) );
  XOR U27461 ( .A(n26059), .B(n26060), .Z(n25716) );
  AND U27462 ( .A(n26061), .B(n26062), .Z(n26059) );
  AND U27463 ( .A(a[19]), .B(b[38]), .Z(n26058) );
  XOR U27464 ( .A(n26063), .B(n25721), .Z(n25723) );
  XOR U27465 ( .A(n26064), .B(n26065), .Z(n25721) );
  AND U27466 ( .A(n26066), .B(n26067), .Z(n26064) );
  AND U27467 ( .A(a[20]), .B(b[37]), .Z(n26063) );
  XOR U27468 ( .A(n26068), .B(n25726), .Z(n25728) );
  XOR U27469 ( .A(n26069), .B(n26070), .Z(n25726) );
  AND U27470 ( .A(n26071), .B(n26072), .Z(n26069) );
  AND U27471 ( .A(a[21]), .B(b[36]), .Z(n26068) );
  XOR U27472 ( .A(n26073), .B(n25731), .Z(n25733) );
  XOR U27473 ( .A(n26074), .B(n26075), .Z(n25731) );
  AND U27474 ( .A(n26076), .B(n26077), .Z(n26074) );
  AND U27475 ( .A(a[22]), .B(b[35]), .Z(n26073) );
  XOR U27476 ( .A(n26078), .B(n25736), .Z(n25738) );
  XOR U27477 ( .A(n26079), .B(n26080), .Z(n25736) );
  AND U27478 ( .A(n26081), .B(n26082), .Z(n26079) );
  AND U27479 ( .A(a[23]), .B(b[34]), .Z(n26078) );
  XOR U27480 ( .A(n26083), .B(n25741), .Z(n25743) );
  XOR U27481 ( .A(n26084), .B(n26085), .Z(n25741) );
  AND U27482 ( .A(n26086), .B(n26087), .Z(n26084) );
  AND U27483 ( .A(a[24]), .B(b[33]), .Z(n26083) );
  XOR U27484 ( .A(n26088), .B(n25746), .Z(n25748) );
  XOR U27485 ( .A(n26089), .B(n26090), .Z(n25746) );
  AND U27486 ( .A(n26091), .B(n26092), .Z(n26089) );
  AND U27487 ( .A(a[25]), .B(b[32]), .Z(n26088) );
  XOR U27488 ( .A(n26093), .B(n25751), .Z(n25753) );
  XOR U27489 ( .A(n26094), .B(n26095), .Z(n25751) );
  AND U27490 ( .A(n26096), .B(n26097), .Z(n26094) );
  AND U27491 ( .A(a[26]), .B(b[31]), .Z(n26093) );
  XOR U27492 ( .A(n26098), .B(n25756), .Z(n25758) );
  XOR U27493 ( .A(n26099), .B(n26100), .Z(n25756) );
  AND U27494 ( .A(n26101), .B(n26102), .Z(n26099) );
  AND U27495 ( .A(a[27]), .B(b[30]), .Z(n26098) );
  XOR U27496 ( .A(n26103), .B(n25761), .Z(n25763) );
  XOR U27497 ( .A(n26104), .B(n26105), .Z(n25761) );
  AND U27498 ( .A(n26106), .B(n26107), .Z(n26104) );
  AND U27499 ( .A(a[28]), .B(b[29]), .Z(n26103) );
  XOR U27500 ( .A(n26108), .B(n25766), .Z(n25768) );
  XOR U27501 ( .A(n26109), .B(n26110), .Z(n25766) );
  AND U27502 ( .A(n26111), .B(n26112), .Z(n26109) );
  AND U27503 ( .A(b[28]), .B(a[29]), .Z(n26108) );
  XOR U27504 ( .A(n26113), .B(n25771), .Z(n25773) );
  XOR U27505 ( .A(n26114), .B(n26115), .Z(n25771) );
  AND U27506 ( .A(n26116), .B(n26117), .Z(n26114) );
  AND U27507 ( .A(b[27]), .B(a[30]), .Z(n26113) );
  XOR U27508 ( .A(n26118), .B(n25776), .Z(n25778) );
  XOR U27509 ( .A(n26119), .B(n26120), .Z(n25776) );
  AND U27510 ( .A(n26121), .B(n26122), .Z(n26119) );
  AND U27511 ( .A(b[26]), .B(a[31]), .Z(n26118) );
  XOR U27512 ( .A(n26123), .B(n25781), .Z(n25783) );
  XOR U27513 ( .A(n26124), .B(n26125), .Z(n25781) );
  AND U27514 ( .A(n26126), .B(n26127), .Z(n26124) );
  AND U27515 ( .A(b[25]), .B(a[32]), .Z(n26123) );
  XOR U27516 ( .A(n26128), .B(n25786), .Z(n25788) );
  XOR U27517 ( .A(n26129), .B(n26130), .Z(n25786) );
  AND U27518 ( .A(n26131), .B(n26132), .Z(n26129) );
  AND U27519 ( .A(b[24]), .B(a[33]), .Z(n26128) );
  XOR U27520 ( .A(n26133), .B(n25791), .Z(n25793) );
  XOR U27521 ( .A(n26134), .B(n26135), .Z(n25791) );
  AND U27522 ( .A(n26136), .B(n26137), .Z(n26134) );
  AND U27523 ( .A(b[23]), .B(a[34]), .Z(n26133) );
  XOR U27524 ( .A(n26138), .B(n25796), .Z(n25798) );
  XOR U27525 ( .A(n26139), .B(n26140), .Z(n25796) );
  AND U27526 ( .A(n26141), .B(n26142), .Z(n26139) );
  AND U27527 ( .A(b[22]), .B(a[35]), .Z(n26138) );
  XOR U27528 ( .A(n26143), .B(n25801), .Z(n25803) );
  XOR U27529 ( .A(n26144), .B(n26145), .Z(n25801) );
  AND U27530 ( .A(n26146), .B(n26147), .Z(n26144) );
  AND U27531 ( .A(b[21]), .B(a[36]), .Z(n26143) );
  XOR U27532 ( .A(n26148), .B(n25806), .Z(n25808) );
  XOR U27533 ( .A(n26149), .B(n26150), .Z(n25806) );
  AND U27534 ( .A(n26151), .B(n26152), .Z(n26149) );
  AND U27535 ( .A(b[20]), .B(a[37]), .Z(n26148) );
  XOR U27536 ( .A(n26153), .B(n25811), .Z(n25813) );
  XOR U27537 ( .A(n26154), .B(n26155), .Z(n25811) );
  AND U27538 ( .A(n26156), .B(n26157), .Z(n26154) );
  AND U27539 ( .A(b[19]), .B(a[38]), .Z(n26153) );
  XOR U27540 ( .A(n26158), .B(n25816), .Z(n25818) );
  XOR U27541 ( .A(n26159), .B(n26160), .Z(n25816) );
  AND U27542 ( .A(n26161), .B(n26162), .Z(n26159) );
  AND U27543 ( .A(b[18]), .B(a[39]), .Z(n26158) );
  XOR U27544 ( .A(n26163), .B(n25821), .Z(n25823) );
  XOR U27545 ( .A(n26164), .B(n26165), .Z(n25821) );
  AND U27546 ( .A(n26166), .B(n26167), .Z(n26164) );
  AND U27547 ( .A(b[17]), .B(a[40]), .Z(n26163) );
  XOR U27548 ( .A(n26168), .B(n25826), .Z(n25828) );
  XOR U27549 ( .A(n26169), .B(n26170), .Z(n25826) );
  AND U27550 ( .A(n26171), .B(n26172), .Z(n26169) );
  AND U27551 ( .A(b[16]), .B(a[41]), .Z(n26168) );
  XOR U27552 ( .A(n26173), .B(n25831), .Z(n25833) );
  XOR U27553 ( .A(n26174), .B(n26175), .Z(n25831) );
  AND U27554 ( .A(n26176), .B(n26177), .Z(n26174) );
  AND U27555 ( .A(b[15]), .B(a[42]), .Z(n26173) );
  XOR U27556 ( .A(n26178), .B(n25836), .Z(n25838) );
  XOR U27557 ( .A(n26179), .B(n26180), .Z(n25836) );
  AND U27558 ( .A(n26181), .B(n26182), .Z(n26179) );
  AND U27559 ( .A(b[14]), .B(a[43]), .Z(n26178) );
  XOR U27560 ( .A(n26183), .B(n25841), .Z(n25843) );
  XOR U27561 ( .A(n26184), .B(n26185), .Z(n25841) );
  AND U27562 ( .A(n26186), .B(n26187), .Z(n26184) );
  AND U27563 ( .A(b[13]), .B(a[44]), .Z(n26183) );
  XOR U27564 ( .A(n26188), .B(n25846), .Z(n25848) );
  XOR U27565 ( .A(n26189), .B(n26190), .Z(n25846) );
  AND U27566 ( .A(n26191), .B(n26192), .Z(n26189) );
  AND U27567 ( .A(b[12]), .B(a[45]), .Z(n26188) );
  XOR U27568 ( .A(n26193), .B(n25851), .Z(n25853) );
  XOR U27569 ( .A(n26194), .B(n26195), .Z(n25851) );
  AND U27570 ( .A(n26196), .B(n26197), .Z(n26194) );
  AND U27571 ( .A(b[11]), .B(a[46]), .Z(n26193) );
  XOR U27572 ( .A(n26198), .B(n25856), .Z(n25858) );
  XOR U27573 ( .A(n26199), .B(n26200), .Z(n25856) );
  AND U27574 ( .A(n26201), .B(n26202), .Z(n26199) );
  AND U27575 ( .A(b[10]), .B(a[47]), .Z(n26198) );
  XOR U27576 ( .A(n26203), .B(n25861), .Z(n25863) );
  XOR U27577 ( .A(n26204), .B(n26205), .Z(n25861) );
  AND U27578 ( .A(n26206), .B(n26207), .Z(n26204) );
  AND U27579 ( .A(b[9]), .B(a[48]), .Z(n26203) );
  XOR U27580 ( .A(n26208), .B(n25866), .Z(n25868) );
  XOR U27581 ( .A(n26209), .B(n26210), .Z(n25866) );
  AND U27582 ( .A(n26211), .B(n26212), .Z(n26209) );
  AND U27583 ( .A(b[8]), .B(a[49]), .Z(n26208) );
  XOR U27584 ( .A(n26213), .B(n25871), .Z(n25873) );
  XOR U27585 ( .A(n26214), .B(n26215), .Z(n25871) );
  AND U27586 ( .A(n26216), .B(n26217), .Z(n26214) );
  AND U27587 ( .A(b[7]), .B(a[50]), .Z(n26213) );
  XOR U27588 ( .A(n26218), .B(n25876), .Z(n25878) );
  XOR U27589 ( .A(n26219), .B(n26220), .Z(n25876) );
  AND U27590 ( .A(n26221), .B(n26222), .Z(n26219) );
  AND U27591 ( .A(b[6]), .B(a[51]), .Z(n26218) );
  XOR U27592 ( .A(n26223), .B(n25881), .Z(n25883) );
  XOR U27593 ( .A(n26224), .B(n26225), .Z(n25881) );
  AND U27594 ( .A(n26226), .B(n26227), .Z(n26224) );
  AND U27595 ( .A(b[5]), .B(a[52]), .Z(n26223) );
  XOR U27596 ( .A(n26228), .B(n25886), .Z(n25888) );
  XOR U27597 ( .A(n26229), .B(n26230), .Z(n25886) );
  AND U27598 ( .A(n26231), .B(n26232), .Z(n26229) );
  AND U27599 ( .A(b[4]), .B(a[53]), .Z(n26228) );
  XNOR U27600 ( .A(n26233), .B(n26234), .Z(n25900) );
  NANDN U27601 ( .A(n26235), .B(n26236), .Z(n26234) );
  XOR U27602 ( .A(n26237), .B(n25891), .Z(n25893) );
  XNOR U27603 ( .A(n26238), .B(n26239), .Z(n25891) );
  AND U27604 ( .A(n26240), .B(n26241), .Z(n26238) );
  AND U27605 ( .A(b[3]), .B(a[54]), .Z(n26237) );
  XOR U27606 ( .A(n25907), .B(n25906), .Z(c[120]) );
  XOR U27607 ( .A(sreg[184]), .B(n25905), .Z(n25906) );
  XOR U27608 ( .A(n25912), .B(n26242), .Z(n25907) );
  XNOR U27609 ( .A(n25911), .B(n25905), .Z(n26242) );
  XOR U27610 ( .A(n26243), .B(n26244), .Z(n25905) );
  NOR U27611 ( .A(n26245), .B(n26246), .Z(n26243) );
  NAND U27612 ( .A(a[56]), .B(b[0]), .Z(n25911) );
  XNOR U27613 ( .A(n26235), .B(n26236), .Z(n25912) );
  XOR U27614 ( .A(n26233), .B(n26247), .Z(n26236) );
  NAND U27615 ( .A(b[1]), .B(a[55]), .Z(n26247) );
  XOR U27616 ( .A(n26241), .B(n26248), .Z(n26235) );
  XOR U27617 ( .A(n26233), .B(n26240), .Z(n26248) );
  XNOR U27618 ( .A(n26249), .B(n26239), .Z(n26240) );
  AND U27619 ( .A(b[2]), .B(a[54]), .Z(n26249) );
  NANDN U27620 ( .A(n26250), .B(n26251), .Z(n26233) );
  XOR U27621 ( .A(n26239), .B(n26231), .Z(n26252) );
  XNOR U27622 ( .A(n26230), .B(n26226), .Z(n26253) );
  XNOR U27623 ( .A(n26225), .B(n26221), .Z(n26254) );
  XNOR U27624 ( .A(n26220), .B(n26216), .Z(n26255) );
  XNOR U27625 ( .A(n26215), .B(n26211), .Z(n26256) );
  XNOR U27626 ( .A(n26210), .B(n26206), .Z(n26257) );
  XNOR U27627 ( .A(n26205), .B(n26201), .Z(n26258) );
  XNOR U27628 ( .A(n26200), .B(n26196), .Z(n26259) );
  XNOR U27629 ( .A(n26195), .B(n26191), .Z(n26260) );
  XNOR U27630 ( .A(n26190), .B(n26186), .Z(n26261) );
  XNOR U27631 ( .A(n26185), .B(n26181), .Z(n26262) );
  XNOR U27632 ( .A(n26180), .B(n26176), .Z(n26263) );
  XNOR U27633 ( .A(n26175), .B(n26171), .Z(n26264) );
  XNOR U27634 ( .A(n26170), .B(n26166), .Z(n26265) );
  XNOR U27635 ( .A(n26165), .B(n26161), .Z(n26266) );
  XNOR U27636 ( .A(n26160), .B(n26156), .Z(n26267) );
  XNOR U27637 ( .A(n26155), .B(n26151), .Z(n26268) );
  XNOR U27638 ( .A(n26150), .B(n26146), .Z(n26269) );
  XNOR U27639 ( .A(n26145), .B(n26141), .Z(n26270) );
  XNOR U27640 ( .A(n26140), .B(n26136), .Z(n26271) );
  XNOR U27641 ( .A(n26135), .B(n26131), .Z(n26272) );
  XNOR U27642 ( .A(n26130), .B(n26126), .Z(n26273) );
  XNOR U27643 ( .A(n26125), .B(n26121), .Z(n26274) );
  XNOR U27644 ( .A(n26120), .B(n26116), .Z(n26275) );
  XNOR U27645 ( .A(n26115), .B(n26111), .Z(n26276) );
  XNOR U27646 ( .A(n26110), .B(n26106), .Z(n26277) );
  XNOR U27647 ( .A(n26105), .B(n26101), .Z(n26278) );
  XNOR U27648 ( .A(n26100), .B(n26096), .Z(n26279) );
  XNOR U27649 ( .A(n26095), .B(n26091), .Z(n26280) );
  XNOR U27650 ( .A(n26090), .B(n26086), .Z(n26281) );
  XNOR U27651 ( .A(n26085), .B(n26081), .Z(n26282) );
  XNOR U27652 ( .A(n26080), .B(n26076), .Z(n26283) );
  XNOR U27653 ( .A(n26075), .B(n26071), .Z(n26284) );
  XNOR U27654 ( .A(n26070), .B(n26066), .Z(n26285) );
  XNOR U27655 ( .A(n26065), .B(n26061), .Z(n26286) );
  XNOR U27656 ( .A(n26060), .B(n26056), .Z(n26287) );
  XNOR U27657 ( .A(n26055), .B(n26051), .Z(n26288) );
  XNOR U27658 ( .A(n26050), .B(n26046), .Z(n26289) );
  XNOR U27659 ( .A(n26045), .B(n26041), .Z(n26290) );
  XNOR U27660 ( .A(n26040), .B(n26036), .Z(n26291) );
  XNOR U27661 ( .A(n26035), .B(n26031), .Z(n26292) );
  XNOR U27662 ( .A(n26030), .B(n26026), .Z(n26293) );
  XNOR U27663 ( .A(n26025), .B(n26021), .Z(n26294) );
  XNOR U27664 ( .A(n26020), .B(n26016), .Z(n26295) );
  XNOR U27665 ( .A(n26015), .B(n26011), .Z(n26296) );
  XNOR U27666 ( .A(n26010), .B(n26006), .Z(n26297) );
  XNOR U27667 ( .A(n26005), .B(n26001), .Z(n26298) );
  XNOR U27668 ( .A(n26000), .B(n25996), .Z(n26299) );
  XNOR U27669 ( .A(n25995), .B(n25991), .Z(n26300) );
  XNOR U27670 ( .A(n25990), .B(n25986), .Z(n26301) );
  XNOR U27671 ( .A(n25985), .B(n25981), .Z(n26302) );
  XNOR U27672 ( .A(n25980), .B(n25976), .Z(n26303) );
  XNOR U27673 ( .A(n25975), .B(n25971), .Z(n26304) );
  XNOR U27674 ( .A(n26305), .B(n25970), .Z(n25971) );
  AND U27675 ( .A(a[0]), .B(b[56]), .Z(n26305) );
  XNOR U27676 ( .A(n26306), .B(n25970), .Z(n25972) );
  XNOR U27677 ( .A(n26307), .B(n26308), .Z(n25970) );
  AND U27678 ( .A(n26309), .B(n26310), .Z(n26307) );
  AND U27679 ( .A(a[1]), .B(b[55]), .Z(n26306) );
  XOR U27680 ( .A(n26311), .B(n25975), .Z(n25977) );
  XOR U27681 ( .A(n26312), .B(n26313), .Z(n25975) );
  AND U27682 ( .A(n26314), .B(n26315), .Z(n26312) );
  AND U27683 ( .A(a[2]), .B(b[54]), .Z(n26311) );
  XOR U27684 ( .A(n26316), .B(n25980), .Z(n25982) );
  XOR U27685 ( .A(n26317), .B(n26318), .Z(n25980) );
  AND U27686 ( .A(n26319), .B(n26320), .Z(n26317) );
  AND U27687 ( .A(a[3]), .B(b[53]), .Z(n26316) );
  XOR U27688 ( .A(n26321), .B(n25985), .Z(n25987) );
  XOR U27689 ( .A(n26322), .B(n26323), .Z(n25985) );
  AND U27690 ( .A(n26324), .B(n26325), .Z(n26322) );
  AND U27691 ( .A(a[4]), .B(b[52]), .Z(n26321) );
  XOR U27692 ( .A(n26326), .B(n25990), .Z(n25992) );
  XOR U27693 ( .A(n26327), .B(n26328), .Z(n25990) );
  AND U27694 ( .A(n26329), .B(n26330), .Z(n26327) );
  AND U27695 ( .A(a[5]), .B(b[51]), .Z(n26326) );
  XOR U27696 ( .A(n26331), .B(n25995), .Z(n25997) );
  XOR U27697 ( .A(n26332), .B(n26333), .Z(n25995) );
  AND U27698 ( .A(n26334), .B(n26335), .Z(n26332) );
  AND U27699 ( .A(a[6]), .B(b[50]), .Z(n26331) );
  XOR U27700 ( .A(n26336), .B(n26000), .Z(n26002) );
  XOR U27701 ( .A(n26337), .B(n26338), .Z(n26000) );
  AND U27702 ( .A(n26339), .B(n26340), .Z(n26337) );
  AND U27703 ( .A(a[7]), .B(b[49]), .Z(n26336) );
  XOR U27704 ( .A(n26341), .B(n26005), .Z(n26007) );
  XOR U27705 ( .A(n26342), .B(n26343), .Z(n26005) );
  AND U27706 ( .A(n26344), .B(n26345), .Z(n26342) );
  AND U27707 ( .A(a[8]), .B(b[48]), .Z(n26341) );
  XOR U27708 ( .A(n26346), .B(n26010), .Z(n26012) );
  XOR U27709 ( .A(n26347), .B(n26348), .Z(n26010) );
  AND U27710 ( .A(n26349), .B(n26350), .Z(n26347) );
  AND U27711 ( .A(a[9]), .B(b[47]), .Z(n26346) );
  XOR U27712 ( .A(n26351), .B(n26015), .Z(n26017) );
  XOR U27713 ( .A(n26352), .B(n26353), .Z(n26015) );
  AND U27714 ( .A(n26354), .B(n26355), .Z(n26352) );
  AND U27715 ( .A(a[10]), .B(b[46]), .Z(n26351) );
  XOR U27716 ( .A(n26356), .B(n26020), .Z(n26022) );
  XOR U27717 ( .A(n26357), .B(n26358), .Z(n26020) );
  AND U27718 ( .A(n26359), .B(n26360), .Z(n26357) );
  AND U27719 ( .A(a[11]), .B(b[45]), .Z(n26356) );
  XOR U27720 ( .A(n26361), .B(n26025), .Z(n26027) );
  XOR U27721 ( .A(n26362), .B(n26363), .Z(n26025) );
  AND U27722 ( .A(n26364), .B(n26365), .Z(n26362) );
  AND U27723 ( .A(a[12]), .B(b[44]), .Z(n26361) );
  XOR U27724 ( .A(n26366), .B(n26030), .Z(n26032) );
  XOR U27725 ( .A(n26367), .B(n26368), .Z(n26030) );
  AND U27726 ( .A(n26369), .B(n26370), .Z(n26367) );
  AND U27727 ( .A(a[13]), .B(b[43]), .Z(n26366) );
  XOR U27728 ( .A(n26371), .B(n26035), .Z(n26037) );
  XOR U27729 ( .A(n26372), .B(n26373), .Z(n26035) );
  AND U27730 ( .A(n26374), .B(n26375), .Z(n26372) );
  AND U27731 ( .A(a[14]), .B(b[42]), .Z(n26371) );
  XOR U27732 ( .A(n26376), .B(n26040), .Z(n26042) );
  XOR U27733 ( .A(n26377), .B(n26378), .Z(n26040) );
  AND U27734 ( .A(n26379), .B(n26380), .Z(n26377) );
  AND U27735 ( .A(a[15]), .B(b[41]), .Z(n26376) );
  XOR U27736 ( .A(n26381), .B(n26045), .Z(n26047) );
  XOR U27737 ( .A(n26382), .B(n26383), .Z(n26045) );
  AND U27738 ( .A(n26384), .B(n26385), .Z(n26382) );
  AND U27739 ( .A(a[16]), .B(b[40]), .Z(n26381) );
  XOR U27740 ( .A(n26386), .B(n26050), .Z(n26052) );
  XOR U27741 ( .A(n26387), .B(n26388), .Z(n26050) );
  AND U27742 ( .A(n26389), .B(n26390), .Z(n26387) );
  AND U27743 ( .A(a[17]), .B(b[39]), .Z(n26386) );
  XOR U27744 ( .A(n26391), .B(n26055), .Z(n26057) );
  XOR U27745 ( .A(n26392), .B(n26393), .Z(n26055) );
  AND U27746 ( .A(n26394), .B(n26395), .Z(n26392) );
  AND U27747 ( .A(a[18]), .B(b[38]), .Z(n26391) );
  XOR U27748 ( .A(n26396), .B(n26060), .Z(n26062) );
  XOR U27749 ( .A(n26397), .B(n26398), .Z(n26060) );
  AND U27750 ( .A(n26399), .B(n26400), .Z(n26397) );
  AND U27751 ( .A(a[19]), .B(b[37]), .Z(n26396) );
  XOR U27752 ( .A(n26401), .B(n26065), .Z(n26067) );
  XOR U27753 ( .A(n26402), .B(n26403), .Z(n26065) );
  AND U27754 ( .A(n26404), .B(n26405), .Z(n26402) );
  AND U27755 ( .A(a[20]), .B(b[36]), .Z(n26401) );
  XOR U27756 ( .A(n26406), .B(n26070), .Z(n26072) );
  XOR U27757 ( .A(n26407), .B(n26408), .Z(n26070) );
  AND U27758 ( .A(n26409), .B(n26410), .Z(n26407) );
  AND U27759 ( .A(a[21]), .B(b[35]), .Z(n26406) );
  XOR U27760 ( .A(n26411), .B(n26075), .Z(n26077) );
  XOR U27761 ( .A(n26412), .B(n26413), .Z(n26075) );
  AND U27762 ( .A(n26414), .B(n26415), .Z(n26412) );
  AND U27763 ( .A(a[22]), .B(b[34]), .Z(n26411) );
  XOR U27764 ( .A(n26416), .B(n26080), .Z(n26082) );
  XOR U27765 ( .A(n26417), .B(n26418), .Z(n26080) );
  AND U27766 ( .A(n26419), .B(n26420), .Z(n26417) );
  AND U27767 ( .A(a[23]), .B(b[33]), .Z(n26416) );
  XOR U27768 ( .A(n26421), .B(n26085), .Z(n26087) );
  XOR U27769 ( .A(n26422), .B(n26423), .Z(n26085) );
  AND U27770 ( .A(n26424), .B(n26425), .Z(n26422) );
  AND U27771 ( .A(a[24]), .B(b[32]), .Z(n26421) );
  XOR U27772 ( .A(n26426), .B(n26090), .Z(n26092) );
  XOR U27773 ( .A(n26427), .B(n26428), .Z(n26090) );
  AND U27774 ( .A(n26429), .B(n26430), .Z(n26427) );
  AND U27775 ( .A(a[25]), .B(b[31]), .Z(n26426) );
  XOR U27776 ( .A(n26431), .B(n26095), .Z(n26097) );
  XOR U27777 ( .A(n26432), .B(n26433), .Z(n26095) );
  AND U27778 ( .A(n26434), .B(n26435), .Z(n26432) );
  AND U27779 ( .A(a[26]), .B(b[30]), .Z(n26431) );
  XOR U27780 ( .A(n26436), .B(n26100), .Z(n26102) );
  XOR U27781 ( .A(n26437), .B(n26438), .Z(n26100) );
  AND U27782 ( .A(n26439), .B(n26440), .Z(n26437) );
  AND U27783 ( .A(a[27]), .B(b[29]), .Z(n26436) );
  XOR U27784 ( .A(n26441), .B(n26105), .Z(n26107) );
  XOR U27785 ( .A(n26442), .B(n26443), .Z(n26105) );
  AND U27786 ( .A(n26444), .B(n26445), .Z(n26442) );
  AND U27787 ( .A(a[28]), .B(b[28]), .Z(n26441) );
  XOR U27788 ( .A(n26446), .B(n26110), .Z(n26112) );
  XOR U27789 ( .A(n26447), .B(n26448), .Z(n26110) );
  AND U27790 ( .A(n26449), .B(n26450), .Z(n26447) );
  AND U27791 ( .A(b[27]), .B(a[29]), .Z(n26446) );
  XOR U27792 ( .A(n26451), .B(n26115), .Z(n26117) );
  XOR U27793 ( .A(n26452), .B(n26453), .Z(n26115) );
  AND U27794 ( .A(n26454), .B(n26455), .Z(n26452) );
  AND U27795 ( .A(b[26]), .B(a[30]), .Z(n26451) );
  XOR U27796 ( .A(n26456), .B(n26120), .Z(n26122) );
  XOR U27797 ( .A(n26457), .B(n26458), .Z(n26120) );
  AND U27798 ( .A(n26459), .B(n26460), .Z(n26457) );
  AND U27799 ( .A(b[25]), .B(a[31]), .Z(n26456) );
  XOR U27800 ( .A(n26461), .B(n26125), .Z(n26127) );
  XOR U27801 ( .A(n26462), .B(n26463), .Z(n26125) );
  AND U27802 ( .A(n26464), .B(n26465), .Z(n26462) );
  AND U27803 ( .A(b[24]), .B(a[32]), .Z(n26461) );
  XOR U27804 ( .A(n26466), .B(n26130), .Z(n26132) );
  XOR U27805 ( .A(n26467), .B(n26468), .Z(n26130) );
  AND U27806 ( .A(n26469), .B(n26470), .Z(n26467) );
  AND U27807 ( .A(b[23]), .B(a[33]), .Z(n26466) );
  XOR U27808 ( .A(n26471), .B(n26135), .Z(n26137) );
  XOR U27809 ( .A(n26472), .B(n26473), .Z(n26135) );
  AND U27810 ( .A(n26474), .B(n26475), .Z(n26472) );
  AND U27811 ( .A(b[22]), .B(a[34]), .Z(n26471) );
  XOR U27812 ( .A(n26476), .B(n26140), .Z(n26142) );
  XOR U27813 ( .A(n26477), .B(n26478), .Z(n26140) );
  AND U27814 ( .A(n26479), .B(n26480), .Z(n26477) );
  AND U27815 ( .A(b[21]), .B(a[35]), .Z(n26476) );
  XOR U27816 ( .A(n26481), .B(n26145), .Z(n26147) );
  XOR U27817 ( .A(n26482), .B(n26483), .Z(n26145) );
  AND U27818 ( .A(n26484), .B(n26485), .Z(n26482) );
  AND U27819 ( .A(b[20]), .B(a[36]), .Z(n26481) );
  XOR U27820 ( .A(n26486), .B(n26150), .Z(n26152) );
  XOR U27821 ( .A(n26487), .B(n26488), .Z(n26150) );
  AND U27822 ( .A(n26489), .B(n26490), .Z(n26487) );
  AND U27823 ( .A(b[19]), .B(a[37]), .Z(n26486) );
  XOR U27824 ( .A(n26491), .B(n26155), .Z(n26157) );
  XOR U27825 ( .A(n26492), .B(n26493), .Z(n26155) );
  AND U27826 ( .A(n26494), .B(n26495), .Z(n26492) );
  AND U27827 ( .A(b[18]), .B(a[38]), .Z(n26491) );
  XOR U27828 ( .A(n26496), .B(n26160), .Z(n26162) );
  XOR U27829 ( .A(n26497), .B(n26498), .Z(n26160) );
  AND U27830 ( .A(n26499), .B(n26500), .Z(n26497) );
  AND U27831 ( .A(b[17]), .B(a[39]), .Z(n26496) );
  XOR U27832 ( .A(n26501), .B(n26165), .Z(n26167) );
  XOR U27833 ( .A(n26502), .B(n26503), .Z(n26165) );
  AND U27834 ( .A(n26504), .B(n26505), .Z(n26502) );
  AND U27835 ( .A(b[16]), .B(a[40]), .Z(n26501) );
  XOR U27836 ( .A(n26506), .B(n26170), .Z(n26172) );
  XOR U27837 ( .A(n26507), .B(n26508), .Z(n26170) );
  AND U27838 ( .A(n26509), .B(n26510), .Z(n26507) );
  AND U27839 ( .A(b[15]), .B(a[41]), .Z(n26506) );
  XOR U27840 ( .A(n26511), .B(n26175), .Z(n26177) );
  XOR U27841 ( .A(n26512), .B(n26513), .Z(n26175) );
  AND U27842 ( .A(n26514), .B(n26515), .Z(n26512) );
  AND U27843 ( .A(b[14]), .B(a[42]), .Z(n26511) );
  XOR U27844 ( .A(n26516), .B(n26180), .Z(n26182) );
  XOR U27845 ( .A(n26517), .B(n26518), .Z(n26180) );
  AND U27846 ( .A(n26519), .B(n26520), .Z(n26517) );
  AND U27847 ( .A(b[13]), .B(a[43]), .Z(n26516) );
  XOR U27848 ( .A(n26521), .B(n26185), .Z(n26187) );
  XOR U27849 ( .A(n26522), .B(n26523), .Z(n26185) );
  AND U27850 ( .A(n26524), .B(n26525), .Z(n26522) );
  AND U27851 ( .A(b[12]), .B(a[44]), .Z(n26521) );
  XOR U27852 ( .A(n26526), .B(n26190), .Z(n26192) );
  XOR U27853 ( .A(n26527), .B(n26528), .Z(n26190) );
  AND U27854 ( .A(n26529), .B(n26530), .Z(n26527) );
  AND U27855 ( .A(b[11]), .B(a[45]), .Z(n26526) );
  XOR U27856 ( .A(n26531), .B(n26195), .Z(n26197) );
  XOR U27857 ( .A(n26532), .B(n26533), .Z(n26195) );
  AND U27858 ( .A(n26534), .B(n26535), .Z(n26532) );
  AND U27859 ( .A(b[10]), .B(a[46]), .Z(n26531) );
  XOR U27860 ( .A(n26536), .B(n26200), .Z(n26202) );
  XOR U27861 ( .A(n26537), .B(n26538), .Z(n26200) );
  AND U27862 ( .A(n26539), .B(n26540), .Z(n26537) );
  AND U27863 ( .A(b[9]), .B(a[47]), .Z(n26536) );
  XOR U27864 ( .A(n26541), .B(n26205), .Z(n26207) );
  XOR U27865 ( .A(n26542), .B(n26543), .Z(n26205) );
  AND U27866 ( .A(n26544), .B(n26545), .Z(n26542) );
  AND U27867 ( .A(b[8]), .B(a[48]), .Z(n26541) );
  XOR U27868 ( .A(n26546), .B(n26210), .Z(n26212) );
  XOR U27869 ( .A(n26547), .B(n26548), .Z(n26210) );
  AND U27870 ( .A(n26549), .B(n26550), .Z(n26547) );
  AND U27871 ( .A(b[7]), .B(a[49]), .Z(n26546) );
  XOR U27872 ( .A(n26551), .B(n26215), .Z(n26217) );
  XOR U27873 ( .A(n26552), .B(n26553), .Z(n26215) );
  AND U27874 ( .A(n26554), .B(n26555), .Z(n26552) );
  AND U27875 ( .A(b[6]), .B(a[50]), .Z(n26551) );
  XOR U27876 ( .A(n26556), .B(n26220), .Z(n26222) );
  XOR U27877 ( .A(n26557), .B(n26558), .Z(n26220) );
  AND U27878 ( .A(n26559), .B(n26560), .Z(n26557) );
  AND U27879 ( .A(b[5]), .B(a[51]), .Z(n26556) );
  XOR U27880 ( .A(n26561), .B(n26225), .Z(n26227) );
  XOR U27881 ( .A(n26562), .B(n26563), .Z(n26225) );
  AND U27882 ( .A(n26564), .B(n26565), .Z(n26562) );
  AND U27883 ( .A(b[4]), .B(a[52]), .Z(n26561) );
  XNOR U27884 ( .A(n26566), .B(n26567), .Z(n26239) );
  NANDN U27885 ( .A(n26568), .B(n26569), .Z(n26567) );
  XOR U27886 ( .A(n26570), .B(n26230), .Z(n26232) );
  XNOR U27887 ( .A(n26571), .B(n26572), .Z(n26230) );
  AND U27888 ( .A(n26573), .B(n26574), .Z(n26571) );
  AND U27889 ( .A(b[3]), .B(a[53]), .Z(n26570) );
  XOR U27890 ( .A(n26246), .B(n26245), .Z(c[119]) );
  XOR U27891 ( .A(sreg[183]), .B(n26244), .Z(n26245) );
  XOR U27892 ( .A(n26251), .B(n26575), .Z(n26246) );
  XNOR U27893 ( .A(n26250), .B(n26244), .Z(n26575) );
  XOR U27894 ( .A(n26576), .B(n26577), .Z(n26244) );
  NOR U27895 ( .A(n26578), .B(n26579), .Z(n26576) );
  NAND U27896 ( .A(a[55]), .B(b[0]), .Z(n26250) );
  XNOR U27897 ( .A(n26568), .B(n26569), .Z(n26251) );
  XOR U27898 ( .A(n26566), .B(n26580), .Z(n26569) );
  NAND U27899 ( .A(b[1]), .B(a[54]), .Z(n26580) );
  XOR U27900 ( .A(n26574), .B(n26581), .Z(n26568) );
  XOR U27901 ( .A(n26566), .B(n26573), .Z(n26581) );
  XNOR U27902 ( .A(n26582), .B(n26572), .Z(n26573) );
  AND U27903 ( .A(b[2]), .B(a[53]), .Z(n26582) );
  NANDN U27904 ( .A(n26583), .B(n26584), .Z(n26566) );
  XOR U27905 ( .A(n26572), .B(n26564), .Z(n26585) );
  XNOR U27906 ( .A(n26563), .B(n26559), .Z(n26586) );
  XNOR U27907 ( .A(n26558), .B(n26554), .Z(n26587) );
  XNOR U27908 ( .A(n26553), .B(n26549), .Z(n26588) );
  XNOR U27909 ( .A(n26548), .B(n26544), .Z(n26589) );
  XNOR U27910 ( .A(n26543), .B(n26539), .Z(n26590) );
  XNOR U27911 ( .A(n26538), .B(n26534), .Z(n26591) );
  XNOR U27912 ( .A(n26533), .B(n26529), .Z(n26592) );
  XNOR U27913 ( .A(n26528), .B(n26524), .Z(n26593) );
  XNOR U27914 ( .A(n26523), .B(n26519), .Z(n26594) );
  XNOR U27915 ( .A(n26518), .B(n26514), .Z(n26595) );
  XNOR U27916 ( .A(n26513), .B(n26509), .Z(n26596) );
  XNOR U27917 ( .A(n26508), .B(n26504), .Z(n26597) );
  XNOR U27918 ( .A(n26503), .B(n26499), .Z(n26598) );
  XNOR U27919 ( .A(n26498), .B(n26494), .Z(n26599) );
  XNOR U27920 ( .A(n26493), .B(n26489), .Z(n26600) );
  XNOR U27921 ( .A(n26488), .B(n26484), .Z(n26601) );
  XNOR U27922 ( .A(n26483), .B(n26479), .Z(n26602) );
  XNOR U27923 ( .A(n26478), .B(n26474), .Z(n26603) );
  XNOR U27924 ( .A(n26473), .B(n26469), .Z(n26604) );
  XNOR U27925 ( .A(n26468), .B(n26464), .Z(n26605) );
  XNOR U27926 ( .A(n26463), .B(n26459), .Z(n26606) );
  XNOR U27927 ( .A(n26458), .B(n26454), .Z(n26607) );
  XNOR U27928 ( .A(n26453), .B(n26449), .Z(n26608) );
  XNOR U27929 ( .A(n26448), .B(n26444), .Z(n26609) );
  XNOR U27930 ( .A(n26443), .B(n26439), .Z(n26610) );
  XNOR U27931 ( .A(n26438), .B(n26434), .Z(n26611) );
  XNOR U27932 ( .A(n26433), .B(n26429), .Z(n26612) );
  XNOR U27933 ( .A(n26428), .B(n26424), .Z(n26613) );
  XNOR U27934 ( .A(n26423), .B(n26419), .Z(n26614) );
  XNOR U27935 ( .A(n26418), .B(n26414), .Z(n26615) );
  XNOR U27936 ( .A(n26413), .B(n26409), .Z(n26616) );
  XNOR U27937 ( .A(n26408), .B(n26404), .Z(n26617) );
  XNOR U27938 ( .A(n26403), .B(n26399), .Z(n26618) );
  XNOR U27939 ( .A(n26398), .B(n26394), .Z(n26619) );
  XNOR U27940 ( .A(n26393), .B(n26389), .Z(n26620) );
  XNOR U27941 ( .A(n26388), .B(n26384), .Z(n26621) );
  XNOR U27942 ( .A(n26383), .B(n26379), .Z(n26622) );
  XNOR U27943 ( .A(n26378), .B(n26374), .Z(n26623) );
  XNOR U27944 ( .A(n26373), .B(n26369), .Z(n26624) );
  XNOR U27945 ( .A(n26368), .B(n26364), .Z(n26625) );
  XNOR U27946 ( .A(n26363), .B(n26359), .Z(n26626) );
  XNOR U27947 ( .A(n26358), .B(n26354), .Z(n26627) );
  XNOR U27948 ( .A(n26353), .B(n26349), .Z(n26628) );
  XNOR U27949 ( .A(n26348), .B(n26344), .Z(n26629) );
  XNOR U27950 ( .A(n26343), .B(n26339), .Z(n26630) );
  XNOR U27951 ( .A(n26338), .B(n26334), .Z(n26631) );
  XNOR U27952 ( .A(n26333), .B(n26329), .Z(n26632) );
  XNOR U27953 ( .A(n26328), .B(n26324), .Z(n26633) );
  XNOR U27954 ( .A(n26323), .B(n26319), .Z(n26634) );
  XNOR U27955 ( .A(n26318), .B(n26314), .Z(n26635) );
  XNOR U27956 ( .A(n26313), .B(n26309), .Z(n26636) );
  XOR U27957 ( .A(n26637), .B(n26308), .Z(n26309) );
  AND U27958 ( .A(a[0]), .B(b[55]), .Z(n26637) );
  XOR U27959 ( .A(n26638), .B(n26308), .Z(n26310) );
  XNOR U27960 ( .A(n26639), .B(n26640), .Z(n26308) );
  AND U27961 ( .A(n26641), .B(n26642), .Z(n26639) );
  AND U27962 ( .A(a[1]), .B(b[54]), .Z(n26638) );
  XOR U27963 ( .A(n26643), .B(n26313), .Z(n26315) );
  XOR U27964 ( .A(n26644), .B(n26645), .Z(n26313) );
  AND U27965 ( .A(n26646), .B(n26647), .Z(n26644) );
  AND U27966 ( .A(a[2]), .B(b[53]), .Z(n26643) );
  XOR U27967 ( .A(n26648), .B(n26318), .Z(n26320) );
  XOR U27968 ( .A(n26649), .B(n26650), .Z(n26318) );
  AND U27969 ( .A(n26651), .B(n26652), .Z(n26649) );
  AND U27970 ( .A(a[3]), .B(b[52]), .Z(n26648) );
  XOR U27971 ( .A(n26653), .B(n26323), .Z(n26325) );
  XOR U27972 ( .A(n26654), .B(n26655), .Z(n26323) );
  AND U27973 ( .A(n26656), .B(n26657), .Z(n26654) );
  AND U27974 ( .A(a[4]), .B(b[51]), .Z(n26653) );
  XOR U27975 ( .A(n26658), .B(n26328), .Z(n26330) );
  XOR U27976 ( .A(n26659), .B(n26660), .Z(n26328) );
  AND U27977 ( .A(n26661), .B(n26662), .Z(n26659) );
  AND U27978 ( .A(a[5]), .B(b[50]), .Z(n26658) );
  XOR U27979 ( .A(n26663), .B(n26333), .Z(n26335) );
  XOR U27980 ( .A(n26664), .B(n26665), .Z(n26333) );
  AND U27981 ( .A(n26666), .B(n26667), .Z(n26664) );
  AND U27982 ( .A(a[6]), .B(b[49]), .Z(n26663) );
  XOR U27983 ( .A(n26668), .B(n26338), .Z(n26340) );
  XOR U27984 ( .A(n26669), .B(n26670), .Z(n26338) );
  AND U27985 ( .A(n26671), .B(n26672), .Z(n26669) );
  AND U27986 ( .A(a[7]), .B(b[48]), .Z(n26668) );
  XOR U27987 ( .A(n26673), .B(n26343), .Z(n26345) );
  XOR U27988 ( .A(n26674), .B(n26675), .Z(n26343) );
  AND U27989 ( .A(n26676), .B(n26677), .Z(n26674) );
  AND U27990 ( .A(a[8]), .B(b[47]), .Z(n26673) );
  XOR U27991 ( .A(n26678), .B(n26348), .Z(n26350) );
  XOR U27992 ( .A(n26679), .B(n26680), .Z(n26348) );
  AND U27993 ( .A(n26681), .B(n26682), .Z(n26679) );
  AND U27994 ( .A(a[9]), .B(b[46]), .Z(n26678) );
  XOR U27995 ( .A(n26683), .B(n26353), .Z(n26355) );
  XOR U27996 ( .A(n26684), .B(n26685), .Z(n26353) );
  AND U27997 ( .A(n26686), .B(n26687), .Z(n26684) );
  AND U27998 ( .A(a[10]), .B(b[45]), .Z(n26683) );
  XOR U27999 ( .A(n26688), .B(n26358), .Z(n26360) );
  XOR U28000 ( .A(n26689), .B(n26690), .Z(n26358) );
  AND U28001 ( .A(n26691), .B(n26692), .Z(n26689) );
  AND U28002 ( .A(a[11]), .B(b[44]), .Z(n26688) );
  XOR U28003 ( .A(n26693), .B(n26363), .Z(n26365) );
  XOR U28004 ( .A(n26694), .B(n26695), .Z(n26363) );
  AND U28005 ( .A(n26696), .B(n26697), .Z(n26694) );
  AND U28006 ( .A(a[12]), .B(b[43]), .Z(n26693) );
  XOR U28007 ( .A(n26698), .B(n26368), .Z(n26370) );
  XOR U28008 ( .A(n26699), .B(n26700), .Z(n26368) );
  AND U28009 ( .A(n26701), .B(n26702), .Z(n26699) );
  AND U28010 ( .A(a[13]), .B(b[42]), .Z(n26698) );
  XOR U28011 ( .A(n26703), .B(n26373), .Z(n26375) );
  XOR U28012 ( .A(n26704), .B(n26705), .Z(n26373) );
  AND U28013 ( .A(n26706), .B(n26707), .Z(n26704) );
  AND U28014 ( .A(a[14]), .B(b[41]), .Z(n26703) );
  XOR U28015 ( .A(n26708), .B(n26378), .Z(n26380) );
  XOR U28016 ( .A(n26709), .B(n26710), .Z(n26378) );
  AND U28017 ( .A(n26711), .B(n26712), .Z(n26709) );
  AND U28018 ( .A(a[15]), .B(b[40]), .Z(n26708) );
  XOR U28019 ( .A(n26713), .B(n26383), .Z(n26385) );
  XOR U28020 ( .A(n26714), .B(n26715), .Z(n26383) );
  AND U28021 ( .A(n26716), .B(n26717), .Z(n26714) );
  AND U28022 ( .A(a[16]), .B(b[39]), .Z(n26713) );
  XOR U28023 ( .A(n26718), .B(n26388), .Z(n26390) );
  XOR U28024 ( .A(n26719), .B(n26720), .Z(n26388) );
  AND U28025 ( .A(n26721), .B(n26722), .Z(n26719) );
  AND U28026 ( .A(a[17]), .B(b[38]), .Z(n26718) );
  XOR U28027 ( .A(n26723), .B(n26393), .Z(n26395) );
  XOR U28028 ( .A(n26724), .B(n26725), .Z(n26393) );
  AND U28029 ( .A(n26726), .B(n26727), .Z(n26724) );
  AND U28030 ( .A(a[18]), .B(b[37]), .Z(n26723) );
  XOR U28031 ( .A(n26728), .B(n26398), .Z(n26400) );
  XOR U28032 ( .A(n26729), .B(n26730), .Z(n26398) );
  AND U28033 ( .A(n26731), .B(n26732), .Z(n26729) );
  AND U28034 ( .A(a[19]), .B(b[36]), .Z(n26728) );
  XOR U28035 ( .A(n26733), .B(n26403), .Z(n26405) );
  XOR U28036 ( .A(n26734), .B(n26735), .Z(n26403) );
  AND U28037 ( .A(n26736), .B(n26737), .Z(n26734) );
  AND U28038 ( .A(a[20]), .B(b[35]), .Z(n26733) );
  XOR U28039 ( .A(n26738), .B(n26408), .Z(n26410) );
  XOR U28040 ( .A(n26739), .B(n26740), .Z(n26408) );
  AND U28041 ( .A(n26741), .B(n26742), .Z(n26739) );
  AND U28042 ( .A(a[21]), .B(b[34]), .Z(n26738) );
  XOR U28043 ( .A(n26743), .B(n26413), .Z(n26415) );
  XOR U28044 ( .A(n26744), .B(n26745), .Z(n26413) );
  AND U28045 ( .A(n26746), .B(n26747), .Z(n26744) );
  AND U28046 ( .A(a[22]), .B(b[33]), .Z(n26743) );
  XOR U28047 ( .A(n26748), .B(n26418), .Z(n26420) );
  XOR U28048 ( .A(n26749), .B(n26750), .Z(n26418) );
  AND U28049 ( .A(n26751), .B(n26752), .Z(n26749) );
  AND U28050 ( .A(a[23]), .B(b[32]), .Z(n26748) );
  XOR U28051 ( .A(n26753), .B(n26423), .Z(n26425) );
  XOR U28052 ( .A(n26754), .B(n26755), .Z(n26423) );
  AND U28053 ( .A(n26756), .B(n26757), .Z(n26754) );
  AND U28054 ( .A(a[24]), .B(b[31]), .Z(n26753) );
  XOR U28055 ( .A(n26758), .B(n26428), .Z(n26430) );
  XOR U28056 ( .A(n26759), .B(n26760), .Z(n26428) );
  AND U28057 ( .A(n26761), .B(n26762), .Z(n26759) );
  AND U28058 ( .A(a[25]), .B(b[30]), .Z(n26758) );
  XOR U28059 ( .A(n26763), .B(n26433), .Z(n26435) );
  XOR U28060 ( .A(n26764), .B(n26765), .Z(n26433) );
  AND U28061 ( .A(n26766), .B(n26767), .Z(n26764) );
  AND U28062 ( .A(a[26]), .B(b[29]), .Z(n26763) );
  XOR U28063 ( .A(n26768), .B(n26438), .Z(n26440) );
  XOR U28064 ( .A(n26769), .B(n26770), .Z(n26438) );
  AND U28065 ( .A(n26771), .B(n26772), .Z(n26769) );
  AND U28066 ( .A(a[27]), .B(b[28]), .Z(n26768) );
  XOR U28067 ( .A(n26773), .B(n26443), .Z(n26445) );
  XOR U28068 ( .A(n26774), .B(n26775), .Z(n26443) );
  AND U28069 ( .A(n26776), .B(n26777), .Z(n26774) );
  AND U28070 ( .A(b[27]), .B(a[28]), .Z(n26773) );
  XOR U28071 ( .A(n26778), .B(n26448), .Z(n26450) );
  XOR U28072 ( .A(n26779), .B(n26780), .Z(n26448) );
  AND U28073 ( .A(n26781), .B(n26782), .Z(n26779) );
  AND U28074 ( .A(b[26]), .B(a[29]), .Z(n26778) );
  XOR U28075 ( .A(n26783), .B(n26453), .Z(n26455) );
  XOR U28076 ( .A(n26784), .B(n26785), .Z(n26453) );
  AND U28077 ( .A(n26786), .B(n26787), .Z(n26784) );
  AND U28078 ( .A(b[25]), .B(a[30]), .Z(n26783) );
  XOR U28079 ( .A(n26788), .B(n26458), .Z(n26460) );
  XOR U28080 ( .A(n26789), .B(n26790), .Z(n26458) );
  AND U28081 ( .A(n26791), .B(n26792), .Z(n26789) );
  AND U28082 ( .A(b[24]), .B(a[31]), .Z(n26788) );
  XOR U28083 ( .A(n26793), .B(n26463), .Z(n26465) );
  XOR U28084 ( .A(n26794), .B(n26795), .Z(n26463) );
  AND U28085 ( .A(n26796), .B(n26797), .Z(n26794) );
  AND U28086 ( .A(b[23]), .B(a[32]), .Z(n26793) );
  XOR U28087 ( .A(n26798), .B(n26468), .Z(n26470) );
  XOR U28088 ( .A(n26799), .B(n26800), .Z(n26468) );
  AND U28089 ( .A(n26801), .B(n26802), .Z(n26799) );
  AND U28090 ( .A(b[22]), .B(a[33]), .Z(n26798) );
  XOR U28091 ( .A(n26803), .B(n26473), .Z(n26475) );
  XOR U28092 ( .A(n26804), .B(n26805), .Z(n26473) );
  AND U28093 ( .A(n26806), .B(n26807), .Z(n26804) );
  AND U28094 ( .A(b[21]), .B(a[34]), .Z(n26803) );
  XOR U28095 ( .A(n26808), .B(n26478), .Z(n26480) );
  XOR U28096 ( .A(n26809), .B(n26810), .Z(n26478) );
  AND U28097 ( .A(n26811), .B(n26812), .Z(n26809) );
  AND U28098 ( .A(b[20]), .B(a[35]), .Z(n26808) );
  XOR U28099 ( .A(n26813), .B(n26483), .Z(n26485) );
  XOR U28100 ( .A(n26814), .B(n26815), .Z(n26483) );
  AND U28101 ( .A(n26816), .B(n26817), .Z(n26814) );
  AND U28102 ( .A(b[19]), .B(a[36]), .Z(n26813) );
  XOR U28103 ( .A(n26818), .B(n26488), .Z(n26490) );
  XOR U28104 ( .A(n26819), .B(n26820), .Z(n26488) );
  AND U28105 ( .A(n26821), .B(n26822), .Z(n26819) );
  AND U28106 ( .A(b[18]), .B(a[37]), .Z(n26818) );
  XOR U28107 ( .A(n26823), .B(n26493), .Z(n26495) );
  XOR U28108 ( .A(n26824), .B(n26825), .Z(n26493) );
  AND U28109 ( .A(n26826), .B(n26827), .Z(n26824) );
  AND U28110 ( .A(b[17]), .B(a[38]), .Z(n26823) );
  XOR U28111 ( .A(n26828), .B(n26498), .Z(n26500) );
  XOR U28112 ( .A(n26829), .B(n26830), .Z(n26498) );
  AND U28113 ( .A(n26831), .B(n26832), .Z(n26829) );
  AND U28114 ( .A(b[16]), .B(a[39]), .Z(n26828) );
  XOR U28115 ( .A(n26833), .B(n26503), .Z(n26505) );
  XOR U28116 ( .A(n26834), .B(n26835), .Z(n26503) );
  AND U28117 ( .A(n26836), .B(n26837), .Z(n26834) );
  AND U28118 ( .A(b[15]), .B(a[40]), .Z(n26833) );
  XOR U28119 ( .A(n26838), .B(n26508), .Z(n26510) );
  XOR U28120 ( .A(n26839), .B(n26840), .Z(n26508) );
  AND U28121 ( .A(n26841), .B(n26842), .Z(n26839) );
  AND U28122 ( .A(b[14]), .B(a[41]), .Z(n26838) );
  XOR U28123 ( .A(n26843), .B(n26513), .Z(n26515) );
  XOR U28124 ( .A(n26844), .B(n26845), .Z(n26513) );
  AND U28125 ( .A(n26846), .B(n26847), .Z(n26844) );
  AND U28126 ( .A(b[13]), .B(a[42]), .Z(n26843) );
  XOR U28127 ( .A(n26848), .B(n26518), .Z(n26520) );
  XOR U28128 ( .A(n26849), .B(n26850), .Z(n26518) );
  AND U28129 ( .A(n26851), .B(n26852), .Z(n26849) );
  AND U28130 ( .A(b[12]), .B(a[43]), .Z(n26848) );
  XOR U28131 ( .A(n26853), .B(n26523), .Z(n26525) );
  XOR U28132 ( .A(n26854), .B(n26855), .Z(n26523) );
  AND U28133 ( .A(n26856), .B(n26857), .Z(n26854) );
  AND U28134 ( .A(b[11]), .B(a[44]), .Z(n26853) );
  XOR U28135 ( .A(n26858), .B(n26528), .Z(n26530) );
  XOR U28136 ( .A(n26859), .B(n26860), .Z(n26528) );
  AND U28137 ( .A(n26861), .B(n26862), .Z(n26859) );
  AND U28138 ( .A(b[10]), .B(a[45]), .Z(n26858) );
  XOR U28139 ( .A(n26863), .B(n26533), .Z(n26535) );
  XOR U28140 ( .A(n26864), .B(n26865), .Z(n26533) );
  AND U28141 ( .A(n26866), .B(n26867), .Z(n26864) );
  AND U28142 ( .A(b[9]), .B(a[46]), .Z(n26863) );
  XOR U28143 ( .A(n26868), .B(n26538), .Z(n26540) );
  XOR U28144 ( .A(n26869), .B(n26870), .Z(n26538) );
  AND U28145 ( .A(n26871), .B(n26872), .Z(n26869) );
  AND U28146 ( .A(b[8]), .B(a[47]), .Z(n26868) );
  XOR U28147 ( .A(n26873), .B(n26543), .Z(n26545) );
  XOR U28148 ( .A(n26874), .B(n26875), .Z(n26543) );
  AND U28149 ( .A(n26876), .B(n26877), .Z(n26874) );
  AND U28150 ( .A(b[7]), .B(a[48]), .Z(n26873) );
  XOR U28151 ( .A(n26878), .B(n26548), .Z(n26550) );
  XOR U28152 ( .A(n26879), .B(n26880), .Z(n26548) );
  AND U28153 ( .A(n26881), .B(n26882), .Z(n26879) );
  AND U28154 ( .A(b[6]), .B(a[49]), .Z(n26878) );
  XOR U28155 ( .A(n26883), .B(n26553), .Z(n26555) );
  XOR U28156 ( .A(n26884), .B(n26885), .Z(n26553) );
  AND U28157 ( .A(n26886), .B(n26887), .Z(n26884) );
  AND U28158 ( .A(b[5]), .B(a[50]), .Z(n26883) );
  XOR U28159 ( .A(n26888), .B(n26558), .Z(n26560) );
  XOR U28160 ( .A(n26889), .B(n26890), .Z(n26558) );
  AND U28161 ( .A(n26891), .B(n26892), .Z(n26889) );
  AND U28162 ( .A(b[4]), .B(a[51]), .Z(n26888) );
  XNOR U28163 ( .A(n26893), .B(n26894), .Z(n26572) );
  NANDN U28164 ( .A(n26895), .B(n26896), .Z(n26894) );
  XOR U28165 ( .A(n26897), .B(n26563), .Z(n26565) );
  XNOR U28166 ( .A(n26898), .B(n26899), .Z(n26563) );
  AND U28167 ( .A(n26900), .B(n26901), .Z(n26898) );
  AND U28168 ( .A(b[3]), .B(a[52]), .Z(n26897) );
  XOR U28169 ( .A(n26579), .B(n26578), .Z(c[118]) );
  XOR U28170 ( .A(sreg[182]), .B(n26577), .Z(n26578) );
  XOR U28171 ( .A(n26584), .B(n26902), .Z(n26579) );
  XNOR U28172 ( .A(n26583), .B(n26577), .Z(n26902) );
  XOR U28173 ( .A(n26903), .B(n26904), .Z(n26577) );
  NOR U28174 ( .A(n26905), .B(n26906), .Z(n26903) );
  NAND U28175 ( .A(a[54]), .B(b[0]), .Z(n26583) );
  XNOR U28176 ( .A(n26895), .B(n26896), .Z(n26584) );
  XOR U28177 ( .A(n26893), .B(n26907), .Z(n26896) );
  NAND U28178 ( .A(b[1]), .B(a[53]), .Z(n26907) );
  XOR U28179 ( .A(n26901), .B(n26908), .Z(n26895) );
  XOR U28180 ( .A(n26893), .B(n26900), .Z(n26908) );
  XNOR U28181 ( .A(n26909), .B(n26899), .Z(n26900) );
  AND U28182 ( .A(b[2]), .B(a[52]), .Z(n26909) );
  NANDN U28183 ( .A(n26910), .B(n26911), .Z(n26893) );
  XOR U28184 ( .A(n26899), .B(n26891), .Z(n26912) );
  XNOR U28185 ( .A(n26890), .B(n26886), .Z(n26913) );
  XNOR U28186 ( .A(n26885), .B(n26881), .Z(n26914) );
  XNOR U28187 ( .A(n26880), .B(n26876), .Z(n26915) );
  XNOR U28188 ( .A(n26875), .B(n26871), .Z(n26916) );
  XNOR U28189 ( .A(n26870), .B(n26866), .Z(n26917) );
  XNOR U28190 ( .A(n26865), .B(n26861), .Z(n26918) );
  XNOR U28191 ( .A(n26860), .B(n26856), .Z(n26919) );
  XNOR U28192 ( .A(n26855), .B(n26851), .Z(n26920) );
  XNOR U28193 ( .A(n26850), .B(n26846), .Z(n26921) );
  XNOR U28194 ( .A(n26845), .B(n26841), .Z(n26922) );
  XNOR U28195 ( .A(n26840), .B(n26836), .Z(n26923) );
  XNOR U28196 ( .A(n26835), .B(n26831), .Z(n26924) );
  XNOR U28197 ( .A(n26830), .B(n26826), .Z(n26925) );
  XNOR U28198 ( .A(n26825), .B(n26821), .Z(n26926) );
  XNOR U28199 ( .A(n26820), .B(n26816), .Z(n26927) );
  XNOR U28200 ( .A(n26815), .B(n26811), .Z(n26928) );
  XNOR U28201 ( .A(n26810), .B(n26806), .Z(n26929) );
  XNOR U28202 ( .A(n26805), .B(n26801), .Z(n26930) );
  XNOR U28203 ( .A(n26800), .B(n26796), .Z(n26931) );
  XNOR U28204 ( .A(n26795), .B(n26791), .Z(n26932) );
  XNOR U28205 ( .A(n26790), .B(n26786), .Z(n26933) );
  XNOR U28206 ( .A(n26785), .B(n26781), .Z(n26934) );
  XNOR U28207 ( .A(n26780), .B(n26776), .Z(n26935) );
  XNOR U28208 ( .A(n26775), .B(n26771), .Z(n26936) );
  XNOR U28209 ( .A(n26770), .B(n26766), .Z(n26937) );
  XNOR U28210 ( .A(n26765), .B(n26761), .Z(n26938) );
  XNOR U28211 ( .A(n26760), .B(n26756), .Z(n26939) );
  XNOR U28212 ( .A(n26755), .B(n26751), .Z(n26940) );
  XNOR U28213 ( .A(n26750), .B(n26746), .Z(n26941) );
  XNOR U28214 ( .A(n26745), .B(n26741), .Z(n26942) );
  XNOR U28215 ( .A(n26740), .B(n26736), .Z(n26943) );
  XNOR U28216 ( .A(n26735), .B(n26731), .Z(n26944) );
  XNOR U28217 ( .A(n26730), .B(n26726), .Z(n26945) );
  XNOR U28218 ( .A(n26725), .B(n26721), .Z(n26946) );
  XNOR U28219 ( .A(n26720), .B(n26716), .Z(n26947) );
  XNOR U28220 ( .A(n26715), .B(n26711), .Z(n26948) );
  XNOR U28221 ( .A(n26710), .B(n26706), .Z(n26949) );
  XNOR U28222 ( .A(n26705), .B(n26701), .Z(n26950) );
  XNOR U28223 ( .A(n26700), .B(n26696), .Z(n26951) );
  XNOR U28224 ( .A(n26695), .B(n26691), .Z(n26952) );
  XNOR U28225 ( .A(n26690), .B(n26686), .Z(n26953) );
  XNOR U28226 ( .A(n26685), .B(n26681), .Z(n26954) );
  XNOR U28227 ( .A(n26680), .B(n26676), .Z(n26955) );
  XNOR U28228 ( .A(n26675), .B(n26671), .Z(n26956) );
  XNOR U28229 ( .A(n26670), .B(n26666), .Z(n26957) );
  XNOR U28230 ( .A(n26665), .B(n26661), .Z(n26958) );
  XNOR U28231 ( .A(n26660), .B(n26656), .Z(n26959) );
  XNOR U28232 ( .A(n26655), .B(n26651), .Z(n26960) );
  XNOR U28233 ( .A(n26650), .B(n26646), .Z(n26961) );
  XNOR U28234 ( .A(n26645), .B(n26641), .Z(n26962) );
  XNOR U28235 ( .A(n26963), .B(n26640), .Z(n26641) );
  AND U28236 ( .A(a[0]), .B(b[54]), .Z(n26963) );
  XNOR U28237 ( .A(n26964), .B(n26640), .Z(n26642) );
  XNOR U28238 ( .A(n26965), .B(n26966), .Z(n26640) );
  AND U28239 ( .A(n26967), .B(n26968), .Z(n26965) );
  AND U28240 ( .A(a[1]), .B(b[53]), .Z(n26964) );
  XOR U28241 ( .A(n26969), .B(n26645), .Z(n26647) );
  XOR U28242 ( .A(n26970), .B(n26971), .Z(n26645) );
  AND U28243 ( .A(n26972), .B(n26973), .Z(n26970) );
  AND U28244 ( .A(a[2]), .B(b[52]), .Z(n26969) );
  XOR U28245 ( .A(n26974), .B(n26650), .Z(n26652) );
  XOR U28246 ( .A(n26975), .B(n26976), .Z(n26650) );
  AND U28247 ( .A(n26977), .B(n26978), .Z(n26975) );
  AND U28248 ( .A(a[3]), .B(b[51]), .Z(n26974) );
  XOR U28249 ( .A(n26979), .B(n26655), .Z(n26657) );
  XOR U28250 ( .A(n26980), .B(n26981), .Z(n26655) );
  AND U28251 ( .A(n26982), .B(n26983), .Z(n26980) );
  AND U28252 ( .A(a[4]), .B(b[50]), .Z(n26979) );
  XOR U28253 ( .A(n26984), .B(n26660), .Z(n26662) );
  XOR U28254 ( .A(n26985), .B(n26986), .Z(n26660) );
  AND U28255 ( .A(n26987), .B(n26988), .Z(n26985) );
  AND U28256 ( .A(a[5]), .B(b[49]), .Z(n26984) );
  XOR U28257 ( .A(n26989), .B(n26665), .Z(n26667) );
  XOR U28258 ( .A(n26990), .B(n26991), .Z(n26665) );
  AND U28259 ( .A(n26992), .B(n26993), .Z(n26990) );
  AND U28260 ( .A(a[6]), .B(b[48]), .Z(n26989) );
  XOR U28261 ( .A(n26994), .B(n26670), .Z(n26672) );
  XOR U28262 ( .A(n26995), .B(n26996), .Z(n26670) );
  AND U28263 ( .A(n26997), .B(n26998), .Z(n26995) );
  AND U28264 ( .A(a[7]), .B(b[47]), .Z(n26994) );
  XOR U28265 ( .A(n26999), .B(n26675), .Z(n26677) );
  XOR U28266 ( .A(n27000), .B(n27001), .Z(n26675) );
  AND U28267 ( .A(n27002), .B(n27003), .Z(n27000) );
  AND U28268 ( .A(a[8]), .B(b[46]), .Z(n26999) );
  XOR U28269 ( .A(n27004), .B(n26680), .Z(n26682) );
  XOR U28270 ( .A(n27005), .B(n27006), .Z(n26680) );
  AND U28271 ( .A(n27007), .B(n27008), .Z(n27005) );
  AND U28272 ( .A(a[9]), .B(b[45]), .Z(n27004) );
  XOR U28273 ( .A(n27009), .B(n26685), .Z(n26687) );
  XOR U28274 ( .A(n27010), .B(n27011), .Z(n26685) );
  AND U28275 ( .A(n27012), .B(n27013), .Z(n27010) );
  AND U28276 ( .A(a[10]), .B(b[44]), .Z(n27009) );
  XOR U28277 ( .A(n27014), .B(n26690), .Z(n26692) );
  XOR U28278 ( .A(n27015), .B(n27016), .Z(n26690) );
  AND U28279 ( .A(n27017), .B(n27018), .Z(n27015) );
  AND U28280 ( .A(a[11]), .B(b[43]), .Z(n27014) );
  XOR U28281 ( .A(n27019), .B(n26695), .Z(n26697) );
  XOR U28282 ( .A(n27020), .B(n27021), .Z(n26695) );
  AND U28283 ( .A(n27022), .B(n27023), .Z(n27020) );
  AND U28284 ( .A(a[12]), .B(b[42]), .Z(n27019) );
  XOR U28285 ( .A(n27024), .B(n26700), .Z(n26702) );
  XOR U28286 ( .A(n27025), .B(n27026), .Z(n26700) );
  AND U28287 ( .A(n27027), .B(n27028), .Z(n27025) );
  AND U28288 ( .A(a[13]), .B(b[41]), .Z(n27024) );
  XOR U28289 ( .A(n27029), .B(n26705), .Z(n26707) );
  XOR U28290 ( .A(n27030), .B(n27031), .Z(n26705) );
  AND U28291 ( .A(n27032), .B(n27033), .Z(n27030) );
  AND U28292 ( .A(a[14]), .B(b[40]), .Z(n27029) );
  XOR U28293 ( .A(n27034), .B(n26710), .Z(n26712) );
  XOR U28294 ( .A(n27035), .B(n27036), .Z(n26710) );
  AND U28295 ( .A(n27037), .B(n27038), .Z(n27035) );
  AND U28296 ( .A(a[15]), .B(b[39]), .Z(n27034) );
  XOR U28297 ( .A(n27039), .B(n26715), .Z(n26717) );
  XOR U28298 ( .A(n27040), .B(n27041), .Z(n26715) );
  AND U28299 ( .A(n27042), .B(n27043), .Z(n27040) );
  AND U28300 ( .A(a[16]), .B(b[38]), .Z(n27039) );
  XOR U28301 ( .A(n27044), .B(n26720), .Z(n26722) );
  XOR U28302 ( .A(n27045), .B(n27046), .Z(n26720) );
  AND U28303 ( .A(n27047), .B(n27048), .Z(n27045) );
  AND U28304 ( .A(a[17]), .B(b[37]), .Z(n27044) );
  XOR U28305 ( .A(n27049), .B(n26725), .Z(n26727) );
  XOR U28306 ( .A(n27050), .B(n27051), .Z(n26725) );
  AND U28307 ( .A(n27052), .B(n27053), .Z(n27050) );
  AND U28308 ( .A(a[18]), .B(b[36]), .Z(n27049) );
  XOR U28309 ( .A(n27054), .B(n26730), .Z(n26732) );
  XOR U28310 ( .A(n27055), .B(n27056), .Z(n26730) );
  AND U28311 ( .A(n27057), .B(n27058), .Z(n27055) );
  AND U28312 ( .A(a[19]), .B(b[35]), .Z(n27054) );
  XOR U28313 ( .A(n27059), .B(n26735), .Z(n26737) );
  XOR U28314 ( .A(n27060), .B(n27061), .Z(n26735) );
  AND U28315 ( .A(n27062), .B(n27063), .Z(n27060) );
  AND U28316 ( .A(a[20]), .B(b[34]), .Z(n27059) );
  XOR U28317 ( .A(n27064), .B(n26740), .Z(n26742) );
  XOR U28318 ( .A(n27065), .B(n27066), .Z(n26740) );
  AND U28319 ( .A(n27067), .B(n27068), .Z(n27065) );
  AND U28320 ( .A(a[21]), .B(b[33]), .Z(n27064) );
  XOR U28321 ( .A(n27069), .B(n26745), .Z(n26747) );
  XOR U28322 ( .A(n27070), .B(n27071), .Z(n26745) );
  AND U28323 ( .A(n27072), .B(n27073), .Z(n27070) );
  AND U28324 ( .A(a[22]), .B(b[32]), .Z(n27069) );
  XOR U28325 ( .A(n27074), .B(n26750), .Z(n26752) );
  XOR U28326 ( .A(n27075), .B(n27076), .Z(n26750) );
  AND U28327 ( .A(n27077), .B(n27078), .Z(n27075) );
  AND U28328 ( .A(a[23]), .B(b[31]), .Z(n27074) );
  XOR U28329 ( .A(n27079), .B(n26755), .Z(n26757) );
  XOR U28330 ( .A(n27080), .B(n27081), .Z(n26755) );
  AND U28331 ( .A(n27082), .B(n27083), .Z(n27080) );
  AND U28332 ( .A(a[24]), .B(b[30]), .Z(n27079) );
  XOR U28333 ( .A(n27084), .B(n26760), .Z(n26762) );
  XOR U28334 ( .A(n27085), .B(n27086), .Z(n26760) );
  AND U28335 ( .A(n27087), .B(n27088), .Z(n27085) );
  AND U28336 ( .A(a[25]), .B(b[29]), .Z(n27084) );
  XOR U28337 ( .A(n27089), .B(n26765), .Z(n26767) );
  XOR U28338 ( .A(n27090), .B(n27091), .Z(n26765) );
  AND U28339 ( .A(n27092), .B(n27093), .Z(n27090) );
  AND U28340 ( .A(a[26]), .B(b[28]), .Z(n27089) );
  XOR U28341 ( .A(n27094), .B(n26770), .Z(n26772) );
  XOR U28342 ( .A(n27095), .B(n27096), .Z(n26770) );
  AND U28343 ( .A(n27097), .B(n27098), .Z(n27095) );
  AND U28344 ( .A(a[27]), .B(b[27]), .Z(n27094) );
  XOR U28345 ( .A(n27099), .B(n26775), .Z(n26777) );
  XOR U28346 ( .A(n27100), .B(n27101), .Z(n26775) );
  AND U28347 ( .A(n27102), .B(n27103), .Z(n27100) );
  AND U28348 ( .A(b[26]), .B(a[28]), .Z(n27099) );
  XOR U28349 ( .A(n27104), .B(n26780), .Z(n26782) );
  XOR U28350 ( .A(n27105), .B(n27106), .Z(n26780) );
  AND U28351 ( .A(n27107), .B(n27108), .Z(n27105) );
  AND U28352 ( .A(b[25]), .B(a[29]), .Z(n27104) );
  XOR U28353 ( .A(n27109), .B(n26785), .Z(n26787) );
  XOR U28354 ( .A(n27110), .B(n27111), .Z(n26785) );
  AND U28355 ( .A(n27112), .B(n27113), .Z(n27110) );
  AND U28356 ( .A(b[24]), .B(a[30]), .Z(n27109) );
  XOR U28357 ( .A(n27114), .B(n26790), .Z(n26792) );
  XOR U28358 ( .A(n27115), .B(n27116), .Z(n26790) );
  AND U28359 ( .A(n27117), .B(n27118), .Z(n27115) );
  AND U28360 ( .A(b[23]), .B(a[31]), .Z(n27114) );
  XOR U28361 ( .A(n27119), .B(n26795), .Z(n26797) );
  XOR U28362 ( .A(n27120), .B(n27121), .Z(n26795) );
  AND U28363 ( .A(n27122), .B(n27123), .Z(n27120) );
  AND U28364 ( .A(b[22]), .B(a[32]), .Z(n27119) );
  XOR U28365 ( .A(n27124), .B(n26800), .Z(n26802) );
  XOR U28366 ( .A(n27125), .B(n27126), .Z(n26800) );
  AND U28367 ( .A(n27127), .B(n27128), .Z(n27125) );
  AND U28368 ( .A(b[21]), .B(a[33]), .Z(n27124) );
  XOR U28369 ( .A(n27129), .B(n26805), .Z(n26807) );
  XOR U28370 ( .A(n27130), .B(n27131), .Z(n26805) );
  AND U28371 ( .A(n27132), .B(n27133), .Z(n27130) );
  AND U28372 ( .A(b[20]), .B(a[34]), .Z(n27129) );
  XOR U28373 ( .A(n27134), .B(n26810), .Z(n26812) );
  XOR U28374 ( .A(n27135), .B(n27136), .Z(n26810) );
  AND U28375 ( .A(n27137), .B(n27138), .Z(n27135) );
  AND U28376 ( .A(b[19]), .B(a[35]), .Z(n27134) );
  XOR U28377 ( .A(n27139), .B(n26815), .Z(n26817) );
  XOR U28378 ( .A(n27140), .B(n27141), .Z(n26815) );
  AND U28379 ( .A(n27142), .B(n27143), .Z(n27140) );
  AND U28380 ( .A(b[18]), .B(a[36]), .Z(n27139) );
  XOR U28381 ( .A(n27144), .B(n26820), .Z(n26822) );
  XOR U28382 ( .A(n27145), .B(n27146), .Z(n26820) );
  AND U28383 ( .A(n27147), .B(n27148), .Z(n27145) );
  AND U28384 ( .A(b[17]), .B(a[37]), .Z(n27144) );
  XOR U28385 ( .A(n27149), .B(n26825), .Z(n26827) );
  XOR U28386 ( .A(n27150), .B(n27151), .Z(n26825) );
  AND U28387 ( .A(n27152), .B(n27153), .Z(n27150) );
  AND U28388 ( .A(b[16]), .B(a[38]), .Z(n27149) );
  XOR U28389 ( .A(n27154), .B(n26830), .Z(n26832) );
  XOR U28390 ( .A(n27155), .B(n27156), .Z(n26830) );
  AND U28391 ( .A(n27157), .B(n27158), .Z(n27155) );
  AND U28392 ( .A(b[15]), .B(a[39]), .Z(n27154) );
  XOR U28393 ( .A(n27159), .B(n26835), .Z(n26837) );
  XOR U28394 ( .A(n27160), .B(n27161), .Z(n26835) );
  AND U28395 ( .A(n27162), .B(n27163), .Z(n27160) );
  AND U28396 ( .A(b[14]), .B(a[40]), .Z(n27159) );
  XOR U28397 ( .A(n27164), .B(n26840), .Z(n26842) );
  XOR U28398 ( .A(n27165), .B(n27166), .Z(n26840) );
  AND U28399 ( .A(n27167), .B(n27168), .Z(n27165) );
  AND U28400 ( .A(b[13]), .B(a[41]), .Z(n27164) );
  XOR U28401 ( .A(n27169), .B(n26845), .Z(n26847) );
  XOR U28402 ( .A(n27170), .B(n27171), .Z(n26845) );
  AND U28403 ( .A(n27172), .B(n27173), .Z(n27170) );
  AND U28404 ( .A(b[12]), .B(a[42]), .Z(n27169) );
  XOR U28405 ( .A(n27174), .B(n26850), .Z(n26852) );
  XOR U28406 ( .A(n27175), .B(n27176), .Z(n26850) );
  AND U28407 ( .A(n27177), .B(n27178), .Z(n27175) );
  AND U28408 ( .A(b[11]), .B(a[43]), .Z(n27174) );
  XOR U28409 ( .A(n27179), .B(n26855), .Z(n26857) );
  XOR U28410 ( .A(n27180), .B(n27181), .Z(n26855) );
  AND U28411 ( .A(n27182), .B(n27183), .Z(n27180) );
  AND U28412 ( .A(b[10]), .B(a[44]), .Z(n27179) );
  XOR U28413 ( .A(n27184), .B(n26860), .Z(n26862) );
  XOR U28414 ( .A(n27185), .B(n27186), .Z(n26860) );
  AND U28415 ( .A(n27187), .B(n27188), .Z(n27185) );
  AND U28416 ( .A(b[9]), .B(a[45]), .Z(n27184) );
  XOR U28417 ( .A(n27189), .B(n26865), .Z(n26867) );
  XOR U28418 ( .A(n27190), .B(n27191), .Z(n26865) );
  AND U28419 ( .A(n27192), .B(n27193), .Z(n27190) );
  AND U28420 ( .A(b[8]), .B(a[46]), .Z(n27189) );
  XOR U28421 ( .A(n27194), .B(n26870), .Z(n26872) );
  XOR U28422 ( .A(n27195), .B(n27196), .Z(n26870) );
  AND U28423 ( .A(n27197), .B(n27198), .Z(n27195) );
  AND U28424 ( .A(b[7]), .B(a[47]), .Z(n27194) );
  XOR U28425 ( .A(n27199), .B(n26875), .Z(n26877) );
  XOR U28426 ( .A(n27200), .B(n27201), .Z(n26875) );
  AND U28427 ( .A(n27202), .B(n27203), .Z(n27200) );
  AND U28428 ( .A(b[6]), .B(a[48]), .Z(n27199) );
  XOR U28429 ( .A(n27204), .B(n26880), .Z(n26882) );
  XOR U28430 ( .A(n27205), .B(n27206), .Z(n26880) );
  AND U28431 ( .A(n27207), .B(n27208), .Z(n27205) );
  AND U28432 ( .A(b[5]), .B(a[49]), .Z(n27204) );
  XOR U28433 ( .A(n27209), .B(n26885), .Z(n26887) );
  XOR U28434 ( .A(n27210), .B(n27211), .Z(n26885) );
  AND U28435 ( .A(n27212), .B(n27213), .Z(n27210) );
  AND U28436 ( .A(b[4]), .B(a[50]), .Z(n27209) );
  XNOR U28437 ( .A(n27214), .B(n27215), .Z(n26899) );
  NANDN U28438 ( .A(n27216), .B(n27217), .Z(n27215) );
  XOR U28439 ( .A(n27218), .B(n26890), .Z(n26892) );
  XNOR U28440 ( .A(n27219), .B(n27220), .Z(n26890) );
  AND U28441 ( .A(n27221), .B(n27222), .Z(n27219) );
  AND U28442 ( .A(b[3]), .B(a[51]), .Z(n27218) );
  XOR U28443 ( .A(n26906), .B(n26905), .Z(c[117]) );
  XOR U28444 ( .A(sreg[181]), .B(n26904), .Z(n26905) );
  XOR U28445 ( .A(n26911), .B(n27223), .Z(n26906) );
  XNOR U28446 ( .A(n26910), .B(n26904), .Z(n27223) );
  XOR U28447 ( .A(n27224), .B(n27225), .Z(n26904) );
  NOR U28448 ( .A(n27226), .B(n27227), .Z(n27224) );
  NAND U28449 ( .A(a[53]), .B(b[0]), .Z(n26910) );
  XNOR U28450 ( .A(n27216), .B(n27217), .Z(n26911) );
  XOR U28451 ( .A(n27214), .B(n27228), .Z(n27217) );
  NAND U28452 ( .A(b[1]), .B(a[52]), .Z(n27228) );
  XOR U28453 ( .A(n27222), .B(n27229), .Z(n27216) );
  XOR U28454 ( .A(n27214), .B(n27221), .Z(n27229) );
  XNOR U28455 ( .A(n27230), .B(n27220), .Z(n27221) );
  AND U28456 ( .A(b[2]), .B(a[51]), .Z(n27230) );
  NANDN U28457 ( .A(n27231), .B(n27232), .Z(n27214) );
  XOR U28458 ( .A(n27220), .B(n27212), .Z(n27233) );
  XNOR U28459 ( .A(n27211), .B(n27207), .Z(n27234) );
  XNOR U28460 ( .A(n27206), .B(n27202), .Z(n27235) );
  XNOR U28461 ( .A(n27201), .B(n27197), .Z(n27236) );
  XNOR U28462 ( .A(n27196), .B(n27192), .Z(n27237) );
  XNOR U28463 ( .A(n27191), .B(n27187), .Z(n27238) );
  XNOR U28464 ( .A(n27186), .B(n27182), .Z(n27239) );
  XNOR U28465 ( .A(n27181), .B(n27177), .Z(n27240) );
  XNOR U28466 ( .A(n27176), .B(n27172), .Z(n27241) );
  XNOR U28467 ( .A(n27171), .B(n27167), .Z(n27242) );
  XNOR U28468 ( .A(n27166), .B(n27162), .Z(n27243) );
  XNOR U28469 ( .A(n27161), .B(n27157), .Z(n27244) );
  XNOR U28470 ( .A(n27156), .B(n27152), .Z(n27245) );
  XNOR U28471 ( .A(n27151), .B(n27147), .Z(n27246) );
  XNOR U28472 ( .A(n27146), .B(n27142), .Z(n27247) );
  XNOR U28473 ( .A(n27141), .B(n27137), .Z(n27248) );
  XNOR U28474 ( .A(n27136), .B(n27132), .Z(n27249) );
  XNOR U28475 ( .A(n27131), .B(n27127), .Z(n27250) );
  XNOR U28476 ( .A(n27126), .B(n27122), .Z(n27251) );
  XNOR U28477 ( .A(n27121), .B(n27117), .Z(n27252) );
  XNOR U28478 ( .A(n27116), .B(n27112), .Z(n27253) );
  XNOR U28479 ( .A(n27111), .B(n27107), .Z(n27254) );
  XNOR U28480 ( .A(n27106), .B(n27102), .Z(n27255) );
  XNOR U28481 ( .A(n27101), .B(n27097), .Z(n27256) );
  XNOR U28482 ( .A(n27096), .B(n27092), .Z(n27257) );
  XNOR U28483 ( .A(n27091), .B(n27087), .Z(n27258) );
  XNOR U28484 ( .A(n27086), .B(n27082), .Z(n27259) );
  XNOR U28485 ( .A(n27081), .B(n27077), .Z(n27260) );
  XNOR U28486 ( .A(n27076), .B(n27072), .Z(n27261) );
  XNOR U28487 ( .A(n27071), .B(n27067), .Z(n27262) );
  XNOR U28488 ( .A(n27066), .B(n27062), .Z(n27263) );
  XNOR U28489 ( .A(n27061), .B(n27057), .Z(n27264) );
  XNOR U28490 ( .A(n27056), .B(n27052), .Z(n27265) );
  XNOR U28491 ( .A(n27051), .B(n27047), .Z(n27266) );
  XNOR U28492 ( .A(n27046), .B(n27042), .Z(n27267) );
  XNOR U28493 ( .A(n27041), .B(n27037), .Z(n27268) );
  XNOR U28494 ( .A(n27036), .B(n27032), .Z(n27269) );
  XNOR U28495 ( .A(n27031), .B(n27027), .Z(n27270) );
  XNOR U28496 ( .A(n27026), .B(n27022), .Z(n27271) );
  XNOR U28497 ( .A(n27021), .B(n27017), .Z(n27272) );
  XNOR U28498 ( .A(n27016), .B(n27012), .Z(n27273) );
  XNOR U28499 ( .A(n27011), .B(n27007), .Z(n27274) );
  XNOR U28500 ( .A(n27006), .B(n27002), .Z(n27275) );
  XNOR U28501 ( .A(n27001), .B(n26997), .Z(n27276) );
  XNOR U28502 ( .A(n26996), .B(n26992), .Z(n27277) );
  XNOR U28503 ( .A(n26991), .B(n26987), .Z(n27278) );
  XNOR U28504 ( .A(n26986), .B(n26982), .Z(n27279) );
  XNOR U28505 ( .A(n26981), .B(n26977), .Z(n27280) );
  XNOR U28506 ( .A(n26976), .B(n26972), .Z(n27281) );
  XNOR U28507 ( .A(n26971), .B(n26967), .Z(n27282) );
  XOR U28508 ( .A(n27283), .B(n26966), .Z(n26967) );
  AND U28509 ( .A(a[0]), .B(b[53]), .Z(n27283) );
  XOR U28510 ( .A(n27284), .B(n26966), .Z(n26968) );
  XNOR U28511 ( .A(n27285), .B(n27286), .Z(n26966) );
  AND U28512 ( .A(n27287), .B(n27288), .Z(n27285) );
  AND U28513 ( .A(a[1]), .B(b[52]), .Z(n27284) );
  XOR U28514 ( .A(n27289), .B(n26971), .Z(n26973) );
  XOR U28515 ( .A(n27290), .B(n27291), .Z(n26971) );
  AND U28516 ( .A(n27292), .B(n27293), .Z(n27290) );
  AND U28517 ( .A(a[2]), .B(b[51]), .Z(n27289) );
  XOR U28518 ( .A(n27294), .B(n26976), .Z(n26978) );
  XOR U28519 ( .A(n27295), .B(n27296), .Z(n26976) );
  AND U28520 ( .A(n27297), .B(n27298), .Z(n27295) );
  AND U28521 ( .A(a[3]), .B(b[50]), .Z(n27294) );
  XOR U28522 ( .A(n27299), .B(n26981), .Z(n26983) );
  XOR U28523 ( .A(n27300), .B(n27301), .Z(n26981) );
  AND U28524 ( .A(n27302), .B(n27303), .Z(n27300) );
  AND U28525 ( .A(a[4]), .B(b[49]), .Z(n27299) );
  XOR U28526 ( .A(n27304), .B(n26986), .Z(n26988) );
  XOR U28527 ( .A(n27305), .B(n27306), .Z(n26986) );
  AND U28528 ( .A(n27307), .B(n27308), .Z(n27305) );
  AND U28529 ( .A(a[5]), .B(b[48]), .Z(n27304) );
  XOR U28530 ( .A(n27309), .B(n26991), .Z(n26993) );
  XOR U28531 ( .A(n27310), .B(n27311), .Z(n26991) );
  AND U28532 ( .A(n27312), .B(n27313), .Z(n27310) );
  AND U28533 ( .A(a[6]), .B(b[47]), .Z(n27309) );
  XOR U28534 ( .A(n27314), .B(n26996), .Z(n26998) );
  XOR U28535 ( .A(n27315), .B(n27316), .Z(n26996) );
  AND U28536 ( .A(n27317), .B(n27318), .Z(n27315) );
  AND U28537 ( .A(a[7]), .B(b[46]), .Z(n27314) );
  XOR U28538 ( .A(n27319), .B(n27001), .Z(n27003) );
  XOR U28539 ( .A(n27320), .B(n27321), .Z(n27001) );
  AND U28540 ( .A(n27322), .B(n27323), .Z(n27320) );
  AND U28541 ( .A(a[8]), .B(b[45]), .Z(n27319) );
  XOR U28542 ( .A(n27324), .B(n27006), .Z(n27008) );
  XOR U28543 ( .A(n27325), .B(n27326), .Z(n27006) );
  AND U28544 ( .A(n27327), .B(n27328), .Z(n27325) );
  AND U28545 ( .A(a[9]), .B(b[44]), .Z(n27324) );
  XOR U28546 ( .A(n27329), .B(n27011), .Z(n27013) );
  XOR U28547 ( .A(n27330), .B(n27331), .Z(n27011) );
  AND U28548 ( .A(n27332), .B(n27333), .Z(n27330) );
  AND U28549 ( .A(a[10]), .B(b[43]), .Z(n27329) );
  XOR U28550 ( .A(n27334), .B(n27016), .Z(n27018) );
  XOR U28551 ( .A(n27335), .B(n27336), .Z(n27016) );
  AND U28552 ( .A(n27337), .B(n27338), .Z(n27335) );
  AND U28553 ( .A(a[11]), .B(b[42]), .Z(n27334) );
  XOR U28554 ( .A(n27339), .B(n27021), .Z(n27023) );
  XOR U28555 ( .A(n27340), .B(n27341), .Z(n27021) );
  AND U28556 ( .A(n27342), .B(n27343), .Z(n27340) );
  AND U28557 ( .A(a[12]), .B(b[41]), .Z(n27339) );
  XOR U28558 ( .A(n27344), .B(n27026), .Z(n27028) );
  XOR U28559 ( .A(n27345), .B(n27346), .Z(n27026) );
  AND U28560 ( .A(n27347), .B(n27348), .Z(n27345) );
  AND U28561 ( .A(a[13]), .B(b[40]), .Z(n27344) );
  XOR U28562 ( .A(n27349), .B(n27031), .Z(n27033) );
  XOR U28563 ( .A(n27350), .B(n27351), .Z(n27031) );
  AND U28564 ( .A(n27352), .B(n27353), .Z(n27350) );
  AND U28565 ( .A(a[14]), .B(b[39]), .Z(n27349) );
  XOR U28566 ( .A(n27354), .B(n27036), .Z(n27038) );
  XOR U28567 ( .A(n27355), .B(n27356), .Z(n27036) );
  AND U28568 ( .A(n27357), .B(n27358), .Z(n27355) );
  AND U28569 ( .A(a[15]), .B(b[38]), .Z(n27354) );
  XOR U28570 ( .A(n27359), .B(n27041), .Z(n27043) );
  XOR U28571 ( .A(n27360), .B(n27361), .Z(n27041) );
  AND U28572 ( .A(n27362), .B(n27363), .Z(n27360) );
  AND U28573 ( .A(a[16]), .B(b[37]), .Z(n27359) );
  XOR U28574 ( .A(n27364), .B(n27046), .Z(n27048) );
  XOR U28575 ( .A(n27365), .B(n27366), .Z(n27046) );
  AND U28576 ( .A(n27367), .B(n27368), .Z(n27365) );
  AND U28577 ( .A(a[17]), .B(b[36]), .Z(n27364) );
  XOR U28578 ( .A(n27369), .B(n27051), .Z(n27053) );
  XOR U28579 ( .A(n27370), .B(n27371), .Z(n27051) );
  AND U28580 ( .A(n27372), .B(n27373), .Z(n27370) );
  AND U28581 ( .A(a[18]), .B(b[35]), .Z(n27369) );
  XOR U28582 ( .A(n27374), .B(n27056), .Z(n27058) );
  XOR U28583 ( .A(n27375), .B(n27376), .Z(n27056) );
  AND U28584 ( .A(n27377), .B(n27378), .Z(n27375) );
  AND U28585 ( .A(a[19]), .B(b[34]), .Z(n27374) );
  XOR U28586 ( .A(n27379), .B(n27061), .Z(n27063) );
  XOR U28587 ( .A(n27380), .B(n27381), .Z(n27061) );
  AND U28588 ( .A(n27382), .B(n27383), .Z(n27380) );
  AND U28589 ( .A(a[20]), .B(b[33]), .Z(n27379) );
  XOR U28590 ( .A(n27384), .B(n27066), .Z(n27068) );
  XOR U28591 ( .A(n27385), .B(n27386), .Z(n27066) );
  AND U28592 ( .A(n27387), .B(n27388), .Z(n27385) );
  AND U28593 ( .A(a[21]), .B(b[32]), .Z(n27384) );
  XOR U28594 ( .A(n27389), .B(n27071), .Z(n27073) );
  XOR U28595 ( .A(n27390), .B(n27391), .Z(n27071) );
  AND U28596 ( .A(n27392), .B(n27393), .Z(n27390) );
  AND U28597 ( .A(a[22]), .B(b[31]), .Z(n27389) );
  XOR U28598 ( .A(n27394), .B(n27076), .Z(n27078) );
  XOR U28599 ( .A(n27395), .B(n27396), .Z(n27076) );
  AND U28600 ( .A(n27397), .B(n27398), .Z(n27395) );
  AND U28601 ( .A(a[23]), .B(b[30]), .Z(n27394) );
  XOR U28602 ( .A(n27399), .B(n27081), .Z(n27083) );
  XOR U28603 ( .A(n27400), .B(n27401), .Z(n27081) );
  AND U28604 ( .A(n27402), .B(n27403), .Z(n27400) );
  AND U28605 ( .A(a[24]), .B(b[29]), .Z(n27399) );
  XOR U28606 ( .A(n27404), .B(n27086), .Z(n27088) );
  XOR U28607 ( .A(n27405), .B(n27406), .Z(n27086) );
  AND U28608 ( .A(n27407), .B(n27408), .Z(n27405) );
  AND U28609 ( .A(a[25]), .B(b[28]), .Z(n27404) );
  XOR U28610 ( .A(n27409), .B(n27091), .Z(n27093) );
  XOR U28611 ( .A(n27410), .B(n27411), .Z(n27091) );
  AND U28612 ( .A(n27412), .B(n27413), .Z(n27410) );
  AND U28613 ( .A(a[26]), .B(b[27]), .Z(n27409) );
  XOR U28614 ( .A(n27414), .B(n27096), .Z(n27098) );
  XOR U28615 ( .A(n27415), .B(n27416), .Z(n27096) );
  AND U28616 ( .A(n27417), .B(n27418), .Z(n27415) );
  AND U28617 ( .A(b[26]), .B(a[27]), .Z(n27414) );
  XOR U28618 ( .A(n27419), .B(n27101), .Z(n27103) );
  XOR U28619 ( .A(n27420), .B(n27421), .Z(n27101) );
  AND U28620 ( .A(n27422), .B(n27423), .Z(n27420) );
  AND U28621 ( .A(b[25]), .B(a[28]), .Z(n27419) );
  XOR U28622 ( .A(n27424), .B(n27106), .Z(n27108) );
  XOR U28623 ( .A(n27425), .B(n27426), .Z(n27106) );
  AND U28624 ( .A(n27427), .B(n27428), .Z(n27425) );
  AND U28625 ( .A(b[24]), .B(a[29]), .Z(n27424) );
  XOR U28626 ( .A(n27429), .B(n27111), .Z(n27113) );
  XOR U28627 ( .A(n27430), .B(n27431), .Z(n27111) );
  AND U28628 ( .A(n27432), .B(n27433), .Z(n27430) );
  AND U28629 ( .A(b[23]), .B(a[30]), .Z(n27429) );
  XOR U28630 ( .A(n27434), .B(n27116), .Z(n27118) );
  XOR U28631 ( .A(n27435), .B(n27436), .Z(n27116) );
  AND U28632 ( .A(n27437), .B(n27438), .Z(n27435) );
  AND U28633 ( .A(b[22]), .B(a[31]), .Z(n27434) );
  XOR U28634 ( .A(n27439), .B(n27121), .Z(n27123) );
  XOR U28635 ( .A(n27440), .B(n27441), .Z(n27121) );
  AND U28636 ( .A(n27442), .B(n27443), .Z(n27440) );
  AND U28637 ( .A(b[21]), .B(a[32]), .Z(n27439) );
  XOR U28638 ( .A(n27444), .B(n27126), .Z(n27128) );
  XOR U28639 ( .A(n27445), .B(n27446), .Z(n27126) );
  AND U28640 ( .A(n27447), .B(n27448), .Z(n27445) );
  AND U28641 ( .A(b[20]), .B(a[33]), .Z(n27444) );
  XOR U28642 ( .A(n27449), .B(n27131), .Z(n27133) );
  XOR U28643 ( .A(n27450), .B(n27451), .Z(n27131) );
  AND U28644 ( .A(n27452), .B(n27453), .Z(n27450) );
  AND U28645 ( .A(b[19]), .B(a[34]), .Z(n27449) );
  XOR U28646 ( .A(n27454), .B(n27136), .Z(n27138) );
  XOR U28647 ( .A(n27455), .B(n27456), .Z(n27136) );
  AND U28648 ( .A(n27457), .B(n27458), .Z(n27455) );
  AND U28649 ( .A(b[18]), .B(a[35]), .Z(n27454) );
  XOR U28650 ( .A(n27459), .B(n27141), .Z(n27143) );
  XOR U28651 ( .A(n27460), .B(n27461), .Z(n27141) );
  AND U28652 ( .A(n27462), .B(n27463), .Z(n27460) );
  AND U28653 ( .A(b[17]), .B(a[36]), .Z(n27459) );
  XOR U28654 ( .A(n27464), .B(n27146), .Z(n27148) );
  XOR U28655 ( .A(n27465), .B(n27466), .Z(n27146) );
  AND U28656 ( .A(n27467), .B(n27468), .Z(n27465) );
  AND U28657 ( .A(b[16]), .B(a[37]), .Z(n27464) );
  XOR U28658 ( .A(n27469), .B(n27151), .Z(n27153) );
  XOR U28659 ( .A(n27470), .B(n27471), .Z(n27151) );
  AND U28660 ( .A(n27472), .B(n27473), .Z(n27470) );
  AND U28661 ( .A(b[15]), .B(a[38]), .Z(n27469) );
  XOR U28662 ( .A(n27474), .B(n27156), .Z(n27158) );
  XOR U28663 ( .A(n27475), .B(n27476), .Z(n27156) );
  AND U28664 ( .A(n27477), .B(n27478), .Z(n27475) );
  AND U28665 ( .A(b[14]), .B(a[39]), .Z(n27474) );
  XOR U28666 ( .A(n27479), .B(n27161), .Z(n27163) );
  XOR U28667 ( .A(n27480), .B(n27481), .Z(n27161) );
  AND U28668 ( .A(n27482), .B(n27483), .Z(n27480) );
  AND U28669 ( .A(b[13]), .B(a[40]), .Z(n27479) );
  XOR U28670 ( .A(n27484), .B(n27166), .Z(n27168) );
  XOR U28671 ( .A(n27485), .B(n27486), .Z(n27166) );
  AND U28672 ( .A(n27487), .B(n27488), .Z(n27485) );
  AND U28673 ( .A(b[12]), .B(a[41]), .Z(n27484) );
  XOR U28674 ( .A(n27489), .B(n27171), .Z(n27173) );
  XOR U28675 ( .A(n27490), .B(n27491), .Z(n27171) );
  AND U28676 ( .A(n27492), .B(n27493), .Z(n27490) );
  AND U28677 ( .A(b[11]), .B(a[42]), .Z(n27489) );
  XOR U28678 ( .A(n27494), .B(n27176), .Z(n27178) );
  XOR U28679 ( .A(n27495), .B(n27496), .Z(n27176) );
  AND U28680 ( .A(n27497), .B(n27498), .Z(n27495) );
  AND U28681 ( .A(b[10]), .B(a[43]), .Z(n27494) );
  XOR U28682 ( .A(n27499), .B(n27181), .Z(n27183) );
  XOR U28683 ( .A(n27500), .B(n27501), .Z(n27181) );
  AND U28684 ( .A(n27502), .B(n27503), .Z(n27500) );
  AND U28685 ( .A(b[9]), .B(a[44]), .Z(n27499) );
  XOR U28686 ( .A(n27504), .B(n27186), .Z(n27188) );
  XOR U28687 ( .A(n27505), .B(n27506), .Z(n27186) );
  AND U28688 ( .A(n27507), .B(n27508), .Z(n27505) );
  AND U28689 ( .A(b[8]), .B(a[45]), .Z(n27504) );
  XOR U28690 ( .A(n27509), .B(n27191), .Z(n27193) );
  XOR U28691 ( .A(n27510), .B(n27511), .Z(n27191) );
  AND U28692 ( .A(n27512), .B(n27513), .Z(n27510) );
  AND U28693 ( .A(b[7]), .B(a[46]), .Z(n27509) );
  XOR U28694 ( .A(n27514), .B(n27196), .Z(n27198) );
  XOR U28695 ( .A(n27515), .B(n27516), .Z(n27196) );
  AND U28696 ( .A(n27517), .B(n27518), .Z(n27515) );
  AND U28697 ( .A(b[6]), .B(a[47]), .Z(n27514) );
  XOR U28698 ( .A(n27519), .B(n27201), .Z(n27203) );
  XOR U28699 ( .A(n27520), .B(n27521), .Z(n27201) );
  AND U28700 ( .A(n27522), .B(n27523), .Z(n27520) );
  AND U28701 ( .A(b[5]), .B(a[48]), .Z(n27519) );
  XOR U28702 ( .A(n27524), .B(n27206), .Z(n27208) );
  XOR U28703 ( .A(n27525), .B(n27526), .Z(n27206) );
  AND U28704 ( .A(n27527), .B(n27528), .Z(n27525) );
  AND U28705 ( .A(b[4]), .B(a[49]), .Z(n27524) );
  XNOR U28706 ( .A(n27529), .B(n27530), .Z(n27220) );
  NANDN U28707 ( .A(n27531), .B(n27532), .Z(n27530) );
  XOR U28708 ( .A(n27533), .B(n27211), .Z(n27213) );
  XNOR U28709 ( .A(n27534), .B(n27535), .Z(n27211) );
  AND U28710 ( .A(n27536), .B(n27537), .Z(n27534) );
  AND U28711 ( .A(b[3]), .B(a[50]), .Z(n27533) );
  XOR U28712 ( .A(n27227), .B(n27226), .Z(c[116]) );
  XOR U28713 ( .A(sreg[180]), .B(n27225), .Z(n27226) );
  XOR U28714 ( .A(n27232), .B(n27538), .Z(n27227) );
  XNOR U28715 ( .A(n27231), .B(n27225), .Z(n27538) );
  XOR U28716 ( .A(n27539), .B(n27540), .Z(n27225) );
  NOR U28717 ( .A(n27541), .B(n27542), .Z(n27539) );
  NAND U28718 ( .A(a[52]), .B(b[0]), .Z(n27231) );
  XNOR U28719 ( .A(n27531), .B(n27532), .Z(n27232) );
  XOR U28720 ( .A(n27529), .B(n27543), .Z(n27532) );
  NAND U28721 ( .A(b[1]), .B(a[51]), .Z(n27543) );
  XOR U28722 ( .A(n27537), .B(n27544), .Z(n27531) );
  XOR U28723 ( .A(n27529), .B(n27536), .Z(n27544) );
  XNOR U28724 ( .A(n27545), .B(n27535), .Z(n27536) );
  AND U28725 ( .A(b[2]), .B(a[50]), .Z(n27545) );
  NANDN U28726 ( .A(n27546), .B(n27547), .Z(n27529) );
  XOR U28727 ( .A(n27535), .B(n27527), .Z(n27548) );
  XNOR U28728 ( .A(n27526), .B(n27522), .Z(n27549) );
  XNOR U28729 ( .A(n27521), .B(n27517), .Z(n27550) );
  XNOR U28730 ( .A(n27516), .B(n27512), .Z(n27551) );
  XNOR U28731 ( .A(n27511), .B(n27507), .Z(n27552) );
  XNOR U28732 ( .A(n27506), .B(n27502), .Z(n27553) );
  XNOR U28733 ( .A(n27501), .B(n27497), .Z(n27554) );
  XNOR U28734 ( .A(n27496), .B(n27492), .Z(n27555) );
  XNOR U28735 ( .A(n27491), .B(n27487), .Z(n27556) );
  XNOR U28736 ( .A(n27486), .B(n27482), .Z(n27557) );
  XNOR U28737 ( .A(n27481), .B(n27477), .Z(n27558) );
  XNOR U28738 ( .A(n27476), .B(n27472), .Z(n27559) );
  XNOR U28739 ( .A(n27471), .B(n27467), .Z(n27560) );
  XNOR U28740 ( .A(n27466), .B(n27462), .Z(n27561) );
  XNOR U28741 ( .A(n27461), .B(n27457), .Z(n27562) );
  XNOR U28742 ( .A(n27456), .B(n27452), .Z(n27563) );
  XNOR U28743 ( .A(n27451), .B(n27447), .Z(n27564) );
  XNOR U28744 ( .A(n27446), .B(n27442), .Z(n27565) );
  XNOR U28745 ( .A(n27441), .B(n27437), .Z(n27566) );
  XNOR U28746 ( .A(n27436), .B(n27432), .Z(n27567) );
  XNOR U28747 ( .A(n27431), .B(n27427), .Z(n27568) );
  XNOR U28748 ( .A(n27426), .B(n27422), .Z(n27569) );
  XNOR U28749 ( .A(n27421), .B(n27417), .Z(n27570) );
  XNOR U28750 ( .A(n27416), .B(n27412), .Z(n27571) );
  XNOR U28751 ( .A(n27411), .B(n27407), .Z(n27572) );
  XNOR U28752 ( .A(n27406), .B(n27402), .Z(n27573) );
  XNOR U28753 ( .A(n27401), .B(n27397), .Z(n27574) );
  XNOR U28754 ( .A(n27396), .B(n27392), .Z(n27575) );
  XNOR U28755 ( .A(n27391), .B(n27387), .Z(n27576) );
  XNOR U28756 ( .A(n27386), .B(n27382), .Z(n27577) );
  XNOR U28757 ( .A(n27381), .B(n27377), .Z(n27578) );
  XNOR U28758 ( .A(n27376), .B(n27372), .Z(n27579) );
  XNOR U28759 ( .A(n27371), .B(n27367), .Z(n27580) );
  XNOR U28760 ( .A(n27366), .B(n27362), .Z(n27581) );
  XNOR U28761 ( .A(n27361), .B(n27357), .Z(n27582) );
  XNOR U28762 ( .A(n27356), .B(n27352), .Z(n27583) );
  XNOR U28763 ( .A(n27351), .B(n27347), .Z(n27584) );
  XNOR U28764 ( .A(n27346), .B(n27342), .Z(n27585) );
  XNOR U28765 ( .A(n27341), .B(n27337), .Z(n27586) );
  XNOR U28766 ( .A(n27336), .B(n27332), .Z(n27587) );
  XNOR U28767 ( .A(n27331), .B(n27327), .Z(n27588) );
  XNOR U28768 ( .A(n27326), .B(n27322), .Z(n27589) );
  XNOR U28769 ( .A(n27321), .B(n27317), .Z(n27590) );
  XNOR U28770 ( .A(n27316), .B(n27312), .Z(n27591) );
  XNOR U28771 ( .A(n27311), .B(n27307), .Z(n27592) );
  XNOR U28772 ( .A(n27306), .B(n27302), .Z(n27593) );
  XNOR U28773 ( .A(n27301), .B(n27297), .Z(n27594) );
  XNOR U28774 ( .A(n27296), .B(n27292), .Z(n27595) );
  XNOR U28775 ( .A(n27291), .B(n27287), .Z(n27596) );
  XNOR U28776 ( .A(n27597), .B(n27286), .Z(n27287) );
  AND U28777 ( .A(a[0]), .B(b[52]), .Z(n27597) );
  XNOR U28778 ( .A(n27598), .B(n27286), .Z(n27288) );
  XNOR U28779 ( .A(n27599), .B(n27600), .Z(n27286) );
  AND U28780 ( .A(n27601), .B(n27602), .Z(n27599) );
  AND U28781 ( .A(a[1]), .B(b[51]), .Z(n27598) );
  XOR U28782 ( .A(n27603), .B(n27291), .Z(n27293) );
  XOR U28783 ( .A(n27604), .B(n27605), .Z(n27291) );
  AND U28784 ( .A(n27606), .B(n27607), .Z(n27604) );
  AND U28785 ( .A(a[2]), .B(b[50]), .Z(n27603) );
  XOR U28786 ( .A(n27608), .B(n27296), .Z(n27298) );
  XOR U28787 ( .A(n27609), .B(n27610), .Z(n27296) );
  AND U28788 ( .A(n27611), .B(n27612), .Z(n27609) );
  AND U28789 ( .A(a[3]), .B(b[49]), .Z(n27608) );
  XOR U28790 ( .A(n27613), .B(n27301), .Z(n27303) );
  XOR U28791 ( .A(n27614), .B(n27615), .Z(n27301) );
  AND U28792 ( .A(n27616), .B(n27617), .Z(n27614) );
  AND U28793 ( .A(a[4]), .B(b[48]), .Z(n27613) );
  XOR U28794 ( .A(n27618), .B(n27306), .Z(n27308) );
  XOR U28795 ( .A(n27619), .B(n27620), .Z(n27306) );
  AND U28796 ( .A(n27621), .B(n27622), .Z(n27619) );
  AND U28797 ( .A(a[5]), .B(b[47]), .Z(n27618) );
  XOR U28798 ( .A(n27623), .B(n27311), .Z(n27313) );
  XOR U28799 ( .A(n27624), .B(n27625), .Z(n27311) );
  AND U28800 ( .A(n27626), .B(n27627), .Z(n27624) );
  AND U28801 ( .A(a[6]), .B(b[46]), .Z(n27623) );
  XOR U28802 ( .A(n27628), .B(n27316), .Z(n27318) );
  XOR U28803 ( .A(n27629), .B(n27630), .Z(n27316) );
  AND U28804 ( .A(n27631), .B(n27632), .Z(n27629) );
  AND U28805 ( .A(a[7]), .B(b[45]), .Z(n27628) );
  XOR U28806 ( .A(n27633), .B(n27321), .Z(n27323) );
  XOR U28807 ( .A(n27634), .B(n27635), .Z(n27321) );
  AND U28808 ( .A(n27636), .B(n27637), .Z(n27634) );
  AND U28809 ( .A(a[8]), .B(b[44]), .Z(n27633) );
  XOR U28810 ( .A(n27638), .B(n27326), .Z(n27328) );
  XOR U28811 ( .A(n27639), .B(n27640), .Z(n27326) );
  AND U28812 ( .A(n27641), .B(n27642), .Z(n27639) );
  AND U28813 ( .A(a[9]), .B(b[43]), .Z(n27638) );
  XOR U28814 ( .A(n27643), .B(n27331), .Z(n27333) );
  XOR U28815 ( .A(n27644), .B(n27645), .Z(n27331) );
  AND U28816 ( .A(n27646), .B(n27647), .Z(n27644) );
  AND U28817 ( .A(a[10]), .B(b[42]), .Z(n27643) );
  XOR U28818 ( .A(n27648), .B(n27336), .Z(n27338) );
  XOR U28819 ( .A(n27649), .B(n27650), .Z(n27336) );
  AND U28820 ( .A(n27651), .B(n27652), .Z(n27649) );
  AND U28821 ( .A(a[11]), .B(b[41]), .Z(n27648) );
  XOR U28822 ( .A(n27653), .B(n27341), .Z(n27343) );
  XOR U28823 ( .A(n27654), .B(n27655), .Z(n27341) );
  AND U28824 ( .A(n27656), .B(n27657), .Z(n27654) );
  AND U28825 ( .A(a[12]), .B(b[40]), .Z(n27653) );
  XOR U28826 ( .A(n27658), .B(n27346), .Z(n27348) );
  XOR U28827 ( .A(n27659), .B(n27660), .Z(n27346) );
  AND U28828 ( .A(n27661), .B(n27662), .Z(n27659) );
  AND U28829 ( .A(a[13]), .B(b[39]), .Z(n27658) );
  XOR U28830 ( .A(n27663), .B(n27351), .Z(n27353) );
  XOR U28831 ( .A(n27664), .B(n27665), .Z(n27351) );
  AND U28832 ( .A(n27666), .B(n27667), .Z(n27664) );
  AND U28833 ( .A(a[14]), .B(b[38]), .Z(n27663) );
  XOR U28834 ( .A(n27668), .B(n27356), .Z(n27358) );
  XOR U28835 ( .A(n27669), .B(n27670), .Z(n27356) );
  AND U28836 ( .A(n27671), .B(n27672), .Z(n27669) );
  AND U28837 ( .A(a[15]), .B(b[37]), .Z(n27668) );
  XOR U28838 ( .A(n27673), .B(n27361), .Z(n27363) );
  XOR U28839 ( .A(n27674), .B(n27675), .Z(n27361) );
  AND U28840 ( .A(n27676), .B(n27677), .Z(n27674) );
  AND U28841 ( .A(a[16]), .B(b[36]), .Z(n27673) );
  XOR U28842 ( .A(n27678), .B(n27366), .Z(n27368) );
  XOR U28843 ( .A(n27679), .B(n27680), .Z(n27366) );
  AND U28844 ( .A(n27681), .B(n27682), .Z(n27679) );
  AND U28845 ( .A(a[17]), .B(b[35]), .Z(n27678) );
  XOR U28846 ( .A(n27683), .B(n27371), .Z(n27373) );
  XOR U28847 ( .A(n27684), .B(n27685), .Z(n27371) );
  AND U28848 ( .A(n27686), .B(n27687), .Z(n27684) );
  AND U28849 ( .A(a[18]), .B(b[34]), .Z(n27683) );
  XOR U28850 ( .A(n27688), .B(n27376), .Z(n27378) );
  XOR U28851 ( .A(n27689), .B(n27690), .Z(n27376) );
  AND U28852 ( .A(n27691), .B(n27692), .Z(n27689) );
  AND U28853 ( .A(a[19]), .B(b[33]), .Z(n27688) );
  XOR U28854 ( .A(n27693), .B(n27381), .Z(n27383) );
  XOR U28855 ( .A(n27694), .B(n27695), .Z(n27381) );
  AND U28856 ( .A(n27696), .B(n27697), .Z(n27694) );
  AND U28857 ( .A(a[20]), .B(b[32]), .Z(n27693) );
  XOR U28858 ( .A(n27698), .B(n27386), .Z(n27388) );
  XOR U28859 ( .A(n27699), .B(n27700), .Z(n27386) );
  AND U28860 ( .A(n27701), .B(n27702), .Z(n27699) );
  AND U28861 ( .A(a[21]), .B(b[31]), .Z(n27698) );
  XOR U28862 ( .A(n27703), .B(n27391), .Z(n27393) );
  XOR U28863 ( .A(n27704), .B(n27705), .Z(n27391) );
  AND U28864 ( .A(n27706), .B(n27707), .Z(n27704) );
  AND U28865 ( .A(a[22]), .B(b[30]), .Z(n27703) );
  XOR U28866 ( .A(n27708), .B(n27396), .Z(n27398) );
  XOR U28867 ( .A(n27709), .B(n27710), .Z(n27396) );
  AND U28868 ( .A(n27711), .B(n27712), .Z(n27709) );
  AND U28869 ( .A(a[23]), .B(b[29]), .Z(n27708) );
  XOR U28870 ( .A(n27713), .B(n27401), .Z(n27403) );
  XOR U28871 ( .A(n27714), .B(n27715), .Z(n27401) );
  AND U28872 ( .A(n27716), .B(n27717), .Z(n27714) );
  AND U28873 ( .A(a[24]), .B(b[28]), .Z(n27713) );
  XOR U28874 ( .A(n27718), .B(n27406), .Z(n27408) );
  XOR U28875 ( .A(n27719), .B(n27720), .Z(n27406) );
  AND U28876 ( .A(n27721), .B(n27722), .Z(n27719) );
  AND U28877 ( .A(a[25]), .B(b[27]), .Z(n27718) );
  XOR U28878 ( .A(n27723), .B(n27411), .Z(n27413) );
  XOR U28879 ( .A(n27724), .B(n27725), .Z(n27411) );
  AND U28880 ( .A(n27726), .B(n27727), .Z(n27724) );
  AND U28881 ( .A(a[26]), .B(b[26]), .Z(n27723) );
  XOR U28882 ( .A(n27728), .B(n27416), .Z(n27418) );
  XOR U28883 ( .A(n27729), .B(n27730), .Z(n27416) );
  AND U28884 ( .A(n27731), .B(n27732), .Z(n27729) );
  AND U28885 ( .A(b[25]), .B(a[27]), .Z(n27728) );
  XOR U28886 ( .A(n27733), .B(n27421), .Z(n27423) );
  XOR U28887 ( .A(n27734), .B(n27735), .Z(n27421) );
  AND U28888 ( .A(n27736), .B(n27737), .Z(n27734) );
  AND U28889 ( .A(b[24]), .B(a[28]), .Z(n27733) );
  XOR U28890 ( .A(n27738), .B(n27426), .Z(n27428) );
  XOR U28891 ( .A(n27739), .B(n27740), .Z(n27426) );
  AND U28892 ( .A(n27741), .B(n27742), .Z(n27739) );
  AND U28893 ( .A(b[23]), .B(a[29]), .Z(n27738) );
  XOR U28894 ( .A(n27743), .B(n27431), .Z(n27433) );
  XOR U28895 ( .A(n27744), .B(n27745), .Z(n27431) );
  AND U28896 ( .A(n27746), .B(n27747), .Z(n27744) );
  AND U28897 ( .A(b[22]), .B(a[30]), .Z(n27743) );
  XOR U28898 ( .A(n27748), .B(n27436), .Z(n27438) );
  XOR U28899 ( .A(n27749), .B(n27750), .Z(n27436) );
  AND U28900 ( .A(n27751), .B(n27752), .Z(n27749) );
  AND U28901 ( .A(b[21]), .B(a[31]), .Z(n27748) );
  XOR U28902 ( .A(n27753), .B(n27441), .Z(n27443) );
  XOR U28903 ( .A(n27754), .B(n27755), .Z(n27441) );
  AND U28904 ( .A(n27756), .B(n27757), .Z(n27754) );
  AND U28905 ( .A(b[20]), .B(a[32]), .Z(n27753) );
  XOR U28906 ( .A(n27758), .B(n27446), .Z(n27448) );
  XOR U28907 ( .A(n27759), .B(n27760), .Z(n27446) );
  AND U28908 ( .A(n27761), .B(n27762), .Z(n27759) );
  AND U28909 ( .A(b[19]), .B(a[33]), .Z(n27758) );
  XOR U28910 ( .A(n27763), .B(n27451), .Z(n27453) );
  XOR U28911 ( .A(n27764), .B(n27765), .Z(n27451) );
  AND U28912 ( .A(n27766), .B(n27767), .Z(n27764) );
  AND U28913 ( .A(b[18]), .B(a[34]), .Z(n27763) );
  XOR U28914 ( .A(n27768), .B(n27456), .Z(n27458) );
  XOR U28915 ( .A(n27769), .B(n27770), .Z(n27456) );
  AND U28916 ( .A(n27771), .B(n27772), .Z(n27769) );
  AND U28917 ( .A(b[17]), .B(a[35]), .Z(n27768) );
  XOR U28918 ( .A(n27773), .B(n27461), .Z(n27463) );
  XOR U28919 ( .A(n27774), .B(n27775), .Z(n27461) );
  AND U28920 ( .A(n27776), .B(n27777), .Z(n27774) );
  AND U28921 ( .A(b[16]), .B(a[36]), .Z(n27773) );
  XOR U28922 ( .A(n27778), .B(n27466), .Z(n27468) );
  XOR U28923 ( .A(n27779), .B(n27780), .Z(n27466) );
  AND U28924 ( .A(n27781), .B(n27782), .Z(n27779) );
  AND U28925 ( .A(b[15]), .B(a[37]), .Z(n27778) );
  XOR U28926 ( .A(n27783), .B(n27471), .Z(n27473) );
  XOR U28927 ( .A(n27784), .B(n27785), .Z(n27471) );
  AND U28928 ( .A(n27786), .B(n27787), .Z(n27784) );
  AND U28929 ( .A(b[14]), .B(a[38]), .Z(n27783) );
  XOR U28930 ( .A(n27788), .B(n27476), .Z(n27478) );
  XOR U28931 ( .A(n27789), .B(n27790), .Z(n27476) );
  AND U28932 ( .A(n27791), .B(n27792), .Z(n27789) );
  AND U28933 ( .A(b[13]), .B(a[39]), .Z(n27788) );
  XOR U28934 ( .A(n27793), .B(n27481), .Z(n27483) );
  XOR U28935 ( .A(n27794), .B(n27795), .Z(n27481) );
  AND U28936 ( .A(n27796), .B(n27797), .Z(n27794) );
  AND U28937 ( .A(b[12]), .B(a[40]), .Z(n27793) );
  XOR U28938 ( .A(n27798), .B(n27486), .Z(n27488) );
  XOR U28939 ( .A(n27799), .B(n27800), .Z(n27486) );
  AND U28940 ( .A(n27801), .B(n27802), .Z(n27799) );
  AND U28941 ( .A(b[11]), .B(a[41]), .Z(n27798) );
  XOR U28942 ( .A(n27803), .B(n27491), .Z(n27493) );
  XOR U28943 ( .A(n27804), .B(n27805), .Z(n27491) );
  AND U28944 ( .A(n27806), .B(n27807), .Z(n27804) );
  AND U28945 ( .A(b[10]), .B(a[42]), .Z(n27803) );
  XOR U28946 ( .A(n27808), .B(n27496), .Z(n27498) );
  XOR U28947 ( .A(n27809), .B(n27810), .Z(n27496) );
  AND U28948 ( .A(n27811), .B(n27812), .Z(n27809) );
  AND U28949 ( .A(b[9]), .B(a[43]), .Z(n27808) );
  XOR U28950 ( .A(n27813), .B(n27501), .Z(n27503) );
  XOR U28951 ( .A(n27814), .B(n27815), .Z(n27501) );
  AND U28952 ( .A(n27816), .B(n27817), .Z(n27814) );
  AND U28953 ( .A(b[8]), .B(a[44]), .Z(n27813) );
  XOR U28954 ( .A(n27818), .B(n27506), .Z(n27508) );
  XOR U28955 ( .A(n27819), .B(n27820), .Z(n27506) );
  AND U28956 ( .A(n27821), .B(n27822), .Z(n27819) );
  AND U28957 ( .A(b[7]), .B(a[45]), .Z(n27818) );
  XOR U28958 ( .A(n27823), .B(n27511), .Z(n27513) );
  XOR U28959 ( .A(n27824), .B(n27825), .Z(n27511) );
  AND U28960 ( .A(n27826), .B(n27827), .Z(n27824) );
  AND U28961 ( .A(b[6]), .B(a[46]), .Z(n27823) );
  XOR U28962 ( .A(n27828), .B(n27516), .Z(n27518) );
  XOR U28963 ( .A(n27829), .B(n27830), .Z(n27516) );
  AND U28964 ( .A(n27831), .B(n27832), .Z(n27829) );
  AND U28965 ( .A(b[5]), .B(a[47]), .Z(n27828) );
  XOR U28966 ( .A(n27833), .B(n27521), .Z(n27523) );
  XOR U28967 ( .A(n27834), .B(n27835), .Z(n27521) );
  AND U28968 ( .A(n27836), .B(n27837), .Z(n27834) );
  AND U28969 ( .A(b[4]), .B(a[48]), .Z(n27833) );
  XNOR U28970 ( .A(n27838), .B(n27839), .Z(n27535) );
  NANDN U28971 ( .A(n27840), .B(n27841), .Z(n27839) );
  XOR U28972 ( .A(n27842), .B(n27526), .Z(n27528) );
  XNOR U28973 ( .A(n27843), .B(n27844), .Z(n27526) );
  AND U28974 ( .A(n27845), .B(n27846), .Z(n27843) );
  AND U28975 ( .A(b[3]), .B(a[49]), .Z(n27842) );
  XOR U28976 ( .A(n27542), .B(n27541), .Z(c[115]) );
  XOR U28977 ( .A(sreg[179]), .B(n27540), .Z(n27541) );
  XOR U28978 ( .A(n27547), .B(n27847), .Z(n27542) );
  XNOR U28979 ( .A(n27546), .B(n27540), .Z(n27847) );
  XOR U28980 ( .A(n27848), .B(n27849), .Z(n27540) );
  NOR U28981 ( .A(n27850), .B(n27851), .Z(n27848) );
  NAND U28982 ( .A(a[51]), .B(b[0]), .Z(n27546) );
  XNOR U28983 ( .A(n27840), .B(n27841), .Z(n27547) );
  XOR U28984 ( .A(n27838), .B(n27852), .Z(n27841) );
  NAND U28985 ( .A(b[1]), .B(a[50]), .Z(n27852) );
  XOR U28986 ( .A(n27846), .B(n27853), .Z(n27840) );
  XOR U28987 ( .A(n27838), .B(n27845), .Z(n27853) );
  XNOR U28988 ( .A(n27854), .B(n27844), .Z(n27845) );
  AND U28989 ( .A(b[2]), .B(a[49]), .Z(n27854) );
  NANDN U28990 ( .A(n27855), .B(n27856), .Z(n27838) );
  XOR U28991 ( .A(n27844), .B(n27836), .Z(n27857) );
  XNOR U28992 ( .A(n27835), .B(n27831), .Z(n27858) );
  XNOR U28993 ( .A(n27830), .B(n27826), .Z(n27859) );
  XNOR U28994 ( .A(n27825), .B(n27821), .Z(n27860) );
  XNOR U28995 ( .A(n27820), .B(n27816), .Z(n27861) );
  XNOR U28996 ( .A(n27815), .B(n27811), .Z(n27862) );
  XNOR U28997 ( .A(n27810), .B(n27806), .Z(n27863) );
  XNOR U28998 ( .A(n27805), .B(n27801), .Z(n27864) );
  XNOR U28999 ( .A(n27800), .B(n27796), .Z(n27865) );
  XNOR U29000 ( .A(n27795), .B(n27791), .Z(n27866) );
  XNOR U29001 ( .A(n27790), .B(n27786), .Z(n27867) );
  XNOR U29002 ( .A(n27785), .B(n27781), .Z(n27868) );
  XNOR U29003 ( .A(n27780), .B(n27776), .Z(n27869) );
  XNOR U29004 ( .A(n27775), .B(n27771), .Z(n27870) );
  XNOR U29005 ( .A(n27770), .B(n27766), .Z(n27871) );
  XNOR U29006 ( .A(n27765), .B(n27761), .Z(n27872) );
  XNOR U29007 ( .A(n27760), .B(n27756), .Z(n27873) );
  XNOR U29008 ( .A(n27755), .B(n27751), .Z(n27874) );
  XNOR U29009 ( .A(n27750), .B(n27746), .Z(n27875) );
  XNOR U29010 ( .A(n27745), .B(n27741), .Z(n27876) );
  XNOR U29011 ( .A(n27740), .B(n27736), .Z(n27877) );
  XNOR U29012 ( .A(n27735), .B(n27731), .Z(n27878) );
  XNOR U29013 ( .A(n27730), .B(n27726), .Z(n27879) );
  XNOR U29014 ( .A(n27725), .B(n27721), .Z(n27880) );
  XNOR U29015 ( .A(n27720), .B(n27716), .Z(n27881) );
  XNOR U29016 ( .A(n27715), .B(n27711), .Z(n27882) );
  XNOR U29017 ( .A(n27710), .B(n27706), .Z(n27883) );
  XNOR U29018 ( .A(n27705), .B(n27701), .Z(n27884) );
  XNOR U29019 ( .A(n27700), .B(n27696), .Z(n27885) );
  XNOR U29020 ( .A(n27695), .B(n27691), .Z(n27886) );
  XNOR U29021 ( .A(n27690), .B(n27686), .Z(n27887) );
  XNOR U29022 ( .A(n27685), .B(n27681), .Z(n27888) );
  XNOR U29023 ( .A(n27680), .B(n27676), .Z(n27889) );
  XNOR U29024 ( .A(n27675), .B(n27671), .Z(n27890) );
  XNOR U29025 ( .A(n27670), .B(n27666), .Z(n27891) );
  XNOR U29026 ( .A(n27665), .B(n27661), .Z(n27892) );
  XNOR U29027 ( .A(n27660), .B(n27656), .Z(n27893) );
  XNOR U29028 ( .A(n27655), .B(n27651), .Z(n27894) );
  XNOR U29029 ( .A(n27650), .B(n27646), .Z(n27895) );
  XNOR U29030 ( .A(n27645), .B(n27641), .Z(n27896) );
  XNOR U29031 ( .A(n27640), .B(n27636), .Z(n27897) );
  XNOR U29032 ( .A(n27635), .B(n27631), .Z(n27898) );
  XNOR U29033 ( .A(n27630), .B(n27626), .Z(n27899) );
  XNOR U29034 ( .A(n27625), .B(n27621), .Z(n27900) );
  XNOR U29035 ( .A(n27620), .B(n27616), .Z(n27901) );
  XNOR U29036 ( .A(n27615), .B(n27611), .Z(n27902) );
  XNOR U29037 ( .A(n27610), .B(n27606), .Z(n27903) );
  XNOR U29038 ( .A(n27605), .B(n27601), .Z(n27904) );
  XOR U29039 ( .A(n27905), .B(n27600), .Z(n27601) );
  AND U29040 ( .A(a[0]), .B(b[51]), .Z(n27905) );
  XOR U29041 ( .A(n27906), .B(n27600), .Z(n27602) );
  XNOR U29042 ( .A(n27907), .B(n27908), .Z(n27600) );
  AND U29043 ( .A(n27909), .B(n27910), .Z(n27907) );
  AND U29044 ( .A(a[1]), .B(b[50]), .Z(n27906) );
  XOR U29045 ( .A(n27911), .B(n27605), .Z(n27607) );
  XOR U29046 ( .A(n27912), .B(n27913), .Z(n27605) );
  AND U29047 ( .A(n27914), .B(n27915), .Z(n27912) );
  AND U29048 ( .A(a[2]), .B(b[49]), .Z(n27911) );
  XOR U29049 ( .A(n27916), .B(n27610), .Z(n27612) );
  XOR U29050 ( .A(n27917), .B(n27918), .Z(n27610) );
  AND U29051 ( .A(n27919), .B(n27920), .Z(n27917) );
  AND U29052 ( .A(a[3]), .B(b[48]), .Z(n27916) );
  XOR U29053 ( .A(n27921), .B(n27615), .Z(n27617) );
  XOR U29054 ( .A(n27922), .B(n27923), .Z(n27615) );
  AND U29055 ( .A(n27924), .B(n27925), .Z(n27922) );
  AND U29056 ( .A(a[4]), .B(b[47]), .Z(n27921) );
  XOR U29057 ( .A(n27926), .B(n27620), .Z(n27622) );
  XOR U29058 ( .A(n27927), .B(n27928), .Z(n27620) );
  AND U29059 ( .A(n27929), .B(n27930), .Z(n27927) );
  AND U29060 ( .A(a[5]), .B(b[46]), .Z(n27926) );
  XOR U29061 ( .A(n27931), .B(n27625), .Z(n27627) );
  XOR U29062 ( .A(n27932), .B(n27933), .Z(n27625) );
  AND U29063 ( .A(n27934), .B(n27935), .Z(n27932) );
  AND U29064 ( .A(a[6]), .B(b[45]), .Z(n27931) );
  XOR U29065 ( .A(n27936), .B(n27630), .Z(n27632) );
  XOR U29066 ( .A(n27937), .B(n27938), .Z(n27630) );
  AND U29067 ( .A(n27939), .B(n27940), .Z(n27937) );
  AND U29068 ( .A(a[7]), .B(b[44]), .Z(n27936) );
  XOR U29069 ( .A(n27941), .B(n27635), .Z(n27637) );
  XOR U29070 ( .A(n27942), .B(n27943), .Z(n27635) );
  AND U29071 ( .A(n27944), .B(n27945), .Z(n27942) );
  AND U29072 ( .A(a[8]), .B(b[43]), .Z(n27941) );
  XOR U29073 ( .A(n27946), .B(n27640), .Z(n27642) );
  XOR U29074 ( .A(n27947), .B(n27948), .Z(n27640) );
  AND U29075 ( .A(n27949), .B(n27950), .Z(n27947) );
  AND U29076 ( .A(a[9]), .B(b[42]), .Z(n27946) );
  XOR U29077 ( .A(n27951), .B(n27645), .Z(n27647) );
  XOR U29078 ( .A(n27952), .B(n27953), .Z(n27645) );
  AND U29079 ( .A(n27954), .B(n27955), .Z(n27952) );
  AND U29080 ( .A(a[10]), .B(b[41]), .Z(n27951) );
  XOR U29081 ( .A(n27956), .B(n27650), .Z(n27652) );
  XOR U29082 ( .A(n27957), .B(n27958), .Z(n27650) );
  AND U29083 ( .A(n27959), .B(n27960), .Z(n27957) );
  AND U29084 ( .A(a[11]), .B(b[40]), .Z(n27956) );
  XOR U29085 ( .A(n27961), .B(n27655), .Z(n27657) );
  XOR U29086 ( .A(n27962), .B(n27963), .Z(n27655) );
  AND U29087 ( .A(n27964), .B(n27965), .Z(n27962) );
  AND U29088 ( .A(a[12]), .B(b[39]), .Z(n27961) );
  XOR U29089 ( .A(n27966), .B(n27660), .Z(n27662) );
  XOR U29090 ( .A(n27967), .B(n27968), .Z(n27660) );
  AND U29091 ( .A(n27969), .B(n27970), .Z(n27967) );
  AND U29092 ( .A(a[13]), .B(b[38]), .Z(n27966) );
  XOR U29093 ( .A(n27971), .B(n27665), .Z(n27667) );
  XOR U29094 ( .A(n27972), .B(n27973), .Z(n27665) );
  AND U29095 ( .A(n27974), .B(n27975), .Z(n27972) );
  AND U29096 ( .A(a[14]), .B(b[37]), .Z(n27971) );
  XOR U29097 ( .A(n27976), .B(n27670), .Z(n27672) );
  XOR U29098 ( .A(n27977), .B(n27978), .Z(n27670) );
  AND U29099 ( .A(n27979), .B(n27980), .Z(n27977) );
  AND U29100 ( .A(a[15]), .B(b[36]), .Z(n27976) );
  XOR U29101 ( .A(n27981), .B(n27675), .Z(n27677) );
  XOR U29102 ( .A(n27982), .B(n27983), .Z(n27675) );
  AND U29103 ( .A(n27984), .B(n27985), .Z(n27982) );
  AND U29104 ( .A(a[16]), .B(b[35]), .Z(n27981) );
  XOR U29105 ( .A(n27986), .B(n27680), .Z(n27682) );
  XOR U29106 ( .A(n27987), .B(n27988), .Z(n27680) );
  AND U29107 ( .A(n27989), .B(n27990), .Z(n27987) );
  AND U29108 ( .A(a[17]), .B(b[34]), .Z(n27986) );
  XOR U29109 ( .A(n27991), .B(n27685), .Z(n27687) );
  XOR U29110 ( .A(n27992), .B(n27993), .Z(n27685) );
  AND U29111 ( .A(n27994), .B(n27995), .Z(n27992) );
  AND U29112 ( .A(a[18]), .B(b[33]), .Z(n27991) );
  XOR U29113 ( .A(n27996), .B(n27690), .Z(n27692) );
  XOR U29114 ( .A(n27997), .B(n27998), .Z(n27690) );
  AND U29115 ( .A(n27999), .B(n28000), .Z(n27997) );
  AND U29116 ( .A(a[19]), .B(b[32]), .Z(n27996) );
  XOR U29117 ( .A(n28001), .B(n27695), .Z(n27697) );
  XOR U29118 ( .A(n28002), .B(n28003), .Z(n27695) );
  AND U29119 ( .A(n28004), .B(n28005), .Z(n28002) );
  AND U29120 ( .A(a[20]), .B(b[31]), .Z(n28001) );
  XOR U29121 ( .A(n28006), .B(n27700), .Z(n27702) );
  XOR U29122 ( .A(n28007), .B(n28008), .Z(n27700) );
  AND U29123 ( .A(n28009), .B(n28010), .Z(n28007) );
  AND U29124 ( .A(a[21]), .B(b[30]), .Z(n28006) );
  XOR U29125 ( .A(n28011), .B(n27705), .Z(n27707) );
  XOR U29126 ( .A(n28012), .B(n28013), .Z(n27705) );
  AND U29127 ( .A(n28014), .B(n28015), .Z(n28012) );
  AND U29128 ( .A(a[22]), .B(b[29]), .Z(n28011) );
  XOR U29129 ( .A(n28016), .B(n27710), .Z(n27712) );
  XOR U29130 ( .A(n28017), .B(n28018), .Z(n27710) );
  AND U29131 ( .A(n28019), .B(n28020), .Z(n28017) );
  AND U29132 ( .A(a[23]), .B(b[28]), .Z(n28016) );
  XOR U29133 ( .A(n28021), .B(n27715), .Z(n27717) );
  XOR U29134 ( .A(n28022), .B(n28023), .Z(n27715) );
  AND U29135 ( .A(n28024), .B(n28025), .Z(n28022) );
  AND U29136 ( .A(a[24]), .B(b[27]), .Z(n28021) );
  XOR U29137 ( .A(n28026), .B(n27720), .Z(n27722) );
  XOR U29138 ( .A(n28027), .B(n28028), .Z(n27720) );
  AND U29139 ( .A(n28029), .B(n28030), .Z(n28027) );
  AND U29140 ( .A(a[25]), .B(b[26]), .Z(n28026) );
  XOR U29141 ( .A(n28031), .B(n27725), .Z(n27727) );
  XOR U29142 ( .A(n28032), .B(n28033), .Z(n27725) );
  AND U29143 ( .A(n28034), .B(n28035), .Z(n28032) );
  AND U29144 ( .A(b[25]), .B(a[26]), .Z(n28031) );
  XOR U29145 ( .A(n28036), .B(n27730), .Z(n27732) );
  XOR U29146 ( .A(n28037), .B(n28038), .Z(n27730) );
  AND U29147 ( .A(n28039), .B(n28040), .Z(n28037) );
  AND U29148 ( .A(b[24]), .B(a[27]), .Z(n28036) );
  XOR U29149 ( .A(n28041), .B(n27735), .Z(n27737) );
  XOR U29150 ( .A(n28042), .B(n28043), .Z(n27735) );
  AND U29151 ( .A(n28044), .B(n28045), .Z(n28042) );
  AND U29152 ( .A(b[23]), .B(a[28]), .Z(n28041) );
  XOR U29153 ( .A(n28046), .B(n27740), .Z(n27742) );
  XOR U29154 ( .A(n28047), .B(n28048), .Z(n27740) );
  AND U29155 ( .A(n28049), .B(n28050), .Z(n28047) );
  AND U29156 ( .A(b[22]), .B(a[29]), .Z(n28046) );
  XOR U29157 ( .A(n28051), .B(n27745), .Z(n27747) );
  XOR U29158 ( .A(n28052), .B(n28053), .Z(n27745) );
  AND U29159 ( .A(n28054), .B(n28055), .Z(n28052) );
  AND U29160 ( .A(b[21]), .B(a[30]), .Z(n28051) );
  XOR U29161 ( .A(n28056), .B(n27750), .Z(n27752) );
  XOR U29162 ( .A(n28057), .B(n28058), .Z(n27750) );
  AND U29163 ( .A(n28059), .B(n28060), .Z(n28057) );
  AND U29164 ( .A(b[20]), .B(a[31]), .Z(n28056) );
  XOR U29165 ( .A(n28061), .B(n27755), .Z(n27757) );
  XOR U29166 ( .A(n28062), .B(n28063), .Z(n27755) );
  AND U29167 ( .A(n28064), .B(n28065), .Z(n28062) );
  AND U29168 ( .A(b[19]), .B(a[32]), .Z(n28061) );
  XOR U29169 ( .A(n28066), .B(n27760), .Z(n27762) );
  XOR U29170 ( .A(n28067), .B(n28068), .Z(n27760) );
  AND U29171 ( .A(n28069), .B(n28070), .Z(n28067) );
  AND U29172 ( .A(b[18]), .B(a[33]), .Z(n28066) );
  XOR U29173 ( .A(n28071), .B(n27765), .Z(n27767) );
  XOR U29174 ( .A(n28072), .B(n28073), .Z(n27765) );
  AND U29175 ( .A(n28074), .B(n28075), .Z(n28072) );
  AND U29176 ( .A(b[17]), .B(a[34]), .Z(n28071) );
  XOR U29177 ( .A(n28076), .B(n27770), .Z(n27772) );
  XOR U29178 ( .A(n28077), .B(n28078), .Z(n27770) );
  AND U29179 ( .A(n28079), .B(n28080), .Z(n28077) );
  AND U29180 ( .A(b[16]), .B(a[35]), .Z(n28076) );
  XOR U29181 ( .A(n28081), .B(n27775), .Z(n27777) );
  XOR U29182 ( .A(n28082), .B(n28083), .Z(n27775) );
  AND U29183 ( .A(n28084), .B(n28085), .Z(n28082) );
  AND U29184 ( .A(b[15]), .B(a[36]), .Z(n28081) );
  XOR U29185 ( .A(n28086), .B(n27780), .Z(n27782) );
  XOR U29186 ( .A(n28087), .B(n28088), .Z(n27780) );
  AND U29187 ( .A(n28089), .B(n28090), .Z(n28087) );
  AND U29188 ( .A(b[14]), .B(a[37]), .Z(n28086) );
  XOR U29189 ( .A(n28091), .B(n27785), .Z(n27787) );
  XOR U29190 ( .A(n28092), .B(n28093), .Z(n27785) );
  AND U29191 ( .A(n28094), .B(n28095), .Z(n28092) );
  AND U29192 ( .A(b[13]), .B(a[38]), .Z(n28091) );
  XOR U29193 ( .A(n28096), .B(n27790), .Z(n27792) );
  XOR U29194 ( .A(n28097), .B(n28098), .Z(n27790) );
  AND U29195 ( .A(n28099), .B(n28100), .Z(n28097) );
  AND U29196 ( .A(b[12]), .B(a[39]), .Z(n28096) );
  XOR U29197 ( .A(n28101), .B(n27795), .Z(n27797) );
  XOR U29198 ( .A(n28102), .B(n28103), .Z(n27795) );
  AND U29199 ( .A(n28104), .B(n28105), .Z(n28102) );
  AND U29200 ( .A(b[11]), .B(a[40]), .Z(n28101) );
  XOR U29201 ( .A(n28106), .B(n27800), .Z(n27802) );
  XOR U29202 ( .A(n28107), .B(n28108), .Z(n27800) );
  AND U29203 ( .A(n28109), .B(n28110), .Z(n28107) );
  AND U29204 ( .A(b[10]), .B(a[41]), .Z(n28106) );
  XOR U29205 ( .A(n28111), .B(n27805), .Z(n27807) );
  XOR U29206 ( .A(n28112), .B(n28113), .Z(n27805) );
  AND U29207 ( .A(n28114), .B(n28115), .Z(n28112) );
  AND U29208 ( .A(b[9]), .B(a[42]), .Z(n28111) );
  XOR U29209 ( .A(n28116), .B(n27810), .Z(n27812) );
  XOR U29210 ( .A(n28117), .B(n28118), .Z(n27810) );
  AND U29211 ( .A(n28119), .B(n28120), .Z(n28117) );
  AND U29212 ( .A(b[8]), .B(a[43]), .Z(n28116) );
  XOR U29213 ( .A(n28121), .B(n27815), .Z(n27817) );
  XOR U29214 ( .A(n28122), .B(n28123), .Z(n27815) );
  AND U29215 ( .A(n28124), .B(n28125), .Z(n28122) );
  AND U29216 ( .A(b[7]), .B(a[44]), .Z(n28121) );
  XOR U29217 ( .A(n28126), .B(n27820), .Z(n27822) );
  XOR U29218 ( .A(n28127), .B(n28128), .Z(n27820) );
  AND U29219 ( .A(n28129), .B(n28130), .Z(n28127) );
  AND U29220 ( .A(b[6]), .B(a[45]), .Z(n28126) );
  XOR U29221 ( .A(n28131), .B(n27825), .Z(n27827) );
  XOR U29222 ( .A(n28132), .B(n28133), .Z(n27825) );
  AND U29223 ( .A(n28134), .B(n28135), .Z(n28132) );
  AND U29224 ( .A(b[5]), .B(a[46]), .Z(n28131) );
  XOR U29225 ( .A(n28136), .B(n27830), .Z(n27832) );
  XOR U29226 ( .A(n28137), .B(n28138), .Z(n27830) );
  AND U29227 ( .A(n28139), .B(n28140), .Z(n28137) );
  AND U29228 ( .A(b[4]), .B(a[47]), .Z(n28136) );
  XNOR U29229 ( .A(n28141), .B(n28142), .Z(n27844) );
  NANDN U29230 ( .A(n28143), .B(n28144), .Z(n28142) );
  XOR U29231 ( .A(n28145), .B(n27835), .Z(n27837) );
  XNOR U29232 ( .A(n28146), .B(n28147), .Z(n27835) );
  AND U29233 ( .A(n28148), .B(n28149), .Z(n28146) );
  AND U29234 ( .A(b[3]), .B(a[48]), .Z(n28145) );
  XOR U29235 ( .A(n27851), .B(n27850), .Z(c[114]) );
  XOR U29236 ( .A(sreg[178]), .B(n27849), .Z(n27850) );
  XOR U29237 ( .A(n27856), .B(n28150), .Z(n27851) );
  XNOR U29238 ( .A(n27855), .B(n27849), .Z(n28150) );
  XOR U29239 ( .A(n28151), .B(n28152), .Z(n27849) );
  NOR U29240 ( .A(n28153), .B(n28154), .Z(n28151) );
  NAND U29241 ( .A(a[50]), .B(b[0]), .Z(n27855) );
  XNOR U29242 ( .A(n28143), .B(n28144), .Z(n27856) );
  XOR U29243 ( .A(n28141), .B(n28155), .Z(n28144) );
  NAND U29244 ( .A(b[1]), .B(a[49]), .Z(n28155) );
  XOR U29245 ( .A(n28149), .B(n28156), .Z(n28143) );
  XOR U29246 ( .A(n28141), .B(n28148), .Z(n28156) );
  XNOR U29247 ( .A(n28157), .B(n28147), .Z(n28148) );
  AND U29248 ( .A(b[2]), .B(a[48]), .Z(n28157) );
  NANDN U29249 ( .A(n28158), .B(n28159), .Z(n28141) );
  XOR U29250 ( .A(n28147), .B(n28139), .Z(n28160) );
  XNOR U29251 ( .A(n28138), .B(n28134), .Z(n28161) );
  XNOR U29252 ( .A(n28133), .B(n28129), .Z(n28162) );
  XNOR U29253 ( .A(n28128), .B(n28124), .Z(n28163) );
  XNOR U29254 ( .A(n28123), .B(n28119), .Z(n28164) );
  XNOR U29255 ( .A(n28118), .B(n28114), .Z(n28165) );
  XNOR U29256 ( .A(n28113), .B(n28109), .Z(n28166) );
  XNOR U29257 ( .A(n28108), .B(n28104), .Z(n28167) );
  XNOR U29258 ( .A(n28103), .B(n28099), .Z(n28168) );
  XNOR U29259 ( .A(n28098), .B(n28094), .Z(n28169) );
  XNOR U29260 ( .A(n28093), .B(n28089), .Z(n28170) );
  XNOR U29261 ( .A(n28088), .B(n28084), .Z(n28171) );
  XNOR U29262 ( .A(n28083), .B(n28079), .Z(n28172) );
  XNOR U29263 ( .A(n28078), .B(n28074), .Z(n28173) );
  XNOR U29264 ( .A(n28073), .B(n28069), .Z(n28174) );
  XNOR U29265 ( .A(n28068), .B(n28064), .Z(n28175) );
  XNOR U29266 ( .A(n28063), .B(n28059), .Z(n28176) );
  XNOR U29267 ( .A(n28058), .B(n28054), .Z(n28177) );
  XNOR U29268 ( .A(n28053), .B(n28049), .Z(n28178) );
  XNOR U29269 ( .A(n28048), .B(n28044), .Z(n28179) );
  XNOR U29270 ( .A(n28043), .B(n28039), .Z(n28180) );
  XNOR U29271 ( .A(n28038), .B(n28034), .Z(n28181) );
  XNOR U29272 ( .A(n28033), .B(n28029), .Z(n28182) );
  XNOR U29273 ( .A(n28028), .B(n28024), .Z(n28183) );
  XNOR U29274 ( .A(n28023), .B(n28019), .Z(n28184) );
  XNOR U29275 ( .A(n28018), .B(n28014), .Z(n28185) );
  XNOR U29276 ( .A(n28013), .B(n28009), .Z(n28186) );
  XNOR U29277 ( .A(n28008), .B(n28004), .Z(n28187) );
  XNOR U29278 ( .A(n28003), .B(n27999), .Z(n28188) );
  XNOR U29279 ( .A(n27998), .B(n27994), .Z(n28189) );
  XNOR U29280 ( .A(n27993), .B(n27989), .Z(n28190) );
  XNOR U29281 ( .A(n27988), .B(n27984), .Z(n28191) );
  XNOR U29282 ( .A(n27983), .B(n27979), .Z(n28192) );
  XNOR U29283 ( .A(n27978), .B(n27974), .Z(n28193) );
  XNOR U29284 ( .A(n27973), .B(n27969), .Z(n28194) );
  XNOR U29285 ( .A(n27968), .B(n27964), .Z(n28195) );
  XNOR U29286 ( .A(n27963), .B(n27959), .Z(n28196) );
  XNOR U29287 ( .A(n27958), .B(n27954), .Z(n28197) );
  XNOR U29288 ( .A(n27953), .B(n27949), .Z(n28198) );
  XNOR U29289 ( .A(n27948), .B(n27944), .Z(n28199) );
  XNOR U29290 ( .A(n27943), .B(n27939), .Z(n28200) );
  XNOR U29291 ( .A(n27938), .B(n27934), .Z(n28201) );
  XNOR U29292 ( .A(n27933), .B(n27929), .Z(n28202) );
  XNOR U29293 ( .A(n27928), .B(n27924), .Z(n28203) );
  XNOR U29294 ( .A(n27923), .B(n27919), .Z(n28204) );
  XNOR U29295 ( .A(n27918), .B(n27914), .Z(n28205) );
  XNOR U29296 ( .A(n27913), .B(n27909), .Z(n28206) );
  XNOR U29297 ( .A(n28207), .B(n27908), .Z(n27909) );
  AND U29298 ( .A(a[0]), .B(b[50]), .Z(n28207) );
  XNOR U29299 ( .A(n28208), .B(n27908), .Z(n27910) );
  XNOR U29300 ( .A(n28209), .B(n28210), .Z(n27908) );
  AND U29301 ( .A(n28211), .B(n28212), .Z(n28209) );
  AND U29302 ( .A(a[1]), .B(b[49]), .Z(n28208) );
  XOR U29303 ( .A(n28213), .B(n27913), .Z(n27915) );
  XOR U29304 ( .A(n28214), .B(n28215), .Z(n27913) );
  AND U29305 ( .A(n28216), .B(n28217), .Z(n28214) );
  AND U29306 ( .A(a[2]), .B(b[48]), .Z(n28213) );
  XOR U29307 ( .A(n28218), .B(n27918), .Z(n27920) );
  XOR U29308 ( .A(n28219), .B(n28220), .Z(n27918) );
  AND U29309 ( .A(n28221), .B(n28222), .Z(n28219) );
  AND U29310 ( .A(a[3]), .B(b[47]), .Z(n28218) );
  XOR U29311 ( .A(n28223), .B(n27923), .Z(n27925) );
  XOR U29312 ( .A(n28224), .B(n28225), .Z(n27923) );
  AND U29313 ( .A(n28226), .B(n28227), .Z(n28224) );
  AND U29314 ( .A(a[4]), .B(b[46]), .Z(n28223) );
  XOR U29315 ( .A(n28228), .B(n27928), .Z(n27930) );
  XOR U29316 ( .A(n28229), .B(n28230), .Z(n27928) );
  AND U29317 ( .A(n28231), .B(n28232), .Z(n28229) );
  AND U29318 ( .A(a[5]), .B(b[45]), .Z(n28228) );
  XOR U29319 ( .A(n28233), .B(n27933), .Z(n27935) );
  XOR U29320 ( .A(n28234), .B(n28235), .Z(n27933) );
  AND U29321 ( .A(n28236), .B(n28237), .Z(n28234) );
  AND U29322 ( .A(a[6]), .B(b[44]), .Z(n28233) );
  XOR U29323 ( .A(n28238), .B(n27938), .Z(n27940) );
  XOR U29324 ( .A(n28239), .B(n28240), .Z(n27938) );
  AND U29325 ( .A(n28241), .B(n28242), .Z(n28239) );
  AND U29326 ( .A(a[7]), .B(b[43]), .Z(n28238) );
  XOR U29327 ( .A(n28243), .B(n27943), .Z(n27945) );
  XOR U29328 ( .A(n28244), .B(n28245), .Z(n27943) );
  AND U29329 ( .A(n28246), .B(n28247), .Z(n28244) );
  AND U29330 ( .A(a[8]), .B(b[42]), .Z(n28243) );
  XOR U29331 ( .A(n28248), .B(n27948), .Z(n27950) );
  XOR U29332 ( .A(n28249), .B(n28250), .Z(n27948) );
  AND U29333 ( .A(n28251), .B(n28252), .Z(n28249) );
  AND U29334 ( .A(a[9]), .B(b[41]), .Z(n28248) );
  XOR U29335 ( .A(n28253), .B(n27953), .Z(n27955) );
  XOR U29336 ( .A(n28254), .B(n28255), .Z(n27953) );
  AND U29337 ( .A(n28256), .B(n28257), .Z(n28254) );
  AND U29338 ( .A(a[10]), .B(b[40]), .Z(n28253) );
  XOR U29339 ( .A(n28258), .B(n27958), .Z(n27960) );
  XOR U29340 ( .A(n28259), .B(n28260), .Z(n27958) );
  AND U29341 ( .A(n28261), .B(n28262), .Z(n28259) );
  AND U29342 ( .A(a[11]), .B(b[39]), .Z(n28258) );
  XOR U29343 ( .A(n28263), .B(n27963), .Z(n27965) );
  XOR U29344 ( .A(n28264), .B(n28265), .Z(n27963) );
  AND U29345 ( .A(n28266), .B(n28267), .Z(n28264) );
  AND U29346 ( .A(a[12]), .B(b[38]), .Z(n28263) );
  XOR U29347 ( .A(n28268), .B(n27968), .Z(n27970) );
  XOR U29348 ( .A(n28269), .B(n28270), .Z(n27968) );
  AND U29349 ( .A(n28271), .B(n28272), .Z(n28269) );
  AND U29350 ( .A(a[13]), .B(b[37]), .Z(n28268) );
  XOR U29351 ( .A(n28273), .B(n27973), .Z(n27975) );
  XOR U29352 ( .A(n28274), .B(n28275), .Z(n27973) );
  AND U29353 ( .A(n28276), .B(n28277), .Z(n28274) );
  AND U29354 ( .A(a[14]), .B(b[36]), .Z(n28273) );
  XOR U29355 ( .A(n28278), .B(n27978), .Z(n27980) );
  XOR U29356 ( .A(n28279), .B(n28280), .Z(n27978) );
  AND U29357 ( .A(n28281), .B(n28282), .Z(n28279) );
  AND U29358 ( .A(a[15]), .B(b[35]), .Z(n28278) );
  XOR U29359 ( .A(n28283), .B(n27983), .Z(n27985) );
  XOR U29360 ( .A(n28284), .B(n28285), .Z(n27983) );
  AND U29361 ( .A(n28286), .B(n28287), .Z(n28284) );
  AND U29362 ( .A(a[16]), .B(b[34]), .Z(n28283) );
  XOR U29363 ( .A(n28288), .B(n27988), .Z(n27990) );
  XOR U29364 ( .A(n28289), .B(n28290), .Z(n27988) );
  AND U29365 ( .A(n28291), .B(n28292), .Z(n28289) );
  AND U29366 ( .A(a[17]), .B(b[33]), .Z(n28288) );
  XOR U29367 ( .A(n28293), .B(n27993), .Z(n27995) );
  XOR U29368 ( .A(n28294), .B(n28295), .Z(n27993) );
  AND U29369 ( .A(n28296), .B(n28297), .Z(n28294) );
  AND U29370 ( .A(a[18]), .B(b[32]), .Z(n28293) );
  XOR U29371 ( .A(n28298), .B(n27998), .Z(n28000) );
  XOR U29372 ( .A(n28299), .B(n28300), .Z(n27998) );
  AND U29373 ( .A(n28301), .B(n28302), .Z(n28299) );
  AND U29374 ( .A(a[19]), .B(b[31]), .Z(n28298) );
  XOR U29375 ( .A(n28303), .B(n28003), .Z(n28005) );
  XOR U29376 ( .A(n28304), .B(n28305), .Z(n28003) );
  AND U29377 ( .A(n28306), .B(n28307), .Z(n28304) );
  AND U29378 ( .A(a[20]), .B(b[30]), .Z(n28303) );
  XOR U29379 ( .A(n28308), .B(n28008), .Z(n28010) );
  XOR U29380 ( .A(n28309), .B(n28310), .Z(n28008) );
  AND U29381 ( .A(n28311), .B(n28312), .Z(n28309) );
  AND U29382 ( .A(a[21]), .B(b[29]), .Z(n28308) );
  XOR U29383 ( .A(n28313), .B(n28013), .Z(n28015) );
  XOR U29384 ( .A(n28314), .B(n28315), .Z(n28013) );
  AND U29385 ( .A(n28316), .B(n28317), .Z(n28314) );
  AND U29386 ( .A(a[22]), .B(b[28]), .Z(n28313) );
  XOR U29387 ( .A(n28318), .B(n28018), .Z(n28020) );
  XOR U29388 ( .A(n28319), .B(n28320), .Z(n28018) );
  AND U29389 ( .A(n28321), .B(n28322), .Z(n28319) );
  AND U29390 ( .A(a[23]), .B(b[27]), .Z(n28318) );
  XOR U29391 ( .A(n28323), .B(n28023), .Z(n28025) );
  XOR U29392 ( .A(n28324), .B(n28325), .Z(n28023) );
  AND U29393 ( .A(n28326), .B(n28327), .Z(n28324) );
  AND U29394 ( .A(a[24]), .B(b[26]), .Z(n28323) );
  XOR U29395 ( .A(n28328), .B(n28028), .Z(n28030) );
  XOR U29396 ( .A(n28329), .B(n28330), .Z(n28028) );
  AND U29397 ( .A(n28331), .B(n28332), .Z(n28329) );
  AND U29398 ( .A(a[25]), .B(b[25]), .Z(n28328) );
  XOR U29399 ( .A(n28333), .B(n28033), .Z(n28035) );
  XOR U29400 ( .A(n28334), .B(n28335), .Z(n28033) );
  AND U29401 ( .A(n28336), .B(n28337), .Z(n28334) );
  AND U29402 ( .A(b[24]), .B(a[26]), .Z(n28333) );
  XOR U29403 ( .A(n28338), .B(n28038), .Z(n28040) );
  XOR U29404 ( .A(n28339), .B(n28340), .Z(n28038) );
  AND U29405 ( .A(n28341), .B(n28342), .Z(n28339) );
  AND U29406 ( .A(b[23]), .B(a[27]), .Z(n28338) );
  XOR U29407 ( .A(n28343), .B(n28043), .Z(n28045) );
  XOR U29408 ( .A(n28344), .B(n28345), .Z(n28043) );
  AND U29409 ( .A(n28346), .B(n28347), .Z(n28344) );
  AND U29410 ( .A(b[22]), .B(a[28]), .Z(n28343) );
  XOR U29411 ( .A(n28348), .B(n28048), .Z(n28050) );
  XOR U29412 ( .A(n28349), .B(n28350), .Z(n28048) );
  AND U29413 ( .A(n28351), .B(n28352), .Z(n28349) );
  AND U29414 ( .A(b[21]), .B(a[29]), .Z(n28348) );
  XOR U29415 ( .A(n28353), .B(n28053), .Z(n28055) );
  XOR U29416 ( .A(n28354), .B(n28355), .Z(n28053) );
  AND U29417 ( .A(n28356), .B(n28357), .Z(n28354) );
  AND U29418 ( .A(b[20]), .B(a[30]), .Z(n28353) );
  XOR U29419 ( .A(n28358), .B(n28058), .Z(n28060) );
  XOR U29420 ( .A(n28359), .B(n28360), .Z(n28058) );
  AND U29421 ( .A(n28361), .B(n28362), .Z(n28359) );
  AND U29422 ( .A(b[19]), .B(a[31]), .Z(n28358) );
  XOR U29423 ( .A(n28363), .B(n28063), .Z(n28065) );
  XOR U29424 ( .A(n28364), .B(n28365), .Z(n28063) );
  AND U29425 ( .A(n28366), .B(n28367), .Z(n28364) );
  AND U29426 ( .A(b[18]), .B(a[32]), .Z(n28363) );
  XOR U29427 ( .A(n28368), .B(n28068), .Z(n28070) );
  XOR U29428 ( .A(n28369), .B(n28370), .Z(n28068) );
  AND U29429 ( .A(n28371), .B(n28372), .Z(n28369) );
  AND U29430 ( .A(b[17]), .B(a[33]), .Z(n28368) );
  XOR U29431 ( .A(n28373), .B(n28073), .Z(n28075) );
  XOR U29432 ( .A(n28374), .B(n28375), .Z(n28073) );
  AND U29433 ( .A(n28376), .B(n28377), .Z(n28374) );
  AND U29434 ( .A(b[16]), .B(a[34]), .Z(n28373) );
  XOR U29435 ( .A(n28378), .B(n28078), .Z(n28080) );
  XOR U29436 ( .A(n28379), .B(n28380), .Z(n28078) );
  AND U29437 ( .A(n28381), .B(n28382), .Z(n28379) );
  AND U29438 ( .A(b[15]), .B(a[35]), .Z(n28378) );
  XOR U29439 ( .A(n28383), .B(n28083), .Z(n28085) );
  XOR U29440 ( .A(n28384), .B(n28385), .Z(n28083) );
  AND U29441 ( .A(n28386), .B(n28387), .Z(n28384) );
  AND U29442 ( .A(b[14]), .B(a[36]), .Z(n28383) );
  XOR U29443 ( .A(n28388), .B(n28088), .Z(n28090) );
  XOR U29444 ( .A(n28389), .B(n28390), .Z(n28088) );
  AND U29445 ( .A(n28391), .B(n28392), .Z(n28389) );
  AND U29446 ( .A(b[13]), .B(a[37]), .Z(n28388) );
  XOR U29447 ( .A(n28393), .B(n28093), .Z(n28095) );
  XOR U29448 ( .A(n28394), .B(n28395), .Z(n28093) );
  AND U29449 ( .A(n28396), .B(n28397), .Z(n28394) );
  AND U29450 ( .A(b[12]), .B(a[38]), .Z(n28393) );
  XOR U29451 ( .A(n28398), .B(n28098), .Z(n28100) );
  XOR U29452 ( .A(n28399), .B(n28400), .Z(n28098) );
  AND U29453 ( .A(n28401), .B(n28402), .Z(n28399) );
  AND U29454 ( .A(b[11]), .B(a[39]), .Z(n28398) );
  XOR U29455 ( .A(n28403), .B(n28103), .Z(n28105) );
  XOR U29456 ( .A(n28404), .B(n28405), .Z(n28103) );
  AND U29457 ( .A(n28406), .B(n28407), .Z(n28404) );
  AND U29458 ( .A(b[10]), .B(a[40]), .Z(n28403) );
  XOR U29459 ( .A(n28408), .B(n28108), .Z(n28110) );
  XOR U29460 ( .A(n28409), .B(n28410), .Z(n28108) );
  AND U29461 ( .A(n28411), .B(n28412), .Z(n28409) );
  AND U29462 ( .A(b[9]), .B(a[41]), .Z(n28408) );
  XOR U29463 ( .A(n28413), .B(n28113), .Z(n28115) );
  XOR U29464 ( .A(n28414), .B(n28415), .Z(n28113) );
  AND U29465 ( .A(n28416), .B(n28417), .Z(n28414) );
  AND U29466 ( .A(b[8]), .B(a[42]), .Z(n28413) );
  XOR U29467 ( .A(n28418), .B(n28118), .Z(n28120) );
  XOR U29468 ( .A(n28419), .B(n28420), .Z(n28118) );
  AND U29469 ( .A(n28421), .B(n28422), .Z(n28419) );
  AND U29470 ( .A(b[7]), .B(a[43]), .Z(n28418) );
  XOR U29471 ( .A(n28423), .B(n28123), .Z(n28125) );
  XOR U29472 ( .A(n28424), .B(n28425), .Z(n28123) );
  AND U29473 ( .A(n28426), .B(n28427), .Z(n28424) );
  AND U29474 ( .A(b[6]), .B(a[44]), .Z(n28423) );
  XOR U29475 ( .A(n28428), .B(n28128), .Z(n28130) );
  XOR U29476 ( .A(n28429), .B(n28430), .Z(n28128) );
  AND U29477 ( .A(n28431), .B(n28432), .Z(n28429) );
  AND U29478 ( .A(b[5]), .B(a[45]), .Z(n28428) );
  XOR U29479 ( .A(n28433), .B(n28133), .Z(n28135) );
  XOR U29480 ( .A(n28434), .B(n28435), .Z(n28133) );
  AND U29481 ( .A(n28436), .B(n28437), .Z(n28434) );
  AND U29482 ( .A(b[4]), .B(a[46]), .Z(n28433) );
  XNOR U29483 ( .A(n28438), .B(n28439), .Z(n28147) );
  NANDN U29484 ( .A(n28440), .B(n28441), .Z(n28439) );
  XOR U29485 ( .A(n28442), .B(n28138), .Z(n28140) );
  XNOR U29486 ( .A(n28443), .B(n28444), .Z(n28138) );
  AND U29487 ( .A(n28445), .B(n28446), .Z(n28443) );
  AND U29488 ( .A(b[3]), .B(a[47]), .Z(n28442) );
  XOR U29489 ( .A(n28154), .B(n28153), .Z(c[113]) );
  XOR U29490 ( .A(sreg[177]), .B(n28152), .Z(n28153) );
  XOR U29491 ( .A(n28159), .B(n28447), .Z(n28154) );
  XNOR U29492 ( .A(n28158), .B(n28152), .Z(n28447) );
  XOR U29493 ( .A(n28448), .B(n28449), .Z(n28152) );
  NOR U29494 ( .A(n28450), .B(n28451), .Z(n28448) );
  NAND U29495 ( .A(a[49]), .B(b[0]), .Z(n28158) );
  XNOR U29496 ( .A(n28440), .B(n28441), .Z(n28159) );
  XOR U29497 ( .A(n28438), .B(n28452), .Z(n28441) );
  NAND U29498 ( .A(b[1]), .B(a[48]), .Z(n28452) );
  XOR U29499 ( .A(n28446), .B(n28453), .Z(n28440) );
  XOR U29500 ( .A(n28438), .B(n28445), .Z(n28453) );
  XNOR U29501 ( .A(n28454), .B(n28444), .Z(n28445) );
  AND U29502 ( .A(b[2]), .B(a[47]), .Z(n28454) );
  NANDN U29503 ( .A(n28455), .B(n28456), .Z(n28438) );
  XOR U29504 ( .A(n28444), .B(n28436), .Z(n28457) );
  XNOR U29505 ( .A(n28435), .B(n28431), .Z(n28458) );
  XNOR U29506 ( .A(n28430), .B(n28426), .Z(n28459) );
  XNOR U29507 ( .A(n28425), .B(n28421), .Z(n28460) );
  XNOR U29508 ( .A(n28420), .B(n28416), .Z(n28461) );
  XNOR U29509 ( .A(n28415), .B(n28411), .Z(n28462) );
  XNOR U29510 ( .A(n28410), .B(n28406), .Z(n28463) );
  XNOR U29511 ( .A(n28405), .B(n28401), .Z(n28464) );
  XNOR U29512 ( .A(n28400), .B(n28396), .Z(n28465) );
  XNOR U29513 ( .A(n28395), .B(n28391), .Z(n28466) );
  XNOR U29514 ( .A(n28390), .B(n28386), .Z(n28467) );
  XNOR U29515 ( .A(n28385), .B(n28381), .Z(n28468) );
  XNOR U29516 ( .A(n28380), .B(n28376), .Z(n28469) );
  XNOR U29517 ( .A(n28375), .B(n28371), .Z(n28470) );
  XNOR U29518 ( .A(n28370), .B(n28366), .Z(n28471) );
  XNOR U29519 ( .A(n28365), .B(n28361), .Z(n28472) );
  XNOR U29520 ( .A(n28360), .B(n28356), .Z(n28473) );
  XNOR U29521 ( .A(n28355), .B(n28351), .Z(n28474) );
  XNOR U29522 ( .A(n28350), .B(n28346), .Z(n28475) );
  XNOR U29523 ( .A(n28345), .B(n28341), .Z(n28476) );
  XNOR U29524 ( .A(n28340), .B(n28336), .Z(n28477) );
  XNOR U29525 ( .A(n28335), .B(n28331), .Z(n28478) );
  XNOR U29526 ( .A(n28330), .B(n28326), .Z(n28479) );
  XNOR U29527 ( .A(n28325), .B(n28321), .Z(n28480) );
  XNOR U29528 ( .A(n28320), .B(n28316), .Z(n28481) );
  XNOR U29529 ( .A(n28315), .B(n28311), .Z(n28482) );
  XNOR U29530 ( .A(n28310), .B(n28306), .Z(n28483) );
  XNOR U29531 ( .A(n28305), .B(n28301), .Z(n28484) );
  XNOR U29532 ( .A(n28300), .B(n28296), .Z(n28485) );
  XNOR U29533 ( .A(n28295), .B(n28291), .Z(n28486) );
  XNOR U29534 ( .A(n28290), .B(n28286), .Z(n28487) );
  XNOR U29535 ( .A(n28285), .B(n28281), .Z(n28488) );
  XNOR U29536 ( .A(n28280), .B(n28276), .Z(n28489) );
  XNOR U29537 ( .A(n28275), .B(n28271), .Z(n28490) );
  XNOR U29538 ( .A(n28270), .B(n28266), .Z(n28491) );
  XNOR U29539 ( .A(n28265), .B(n28261), .Z(n28492) );
  XNOR U29540 ( .A(n28260), .B(n28256), .Z(n28493) );
  XNOR U29541 ( .A(n28255), .B(n28251), .Z(n28494) );
  XNOR U29542 ( .A(n28250), .B(n28246), .Z(n28495) );
  XNOR U29543 ( .A(n28245), .B(n28241), .Z(n28496) );
  XNOR U29544 ( .A(n28240), .B(n28236), .Z(n28497) );
  XNOR U29545 ( .A(n28235), .B(n28231), .Z(n28498) );
  XNOR U29546 ( .A(n28230), .B(n28226), .Z(n28499) );
  XNOR U29547 ( .A(n28225), .B(n28221), .Z(n28500) );
  XNOR U29548 ( .A(n28220), .B(n28216), .Z(n28501) );
  XNOR U29549 ( .A(n28215), .B(n28211), .Z(n28502) );
  XOR U29550 ( .A(n28503), .B(n28210), .Z(n28211) );
  AND U29551 ( .A(a[0]), .B(b[49]), .Z(n28503) );
  XOR U29552 ( .A(n28504), .B(n28210), .Z(n28212) );
  XNOR U29553 ( .A(n28505), .B(n28506), .Z(n28210) );
  AND U29554 ( .A(n28507), .B(n28508), .Z(n28505) );
  AND U29555 ( .A(a[1]), .B(b[48]), .Z(n28504) );
  XOR U29556 ( .A(n28509), .B(n28215), .Z(n28217) );
  XOR U29557 ( .A(n28510), .B(n28511), .Z(n28215) );
  AND U29558 ( .A(n28512), .B(n28513), .Z(n28510) );
  AND U29559 ( .A(a[2]), .B(b[47]), .Z(n28509) );
  XOR U29560 ( .A(n28514), .B(n28220), .Z(n28222) );
  XOR U29561 ( .A(n28515), .B(n28516), .Z(n28220) );
  AND U29562 ( .A(n28517), .B(n28518), .Z(n28515) );
  AND U29563 ( .A(a[3]), .B(b[46]), .Z(n28514) );
  XOR U29564 ( .A(n28519), .B(n28225), .Z(n28227) );
  XOR U29565 ( .A(n28520), .B(n28521), .Z(n28225) );
  AND U29566 ( .A(n28522), .B(n28523), .Z(n28520) );
  AND U29567 ( .A(a[4]), .B(b[45]), .Z(n28519) );
  XOR U29568 ( .A(n28524), .B(n28230), .Z(n28232) );
  XOR U29569 ( .A(n28525), .B(n28526), .Z(n28230) );
  AND U29570 ( .A(n28527), .B(n28528), .Z(n28525) );
  AND U29571 ( .A(a[5]), .B(b[44]), .Z(n28524) );
  XOR U29572 ( .A(n28529), .B(n28235), .Z(n28237) );
  XOR U29573 ( .A(n28530), .B(n28531), .Z(n28235) );
  AND U29574 ( .A(n28532), .B(n28533), .Z(n28530) );
  AND U29575 ( .A(a[6]), .B(b[43]), .Z(n28529) );
  XOR U29576 ( .A(n28534), .B(n28240), .Z(n28242) );
  XOR U29577 ( .A(n28535), .B(n28536), .Z(n28240) );
  AND U29578 ( .A(n28537), .B(n28538), .Z(n28535) );
  AND U29579 ( .A(a[7]), .B(b[42]), .Z(n28534) );
  XOR U29580 ( .A(n28539), .B(n28245), .Z(n28247) );
  XOR U29581 ( .A(n28540), .B(n28541), .Z(n28245) );
  AND U29582 ( .A(n28542), .B(n28543), .Z(n28540) );
  AND U29583 ( .A(a[8]), .B(b[41]), .Z(n28539) );
  XOR U29584 ( .A(n28544), .B(n28250), .Z(n28252) );
  XOR U29585 ( .A(n28545), .B(n28546), .Z(n28250) );
  AND U29586 ( .A(n28547), .B(n28548), .Z(n28545) );
  AND U29587 ( .A(a[9]), .B(b[40]), .Z(n28544) );
  XOR U29588 ( .A(n28549), .B(n28255), .Z(n28257) );
  XOR U29589 ( .A(n28550), .B(n28551), .Z(n28255) );
  AND U29590 ( .A(n28552), .B(n28553), .Z(n28550) );
  AND U29591 ( .A(a[10]), .B(b[39]), .Z(n28549) );
  XOR U29592 ( .A(n28554), .B(n28260), .Z(n28262) );
  XOR U29593 ( .A(n28555), .B(n28556), .Z(n28260) );
  AND U29594 ( .A(n28557), .B(n28558), .Z(n28555) );
  AND U29595 ( .A(a[11]), .B(b[38]), .Z(n28554) );
  XOR U29596 ( .A(n28559), .B(n28265), .Z(n28267) );
  XOR U29597 ( .A(n28560), .B(n28561), .Z(n28265) );
  AND U29598 ( .A(n28562), .B(n28563), .Z(n28560) );
  AND U29599 ( .A(a[12]), .B(b[37]), .Z(n28559) );
  XOR U29600 ( .A(n28564), .B(n28270), .Z(n28272) );
  XOR U29601 ( .A(n28565), .B(n28566), .Z(n28270) );
  AND U29602 ( .A(n28567), .B(n28568), .Z(n28565) );
  AND U29603 ( .A(a[13]), .B(b[36]), .Z(n28564) );
  XOR U29604 ( .A(n28569), .B(n28275), .Z(n28277) );
  XOR U29605 ( .A(n28570), .B(n28571), .Z(n28275) );
  AND U29606 ( .A(n28572), .B(n28573), .Z(n28570) );
  AND U29607 ( .A(a[14]), .B(b[35]), .Z(n28569) );
  XOR U29608 ( .A(n28574), .B(n28280), .Z(n28282) );
  XOR U29609 ( .A(n28575), .B(n28576), .Z(n28280) );
  AND U29610 ( .A(n28577), .B(n28578), .Z(n28575) );
  AND U29611 ( .A(a[15]), .B(b[34]), .Z(n28574) );
  XOR U29612 ( .A(n28579), .B(n28285), .Z(n28287) );
  XOR U29613 ( .A(n28580), .B(n28581), .Z(n28285) );
  AND U29614 ( .A(n28582), .B(n28583), .Z(n28580) );
  AND U29615 ( .A(a[16]), .B(b[33]), .Z(n28579) );
  XOR U29616 ( .A(n28584), .B(n28290), .Z(n28292) );
  XOR U29617 ( .A(n28585), .B(n28586), .Z(n28290) );
  AND U29618 ( .A(n28587), .B(n28588), .Z(n28585) );
  AND U29619 ( .A(a[17]), .B(b[32]), .Z(n28584) );
  XOR U29620 ( .A(n28589), .B(n28295), .Z(n28297) );
  XOR U29621 ( .A(n28590), .B(n28591), .Z(n28295) );
  AND U29622 ( .A(n28592), .B(n28593), .Z(n28590) );
  AND U29623 ( .A(a[18]), .B(b[31]), .Z(n28589) );
  XOR U29624 ( .A(n28594), .B(n28300), .Z(n28302) );
  XOR U29625 ( .A(n28595), .B(n28596), .Z(n28300) );
  AND U29626 ( .A(n28597), .B(n28598), .Z(n28595) );
  AND U29627 ( .A(a[19]), .B(b[30]), .Z(n28594) );
  XOR U29628 ( .A(n28599), .B(n28305), .Z(n28307) );
  XOR U29629 ( .A(n28600), .B(n28601), .Z(n28305) );
  AND U29630 ( .A(n28602), .B(n28603), .Z(n28600) );
  AND U29631 ( .A(a[20]), .B(b[29]), .Z(n28599) );
  XOR U29632 ( .A(n28604), .B(n28310), .Z(n28312) );
  XOR U29633 ( .A(n28605), .B(n28606), .Z(n28310) );
  AND U29634 ( .A(n28607), .B(n28608), .Z(n28605) );
  AND U29635 ( .A(a[21]), .B(b[28]), .Z(n28604) );
  XOR U29636 ( .A(n28609), .B(n28315), .Z(n28317) );
  XOR U29637 ( .A(n28610), .B(n28611), .Z(n28315) );
  AND U29638 ( .A(n28612), .B(n28613), .Z(n28610) );
  AND U29639 ( .A(a[22]), .B(b[27]), .Z(n28609) );
  XOR U29640 ( .A(n28614), .B(n28320), .Z(n28322) );
  XOR U29641 ( .A(n28615), .B(n28616), .Z(n28320) );
  AND U29642 ( .A(n28617), .B(n28618), .Z(n28615) );
  AND U29643 ( .A(a[23]), .B(b[26]), .Z(n28614) );
  XOR U29644 ( .A(n28619), .B(n28325), .Z(n28327) );
  XOR U29645 ( .A(n28620), .B(n28621), .Z(n28325) );
  AND U29646 ( .A(n28622), .B(n28623), .Z(n28620) );
  AND U29647 ( .A(a[24]), .B(b[25]), .Z(n28619) );
  XOR U29648 ( .A(n28624), .B(n28330), .Z(n28332) );
  XOR U29649 ( .A(n28625), .B(n28626), .Z(n28330) );
  AND U29650 ( .A(n28627), .B(n28628), .Z(n28625) );
  AND U29651 ( .A(b[24]), .B(a[25]), .Z(n28624) );
  XOR U29652 ( .A(n28629), .B(n28335), .Z(n28337) );
  XOR U29653 ( .A(n28630), .B(n28631), .Z(n28335) );
  AND U29654 ( .A(n28632), .B(n28633), .Z(n28630) );
  AND U29655 ( .A(b[23]), .B(a[26]), .Z(n28629) );
  XOR U29656 ( .A(n28634), .B(n28340), .Z(n28342) );
  XOR U29657 ( .A(n28635), .B(n28636), .Z(n28340) );
  AND U29658 ( .A(n28637), .B(n28638), .Z(n28635) );
  AND U29659 ( .A(b[22]), .B(a[27]), .Z(n28634) );
  XOR U29660 ( .A(n28639), .B(n28345), .Z(n28347) );
  XOR U29661 ( .A(n28640), .B(n28641), .Z(n28345) );
  AND U29662 ( .A(n28642), .B(n28643), .Z(n28640) );
  AND U29663 ( .A(b[21]), .B(a[28]), .Z(n28639) );
  XOR U29664 ( .A(n28644), .B(n28350), .Z(n28352) );
  XOR U29665 ( .A(n28645), .B(n28646), .Z(n28350) );
  AND U29666 ( .A(n28647), .B(n28648), .Z(n28645) );
  AND U29667 ( .A(b[20]), .B(a[29]), .Z(n28644) );
  XOR U29668 ( .A(n28649), .B(n28355), .Z(n28357) );
  XOR U29669 ( .A(n28650), .B(n28651), .Z(n28355) );
  AND U29670 ( .A(n28652), .B(n28653), .Z(n28650) );
  AND U29671 ( .A(b[19]), .B(a[30]), .Z(n28649) );
  XOR U29672 ( .A(n28654), .B(n28360), .Z(n28362) );
  XOR U29673 ( .A(n28655), .B(n28656), .Z(n28360) );
  AND U29674 ( .A(n28657), .B(n28658), .Z(n28655) );
  AND U29675 ( .A(b[18]), .B(a[31]), .Z(n28654) );
  XOR U29676 ( .A(n28659), .B(n28365), .Z(n28367) );
  XOR U29677 ( .A(n28660), .B(n28661), .Z(n28365) );
  AND U29678 ( .A(n28662), .B(n28663), .Z(n28660) );
  AND U29679 ( .A(b[17]), .B(a[32]), .Z(n28659) );
  XOR U29680 ( .A(n28664), .B(n28370), .Z(n28372) );
  XOR U29681 ( .A(n28665), .B(n28666), .Z(n28370) );
  AND U29682 ( .A(n28667), .B(n28668), .Z(n28665) );
  AND U29683 ( .A(b[16]), .B(a[33]), .Z(n28664) );
  XOR U29684 ( .A(n28669), .B(n28375), .Z(n28377) );
  XOR U29685 ( .A(n28670), .B(n28671), .Z(n28375) );
  AND U29686 ( .A(n28672), .B(n28673), .Z(n28670) );
  AND U29687 ( .A(b[15]), .B(a[34]), .Z(n28669) );
  XOR U29688 ( .A(n28674), .B(n28380), .Z(n28382) );
  XOR U29689 ( .A(n28675), .B(n28676), .Z(n28380) );
  AND U29690 ( .A(n28677), .B(n28678), .Z(n28675) );
  AND U29691 ( .A(b[14]), .B(a[35]), .Z(n28674) );
  XOR U29692 ( .A(n28679), .B(n28385), .Z(n28387) );
  XOR U29693 ( .A(n28680), .B(n28681), .Z(n28385) );
  AND U29694 ( .A(n28682), .B(n28683), .Z(n28680) );
  AND U29695 ( .A(b[13]), .B(a[36]), .Z(n28679) );
  XOR U29696 ( .A(n28684), .B(n28390), .Z(n28392) );
  XOR U29697 ( .A(n28685), .B(n28686), .Z(n28390) );
  AND U29698 ( .A(n28687), .B(n28688), .Z(n28685) );
  AND U29699 ( .A(b[12]), .B(a[37]), .Z(n28684) );
  XOR U29700 ( .A(n28689), .B(n28395), .Z(n28397) );
  XOR U29701 ( .A(n28690), .B(n28691), .Z(n28395) );
  AND U29702 ( .A(n28692), .B(n28693), .Z(n28690) );
  AND U29703 ( .A(b[11]), .B(a[38]), .Z(n28689) );
  XOR U29704 ( .A(n28694), .B(n28400), .Z(n28402) );
  XOR U29705 ( .A(n28695), .B(n28696), .Z(n28400) );
  AND U29706 ( .A(n28697), .B(n28698), .Z(n28695) );
  AND U29707 ( .A(b[10]), .B(a[39]), .Z(n28694) );
  XOR U29708 ( .A(n28699), .B(n28405), .Z(n28407) );
  XOR U29709 ( .A(n28700), .B(n28701), .Z(n28405) );
  AND U29710 ( .A(n28702), .B(n28703), .Z(n28700) );
  AND U29711 ( .A(b[9]), .B(a[40]), .Z(n28699) );
  XOR U29712 ( .A(n28704), .B(n28410), .Z(n28412) );
  XOR U29713 ( .A(n28705), .B(n28706), .Z(n28410) );
  AND U29714 ( .A(n28707), .B(n28708), .Z(n28705) );
  AND U29715 ( .A(b[8]), .B(a[41]), .Z(n28704) );
  XOR U29716 ( .A(n28709), .B(n28415), .Z(n28417) );
  XOR U29717 ( .A(n28710), .B(n28711), .Z(n28415) );
  AND U29718 ( .A(n28712), .B(n28713), .Z(n28710) );
  AND U29719 ( .A(b[7]), .B(a[42]), .Z(n28709) );
  XOR U29720 ( .A(n28714), .B(n28420), .Z(n28422) );
  XOR U29721 ( .A(n28715), .B(n28716), .Z(n28420) );
  AND U29722 ( .A(n28717), .B(n28718), .Z(n28715) );
  AND U29723 ( .A(b[6]), .B(a[43]), .Z(n28714) );
  XOR U29724 ( .A(n28719), .B(n28425), .Z(n28427) );
  XOR U29725 ( .A(n28720), .B(n28721), .Z(n28425) );
  AND U29726 ( .A(n28722), .B(n28723), .Z(n28720) );
  AND U29727 ( .A(b[5]), .B(a[44]), .Z(n28719) );
  XOR U29728 ( .A(n28724), .B(n28430), .Z(n28432) );
  XOR U29729 ( .A(n28725), .B(n28726), .Z(n28430) );
  AND U29730 ( .A(n28727), .B(n28728), .Z(n28725) );
  AND U29731 ( .A(b[4]), .B(a[45]), .Z(n28724) );
  XNOR U29732 ( .A(n28729), .B(n28730), .Z(n28444) );
  NANDN U29733 ( .A(n28731), .B(n28732), .Z(n28730) );
  XOR U29734 ( .A(n28733), .B(n28435), .Z(n28437) );
  XNOR U29735 ( .A(n28734), .B(n28735), .Z(n28435) );
  AND U29736 ( .A(n28736), .B(n28737), .Z(n28734) );
  AND U29737 ( .A(b[3]), .B(a[46]), .Z(n28733) );
  XOR U29738 ( .A(n28451), .B(n28450), .Z(c[112]) );
  XOR U29739 ( .A(sreg[176]), .B(n28449), .Z(n28450) );
  XOR U29740 ( .A(n28456), .B(n28738), .Z(n28451) );
  XNOR U29741 ( .A(n28455), .B(n28449), .Z(n28738) );
  XOR U29742 ( .A(n28739), .B(n28740), .Z(n28449) );
  NOR U29743 ( .A(n28741), .B(n28742), .Z(n28739) );
  NAND U29744 ( .A(a[48]), .B(b[0]), .Z(n28455) );
  XNOR U29745 ( .A(n28731), .B(n28732), .Z(n28456) );
  XOR U29746 ( .A(n28729), .B(n28743), .Z(n28732) );
  NAND U29747 ( .A(b[1]), .B(a[47]), .Z(n28743) );
  XOR U29748 ( .A(n28737), .B(n28744), .Z(n28731) );
  XOR U29749 ( .A(n28729), .B(n28736), .Z(n28744) );
  XNOR U29750 ( .A(n28745), .B(n28735), .Z(n28736) );
  AND U29751 ( .A(b[2]), .B(a[46]), .Z(n28745) );
  NANDN U29752 ( .A(n28746), .B(n28747), .Z(n28729) );
  XOR U29753 ( .A(n28735), .B(n28727), .Z(n28748) );
  XNOR U29754 ( .A(n28726), .B(n28722), .Z(n28749) );
  XNOR U29755 ( .A(n28721), .B(n28717), .Z(n28750) );
  XNOR U29756 ( .A(n28716), .B(n28712), .Z(n28751) );
  XNOR U29757 ( .A(n28711), .B(n28707), .Z(n28752) );
  XNOR U29758 ( .A(n28706), .B(n28702), .Z(n28753) );
  XNOR U29759 ( .A(n28701), .B(n28697), .Z(n28754) );
  XNOR U29760 ( .A(n28696), .B(n28692), .Z(n28755) );
  XNOR U29761 ( .A(n28691), .B(n28687), .Z(n28756) );
  XNOR U29762 ( .A(n28686), .B(n28682), .Z(n28757) );
  XNOR U29763 ( .A(n28681), .B(n28677), .Z(n28758) );
  XNOR U29764 ( .A(n28676), .B(n28672), .Z(n28759) );
  XNOR U29765 ( .A(n28671), .B(n28667), .Z(n28760) );
  XNOR U29766 ( .A(n28666), .B(n28662), .Z(n28761) );
  XNOR U29767 ( .A(n28661), .B(n28657), .Z(n28762) );
  XNOR U29768 ( .A(n28656), .B(n28652), .Z(n28763) );
  XNOR U29769 ( .A(n28651), .B(n28647), .Z(n28764) );
  XNOR U29770 ( .A(n28646), .B(n28642), .Z(n28765) );
  XNOR U29771 ( .A(n28641), .B(n28637), .Z(n28766) );
  XNOR U29772 ( .A(n28636), .B(n28632), .Z(n28767) );
  XNOR U29773 ( .A(n28631), .B(n28627), .Z(n28768) );
  XNOR U29774 ( .A(n28626), .B(n28622), .Z(n28769) );
  XNOR U29775 ( .A(n28621), .B(n28617), .Z(n28770) );
  XNOR U29776 ( .A(n28616), .B(n28612), .Z(n28771) );
  XNOR U29777 ( .A(n28611), .B(n28607), .Z(n28772) );
  XNOR U29778 ( .A(n28606), .B(n28602), .Z(n28773) );
  XNOR U29779 ( .A(n28601), .B(n28597), .Z(n28774) );
  XNOR U29780 ( .A(n28596), .B(n28592), .Z(n28775) );
  XNOR U29781 ( .A(n28591), .B(n28587), .Z(n28776) );
  XNOR U29782 ( .A(n28586), .B(n28582), .Z(n28777) );
  XNOR U29783 ( .A(n28581), .B(n28577), .Z(n28778) );
  XNOR U29784 ( .A(n28576), .B(n28572), .Z(n28779) );
  XNOR U29785 ( .A(n28571), .B(n28567), .Z(n28780) );
  XNOR U29786 ( .A(n28566), .B(n28562), .Z(n28781) );
  XNOR U29787 ( .A(n28561), .B(n28557), .Z(n28782) );
  XNOR U29788 ( .A(n28556), .B(n28552), .Z(n28783) );
  XNOR U29789 ( .A(n28551), .B(n28547), .Z(n28784) );
  XNOR U29790 ( .A(n28546), .B(n28542), .Z(n28785) );
  XNOR U29791 ( .A(n28541), .B(n28537), .Z(n28786) );
  XNOR U29792 ( .A(n28536), .B(n28532), .Z(n28787) );
  XNOR U29793 ( .A(n28531), .B(n28527), .Z(n28788) );
  XNOR U29794 ( .A(n28526), .B(n28522), .Z(n28789) );
  XNOR U29795 ( .A(n28521), .B(n28517), .Z(n28790) );
  XNOR U29796 ( .A(n28516), .B(n28512), .Z(n28791) );
  XNOR U29797 ( .A(n28511), .B(n28507), .Z(n28792) );
  XNOR U29798 ( .A(n28793), .B(n28506), .Z(n28507) );
  AND U29799 ( .A(a[0]), .B(b[48]), .Z(n28793) );
  XNOR U29800 ( .A(n28794), .B(n28506), .Z(n28508) );
  XNOR U29801 ( .A(n28795), .B(n28796), .Z(n28506) );
  AND U29802 ( .A(n28797), .B(n28798), .Z(n28795) );
  AND U29803 ( .A(a[1]), .B(b[47]), .Z(n28794) );
  XOR U29804 ( .A(n28799), .B(n28511), .Z(n28513) );
  XOR U29805 ( .A(n28800), .B(n28801), .Z(n28511) );
  AND U29806 ( .A(n28802), .B(n28803), .Z(n28800) );
  AND U29807 ( .A(a[2]), .B(b[46]), .Z(n28799) );
  XOR U29808 ( .A(n28804), .B(n28516), .Z(n28518) );
  XOR U29809 ( .A(n28805), .B(n28806), .Z(n28516) );
  AND U29810 ( .A(n28807), .B(n28808), .Z(n28805) );
  AND U29811 ( .A(a[3]), .B(b[45]), .Z(n28804) );
  XOR U29812 ( .A(n28809), .B(n28521), .Z(n28523) );
  XOR U29813 ( .A(n28810), .B(n28811), .Z(n28521) );
  AND U29814 ( .A(n28812), .B(n28813), .Z(n28810) );
  AND U29815 ( .A(a[4]), .B(b[44]), .Z(n28809) );
  XOR U29816 ( .A(n28814), .B(n28526), .Z(n28528) );
  XOR U29817 ( .A(n28815), .B(n28816), .Z(n28526) );
  AND U29818 ( .A(n28817), .B(n28818), .Z(n28815) );
  AND U29819 ( .A(a[5]), .B(b[43]), .Z(n28814) );
  XOR U29820 ( .A(n28819), .B(n28531), .Z(n28533) );
  XOR U29821 ( .A(n28820), .B(n28821), .Z(n28531) );
  AND U29822 ( .A(n28822), .B(n28823), .Z(n28820) );
  AND U29823 ( .A(a[6]), .B(b[42]), .Z(n28819) );
  XOR U29824 ( .A(n28824), .B(n28536), .Z(n28538) );
  XOR U29825 ( .A(n28825), .B(n28826), .Z(n28536) );
  AND U29826 ( .A(n28827), .B(n28828), .Z(n28825) );
  AND U29827 ( .A(a[7]), .B(b[41]), .Z(n28824) );
  XOR U29828 ( .A(n28829), .B(n28541), .Z(n28543) );
  XOR U29829 ( .A(n28830), .B(n28831), .Z(n28541) );
  AND U29830 ( .A(n28832), .B(n28833), .Z(n28830) );
  AND U29831 ( .A(a[8]), .B(b[40]), .Z(n28829) );
  XOR U29832 ( .A(n28834), .B(n28546), .Z(n28548) );
  XOR U29833 ( .A(n28835), .B(n28836), .Z(n28546) );
  AND U29834 ( .A(n28837), .B(n28838), .Z(n28835) );
  AND U29835 ( .A(a[9]), .B(b[39]), .Z(n28834) );
  XOR U29836 ( .A(n28839), .B(n28551), .Z(n28553) );
  XOR U29837 ( .A(n28840), .B(n28841), .Z(n28551) );
  AND U29838 ( .A(n28842), .B(n28843), .Z(n28840) );
  AND U29839 ( .A(a[10]), .B(b[38]), .Z(n28839) );
  XOR U29840 ( .A(n28844), .B(n28556), .Z(n28558) );
  XOR U29841 ( .A(n28845), .B(n28846), .Z(n28556) );
  AND U29842 ( .A(n28847), .B(n28848), .Z(n28845) );
  AND U29843 ( .A(a[11]), .B(b[37]), .Z(n28844) );
  XOR U29844 ( .A(n28849), .B(n28561), .Z(n28563) );
  XOR U29845 ( .A(n28850), .B(n28851), .Z(n28561) );
  AND U29846 ( .A(n28852), .B(n28853), .Z(n28850) );
  AND U29847 ( .A(a[12]), .B(b[36]), .Z(n28849) );
  XOR U29848 ( .A(n28854), .B(n28566), .Z(n28568) );
  XOR U29849 ( .A(n28855), .B(n28856), .Z(n28566) );
  AND U29850 ( .A(n28857), .B(n28858), .Z(n28855) );
  AND U29851 ( .A(a[13]), .B(b[35]), .Z(n28854) );
  XOR U29852 ( .A(n28859), .B(n28571), .Z(n28573) );
  XOR U29853 ( .A(n28860), .B(n28861), .Z(n28571) );
  AND U29854 ( .A(n28862), .B(n28863), .Z(n28860) );
  AND U29855 ( .A(a[14]), .B(b[34]), .Z(n28859) );
  XOR U29856 ( .A(n28864), .B(n28576), .Z(n28578) );
  XOR U29857 ( .A(n28865), .B(n28866), .Z(n28576) );
  AND U29858 ( .A(n28867), .B(n28868), .Z(n28865) );
  AND U29859 ( .A(a[15]), .B(b[33]), .Z(n28864) );
  XOR U29860 ( .A(n28869), .B(n28581), .Z(n28583) );
  XOR U29861 ( .A(n28870), .B(n28871), .Z(n28581) );
  AND U29862 ( .A(n28872), .B(n28873), .Z(n28870) );
  AND U29863 ( .A(a[16]), .B(b[32]), .Z(n28869) );
  XOR U29864 ( .A(n28874), .B(n28586), .Z(n28588) );
  XOR U29865 ( .A(n28875), .B(n28876), .Z(n28586) );
  AND U29866 ( .A(n28877), .B(n28878), .Z(n28875) );
  AND U29867 ( .A(a[17]), .B(b[31]), .Z(n28874) );
  XOR U29868 ( .A(n28879), .B(n28591), .Z(n28593) );
  XOR U29869 ( .A(n28880), .B(n28881), .Z(n28591) );
  AND U29870 ( .A(n28882), .B(n28883), .Z(n28880) );
  AND U29871 ( .A(a[18]), .B(b[30]), .Z(n28879) );
  XOR U29872 ( .A(n28884), .B(n28596), .Z(n28598) );
  XOR U29873 ( .A(n28885), .B(n28886), .Z(n28596) );
  AND U29874 ( .A(n28887), .B(n28888), .Z(n28885) );
  AND U29875 ( .A(a[19]), .B(b[29]), .Z(n28884) );
  XOR U29876 ( .A(n28889), .B(n28601), .Z(n28603) );
  XOR U29877 ( .A(n28890), .B(n28891), .Z(n28601) );
  AND U29878 ( .A(n28892), .B(n28893), .Z(n28890) );
  AND U29879 ( .A(a[20]), .B(b[28]), .Z(n28889) );
  XOR U29880 ( .A(n28894), .B(n28606), .Z(n28608) );
  XOR U29881 ( .A(n28895), .B(n28896), .Z(n28606) );
  AND U29882 ( .A(n28897), .B(n28898), .Z(n28895) );
  AND U29883 ( .A(a[21]), .B(b[27]), .Z(n28894) );
  XOR U29884 ( .A(n28899), .B(n28611), .Z(n28613) );
  XOR U29885 ( .A(n28900), .B(n28901), .Z(n28611) );
  AND U29886 ( .A(n28902), .B(n28903), .Z(n28900) );
  AND U29887 ( .A(a[22]), .B(b[26]), .Z(n28899) );
  XOR U29888 ( .A(n28904), .B(n28616), .Z(n28618) );
  XOR U29889 ( .A(n28905), .B(n28906), .Z(n28616) );
  AND U29890 ( .A(n28907), .B(n28908), .Z(n28905) );
  AND U29891 ( .A(a[23]), .B(b[25]), .Z(n28904) );
  XOR U29892 ( .A(n28909), .B(n28621), .Z(n28623) );
  XOR U29893 ( .A(n28910), .B(n28911), .Z(n28621) );
  AND U29894 ( .A(n28912), .B(n28913), .Z(n28910) );
  AND U29895 ( .A(a[24]), .B(b[24]), .Z(n28909) );
  XOR U29896 ( .A(n28914), .B(n28626), .Z(n28628) );
  XOR U29897 ( .A(n28915), .B(n28916), .Z(n28626) );
  AND U29898 ( .A(n28917), .B(n28918), .Z(n28915) );
  AND U29899 ( .A(b[23]), .B(a[25]), .Z(n28914) );
  XOR U29900 ( .A(n28919), .B(n28631), .Z(n28633) );
  XOR U29901 ( .A(n28920), .B(n28921), .Z(n28631) );
  AND U29902 ( .A(n28922), .B(n28923), .Z(n28920) );
  AND U29903 ( .A(b[22]), .B(a[26]), .Z(n28919) );
  XOR U29904 ( .A(n28924), .B(n28636), .Z(n28638) );
  XOR U29905 ( .A(n28925), .B(n28926), .Z(n28636) );
  AND U29906 ( .A(n28927), .B(n28928), .Z(n28925) );
  AND U29907 ( .A(b[21]), .B(a[27]), .Z(n28924) );
  XOR U29908 ( .A(n28929), .B(n28641), .Z(n28643) );
  XOR U29909 ( .A(n28930), .B(n28931), .Z(n28641) );
  AND U29910 ( .A(n28932), .B(n28933), .Z(n28930) );
  AND U29911 ( .A(b[20]), .B(a[28]), .Z(n28929) );
  XOR U29912 ( .A(n28934), .B(n28646), .Z(n28648) );
  XOR U29913 ( .A(n28935), .B(n28936), .Z(n28646) );
  AND U29914 ( .A(n28937), .B(n28938), .Z(n28935) );
  AND U29915 ( .A(b[19]), .B(a[29]), .Z(n28934) );
  XOR U29916 ( .A(n28939), .B(n28651), .Z(n28653) );
  XOR U29917 ( .A(n28940), .B(n28941), .Z(n28651) );
  AND U29918 ( .A(n28942), .B(n28943), .Z(n28940) );
  AND U29919 ( .A(b[18]), .B(a[30]), .Z(n28939) );
  XOR U29920 ( .A(n28944), .B(n28656), .Z(n28658) );
  XOR U29921 ( .A(n28945), .B(n28946), .Z(n28656) );
  AND U29922 ( .A(n28947), .B(n28948), .Z(n28945) );
  AND U29923 ( .A(b[17]), .B(a[31]), .Z(n28944) );
  XOR U29924 ( .A(n28949), .B(n28661), .Z(n28663) );
  XOR U29925 ( .A(n28950), .B(n28951), .Z(n28661) );
  AND U29926 ( .A(n28952), .B(n28953), .Z(n28950) );
  AND U29927 ( .A(b[16]), .B(a[32]), .Z(n28949) );
  XOR U29928 ( .A(n28954), .B(n28666), .Z(n28668) );
  XOR U29929 ( .A(n28955), .B(n28956), .Z(n28666) );
  AND U29930 ( .A(n28957), .B(n28958), .Z(n28955) );
  AND U29931 ( .A(b[15]), .B(a[33]), .Z(n28954) );
  XOR U29932 ( .A(n28959), .B(n28671), .Z(n28673) );
  XOR U29933 ( .A(n28960), .B(n28961), .Z(n28671) );
  AND U29934 ( .A(n28962), .B(n28963), .Z(n28960) );
  AND U29935 ( .A(b[14]), .B(a[34]), .Z(n28959) );
  XOR U29936 ( .A(n28964), .B(n28676), .Z(n28678) );
  XOR U29937 ( .A(n28965), .B(n28966), .Z(n28676) );
  AND U29938 ( .A(n28967), .B(n28968), .Z(n28965) );
  AND U29939 ( .A(b[13]), .B(a[35]), .Z(n28964) );
  XOR U29940 ( .A(n28969), .B(n28681), .Z(n28683) );
  XOR U29941 ( .A(n28970), .B(n28971), .Z(n28681) );
  AND U29942 ( .A(n28972), .B(n28973), .Z(n28970) );
  AND U29943 ( .A(b[12]), .B(a[36]), .Z(n28969) );
  XOR U29944 ( .A(n28974), .B(n28686), .Z(n28688) );
  XOR U29945 ( .A(n28975), .B(n28976), .Z(n28686) );
  AND U29946 ( .A(n28977), .B(n28978), .Z(n28975) );
  AND U29947 ( .A(b[11]), .B(a[37]), .Z(n28974) );
  XOR U29948 ( .A(n28979), .B(n28691), .Z(n28693) );
  XOR U29949 ( .A(n28980), .B(n28981), .Z(n28691) );
  AND U29950 ( .A(n28982), .B(n28983), .Z(n28980) );
  AND U29951 ( .A(b[10]), .B(a[38]), .Z(n28979) );
  XOR U29952 ( .A(n28984), .B(n28696), .Z(n28698) );
  XOR U29953 ( .A(n28985), .B(n28986), .Z(n28696) );
  AND U29954 ( .A(n28987), .B(n28988), .Z(n28985) );
  AND U29955 ( .A(b[9]), .B(a[39]), .Z(n28984) );
  XOR U29956 ( .A(n28989), .B(n28701), .Z(n28703) );
  XOR U29957 ( .A(n28990), .B(n28991), .Z(n28701) );
  AND U29958 ( .A(n28992), .B(n28993), .Z(n28990) );
  AND U29959 ( .A(b[8]), .B(a[40]), .Z(n28989) );
  XOR U29960 ( .A(n28994), .B(n28706), .Z(n28708) );
  XOR U29961 ( .A(n28995), .B(n28996), .Z(n28706) );
  AND U29962 ( .A(n28997), .B(n28998), .Z(n28995) );
  AND U29963 ( .A(b[7]), .B(a[41]), .Z(n28994) );
  XOR U29964 ( .A(n28999), .B(n28711), .Z(n28713) );
  XOR U29965 ( .A(n29000), .B(n29001), .Z(n28711) );
  AND U29966 ( .A(n29002), .B(n29003), .Z(n29000) );
  AND U29967 ( .A(b[6]), .B(a[42]), .Z(n28999) );
  XOR U29968 ( .A(n29004), .B(n28716), .Z(n28718) );
  XOR U29969 ( .A(n29005), .B(n29006), .Z(n28716) );
  AND U29970 ( .A(n29007), .B(n29008), .Z(n29005) );
  AND U29971 ( .A(b[5]), .B(a[43]), .Z(n29004) );
  XOR U29972 ( .A(n29009), .B(n28721), .Z(n28723) );
  XOR U29973 ( .A(n29010), .B(n29011), .Z(n28721) );
  AND U29974 ( .A(n29012), .B(n29013), .Z(n29010) );
  AND U29975 ( .A(b[4]), .B(a[44]), .Z(n29009) );
  XNOR U29976 ( .A(n29014), .B(n29015), .Z(n28735) );
  NANDN U29977 ( .A(n29016), .B(n29017), .Z(n29015) );
  XOR U29978 ( .A(n29018), .B(n28726), .Z(n28728) );
  XNOR U29979 ( .A(n29019), .B(n29020), .Z(n28726) );
  AND U29980 ( .A(n29021), .B(n29022), .Z(n29019) );
  AND U29981 ( .A(b[3]), .B(a[45]), .Z(n29018) );
  XOR U29982 ( .A(n28742), .B(n28741), .Z(c[111]) );
  XOR U29983 ( .A(sreg[175]), .B(n28740), .Z(n28741) );
  XOR U29984 ( .A(n28747), .B(n29023), .Z(n28742) );
  XNOR U29985 ( .A(n28746), .B(n28740), .Z(n29023) );
  XOR U29986 ( .A(n29024), .B(n29025), .Z(n28740) );
  NOR U29987 ( .A(n29026), .B(n29027), .Z(n29024) );
  NAND U29988 ( .A(a[47]), .B(b[0]), .Z(n28746) );
  XNOR U29989 ( .A(n29016), .B(n29017), .Z(n28747) );
  XOR U29990 ( .A(n29014), .B(n29028), .Z(n29017) );
  NAND U29991 ( .A(b[1]), .B(a[46]), .Z(n29028) );
  XOR U29992 ( .A(n29022), .B(n29029), .Z(n29016) );
  XOR U29993 ( .A(n29014), .B(n29021), .Z(n29029) );
  XNOR U29994 ( .A(n29030), .B(n29020), .Z(n29021) );
  AND U29995 ( .A(b[2]), .B(a[45]), .Z(n29030) );
  NANDN U29996 ( .A(n29031), .B(n29032), .Z(n29014) );
  XOR U29997 ( .A(n29020), .B(n29012), .Z(n29033) );
  XNOR U29998 ( .A(n29011), .B(n29007), .Z(n29034) );
  XNOR U29999 ( .A(n29006), .B(n29002), .Z(n29035) );
  XNOR U30000 ( .A(n29001), .B(n28997), .Z(n29036) );
  XNOR U30001 ( .A(n28996), .B(n28992), .Z(n29037) );
  XNOR U30002 ( .A(n28991), .B(n28987), .Z(n29038) );
  XNOR U30003 ( .A(n28986), .B(n28982), .Z(n29039) );
  XNOR U30004 ( .A(n28981), .B(n28977), .Z(n29040) );
  XNOR U30005 ( .A(n28976), .B(n28972), .Z(n29041) );
  XNOR U30006 ( .A(n28971), .B(n28967), .Z(n29042) );
  XNOR U30007 ( .A(n28966), .B(n28962), .Z(n29043) );
  XNOR U30008 ( .A(n28961), .B(n28957), .Z(n29044) );
  XNOR U30009 ( .A(n28956), .B(n28952), .Z(n29045) );
  XNOR U30010 ( .A(n28951), .B(n28947), .Z(n29046) );
  XNOR U30011 ( .A(n28946), .B(n28942), .Z(n29047) );
  XNOR U30012 ( .A(n28941), .B(n28937), .Z(n29048) );
  XNOR U30013 ( .A(n28936), .B(n28932), .Z(n29049) );
  XNOR U30014 ( .A(n28931), .B(n28927), .Z(n29050) );
  XNOR U30015 ( .A(n28926), .B(n28922), .Z(n29051) );
  XNOR U30016 ( .A(n28921), .B(n28917), .Z(n29052) );
  XNOR U30017 ( .A(n28916), .B(n28912), .Z(n29053) );
  XNOR U30018 ( .A(n28911), .B(n28907), .Z(n29054) );
  XNOR U30019 ( .A(n28906), .B(n28902), .Z(n29055) );
  XNOR U30020 ( .A(n28901), .B(n28897), .Z(n29056) );
  XNOR U30021 ( .A(n28896), .B(n28892), .Z(n29057) );
  XNOR U30022 ( .A(n28891), .B(n28887), .Z(n29058) );
  XNOR U30023 ( .A(n28886), .B(n28882), .Z(n29059) );
  XNOR U30024 ( .A(n28881), .B(n28877), .Z(n29060) );
  XNOR U30025 ( .A(n28876), .B(n28872), .Z(n29061) );
  XNOR U30026 ( .A(n28871), .B(n28867), .Z(n29062) );
  XNOR U30027 ( .A(n28866), .B(n28862), .Z(n29063) );
  XNOR U30028 ( .A(n28861), .B(n28857), .Z(n29064) );
  XNOR U30029 ( .A(n28856), .B(n28852), .Z(n29065) );
  XNOR U30030 ( .A(n28851), .B(n28847), .Z(n29066) );
  XNOR U30031 ( .A(n28846), .B(n28842), .Z(n29067) );
  XNOR U30032 ( .A(n28841), .B(n28837), .Z(n29068) );
  XNOR U30033 ( .A(n28836), .B(n28832), .Z(n29069) );
  XNOR U30034 ( .A(n28831), .B(n28827), .Z(n29070) );
  XNOR U30035 ( .A(n28826), .B(n28822), .Z(n29071) );
  XNOR U30036 ( .A(n28821), .B(n28817), .Z(n29072) );
  XNOR U30037 ( .A(n28816), .B(n28812), .Z(n29073) );
  XNOR U30038 ( .A(n28811), .B(n28807), .Z(n29074) );
  XNOR U30039 ( .A(n28806), .B(n28802), .Z(n29075) );
  XNOR U30040 ( .A(n28801), .B(n28797), .Z(n29076) );
  XOR U30041 ( .A(n29077), .B(n28796), .Z(n28797) );
  AND U30042 ( .A(a[0]), .B(b[47]), .Z(n29077) );
  XOR U30043 ( .A(n29078), .B(n28796), .Z(n28798) );
  XNOR U30044 ( .A(n29079), .B(n29080), .Z(n28796) );
  AND U30045 ( .A(n29081), .B(n29082), .Z(n29079) );
  AND U30046 ( .A(a[1]), .B(b[46]), .Z(n29078) );
  XOR U30047 ( .A(n29083), .B(n28801), .Z(n28803) );
  XOR U30048 ( .A(n29084), .B(n29085), .Z(n28801) );
  AND U30049 ( .A(n29086), .B(n29087), .Z(n29084) );
  AND U30050 ( .A(a[2]), .B(b[45]), .Z(n29083) );
  XOR U30051 ( .A(n29088), .B(n28806), .Z(n28808) );
  XOR U30052 ( .A(n29089), .B(n29090), .Z(n28806) );
  AND U30053 ( .A(n29091), .B(n29092), .Z(n29089) );
  AND U30054 ( .A(a[3]), .B(b[44]), .Z(n29088) );
  XOR U30055 ( .A(n29093), .B(n28811), .Z(n28813) );
  XOR U30056 ( .A(n29094), .B(n29095), .Z(n28811) );
  AND U30057 ( .A(n29096), .B(n29097), .Z(n29094) );
  AND U30058 ( .A(a[4]), .B(b[43]), .Z(n29093) );
  XOR U30059 ( .A(n29098), .B(n28816), .Z(n28818) );
  XOR U30060 ( .A(n29099), .B(n29100), .Z(n28816) );
  AND U30061 ( .A(n29101), .B(n29102), .Z(n29099) );
  AND U30062 ( .A(a[5]), .B(b[42]), .Z(n29098) );
  XOR U30063 ( .A(n29103), .B(n28821), .Z(n28823) );
  XOR U30064 ( .A(n29104), .B(n29105), .Z(n28821) );
  AND U30065 ( .A(n29106), .B(n29107), .Z(n29104) );
  AND U30066 ( .A(a[6]), .B(b[41]), .Z(n29103) );
  XOR U30067 ( .A(n29108), .B(n28826), .Z(n28828) );
  XOR U30068 ( .A(n29109), .B(n29110), .Z(n28826) );
  AND U30069 ( .A(n29111), .B(n29112), .Z(n29109) );
  AND U30070 ( .A(a[7]), .B(b[40]), .Z(n29108) );
  XOR U30071 ( .A(n29113), .B(n28831), .Z(n28833) );
  XOR U30072 ( .A(n29114), .B(n29115), .Z(n28831) );
  AND U30073 ( .A(n29116), .B(n29117), .Z(n29114) );
  AND U30074 ( .A(a[8]), .B(b[39]), .Z(n29113) );
  XOR U30075 ( .A(n29118), .B(n28836), .Z(n28838) );
  XOR U30076 ( .A(n29119), .B(n29120), .Z(n28836) );
  AND U30077 ( .A(n29121), .B(n29122), .Z(n29119) );
  AND U30078 ( .A(a[9]), .B(b[38]), .Z(n29118) );
  XOR U30079 ( .A(n29123), .B(n28841), .Z(n28843) );
  XOR U30080 ( .A(n29124), .B(n29125), .Z(n28841) );
  AND U30081 ( .A(n29126), .B(n29127), .Z(n29124) );
  AND U30082 ( .A(a[10]), .B(b[37]), .Z(n29123) );
  XOR U30083 ( .A(n29128), .B(n28846), .Z(n28848) );
  XOR U30084 ( .A(n29129), .B(n29130), .Z(n28846) );
  AND U30085 ( .A(n29131), .B(n29132), .Z(n29129) );
  AND U30086 ( .A(a[11]), .B(b[36]), .Z(n29128) );
  XOR U30087 ( .A(n29133), .B(n28851), .Z(n28853) );
  XOR U30088 ( .A(n29134), .B(n29135), .Z(n28851) );
  AND U30089 ( .A(n29136), .B(n29137), .Z(n29134) );
  AND U30090 ( .A(a[12]), .B(b[35]), .Z(n29133) );
  XOR U30091 ( .A(n29138), .B(n28856), .Z(n28858) );
  XOR U30092 ( .A(n29139), .B(n29140), .Z(n28856) );
  AND U30093 ( .A(n29141), .B(n29142), .Z(n29139) );
  AND U30094 ( .A(a[13]), .B(b[34]), .Z(n29138) );
  XOR U30095 ( .A(n29143), .B(n28861), .Z(n28863) );
  XOR U30096 ( .A(n29144), .B(n29145), .Z(n28861) );
  AND U30097 ( .A(n29146), .B(n29147), .Z(n29144) );
  AND U30098 ( .A(a[14]), .B(b[33]), .Z(n29143) );
  XOR U30099 ( .A(n29148), .B(n28866), .Z(n28868) );
  XOR U30100 ( .A(n29149), .B(n29150), .Z(n28866) );
  AND U30101 ( .A(n29151), .B(n29152), .Z(n29149) );
  AND U30102 ( .A(a[15]), .B(b[32]), .Z(n29148) );
  XOR U30103 ( .A(n29153), .B(n28871), .Z(n28873) );
  XOR U30104 ( .A(n29154), .B(n29155), .Z(n28871) );
  AND U30105 ( .A(n29156), .B(n29157), .Z(n29154) );
  AND U30106 ( .A(a[16]), .B(b[31]), .Z(n29153) );
  XOR U30107 ( .A(n29158), .B(n28876), .Z(n28878) );
  XOR U30108 ( .A(n29159), .B(n29160), .Z(n28876) );
  AND U30109 ( .A(n29161), .B(n29162), .Z(n29159) );
  AND U30110 ( .A(a[17]), .B(b[30]), .Z(n29158) );
  XOR U30111 ( .A(n29163), .B(n28881), .Z(n28883) );
  XOR U30112 ( .A(n29164), .B(n29165), .Z(n28881) );
  AND U30113 ( .A(n29166), .B(n29167), .Z(n29164) );
  AND U30114 ( .A(a[18]), .B(b[29]), .Z(n29163) );
  XOR U30115 ( .A(n29168), .B(n28886), .Z(n28888) );
  XOR U30116 ( .A(n29169), .B(n29170), .Z(n28886) );
  AND U30117 ( .A(n29171), .B(n29172), .Z(n29169) );
  AND U30118 ( .A(a[19]), .B(b[28]), .Z(n29168) );
  XOR U30119 ( .A(n29173), .B(n28891), .Z(n28893) );
  XOR U30120 ( .A(n29174), .B(n29175), .Z(n28891) );
  AND U30121 ( .A(n29176), .B(n29177), .Z(n29174) );
  AND U30122 ( .A(a[20]), .B(b[27]), .Z(n29173) );
  XOR U30123 ( .A(n29178), .B(n28896), .Z(n28898) );
  XOR U30124 ( .A(n29179), .B(n29180), .Z(n28896) );
  AND U30125 ( .A(n29181), .B(n29182), .Z(n29179) );
  AND U30126 ( .A(a[21]), .B(b[26]), .Z(n29178) );
  XOR U30127 ( .A(n29183), .B(n28901), .Z(n28903) );
  XOR U30128 ( .A(n29184), .B(n29185), .Z(n28901) );
  AND U30129 ( .A(n29186), .B(n29187), .Z(n29184) );
  AND U30130 ( .A(a[22]), .B(b[25]), .Z(n29183) );
  XOR U30131 ( .A(n29188), .B(n28906), .Z(n28908) );
  XOR U30132 ( .A(n29189), .B(n29190), .Z(n28906) );
  AND U30133 ( .A(n29191), .B(n29192), .Z(n29189) );
  AND U30134 ( .A(a[23]), .B(b[24]), .Z(n29188) );
  XOR U30135 ( .A(n29193), .B(n28911), .Z(n28913) );
  XOR U30136 ( .A(n29194), .B(n29195), .Z(n28911) );
  AND U30137 ( .A(n29196), .B(n29197), .Z(n29194) );
  AND U30138 ( .A(b[23]), .B(a[24]), .Z(n29193) );
  XOR U30139 ( .A(n29198), .B(n28916), .Z(n28918) );
  XOR U30140 ( .A(n29199), .B(n29200), .Z(n28916) );
  AND U30141 ( .A(n29201), .B(n29202), .Z(n29199) );
  AND U30142 ( .A(b[22]), .B(a[25]), .Z(n29198) );
  XOR U30143 ( .A(n29203), .B(n28921), .Z(n28923) );
  XOR U30144 ( .A(n29204), .B(n29205), .Z(n28921) );
  AND U30145 ( .A(n29206), .B(n29207), .Z(n29204) );
  AND U30146 ( .A(b[21]), .B(a[26]), .Z(n29203) );
  XOR U30147 ( .A(n29208), .B(n28926), .Z(n28928) );
  XOR U30148 ( .A(n29209), .B(n29210), .Z(n28926) );
  AND U30149 ( .A(n29211), .B(n29212), .Z(n29209) );
  AND U30150 ( .A(b[20]), .B(a[27]), .Z(n29208) );
  XOR U30151 ( .A(n29213), .B(n28931), .Z(n28933) );
  XOR U30152 ( .A(n29214), .B(n29215), .Z(n28931) );
  AND U30153 ( .A(n29216), .B(n29217), .Z(n29214) );
  AND U30154 ( .A(b[19]), .B(a[28]), .Z(n29213) );
  XOR U30155 ( .A(n29218), .B(n28936), .Z(n28938) );
  XOR U30156 ( .A(n29219), .B(n29220), .Z(n28936) );
  AND U30157 ( .A(n29221), .B(n29222), .Z(n29219) );
  AND U30158 ( .A(b[18]), .B(a[29]), .Z(n29218) );
  XOR U30159 ( .A(n29223), .B(n28941), .Z(n28943) );
  XOR U30160 ( .A(n29224), .B(n29225), .Z(n28941) );
  AND U30161 ( .A(n29226), .B(n29227), .Z(n29224) );
  AND U30162 ( .A(b[17]), .B(a[30]), .Z(n29223) );
  XOR U30163 ( .A(n29228), .B(n28946), .Z(n28948) );
  XOR U30164 ( .A(n29229), .B(n29230), .Z(n28946) );
  AND U30165 ( .A(n29231), .B(n29232), .Z(n29229) );
  AND U30166 ( .A(b[16]), .B(a[31]), .Z(n29228) );
  XOR U30167 ( .A(n29233), .B(n28951), .Z(n28953) );
  XOR U30168 ( .A(n29234), .B(n29235), .Z(n28951) );
  AND U30169 ( .A(n29236), .B(n29237), .Z(n29234) );
  AND U30170 ( .A(b[15]), .B(a[32]), .Z(n29233) );
  XOR U30171 ( .A(n29238), .B(n28956), .Z(n28958) );
  XOR U30172 ( .A(n29239), .B(n29240), .Z(n28956) );
  AND U30173 ( .A(n29241), .B(n29242), .Z(n29239) );
  AND U30174 ( .A(b[14]), .B(a[33]), .Z(n29238) );
  XOR U30175 ( .A(n29243), .B(n28961), .Z(n28963) );
  XOR U30176 ( .A(n29244), .B(n29245), .Z(n28961) );
  AND U30177 ( .A(n29246), .B(n29247), .Z(n29244) );
  AND U30178 ( .A(b[13]), .B(a[34]), .Z(n29243) );
  XOR U30179 ( .A(n29248), .B(n28966), .Z(n28968) );
  XOR U30180 ( .A(n29249), .B(n29250), .Z(n28966) );
  AND U30181 ( .A(n29251), .B(n29252), .Z(n29249) );
  AND U30182 ( .A(b[12]), .B(a[35]), .Z(n29248) );
  XOR U30183 ( .A(n29253), .B(n28971), .Z(n28973) );
  XOR U30184 ( .A(n29254), .B(n29255), .Z(n28971) );
  AND U30185 ( .A(n29256), .B(n29257), .Z(n29254) );
  AND U30186 ( .A(b[11]), .B(a[36]), .Z(n29253) );
  XOR U30187 ( .A(n29258), .B(n28976), .Z(n28978) );
  XOR U30188 ( .A(n29259), .B(n29260), .Z(n28976) );
  AND U30189 ( .A(n29261), .B(n29262), .Z(n29259) );
  AND U30190 ( .A(b[10]), .B(a[37]), .Z(n29258) );
  XOR U30191 ( .A(n29263), .B(n28981), .Z(n28983) );
  XOR U30192 ( .A(n29264), .B(n29265), .Z(n28981) );
  AND U30193 ( .A(n29266), .B(n29267), .Z(n29264) );
  AND U30194 ( .A(b[9]), .B(a[38]), .Z(n29263) );
  XOR U30195 ( .A(n29268), .B(n28986), .Z(n28988) );
  XOR U30196 ( .A(n29269), .B(n29270), .Z(n28986) );
  AND U30197 ( .A(n29271), .B(n29272), .Z(n29269) );
  AND U30198 ( .A(b[8]), .B(a[39]), .Z(n29268) );
  XOR U30199 ( .A(n29273), .B(n28991), .Z(n28993) );
  XOR U30200 ( .A(n29274), .B(n29275), .Z(n28991) );
  AND U30201 ( .A(n29276), .B(n29277), .Z(n29274) );
  AND U30202 ( .A(b[7]), .B(a[40]), .Z(n29273) );
  XOR U30203 ( .A(n29278), .B(n28996), .Z(n28998) );
  XOR U30204 ( .A(n29279), .B(n29280), .Z(n28996) );
  AND U30205 ( .A(n29281), .B(n29282), .Z(n29279) );
  AND U30206 ( .A(b[6]), .B(a[41]), .Z(n29278) );
  XOR U30207 ( .A(n29283), .B(n29001), .Z(n29003) );
  XOR U30208 ( .A(n29284), .B(n29285), .Z(n29001) );
  AND U30209 ( .A(n29286), .B(n29287), .Z(n29284) );
  AND U30210 ( .A(b[5]), .B(a[42]), .Z(n29283) );
  XOR U30211 ( .A(n29288), .B(n29006), .Z(n29008) );
  XOR U30212 ( .A(n29289), .B(n29290), .Z(n29006) );
  AND U30213 ( .A(n29291), .B(n29292), .Z(n29289) );
  AND U30214 ( .A(b[4]), .B(a[43]), .Z(n29288) );
  XNOR U30215 ( .A(n29293), .B(n29294), .Z(n29020) );
  NANDN U30216 ( .A(n29295), .B(n29296), .Z(n29294) );
  XOR U30217 ( .A(n29297), .B(n29011), .Z(n29013) );
  XNOR U30218 ( .A(n29298), .B(n29299), .Z(n29011) );
  AND U30219 ( .A(n29300), .B(n29301), .Z(n29298) );
  AND U30220 ( .A(b[3]), .B(a[44]), .Z(n29297) );
  XOR U30221 ( .A(n29027), .B(n29026), .Z(c[110]) );
  XOR U30222 ( .A(sreg[174]), .B(n29025), .Z(n29026) );
  XOR U30223 ( .A(n29032), .B(n29302), .Z(n29027) );
  XNOR U30224 ( .A(n29031), .B(n29025), .Z(n29302) );
  XOR U30225 ( .A(n29303), .B(n29304), .Z(n29025) );
  NOR U30226 ( .A(n29305), .B(n29306), .Z(n29303) );
  NAND U30227 ( .A(a[46]), .B(b[0]), .Z(n29031) );
  XNOR U30228 ( .A(n29295), .B(n29296), .Z(n29032) );
  XOR U30229 ( .A(n29293), .B(n29307), .Z(n29296) );
  NAND U30230 ( .A(b[1]), .B(a[45]), .Z(n29307) );
  XOR U30231 ( .A(n29301), .B(n29308), .Z(n29295) );
  XOR U30232 ( .A(n29293), .B(n29300), .Z(n29308) );
  XNOR U30233 ( .A(n29309), .B(n29299), .Z(n29300) );
  AND U30234 ( .A(b[2]), .B(a[44]), .Z(n29309) );
  NANDN U30235 ( .A(n29310), .B(n29311), .Z(n29293) );
  XOR U30236 ( .A(n29299), .B(n29291), .Z(n29312) );
  XNOR U30237 ( .A(n29290), .B(n29286), .Z(n29313) );
  XNOR U30238 ( .A(n29285), .B(n29281), .Z(n29314) );
  XNOR U30239 ( .A(n29280), .B(n29276), .Z(n29315) );
  XNOR U30240 ( .A(n29275), .B(n29271), .Z(n29316) );
  XNOR U30241 ( .A(n29270), .B(n29266), .Z(n29317) );
  XNOR U30242 ( .A(n29265), .B(n29261), .Z(n29318) );
  XNOR U30243 ( .A(n29260), .B(n29256), .Z(n29319) );
  XNOR U30244 ( .A(n29255), .B(n29251), .Z(n29320) );
  XNOR U30245 ( .A(n29250), .B(n29246), .Z(n29321) );
  XNOR U30246 ( .A(n29245), .B(n29241), .Z(n29322) );
  XNOR U30247 ( .A(n29240), .B(n29236), .Z(n29323) );
  XNOR U30248 ( .A(n29235), .B(n29231), .Z(n29324) );
  XNOR U30249 ( .A(n29230), .B(n29226), .Z(n29325) );
  XNOR U30250 ( .A(n29225), .B(n29221), .Z(n29326) );
  XNOR U30251 ( .A(n29220), .B(n29216), .Z(n29327) );
  XNOR U30252 ( .A(n29215), .B(n29211), .Z(n29328) );
  XNOR U30253 ( .A(n29210), .B(n29206), .Z(n29329) );
  XNOR U30254 ( .A(n29205), .B(n29201), .Z(n29330) );
  XNOR U30255 ( .A(n29200), .B(n29196), .Z(n29331) );
  XNOR U30256 ( .A(n29195), .B(n29191), .Z(n29332) );
  XNOR U30257 ( .A(n29190), .B(n29186), .Z(n29333) );
  XNOR U30258 ( .A(n29185), .B(n29181), .Z(n29334) );
  XNOR U30259 ( .A(n29180), .B(n29176), .Z(n29335) );
  XNOR U30260 ( .A(n29175), .B(n29171), .Z(n29336) );
  XNOR U30261 ( .A(n29170), .B(n29166), .Z(n29337) );
  XNOR U30262 ( .A(n29165), .B(n29161), .Z(n29338) );
  XNOR U30263 ( .A(n29160), .B(n29156), .Z(n29339) );
  XNOR U30264 ( .A(n29155), .B(n29151), .Z(n29340) );
  XNOR U30265 ( .A(n29150), .B(n29146), .Z(n29341) );
  XNOR U30266 ( .A(n29145), .B(n29141), .Z(n29342) );
  XNOR U30267 ( .A(n29140), .B(n29136), .Z(n29343) );
  XNOR U30268 ( .A(n29135), .B(n29131), .Z(n29344) );
  XNOR U30269 ( .A(n29130), .B(n29126), .Z(n29345) );
  XNOR U30270 ( .A(n29125), .B(n29121), .Z(n29346) );
  XNOR U30271 ( .A(n29120), .B(n29116), .Z(n29347) );
  XNOR U30272 ( .A(n29115), .B(n29111), .Z(n29348) );
  XNOR U30273 ( .A(n29110), .B(n29106), .Z(n29349) );
  XNOR U30274 ( .A(n29105), .B(n29101), .Z(n29350) );
  XNOR U30275 ( .A(n29100), .B(n29096), .Z(n29351) );
  XNOR U30276 ( .A(n29095), .B(n29091), .Z(n29352) );
  XNOR U30277 ( .A(n29090), .B(n29086), .Z(n29353) );
  XNOR U30278 ( .A(n29085), .B(n29081), .Z(n29354) );
  XNOR U30279 ( .A(n29355), .B(n29080), .Z(n29081) );
  AND U30280 ( .A(a[0]), .B(b[46]), .Z(n29355) );
  XNOR U30281 ( .A(n29356), .B(n29080), .Z(n29082) );
  XNOR U30282 ( .A(n29357), .B(n29358), .Z(n29080) );
  AND U30283 ( .A(n29359), .B(n29360), .Z(n29357) );
  AND U30284 ( .A(a[1]), .B(b[45]), .Z(n29356) );
  XOR U30285 ( .A(n29361), .B(n29085), .Z(n29087) );
  XOR U30286 ( .A(n29362), .B(n29363), .Z(n29085) );
  AND U30287 ( .A(n29364), .B(n29365), .Z(n29362) );
  AND U30288 ( .A(a[2]), .B(b[44]), .Z(n29361) );
  XOR U30289 ( .A(n29366), .B(n29090), .Z(n29092) );
  XOR U30290 ( .A(n29367), .B(n29368), .Z(n29090) );
  AND U30291 ( .A(n29369), .B(n29370), .Z(n29367) );
  AND U30292 ( .A(a[3]), .B(b[43]), .Z(n29366) );
  XOR U30293 ( .A(n29371), .B(n29095), .Z(n29097) );
  XOR U30294 ( .A(n29372), .B(n29373), .Z(n29095) );
  AND U30295 ( .A(n29374), .B(n29375), .Z(n29372) );
  AND U30296 ( .A(a[4]), .B(b[42]), .Z(n29371) );
  XOR U30297 ( .A(n29376), .B(n29100), .Z(n29102) );
  XOR U30298 ( .A(n29377), .B(n29378), .Z(n29100) );
  AND U30299 ( .A(n29379), .B(n29380), .Z(n29377) );
  AND U30300 ( .A(a[5]), .B(b[41]), .Z(n29376) );
  XOR U30301 ( .A(n29381), .B(n29105), .Z(n29107) );
  XOR U30302 ( .A(n29382), .B(n29383), .Z(n29105) );
  AND U30303 ( .A(n29384), .B(n29385), .Z(n29382) );
  AND U30304 ( .A(a[6]), .B(b[40]), .Z(n29381) );
  XOR U30305 ( .A(n29386), .B(n29110), .Z(n29112) );
  XOR U30306 ( .A(n29387), .B(n29388), .Z(n29110) );
  AND U30307 ( .A(n29389), .B(n29390), .Z(n29387) );
  AND U30308 ( .A(a[7]), .B(b[39]), .Z(n29386) );
  XOR U30309 ( .A(n29391), .B(n29115), .Z(n29117) );
  XOR U30310 ( .A(n29392), .B(n29393), .Z(n29115) );
  AND U30311 ( .A(n29394), .B(n29395), .Z(n29392) );
  AND U30312 ( .A(a[8]), .B(b[38]), .Z(n29391) );
  XOR U30313 ( .A(n29396), .B(n29120), .Z(n29122) );
  XOR U30314 ( .A(n29397), .B(n29398), .Z(n29120) );
  AND U30315 ( .A(n29399), .B(n29400), .Z(n29397) );
  AND U30316 ( .A(a[9]), .B(b[37]), .Z(n29396) );
  XOR U30317 ( .A(n29401), .B(n29125), .Z(n29127) );
  XOR U30318 ( .A(n29402), .B(n29403), .Z(n29125) );
  AND U30319 ( .A(n29404), .B(n29405), .Z(n29402) );
  AND U30320 ( .A(a[10]), .B(b[36]), .Z(n29401) );
  XOR U30321 ( .A(n29406), .B(n29130), .Z(n29132) );
  XOR U30322 ( .A(n29407), .B(n29408), .Z(n29130) );
  AND U30323 ( .A(n29409), .B(n29410), .Z(n29407) );
  AND U30324 ( .A(a[11]), .B(b[35]), .Z(n29406) );
  XOR U30325 ( .A(n29411), .B(n29135), .Z(n29137) );
  XOR U30326 ( .A(n29412), .B(n29413), .Z(n29135) );
  AND U30327 ( .A(n29414), .B(n29415), .Z(n29412) );
  AND U30328 ( .A(a[12]), .B(b[34]), .Z(n29411) );
  XOR U30329 ( .A(n29416), .B(n29140), .Z(n29142) );
  XOR U30330 ( .A(n29417), .B(n29418), .Z(n29140) );
  AND U30331 ( .A(n29419), .B(n29420), .Z(n29417) );
  AND U30332 ( .A(a[13]), .B(b[33]), .Z(n29416) );
  XOR U30333 ( .A(n29421), .B(n29145), .Z(n29147) );
  XOR U30334 ( .A(n29422), .B(n29423), .Z(n29145) );
  AND U30335 ( .A(n29424), .B(n29425), .Z(n29422) );
  AND U30336 ( .A(a[14]), .B(b[32]), .Z(n29421) );
  XOR U30337 ( .A(n29426), .B(n29150), .Z(n29152) );
  XOR U30338 ( .A(n29427), .B(n29428), .Z(n29150) );
  AND U30339 ( .A(n29429), .B(n29430), .Z(n29427) );
  AND U30340 ( .A(a[15]), .B(b[31]), .Z(n29426) );
  XOR U30341 ( .A(n29431), .B(n29155), .Z(n29157) );
  XOR U30342 ( .A(n29432), .B(n29433), .Z(n29155) );
  AND U30343 ( .A(n29434), .B(n29435), .Z(n29432) );
  AND U30344 ( .A(a[16]), .B(b[30]), .Z(n29431) );
  XOR U30345 ( .A(n29436), .B(n29160), .Z(n29162) );
  XOR U30346 ( .A(n29437), .B(n29438), .Z(n29160) );
  AND U30347 ( .A(n29439), .B(n29440), .Z(n29437) );
  AND U30348 ( .A(a[17]), .B(b[29]), .Z(n29436) );
  XOR U30349 ( .A(n29441), .B(n29165), .Z(n29167) );
  XOR U30350 ( .A(n29442), .B(n29443), .Z(n29165) );
  AND U30351 ( .A(n29444), .B(n29445), .Z(n29442) );
  AND U30352 ( .A(a[18]), .B(b[28]), .Z(n29441) );
  XOR U30353 ( .A(n29446), .B(n29170), .Z(n29172) );
  XOR U30354 ( .A(n29447), .B(n29448), .Z(n29170) );
  AND U30355 ( .A(n29449), .B(n29450), .Z(n29447) );
  AND U30356 ( .A(a[19]), .B(b[27]), .Z(n29446) );
  XOR U30357 ( .A(n29451), .B(n29175), .Z(n29177) );
  XOR U30358 ( .A(n29452), .B(n29453), .Z(n29175) );
  AND U30359 ( .A(n29454), .B(n29455), .Z(n29452) );
  AND U30360 ( .A(a[20]), .B(b[26]), .Z(n29451) );
  XOR U30361 ( .A(n29456), .B(n29180), .Z(n29182) );
  XOR U30362 ( .A(n29457), .B(n29458), .Z(n29180) );
  AND U30363 ( .A(n29459), .B(n29460), .Z(n29457) );
  AND U30364 ( .A(a[21]), .B(b[25]), .Z(n29456) );
  XOR U30365 ( .A(n29461), .B(n29185), .Z(n29187) );
  XOR U30366 ( .A(n29462), .B(n29463), .Z(n29185) );
  AND U30367 ( .A(n29464), .B(n29465), .Z(n29462) );
  AND U30368 ( .A(a[22]), .B(b[24]), .Z(n29461) );
  XOR U30369 ( .A(n29466), .B(n29190), .Z(n29192) );
  XOR U30370 ( .A(n29467), .B(n29468), .Z(n29190) );
  AND U30371 ( .A(n29469), .B(n29470), .Z(n29467) );
  AND U30372 ( .A(a[23]), .B(b[23]), .Z(n29466) );
  XOR U30373 ( .A(n29471), .B(n29195), .Z(n29197) );
  XOR U30374 ( .A(n29472), .B(n29473), .Z(n29195) );
  AND U30375 ( .A(n29474), .B(n29475), .Z(n29472) );
  AND U30376 ( .A(b[22]), .B(a[24]), .Z(n29471) );
  XOR U30377 ( .A(n29476), .B(n29200), .Z(n29202) );
  XOR U30378 ( .A(n29477), .B(n29478), .Z(n29200) );
  AND U30379 ( .A(n29479), .B(n29480), .Z(n29477) );
  AND U30380 ( .A(b[21]), .B(a[25]), .Z(n29476) );
  XOR U30381 ( .A(n29481), .B(n29205), .Z(n29207) );
  XOR U30382 ( .A(n29482), .B(n29483), .Z(n29205) );
  AND U30383 ( .A(n29484), .B(n29485), .Z(n29482) );
  AND U30384 ( .A(b[20]), .B(a[26]), .Z(n29481) );
  XOR U30385 ( .A(n29486), .B(n29210), .Z(n29212) );
  XOR U30386 ( .A(n29487), .B(n29488), .Z(n29210) );
  AND U30387 ( .A(n29489), .B(n29490), .Z(n29487) );
  AND U30388 ( .A(b[19]), .B(a[27]), .Z(n29486) );
  XOR U30389 ( .A(n29491), .B(n29215), .Z(n29217) );
  XOR U30390 ( .A(n29492), .B(n29493), .Z(n29215) );
  AND U30391 ( .A(n29494), .B(n29495), .Z(n29492) );
  AND U30392 ( .A(b[18]), .B(a[28]), .Z(n29491) );
  XOR U30393 ( .A(n29496), .B(n29220), .Z(n29222) );
  XOR U30394 ( .A(n29497), .B(n29498), .Z(n29220) );
  AND U30395 ( .A(n29499), .B(n29500), .Z(n29497) );
  AND U30396 ( .A(b[17]), .B(a[29]), .Z(n29496) );
  XOR U30397 ( .A(n29501), .B(n29225), .Z(n29227) );
  XOR U30398 ( .A(n29502), .B(n29503), .Z(n29225) );
  AND U30399 ( .A(n29504), .B(n29505), .Z(n29502) );
  AND U30400 ( .A(b[16]), .B(a[30]), .Z(n29501) );
  XOR U30401 ( .A(n29506), .B(n29230), .Z(n29232) );
  XOR U30402 ( .A(n29507), .B(n29508), .Z(n29230) );
  AND U30403 ( .A(n29509), .B(n29510), .Z(n29507) );
  AND U30404 ( .A(b[15]), .B(a[31]), .Z(n29506) );
  XOR U30405 ( .A(n29511), .B(n29235), .Z(n29237) );
  XOR U30406 ( .A(n29512), .B(n29513), .Z(n29235) );
  AND U30407 ( .A(n29514), .B(n29515), .Z(n29512) );
  AND U30408 ( .A(b[14]), .B(a[32]), .Z(n29511) );
  XOR U30409 ( .A(n29516), .B(n29240), .Z(n29242) );
  XOR U30410 ( .A(n29517), .B(n29518), .Z(n29240) );
  AND U30411 ( .A(n29519), .B(n29520), .Z(n29517) );
  AND U30412 ( .A(b[13]), .B(a[33]), .Z(n29516) );
  XOR U30413 ( .A(n29521), .B(n29245), .Z(n29247) );
  XOR U30414 ( .A(n29522), .B(n29523), .Z(n29245) );
  AND U30415 ( .A(n29524), .B(n29525), .Z(n29522) );
  AND U30416 ( .A(b[12]), .B(a[34]), .Z(n29521) );
  XOR U30417 ( .A(n29526), .B(n29250), .Z(n29252) );
  XOR U30418 ( .A(n29527), .B(n29528), .Z(n29250) );
  AND U30419 ( .A(n29529), .B(n29530), .Z(n29527) );
  AND U30420 ( .A(b[11]), .B(a[35]), .Z(n29526) );
  XOR U30421 ( .A(n29531), .B(n29255), .Z(n29257) );
  XOR U30422 ( .A(n29532), .B(n29533), .Z(n29255) );
  AND U30423 ( .A(n29534), .B(n29535), .Z(n29532) );
  AND U30424 ( .A(b[10]), .B(a[36]), .Z(n29531) );
  XOR U30425 ( .A(n29536), .B(n29260), .Z(n29262) );
  XOR U30426 ( .A(n29537), .B(n29538), .Z(n29260) );
  AND U30427 ( .A(n29539), .B(n29540), .Z(n29537) );
  AND U30428 ( .A(b[9]), .B(a[37]), .Z(n29536) );
  XOR U30429 ( .A(n29541), .B(n29265), .Z(n29267) );
  XOR U30430 ( .A(n29542), .B(n29543), .Z(n29265) );
  AND U30431 ( .A(n29544), .B(n29545), .Z(n29542) );
  AND U30432 ( .A(b[8]), .B(a[38]), .Z(n29541) );
  XOR U30433 ( .A(n29546), .B(n29270), .Z(n29272) );
  XOR U30434 ( .A(n29547), .B(n29548), .Z(n29270) );
  AND U30435 ( .A(n29549), .B(n29550), .Z(n29547) );
  AND U30436 ( .A(b[7]), .B(a[39]), .Z(n29546) );
  XOR U30437 ( .A(n29551), .B(n29275), .Z(n29277) );
  XOR U30438 ( .A(n29552), .B(n29553), .Z(n29275) );
  AND U30439 ( .A(n29554), .B(n29555), .Z(n29552) );
  AND U30440 ( .A(b[6]), .B(a[40]), .Z(n29551) );
  XOR U30441 ( .A(n29556), .B(n29280), .Z(n29282) );
  XOR U30442 ( .A(n29557), .B(n29558), .Z(n29280) );
  AND U30443 ( .A(n29559), .B(n29560), .Z(n29557) );
  AND U30444 ( .A(b[5]), .B(a[41]), .Z(n29556) );
  XOR U30445 ( .A(n29561), .B(n29285), .Z(n29287) );
  XOR U30446 ( .A(n29562), .B(n29563), .Z(n29285) );
  AND U30447 ( .A(n29564), .B(n29565), .Z(n29562) );
  AND U30448 ( .A(b[4]), .B(a[42]), .Z(n29561) );
  XNOR U30449 ( .A(n29566), .B(n29567), .Z(n29299) );
  NANDN U30450 ( .A(n29568), .B(n29569), .Z(n29567) );
  XOR U30451 ( .A(n29570), .B(n29290), .Z(n29292) );
  XNOR U30452 ( .A(n29571), .B(n29572), .Z(n29290) );
  AND U30453 ( .A(n29573), .B(n29574), .Z(n29571) );
  AND U30454 ( .A(b[3]), .B(a[43]), .Z(n29570) );
  XOR U30455 ( .A(n29306), .B(n29305), .Z(c[109]) );
  XOR U30456 ( .A(sreg[173]), .B(n29304), .Z(n29305) );
  XOR U30457 ( .A(n29311), .B(n29575), .Z(n29306) );
  XNOR U30458 ( .A(n29310), .B(n29304), .Z(n29575) );
  XOR U30459 ( .A(n29576), .B(n29577), .Z(n29304) );
  NOR U30460 ( .A(n29578), .B(n29579), .Z(n29576) );
  NAND U30461 ( .A(a[45]), .B(b[0]), .Z(n29310) );
  XNOR U30462 ( .A(n29568), .B(n29569), .Z(n29311) );
  XOR U30463 ( .A(n29566), .B(n29580), .Z(n29569) );
  NAND U30464 ( .A(b[1]), .B(a[44]), .Z(n29580) );
  XOR U30465 ( .A(n29574), .B(n29581), .Z(n29568) );
  XOR U30466 ( .A(n29566), .B(n29573), .Z(n29581) );
  XNOR U30467 ( .A(n29582), .B(n29572), .Z(n29573) );
  AND U30468 ( .A(b[2]), .B(a[43]), .Z(n29582) );
  NANDN U30469 ( .A(n29583), .B(n29584), .Z(n29566) );
  XOR U30470 ( .A(n29572), .B(n29564), .Z(n29585) );
  XNOR U30471 ( .A(n29563), .B(n29559), .Z(n29586) );
  XNOR U30472 ( .A(n29558), .B(n29554), .Z(n29587) );
  XNOR U30473 ( .A(n29553), .B(n29549), .Z(n29588) );
  XNOR U30474 ( .A(n29548), .B(n29544), .Z(n29589) );
  XNOR U30475 ( .A(n29543), .B(n29539), .Z(n29590) );
  XNOR U30476 ( .A(n29538), .B(n29534), .Z(n29591) );
  XNOR U30477 ( .A(n29533), .B(n29529), .Z(n29592) );
  XNOR U30478 ( .A(n29528), .B(n29524), .Z(n29593) );
  XNOR U30479 ( .A(n29523), .B(n29519), .Z(n29594) );
  XNOR U30480 ( .A(n29518), .B(n29514), .Z(n29595) );
  XNOR U30481 ( .A(n29513), .B(n29509), .Z(n29596) );
  XNOR U30482 ( .A(n29508), .B(n29504), .Z(n29597) );
  XNOR U30483 ( .A(n29503), .B(n29499), .Z(n29598) );
  XNOR U30484 ( .A(n29498), .B(n29494), .Z(n29599) );
  XNOR U30485 ( .A(n29493), .B(n29489), .Z(n29600) );
  XNOR U30486 ( .A(n29488), .B(n29484), .Z(n29601) );
  XNOR U30487 ( .A(n29483), .B(n29479), .Z(n29602) );
  XNOR U30488 ( .A(n29478), .B(n29474), .Z(n29603) );
  XNOR U30489 ( .A(n29473), .B(n29469), .Z(n29604) );
  XNOR U30490 ( .A(n29468), .B(n29464), .Z(n29605) );
  XNOR U30491 ( .A(n29463), .B(n29459), .Z(n29606) );
  XNOR U30492 ( .A(n29458), .B(n29454), .Z(n29607) );
  XNOR U30493 ( .A(n29453), .B(n29449), .Z(n29608) );
  XNOR U30494 ( .A(n29448), .B(n29444), .Z(n29609) );
  XNOR U30495 ( .A(n29443), .B(n29439), .Z(n29610) );
  XNOR U30496 ( .A(n29438), .B(n29434), .Z(n29611) );
  XNOR U30497 ( .A(n29433), .B(n29429), .Z(n29612) );
  XNOR U30498 ( .A(n29428), .B(n29424), .Z(n29613) );
  XNOR U30499 ( .A(n29423), .B(n29419), .Z(n29614) );
  XNOR U30500 ( .A(n29418), .B(n29414), .Z(n29615) );
  XNOR U30501 ( .A(n29413), .B(n29409), .Z(n29616) );
  XNOR U30502 ( .A(n29408), .B(n29404), .Z(n29617) );
  XNOR U30503 ( .A(n29403), .B(n29399), .Z(n29618) );
  XNOR U30504 ( .A(n29398), .B(n29394), .Z(n29619) );
  XNOR U30505 ( .A(n29393), .B(n29389), .Z(n29620) );
  XNOR U30506 ( .A(n29388), .B(n29384), .Z(n29621) );
  XNOR U30507 ( .A(n29383), .B(n29379), .Z(n29622) );
  XNOR U30508 ( .A(n29378), .B(n29374), .Z(n29623) );
  XNOR U30509 ( .A(n29373), .B(n29369), .Z(n29624) );
  XNOR U30510 ( .A(n29368), .B(n29364), .Z(n29625) );
  XNOR U30511 ( .A(n29363), .B(n29359), .Z(n29626) );
  XOR U30512 ( .A(n29627), .B(n29358), .Z(n29359) );
  AND U30513 ( .A(a[0]), .B(b[45]), .Z(n29627) );
  XOR U30514 ( .A(n29628), .B(n29358), .Z(n29360) );
  XNOR U30515 ( .A(n29629), .B(n29630), .Z(n29358) );
  AND U30516 ( .A(n29631), .B(n29632), .Z(n29629) );
  AND U30517 ( .A(a[1]), .B(b[44]), .Z(n29628) );
  XOR U30518 ( .A(n29633), .B(n29363), .Z(n29365) );
  XOR U30519 ( .A(n29634), .B(n29635), .Z(n29363) );
  AND U30520 ( .A(n29636), .B(n29637), .Z(n29634) );
  AND U30521 ( .A(a[2]), .B(b[43]), .Z(n29633) );
  XOR U30522 ( .A(n29638), .B(n29368), .Z(n29370) );
  XOR U30523 ( .A(n29639), .B(n29640), .Z(n29368) );
  AND U30524 ( .A(n29641), .B(n29642), .Z(n29639) );
  AND U30525 ( .A(a[3]), .B(b[42]), .Z(n29638) );
  XOR U30526 ( .A(n29643), .B(n29373), .Z(n29375) );
  XOR U30527 ( .A(n29644), .B(n29645), .Z(n29373) );
  AND U30528 ( .A(n29646), .B(n29647), .Z(n29644) );
  AND U30529 ( .A(a[4]), .B(b[41]), .Z(n29643) );
  XOR U30530 ( .A(n29648), .B(n29378), .Z(n29380) );
  XOR U30531 ( .A(n29649), .B(n29650), .Z(n29378) );
  AND U30532 ( .A(n29651), .B(n29652), .Z(n29649) );
  AND U30533 ( .A(a[5]), .B(b[40]), .Z(n29648) );
  XOR U30534 ( .A(n29653), .B(n29383), .Z(n29385) );
  XOR U30535 ( .A(n29654), .B(n29655), .Z(n29383) );
  AND U30536 ( .A(n29656), .B(n29657), .Z(n29654) );
  AND U30537 ( .A(a[6]), .B(b[39]), .Z(n29653) );
  XOR U30538 ( .A(n29658), .B(n29388), .Z(n29390) );
  XOR U30539 ( .A(n29659), .B(n29660), .Z(n29388) );
  AND U30540 ( .A(n29661), .B(n29662), .Z(n29659) );
  AND U30541 ( .A(a[7]), .B(b[38]), .Z(n29658) );
  XOR U30542 ( .A(n29663), .B(n29393), .Z(n29395) );
  XOR U30543 ( .A(n29664), .B(n29665), .Z(n29393) );
  AND U30544 ( .A(n29666), .B(n29667), .Z(n29664) );
  AND U30545 ( .A(a[8]), .B(b[37]), .Z(n29663) );
  XOR U30546 ( .A(n29668), .B(n29398), .Z(n29400) );
  XOR U30547 ( .A(n29669), .B(n29670), .Z(n29398) );
  AND U30548 ( .A(n29671), .B(n29672), .Z(n29669) );
  AND U30549 ( .A(a[9]), .B(b[36]), .Z(n29668) );
  XOR U30550 ( .A(n29673), .B(n29403), .Z(n29405) );
  XOR U30551 ( .A(n29674), .B(n29675), .Z(n29403) );
  AND U30552 ( .A(n29676), .B(n29677), .Z(n29674) );
  AND U30553 ( .A(a[10]), .B(b[35]), .Z(n29673) );
  XOR U30554 ( .A(n29678), .B(n29408), .Z(n29410) );
  XOR U30555 ( .A(n29679), .B(n29680), .Z(n29408) );
  AND U30556 ( .A(n29681), .B(n29682), .Z(n29679) );
  AND U30557 ( .A(a[11]), .B(b[34]), .Z(n29678) );
  XOR U30558 ( .A(n29683), .B(n29413), .Z(n29415) );
  XOR U30559 ( .A(n29684), .B(n29685), .Z(n29413) );
  AND U30560 ( .A(n29686), .B(n29687), .Z(n29684) );
  AND U30561 ( .A(a[12]), .B(b[33]), .Z(n29683) );
  XOR U30562 ( .A(n29688), .B(n29418), .Z(n29420) );
  XOR U30563 ( .A(n29689), .B(n29690), .Z(n29418) );
  AND U30564 ( .A(n29691), .B(n29692), .Z(n29689) );
  AND U30565 ( .A(a[13]), .B(b[32]), .Z(n29688) );
  XOR U30566 ( .A(n29693), .B(n29423), .Z(n29425) );
  XOR U30567 ( .A(n29694), .B(n29695), .Z(n29423) );
  AND U30568 ( .A(n29696), .B(n29697), .Z(n29694) );
  AND U30569 ( .A(a[14]), .B(b[31]), .Z(n29693) );
  XOR U30570 ( .A(n29698), .B(n29428), .Z(n29430) );
  XOR U30571 ( .A(n29699), .B(n29700), .Z(n29428) );
  AND U30572 ( .A(n29701), .B(n29702), .Z(n29699) );
  AND U30573 ( .A(a[15]), .B(b[30]), .Z(n29698) );
  XOR U30574 ( .A(n29703), .B(n29433), .Z(n29435) );
  XOR U30575 ( .A(n29704), .B(n29705), .Z(n29433) );
  AND U30576 ( .A(n29706), .B(n29707), .Z(n29704) );
  AND U30577 ( .A(a[16]), .B(b[29]), .Z(n29703) );
  XOR U30578 ( .A(n29708), .B(n29438), .Z(n29440) );
  XOR U30579 ( .A(n29709), .B(n29710), .Z(n29438) );
  AND U30580 ( .A(n29711), .B(n29712), .Z(n29709) );
  AND U30581 ( .A(a[17]), .B(b[28]), .Z(n29708) );
  XOR U30582 ( .A(n29713), .B(n29443), .Z(n29445) );
  XOR U30583 ( .A(n29714), .B(n29715), .Z(n29443) );
  AND U30584 ( .A(n29716), .B(n29717), .Z(n29714) );
  AND U30585 ( .A(a[18]), .B(b[27]), .Z(n29713) );
  XOR U30586 ( .A(n29718), .B(n29448), .Z(n29450) );
  XOR U30587 ( .A(n29719), .B(n29720), .Z(n29448) );
  AND U30588 ( .A(n29721), .B(n29722), .Z(n29719) );
  AND U30589 ( .A(a[19]), .B(b[26]), .Z(n29718) );
  XOR U30590 ( .A(n29723), .B(n29453), .Z(n29455) );
  XOR U30591 ( .A(n29724), .B(n29725), .Z(n29453) );
  AND U30592 ( .A(n29726), .B(n29727), .Z(n29724) );
  AND U30593 ( .A(a[20]), .B(b[25]), .Z(n29723) );
  XOR U30594 ( .A(n29728), .B(n29458), .Z(n29460) );
  XOR U30595 ( .A(n29729), .B(n29730), .Z(n29458) );
  AND U30596 ( .A(n29731), .B(n29732), .Z(n29729) );
  AND U30597 ( .A(a[21]), .B(b[24]), .Z(n29728) );
  XOR U30598 ( .A(n29733), .B(n29463), .Z(n29465) );
  XOR U30599 ( .A(n29734), .B(n29735), .Z(n29463) );
  AND U30600 ( .A(n29736), .B(n29737), .Z(n29734) );
  AND U30601 ( .A(a[22]), .B(b[23]), .Z(n29733) );
  XOR U30602 ( .A(n29738), .B(n29468), .Z(n29470) );
  XOR U30603 ( .A(n29739), .B(n29740), .Z(n29468) );
  AND U30604 ( .A(n29741), .B(n29742), .Z(n29739) );
  AND U30605 ( .A(b[22]), .B(a[23]), .Z(n29738) );
  XOR U30606 ( .A(n29743), .B(n29473), .Z(n29475) );
  XOR U30607 ( .A(n29744), .B(n29745), .Z(n29473) );
  AND U30608 ( .A(n29746), .B(n29747), .Z(n29744) );
  AND U30609 ( .A(b[21]), .B(a[24]), .Z(n29743) );
  XOR U30610 ( .A(n29748), .B(n29478), .Z(n29480) );
  XOR U30611 ( .A(n29749), .B(n29750), .Z(n29478) );
  AND U30612 ( .A(n29751), .B(n29752), .Z(n29749) );
  AND U30613 ( .A(b[20]), .B(a[25]), .Z(n29748) );
  XOR U30614 ( .A(n29753), .B(n29483), .Z(n29485) );
  XOR U30615 ( .A(n29754), .B(n29755), .Z(n29483) );
  AND U30616 ( .A(n29756), .B(n29757), .Z(n29754) );
  AND U30617 ( .A(b[19]), .B(a[26]), .Z(n29753) );
  XOR U30618 ( .A(n29758), .B(n29488), .Z(n29490) );
  XOR U30619 ( .A(n29759), .B(n29760), .Z(n29488) );
  AND U30620 ( .A(n29761), .B(n29762), .Z(n29759) );
  AND U30621 ( .A(b[18]), .B(a[27]), .Z(n29758) );
  XOR U30622 ( .A(n29763), .B(n29493), .Z(n29495) );
  XOR U30623 ( .A(n29764), .B(n29765), .Z(n29493) );
  AND U30624 ( .A(n29766), .B(n29767), .Z(n29764) );
  AND U30625 ( .A(b[17]), .B(a[28]), .Z(n29763) );
  XOR U30626 ( .A(n29768), .B(n29498), .Z(n29500) );
  XOR U30627 ( .A(n29769), .B(n29770), .Z(n29498) );
  AND U30628 ( .A(n29771), .B(n29772), .Z(n29769) );
  AND U30629 ( .A(b[16]), .B(a[29]), .Z(n29768) );
  XOR U30630 ( .A(n29773), .B(n29503), .Z(n29505) );
  XOR U30631 ( .A(n29774), .B(n29775), .Z(n29503) );
  AND U30632 ( .A(n29776), .B(n29777), .Z(n29774) );
  AND U30633 ( .A(b[15]), .B(a[30]), .Z(n29773) );
  XOR U30634 ( .A(n29778), .B(n29508), .Z(n29510) );
  XOR U30635 ( .A(n29779), .B(n29780), .Z(n29508) );
  AND U30636 ( .A(n29781), .B(n29782), .Z(n29779) );
  AND U30637 ( .A(b[14]), .B(a[31]), .Z(n29778) );
  XOR U30638 ( .A(n29783), .B(n29513), .Z(n29515) );
  XOR U30639 ( .A(n29784), .B(n29785), .Z(n29513) );
  AND U30640 ( .A(n29786), .B(n29787), .Z(n29784) );
  AND U30641 ( .A(b[13]), .B(a[32]), .Z(n29783) );
  XOR U30642 ( .A(n29788), .B(n29518), .Z(n29520) );
  XOR U30643 ( .A(n29789), .B(n29790), .Z(n29518) );
  AND U30644 ( .A(n29791), .B(n29792), .Z(n29789) );
  AND U30645 ( .A(b[12]), .B(a[33]), .Z(n29788) );
  XOR U30646 ( .A(n29793), .B(n29523), .Z(n29525) );
  XOR U30647 ( .A(n29794), .B(n29795), .Z(n29523) );
  AND U30648 ( .A(n29796), .B(n29797), .Z(n29794) );
  AND U30649 ( .A(b[11]), .B(a[34]), .Z(n29793) );
  XOR U30650 ( .A(n29798), .B(n29528), .Z(n29530) );
  XOR U30651 ( .A(n29799), .B(n29800), .Z(n29528) );
  AND U30652 ( .A(n29801), .B(n29802), .Z(n29799) );
  AND U30653 ( .A(b[10]), .B(a[35]), .Z(n29798) );
  XOR U30654 ( .A(n29803), .B(n29533), .Z(n29535) );
  XOR U30655 ( .A(n29804), .B(n29805), .Z(n29533) );
  AND U30656 ( .A(n29806), .B(n29807), .Z(n29804) );
  AND U30657 ( .A(b[9]), .B(a[36]), .Z(n29803) );
  XOR U30658 ( .A(n29808), .B(n29538), .Z(n29540) );
  XOR U30659 ( .A(n29809), .B(n29810), .Z(n29538) );
  AND U30660 ( .A(n29811), .B(n29812), .Z(n29809) );
  AND U30661 ( .A(b[8]), .B(a[37]), .Z(n29808) );
  XOR U30662 ( .A(n29813), .B(n29543), .Z(n29545) );
  XOR U30663 ( .A(n29814), .B(n29815), .Z(n29543) );
  AND U30664 ( .A(n29816), .B(n29817), .Z(n29814) );
  AND U30665 ( .A(b[7]), .B(a[38]), .Z(n29813) );
  XOR U30666 ( .A(n29818), .B(n29548), .Z(n29550) );
  XOR U30667 ( .A(n29819), .B(n29820), .Z(n29548) );
  AND U30668 ( .A(n29821), .B(n29822), .Z(n29819) );
  AND U30669 ( .A(b[6]), .B(a[39]), .Z(n29818) );
  XOR U30670 ( .A(n29823), .B(n29553), .Z(n29555) );
  XOR U30671 ( .A(n29824), .B(n29825), .Z(n29553) );
  AND U30672 ( .A(n29826), .B(n29827), .Z(n29824) );
  AND U30673 ( .A(b[5]), .B(a[40]), .Z(n29823) );
  XOR U30674 ( .A(n29828), .B(n29558), .Z(n29560) );
  XOR U30675 ( .A(n29829), .B(n29830), .Z(n29558) );
  AND U30676 ( .A(n29831), .B(n29832), .Z(n29829) );
  AND U30677 ( .A(b[4]), .B(a[41]), .Z(n29828) );
  XNOR U30678 ( .A(n29833), .B(n29834), .Z(n29572) );
  NANDN U30679 ( .A(n29835), .B(n29836), .Z(n29834) );
  XOR U30680 ( .A(n29837), .B(n29563), .Z(n29565) );
  XNOR U30681 ( .A(n29838), .B(n29839), .Z(n29563) );
  AND U30682 ( .A(n29840), .B(n29841), .Z(n29838) );
  AND U30683 ( .A(b[3]), .B(a[42]), .Z(n29837) );
  XOR U30684 ( .A(n29579), .B(n29578), .Z(c[108]) );
  XOR U30685 ( .A(sreg[172]), .B(n29577), .Z(n29578) );
  XOR U30686 ( .A(n29584), .B(n29842), .Z(n29579) );
  XNOR U30687 ( .A(n29583), .B(n29577), .Z(n29842) );
  XOR U30688 ( .A(n29843), .B(n29844), .Z(n29577) );
  NOR U30689 ( .A(n29845), .B(n29846), .Z(n29843) );
  NAND U30690 ( .A(a[44]), .B(b[0]), .Z(n29583) );
  XNOR U30691 ( .A(n29835), .B(n29836), .Z(n29584) );
  XOR U30692 ( .A(n29833), .B(n29847), .Z(n29836) );
  NAND U30693 ( .A(b[1]), .B(a[43]), .Z(n29847) );
  XOR U30694 ( .A(n29841), .B(n29848), .Z(n29835) );
  XOR U30695 ( .A(n29833), .B(n29840), .Z(n29848) );
  XNOR U30696 ( .A(n29849), .B(n29839), .Z(n29840) );
  AND U30697 ( .A(b[2]), .B(a[42]), .Z(n29849) );
  NANDN U30698 ( .A(n29850), .B(n29851), .Z(n29833) );
  XOR U30699 ( .A(n29839), .B(n29831), .Z(n29852) );
  XNOR U30700 ( .A(n29830), .B(n29826), .Z(n29853) );
  XNOR U30701 ( .A(n29825), .B(n29821), .Z(n29854) );
  XNOR U30702 ( .A(n29820), .B(n29816), .Z(n29855) );
  XNOR U30703 ( .A(n29815), .B(n29811), .Z(n29856) );
  XNOR U30704 ( .A(n29810), .B(n29806), .Z(n29857) );
  XNOR U30705 ( .A(n29805), .B(n29801), .Z(n29858) );
  XNOR U30706 ( .A(n29800), .B(n29796), .Z(n29859) );
  XNOR U30707 ( .A(n29795), .B(n29791), .Z(n29860) );
  XNOR U30708 ( .A(n29790), .B(n29786), .Z(n29861) );
  XNOR U30709 ( .A(n29785), .B(n29781), .Z(n29862) );
  XNOR U30710 ( .A(n29780), .B(n29776), .Z(n29863) );
  XNOR U30711 ( .A(n29775), .B(n29771), .Z(n29864) );
  XNOR U30712 ( .A(n29770), .B(n29766), .Z(n29865) );
  XNOR U30713 ( .A(n29765), .B(n29761), .Z(n29866) );
  XNOR U30714 ( .A(n29760), .B(n29756), .Z(n29867) );
  XNOR U30715 ( .A(n29755), .B(n29751), .Z(n29868) );
  XNOR U30716 ( .A(n29750), .B(n29746), .Z(n29869) );
  XNOR U30717 ( .A(n29745), .B(n29741), .Z(n29870) );
  XNOR U30718 ( .A(n29740), .B(n29736), .Z(n29871) );
  XNOR U30719 ( .A(n29735), .B(n29731), .Z(n29872) );
  XNOR U30720 ( .A(n29730), .B(n29726), .Z(n29873) );
  XNOR U30721 ( .A(n29725), .B(n29721), .Z(n29874) );
  XNOR U30722 ( .A(n29720), .B(n29716), .Z(n29875) );
  XNOR U30723 ( .A(n29715), .B(n29711), .Z(n29876) );
  XNOR U30724 ( .A(n29710), .B(n29706), .Z(n29877) );
  XNOR U30725 ( .A(n29705), .B(n29701), .Z(n29878) );
  XNOR U30726 ( .A(n29700), .B(n29696), .Z(n29879) );
  XNOR U30727 ( .A(n29695), .B(n29691), .Z(n29880) );
  XNOR U30728 ( .A(n29690), .B(n29686), .Z(n29881) );
  XNOR U30729 ( .A(n29685), .B(n29681), .Z(n29882) );
  XNOR U30730 ( .A(n29680), .B(n29676), .Z(n29883) );
  XNOR U30731 ( .A(n29675), .B(n29671), .Z(n29884) );
  XNOR U30732 ( .A(n29670), .B(n29666), .Z(n29885) );
  XNOR U30733 ( .A(n29665), .B(n29661), .Z(n29886) );
  XNOR U30734 ( .A(n29660), .B(n29656), .Z(n29887) );
  XNOR U30735 ( .A(n29655), .B(n29651), .Z(n29888) );
  XNOR U30736 ( .A(n29650), .B(n29646), .Z(n29889) );
  XNOR U30737 ( .A(n29645), .B(n29641), .Z(n29890) );
  XNOR U30738 ( .A(n29640), .B(n29636), .Z(n29891) );
  XNOR U30739 ( .A(n29635), .B(n29631), .Z(n29892) );
  XNOR U30740 ( .A(n29893), .B(n29630), .Z(n29631) );
  AND U30741 ( .A(a[0]), .B(b[44]), .Z(n29893) );
  XNOR U30742 ( .A(n29894), .B(n29630), .Z(n29632) );
  XNOR U30743 ( .A(n29895), .B(n29896), .Z(n29630) );
  AND U30744 ( .A(n29897), .B(n29898), .Z(n29895) );
  AND U30745 ( .A(a[1]), .B(b[43]), .Z(n29894) );
  XOR U30746 ( .A(n29899), .B(n29635), .Z(n29637) );
  XOR U30747 ( .A(n29900), .B(n29901), .Z(n29635) );
  AND U30748 ( .A(n29902), .B(n29903), .Z(n29900) );
  AND U30749 ( .A(a[2]), .B(b[42]), .Z(n29899) );
  XOR U30750 ( .A(n29904), .B(n29640), .Z(n29642) );
  XOR U30751 ( .A(n29905), .B(n29906), .Z(n29640) );
  AND U30752 ( .A(n29907), .B(n29908), .Z(n29905) );
  AND U30753 ( .A(a[3]), .B(b[41]), .Z(n29904) );
  XOR U30754 ( .A(n29909), .B(n29645), .Z(n29647) );
  XOR U30755 ( .A(n29910), .B(n29911), .Z(n29645) );
  AND U30756 ( .A(n29912), .B(n29913), .Z(n29910) );
  AND U30757 ( .A(a[4]), .B(b[40]), .Z(n29909) );
  XOR U30758 ( .A(n29914), .B(n29650), .Z(n29652) );
  XOR U30759 ( .A(n29915), .B(n29916), .Z(n29650) );
  AND U30760 ( .A(n29917), .B(n29918), .Z(n29915) );
  AND U30761 ( .A(a[5]), .B(b[39]), .Z(n29914) );
  XOR U30762 ( .A(n29919), .B(n29655), .Z(n29657) );
  XOR U30763 ( .A(n29920), .B(n29921), .Z(n29655) );
  AND U30764 ( .A(n29922), .B(n29923), .Z(n29920) );
  AND U30765 ( .A(a[6]), .B(b[38]), .Z(n29919) );
  XOR U30766 ( .A(n29924), .B(n29660), .Z(n29662) );
  XOR U30767 ( .A(n29925), .B(n29926), .Z(n29660) );
  AND U30768 ( .A(n29927), .B(n29928), .Z(n29925) );
  AND U30769 ( .A(a[7]), .B(b[37]), .Z(n29924) );
  XOR U30770 ( .A(n29929), .B(n29665), .Z(n29667) );
  XOR U30771 ( .A(n29930), .B(n29931), .Z(n29665) );
  AND U30772 ( .A(n29932), .B(n29933), .Z(n29930) );
  AND U30773 ( .A(a[8]), .B(b[36]), .Z(n29929) );
  XOR U30774 ( .A(n29934), .B(n29670), .Z(n29672) );
  XOR U30775 ( .A(n29935), .B(n29936), .Z(n29670) );
  AND U30776 ( .A(n29937), .B(n29938), .Z(n29935) );
  AND U30777 ( .A(a[9]), .B(b[35]), .Z(n29934) );
  XOR U30778 ( .A(n29939), .B(n29675), .Z(n29677) );
  XOR U30779 ( .A(n29940), .B(n29941), .Z(n29675) );
  AND U30780 ( .A(n29942), .B(n29943), .Z(n29940) );
  AND U30781 ( .A(a[10]), .B(b[34]), .Z(n29939) );
  XOR U30782 ( .A(n29944), .B(n29680), .Z(n29682) );
  XOR U30783 ( .A(n29945), .B(n29946), .Z(n29680) );
  AND U30784 ( .A(n29947), .B(n29948), .Z(n29945) );
  AND U30785 ( .A(a[11]), .B(b[33]), .Z(n29944) );
  XOR U30786 ( .A(n29949), .B(n29685), .Z(n29687) );
  XOR U30787 ( .A(n29950), .B(n29951), .Z(n29685) );
  AND U30788 ( .A(n29952), .B(n29953), .Z(n29950) );
  AND U30789 ( .A(a[12]), .B(b[32]), .Z(n29949) );
  XOR U30790 ( .A(n29954), .B(n29690), .Z(n29692) );
  XOR U30791 ( .A(n29955), .B(n29956), .Z(n29690) );
  AND U30792 ( .A(n29957), .B(n29958), .Z(n29955) );
  AND U30793 ( .A(a[13]), .B(b[31]), .Z(n29954) );
  XOR U30794 ( .A(n29959), .B(n29695), .Z(n29697) );
  XOR U30795 ( .A(n29960), .B(n29961), .Z(n29695) );
  AND U30796 ( .A(n29962), .B(n29963), .Z(n29960) );
  AND U30797 ( .A(a[14]), .B(b[30]), .Z(n29959) );
  XOR U30798 ( .A(n29964), .B(n29700), .Z(n29702) );
  XOR U30799 ( .A(n29965), .B(n29966), .Z(n29700) );
  AND U30800 ( .A(n29967), .B(n29968), .Z(n29965) );
  AND U30801 ( .A(a[15]), .B(b[29]), .Z(n29964) );
  XOR U30802 ( .A(n29969), .B(n29705), .Z(n29707) );
  XOR U30803 ( .A(n29970), .B(n29971), .Z(n29705) );
  AND U30804 ( .A(n29972), .B(n29973), .Z(n29970) );
  AND U30805 ( .A(a[16]), .B(b[28]), .Z(n29969) );
  XOR U30806 ( .A(n29974), .B(n29710), .Z(n29712) );
  XOR U30807 ( .A(n29975), .B(n29976), .Z(n29710) );
  AND U30808 ( .A(n29977), .B(n29978), .Z(n29975) );
  AND U30809 ( .A(a[17]), .B(b[27]), .Z(n29974) );
  XOR U30810 ( .A(n29979), .B(n29715), .Z(n29717) );
  XOR U30811 ( .A(n29980), .B(n29981), .Z(n29715) );
  AND U30812 ( .A(n29982), .B(n29983), .Z(n29980) );
  AND U30813 ( .A(a[18]), .B(b[26]), .Z(n29979) );
  XOR U30814 ( .A(n29984), .B(n29720), .Z(n29722) );
  XOR U30815 ( .A(n29985), .B(n29986), .Z(n29720) );
  AND U30816 ( .A(n29987), .B(n29988), .Z(n29985) );
  AND U30817 ( .A(a[19]), .B(b[25]), .Z(n29984) );
  XOR U30818 ( .A(n29989), .B(n29725), .Z(n29727) );
  XOR U30819 ( .A(n29990), .B(n29991), .Z(n29725) );
  AND U30820 ( .A(n29992), .B(n29993), .Z(n29990) );
  AND U30821 ( .A(a[20]), .B(b[24]), .Z(n29989) );
  XOR U30822 ( .A(n29994), .B(n29730), .Z(n29732) );
  XOR U30823 ( .A(n29995), .B(n29996), .Z(n29730) );
  AND U30824 ( .A(n29997), .B(n29998), .Z(n29995) );
  AND U30825 ( .A(a[21]), .B(b[23]), .Z(n29994) );
  XOR U30826 ( .A(n29999), .B(n29735), .Z(n29737) );
  XOR U30827 ( .A(n30000), .B(n30001), .Z(n29735) );
  AND U30828 ( .A(n30002), .B(n30003), .Z(n30000) );
  AND U30829 ( .A(a[22]), .B(b[22]), .Z(n29999) );
  XOR U30830 ( .A(n30004), .B(n29740), .Z(n29742) );
  XOR U30831 ( .A(n30005), .B(n30006), .Z(n29740) );
  AND U30832 ( .A(n30007), .B(n30008), .Z(n30005) );
  AND U30833 ( .A(b[21]), .B(a[23]), .Z(n30004) );
  XOR U30834 ( .A(n30009), .B(n29745), .Z(n29747) );
  XOR U30835 ( .A(n30010), .B(n30011), .Z(n29745) );
  AND U30836 ( .A(n30012), .B(n30013), .Z(n30010) );
  AND U30837 ( .A(b[20]), .B(a[24]), .Z(n30009) );
  XOR U30838 ( .A(n30014), .B(n29750), .Z(n29752) );
  XOR U30839 ( .A(n30015), .B(n30016), .Z(n29750) );
  AND U30840 ( .A(n30017), .B(n30018), .Z(n30015) );
  AND U30841 ( .A(b[19]), .B(a[25]), .Z(n30014) );
  XOR U30842 ( .A(n30019), .B(n29755), .Z(n29757) );
  XOR U30843 ( .A(n30020), .B(n30021), .Z(n29755) );
  AND U30844 ( .A(n30022), .B(n30023), .Z(n30020) );
  AND U30845 ( .A(b[18]), .B(a[26]), .Z(n30019) );
  XOR U30846 ( .A(n30024), .B(n29760), .Z(n29762) );
  XOR U30847 ( .A(n30025), .B(n30026), .Z(n29760) );
  AND U30848 ( .A(n30027), .B(n30028), .Z(n30025) );
  AND U30849 ( .A(b[17]), .B(a[27]), .Z(n30024) );
  XOR U30850 ( .A(n30029), .B(n29765), .Z(n29767) );
  XOR U30851 ( .A(n30030), .B(n30031), .Z(n29765) );
  AND U30852 ( .A(n30032), .B(n30033), .Z(n30030) );
  AND U30853 ( .A(b[16]), .B(a[28]), .Z(n30029) );
  XOR U30854 ( .A(n30034), .B(n29770), .Z(n29772) );
  XOR U30855 ( .A(n30035), .B(n30036), .Z(n29770) );
  AND U30856 ( .A(n30037), .B(n30038), .Z(n30035) );
  AND U30857 ( .A(b[15]), .B(a[29]), .Z(n30034) );
  XOR U30858 ( .A(n30039), .B(n29775), .Z(n29777) );
  XOR U30859 ( .A(n30040), .B(n30041), .Z(n29775) );
  AND U30860 ( .A(n30042), .B(n30043), .Z(n30040) );
  AND U30861 ( .A(b[14]), .B(a[30]), .Z(n30039) );
  XOR U30862 ( .A(n30044), .B(n29780), .Z(n29782) );
  XOR U30863 ( .A(n30045), .B(n30046), .Z(n29780) );
  AND U30864 ( .A(n30047), .B(n30048), .Z(n30045) );
  AND U30865 ( .A(b[13]), .B(a[31]), .Z(n30044) );
  XOR U30866 ( .A(n30049), .B(n29785), .Z(n29787) );
  XOR U30867 ( .A(n30050), .B(n30051), .Z(n29785) );
  AND U30868 ( .A(n30052), .B(n30053), .Z(n30050) );
  AND U30869 ( .A(b[12]), .B(a[32]), .Z(n30049) );
  XOR U30870 ( .A(n30054), .B(n29790), .Z(n29792) );
  XOR U30871 ( .A(n30055), .B(n30056), .Z(n29790) );
  AND U30872 ( .A(n30057), .B(n30058), .Z(n30055) );
  AND U30873 ( .A(b[11]), .B(a[33]), .Z(n30054) );
  XOR U30874 ( .A(n30059), .B(n29795), .Z(n29797) );
  XOR U30875 ( .A(n30060), .B(n30061), .Z(n29795) );
  AND U30876 ( .A(n30062), .B(n30063), .Z(n30060) );
  AND U30877 ( .A(b[10]), .B(a[34]), .Z(n30059) );
  XOR U30878 ( .A(n30064), .B(n29800), .Z(n29802) );
  XOR U30879 ( .A(n30065), .B(n30066), .Z(n29800) );
  AND U30880 ( .A(n30067), .B(n30068), .Z(n30065) );
  AND U30881 ( .A(b[9]), .B(a[35]), .Z(n30064) );
  XOR U30882 ( .A(n30069), .B(n29805), .Z(n29807) );
  XOR U30883 ( .A(n30070), .B(n30071), .Z(n29805) );
  AND U30884 ( .A(n30072), .B(n30073), .Z(n30070) );
  AND U30885 ( .A(b[8]), .B(a[36]), .Z(n30069) );
  XOR U30886 ( .A(n30074), .B(n29810), .Z(n29812) );
  XOR U30887 ( .A(n30075), .B(n30076), .Z(n29810) );
  AND U30888 ( .A(n30077), .B(n30078), .Z(n30075) );
  AND U30889 ( .A(b[7]), .B(a[37]), .Z(n30074) );
  XOR U30890 ( .A(n30079), .B(n29815), .Z(n29817) );
  XOR U30891 ( .A(n30080), .B(n30081), .Z(n29815) );
  AND U30892 ( .A(n30082), .B(n30083), .Z(n30080) );
  AND U30893 ( .A(b[6]), .B(a[38]), .Z(n30079) );
  XOR U30894 ( .A(n30084), .B(n29820), .Z(n29822) );
  XOR U30895 ( .A(n30085), .B(n30086), .Z(n29820) );
  AND U30896 ( .A(n30087), .B(n30088), .Z(n30085) );
  AND U30897 ( .A(b[5]), .B(a[39]), .Z(n30084) );
  XOR U30898 ( .A(n30089), .B(n29825), .Z(n29827) );
  XOR U30899 ( .A(n30090), .B(n30091), .Z(n29825) );
  AND U30900 ( .A(n30092), .B(n30093), .Z(n30090) );
  AND U30901 ( .A(b[4]), .B(a[40]), .Z(n30089) );
  XNOR U30902 ( .A(n30094), .B(n30095), .Z(n29839) );
  NANDN U30903 ( .A(n30096), .B(n30097), .Z(n30095) );
  XOR U30904 ( .A(n30098), .B(n29830), .Z(n29832) );
  XNOR U30905 ( .A(n30099), .B(n30100), .Z(n29830) );
  AND U30906 ( .A(n30101), .B(n30102), .Z(n30099) );
  AND U30907 ( .A(b[3]), .B(a[41]), .Z(n30098) );
  XOR U30908 ( .A(n29846), .B(n29845), .Z(c[107]) );
  XOR U30909 ( .A(sreg[171]), .B(n29844), .Z(n29845) );
  XOR U30910 ( .A(n29851), .B(n30103), .Z(n29846) );
  XNOR U30911 ( .A(n29850), .B(n29844), .Z(n30103) );
  XOR U30912 ( .A(n30104), .B(n30105), .Z(n29844) );
  NOR U30913 ( .A(n30106), .B(n30107), .Z(n30104) );
  NAND U30914 ( .A(a[43]), .B(b[0]), .Z(n29850) );
  XNOR U30915 ( .A(n30096), .B(n30097), .Z(n29851) );
  XOR U30916 ( .A(n30094), .B(n30108), .Z(n30097) );
  NAND U30917 ( .A(b[1]), .B(a[42]), .Z(n30108) );
  XOR U30918 ( .A(n30102), .B(n30109), .Z(n30096) );
  XOR U30919 ( .A(n30094), .B(n30101), .Z(n30109) );
  XNOR U30920 ( .A(n30110), .B(n30100), .Z(n30101) );
  AND U30921 ( .A(b[2]), .B(a[41]), .Z(n30110) );
  NANDN U30922 ( .A(n30111), .B(n30112), .Z(n30094) );
  XOR U30923 ( .A(n30100), .B(n30092), .Z(n30113) );
  XNOR U30924 ( .A(n30091), .B(n30087), .Z(n30114) );
  XNOR U30925 ( .A(n30086), .B(n30082), .Z(n30115) );
  XNOR U30926 ( .A(n30081), .B(n30077), .Z(n30116) );
  XNOR U30927 ( .A(n30076), .B(n30072), .Z(n30117) );
  XNOR U30928 ( .A(n30071), .B(n30067), .Z(n30118) );
  XNOR U30929 ( .A(n30066), .B(n30062), .Z(n30119) );
  XNOR U30930 ( .A(n30061), .B(n30057), .Z(n30120) );
  XNOR U30931 ( .A(n30056), .B(n30052), .Z(n30121) );
  XNOR U30932 ( .A(n30051), .B(n30047), .Z(n30122) );
  XNOR U30933 ( .A(n30046), .B(n30042), .Z(n30123) );
  XNOR U30934 ( .A(n30041), .B(n30037), .Z(n30124) );
  XNOR U30935 ( .A(n30036), .B(n30032), .Z(n30125) );
  XNOR U30936 ( .A(n30031), .B(n30027), .Z(n30126) );
  XNOR U30937 ( .A(n30026), .B(n30022), .Z(n30127) );
  XNOR U30938 ( .A(n30021), .B(n30017), .Z(n30128) );
  XNOR U30939 ( .A(n30016), .B(n30012), .Z(n30129) );
  XNOR U30940 ( .A(n30011), .B(n30007), .Z(n30130) );
  XNOR U30941 ( .A(n30006), .B(n30002), .Z(n30131) );
  XNOR U30942 ( .A(n30001), .B(n29997), .Z(n30132) );
  XNOR U30943 ( .A(n29996), .B(n29992), .Z(n30133) );
  XNOR U30944 ( .A(n29991), .B(n29987), .Z(n30134) );
  XNOR U30945 ( .A(n29986), .B(n29982), .Z(n30135) );
  XNOR U30946 ( .A(n29981), .B(n29977), .Z(n30136) );
  XNOR U30947 ( .A(n29976), .B(n29972), .Z(n30137) );
  XNOR U30948 ( .A(n29971), .B(n29967), .Z(n30138) );
  XNOR U30949 ( .A(n29966), .B(n29962), .Z(n30139) );
  XNOR U30950 ( .A(n29961), .B(n29957), .Z(n30140) );
  XNOR U30951 ( .A(n29956), .B(n29952), .Z(n30141) );
  XNOR U30952 ( .A(n29951), .B(n29947), .Z(n30142) );
  XNOR U30953 ( .A(n29946), .B(n29942), .Z(n30143) );
  XNOR U30954 ( .A(n29941), .B(n29937), .Z(n30144) );
  XNOR U30955 ( .A(n29936), .B(n29932), .Z(n30145) );
  XNOR U30956 ( .A(n29931), .B(n29927), .Z(n30146) );
  XNOR U30957 ( .A(n29926), .B(n29922), .Z(n30147) );
  XNOR U30958 ( .A(n29921), .B(n29917), .Z(n30148) );
  XNOR U30959 ( .A(n29916), .B(n29912), .Z(n30149) );
  XNOR U30960 ( .A(n29911), .B(n29907), .Z(n30150) );
  XNOR U30961 ( .A(n29906), .B(n29902), .Z(n30151) );
  XNOR U30962 ( .A(n29901), .B(n29897), .Z(n30152) );
  XOR U30963 ( .A(n30153), .B(n29896), .Z(n29897) );
  AND U30964 ( .A(a[0]), .B(b[43]), .Z(n30153) );
  XOR U30965 ( .A(n30154), .B(n29896), .Z(n29898) );
  XNOR U30966 ( .A(n30155), .B(n30156), .Z(n29896) );
  AND U30967 ( .A(n30157), .B(n30158), .Z(n30155) );
  AND U30968 ( .A(a[1]), .B(b[42]), .Z(n30154) );
  XOR U30969 ( .A(n30159), .B(n29901), .Z(n29903) );
  XOR U30970 ( .A(n30160), .B(n30161), .Z(n29901) );
  AND U30971 ( .A(n30162), .B(n30163), .Z(n30160) );
  AND U30972 ( .A(a[2]), .B(b[41]), .Z(n30159) );
  XOR U30973 ( .A(n30164), .B(n29906), .Z(n29908) );
  XOR U30974 ( .A(n30165), .B(n30166), .Z(n29906) );
  AND U30975 ( .A(n30167), .B(n30168), .Z(n30165) );
  AND U30976 ( .A(a[3]), .B(b[40]), .Z(n30164) );
  XOR U30977 ( .A(n30169), .B(n29911), .Z(n29913) );
  XOR U30978 ( .A(n30170), .B(n30171), .Z(n29911) );
  AND U30979 ( .A(n30172), .B(n30173), .Z(n30170) );
  AND U30980 ( .A(a[4]), .B(b[39]), .Z(n30169) );
  XOR U30981 ( .A(n30174), .B(n29916), .Z(n29918) );
  XOR U30982 ( .A(n30175), .B(n30176), .Z(n29916) );
  AND U30983 ( .A(n30177), .B(n30178), .Z(n30175) );
  AND U30984 ( .A(a[5]), .B(b[38]), .Z(n30174) );
  XOR U30985 ( .A(n30179), .B(n29921), .Z(n29923) );
  XOR U30986 ( .A(n30180), .B(n30181), .Z(n29921) );
  AND U30987 ( .A(n30182), .B(n30183), .Z(n30180) );
  AND U30988 ( .A(a[6]), .B(b[37]), .Z(n30179) );
  XOR U30989 ( .A(n30184), .B(n29926), .Z(n29928) );
  XOR U30990 ( .A(n30185), .B(n30186), .Z(n29926) );
  AND U30991 ( .A(n30187), .B(n30188), .Z(n30185) );
  AND U30992 ( .A(a[7]), .B(b[36]), .Z(n30184) );
  XOR U30993 ( .A(n30189), .B(n29931), .Z(n29933) );
  XOR U30994 ( .A(n30190), .B(n30191), .Z(n29931) );
  AND U30995 ( .A(n30192), .B(n30193), .Z(n30190) );
  AND U30996 ( .A(a[8]), .B(b[35]), .Z(n30189) );
  XOR U30997 ( .A(n30194), .B(n29936), .Z(n29938) );
  XOR U30998 ( .A(n30195), .B(n30196), .Z(n29936) );
  AND U30999 ( .A(n30197), .B(n30198), .Z(n30195) );
  AND U31000 ( .A(a[9]), .B(b[34]), .Z(n30194) );
  XOR U31001 ( .A(n30199), .B(n29941), .Z(n29943) );
  XOR U31002 ( .A(n30200), .B(n30201), .Z(n29941) );
  AND U31003 ( .A(n30202), .B(n30203), .Z(n30200) );
  AND U31004 ( .A(a[10]), .B(b[33]), .Z(n30199) );
  XOR U31005 ( .A(n30204), .B(n29946), .Z(n29948) );
  XOR U31006 ( .A(n30205), .B(n30206), .Z(n29946) );
  AND U31007 ( .A(n30207), .B(n30208), .Z(n30205) );
  AND U31008 ( .A(a[11]), .B(b[32]), .Z(n30204) );
  XOR U31009 ( .A(n30209), .B(n29951), .Z(n29953) );
  XOR U31010 ( .A(n30210), .B(n30211), .Z(n29951) );
  AND U31011 ( .A(n30212), .B(n30213), .Z(n30210) );
  AND U31012 ( .A(a[12]), .B(b[31]), .Z(n30209) );
  XOR U31013 ( .A(n30214), .B(n29956), .Z(n29958) );
  XOR U31014 ( .A(n30215), .B(n30216), .Z(n29956) );
  AND U31015 ( .A(n30217), .B(n30218), .Z(n30215) );
  AND U31016 ( .A(a[13]), .B(b[30]), .Z(n30214) );
  XOR U31017 ( .A(n30219), .B(n29961), .Z(n29963) );
  XOR U31018 ( .A(n30220), .B(n30221), .Z(n29961) );
  AND U31019 ( .A(n30222), .B(n30223), .Z(n30220) );
  AND U31020 ( .A(a[14]), .B(b[29]), .Z(n30219) );
  XOR U31021 ( .A(n30224), .B(n29966), .Z(n29968) );
  XOR U31022 ( .A(n30225), .B(n30226), .Z(n29966) );
  AND U31023 ( .A(n30227), .B(n30228), .Z(n30225) );
  AND U31024 ( .A(a[15]), .B(b[28]), .Z(n30224) );
  XOR U31025 ( .A(n30229), .B(n29971), .Z(n29973) );
  XOR U31026 ( .A(n30230), .B(n30231), .Z(n29971) );
  AND U31027 ( .A(n30232), .B(n30233), .Z(n30230) );
  AND U31028 ( .A(a[16]), .B(b[27]), .Z(n30229) );
  XOR U31029 ( .A(n30234), .B(n29976), .Z(n29978) );
  XOR U31030 ( .A(n30235), .B(n30236), .Z(n29976) );
  AND U31031 ( .A(n30237), .B(n30238), .Z(n30235) );
  AND U31032 ( .A(a[17]), .B(b[26]), .Z(n30234) );
  XOR U31033 ( .A(n30239), .B(n29981), .Z(n29983) );
  XOR U31034 ( .A(n30240), .B(n30241), .Z(n29981) );
  AND U31035 ( .A(n30242), .B(n30243), .Z(n30240) );
  AND U31036 ( .A(a[18]), .B(b[25]), .Z(n30239) );
  XOR U31037 ( .A(n30244), .B(n29986), .Z(n29988) );
  XOR U31038 ( .A(n30245), .B(n30246), .Z(n29986) );
  AND U31039 ( .A(n30247), .B(n30248), .Z(n30245) );
  AND U31040 ( .A(a[19]), .B(b[24]), .Z(n30244) );
  XOR U31041 ( .A(n30249), .B(n29991), .Z(n29993) );
  XOR U31042 ( .A(n30250), .B(n30251), .Z(n29991) );
  AND U31043 ( .A(n30252), .B(n30253), .Z(n30250) );
  AND U31044 ( .A(a[20]), .B(b[23]), .Z(n30249) );
  XOR U31045 ( .A(n30254), .B(n29996), .Z(n29998) );
  XOR U31046 ( .A(n30255), .B(n30256), .Z(n29996) );
  AND U31047 ( .A(n30257), .B(n30258), .Z(n30255) );
  AND U31048 ( .A(a[21]), .B(b[22]), .Z(n30254) );
  XOR U31049 ( .A(n30259), .B(n30001), .Z(n30003) );
  XOR U31050 ( .A(n30260), .B(n30261), .Z(n30001) );
  AND U31051 ( .A(n30262), .B(n30263), .Z(n30260) );
  AND U31052 ( .A(b[21]), .B(a[22]), .Z(n30259) );
  XOR U31053 ( .A(n30264), .B(n30006), .Z(n30008) );
  XOR U31054 ( .A(n30265), .B(n30266), .Z(n30006) );
  AND U31055 ( .A(n30267), .B(n30268), .Z(n30265) );
  AND U31056 ( .A(b[20]), .B(a[23]), .Z(n30264) );
  XOR U31057 ( .A(n30269), .B(n30011), .Z(n30013) );
  XOR U31058 ( .A(n30270), .B(n30271), .Z(n30011) );
  AND U31059 ( .A(n30272), .B(n30273), .Z(n30270) );
  AND U31060 ( .A(b[19]), .B(a[24]), .Z(n30269) );
  XOR U31061 ( .A(n30274), .B(n30016), .Z(n30018) );
  XOR U31062 ( .A(n30275), .B(n30276), .Z(n30016) );
  AND U31063 ( .A(n30277), .B(n30278), .Z(n30275) );
  AND U31064 ( .A(b[18]), .B(a[25]), .Z(n30274) );
  XOR U31065 ( .A(n30279), .B(n30021), .Z(n30023) );
  XOR U31066 ( .A(n30280), .B(n30281), .Z(n30021) );
  AND U31067 ( .A(n30282), .B(n30283), .Z(n30280) );
  AND U31068 ( .A(b[17]), .B(a[26]), .Z(n30279) );
  XOR U31069 ( .A(n30284), .B(n30026), .Z(n30028) );
  XOR U31070 ( .A(n30285), .B(n30286), .Z(n30026) );
  AND U31071 ( .A(n30287), .B(n30288), .Z(n30285) );
  AND U31072 ( .A(b[16]), .B(a[27]), .Z(n30284) );
  XOR U31073 ( .A(n30289), .B(n30031), .Z(n30033) );
  XOR U31074 ( .A(n30290), .B(n30291), .Z(n30031) );
  AND U31075 ( .A(n30292), .B(n30293), .Z(n30290) );
  AND U31076 ( .A(b[15]), .B(a[28]), .Z(n30289) );
  XOR U31077 ( .A(n30294), .B(n30036), .Z(n30038) );
  XOR U31078 ( .A(n30295), .B(n30296), .Z(n30036) );
  AND U31079 ( .A(n30297), .B(n30298), .Z(n30295) );
  AND U31080 ( .A(b[14]), .B(a[29]), .Z(n30294) );
  XOR U31081 ( .A(n30299), .B(n30041), .Z(n30043) );
  XOR U31082 ( .A(n30300), .B(n30301), .Z(n30041) );
  AND U31083 ( .A(n30302), .B(n30303), .Z(n30300) );
  AND U31084 ( .A(b[13]), .B(a[30]), .Z(n30299) );
  XOR U31085 ( .A(n30304), .B(n30046), .Z(n30048) );
  XOR U31086 ( .A(n30305), .B(n30306), .Z(n30046) );
  AND U31087 ( .A(n30307), .B(n30308), .Z(n30305) );
  AND U31088 ( .A(b[12]), .B(a[31]), .Z(n30304) );
  XOR U31089 ( .A(n30309), .B(n30051), .Z(n30053) );
  XOR U31090 ( .A(n30310), .B(n30311), .Z(n30051) );
  AND U31091 ( .A(n30312), .B(n30313), .Z(n30310) );
  AND U31092 ( .A(b[11]), .B(a[32]), .Z(n30309) );
  XOR U31093 ( .A(n30314), .B(n30056), .Z(n30058) );
  XOR U31094 ( .A(n30315), .B(n30316), .Z(n30056) );
  AND U31095 ( .A(n30317), .B(n30318), .Z(n30315) );
  AND U31096 ( .A(b[10]), .B(a[33]), .Z(n30314) );
  XOR U31097 ( .A(n30319), .B(n30061), .Z(n30063) );
  XOR U31098 ( .A(n30320), .B(n30321), .Z(n30061) );
  AND U31099 ( .A(n30322), .B(n30323), .Z(n30320) );
  AND U31100 ( .A(b[9]), .B(a[34]), .Z(n30319) );
  XOR U31101 ( .A(n30324), .B(n30066), .Z(n30068) );
  XOR U31102 ( .A(n30325), .B(n30326), .Z(n30066) );
  AND U31103 ( .A(n30327), .B(n30328), .Z(n30325) );
  AND U31104 ( .A(b[8]), .B(a[35]), .Z(n30324) );
  XOR U31105 ( .A(n30329), .B(n30071), .Z(n30073) );
  XOR U31106 ( .A(n30330), .B(n30331), .Z(n30071) );
  AND U31107 ( .A(n30332), .B(n30333), .Z(n30330) );
  AND U31108 ( .A(b[7]), .B(a[36]), .Z(n30329) );
  XOR U31109 ( .A(n30334), .B(n30076), .Z(n30078) );
  XOR U31110 ( .A(n30335), .B(n30336), .Z(n30076) );
  AND U31111 ( .A(n30337), .B(n30338), .Z(n30335) );
  AND U31112 ( .A(b[6]), .B(a[37]), .Z(n30334) );
  XOR U31113 ( .A(n30339), .B(n30081), .Z(n30083) );
  XOR U31114 ( .A(n30340), .B(n30341), .Z(n30081) );
  AND U31115 ( .A(n30342), .B(n30343), .Z(n30340) );
  AND U31116 ( .A(b[5]), .B(a[38]), .Z(n30339) );
  XOR U31117 ( .A(n30344), .B(n30086), .Z(n30088) );
  XOR U31118 ( .A(n30345), .B(n30346), .Z(n30086) );
  AND U31119 ( .A(n30347), .B(n30348), .Z(n30345) );
  AND U31120 ( .A(b[4]), .B(a[39]), .Z(n30344) );
  XNOR U31121 ( .A(n30349), .B(n30350), .Z(n30100) );
  NANDN U31122 ( .A(n30351), .B(n30352), .Z(n30350) );
  XOR U31123 ( .A(n30353), .B(n30091), .Z(n30093) );
  XNOR U31124 ( .A(n30354), .B(n30355), .Z(n30091) );
  AND U31125 ( .A(n30356), .B(n30357), .Z(n30354) );
  AND U31126 ( .A(b[3]), .B(a[40]), .Z(n30353) );
  XOR U31127 ( .A(n30107), .B(n30106), .Z(c[106]) );
  XOR U31128 ( .A(sreg[170]), .B(n30105), .Z(n30106) );
  XOR U31129 ( .A(n30112), .B(n30358), .Z(n30107) );
  XNOR U31130 ( .A(n30111), .B(n30105), .Z(n30358) );
  XOR U31131 ( .A(n30359), .B(n30360), .Z(n30105) );
  NOR U31132 ( .A(n30361), .B(n30362), .Z(n30359) );
  NAND U31133 ( .A(a[42]), .B(b[0]), .Z(n30111) );
  XNOR U31134 ( .A(n30351), .B(n30352), .Z(n30112) );
  XOR U31135 ( .A(n30349), .B(n30363), .Z(n30352) );
  NAND U31136 ( .A(b[1]), .B(a[41]), .Z(n30363) );
  XOR U31137 ( .A(n30357), .B(n30364), .Z(n30351) );
  XOR U31138 ( .A(n30349), .B(n30356), .Z(n30364) );
  XNOR U31139 ( .A(n30365), .B(n30355), .Z(n30356) );
  AND U31140 ( .A(b[2]), .B(a[40]), .Z(n30365) );
  NANDN U31141 ( .A(n30366), .B(n30367), .Z(n30349) );
  XOR U31142 ( .A(n30355), .B(n30347), .Z(n30368) );
  XNOR U31143 ( .A(n30346), .B(n30342), .Z(n30369) );
  XNOR U31144 ( .A(n30341), .B(n30337), .Z(n30370) );
  XNOR U31145 ( .A(n30336), .B(n30332), .Z(n30371) );
  XNOR U31146 ( .A(n30331), .B(n30327), .Z(n30372) );
  XNOR U31147 ( .A(n30326), .B(n30322), .Z(n30373) );
  XNOR U31148 ( .A(n30321), .B(n30317), .Z(n30374) );
  XNOR U31149 ( .A(n30316), .B(n30312), .Z(n30375) );
  XNOR U31150 ( .A(n30311), .B(n30307), .Z(n30376) );
  XNOR U31151 ( .A(n30306), .B(n30302), .Z(n30377) );
  XNOR U31152 ( .A(n30301), .B(n30297), .Z(n30378) );
  XNOR U31153 ( .A(n30296), .B(n30292), .Z(n30379) );
  XNOR U31154 ( .A(n30291), .B(n30287), .Z(n30380) );
  XNOR U31155 ( .A(n30286), .B(n30282), .Z(n30381) );
  XNOR U31156 ( .A(n30281), .B(n30277), .Z(n30382) );
  XNOR U31157 ( .A(n30276), .B(n30272), .Z(n30383) );
  XNOR U31158 ( .A(n30271), .B(n30267), .Z(n30384) );
  XNOR U31159 ( .A(n30266), .B(n30262), .Z(n30385) );
  XNOR U31160 ( .A(n30261), .B(n30257), .Z(n30386) );
  XNOR U31161 ( .A(n30256), .B(n30252), .Z(n30387) );
  XNOR U31162 ( .A(n30251), .B(n30247), .Z(n30388) );
  XNOR U31163 ( .A(n30246), .B(n30242), .Z(n30389) );
  XNOR U31164 ( .A(n30241), .B(n30237), .Z(n30390) );
  XNOR U31165 ( .A(n30236), .B(n30232), .Z(n30391) );
  XNOR U31166 ( .A(n30231), .B(n30227), .Z(n30392) );
  XNOR U31167 ( .A(n30226), .B(n30222), .Z(n30393) );
  XNOR U31168 ( .A(n30221), .B(n30217), .Z(n30394) );
  XNOR U31169 ( .A(n30216), .B(n30212), .Z(n30395) );
  XNOR U31170 ( .A(n30211), .B(n30207), .Z(n30396) );
  XNOR U31171 ( .A(n30206), .B(n30202), .Z(n30397) );
  XNOR U31172 ( .A(n30201), .B(n30197), .Z(n30398) );
  XNOR U31173 ( .A(n30196), .B(n30192), .Z(n30399) );
  XNOR U31174 ( .A(n30191), .B(n30187), .Z(n30400) );
  XNOR U31175 ( .A(n30186), .B(n30182), .Z(n30401) );
  XNOR U31176 ( .A(n30181), .B(n30177), .Z(n30402) );
  XNOR U31177 ( .A(n30176), .B(n30172), .Z(n30403) );
  XNOR U31178 ( .A(n30171), .B(n30167), .Z(n30404) );
  XNOR U31179 ( .A(n30166), .B(n30162), .Z(n30405) );
  XNOR U31180 ( .A(n30161), .B(n30157), .Z(n30406) );
  XNOR U31181 ( .A(n30407), .B(n30156), .Z(n30157) );
  AND U31182 ( .A(a[0]), .B(b[42]), .Z(n30407) );
  XNOR U31183 ( .A(n30408), .B(n30156), .Z(n30158) );
  XNOR U31184 ( .A(n30409), .B(n30410), .Z(n30156) );
  AND U31185 ( .A(n30411), .B(n30412), .Z(n30409) );
  AND U31186 ( .A(a[1]), .B(b[41]), .Z(n30408) );
  XOR U31187 ( .A(n30413), .B(n30161), .Z(n30163) );
  XOR U31188 ( .A(n30414), .B(n30415), .Z(n30161) );
  AND U31189 ( .A(n30416), .B(n30417), .Z(n30414) );
  AND U31190 ( .A(a[2]), .B(b[40]), .Z(n30413) );
  XOR U31191 ( .A(n30418), .B(n30166), .Z(n30168) );
  XOR U31192 ( .A(n30419), .B(n30420), .Z(n30166) );
  AND U31193 ( .A(n30421), .B(n30422), .Z(n30419) );
  AND U31194 ( .A(a[3]), .B(b[39]), .Z(n30418) );
  XOR U31195 ( .A(n30423), .B(n30171), .Z(n30173) );
  XOR U31196 ( .A(n30424), .B(n30425), .Z(n30171) );
  AND U31197 ( .A(n30426), .B(n30427), .Z(n30424) );
  AND U31198 ( .A(a[4]), .B(b[38]), .Z(n30423) );
  XOR U31199 ( .A(n30428), .B(n30176), .Z(n30178) );
  XOR U31200 ( .A(n30429), .B(n30430), .Z(n30176) );
  AND U31201 ( .A(n30431), .B(n30432), .Z(n30429) );
  AND U31202 ( .A(a[5]), .B(b[37]), .Z(n30428) );
  XOR U31203 ( .A(n30433), .B(n30181), .Z(n30183) );
  XOR U31204 ( .A(n30434), .B(n30435), .Z(n30181) );
  AND U31205 ( .A(n30436), .B(n30437), .Z(n30434) );
  AND U31206 ( .A(a[6]), .B(b[36]), .Z(n30433) );
  XOR U31207 ( .A(n30438), .B(n30186), .Z(n30188) );
  XOR U31208 ( .A(n30439), .B(n30440), .Z(n30186) );
  AND U31209 ( .A(n30441), .B(n30442), .Z(n30439) );
  AND U31210 ( .A(a[7]), .B(b[35]), .Z(n30438) );
  XOR U31211 ( .A(n30443), .B(n30191), .Z(n30193) );
  XOR U31212 ( .A(n30444), .B(n30445), .Z(n30191) );
  AND U31213 ( .A(n30446), .B(n30447), .Z(n30444) );
  AND U31214 ( .A(a[8]), .B(b[34]), .Z(n30443) );
  XOR U31215 ( .A(n30448), .B(n30196), .Z(n30198) );
  XOR U31216 ( .A(n30449), .B(n30450), .Z(n30196) );
  AND U31217 ( .A(n30451), .B(n30452), .Z(n30449) );
  AND U31218 ( .A(a[9]), .B(b[33]), .Z(n30448) );
  XOR U31219 ( .A(n30453), .B(n30201), .Z(n30203) );
  XOR U31220 ( .A(n30454), .B(n30455), .Z(n30201) );
  AND U31221 ( .A(n30456), .B(n30457), .Z(n30454) );
  AND U31222 ( .A(a[10]), .B(b[32]), .Z(n30453) );
  XOR U31223 ( .A(n30458), .B(n30206), .Z(n30208) );
  XOR U31224 ( .A(n30459), .B(n30460), .Z(n30206) );
  AND U31225 ( .A(n30461), .B(n30462), .Z(n30459) );
  AND U31226 ( .A(a[11]), .B(b[31]), .Z(n30458) );
  XOR U31227 ( .A(n30463), .B(n30211), .Z(n30213) );
  XOR U31228 ( .A(n30464), .B(n30465), .Z(n30211) );
  AND U31229 ( .A(n30466), .B(n30467), .Z(n30464) );
  AND U31230 ( .A(a[12]), .B(b[30]), .Z(n30463) );
  XOR U31231 ( .A(n30468), .B(n30216), .Z(n30218) );
  XOR U31232 ( .A(n30469), .B(n30470), .Z(n30216) );
  AND U31233 ( .A(n30471), .B(n30472), .Z(n30469) );
  AND U31234 ( .A(a[13]), .B(b[29]), .Z(n30468) );
  XOR U31235 ( .A(n30473), .B(n30221), .Z(n30223) );
  XOR U31236 ( .A(n30474), .B(n30475), .Z(n30221) );
  AND U31237 ( .A(n30476), .B(n30477), .Z(n30474) );
  AND U31238 ( .A(a[14]), .B(b[28]), .Z(n30473) );
  XOR U31239 ( .A(n30478), .B(n30226), .Z(n30228) );
  XOR U31240 ( .A(n30479), .B(n30480), .Z(n30226) );
  AND U31241 ( .A(n30481), .B(n30482), .Z(n30479) );
  AND U31242 ( .A(a[15]), .B(b[27]), .Z(n30478) );
  XOR U31243 ( .A(n30483), .B(n30231), .Z(n30233) );
  XOR U31244 ( .A(n30484), .B(n30485), .Z(n30231) );
  AND U31245 ( .A(n30486), .B(n30487), .Z(n30484) );
  AND U31246 ( .A(a[16]), .B(b[26]), .Z(n30483) );
  XOR U31247 ( .A(n30488), .B(n30236), .Z(n30238) );
  XOR U31248 ( .A(n30489), .B(n30490), .Z(n30236) );
  AND U31249 ( .A(n30491), .B(n30492), .Z(n30489) );
  AND U31250 ( .A(a[17]), .B(b[25]), .Z(n30488) );
  XOR U31251 ( .A(n30493), .B(n30241), .Z(n30243) );
  XOR U31252 ( .A(n30494), .B(n30495), .Z(n30241) );
  AND U31253 ( .A(n30496), .B(n30497), .Z(n30494) );
  AND U31254 ( .A(a[18]), .B(b[24]), .Z(n30493) );
  XOR U31255 ( .A(n30498), .B(n30246), .Z(n30248) );
  XOR U31256 ( .A(n30499), .B(n30500), .Z(n30246) );
  AND U31257 ( .A(n30501), .B(n30502), .Z(n30499) );
  AND U31258 ( .A(a[19]), .B(b[23]), .Z(n30498) );
  XOR U31259 ( .A(n30503), .B(n30251), .Z(n30253) );
  XOR U31260 ( .A(n30504), .B(n30505), .Z(n30251) );
  AND U31261 ( .A(n30506), .B(n30507), .Z(n30504) );
  AND U31262 ( .A(a[20]), .B(b[22]), .Z(n30503) );
  XOR U31263 ( .A(n30508), .B(n30256), .Z(n30258) );
  XOR U31264 ( .A(n30509), .B(n30510), .Z(n30256) );
  AND U31265 ( .A(n30511), .B(n30512), .Z(n30509) );
  AND U31266 ( .A(a[21]), .B(b[21]), .Z(n30508) );
  XOR U31267 ( .A(n30513), .B(n30261), .Z(n30263) );
  XOR U31268 ( .A(n30514), .B(n30515), .Z(n30261) );
  AND U31269 ( .A(n30516), .B(n30517), .Z(n30514) );
  AND U31270 ( .A(b[20]), .B(a[22]), .Z(n30513) );
  XOR U31271 ( .A(n30518), .B(n30266), .Z(n30268) );
  XOR U31272 ( .A(n30519), .B(n30520), .Z(n30266) );
  AND U31273 ( .A(n30521), .B(n30522), .Z(n30519) );
  AND U31274 ( .A(b[19]), .B(a[23]), .Z(n30518) );
  XOR U31275 ( .A(n30523), .B(n30271), .Z(n30273) );
  XOR U31276 ( .A(n30524), .B(n30525), .Z(n30271) );
  AND U31277 ( .A(n30526), .B(n30527), .Z(n30524) );
  AND U31278 ( .A(b[18]), .B(a[24]), .Z(n30523) );
  XOR U31279 ( .A(n30528), .B(n30276), .Z(n30278) );
  XOR U31280 ( .A(n30529), .B(n30530), .Z(n30276) );
  AND U31281 ( .A(n30531), .B(n30532), .Z(n30529) );
  AND U31282 ( .A(b[17]), .B(a[25]), .Z(n30528) );
  XOR U31283 ( .A(n30533), .B(n30281), .Z(n30283) );
  XOR U31284 ( .A(n30534), .B(n30535), .Z(n30281) );
  AND U31285 ( .A(n30536), .B(n30537), .Z(n30534) );
  AND U31286 ( .A(b[16]), .B(a[26]), .Z(n30533) );
  XOR U31287 ( .A(n30538), .B(n30286), .Z(n30288) );
  XOR U31288 ( .A(n30539), .B(n30540), .Z(n30286) );
  AND U31289 ( .A(n30541), .B(n30542), .Z(n30539) );
  AND U31290 ( .A(b[15]), .B(a[27]), .Z(n30538) );
  XOR U31291 ( .A(n30543), .B(n30291), .Z(n30293) );
  XOR U31292 ( .A(n30544), .B(n30545), .Z(n30291) );
  AND U31293 ( .A(n30546), .B(n30547), .Z(n30544) );
  AND U31294 ( .A(b[14]), .B(a[28]), .Z(n30543) );
  XOR U31295 ( .A(n30548), .B(n30296), .Z(n30298) );
  XOR U31296 ( .A(n30549), .B(n30550), .Z(n30296) );
  AND U31297 ( .A(n30551), .B(n30552), .Z(n30549) );
  AND U31298 ( .A(b[13]), .B(a[29]), .Z(n30548) );
  XOR U31299 ( .A(n30553), .B(n30301), .Z(n30303) );
  XOR U31300 ( .A(n30554), .B(n30555), .Z(n30301) );
  AND U31301 ( .A(n30556), .B(n30557), .Z(n30554) );
  AND U31302 ( .A(b[12]), .B(a[30]), .Z(n30553) );
  XOR U31303 ( .A(n30558), .B(n30306), .Z(n30308) );
  XOR U31304 ( .A(n30559), .B(n30560), .Z(n30306) );
  AND U31305 ( .A(n30561), .B(n30562), .Z(n30559) );
  AND U31306 ( .A(b[11]), .B(a[31]), .Z(n30558) );
  XOR U31307 ( .A(n30563), .B(n30311), .Z(n30313) );
  XOR U31308 ( .A(n30564), .B(n30565), .Z(n30311) );
  AND U31309 ( .A(n30566), .B(n30567), .Z(n30564) );
  AND U31310 ( .A(b[10]), .B(a[32]), .Z(n30563) );
  XOR U31311 ( .A(n30568), .B(n30316), .Z(n30318) );
  XOR U31312 ( .A(n30569), .B(n30570), .Z(n30316) );
  AND U31313 ( .A(n30571), .B(n30572), .Z(n30569) );
  AND U31314 ( .A(b[9]), .B(a[33]), .Z(n30568) );
  XOR U31315 ( .A(n30573), .B(n30321), .Z(n30323) );
  XOR U31316 ( .A(n30574), .B(n30575), .Z(n30321) );
  AND U31317 ( .A(n30576), .B(n30577), .Z(n30574) );
  AND U31318 ( .A(b[8]), .B(a[34]), .Z(n30573) );
  XOR U31319 ( .A(n30578), .B(n30326), .Z(n30328) );
  XOR U31320 ( .A(n30579), .B(n30580), .Z(n30326) );
  AND U31321 ( .A(n30581), .B(n30582), .Z(n30579) );
  AND U31322 ( .A(b[7]), .B(a[35]), .Z(n30578) );
  XOR U31323 ( .A(n30583), .B(n30331), .Z(n30333) );
  XOR U31324 ( .A(n30584), .B(n30585), .Z(n30331) );
  AND U31325 ( .A(n30586), .B(n30587), .Z(n30584) );
  AND U31326 ( .A(b[6]), .B(a[36]), .Z(n30583) );
  XOR U31327 ( .A(n30588), .B(n30336), .Z(n30338) );
  XOR U31328 ( .A(n30589), .B(n30590), .Z(n30336) );
  AND U31329 ( .A(n30591), .B(n30592), .Z(n30589) );
  AND U31330 ( .A(b[5]), .B(a[37]), .Z(n30588) );
  XOR U31331 ( .A(n30593), .B(n30341), .Z(n30343) );
  XOR U31332 ( .A(n30594), .B(n30595), .Z(n30341) );
  AND U31333 ( .A(n30596), .B(n30597), .Z(n30594) );
  AND U31334 ( .A(b[4]), .B(a[38]), .Z(n30593) );
  XNOR U31335 ( .A(n30598), .B(n30599), .Z(n30355) );
  NANDN U31336 ( .A(n30600), .B(n30601), .Z(n30599) );
  XOR U31337 ( .A(n30602), .B(n30346), .Z(n30348) );
  XNOR U31338 ( .A(n30603), .B(n30604), .Z(n30346) );
  AND U31339 ( .A(n30605), .B(n30606), .Z(n30603) );
  AND U31340 ( .A(b[3]), .B(a[39]), .Z(n30602) );
  XOR U31341 ( .A(n30362), .B(n30361), .Z(c[105]) );
  XOR U31342 ( .A(sreg[169]), .B(n30360), .Z(n30361) );
  XOR U31343 ( .A(n30367), .B(n30607), .Z(n30362) );
  XNOR U31344 ( .A(n30366), .B(n30360), .Z(n30607) );
  XOR U31345 ( .A(n30608), .B(n30609), .Z(n30360) );
  NOR U31346 ( .A(n30610), .B(n30611), .Z(n30608) );
  NAND U31347 ( .A(a[41]), .B(b[0]), .Z(n30366) );
  XNOR U31348 ( .A(n30600), .B(n30601), .Z(n30367) );
  XOR U31349 ( .A(n30598), .B(n30612), .Z(n30601) );
  NAND U31350 ( .A(b[1]), .B(a[40]), .Z(n30612) );
  XOR U31351 ( .A(n30606), .B(n30613), .Z(n30600) );
  XOR U31352 ( .A(n30598), .B(n30605), .Z(n30613) );
  XNOR U31353 ( .A(n30614), .B(n30604), .Z(n30605) );
  AND U31354 ( .A(b[2]), .B(a[39]), .Z(n30614) );
  NANDN U31355 ( .A(n30615), .B(n30616), .Z(n30598) );
  XOR U31356 ( .A(n30604), .B(n30596), .Z(n30617) );
  XNOR U31357 ( .A(n30595), .B(n30591), .Z(n30618) );
  XNOR U31358 ( .A(n30590), .B(n30586), .Z(n30619) );
  XNOR U31359 ( .A(n30585), .B(n30581), .Z(n30620) );
  XNOR U31360 ( .A(n30580), .B(n30576), .Z(n30621) );
  XNOR U31361 ( .A(n30575), .B(n30571), .Z(n30622) );
  XNOR U31362 ( .A(n30570), .B(n30566), .Z(n30623) );
  XNOR U31363 ( .A(n30565), .B(n30561), .Z(n30624) );
  XNOR U31364 ( .A(n30560), .B(n30556), .Z(n30625) );
  XNOR U31365 ( .A(n30555), .B(n30551), .Z(n30626) );
  XNOR U31366 ( .A(n30550), .B(n30546), .Z(n30627) );
  XNOR U31367 ( .A(n30545), .B(n30541), .Z(n30628) );
  XNOR U31368 ( .A(n30540), .B(n30536), .Z(n30629) );
  XNOR U31369 ( .A(n30535), .B(n30531), .Z(n30630) );
  XNOR U31370 ( .A(n30530), .B(n30526), .Z(n30631) );
  XNOR U31371 ( .A(n30525), .B(n30521), .Z(n30632) );
  XNOR U31372 ( .A(n30520), .B(n30516), .Z(n30633) );
  XNOR U31373 ( .A(n30515), .B(n30511), .Z(n30634) );
  XNOR U31374 ( .A(n30510), .B(n30506), .Z(n30635) );
  XNOR U31375 ( .A(n30505), .B(n30501), .Z(n30636) );
  XNOR U31376 ( .A(n30500), .B(n30496), .Z(n30637) );
  XNOR U31377 ( .A(n30495), .B(n30491), .Z(n30638) );
  XNOR U31378 ( .A(n30490), .B(n30486), .Z(n30639) );
  XNOR U31379 ( .A(n30485), .B(n30481), .Z(n30640) );
  XNOR U31380 ( .A(n30480), .B(n30476), .Z(n30641) );
  XNOR U31381 ( .A(n30475), .B(n30471), .Z(n30642) );
  XNOR U31382 ( .A(n30470), .B(n30466), .Z(n30643) );
  XNOR U31383 ( .A(n30465), .B(n30461), .Z(n30644) );
  XNOR U31384 ( .A(n30460), .B(n30456), .Z(n30645) );
  XNOR U31385 ( .A(n30455), .B(n30451), .Z(n30646) );
  XNOR U31386 ( .A(n30450), .B(n30446), .Z(n30647) );
  XNOR U31387 ( .A(n30445), .B(n30441), .Z(n30648) );
  XNOR U31388 ( .A(n30440), .B(n30436), .Z(n30649) );
  XNOR U31389 ( .A(n30435), .B(n30431), .Z(n30650) );
  XNOR U31390 ( .A(n30430), .B(n30426), .Z(n30651) );
  XNOR U31391 ( .A(n30425), .B(n30421), .Z(n30652) );
  XNOR U31392 ( .A(n30420), .B(n30416), .Z(n30653) );
  XNOR U31393 ( .A(n30415), .B(n30411), .Z(n30654) );
  XOR U31394 ( .A(n30655), .B(n30410), .Z(n30411) );
  AND U31395 ( .A(a[0]), .B(b[41]), .Z(n30655) );
  XOR U31396 ( .A(n30656), .B(n30410), .Z(n30412) );
  XNOR U31397 ( .A(n30657), .B(n30658), .Z(n30410) );
  AND U31398 ( .A(n30659), .B(n30660), .Z(n30657) );
  AND U31399 ( .A(a[1]), .B(b[40]), .Z(n30656) );
  XOR U31400 ( .A(n30661), .B(n30415), .Z(n30417) );
  XOR U31401 ( .A(n30662), .B(n30663), .Z(n30415) );
  AND U31402 ( .A(n30664), .B(n30665), .Z(n30662) );
  AND U31403 ( .A(a[2]), .B(b[39]), .Z(n30661) );
  XOR U31404 ( .A(n30666), .B(n30420), .Z(n30422) );
  XOR U31405 ( .A(n30667), .B(n30668), .Z(n30420) );
  AND U31406 ( .A(n30669), .B(n30670), .Z(n30667) );
  AND U31407 ( .A(a[3]), .B(b[38]), .Z(n30666) );
  XOR U31408 ( .A(n30671), .B(n30425), .Z(n30427) );
  XOR U31409 ( .A(n30672), .B(n30673), .Z(n30425) );
  AND U31410 ( .A(n30674), .B(n30675), .Z(n30672) );
  AND U31411 ( .A(a[4]), .B(b[37]), .Z(n30671) );
  XOR U31412 ( .A(n30676), .B(n30430), .Z(n30432) );
  XOR U31413 ( .A(n30677), .B(n30678), .Z(n30430) );
  AND U31414 ( .A(n30679), .B(n30680), .Z(n30677) );
  AND U31415 ( .A(a[5]), .B(b[36]), .Z(n30676) );
  XOR U31416 ( .A(n30681), .B(n30435), .Z(n30437) );
  XOR U31417 ( .A(n30682), .B(n30683), .Z(n30435) );
  AND U31418 ( .A(n30684), .B(n30685), .Z(n30682) );
  AND U31419 ( .A(a[6]), .B(b[35]), .Z(n30681) );
  XOR U31420 ( .A(n30686), .B(n30440), .Z(n30442) );
  XOR U31421 ( .A(n30687), .B(n30688), .Z(n30440) );
  AND U31422 ( .A(n30689), .B(n30690), .Z(n30687) );
  AND U31423 ( .A(a[7]), .B(b[34]), .Z(n30686) );
  XOR U31424 ( .A(n30691), .B(n30445), .Z(n30447) );
  XOR U31425 ( .A(n30692), .B(n30693), .Z(n30445) );
  AND U31426 ( .A(n30694), .B(n30695), .Z(n30692) );
  AND U31427 ( .A(a[8]), .B(b[33]), .Z(n30691) );
  XOR U31428 ( .A(n30696), .B(n30450), .Z(n30452) );
  XOR U31429 ( .A(n30697), .B(n30698), .Z(n30450) );
  AND U31430 ( .A(n30699), .B(n30700), .Z(n30697) );
  AND U31431 ( .A(a[9]), .B(b[32]), .Z(n30696) );
  XOR U31432 ( .A(n30701), .B(n30455), .Z(n30457) );
  XOR U31433 ( .A(n30702), .B(n30703), .Z(n30455) );
  AND U31434 ( .A(n30704), .B(n30705), .Z(n30702) );
  AND U31435 ( .A(a[10]), .B(b[31]), .Z(n30701) );
  XOR U31436 ( .A(n30706), .B(n30460), .Z(n30462) );
  XOR U31437 ( .A(n30707), .B(n30708), .Z(n30460) );
  AND U31438 ( .A(n30709), .B(n30710), .Z(n30707) );
  AND U31439 ( .A(a[11]), .B(b[30]), .Z(n30706) );
  XOR U31440 ( .A(n30711), .B(n30465), .Z(n30467) );
  XOR U31441 ( .A(n30712), .B(n30713), .Z(n30465) );
  AND U31442 ( .A(n30714), .B(n30715), .Z(n30712) );
  AND U31443 ( .A(a[12]), .B(b[29]), .Z(n30711) );
  XOR U31444 ( .A(n30716), .B(n30470), .Z(n30472) );
  XOR U31445 ( .A(n30717), .B(n30718), .Z(n30470) );
  AND U31446 ( .A(n30719), .B(n30720), .Z(n30717) );
  AND U31447 ( .A(a[13]), .B(b[28]), .Z(n30716) );
  XOR U31448 ( .A(n30721), .B(n30475), .Z(n30477) );
  XOR U31449 ( .A(n30722), .B(n30723), .Z(n30475) );
  AND U31450 ( .A(n30724), .B(n30725), .Z(n30722) );
  AND U31451 ( .A(a[14]), .B(b[27]), .Z(n30721) );
  XOR U31452 ( .A(n30726), .B(n30480), .Z(n30482) );
  XOR U31453 ( .A(n30727), .B(n30728), .Z(n30480) );
  AND U31454 ( .A(n30729), .B(n30730), .Z(n30727) );
  AND U31455 ( .A(a[15]), .B(b[26]), .Z(n30726) );
  XOR U31456 ( .A(n30731), .B(n30485), .Z(n30487) );
  XOR U31457 ( .A(n30732), .B(n30733), .Z(n30485) );
  AND U31458 ( .A(n30734), .B(n30735), .Z(n30732) );
  AND U31459 ( .A(a[16]), .B(b[25]), .Z(n30731) );
  XOR U31460 ( .A(n30736), .B(n30490), .Z(n30492) );
  XOR U31461 ( .A(n30737), .B(n30738), .Z(n30490) );
  AND U31462 ( .A(n30739), .B(n30740), .Z(n30737) );
  AND U31463 ( .A(a[17]), .B(b[24]), .Z(n30736) );
  XOR U31464 ( .A(n30741), .B(n30495), .Z(n30497) );
  XOR U31465 ( .A(n30742), .B(n30743), .Z(n30495) );
  AND U31466 ( .A(n30744), .B(n30745), .Z(n30742) );
  AND U31467 ( .A(a[18]), .B(b[23]), .Z(n30741) );
  XOR U31468 ( .A(n30746), .B(n30500), .Z(n30502) );
  XOR U31469 ( .A(n30747), .B(n30748), .Z(n30500) );
  AND U31470 ( .A(n30749), .B(n30750), .Z(n30747) );
  AND U31471 ( .A(a[19]), .B(b[22]), .Z(n30746) );
  XOR U31472 ( .A(n30751), .B(n30505), .Z(n30507) );
  XOR U31473 ( .A(n30752), .B(n30753), .Z(n30505) );
  AND U31474 ( .A(n30754), .B(n30755), .Z(n30752) );
  AND U31475 ( .A(a[20]), .B(b[21]), .Z(n30751) );
  XOR U31476 ( .A(n30756), .B(n30510), .Z(n30512) );
  XOR U31477 ( .A(n30757), .B(n30758), .Z(n30510) );
  AND U31478 ( .A(n30759), .B(n30760), .Z(n30757) );
  AND U31479 ( .A(b[20]), .B(a[21]), .Z(n30756) );
  XOR U31480 ( .A(n30761), .B(n30515), .Z(n30517) );
  XOR U31481 ( .A(n30762), .B(n30763), .Z(n30515) );
  AND U31482 ( .A(n30764), .B(n30765), .Z(n30762) );
  AND U31483 ( .A(b[19]), .B(a[22]), .Z(n30761) );
  XOR U31484 ( .A(n30766), .B(n30520), .Z(n30522) );
  XOR U31485 ( .A(n30767), .B(n30768), .Z(n30520) );
  AND U31486 ( .A(n30769), .B(n30770), .Z(n30767) );
  AND U31487 ( .A(b[18]), .B(a[23]), .Z(n30766) );
  XOR U31488 ( .A(n30771), .B(n30525), .Z(n30527) );
  XOR U31489 ( .A(n30772), .B(n30773), .Z(n30525) );
  AND U31490 ( .A(n30774), .B(n30775), .Z(n30772) );
  AND U31491 ( .A(b[17]), .B(a[24]), .Z(n30771) );
  XOR U31492 ( .A(n30776), .B(n30530), .Z(n30532) );
  XOR U31493 ( .A(n30777), .B(n30778), .Z(n30530) );
  AND U31494 ( .A(n30779), .B(n30780), .Z(n30777) );
  AND U31495 ( .A(b[16]), .B(a[25]), .Z(n30776) );
  XOR U31496 ( .A(n30781), .B(n30535), .Z(n30537) );
  XOR U31497 ( .A(n30782), .B(n30783), .Z(n30535) );
  AND U31498 ( .A(n30784), .B(n30785), .Z(n30782) );
  AND U31499 ( .A(b[15]), .B(a[26]), .Z(n30781) );
  XOR U31500 ( .A(n30786), .B(n30540), .Z(n30542) );
  XOR U31501 ( .A(n30787), .B(n30788), .Z(n30540) );
  AND U31502 ( .A(n30789), .B(n30790), .Z(n30787) );
  AND U31503 ( .A(b[14]), .B(a[27]), .Z(n30786) );
  XOR U31504 ( .A(n30791), .B(n30545), .Z(n30547) );
  XOR U31505 ( .A(n30792), .B(n30793), .Z(n30545) );
  AND U31506 ( .A(n30794), .B(n30795), .Z(n30792) );
  AND U31507 ( .A(b[13]), .B(a[28]), .Z(n30791) );
  XOR U31508 ( .A(n30796), .B(n30550), .Z(n30552) );
  XOR U31509 ( .A(n30797), .B(n30798), .Z(n30550) );
  AND U31510 ( .A(n30799), .B(n30800), .Z(n30797) );
  AND U31511 ( .A(b[12]), .B(a[29]), .Z(n30796) );
  XOR U31512 ( .A(n30801), .B(n30555), .Z(n30557) );
  XOR U31513 ( .A(n30802), .B(n30803), .Z(n30555) );
  AND U31514 ( .A(n30804), .B(n30805), .Z(n30802) );
  AND U31515 ( .A(b[11]), .B(a[30]), .Z(n30801) );
  XOR U31516 ( .A(n30806), .B(n30560), .Z(n30562) );
  XOR U31517 ( .A(n30807), .B(n30808), .Z(n30560) );
  AND U31518 ( .A(n30809), .B(n30810), .Z(n30807) );
  AND U31519 ( .A(b[10]), .B(a[31]), .Z(n30806) );
  XOR U31520 ( .A(n30811), .B(n30565), .Z(n30567) );
  XOR U31521 ( .A(n30812), .B(n30813), .Z(n30565) );
  AND U31522 ( .A(n30814), .B(n30815), .Z(n30812) );
  AND U31523 ( .A(b[9]), .B(a[32]), .Z(n30811) );
  XOR U31524 ( .A(n30816), .B(n30570), .Z(n30572) );
  XOR U31525 ( .A(n30817), .B(n30818), .Z(n30570) );
  AND U31526 ( .A(n30819), .B(n30820), .Z(n30817) );
  AND U31527 ( .A(b[8]), .B(a[33]), .Z(n30816) );
  XOR U31528 ( .A(n30821), .B(n30575), .Z(n30577) );
  XOR U31529 ( .A(n30822), .B(n30823), .Z(n30575) );
  AND U31530 ( .A(n30824), .B(n30825), .Z(n30822) );
  AND U31531 ( .A(b[7]), .B(a[34]), .Z(n30821) );
  XOR U31532 ( .A(n30826), .B(n30580), .Z(n30582) );
  XOR U31533 ( .A(n30827), .B(n30828), .Z(n30580) );
  AND U31534 ( .A(n30829), .B(n30830), .Z(n30827) );
  AND U31535 ( .A(b[6]), .B(a[35]), .Z(n30826) );
  XOR U31536 ( .A(n30831), .B(n30585), .Z(n30587) );
  XOR U31537 ( .A(n30832), .B(n30833), .Z(n30585) );
  AND U31538 ( .A(n30834), .B(n30835), .Z(n30832) );
  AND U31539 ( .A(b[5]), .B(a[36]), .Z(n30831) );
  XOR U31540 ( .A(n30836), .B(n30590), .Z(n30592) );
  XOR U31541 ( .A(n30837), .B(n30838), .Z(n30590) );
  AND U31542 ( .A(n30839), .B(n30840), .Z(n30837) );
  AND U31543 ( .A(b[4]), .B(a[37]), .Z(n30836) );
  XNOR U31544 ( .A(n30841), .B(n30842), .Z(n30604) );
  NANDN U31545 ( .A(n30843), .B(n30844), .Z(n30842) );
  XOR U31546 ( .A(n30845), .B(n30595), .Z(n30597) );
  XNOR U31547 ( .A(n30846), .B(n30847), .Z(n30595) );
  AND U31548 ( .A(n30848), .B(n30849), .Z(n30846) );
  AND U31549 ( .A(b[3]), .B(a[38]), .Z(n30845) );
  XOR U31550 ( .A(n30611), .B(n30610), .Z(c[104]) );
  XOR U31551 ( .A(sreg[168]), .B(n30609), .Z(n30610) );
  XOR U31552 ( .A(n30616), .B(n30850), .Z(n30611) );
  XNOR U31553 ( .A(n30615), .B(n30609), .Z(n30850) );
  XOR U31554 ( .A(n30851), .B(n30852), .Z(n30609) );
  NOR U31555 ( .A(n30853), .B(n30854), .Z(n30851) );
  NAND U31556 ( .A(a[40]), .B(b[0]), .Z(n30615) );
  XNOR U31557 ( .A(n30843), .B(n30844), .Z(n30616) );
  XOR U31558 ( .A(n30841), .B(n30855), .Z(n30844) );
  NAND U31559 ( .A(b[1]), .B(a[39]), .Z(n30855) );
  XOR U31560 ( .A(n30849), .B(n30856), .Z(n30843) );
  XOR U31561 ( .A(n30841), .B(n30848), .Z(n30856) );
  XNOR U31562 ( .A(n30857), .B(n30847), .Z(n30848) );
  AND U31563 ( .A(b[2]), .B(a[38]), .Z(n30857) );
  NANDN U31564 ( .A(n30858), .B(n30859), .Z(n30841) );
  XOR U31565 ( .A(n30847), .B(n30839), .Z(n30860) );
  XNOR U31566 ( .A(n30838), .B(n30834), .Z(n30861) );
  XNOR U31567 ( .A(n30833), .B(n30829), .Z(n30862) );
  XNOR U31568 ( .A(n30828), .B(n30824), .Z(n30863) );
  XNOR U31569 ( .A(n30823), .B(n30819), .Z(n30864) );
  XNOR U31570 ( .A(n30818), .B(n30814), .Z(n30865) );
  XNOR U31571 ( .A(n30813), .B(n30809), .Z(n30866) );
  XNOR U31572 ( .A(n30808), .B(n30804), .Z(n30867) );
  XNOR U31573 ( .A(n30803), .B(n30799), .Z(n30868) );
  XNOR U31574 ( .A(n30798), .B(n30794), .Z(n30869) );
  XNOR U31575 ( .A(n30793), .B(n30789), .Z(n30870) );
  XNOR U31576 ( .A(n30788), .B(n30784), .Z(n30871) );
  XNOR U31577 ( .A(n30783), .B(n30779), .Z(n30872) );
  XNOR U31578 ( .A(n30778), .B(n30774), .Z(n30873) );
  XNOR U31579 ( .A(n30773), .B(n30769), .Z(n30874) );
  XNOR U31580 ( .A(n30768), .B(n30764), .Z(n30875) );
  XNOR U31581 ( .A(n30763), .B(n30759), .Z(n30876) );
  XNOR U31582 ( .A(n30758), .B(n30754), .Z(n30877) );
  XNOR U31583 ( .A(n30753), .B(n30749), .Z(n30878) );
  XNOR U31584 ( .A(n30748), .B(n30744), .Z(n30879) );
  XNOR U31585 ( .A(n30743), .B(n30739), .Z(n30880) );
  XNOR U31586 ( .A(n30738), .B(n30734), .Z(n30881) );
  XNOR U31587 ( .A(n30733), .B(n30729), .Z(n30882) );
  XNOR U31588 ( .A(n30728), .B(n30724), .Z(n30883) );
  XNOR U31589 ( .A(n30723), .B(n30719), .Z(n30884) );
  XNOR U31590 ( .A(n30718), .B(n30714), .Z(n30885) );
  XNOR U31591 ( .A(n30713), .B(n30709), .Z(n30886) );
  XNOR U31592 ( .A(n30708), .B(n30704), .Z(n30887) );
  XNOR U31593 ( .A(n30703), .B(n30699), .Z(n30888) );
  XNOR U31594 ( .A(n30698), .B(n30694), .Z(n30889) );
  XNOR U31595 ( .A(n30693), .B(n30689), .Z(n30890) );
  XNOR U31596 ( .A(n30688), .B(n30684), .Z(n30891) );
  XNOR U31597 ( .A(n30683), .B(n30679), .Z(n30892) );
  XNOR U31598 ( .A(n30678), .B(n30674), .Z(n30893) );
  XNOR U31599 ( .A(n30673), .B(n30669), .Z(n30894) );
  XNOR U31600 ( .A(n30668), .B(n30664), .Z(n30895) );
  XNOR U31601 ( .A(n30663), .B(n30659), .Z(n30896) );
  XNOR U31602 ( .A(n30897), .B(n30658), .Z(n30659) );
  AND U31603 ( .A(a[0]), .B(b[40]), .Z(n30897) );
  XNOR U31604 ( .A(n30898), .B(n30658), .Z(n30660) );
  XNOR U31605 ( .A(n30899), .B(n30900), .Z(n30658) );
  AND U31606 ( .A(n30901), .B(n30902), .Z(n30899) );
  AND U31607 ( .A(a[1]), .B(b[39]), .Z(n30898) );
  XOR U31608 ( .A(n30903), .B(n30663), .Z(n30665) );
  XOR U31609 ( .A(n30904), .B(n30905), .Z(n30663) );
  AND U31610 ( .A(n30906), .B(n30907), .Z(n30904) );
  AND U31611 ( .A(a[2]), .B(b[38]), .Z(n30903) );
  XOR U31612 ( .A(n30908), .B(n30668), .Z(n30670) );
  XOR U31613 ( .A(n30909), .B(n30910), .Z(n30668) );
  AND U31614 ( .A(n30911), .B(n30912), .Z(n30909) );
  AND U31615 ( .A(a[3]), .B(b[37]), .Z(n30908) );
  XOR U31616 ( .A(n30913), .B(n30673), .Z(n30675) );
  XOR U31617 ( .A(n30914), .B(n30915), .Z(n30673) );
  AND U31618 ( .A(n30916), .B(n30917), .Z(n30914) );
  AND U31619 ( .A(a[4]), .B(b[36]), .Z(n30913) );
  XOR U31620 ( .A(n30918), .B(n30678), .Z(n30680) );
  XOR U31621 ( .A(n30919), .B(n30920), .Z(n30678) );
  AND U31622 ( .A(n30921), .B(n30922), .Z(n30919) );
  AND U31623 ( .A(a[5]), .B(b[35]), .Z(n30918) );
  XOR U31624 ( .A(n30923), .B(n30683), .Z(n30685) );
  XOR U31625 ( .A(n30924), .B(n30925), .Z(n30683) );
  AND U31626 ( .A(n30926), .B(n30927), .Z(n30924) );
  AND U31627 ( .A(a[6]), .B(b[34]), .Z(n30923) );
  XOR U31628 ( .A(n30928), .B(n30688), .Z(n30690) );
  XOR U31629 ( .A(n30929), .B(n30930), .Z(n30688) );
  AND U31630 ( .A(n30931), .B(n30932), .Z(n30929) );
  AND U31631 ( .A(a[7]), .B(b[33]), .Z(n30928) );
  XOR U31632 ( .A(n30933), .B(n30693), .Z(n30695) );
  XOR U31633 ( .A(n30934), .B(n30935), .Z(n30693) );
  AND U31634 ( .A(n30936), .B(n30937), .Z(n30934) );
  AND U31635 ( .A(a[8]), .B(b[32]), .Z(n30933) );
  XOR U31636 ( .A(n30938), .B(n30698), .Z(n30700) );
  XOR U31637 ( .A(n30939), .B(n30940), .Z(n30698) );
  AND U31638 ( .A(n30941), .B(n30942), .Z(n30939) );
  AND U31639 ( .A(a[9]), .B(b[31]), .Z(n30938) );
  XOR U31640 ( .A(n30943), .B(n30703), .Z(n30705) );
  XOR U31641 ( .A(n30944), .B(n30945), .Z(n30703) );
  AND U31642 ( .A(n30946), .B(n30947), .Z(n30944) );
  AND U31643 ( .A(a[10]), .B(b[30]), .Z(n30943) );
  XOR U31644 ( .A(n30948), .B(n30708), .Z(n30710) );
  XOR U31645 ( .A(n30949), .B(n30950), .Z(n30708) );
  AND U31646 ( .A(n30951), .B(n30952), .Z(n30949) );
  AND U31647 ( .A(a[11]), .B(b[29]), .Z(n30948) );
  XOR U31648 ( .A(n30953), .B(n30713), .Z(n30715) );
  XOR U31649 ( .A(n30954), .B(n30955), .Z(n30713) );
  AND U31650 ( .A(n30956), .B(n30957), .Z(n30954) );
  AND U31651 ( .A(a[12]), .B(b[28]), .Z(n30953) );
  XOR U31652 ( .A(n30958), .B(n30718), .Z(n30720) );
  XOR U31653 ( .A(n30959), .B(n30960), .Z(n30718) );
  AND U31654 ( .A(n30961), .B(n30962), .Z(n30959) );
  AND U31655 ( .A(a[13]), .B(b[27]), .Z(n30958) );
  XOR U31656 ( .A(n30963), .B(n30723), .Z(n30725) );
  XOR U31657 ( .A(n30964), .B(n30965), .Z(n30723) );
  AND U31658 ( .A(n30966), .B(n30967), .Z(n30964) );
  AND U31659 ( .A(a[14]), .B(b[26]), .Z(n30963) );
  XOR U31660 ( .A(n30968), .B(n30728), .Z(n30730) );
  XOR U31661 ( .A(n30969), .B(n30970), .Z(n30728) );
  AND U31662 ( .A(n30971), .B(n30972), .Z(n30969) );
  AND U31663 ( .A(a[15]), .B(b[25]), .Z(n30968) );
  XOR U31664 ( .A(n30973), .B(n30733), .Z(n30735) );
  XOR U31665 ( .A(n30974), .B(n30975), .Z(n30733) );
  AND U31666 ( .A(n30976), .B(n30977), .Z(n30974) );
  AND U31667 ( .A(a[16]), .B(b[24]), .Z(n30973) );
  XOR U31668 ( .A(n30978), .B(n30738), .Z(n30740) );
  XOR U31669 ( .A(n30979), .B(n30980), .Z(n30738) );
  AND U31670 ( .A(n30981), .B(n30982), .Z(n30979) );
  AND U31671 ( .A(a[17]), .B(b[23]), .Z(n30978) );
  XOR U31672 ( .A(n30983), .B(n30743), .Z(n30745) );
  XOR U31673 ( .A(n30984), .B(n30985), .Z(n30743) );
  AND U31674 ( .A(n30986), .B(n30987), .Z(n30984) );
  AND U31675 ( .A(a[18]), .B(b[22]), .Z(n30983) );
  XOR U31676 ( .A(n30988), .B(n30748), .Z(n30750) );
  XOR U31677 ( .A(n30989), .B(n30990), .Z(n30748) );
  AND U31678 ( .A(n30991), .B(n30992), .Z(n30989) );
  AND U31679 ( .A(a[19]), .B(b[21]), .Z(n30988) );
  XOR U31680 ( .A(n30993), .B(n30753), .Z(n30755) );
  XOR U31681 ( .A(n30994), .B(n30995), .Z(n30753) );
  AND U31682 ( .A(n30996), .B(n30997), .Z(n30994) );
  AND U31683 ( .A(a[20]), .B(b[20]), .Z(n30993) );
  XOR U31684 ( .A(n30998), .B(n30758), .Z(n30760) );
  XOR U31685 ( .A(n30999), .B(n31000), .Z(n30758) );
  AND U31686 ( .A(n31001), .B(n31002), .Z(n30999) );
  AND U31687 ( .A(b[19]), .B(a[21]), .Z(n30998) );
  XOR U31688 ( .A(n31003), .B(n30763), .Z(n30765) );
  XOR U31689 ( .A(n31004), .B(n31005), .Z(n30763) );
  AND U31690 ( .A(n31006), .B(n31007), .Z(n31004) );
  AND U31691 ( .A(b[18]), .B(a[22]), .Z(n31003) );
  XOR U31692 ( .A(n31008), .B(n30768), .Z(n30770) );
  XOR U31693 ( .A(n31009), .B(n31010), .Z(n30768) );
  AND U31694 ( .A(n31011), .B(n31012), .Z(n31009) );
  AND U31695 ( .A(b[17]), .B(a[23]), .Z(n31008) );
  XOR U31696 ( .A(n31013), .B(n30773), .Z(n30775) );
  XOR U31697 ( .A(n31014), .B(n31015), .Z(n30773) );
  AND U31698 ( .A(n31016), .B(n31017), .Z(n31014) );
  AND U31699 ( .A(b[16]), .B(a[24]), .Z(n31013) );
  XOR U31700 ( .A(n31018), .B(n30778), .Z(n30780) );
  XOR U31701 ( .A(n31019), .B(n31020), .Z(n30778) );
  AND U31702 ( .A(n31021), .B(n31022), .Z(n31019) );
  AND U31703 ( .A(b[15]), .B(a[25]), .Z(n31018) );
  XOR U31704 ( .A(n31023), .B(n30783), .Z(n30785) );
  XOR U31705 ( .A(n31024), .B(n31025), .Z(n30783) );
  AND U31706 ( .A(n31026), .B(n31027), .Z(n31024) );
  AND U31707 ( .A(b[14]), .B(a[26]), .Z(n31023) );
  XOR U31708 ( .A(n31028), .B(n30788), .Z(n30790) );
  XOR U31709 ( .A(n31029), .B(n31030), .Z(n30788) );
  AND U31710 ( .A(n31031), .B(n31032), .Z(n31029) );
  AND U31711 ( .A(b[13]), .B(a[27]), .Z(n31028) );
  XOR U31712 ( .A(n31033), .B(n30793), .Z(n30795) );
  XOR U31713 ( .A(n31034), .B(n31035), .Z(n30793) );
  AND U31714 ( .A(n31036), .B(n31037), .Z(n31034) );
  AND U31715 ( .A(b[12]), .B(a[28]), .Z(n31033) );
  XOR U31716 ( .A(n31038), .B(n30798), .Z(n30800) );
  XOR U31717 ( .A(n31039), .B(n31040), .Z(n30798) );
  AND U31718 ( .A(n31041), .B(n31042), .Z(n31039) );
  AND U31719 ( .A(b[11]), .B(a[29]), .Z(n31038) );
  XOR U31720 ( .A(n31043), .B(n30803), .Z(n30805) );
  XOR U31721 ( .A(n31044), .B(n31045), .Z(n30803) );
  AND U31722 ( .A(n31046), .B(n31047), .Z(n31044) );
  AND U31723 ( .A(b[10]), .B(a[30]), .Z(n31043) );
  XOR U31724 ( .A(n31048), .B(n30808), .Z(n30810) );
  XOR U31725 ( .A(n31049), .B(n31050), .Z(n30808) );
  AND U31726 ( .A(n31051), .B(n31052), .Z(n31049) );
  AND U31727 ( .A(b[9]), .B(a[31]), .Z(n31048) );
  XOR U31728 ( .A(n31053), .B(n30813), .Z(n30815) );
  XOR U31729 ( .A(n31054), .B(n31055), .Z(n30813) );
  AND U31730 ( .A(n31056), .B(n31057), .Z(n31054) );
  AND U31731 ( .A(b[8]), .B(a[32]), .Z(n31053) );
  XOR U31732 ( .A(n31058), .B(n30818), .Z(n30820) );
  XOR U31733 ( .A(n31059), .B(n31060), .Z(n30818) );
  AND U31734 ( .A(n31061), .B(n31062), .Z(n31059) );
  AND U31735 ( .A(b[7]), .B(a[33]), .Z(n31058) );
  XOR U31736 ( .A(n31063), .B(n30823), .Z(n30825) );
  XOR U31737 ( .A(n31064), .B(n31065), .Z(n30823) );
  AND U31738 ( .A(n31066), .B(n31067), .Z(n31064) );
  AND U31739 ( .A(b[6]), .B(a[34]), .Z(n31063) );
  XOR U31740 ( .A(n31068), .B(n30828), .Z(n30830) );
  XOR U31741 ( .A(n31069), .B(n31070), .Z(n30828) );
  AND U31742 ( .A(n31071), .B(n31072), .Z(n31069) );
  AND U31743 ( .A(b[5]), .B(a[35]), .Z(n31068) );
  XOR U31744 ( .A(n31073), .B(n30833), .Z(n30835) );
  XOR U31745 ( .A(n31074), .B(n31075), .Z(n30833) );
  AND U31746 ( .A(n31076), .B(n31077), .Z(n31074) );
  AND U31747 ( .A(b[4]), .B(a[36]), .Z(n31073) );
  XNOR U31748 ( .A(n31078), .B(n31079), .Z(n30847) );
  NANDN U31749 ( .A(n31080), .B(n31081), .Z(n31079) );
  XOR U31750 ( .A(n31082), .B(n30838), .Z(n30840) );
  XNOR U31751 ( .A(n31083), .B(n31084), .Z(n30838) );
  AND U31752 ( .A(n31085), .B(n31086), .Z(n31083) );
  AND U31753 ( .A(b[3]), .B(a[37]), .Z(n31082) );
  XOR U31754 ( .A(n30854), .B(n30853), .Z(c[103]) );
  XOR U31755 ( .A(sreg[167]), .B(n30852), .Z(n30853) );
  XOR U31756 ( .A(n30859), .B(n31087), .Z(n30854) );
  XNOR U31757 ( .A(n30858), .B(n30852), .Z(n31087) );
  XOR U31758 ( .A(n31088), .B(n31089), .Z(n30852) );
  NOR U31759 ( .A(n31090), .B(n31091), .Z(n31088) );
  NAND U31760 ( .A(a[39]), .B(b[0]), .Z(n30858) );
  XNOR U31761 ( .A(n31080), .B(n31081), .Z(n30859) );
  XOR U31762 ( .A(n31078), .B(n31092), .Z(n31081) );
  NAND U31763 ( .A(b[1]), .B(a[38]), .Z(n31092) );
  XOR U31764 ( .A(n31086), .B(n31093), .Z(n31080) );
  XOR U31765 ( .A(n31078), .B(n31085), .Z(n31093) );
  XNOR U31766 ( .A(n31094), .B(n31084), .Z(n31085) );
  AND U31767 ( .A(b[2]), .B(a[37]), .Z(n31094) );
  NANDN U31768 ( .A(n31095), .B(n31096), .Z(n31078) );
  XOR U31769 ( .A(n31084), .B(n31076), .Z(n31097) );
  XNOR U31770 ( .A(n31075), .B(n31071), .Z(n31098) );
  XNOR U31771 ( .A(n31070), .B(n31066), .Z(n31099) );
  XNOR U31772 ( .A(n31065), .B(n31061), .Z(n31100) );
  XNOR U31773 ( .A(n31060), .B(n31056), .Z(n31101) );
  XNOR U31774 ( .A(n31055), .B(n31051), .Z(n31102) );
  XNOR U31775 ( .A(n31050), .B(n31046), .Z(n31103) );
  XNOR U31776 ( .A(n31045), .B(n31041), .Z(n31104) );
  XNOR U31777 ( .A(n31040), .B(n31036), .Z(n31105) );
  XNOR U31778 ( .A(n31035), .B(n31031), .Z(n31106) );
  XNOR U31779 ( .A(n31030), .B(n31026), .Z(n31107) );
  XNOR U31780 ( .A(n31025), .B(n31021), .Z(n31108) );
  XNOR U31781 ( .A(n31020), .B(n31016), .Z(n31109) );
  XNOR U31782 ( .A(n31015), .B(n31011), .Z(n31110) );
  XNOR U31783 ( .A(n31010), .B(n31006), .Z(n31111) );
  XNOR U31784 ( .A(n31005), .B(n31001), .Z(n31112) );
  XNOR U31785 ( .A(n31000), .B(n30996), .Z(n31113) );
  XNOR U31786 ( .A(n30995), .B(n30991), .Z(n31114) );
  XNOR U31787 ( .A(n30990), .B(n30986), .Z(n31115) );
  XNOR U31788 ( .A(n30985), .B(n30981), .Z(n31116) );
  XNOR U31789 ( .A(n30980), .B(n30976), .Z(n31117) );
  XNOR U31790 ( .A(n30975), .B(n30971), .Z(n31118) );
  XNOR U31791 ( .A(n30970), .B(n30966), .Z(n31119) );
  XNOR U31792 ( .A(n30965), .B(n30961), .Z(n31120) );
  XNOR U31793 ( .A(n30960), .B(n30956), .Z(n31121) );
  XNOR U31794 ( .A(n30955), .B(n30951), .Z(n31122) );
  XNOR U31795 ( .A(n30950), .B(n30946), .Z(n31123) );
  XNOR U31796 ( .A(n30945), .B(n30941), .Z(n31124) );
  XNOR U31797 ( .A(n30940), .B(n30936), .Z(n31125) );
  XNOR U31798 ( .A(n30935), .B(n30931), .Z(n31126) );
  XNOR U31799 ( .A(n30930), .B(n30926), .Z(n31127) );
  XNOR U31800 ( .A(n30925), .B(n30921), .Z(n31128) );
  XNOR U31801 ( .A(n30920), .B(n30916), .Z(n31129) );
  XNOR U31802 ( .A(n30915), .B(n30911), .Z(n31130) );
  XNOR U31803 ( .A(n30910), .B(n30906), .Z(n31131) );
  XNOR U31804 ( .A(n30905), .B(n30901), .Z(n31132) );
  XOR U31805 ( .A(n31133), .B(n30900), .Z(n30901) );
  AND U31806 ( .A(a[0]), .B(b[39]), .Z(n31133) );
  XOR U31807 ( .A(n31134), .B(n30900), .Z(n30902) );
  XNOR U31808 ( .A(n31135), .B(n31136), .Z(n30900) );
  AND U31809 ( .A(n31137), .B(n31138), .Z(n31135) );
  AND U31810 ( .A(a[1]), .B(b[38]), .Z(n31134) );
  XOR U31811 ( .A(n31139), .B(n30905), .Z(n30907) );
  XOR U31812 ( .A(n31140), .B(n31141), .Z(n30905) );
  AND U31813 ( .A(n31142), .B(n31143), .Z(n31140) );
  AND U31814 ( .A(a[2]), .B(b[37]), .Z(n31139) );
  XOR U31815 ( .A(n31144), .B(n30910), .Z(n30912) );
  XOR U31816 ( .A(n31145), .B(n31146), .Z(n30910) );
  AND U31817 ( .A(n31147), .B(n31148), .Z(n31145) );
  AND U31818 ( .A(a[3]), .B(b[36]), .Z(n31144) );
  XOR U31819 ( .A(n31149), .B(n30915), .Z(n30917) );
  XOR U31820 ( .A(n31150), .B(n31151), .Z(n30915) );
  AND U31821 ( .A(n31152), .B(n31153), .Z(n31150) );
  AND U31822 ( .A(a[4]), .B(b[35]), .Z(n31149) );
  XOR U31823 ( .A(n31154), .B(n30920), .Z(n30922) );
  XOR U31824 ( .A(n31155), .B(n31156), .Z(n30920) );
  AND U31825 ( .A(n31157), .B(n31158), .Z(n31155) );
  AND U31826 ( .A(a[5]), .B(b[34]), .Z(n31154) );
  XOR U31827 ( .A(n31159), .B(n30925), .Z(n30927) );
  XOR U31828 ( .A(n31160), .B(n31161), .Z(n30925) );
  AND U31829 ( .A(n31162), .B(n31163), .Z(n31160) );
  AND U31830 ( .A(a[6]), .B(b[33]), .Z(n31159) );
  XOR U31831 ( .A(n31164), .B(n30930), .Z(n30932) );
  XOR U31832 ( .A(n31165), .B(n31166), .Z(n30930) );
  AND U31833 ( .A(n31167), .B(n31168), .Z(n31165) );
  AND U31834 ( .A(a[7]), .B(b[32]), .Z(n31164) );
  XOR U31835 ( .A(n31169), .B(n30935), .Z(n30937) );
  XOR U31836 ( .A(n31170), .B(n31171), .Z(n30935) );
  AND U31837 ( .A(n31172), .B(n31173), .Z(n31170) );
  AND U31838 ( .A(a[8]), .B(b[31]), .Z(n31169) );
  XOR U31839 ( .A(n31174), .B(n30940), .Z(n30942) );
  XOR U31840 ( .A(n31175), .B(n31176), .Z(n30940) );
  AND U31841 ( .A(n31177), .B(n31178), .Z(n31175) );
  AND U31842 ( .A(a[9]), .B(b[30]), .Z(n31174) );
  XOR U31843 ( .A(n31179), .B(n30945), .Z(n30947) );
  XOR U31844 ( .A(n31180), .B(n31181), .Z(n30945) );
  AND U31845 ( .A(n31182), .B(n31183), .Z(n31180) );
  AND U31846 ( .A(a[10]), .B(b[29]), .Z(n31179) );
  XOR U31847 ( .A(n31184), .B(n30950), .Z(n30952) );
  XOR U31848 ( .A(n31185), .B(n31186), .Z(n30950) );
  AND U31849 ( .A(n31187), .B(n31188), .Z(n31185) );
  AND U31850 ( .A(a[11]), .B(b[28]), .Z(n31184) );
  XOR U31851 ( .A(n31189), .B(n30955), .Z(n30957) );
  XOR U31852 ( .A(n31190), .B(n31191), .Z(n30955) );
  AND U31853 ( .A(n31192), .B(n31193), .Z(n31190) );
  AND U31854 ( .A(a[12]), .B(b[27]), .Z(n31189) );
  XOR U31855 ( .A(n31194), .B(n30960), .Z(n30962) );
  XOR U31856 ( .A(n31195), .B(n31196), .Z(n30960) );
  AND U31857 ( .A(n31197), .B(n31198), .Z(n31195) );
  AND U31858 ( .A(a[13]), .B(b[26]), .Z(n31194) );
  XOR U31859 ( .A(n31199), .B(n30965), .Z(n30967) );
  XOR U31860 ( .A(n31200), .B(n31201), .Z(n30965) );
  AND U31861 ( .A(n31202), .B(n31203), .Z(n31200) );
  AND U31862 ( .A(a[14]), .B(b[25]), .Z(n31199) );
  XOR U31863 ( .A(n31204), .B(n30970), .Z(n30972) );
  XOR U31864 ( .A(n31205), .B(n31206), .Z(n30970) );
  AND U31865 ( .A(n31207), .B(n31208), .Z(n31205) );
  AND U31866 ( .A(a[15]), .B(b[24]), .Z(n31204) );
  XOR U31867 ( .A(n31209), .B(n30975), .Z(n30977) );
  XOR U31868 ( .A(n31210), .B(n31211), .Z(n30975) );
  AND U31869 ( .A(n31212), .B(n31213), .Z(n31210) );
  AND U31870 ( .A(a[16]), .B(b[23]), .Z(n31209) );
  XOR U31871 ( .A(n31214), .B(n30980), .Z(n30982) );
  XOR U31872 ( .A(n31215), .B(n31216), .Z(n30980) );
  AND U31873 ( .A(n31217), .B(n31218), .Z(n31215) );
  AND U31874 ( .A(a[17]), .B(b[22]), .Z(n31214) );
  XOR U31875 ( .A(n31219), .B(n30985), .Z(n30987) );
  XOR U31876 ( .A(n31220), .B(n31221), .Z(n30985) );
  AND U31877 ( .A(n31222), .B(n31223), .Z(n31220) );
  AND U31878 ( .A(a[18]), .B(b[21]), .Z(n31219) );
  XOR U31879 ( .A(n31224), .B(n30990), .Z(n30992) );
  XOR U31880 ( .A(n31225), .B(n31226), .Z(n30990) );
  AND U31881 ( .A(n31227), .B(n31228), .Z(n31225) );
  AND U31882 ( .A(a[19]), .B(b[20]), .Z(n31224) );
  XOR U31883 ( .A(n31229), .B(n30995), .Z(n30997) );
  XOR U31884 ( .A(n31230), .B(n31231), .Z(n30995) );
  AND U31885 ( .A(n31232), .B(n31233), .Z(n31230) );
  AND U31886 ( .A(b[19]), .B(a[20]), .Z(n31229) );
  XOR U31887 ( .A(n31234), .B(n31000), .Z(n31002) );
  XOR U31888 ( .A(n31235), .B(n31236), .Z(n31000) );
  AND U31889 ( .A(n31237), .B(n31238), .Z(n31235) );
  AND U31890 ( .A(b[18]), .B(a[21]), .Z(n31234) );
  XOR U31891 ( .A(n31239), .B(n31005), .Z(n31007) );
  XOR U31892 ( .A(n31240), .B(n31241), .Z(n31005) );
  AND U31893 ( .A(n31242), .B(n31243), .Z(n31240) );
  AND U31894 ( .A(b[17]), .B(a[22]), .Z(n31239) );
  XOR U31895 ( .A(n31244), .B(n31010), .Z(n31012) );
  XOR U31896 ( .A(n31245), .B(n31246), .Z(n31010) );
  AND U31897 ( .A(n31247), .B(n31248), .Z(n31245) );
  AND U31898 ( .A(b[16]), .B(a[23]), .Z(n31244) );
  XOR U31899 ( .A(n31249), .B(n31015), .Z(n31017) );
  XOR U31900 ( .A(n31250), .B(n31251), .Z(n31015) );
  AND U31901 ( .A(n31252), .B(n31253), .Z(n31250) );
  AND U31902 ( .A(b[15]), .B(a[24]), .Z(n31249) );
  XOR U31903 ( .A(n31254), .B(n31020), .Z(n31022) );
  XOR U31904 ( .A(n31255), .B(n31256), .Z(n31020) );
  AND U31905 ( .A(n31257), .B(n31258), .Z(n31255) );
  AND U31906 ( .A(b[14]), .B(a[25]), .Z(n31254) );
  XOR U31907 ( .A(n31259), .B(n31025), .Z(n31027) );
  XOR U31908 ( .A(n31260), .B(n31261), .Z(n31025) );
  AND U31909 ( .A(n31262), .B(n31263), .Z(n31260) );
  AND U31910 ( .A(b[13]), .B(a[26]), .Z(n31259) );
  XOR U31911 ( .A(n31264), .B(n31030), .Z(n31032) );
  XOR U31912 ( .A(n31265), .B(n31266), .Z(n31030) );
  AND U31913 ( .A(n31267), .B(n31268), .Z(n31265) );
  AND U31914 ( .A(b[12]), .B(a[27]), .Z(n31264) );
  XOR U31915 ( .A(n31269), .B(n31035), .Z(n31037) );
  XOR U31916 ( .A(n31270), .B(n31271), .Z(n31035) );
  AND U31917 ( .A(n31272), .B(n31273), .Z(n31270) );
  AND U31918 ( .A(b[11]), .B(a[28]), .Z(n31269) );
  XOR U31919 ( .A(n31274), .B(n31040), .Z(n31042) );
  XOR U31920 ( .A(n31275), .B(n31276), .Z(n31040) );
  AND U31921 ( .A(n31277), .B(n31278), .Z(n31275) );
  AND U31922 ( .A(b[10]), .B(a[29]), .Z(n31274) );
  XOR U31923 ( .A(n31279), .B(n31045), .Z(n31047) );
  XOR U31924 ( .A(n31280), .B(n31281), .Z(n31045) );
  AND U31925 ( .A(n31282), .B(n31283), .Z(n31280) );
  AND U31926 ( .A(b[9]), .B(a[30]), .Z(n31279) );
  XOR U31927 ( .A(n31284), .B(n31050), .Z(n31052) );
  XOR U31928 ( .A(n31285), .B(n31286), .Z(n31050) );
  AND U31929 ( .A(n31287), .B(n31288), .Z(n31285) );
  AND U31930 ( .A(b[8]), .B(a[31]), .Z(n31284) );
  XOR U31931 ( .A(n31289), .B(n31055), .Z(n31057) );
  XOR U31932 ( .A(n31290), .B(n31291), .Z(n31055) );
  AND U31933 ( .A(n31292), .B(n31293), .Z(n31290) );
  AND U31934 ( .A(b[7]), .B(a[32]), .Z(n31289) );
  XOR U31935 ( .A(n31294), .B(n31060), .Z(n31062) );
  XOR U31936 ( .A(n31295), .B(n31296), .Z(n31060) );
  AND U31937 ( .A(n31297), .B(n31298), .Z(n31295) );
  AND U31938 ( .A(b[6]), .B(a[33]), .Z(n31294) );
  XOR U31939 ( .A(n31299), .B(n31065), .Z(n31067) );
  XOR U31940 ( .A(n31300), .B(n31301), .Z(n31065) );
  AND U31941 ( .A(n31302), .B(n31303), .Z(n31300) );
  AND U31942 ( .A(b[5]), .B(a[34]), .Z(n31299) );
  XOR U31943 ( .A(n31304), .B(n31070), .Z(n31072) );
  XOR U31944 ( .A(n31305), .B(n31306), .Z(n31070) );
  AND U31945 ( .A(n31307), .B(n31308), .Z(n31305) );
  AND U31946 ( .A(b[4]), .B(a[35]), .Z(n31304) );
  XNOR U31947 ( .A(n31309), .B(n31310), .Z(n31084) );
  NANDN U31948 ( .A(n31311), .B(n31312), .Z(n31310) );
  XOR U31949 ( .A(n31313), .B(n31075), .Z(n31077) );
  XNOR U31950 ( .A(n31314), .B(n31315), .Z(n31075) );
  AND U31951 ( .A(n31316), .B(n31317), .Z(n31314) );
  AND U31952 ( .A(b[3]), .B(a[36]), .Z(n31313) );
  XOR U31953 ( .A(n31091), .B(n31090), .Z(c[102]) );
  XOR U31954 ( .A(sreg[166]), .B(n31089), .Z(n31090) );
  XOR U31955 ( .A(n31096), .B(n31318), .Z(n31091) );
  XNOR U31956 ( .A(n31095), .B(n31089), .Z(n31318) );
  XOR U31957 ( .A(n31319), .B(n31320), .Z(n31089) );
  NOR U31958 ( .A(n31321), .B(n31322), .Z(n31319) );
  NAND U31959 ( .A(a[38]), .B(b[0]), .Z(n31095) );
  XNOR U31960 ( .A(n31311), .B(n31312), .Z(n31096) );
  XOR U31961 ( .A(n31309), .B(n31323), .Z(n31312) );
  NAND U31962 ( .A(b[1]), .B(a[37]), .Z(n31323) );
  XOR U31963 ( .A(n31317), .B(n31324), .Z(n31311) );
  XOR U31964 ( .A(n31309), .B(n31316), .Z(n31324) );
  XNOR U31965 ( .A(n31325), .B(n31315), .Z(n31316) );
  AND U31966 ( .A(b[2]), .B(a[36]), .Z(n31325) );
  NANDN U31967 ( .A(n31326), .B(n31327), .Z(n31309) );
  XOR U31968 ( .A(n31315), .B(n31307), .Z(n31328) );
  XNOR U31969 ( .A(n31306), .B(n31302), .Z(n31329) );
  XNOR U31970 ( .A(n31301), .B(n31297), .Z(n31330) );
  XNOR U31971 ( .A(n31296), .B(n31292), .Z(n31331) );
  XNOR U31972 ( .A(n31291), .B(n31287), .Z(n31332) );
  XNOR U31973 ( .A(n31286), .B(n31282), .Z(n31333) );
  XNOR U31974 ( .A(n31281), .B(n31277), .Z(n31334) );
  XNOR U31975 ( .A(n31276), .B(n31272), .Z(n31335) );
  XNOR U31976 ( .A(n31271), .B(n31267), .Z(n31336) );
  XNOR U31977 ( .A(n31266), .B(n31262), .Z(n31337) );
  XNOR U31978 ( .A(n31261), .B(n31257), .Z(n31338) );
  XNOR U31979 ( .A(n31256), .B(n31252), .Z(n31339) );
  XNOR U31980 ( .A(n31251), .B(n31247), .Z(n31340) );
  XNOR U31981 ( .A(n31246), .B(n31242), .Z(n31341) );
  XNOR U31982 ( .A(n31241), .B(n31237), .Z(n31342) );
  XNOR U31983 ( .A(n31236), .B(n31232), .Z(n31343) );
  XNOR U31984 ( .A(n31231), .B(n31227), .Z(n31344) );
  XNOR U31985 ( .A(n31226), .B(n31222), .Z(n31345) );
  XNOR U31986 ( .A(n31221), .B(n31217), .Z(n31346) );
  XNOR U31987 ( .A(n31216), .B(n31212), .Z(n31347) );
  XNOR U31988 ( .A(n31211), .B(n31207), .Z(n31348) );
  XNOR U31989 ( .A(n31206), .B(n31202), .Z(n31349) );
  XNOR U31990 ( .A(n31201), .B(n31197), .Z(n31350) );
  XNOR U31991 ( .A(n31196), .B(n31192), .Z(n31351) );
  XNOR U31992 ( .A(n31191), .B(n31187), .Z(n31352) );
  XNOR U31993 ( .A(n31186), .B(n31182), .Z(n31353) );
  XNOR U31994 ( .A(n31181), .B(n31177), .Z(n31354) );
  XNOR U31995 ( .A(n31176), .B(n31172), .Z(n31355) );
  XNOR U31996 ( .A(n31171), .B(n31167), .Z(n31356) );
  XNOR U31997 ( .A(n31166), .B(n31162), .Z(n31357) );
  XNOR U31998 ( .A(n31161), .B(n31157), .Z(n31358) );
  XNOR U31999 ( .A(n31156), .B(n31152), .Z(n31359) );
  XNOR U32000 ( .A(n31151), .B(n31147), .Z(n31360) );
  XNOR U32001 ( .A(n31146), .B(n31142), .Z(n31361) );
  XNOR U32002 ( .A(n31141), .B(n31137), .Z(n31362) );
  XNOR U32003 ( .A(n31363), .B(n31136), .Z(n31137) );
  AND U32004 ( .A(a[0]), .B(b[38]), .Z(n31363) );
  XNOR U32005 ( .A(n31364), .B(n31136), .Z(n31138) );
  XNOR U32006 ( .A(n31365), .B(n31366), .Z(n31136) );
  AND U32007 ( .A(n31367), .B(n31368), .Z(n31365) );
  AND U32008 ( .A(a[1]), .B(b[37]), .Z(n31364) );
  XOR U32009 ( .A(n31369), .B(n31141), .Z(n31143) );
  XOR U32010 ( .A(n31370), .B(n31371), .Z(n31141) );
  AND U32011 ( .A(n31372), .B(n31373), .Z(n31370) );
  AND U32012 ( .A(a[2]), .B(b[36]), .Z(n31369) );
  XOR U32013 ( .A(n31374), .B(n31146), .Z(n31148) );
  XOR U32014 ( .A(n31375), .B(n31376), .Z(n31146) );
  AND U32015 ( .A(n31377), .B(n31378), .Z(n31375) );
  AND U32016 ( .A(a[3]), .B(b[35]), .Z(n31374) );
  XOR U32017 ( .A(n31379), .B(n31151), .Z(n31153) );
  XOR U32018 ( .A(n31380), .B(n31381), .Z(n31151) );
  AND U32019 ( .A(n31382), .B(n31383), .Z(n31380) );
  AND U32020 ( .A(a[4]), .B(b[34]), .Z(n31379) );
  XOR U32021 ( .A(n31384), .B(n31156), .Z(n31158) );
  XOR U32022 ( .A(n31385), .B(n31386), .Z(n31156) );
  AND U32023 ( .A(n31387), .B(n31388), .Z(n31385) );
  AND U32024 ( .A(a[5]), .B(b[33]), .Z(n31384) );
  XOR U32025 ( .A(n31389), .B(n31161), .Z(n31163) );
  XOR U32026 ( .A(n31390), .B(n31391), .Z(n31161) );
  AND U32027 ( .A(n31392), .B(n31393), .Z(n31390) );
  AND U32028 ( .A(a[6]), .B(b[32]), .Z(n31389) );
  XOR U32029 ( .A(n31394), .B(n31166), .Z(n31168) );
  XOR U32030 ( .A(n31395), .B(n31396), .Z(n31166) );
  AND U32031 ( .A(n31397), .B(n31398), .Z(n31395) );
  AND U32032 ( .A(a[7]), .B(b[31]), .Z(n31394) );
  XOR U32033 ( .A(n31399), .B(n31171), .Z(n31173) );
  XOR U32034 ( .A(n31400), .B(n31401), .Z(n31171) );
  AND U32035 ( .A(n31402), .B(n31403), .Z(n31400) );
  AND U32036 ( .A(a[8]), .B(b[30]), .Z(n31399) );
  XOR U32037 ( .A(n31404), .B(n31176), .Z(n31178) );
  XOR U32038 ( .A(n31405), .B(n31406), .Z(n31176) );
  AND U32039 ( .A(n31407), .B(n31408), .Z(n31405) );
  AND U32040 ( .A(a[9]), .B(b[29]), .Z(n31404) );
  XOR U32041 ( .A(n31409), .B(n31181), .Z(n31183) );
  XOR U32042 ( .A(n31410), .B(n31411), .Z(n31181) );
  AND U32043 ( .A(n31412), .B(n31413), .Z(n31410) );
  AND U32044 ( .A(a[10]), .B(b[28]), .Z(n31409) );
  XOR U32045 ( .A(n31414), .B(n31186), .Z(n31188) );
  XOR U32046 ( .A(n31415), .B(n31416), .Z(n31186) );
  AND U32047 ( .A(n31417), .B(n31418), .Z(n31415) );
  AND U32048 ( .A(a[11]), .B(b[27]), .Z(n31414) );
  XOR U32049 ( .A(n31419), .B(n31191), .Z(n31193) );
  XOR U32050 ( .A(n31420), .B(n31421), .Z(n31191) );
  AND U32051 ( .A(n31422), .B(n31423), .Z(n31420) );
  AND U32052 ( .A(a[12]), .B(b[26]), .Z(n31419) );
  XOR U32053 ( .A(n31424), .B(n31196), .Z(n31198) );
  XOR U32054 ( .A(n31425), .B(n31426), .Z(n31196) );
  AND U32055 ( .A(n31427), .B(n31428), .Z(n31425) );
  AND U32056 ( .A(a[13]), .B(b[25]), .Z(n31424) );
  XOR U32057 ( .A(n31429), .B(n31201), .Z(n31203) );
  XOR U32058 ( .A(n31430), .B(n31431), .Z(n31201) );
  AND U32059 ( .A(n31432), .B(n31433), .Z(n31430) );
  AND U32060 ( .A(a[14]), .B(b[24]), .Z(n31429) );
  XOR U32061 ( .A(n31434), .B(n31206), .Z(n31208) );
  XOR U32062 ( .A(n31435), .B(n31436), .Z(n31206) );
  AND U32063 ( .A(n31437), .B(n31438), .Z(n31435) );
  AND U32064 ( .A(a[15]), .B(b[23]), .Z(n31434) );
  XOR U32065 ( .A(n31439), .B(n31211), .Z(n31213) );
  XOR U32066 ( .A(n31440), .B(n31441), .Z(n31211) );
  AND U32067 ( .A(n31442), .B(n31443), .Z(n31440) );
  AND U32068 ( .A(a[16]), .B(b[22]), .Z(n31439) );
  XOR U32069 ( .A(n31444), .B(n31216), .Z(n31218) );
  XOR U32070 ( .A(n31445), .B(n31446), .Z(n31216) );
  AND U32071 ( .A(n31447), .B(n31448), .Z(n31445) );
  AND U32072 ( .A(a[17]), .B(b[21]), .Z(n31444) );
  XOR U32073 ( .A(n31449), .B(n31221), .Z(n31223) );
  XOR U32074 ( .A(n31450), .B(n31451), .Z(n31221) );
  AND U32075 ( .A(n31452), .B(n31453), .Z(n31450) );
  AND U32076 ( .A(a[18]), .B(b[20]), .Z(n31449) );
  XOR U32077 ( .A(n31454), .B(n31226), .Z(n31228) );
  XOR U32078 ( .A(n31455), .B(n31456), .Z(n31226) );
  AND U32079 ( .A(n31457), .B(n31458), .Z(n31455) );
  AND U32080 ( .A(a[19]), .B(b[19]), .Z(n31454) );
  XOR U32081 ( .A(n31459), .B(n31231), .Z(n31233) );
  XOR U32082 ( .A(n31460), .B(n31461), .Z(n31231) );
  AND U32083 ( .A(n31462), .B(n31463), .Z(n31460) );
  AND U32084 ( .A(b[18]), .B(a[20]), .Z(n31459) );
  XOR U32085 ( .A(n31464), .B(n31236), .Z(n31238) );
  XOR U32086 ( .A(n31465), .B(n31466), .Z(n31236) );
  AND U32087 ( .A(n31467), .B(n31468), .Z(n31465) );
  AND U32088 ( .A(b[17]), .B(a[21]), .Z(n31464) );
  XOR U32089 ( .A(n31469), .B(n31241), .Z(n31243) );
  XOR U32090 ( .A(n31470), .B(n31471), .Z(n31241) );
  AND U32091 ( .A(n31472), .B(n31473), .Z(n31470) );
  AND U32092 ( .A(b[16]), .B(a[22]), .Z(n31469) );
  XOR U32093 ( .A(n31474), .B(n31246), .Z(n31248) );
  XOR U32094 ( .A(n31475), .B(n31476), .Z(n31246) );
  AND U32095 ( .A(n31477), .B(n31478), .Z(n31475) );
  AND U32096 ( .A(b[15]), .B(a[23]), .Z(n31474) );
  XOR U32097 ( .A(n31479), .B(n31251), .Z(n31253) );
  XOR U32098 ( .A(n31480), .B(n31481), .Z(n31251) );
  AND U32099 ( .A(n31482), .B(n31483), .Z(n31480) );
  AND U32100 ( .A(b[14]), .B(a[24]), .Z(n31479) );
  XOR U32101 ( .A(n31484), .B(n31256), .Z(n31258) );
  XOR U32102 ( .A(n31485), .B(n31486), .Z(n31256) );
  AND U32103 ( .A(n31487), .B(n31488), .Z(n31485) );
  AND U32104 ( .A(b[13]), .B(a[25]), .Z(n31484) );
  XOR U32105 ( .A(n31489), .B(n31261), .Z(n31263) );
  XOR U32106 ( .A(n31490), .B(n31491), .Z(n31261) );
  AND U32107 ( .A(n31492), .B(n31493), .Z(n31490) );
  AND U32108 ( .A(b[12]), .B(a[26]), .Z(n31489) );
  XOR U32109 ( .A(n31494), .B(n31266), .Z(n31268) );
  XOR U32110 ( .A(n31495), .B(n31496), .Z(n31266) );
  AND U32111 ( .A(n31497), .B(n31498), .Z(n31495) );
  AND U32112 ( .A(b[11]), .B(a[27]), .Z(n31494) );
  XOR U32113 ( .A(n31499), .B(n31271), .Z(n31273) );
  XOR U32114 ( .A(n31500), .B(n31501), .Z(n31271) );
  AND U32115 ( .A(n31502), .B(n31503), .Z(n31500) );
  AND U32116 ( .A(b[10]), .B(a[28]), .Z(n31499) );
  XOR U32117 ( .A(n31504), .B(n31276), .Z(n31278) );
  XOR U32118 ( .A(n31505), .B(n31506), .Z(n31276) );
  AND U32119 ( .A(n31507), .B(n31508), .Z(n31505) );
  AND U32120 ( .A(b[9]), .B(a[29]), .Z(n31504) );
  XOR U32121 ( .A(n31509), .B(n31281), .Z(n31283) );
  XOR U32122 ( .A(n31510), .B(n31511), .Z(n31281) );
  AND U32123 ( .A(n31512), .B(n31513), .Z(n31510) );
  AND U32124 ( .A(b[8]), .B(a[30]), .Z(n31509) );
  XOR U32125 ( .A(n31514), .B(n31286), .Z(n31288) );
  XOR U32126 ( .A(n31515), .B(n31516), .Z(n31286) );
  AND U32127 ( .A(n31517), .B(n31518), .Z(n31515) );
  AND U32128 ( .A(b[7]), .B(a[31]), .Z(n31514) );
  XOR U32129 ( .A(n31519), .B(n31291), .Z(n31293) );
  XOR U32130 ( .A(n31520), .B(n31521), .Z(n31291) );
  AND U32131 ( .A(n31522), .B(n31523), .Z(n31520) );
  AND U32132 ( .A(b[6]), .B(a[32]), .Z(n31519) );
  XOR U32133 ( .A(n31524), .B(n31296), .Z(n31298) );
  XOR U32134 ( .A(n31525), .B(n31526), .Z(n31296) );
  AND U32135 ( .A(n31527), .B(n31528), .Z(n31525) );
  AND U32136 ( .A(b[5]), .B(a[33]), .Z(n31524) );
  XOR U32137 ( .A(n31529), .B(n31301), .Z(n31303) );
  XOR U32138 ( .A(n31530), .B(n31531), .Z(n31301) );
  AND U32139 ( .A(n31532), .B(n31533), .Z(n31530) );
  AND U32140 ( .A(b[4]), .B(a[34]), .Z(n31529) );
  XNOR U32141 ( .A(n31534), .B(n31535), .Z(n31315) );
  NANDN U32142 ( .A(n31536), .B(n31537), .Z(n31535) );
  XOR U32143 ( .A(n31538), .B(n31306), .Z(n31308) );
  XNOR U32144 ( .A(n31539), .B(n31540), .Z(n31306) );
  AND U32145 ( .A(n31541), .B(n31542), .Z(n31539) );
  AND U32146 ( .A(b[3]), .B(a[35]), .Z(n31538) );
  XOR U32147 ( .A(n31322), .B(n31321), .Z(c[101]) );
  XOR U32148 ( .A(sreg[165]), .B(n31320), .Z(n31321) );
  XOR U32149 ( .A(n31327), .B(n31543), .Z(n31322) );
  XNOR U32150 ( .A(n31326), .B(n31320), .Z(n31543) );
  XOR U32151 ( .A(n31544), .B(n31545), .Z(n31320) );
  NOR U32152 ( .A(n31546), .B(n31547), .Z(n31544) );
  NAND U32153 ( .A(a[37]), .B(b[0]), .Z(n31326) );
  XNOR U32154 ( .A(n31536), .B(n31537), .Z(n31327) );
  XOR U32155 ( .A(n31534), .B(n31548), .Z(n31537) );
  NAND U32156 ( .A(b[1]), .B(a[36]), .Z(n31548) );
  XOR U32157 ( .A(n31542), .B(n31549), .Z(n31536) );
  XOR U32158 ( .A(n31534), .B(n31541), .Z(n31549) );
  XNOR U32159 ( .A(n31550), .B(n31540), .Z(n31541) );
  AND U32160 ( .A(b[2]), .B(a[35]), .Z(n31550) );
  NANDN U32161 ( .A(n31551), .B(n31552), .Z(n31534) );
  XOR U32162 ( .A(n31540), .B(n31532), .Z(n31553) );
  XNOR U32163 ( .A(n31531), .B(n31527), .Z(n31554) );
  XNOR U32164 ( .A(n31526), .B(n31522), .Z(n31555) );
  XNOR U32165 ( .A(n31521), .B(n31517), .Z(n31556) );
  XNOR U32166 ( .A(n31516), .B(n31512), .Z(n31557) );
  XNOR U32167 ( .A(n31511), .B(n31507), .Z(n31558) );
  XNOR U32168 ( .A(n31506), .B(n31502), .Z(n31559) );
  XNOR U32169 ( .A(n31501), .B(n31497), .Z(n31560) );
  XNOR U32170 ( .A(n31496), .B(n31492), .Z(n31561) );
  XNOR U32171 ( .A(n31491), .B(n31487), .Z(n31562) );
  XNOR U32172 ( .A(n31486), .B(n31482), .Z(n31563) );
  XNOR U32173 ( .A(n31481), .B(n31477), .Z(n31564) );
  XNOR U32174 ( .A(n31476), .B(n31472), .Z(n31565) );
  XNOR U32175 ( .A(n31471), .B(n31467), .Z(n31566) );
  XNOR U32176 ( .A(n31466), .B(n31462), .Z(n31567) );
  XNOR U32177 ( .A(n31461), .B(n31457), .Z(n31568) );
  XNOR U32178 ( .A(n31456), .B(n31452), .Z(n31569) );
  XNOR U32179 ( .A(n31451), .B(n31447), .Z(n31570) );
  XNOR U32180 ( .A(n31446), .B(n31442), .Z(n31571) );
  XNOR U32181 ( .A(n31441), .B(n31437), .Z(n31572) );
  XNOR U32182 ( .A(n31436), .B(n31432), .Z(n31573) );
  XNOR U32183 ( .A(n31431), .B(n31427), .Z(n31574) );
  XNOR U32184 ( .A(n31426), .B(n31422), .Z(n31575) );
  XNOR U32185 ( .A(n31421), .B(n31417), .Z(n31576) );
  XNOR U32186 ( .A(n31416), .B(n31412), .Z(n31577) );
  XNOR U32187 ( .A(n31411), .B(n31407), .Z(n31578) );
  XNOR U32188 ( .A(n31406), .B(n31402), .Z(n31579) );
  XNOR U32189 ( .A(n31401), .B(n31397), .Z(n31580) );
  XNOR U32190 ( .A(n31396), .B(n31392), .Z(n31581) );
  XNOR U32191 ( .A(n31391), .B(n31387), .Z(n31582) );
  XNOR U32192 ( .A(n31386), .B(n31382), .Z(n31583) );
  XNOR U32193 ( .A(n31381), .B(n31377), .Z(n31584) );
  XNOR U32194 ( .A(n31376), .B(n31372), .Z(n31585) );
  XNOR U32195 ( .A(n31371), .B(n31367), .Z(n31586) );
  XOR U32196 ( .A(n31587), .B(n31366), .Z(n31367) );
  AND U32197 ( .A(a[0]), .B(b[37]), .Z(n31587) );
  XOR U32198 ( .A(n31588), .B(n31366), .Z(n31368) );
  XNOR U32199 ( .A(n31589), .B(n31590), .Z(n31366) );
  AND U32200 ( .A(n31591), .B(n31592), .Z(n31589) );
  AND U32201 ( .A(a[1]), .B(b[36]), .Z(n31588) );
  XOR U32202 ( .A(n31593), .B(n31371), .Z(n31373) );
  XOR U32203 ( .A(n31594), .B(n31595), .Z(n31371) );
  AND U32204 ( .A(n31596), .B(n31597), .Z(n31594) );
  AND U32205 ( .A(a[2]), .B(b[35]), .Z(n31593) );
  XOR U32206 ( .A(n31598), .B(n31376), .Z(n31378) );
  XOR U32207 ( .A(n31599), .B(n31600), .Z(n31376) );
  AND U32208 ( .A(n31601), .B(n31602), .Z(n31599) );
  AND U32209 ( .A(a[3]), .B(b[34]), .Z(n31598) );
  XOR U32210 ( .A(n31603), .B(n31381), .Z(n31383) );
  XOR U32211 ( .A(n31604), .B(n31605), .Z(n31381) );
  AND U32212 ( .A(n31606), .B(n31607), .Z(n31604) );
  AND U32213 ( .A(a[4]), .B(b[33]), .Z(n31603) );
  XOR U32214 ( .A(n31608), .B(n31386), .Z(n31388) );
  XOR U32215 ( .A(n31609), .B(n31610), .Z(n31386) );
  AND U32216 ( .A(n31611), .B(n31612), .Z(n31609) );
  AND U32217 ( .A(a[5]), .B(b[32]), .Z(n31608) );
  XOR U32218 ( .A(n31613), .B(n31391), .Z(n31393) );
  XOR U32219 ( .A(n31614), .B(n31615), .Z(n31391) );
  AND U32220 ( .A(n31616), .B(n31617), .Z(n31614) );
  AND U32221 ( .A(a[6]), .B(b[31]), .Z(n31613) );
  XOR U32222 ( .A(n31618), .B(n31396), .Z(n31398) );
  XOR U32223 ( .A(n31619), .B(n31620), .Z(n31396) );
  AND U32224 ( .A(n31621), .B(n31622), .Z(n31619) );
  AND U32225 ( .A(a[7]), .B(b[30]), .Z(n31618) );
  XOR U32226 ( .A(n31623), .B(n31401), .Z(n31403) );
  XOR U32227 ( .A(n31624), .B(n31625), .Z(n31401) );
  AND U32228 ( .A(n31626), .B(n31627), .Z(n31624) );
  AND U32229 ( .A(a[8]), .B(b[29]), .Z(n31623) );
  XOR U32230 ( .A(n31628), .B(n31406), .Z(n31408) );
  XOR U32231 ( .A(n31629), .B(n31630), .Z(n31406) );
  AND U32232 ( .A(n31631), .B(n31632), .Z(n31629) );
  AND U32233 ( .A(a[9]), .B(b[28]), .Z(n31628) );
  XOR U32234 ( .A(n31633), .B(n31411), .Z(n31413) );
  XOR U32235 ( .A(n31634), .B(n31635), .Z(n31411) );
  AND U32236 ( .A(n31636), .B(n31637), .Z(n31634) );
  AND U32237 ( .A(a[10]), .B(b[27]), .Z(n31633) );
  XOR U32238 ( .A(n31638), .B(n31416), .Z(n31418) );
  XOR U32239 ( .A(n31639), .B(n31640), .Z(n31416) );
  AND U32240 ( .A(n31641), .B(n31642), .Z(n31639) );
  AND U32241 ( .A(a[11]), .B(b[26]), .Z(n31638) );
  XOR U32242 ( .A(n31643), .B(n31421), .Z(n31423) );
  XOR U32243 ( .A(n31644), .B(n31645), .Z(n31421) );
  AND U32244 ( .A(n31646), .B(n31647), .Z(n31644) );
  AND U32245 ( .A(a[12]), .B(b[25]), .Z(n31643) );
  XOR U32246 ( .A(n31648), .B(n31426), .Z(n31428) );
  XOR U32247 ( .A(n31649), .B(n31650), .Z(n31426) );
  AND U32248 ( .A(n31651), .B(n31652), .Z(n31649) );
  AND U32249 ( .A(a[13]), .B(b[24]), .Z(n31648) );
  XOR U32250 ( .A(n31653), .B(n31431), .Z(n31433) );
  XOR U32251 ( .A(n31654), .B(n31655), .Z(n31431) );
  AND U32252 ( .A(n31656), .B(n31657), .Z(n31654) );
  AND U32253 ( .A(a[14]), .B(b[23]), .Z(n31653) );
  XOR U32254 ( .A(n31658), .B(n31436), .Z(n31438) );
  XOR U32255 ( .A(n31659), .B(n31660), .Z(n31436) );
  AND U32256 ( .A(n31661), .B(n31662), .Z(n31659) );
  AND U32257 ( .A(a[15]), .B(b[22]), .Z(n31658) );
  XOR U32258 ( .A(n31663), .B(n31441), .Z(n31443) );
  XOR U32259 ( .A(n31664), .B(n31665), .Z(n31441) );
  AND U32260 ( .A(n31666), .B(n31667), .Z(n31664) );
  AND U32261 ( .A(a[16]), .B(b[21]), .Z(n31663) );
  XOR U32262 ( .A(n31668), .B(n31446), .Z(n31448) );
  XOR U32263 ( .A(n31669), .B(n31670), .Z(n31446) );
  AND U32264 ( .A(n31671), .B(n31672), .Z(n31669) );
  AND U32265 ( .A(a[17]), .B(b[20]), .Z(n31668) );
  XOR U32266 ( .A(n31673), .B(n31451), .Z(n31453) );
  XOR U32267 ( .A(n31674), .B(n31675), .Z(n31451) );
  AND U32268 ( .A(n31676), .B(n31677), .Z(n31674) );
  AND U32269 ( .A(a[18]), .B(b[19]), .Z(n31673) );
  XOR U32270 ( .A(n31678), .B(n31456), .Z(n31458) );
  XOR U32271 ( .A(n31679), .B(n31680), .Z(n31456) );
  AND U32272 ( .A(n31681), .B(n31682), .Z(n31679) );
  AND U32273 ( .A(b[18]), .B(a[19]), .Z(n31678) );
  XOR U32274 ( .A(n31683), .B(n31461), .Z(n31463) );
  XOR U32275 ( .A(n31684), .B(n31685), .Z(n31461) );
  AND U32276 ( .A(n31686), .B(n31687), .Z(n31684) );
  AND U32277 ( .A(b[17]), .B(a[20]), .Z(n31683) );
  XOR U32278 ( .A(n31688), .B(n31466), .Z(n31468) );
  XOR U32279 ( .A(n31689), .B(n31690), .Z(n31466) );
  AND U32280 ( .A(n31691), .B(n31692), .Z(n31689) );
  AND U32281 ( .A(b[16]), .B(a[21]), .Z(n31688) );
  XOR U32282 ( .A(n31693), .B(n31471), .Z(n31473) );
  XOR U32283 ( .A(n31694), .B(n31695), .Z(n31471) );
  AND U32284 ( .A(n31696), .B(n31697), .Z(n31694) );
  AND U32285 ( .A(b[15]), .B(a[22]), .Z(n31693) );
  XOR U32286 ( .A(n31698), .B(n31476), .Z(n31478) );
  XOR U32287 ( .A(n31699), .B(n31700), .Z(n31476) );
  AND U32288 ( .A(n31701), .B(n31702), .Z(n31699) );
  AND U32289 ( .A(b[14]), .B(a[23]), .Z(n31698) );
  XOR U32290 ( .A(n31703), .B(n31481), .Z(n31483) );
  XOR U32291 ( .A(n31704), .B(n31705), .Z(n31481) );
  AND U32292 ( .A(n31706), .B(n31707), .Z(n31704) );
  AND U32293 ( .A(b[13]), .B(a[24]), .Z(n31703) );
  XOR U32294 ( .A(n31708), .B(n31486), .Z(n31488) );
  XOR U32295 ( .A(n31709), .B(n31710), .Z(n31486) );
  AND U32296 ( .A(n31711), .B(n31712), .Z(n31709) );
  AND U32297 ( .A(b[12]), .B(a[25]), .Z(n31708) );
  XOR U32298 ( .A(n31713), .B(n31491), .Z(n31493) );
  XOR U32299 ( .A(n31714), .B(n31715), .Z(n31491) );
  AND U32300 ( .A(n31716), .B(n31717), .Z(n31714) );
  AND U32301 ( .A(b[11]), .B(a[26]), .Z(n31713) );
  XOR U32302 ( .A(n31718), .B(n31496), .Z(n31498) );
  XOR U32303 ( .A(n31719), .B(n31720), .Z(n31496) );
  AND U32304 ( .A(n31721), .B(n31722), .Z(n31719) );
  AND U32305 ( .A(b[10]), .B(a[27]), .Z(n31718) );
  XOR U32306 ( .A(n31723), .B(n31501), .Z(n31503) );
  XOR U32307 ( .A(n31724), .B(n31725), .Z(n31501) );
  AND U32308 ( .A(n31726), .B(n31727), .Z(n31724) );
  AND U32309 ( .A(b[9]), .B(a[28]), .Z(n31723) );
  XOR U32310 ( .A(n31728), .B(n31506), .Z(n31508) );
  XOR U32311 ( .A(n31729), .B(n31730), .Z(n31506) );
  AND U32312 ( .A(n31731), .B(n31732), .Z(n31729) );
  AND U32313 ( .A(b[8]), .B(a[29]), .Z(n31728) );
  XOR U32314 ( .A(n31733), .B(n31511), .Z(n31513) );
  XOR U32315 ( .A(n31734), .B(n31735), .Z(n31511) );
  AND U32316 ( .A(n31736), .B(n31737), .Z(n31734) );
  AND U32317 ( .A(b[7]), .B(a[30]), .Z(n31733) );
  XOR U32318 ( .A(n31738), .B(n31516), .Z(n31518) );
  XOR U32319 ( .A(n31739), .B(n31740), .Z(n31516) );
  AND U32320 ( .A(n31741), .B(n31742), .Z(n31739) );
  AND U32321 ( .A(b[6]), .B(a[31]), .Z(n31738) );
  XOR U32322 ( .A(n31743), .B(n31521), .Z(n31523) );
  XOR U32323 ( .A(n31744), .B(n31745), .Z(n31521) );
  AND U32324 ( .A(n31746), .B(n31747), .Z(n31744) );
  AND U32325 ( .A(b[5]), .B(a[32]), .Z(n31743) );
  XOR U32326 ( .A(n31748), .B(n31526), .Z(n31528) );
  XOR U32327 ( .A(n31749), .B(n31750), .Z(n31526) );
  AND U32328 ( .A(n31751), .B(n31752), .Z(n31749) );
  AND U32329 ( .A(b[4]), .B(a[33]), .Z(n31748) );
  XNOR U32330 ( .A(n31753), .B(n31754), .Z(n31540) );
  NANDN U32331 ( .A(n31755), .B(n31756), .Z(n31754) );
  XOR U32332 ( .A(n31757), .B(n31531), .Z(n31533) );
  XNOR U32333 ( .A(n31758), .B(n31759), .Z(n31531) );
  AND U32334 ( .A(n31760), .B(n31761), .Z(n31758) );
  AND U32335 ( .A(b[3]), .B(a[34]), .Z(n31757) );
  XOR U32336 ( .A(n31547), .B(n31546), .Z(c[100]) );
  XOR U32337 ( .A(sreg[164]), .B(n31545), .Z(n31546) );
  XOR U32338 ( .A(n31552), .B(n31762), .Z(n31547) );
  XNOR U32339 ( .A(n31551), .B(n31545), .Z(n31762) );
  XOR U32340 ( .A(n31763), .B(n31764), .Z(n31545) );
  NOR U32341 ( .A(n23671), .B(n23670), .Z(n31763) );
  XOR U32342 ( .A(n31765), .B(n31766), .Z(n23670) );
  XNOR U32343 ( .A(n31767), .B(n31764), .Z(n31766) );
  XOR U32344 ( .A(sreg[163]), .B(n31764), .Z(n23671) );
  XOR U32345 ( .A(n31768), .B(n31769), .Z(n31764) );
  NOR U32346 ( .A(n23673), .B(n23672), .Z(n31768) );
  XOR U32347 ( .A(n31770), .B(n31771), .Z(n23672) );
  XNOR U32348 ( .A(n31772), .B(n31769), .Z(n31771) );
  XOR U32349 ( .A(sreg[162]), .B(n31769), .Z(n23673) );
  XOR U32350 ( .A(n31773), .B(n31774), .Z(n31769) );
  NOR U32351 ( .A(n23675), .B(n23674), .Z(n31773) );
  XOR U32352 ( .A(n31775), .B(n31776), .Z(n23674) );
  XNOR U32353 ( .A(n31777), .B(n31774), .Z(n31776) );
  XOR U32354 ( .A(sreg[161]), .B(n31774), .Z(n23675) );
  XOR U32355 ( .A(n31778), .B(n31779), .Z(n31774) );
  NOR U32356 ( .A(n23677), .B(n23676), .Z(n31778) );
  XOR U32357 ( .A(n31780), .B(n31781), .Z(n23676) );
  XNOR U32358 ( .A(n31782), .B(n31779), .Z(n31781) );
  XOR U32359 ( .A(sreg[160]), .B(n31779), .Z(n23677) );
  XOR U32360 ( .A(n31783), .B(n31784), .Z(n31779) );
  NOR U32361 ( .A(n23679), .B(n23678), .Z(n31783) );
  XOR U32362 ( .A(n31785), .B(n31786), .Z(n23678) );
  XNOR U32363 ( .A(n31787), .B(n31784), .Z(n31786) );
  XOR U32364 ( .A(sreg[159]), .B(n31784), .Z(n23679) );
  XOR U32365 ( .A(n31788), .B(n31789), .Z(n31784) );
  NOR U32366 ( .A(n23681), .B(n23680), .Z(n31788) );
  XOR U32367 ( .A(n31790), .B(n31791), .Z(n23680) );
  XNOR U32368 ( .A(n31792), .B(n31789), .Z(n31791) );
  XOR U32369 ( .A(sreg[158]), .B(n31789), .Z(n23681) );
  XOR U32370 ( .A(n31793), .B(n31794), .Z(n31789) );
  NOR U32371 ( .A(n23683), .B(n23682), .Z(n31793) );
  XOR U32372 ( .A(n31795), .B(n31796), .Z(n23682) );
  XNOR U32373 ( .A(n31797), .B(n31794), .Z(n31796) );
  XOR U32374 ( .A(sreg[157]), .B(n31794), .Z(n23683) );
  XOR U32375 ( .A(n31798), .B(n31799), .Z(n31794) );
  NOR U32376 ( .A(n23685), .B(n23684), .Z(n31798) );
  XOR U32377 ( .A(n31800), .B(n31801), .Z(n23684) );
  XNOR U32378 ( .A(n31802), .B(n31799), .Z(n31801) );
  XOR U32379 ( .A(sreg[156]), .B(n31799), .Z(n23685) );
  XOR U32380 ( .A(n31803), .B(n31804), .Z(n31799) );
  NOR U32381 ( .A(n23687), .B(n23686), .Z(n31803) );
  XOR U32382 ( .A(n31805), .B(n31806), .Z(n23686) );
  XNOR U32383 ( .A(n31807), .B(n31804), .Z(n31806) );
  XOR U32384 ( .A(sreg[155]), .B(n31804), .Z(n23687) );
  XOR U32385 ( .A(n31808), .B(n31809), .Z(n31804) );
  NOR U32386 ( .A(n23689), .B(n23688), .Z(n31808) );
  XOR U32387 ( .A(n31810), .B(n31811), .Z(n23688) );
  XNOR U32388 ( .A(n31812), .B(n31809), .Z(n31811) );
  XOR U32389 ( .A(sreg[154]), .B(n31809), .Z(n23689) );
  XOR U32390 ( .A(n31813), .B(n31814), .Z(n31809) );
  NOR U32391 ( .A(n23691), .B(n23690), .Z(n31813) );
  XOR U32392 ( .A(n31815), .B(n31816), .Z(n23690) );
  XNOR U32393 ( .A(n31817), .B(n31814), .Z(n31816) );
  XOR U32394 ( .A(sreg[153]), .B(n31814), .Z(n23691) );
  XOR U32395 ( .A(n31818), .B(n31819), .Z(n31814) );
  NOR U32396 ( .A(n23693), .B(n23692), .Z(n31818) );
  XOR U32397 ( .A(n31820), .B(n31821), .Z(n23692) );
  XNOR U32398 ( .A(n31822), .B(n31819), .Z(n31821) );
  XOR U32399 ( .A(sreg[152]), .B(n31819), .Z(n23693) );
  XOR U32400 ( .A(n31823), .B(n31824), .Z(n31819) );
  NOR U32401 ( .A(n23695), .B(n23694), .Z(n31823) );
  XOR U32402 ( .A(n31825), .B(n31826), .Z(n23694) );
  XNOR U32403 ( .A(n31827), .B(n31824), .Z(n31826) );
  XOR U32404 ( .A(sreg[151]), .B(n31824), .Z(n23695) );
  XOR U32405 ( .A(n31828), .B(n31829), .Z(n31824) );
  NOR U32406 ( .A(n23697), .B(n23696), .Z(n31828) );
  XOR U32407 ( .A(n31830), .B(n31831), .Z(n23696) );
  XNOR U32408 ( .A(n31832), .B(n31829), .Z(n31831) );
  XOR U32409 ( .A(sreg[150]), .B(n31829), .Z(n23697) );
  XOR U32410 ( .A(n31833), .B(n31834), .Z(n31829) );
  NOR U32411 ( .A(n23699), .B(n23698), .Z(n31833) );
  XOR U32412 ( .A(n31835), .B(n31836), .Z(n23698) );
  XNOR U32413 ( .A(n31837), .B(n31834), .Z(n31836) );
  XOR U32414 ( .A(sreg[149]), .B(n31834), .Z(n23699) );
  XOR U32415 ( .A(n31838), .B(n31839), .Z(n31834) );
  NOR U32416 ( .A(n23701), .B(n23700), .Z(n31838) );
  XOR U32417 ( .A(n31840), .B(n31841), .Z(n23700) );
  XNOR U32418 ( .A(n31842), .B(n31839), .Z(n31841) );
  XOR U32419 ( .A(sreg[148]), .B(n31839), .Z(n23701) );
  XOR U32420 ( .A(n31843), .B(n31844), .Z(n31839) );
  NOR U32421 ( .A(n23703), .B(n23702), .Z(n31843) );
  XOR U32422 ( .A(n31845), .B(n31846), .Z(n23702) );
  XNOR U32423 ( .A(n31847), .B(n31844), .Z(n31846) );
  XOR U32424 ( .A(sreg[147]), .B(n31844), .Z(n23703) );
  XOR U32425 ( .A(n31848), .B(n31849), .Z(n31844) );
  NOR U32426 ( .A(n23705), .B(n23704), .Z(n31848) );
  XOR U32427 ( .A(n31850), .B(n31851), .Z(n23704) );
  XNOR U32428 ( .A(n31852), .B(n31849), .Z(n31851) );
  XOR U32429 ( .A(sreg[146]), .B(n31849), .Z(n23705) );
  XOR U32430 ( .A(n31853), .B(n31854), .Z(n31849) );
  NOR U32431 ( .A(n23707), .B(n23706), .Z(n31853) );
  XOR U32432 ( .A(n31855), .B(n31856), .Z(n23706) );
  XNOR U32433 ( .A(n31857), .B(n31854), .Z(n31856) );
  XOR U32434 ( .A(sreg[145]), .B(n31854), .Z(n23707) );
  XOR U32435 ( .A(n31858), .B(n31859), .Z(n31854) );
  NOR U32436 ( .A(n23709), .B(n23708), .Z(n31858) );
  XOR U32437 ( .A(n31860), .B(n31861), .Z(n23708) );
  XNOR U32438 ( .A(n31862), .B(n31859), .Z(n31861) );
  XOR U32439 ( .A(sreg[144]), .B(n31859), .Z(n23709) );
  XOR U32440 ( .A(n31863), .B(n31864), .Z(n31859) );
  NOR U32441 ( .A(n23711), .B(n23710), .Z(n31863) );
  XOR U32442 ( .A(n31865), .B(n31866), .Z(n23710) );
  XNOR U32443 ( .A(n31867), .B(n31864), .Z(n31866) );
  XOR U32444 ( .A(sreg[143]), .B(n31864), .Z(n23711) );
  XOR U32445 ( .A(n31868), .B(n31869), .Z(n31864) );
  NOR U32446 ( .A(n23713), .B(n23712), .Z(n31868) );
  XOR U32447 ( .A(n31870), .B(n31871), .Z(n23712) );
  XNOR U32448 ( .A(n31872), .B(n31869), .Z(n31871) );
  XOR U32449 ( .A(sreg[142]), .B(n31869), .Z(n23713) );
  XOR U32450 ( .A(n31873), .B(n31874), .Z(n31869) );
  NOR U32451 ( .A(n23715), .B(n23714), .Z(n31873) );
  XOR U32452 ( .A(n31875), .B(n31876), .Z(n23714) );
  XNOR U32453 ( .A(n31877), .B(n31874), .Z(n31876) );
  XOR U32454 ( .A(sreg[141]), .B(n31874), .Z(n23715) );
  XOR U32455 ( .A(n31878), .B(n31879), .Z(n31874) );
  NOR U32456 ( .A(n23717), .B(n23716), .Z(n31878) );
  XOR U32457 ( .A(n31880), .B(n31881), .Z(n23716) );
  XNOR U32458 ( .A(n31882), .B(n31879), .Z(n31881) );
  XOR U32459 ( .A(sreg[140]), .B(n31879), .Z(n23717) );
  XOR U32460 ( .A(n31883), .B(n31884), .Z(n31879) );
  NOR U32461 ( .A(n23719), .B(n23718), .Z(n31883) );
  XOR U32462 ( .A(n31885), .B(n31886), .Z(n23718) );
  XNOR U32463 ( .A(n31887), .B(n31884), .Z(n31886) );
  XOR U32464 ( .A(sreg[139]), .B(n31884), .Z(n23719) );
  XOR U32465 ( .A(n31888), .B(n31889), .Z(n31884) );
  NOR U32466 ( .A(n23721), .B(n23720), .Z(n31888) );
  XOR U32467 ( .A(n31890), .B(n31891), .Z(n23720) );
  XNOR U32468 ( .A(n31892), .B(n31889), .Z(n31891) );
  XOR U32469 ( .A(sreg[138]), .B(n31889), .Z(n23721) );
  XOR U32470 ( .A(n31893), .B(n31894), .Z(n31889) );
  NOR U32471 ( .A(n23723), .B(n23722), .Z(n31893) );
  XOR U32472 ( .A(n31895), .B(n31896), .Z(n23722) );
  XNOR U32473 ( .A(n31897), .B(n31894), .Z(n31896) );
  XOR U32474 ( .A(sreg[137]), .B(n31894), .Z(n23723) );
  XOR U32475 ( .A(n31898), .B(n31899), .Z(n31894) );
  NOR U32476 ( .A(n23725), .B(n23724), .Z(n31898) );
  XOR U32477 ( .A(n31900), .B(n31901), .Z(n23724) );
  XNOR U32478 ( .A(n31902), .B(n31899), .Z(n31901) );
  XOR U32479 ( .A(sreg[136]), .B(n31899), .Z(n23725) );
  XOR U32480 ( .A(n31903), .B(n31904), .Z(n31899) );
  NOR U32481 ( .A(n23727), .B(n23726), .Z(n31903) );
  XOR U32482 ( .A(n31905), .B(n31906), .Z(n23726) );
  XNOR U32483 ( .A(n31907), .B(n31904), .Z(n31906) );
  XOR U32484 ( .A(sreg[135]), .B(n31904), .Z(n23727) );
  XOR U32485 ( .A(n31908), .B(n31909), .Z(n31904) );
  NOR U32486 ( .A(n23729), .B(n23728), .Z(n31908) );
  XOR U32487 ( .A(n31910), .B(n31911), .Z(n23728) );
  XNOR U32488 ( .A(n31912), .B(n31909), .Z(n31911) );
  XOR U32489 ( .A(sreg[134]), .B(n31909), .Z(n23729) );
  XOR U32490 ( .A(n31913), .B(n31914), .Z(n31909) );
  NOR U32491 ( .A(n23731), .B(n23730), .Z(n31913) );
  XOR U32492 ( .A(n31915), .B(n31916), .Z(n23730) );
  XNOR U32493 ( .A(n31917), .B(n31914), .Z(n31916) );
  XOR U32494 ( .A(sreg[133]), .B(n31914), .Z(n23731) );
  XOR U32495 ( .A(n31918), .B(n31919), .Z(n31914) );
  NOR U32496 ( .A(n23733), .B(n23732), .Z(n31918) );
  XOR U32497 ( .A(n31920), .B(n31921), .Z(n23732) );
  XNOR U32498 ( .A(n31922), .B(n31919), .Z(n31921) );
  XOR U32499 ( .A(sreg[132]), .B(n31919), .Z(n23733) );
  XOR U32500 ( .A(n31923), .B(n31924), .Z(n31919) );
  NOR U32501 ( .A(n23735), .B(n23734), .Z(n31923) );
  XOR U32502 ( .A(n31925), .B(n31926), .Z(n23734) );
  XNOR U32503 ( .A(n31927), .B(n31924), .Z(n31926) );
  XOR U32504 ( .A(sreg[131]), .B(n31924), .Z(n23735) );
  XOR U32505 ( .A(n31928), .B(n31929), .Z(n31924) );
  NOR U32506 ( .A(n23737), .B(n23736), .Z(n31928) );
  XOR U32507 ( .A(n31930), .B(n31931), .Z(n23736) );
  XOR U32508 ( .A(sreg[130]), .B(n31929), .Z(n23737) );
  XOR U32509 ( .A(n31933), .B(n31934), .Z(n31929) );
  NAND U32510 ( .A(n23738), .B(n23739), .Z(n31934) );
  XOR U32511 ( .A(sreg[129]), .B(n31933), .Z(n23739) );
  XNOR U32512 ( .A(n31933), .B(n31935), .Z(n23738) );
  XNOR U32513 ( .A(n31936), .B(n31937), .Z(n31935) );
  ANDN U32514 ( .B(sreg[128]), .A(n23740), .Z(n31933) );
  NAND U32515 ( .A(b[0]), .B(a[0]), .Z(n23740) );
  NAND U32516 ( .A(a[36]), .B(b[0]), .Z(n31551) );
  XNOR U32517 ( .A(n31755), .B(n31756), .Z(n31552) );
  XOR U32518 ( .A(n31753), .B(n31938), .Z(n31756) );
  NAND U32519 ( .A(b[1]), .B(a[35]), .Z(n31938) );
  XOR U32520 ( .A(n31761), .B(n31939), .Z(n31755) );
  XOR U32521 ( .A(n31753), .B(n31760), .Z(n31939) );
  XNOR U32522 ( .A(n31940), .B(n31759), .Z(n31760) );
  AND U32523 ( .A(b[2]), .B(a[34]), .Z(n31940) );
  NANDN U32524 ( .A(n31767), .B(n31765), .Z(n31753) );
  XNOR U32525 ( .A(n31941), .B(n31942), .Z(n31765) );
  NAND U32526 ( .A(a[35]), .B(b[0]), .Z(n31767) );
  XOR U32527 ( .A(n31759), .B(n31751), .Z(n31943) );
  XNOR U32528 ( .A(n31750), .B(n31746), .Z(n31944) );
  XNOR U32529 ( .A(n31745), .B(n31741), .Z(n31945) );
  XNOR U32530 ( .A(n31740), .B(n31736), .Z(n31946) );
  XNOR U32531 ( .A(n31735), .B(n31731), .Z(n31947) );
  XNOR U32532 ( .A(n31730), .B(n31726), .Z(n31948) );
  XNOR U32533 ( .A(n31725), .B(n31721), .Z(n31949) );
  XNOR U32534 ( .A(n31720), .B(n31716), .Z(n31950) );
  XNOR U32535 ( .A(n31715), .B(n31711), .Z(n31951) );
  XNOR U32536 ( .A(n31710), .B(n31706), .Z(n31952) );
  XNOR U32537 ( .A(n31705), .B(n31701), .Z(n31953) );
  XNOR U32538 ( .A(n31700), .B(n31696), .Z(n31954) );
  XNOR U32539 ( .A(n31695), .B(n31691), .Z(n31955) );
  XNOR U32540 ( .A(n31690), .B(n31686), .Z(n31956) );
  XNOR U32541 ( .A(n31685), .B(n31681), .Z(n31957) );
  XNOR U32542 ( .A(n31680), .B(n31676), .Z(n31958) );
  XNOR U32543 ( .A(n31675), .B(n31671), .Z(n31959) );
  XNOR U32544 ( .A(n31670), .B(n31666), .Z(n31960) );
  XNOR U32545 ( .A(n31665), .B(n31661), .Z(n31961) );
  XNOR U32546 ( .A(n31660), .B(n31656), .Z(n31962) );
  XNOR U32547 ( .A(n31655), .B(n31651), .Z(n31963) );
  XNOR U32548 ( .A(n31650), .B(n31646), .Z(n31964) );
  XNOR U32549 ( .A(n31645), .B(n31641), .Z(n31965) );
  XNOR U32550 ( .A(n31640), .B(n31636), .Z(n31966) );
  XNOR U32551 ( .A(n31635), .B(n31631), .Z(n31967) );
  XNOR U32552 ( .A(n31630), .B(n31626), .Z(n31968) );
  XNOR U32553 ( .A(n31625), .B(n31621), .Z(n31969) );
  XNOR U32554 ( .A(n31620), .B(n31616), .Z(n31970) );
  XNOR U32555 ( .A(n31615), .B(n31611), .Z(n31971) );
  XNOR U32556 ( .A(n31610), .B(n31606), .Z(n31972) );
  XNOR U32557 ( .A(n31605), .B(n31601), .Z(n31973) );
  XNOR U32558 ( .A(n31600), .B(n31596), .Z(n31974) );
  XNOR U32559 ( .A(n31595), .B(n31591), .Z(n31975) );
  XNOR U32560 ( .A(n31976), .B(n31590), .Z(n31591) );
  AND U32561 ( .A(a[0]), .B(b[36]), .Z(n31976) );
  XNOR U32562 ( .A(n31977), .B(n31590), .Z(n31592) );
  XNOR U32563 ( .A(n31978), .B(n31979), .Z(n31590) );
  AND U32564 ( .A(n31980), .B(n31981), .Z(n31978) );
  AND U32565 ( .A(a[1]), .B(b[35]), .Z(n31977) );
  XOR U32566 ( .A(n31982), .B(n31595), .Z(n31597) );
  XOR U32567 ( .A(n31983), .B(n31984), .Z(n31595) );
  AND U32568 ( .A(n31985), .B(n31986), .Z(n31983) );
  AND U32569 ( .A(a[2]), .B(b[34]), .Z(n31982) );
  XOR U32570 ( .A(n31987), .B(n31600), .Z(n31602) );
  XOR U32571 ( .A(n31988), .B(n31989), .Z(n31600) );
  AND U32572 ( .A(n31990), .B(n31991), .Z(n31988) );
  AND U32573 ( .A(a[3]), .B(b[33]), .Z(n31987) );
  XOR U32574 ( .A(n31992), .B(n31605), .Z(n31607) );
  XOR U32575 ( .A(n31993), .B(n31994), .Z(n31605) );
  AND U32576 ( .A(n31995), .B(n31996), .Z(n31993) );
  AND U32577 ( .A(a[4]), .B(b[32]), .Z(n31992) );
  XOR U32578 ( .A(n31997), .B(n31610), .Z(n31612) );
  XOR U32579 ( .A(n31998), .B(n31999), .Z(n31610) );
  AND U32580 ( .A(n32000), .B(n32001), .Z(n31998) );
  AND U32581 ( .A(a[5]), .B(b[31]), .Z(n31997) );
  XOR U32582 ( .A(n32002), .B(n31615), .Z(n31617) );
  XOR U32583 ( .A(n32003), .B(n32004), .Z(n31615) );
  AND U32584 ( .A(n32005), .B(n32006), .Z(n32003) );
  AND U32585 ( .A(a[6]), .B(b[30]), .Z(n32002) );
  XOR U32586 ( .A(n32007), .B(n31620), .Z(n31622) );
  XOR U32587 ( .A(n32008), .B(n32009), .Z(n31620) );
  AND U32588 ( .A(n32010), .B(n32011), .Z(n32008) );
  AND U32589 ( .A(a[7]), .B(b[29]), .Z(n32007) );
  XOR U32590 ( .A(n32012), .B(n31625), .Z(n31627) );
  XOR U32591 ( .A(n32013), .B(n32014), .Z(n31625) );
  AND U32592 ( .A(n32015), .B(n32016), .Z(n32013) );
  AND U32593 ( .A(a[8]), .B(b[28]), .Z(n32012) );
  XOR U32594 ( .A(n32017), .B(n31630), .Z(n31632) );
  XOR U32595 ( .A(n32018), .B(n32019), .Z(n31630) );
  AND U32596 ( .A(n32020), .B(n32021), .Z(n32018) );
  AND U32597 ( .A(a[9]), .B(b[27]), .Z(n32017) );
  XOR U32598 ( .A(n32022), .B(n31635), .Z(n31637) );
  XOR U32599 ( .A(n32023), .B(n32024), .Z(n31635) );
  AND U32600 ( .A(n32025), .B(n32026), .Z(n32023) );
  AND U32601 ( .A(a[10]), .B(b[26]), .Z(n32022) );
  XOR U32602 ( .A(n32027), .B(n31640), .Z(n31642) );
  XOR U32603 ( .A(n32028), .B(n32029), .Z(n31640) );
  AND U32604 ( .A(n32030), .B(n32031), .Z(n32028) );
  AND U32605 ( .A(a[11]), .B(b[25]), .Z(n32027) );
  XOR U32606 ( .A(n32032), .B(n31645), .Z(n31647) );
  XOR U32607 ( .A(n32033), .B(n32034), .Z(n31645) );
  AND U32608 ( .A(n32035), .B(n32036), .Z(n32033) );
  AND U32609 ( .A(a[12]), .B(b[24]), .Z(n32032) );
  XOR U32610 ( .A(n32037), .B(n31650), .Z(n31652) );
  XOR U32611 ( .A(n32038), .B(n32039), .Z(n31650) );
  AND U32612 ( .A(n32040), .B(n32041), .Z(n32038) );
  AND U32613 ( .A(a[13]), .B(b[23]), .Z(n32037) );
  XOR U32614 ( .A(n32042), .B(n31655), .Z(n31657) );
  XOR U32615 ( .A(n32043), .B(n32044), .Z(n31655) );
  AND U32616 ( .A(n32045), .B(n32046), .Z(n32043) );
  AND U32617 ( .A(a[14]), .B(b[22]), .Z(n32042) );
  XOR U32618 ( .A(n32047), .B(n31660), .Z(n31662) );
  XOR U32619 ( .A(n32048), .B(n32049), .Z(n31660) );
  AND U32620 ( .A(n32050), .B(n32051), .Z(n32048) );
  AND U32621 ( .A(a[15]), .B(b[21]), .Z(n32047) );
  XOR U32622 ( .A(n32052), .B(n31665), .Z(n31667) );
  XOR U32623 ( .A(n32053), .B(n32054), .Z(n31665) );
  AND U32624 ( .A(n32055), .B(n32056), .Z(n32053) );
  AND U32625 ( .A(a[16]), .B(b[20]), .Z(n32052) );
  XOR U32626 ( .A(n32057), .B(n31670), .Z(n31672) );
  XOR U32627 ( .A(n32058), .B(n32059), .Z(n31670) );
  AND U32628 ( .A(n32060), .B(n32061), .Z(n32058) );
  AND U32629 ( .A(a[17]), .B(b[19]), .Z(n32057) );
  XOR U32630 ( .A(n32062), .B(n31675), .Z(n31677) );
  XOR U32631 ( .A(n32063), .B(n32064), .Z(n31675) );
  AND U32632 ( .A(n32065), .B(n32066), .Z(n32063) );
  AND U32633 ( .A(a[18]), .B(b[18]), .Z(n32062) );
  XOR U32634 ( .A(n32067), .B(n31680), .Z(n31682) );
  XOR U32635 ( .A(n32068), .B(n32069), .Z(n31680) );
  AND U32636 ( .A(n32070), .B(n32071), .Z(n32068) );
  AND U32637 ( .A(b[17]), .B(a[19]), .Z(n32067) );
  XOR U32638 ( .A(n32072), .B(n31685), .Z(n31687) );
  XOR U32639 ( .A(n32073), .B(n32074), .Z(n31685) );
  AND U32640 ( .A(n32075), .B(n32076), .Z(n32073) );
  AND U32641 ( .A(b[16]), .B(a[20]), .Z(n32072) );
  XOR U32642 ( .A(n32077), .B(n31690), .Z(n31692) );
  XOR U32643 ( .A(n32078), .B(n32079), .Z(n31690) );
  AND U32644 ( .A(n32080), .B(n32081), .Z(n32078) );
  AND U32645 ( .A(b[15]), .B(a[21]), .Z(n32077) );
  XOR U32646 ( .A(n32082), .B(n31695), .Z(n31697) );
  XOR U32647 ( .A(n32083), .B(n32084), .Z(n31695) );
  AND U32648 ( .A(n32085), .B(n32086), .Z(n32083) );
  AND U32649 ( .A(b[14]), .B(a[22]), .Z(n32082) );
  XOR U32650 ( .A(n32087), .B(n31700), .Z(n31702) );
  XOR U32651 ( .A(n32088), .B(n32089), .Z(n31700) );
  AND U32652 ( .A(n32090), .B(n32091), .Z(n32088) );
  AND U32653 ( .A(b[13]), .B(a[23]), .Z(n32087) );
  XOR U32654 ( .A(n32092), .B(n31705), .Z(n31707) );
  XOR U32655 ( .A(n32093), .B(n32094), .Z(n31705) );
  AND U32656 ( .A(n32095), .B(n32096), .Z(n32093) );
  AND U32657 ( .A(b[12]), .B(a[24]), .Z(n32092) );
  XOR U32658 ( .A(n32097), .B(n31710), .Z(n31712) );
  XOR U32659 ( .A(n32098), .B(n32099), .Z(n31710) );
  AND U32660 ( .A(n32100), .B(n32101), .Z(n32098) );
  AND U32661 ( .A(b[11]), .B(a[25]), .Z(n32097) );
  XOR U32662 ( .A(n32102), .B(n31715), .Z(n31717) );
  XOR U32663 ( .A(n32103), .B(n32104), .Z(n31715) );
  AND U32664 ( .A(n32105), .B(n32106), .Z(n32103) );
  AND U32665 ( .A(b[10]), .B(a[26]), .Z(n32102) );
  XOR U32666 ( .A(n32107), .B(n31720), .Z(n31722) );
  XOR U32667 ( .A(n32108), .B(n32109), .Z(n31720) );
  AND U32668 ( .A(n32110), .B(n32111), .Z(n32108) );
  AND U32669 ( .A(b[9]), .B(a[27]), .Z(n32107) );
  XOR U32670 ( .A(n32112), .B(n31725), .Z(n31727) );
  XOR U32671 ( .A(n32113), .B(n32114), .Z(n31725) );
  AND U32672 ( .A(n32115), .B(n32116), .Z(n32113) );
  AND U32673 ( .A(b[8]), .B(a[28]), .Z(n32112) );
  XOR U32674 ( .A(n32117), .B(n31730), .Z(n31732) );
  XOR U32675 ( .A(n32118), .B(n32119), .Z(n31730) );
  AND U32676 ( .A(n32120), .B(n32121), .Z(n32118) );
  AND U32677 ( .A(b[7]), .B(a[29]), .Z(n32117) );
  XOR U32678 ( .A(n32122), .B(n31735), .Z(n31737) );
  XOR U32679 ( .A(n32123), .B(n32124), .Z(n31735) );
  AND U32680 ( .A(n32125), .B(n32126), .Z(n32123) );
  AND U32681 ( .A(b[6]), .B(a[30]), .Z(n32122) );
  XOR U32682 ( .A(n32127), .B(n31740), .Z(n31742) );
  XOR U32683 ( .A(n32128), .B(n32129), .Z(n31740) );
  AND U32684 ( .A(n32130), .B(n32131), .Z(n32128) );
  AND U32685 ( .A(b[5]), .B(a[31]), .Z(n32127) );
  XOR U32686 ( .A(n32132), .B(n31745), .Z(n31747) );
  XOR U32687 ( .A(n32133), .B(n32134), .Z(n31745) );
  AND U32688 ( .A(n32135), .B(n32136), .Z(n32133) );
  AND U32689 ( .A(b[4]), .B(a[32]), .Z(n32132) );
  XNOR U32690 ( .A(n32137), .B(n32138), .Z(n31759) );
  NANDN U32691 ( .A(n31941), .B(n31942), .Z(n32138) );
  XOR U32692 ( .A(n32137), .B(n32139), .Z(n31942) );
  NAND U32693 ( .A(b[1]), .B(a[34]), .Z(n32139) );
  XOR U32694 ( .A(n32140), .B(n32141), .Z(n31941) );
  XOR U32695 ( .A(n32137), .B(n32142), .Z(n32141) );
  NANDN U32696 ( .A(n31772), .B(n31770), .Z(n32137) );
  XNOR U32697 ( .A(n32143), .B(n32144), .Z(n31770) );
  NAND U32698 ( .A(a[34]), .B(b[0]), .Z(n31772) );
  XOR U32699 ( .A(n32145), .B(n31750), .Z(n31752) );
  XNOR U32700 ( .A(n32146), .B(n32147), .Z(n31750) );
  AND U32701 ( .A(n32142), .B(n32140), .Z(n32146) );
  XOR U32702 ( .A(n32147), .B(n32135), .Z(n32148) );
  XNOR U32703 ( .A(n32134), .B(n32130), .Z(n32149) );
  XNOR U32704 ( .A(n32129), .B(n32125), .Z(n32150) );
  XNOR U32705 ( .A(n32124), .B(n32120), .Z(n32151) );
  XNOR U32706 ( .A(n32119), .B(n32115), .Z(n32152) );
  XNOR U32707 ( .A(n32114), .B(n32110), .Z(n32153) );
  XNOR U32708 ( .A(n32109), .B(n32105), .Z(n32154) );
  XNOR U32709 ( .A(n32104), .B(n32100), .Z(n32155) );
  XNOR U32710 ( .A(n32099), .B(n32095), .Z(n32156) );
  XNOR U32711 ( .A(n32094), .B(n32090), .Z(n32157) );
  XNOR U32712 ( .A(n32089), .B(n32085), .Z(n32158) );
  XNOR U32713 ( .A(n32084), .B(n32080), .Z(n32159) );
  XNOR U32714 ( .A(n32079), .B(n32075), .Z(n32160) );
  XNOR U32715 ( .A(n32074), .B(n32070), .Z(n32161) );
  XNOR U32716 ( .A(n32069), .B(n32065), .Z(n32162) );
  XNOR U32717 ( .A(n32064), .B(n32060), .Z(n32163) );
  XNOR U32718 ( .A(n32059), .B(n32055), .Z(n32164) );
  XNOR U32719 ( .A(n32054), .B(n32050), .Z(n32165) );
  XNOR U32720 ( .A(n32049), .B(n32045), .Z(n32166) );
  XNOR U32721 ( .A(n32044), .B(n32040), .Z(n32167) );
  XNOR U32722 ( .A(n32039), .B(n32035), .Z(n32168) );
  XNOR U32723 ( .A(n32034), .B(n32030), .Z(n32169) );
  XNOR U32724 ( .A(n32029), .B(n32025), .Z(n32170) );
  XNOR U32725 ( .A(n32024), .B(n32020), .Z(n32171) );
  XNOR U32726 ( .A(n32019), .B(n32015), .Z(n32172) );
  XNOR U32727 ( .A(n32014), .B(n32010), .Z(n32173) );
  XNOR U32728 ( .A(n32009), .B(n32005), .Z(n32174) );
  XNOR U32729 ( .A(n32004), .B(n32000), .Z(n32175) );
  XNOR U32730 ( .A(n31999), .B(n31995), .Z(n32176) );
  XNOR U32731 ( .A(n31994), .B(n31990), .Z(n32177) );
  XNOR U32732 ( .A(n31989), .B(n31985), .Z(n32178) );
  XNOR U32733 ( .A(n31984), .B(n31980), .Z(n32179) );
  XOR U32734 ( .A(n32180), .B(n31979), .Z(n31980) );
  AND U32735 ( .A(a[0]), .B(b[35]), .Z(n32180) );
  XOR U32736 ( .A(n32181), .B(n31979), .Z(n31981) );
  XNOR U32737 ( .A(n32182), .B(n32183), .Z(n31979) );
  AND U32738 ( .A(n32184), .B(n32185), .Z(n32182) );
  AND U32739 ( .A(a[1]), .B(b[34]), .Z(n32181) );
  XOR U32740 ( .A(n32186), .B(n31984), .Z(n31986) );
  XOR U32741 ( .A(n32187), .B(n32188), .Z(n31984) );
  AND U32742 ( .A(n32189), .B(n32190), .Z(n32187) );
  AND U32743 ( .A(a[2]), .B(b[33]), .Z(n32186) );
  XOR U32744 ( .A(n32191), .B(n31989), .Z(n31991) );
  XOR U32745 ( .A(n32192), .B(n32193), .Z(n31989) );
  AND U32746 ( .A(n32194), .B(n32195), .Z(n32192) );
  AND U32747 ( .A(a[3]), .B(b[32]), .Z(n32191) );
  XOR U32748 ( .A(n32196), .B(n31994), .Z(n31996) );
  XOR U32749 ( .A(n32197), .B(n32198), .Z(n31994) );
  AND U32750 ( .A(n32199), .B(n32200), .Z(n32197) );
  AND U32751 ( .A(a[4]), .B(b[31]), .Z(n32196) );
  XOR U32752 ( .A(n32201), .B(n31999), .Z(n32001) );
  XOR U32753 ( .A(n32202), .B(n32203), .Z(n31999) );
  AND U32754 ( .A(n32204), .B(n32205), .Z(n32202) );
  AND U32755 ( .A(a[5]), .B(b[30]), .Z(n32201) );
  XOR U32756 ( .A(n32206), .B(n32004), .Z(n32006) );
  XOR U32757 ( .A(n32207), .B(n32208), .Z(n32004) );
  AND U32758 ( .A(n32209), .B(n32210), .Z(n32207) );
  AND U32759 ( .A(a[6]), .B(b[29]), .Z(n32206) );
  XOR U32760 ( .A(n32211), .B(n32009), .Z(n32011) );
  XOR U32761 ( .A(n32212), .B(n32213), .Z(n32009) );
  AND U32762 ( .A(n32214), .B(n32215), .Z(n32212) );
  AND U32763 ( .A(a[7]), .B(b[28]), .Z(n32211) );
  XOR U32764 ( .A(n32216), .B(n32014), .Z(n32016) );
  XOR U32765 ( .A(n32217), .B(n32218), .Z(n32014) );
  AND U32766 ( .A(n32219), .B(n32220), .Z(n32217) );
  AND U32767 ( .A(a[8]), .B(b[27]), .Z(n32216) );
  XOR U32768 ( .A(n32221), .B(n32019), .Z(n32021) );
  XOR U32769 ( .A(n32222), .B(n32223), .Z(n32019) );
  AND U32770 ( .A(n32224), .B(n32225), .Z(n32222) );
  AND U32771 ( .A(a[9]), .B(b[26]), .Z(n32221) );
  XOR U32772 ( .A(n32226), .B(n32024), .Z(n32026) );
  XOR U32773 ( .A(n32227), .B(n32228), .Z(n32024) );
  AND U32774 ( .A(n32229), .B(n32230), .Z(n32227) );
  AND U32775 ( .A(a[10]), .B(b[25]), .Z(n32226) );
  XOR U32776 ( .A(n32231), .B(n32029), .Z(n32031) );
  XOR U32777 ( .A(n32232), .B(n32233), .Z(n32029) );
  AND U32778 ( .A(n32234), .B(n32235), .Z(n32232) );
  AND U32779 ( .A(a[11]), .B(b[24]), .Z(n32231) );
  XOR U32780 ( .A(n32236), .B(n32034), .Z(n32036) );
  XOR U32781 ( .A(n32237), .B(n32238), .Z(n32034) );
  AND U32782 ( .A(n32239), .B(n32240), .Z(n32237) );
  AND U32783 ( .A(a[12]), .B(b[23]), .Z(n32236) );
  XOR U32784 ( .A(n32241), .B(n32039), .Z(n32041) );
  XOR U32785 ( .A(n32242), .B(n32243), .Z(n32039) );
  AND U32786 ( .A(n32244), .B(n32245), .Z(n32242) );
  AND U32787 ( .A(a[13]), .B(b[22]), .Z(n32241) );
  XOR U32788 ( .A(n32246), .B(n32044), .Z(n32046) );
  XOR U32789 ( .A(n32247), .B(n32248), .Z(n32044) );
  AND U32790 ( .A(n32249), .B(n32250), .Z(n32247) );
  AND U32791 ( .A(a[14]), .B(b[21]), .Z(n32246) );
  XOR U32792 ( .A(n32251), .B(n32049), .Z(n32051) );
  XOR U32793 ( .A(n32252), .B(n32253), .Z(n32049) );
  AND U32794 ( .A(n32254), .B(n32255), .Z(n32252) );
  AND U32795 ( .A(a[15]), .B(b[20]), .Z(n32251) );
  XOR U32796 ( .A(n32256), .B(n32054), .Z(n32056) );
  XOR U32797 ( .A(n32257), .B(n32258), .Z(n32054) );
  AND U32798 ( .A(n32259), .B(n32260), .Z(n32257) );
  AND U32799 ( .A(a[16]), .B(b[19]), .Z(n32256) );
  XOR U32800 ( .A(n32261), .B(n32059), .Z(n32061) );
  XOR U32801 ( .A(n32262), .B(n32263), .Z(n32059) );
  AND U32802 ( .A(n32264), .B(n32265), .Z(n32262) );
  AND U32803 ( .A(a[17]), .B(b[18]), .Z(n32261) );
  XOR U32804 ( .A(n32266), .B(n32064), .Z(n32066) );
  XOR U32805 ( .A(n32267), .B(n32268), .Z(n32064) );
  AND U32806 ( .A(n32269), .B(n32270), .Z(n32267) );
  AND U32807 ( .A(b[17]), .B(a[18]), .Z(n32266) );
  XOR U32808 ( .A(n32271), .B(n32069), .Z(n32071) );
  XOR U32809 ( .A(n32272), .B(n32273), .Z(n32069) );
  AND U32810 ( .A(n32274), .B(n32275), .Z(n32272) );
  AND U32811 ( .A(b[16]), .B(a[19]), .Z(n32271) );
  XOR U32812 ( .A(n32276), .B(n32074), .Z(n32076) );
  XOR U32813 ( .A(n32277), .B(n32278), .Z(n32074) );
  AND U32814 ( .A(n32279), .B(n32280), .Z(n32277) );
  AND U32815 ( .A(b[15]), .B(a[20]), .Z(n32276) );
  XOR U32816 ( .A(n32281), .B(n32079), .Z(n32081) );
  XOR U32817 ( .A(n32282), .B(n32283), .Z(n32079) );
  AND U32818 ( .A(n32284), .B(n32285), .Z(n32282) );
  AND U32819 ( .A(b[14]), .B(a[21]), .Z(n32281) );
  XOR U32820 ( .A(n32286), .B(n32084), .Z(n32086) );
  XOR U32821 ( .A(n32287), .B(n32288), .Z(n32084) );
  AND U32822 ( .A(n32289), .B(n32290), .Z(n32287) );
  AND U32823 ( .A(b[13]), .B(a[22]), .Z(n32286) );
  XOR U32824 ( .A(n32291), .B(n32089), .Z(n32091) );
  XOR U32825 ( .A(n32292), .B(n32293), .Z(n32089) );
  AND U32826 ( .A(n32294), .B(n32295), .Z(n32292) );
  AND U32827 ( .A(b[12]), .B(a[23]), .Z(n32291) );
  XOR U32828 ( .A(n32296), .B(n32094), .Z(n32096) );
  XOR U32829 ( .A(n32297), .B(n32298), .Z(n32094) );
  AND U32830 ( .A(n32299), .B(n32300), .Z(n32297) );
  AND U32831 ( .A(b[11]), .B(a[24]), .Z(n32296) );
  XOR U32832 ( .A(n32301), .B(n32099), .Z(n32101) );
  XOR U32833 ( .A(n32302), .B(n32303), .Z(n32099) );
  AND U32834 ( .A(n32304), .B(n32305), .Z(n32302) );
  AND U32835 ( .A(b[10]), .B(a[25]), .Z(n32301) );
  XOR U32836 ( .A(n32306), .B(n32104), .Z(n32106) );
  XOR U32837 ( .A(n32307), .B(n32308), .Z(n32104) );
  AND U32838 ( .A(n32309), .B(n32310), .Z(n32307) );
  AND U32839 ( .A(b[9]), .B(a[26]), .Z(n32306) );
  XOR U32840 ( .A(n32311), .B(n32109), .Z(n32111) );
  XOR U32841 ( .A(n32312), .B(n32313), .Z(n32109) );
  AND U32842 ( .A(n32314), .B(n32315), .Z(n32312) );
  AND U32843 ( .A(b[8]), .B(a[27]), .Z(n32311) );
  XOR U32844 ( .A(n32316), .B(n32114), .Z(n32116) );
  XOR U32845 ( .A(n32317), .B(n32318), .Z(n32114) );
  AND U32846 ( .A(n32319), .B(n32320), .Z(n32317) );
  AND U32847 ( .A(b[7]), .B(a[28]), .Z(n32316) );
  XOR U32848 ( .A(n32321), .B(n32119), .Z(n32121) );
  XOR U32849 ( .A(n32322), .B(n32323), .Z(n32119) );
  AND U32850 ( .A(n32324), .B(n32325), .Z(n32322) );
  AND U32851 ( .A(b[6]), .B(a[29]), .Z(n32321) );
  XOR U32852 ( .A(n32326), .B(n32124), .Z(n32126) );
  XOR U32853 ( .A(n32327), .B(n32328), .Z(n32124) );
  AND U32854 ( .A(n32329), .B(n32330), .Z(n32327) );
  AND U32855 ( .A(b[5]), .B(a[30]), .Z(n32326) );
  XOR U32856 ( .A(n32331), .B(n32129), .Z(n32131) );
  XOR U32857 ( .A(n32332), .B(n32333), .Z(n32129) );
  AND U32858 ( .A(n32334), .B(n32335), .Z(n32332) );
  AND U32859 ( .A(b[4]), .B(a[31]), .Z(n32331) );
  XOR U32860 ( .A(n32336), .B(n32134), .Z(n32136) );
  XNOR U32861 ( .A(n32337), .B(n32338), .Z(n32134) );
  AND U32862 ( .A(n32339), .B(n32340), .Z(n32337) );
  AND U32863 ( .A(b[3]), .B(a[32]), .Z(n32336) );
  XNOR U32864 ( .A(n32341), .B(n32147), .Z(n32142) );
  XNOR U32865 ( .A(n32342), .B(n32343), .Z(n32147) );
  NANDN U32866 ( .A(n32143), .B(n32144), .Z(n32343) );
  XOR U32867 ( .A(n32342), .B(n32344), .Z(n32144) );
  NAND U32868 ( .A(b[1]), .B(a[33]), .Z(n32344) );
  XOR U32869 ( .A(n32340), .B(n32345), .Z(n32143) );
  XOR U32870 ( .A(n32342), .B(n32339), .Z(n32345) );
  XNOR U32871 ( .A(n32346), .B(n32338), .Z(n32339) );
  AND U32872 ( .A(b[2]), .B(a[32]), .Z(n32346) );
  XOR U32873 ( .A(n32338), .B(n32334), .Z(n32347) );
  XNOR U32874 ( .A(n32333), .B(n32329), .Z(n32348) );
  XNOR U32875 ( .A(n32328), .B(n32324), .Z(n32349) );
  XNOR U32876 ( .A(n32323), .B(n32319), .Z(n32350) );
  XNOR U32877 ( .A(n32318), .B(n32314), .Z(n32351) );
  XNOR U32878 ( .A(n32313), .B(n32309), .Z(n32352) );
  XNOR U32879 ( .A(n32308), .B(n32304), .Z(n32353) );
  XNOR U32880 ( .A(n32303), .B(n32299), .Z(n32354) );
  XNOR U32881 ( .A(n32298), .B(n32294), .Z(n32355) );
  XNOR U32882 ( .A(n32293), .B(n32289), .Z(n32356) );
  XNOR U32883 ( .A(n32288), .B(n32284), .Z(n32357) );
  XNOR U32884 ( .A(n32283), .B(n32279), .Z(n32358) );
  XNOR U32885 ( .A(n32278), .B(n32274), .Z(n32359) );
  XNOR U32886 ( .A(n32273), .B(n32269), .Z(n32360) );
  XNOR U32887 ( .A(n32268), .B(n32264), .Z(n32361) );
  XNOR U32888 ( .A(n32263), .B(n32259), .Z(n32362) );
  XNOR U32889 ( .A(n32258), .B(n32254), .Z(n32363) );
  XNOR U32890 ( .A(n32253), .B(n32249), .Z(n32364) );
  XNOR U32891 ( .A(n32248), .B(n32244), .Z(n32365) );
  XNOR U32892 ( .A(n32243), .B(n32239), .Z(n32366) );
  XNOR U32893 ( .A(n32238), .B(n32234), .Z(n32367) );
  XNOR U32894 ( .A(n32233), .B(n32229), .Z(n32368) );
  XNOR U32895 ( .A(n32228), .B(n32224), .Z(n32369) );
  XNOR U32896 ( .A(n32223), .B(n32219), .Z(n32370) );
  XNOR U32897 ( .A(n32218), .B(n32214), .Z(n32371) );
  XNOR U32898 ( .A(n32213), .B(n32209), .Z(n32372) );
  XNOR U32899 ( .A(n32208), .B(n32204), .Z(n32373) );
  XNOR U32900 ( .A(n32203), .B(n32199), .Z(n32374) );
  XNOR U32901 ( .A(n32198), .B(n32194), .Z(n32375) );
  XNOR U32902 ( .A(n32193), .B(n32189), .Z(n32376) );
  XNOR U32903 ( .A(n32188), .B(n32184), .Z(n32377) );
  XNOR U32904 ( .A(n32378), .B(n32183), .Z(n32184) );
  AND U32905 ( .A(a[0]), .B(b[34]), .Z(n32378) );
  XNOR U32906 ( .A(n32379), .B(n32183), .Z(n32185) );
  XNOR U32907 ( .A(n32380), .B(n32381), .Z(n32183) );
  AND U32908 ( .A(n32382), .B(n32383), .Z(n32380) );
  AND U32909 ( .A(a[1]), .B(b[33]), .Z(n32379) );
  XOR U32910 ( .A(n32384), .B(n32188), .Z(n32190) );
  XOR U32911 ( .A(n32385), .B(n32386), .Z(n32188) );
  AND U32912 ( .A(n32387), .B(n32388), .Z(n32385) );
  AND U32913 ( .A(a[2]), .B(b[32]), .Z(n32384) );
  XOR U32914 ( .A(n32389), .B(n32193), .Z(n32195) );
  XOR U32915 ( .A(n32390), .B(n32391), .Z(n32193) );
  AND U32916 ( .A(n32392), .B(n32393), .Z(n32390) );
  AND U32917 ( .A(a[3]), .B(b[31]), .Z(n32389) );
  XOR U32918 ( .A(n32394), .B(n32198), .Z(n32200) );
  XOR U32919 ( .A(n32395), .B(n32396), .Z(n32198) );
  AND U32920 ( .A(n32397), .B(n32398), .Z(n32395) );
  AND U32921 ( .A(a[4]), .B(b[30]), .Z(n32394) );
  XOR U32922 ( .A(n32399), .B(n32203), .Z(n32205) );
  XOR U32923 ( .A(n32400), .B(n32401), .Z(n32203) );
  AND U32924 ( .A(n32402), .B(n32403), .Z(n32400) );
  AND U32925 ( .A(a[5]), .B(b[29]), .Z(n32399) );
  XOR U32926 ( .A(n32404), .B(n32208), .Z(n32210) );
  XOR U32927 ( .A(n32405), .B(n32406), .Z(n32208) );
  AND U32928 ( .A(n32407), .B(n32408), .Z(n32405) );
  AND U32929 ( .A(a[6]), .B(b[28]), .Z(n32404) );
  XOR U32930 ( .A(n32409), .B(n32213), .Z(n32215) );
  XOR U32931 ( .A(n32410), .B(n32411), .Z(n32213) );
  AND U32932 ( .A(n32412), .B(n32413), .Z(n32410) );
  AND U32933 ( .A(a[7]), .B(b[27]), .Z(n32409) );
  XOR U32934 ( .A(n32414), .B(n32218), .Z(n32220) );
  XOR U32935 ( .A(n32415), .B(n32416), .Z(n32218) );
  AND U32936 ( .A(n32417), .B(n32418), .Z(n32415) );
  AND U32937 ( .A(a[8]), .B(b[26]), .Z(n32414) );
  XOR U32938 ( .A(n32419), .B(n32223), .Z(n32225) );
  XOR U32939 ( .A(n32420), .B(n32421), .Z(n32223) );
  AND U32940 ( .A(n32422), .B(n32423), .Z(n32420) );
  AND U32941 ( .A(a[9]), .B(b[25]), .Z(n32419) );
  XOR U32942 ( .A(n32424), .B(n32228), .Z(n32230) );
  XOR U32943 ( .A(n32425), .B(n32426), .Z(n32228) );
  AND U32944 ( .A(n32427), .B(n32428), .Z(n32425) );
  AND U32945 ( .A(a[10]), .B(b[24]), .Z(n32424) );
  XOR U32946 ( .A(n32429), .B(n32233), .Z(n32235) );
  XOR U32947 ( .A(n32430), .B(n32431), .Z(n32233) );
  AND U32948 ( .A(n32432), .B(n32433), .Z(n32430) );
  AND U32949 ( .A(a[11]), .B(b[23]), .Z(n32429) );
  XOR U32950 ( .A(n32434), .B(n32238), .Z(n32240) );
  XOR U32951 ( .A(n32435), .B(n32436), .Z(n32238) );
  AND U32952 ( .A(n32437), .B(n32438), .Z(n32435) );
  AND U32953 ( .A(a[12]), .B(b[22]), .Z(n32434) );
  XOR U32954 ( .A(n32439), .B(n32243), .Z(n32245) );
  XOR U32955 ( .A(n32440), .B(n32441), .Z(n32243) );
  AND U32956 ( .A(n32442), .B(n32443), .Z(n32440) );
  AND U32957 ( .A(a[13]), .B(b[21]), .Z(n32439) );
  XOR U32958 ( .A(n32444), .B(n32248), .Z(n32250) );
  XOR U32959 ( .A(n32445), .B(n32446), .Z(n32248) );
  AND U32960 ( .A(n32447), .B(n32448), .Z(n32445) );
  AND U32961 ( .A(a[14]), .B(b[20]), .Z(n32444) );
  XOR U32962 ( .A(n32449), .B(n32253), .Z(n32255) );
  XOR U32963 ( .A(n32450), .B(n32451), .Z(n32253) );
  AND U32964 ( .A(n32452), .B(n32453), .Z(n32450) );
  AND U32965 ( .A(a[15]), .B(b[19]), .Z(n32449) );
  XOR U32966 ( .A(n32454), .B(n32258), .Z(n32260) );
  XOR U32967 ( .A(n32455), .B(n32456), .Z(n32258) );
  AND U32968 ( .A(n32457), .B(n32458), .Z(n32455) );
  AND U32969 ( .A(a[16]), .B(b[18]), .Z(n32454) );
  XOR U32970 ( .A(n32459), .B(n32263), .Z(n32265) );
  XOR U32971 ( .A(n32460), .B(n32461), .Z(n32263) );
  AND U32972 ( .A(n32462), .B(n32463), .Z(n32460) );
  AND U32973 ( .A(a[17]), .B(b[17]), .Z(n32459) );
  XOR U32974 ( .A(n32464), .B(n32268), .Z(n32270) );
  XOR U32975 ( .A(n32465), .B(n32466), .Z(n32268) );
  AND U32976 ( .A(n32467), .B(n32468), .Z(n32465) );
  AND U32977 ( .A(b[16]), .B(a[18]), .Z(n32464) );
  XOR U32978 ( .A(n32469), .B(n32273), .Z(n32275) );
  XOR U32979 ( .A(n32470), .B(n32471), .Z(n32273) );
  AND U32980 ( .A(n32472), .B(n32473), .Z(n32470) );
  AND U32981 ( .A(b[15]), .B(a[19]), .Z(n32469) );
  XOR U32982 ( .A(n32474), .B(n32278), .Z(n32280) );
  XOR U32983 ( .A(n32475), .B(n32476), .Z(n32278) );
  AND U32984 ( .A(n32477), .B(n32478), .Z(n32475) );
  AND U32985 ( .A(b[14]), .B(a[20]), .Z(n32474) );
  XOR U32986 ( .A(n32479), .B(n32283), .Z(n32285) );
  XOR U32987 ( .A(n32480), .B(n32481), .Z(n32283) );
  AND U32988 ( .A(n32482), .B(n32483), .Z(n32480) );
  AND U32989 ( .A(b[13]), .B(a[21]), .Z(n32479) );
  XOR U32990 ( .A(n32484), .B(n32288), .Z(n32290) );
  XOR U32991 ( .A(n32485), .B(n32486), .Z(n32288) );
  AND U32992 ( .A(n32487), .B(n32488), .Z(n32485) );
  AND U32993 ( .A(b[12]), .B(a[22]), .Z(n32484) );
  XOR U32994 ( .A(n32489), .B(n32293), .Z(n32295) );
  XOR U32995 ( .A(n32490), .B(n32491), .Z(n32293) );
  AND U32996 ( .A(n32492), .B(n32493), .Z(n32490) );
  AND U32997 ( .A(b[11]), .B(a[23]), .Z(n32489) );
  XOR U32998 ( .A(n32494), .B(n32298), .Z(n32300) );
  XOR U32999 ( .A(n32495), .B(n32496), .Z(n32298) );
  AND U33000 ( .A(n32497), .B(n32498), .Z(n32495) );
  AND U33001 ( .A(b[10]), .B(a[24]), .Z(n32494) );
  XOR U33002 ( .A(n32499), .B(n32303), .Z(n32305) );
  XOR U33003 ( .A(n32500), .B(n32501), .Z(n32303) );
  AND U33004 ( .A(n32502), .B(n32503), .Z(n32500) );
  AND U33005 ( .A(b[9]), .B(a[25]), .Z(n32499) );
  XOR U33006 ( .A(n32504), .B(n32308), .Z(n32310) );
  XOR U33007 ( .A(n32505), .B(n32506), .Z(n32308) );
  AND U33008 ( .A(n32507), .B(n32508), .Z(n32505) );
  AND U33009 ( .A(b[8]), .B(a[26]), .Z(n32504) );
  XOR U33010 ( .A(n32509), .B(n32313), .Z(n32315) );
  XOR U33011 ( .A(n32510), .B(n32511), .Z(n32313) );
  AND U33012 ( .A(n32512), .B(n32513), .Z(n32510) );
  AND U33013 ( .A(b[7]), .B(a[27]), .Z(n32509) );
  XOR U33014 ( .A(n32514), .B(n32318), .Z(n32320) );
  XOR U33015 ( .A(n32515), .B(n32516), .Z(n32318) );
  AND U33016 ( .A(n32517), .B(n32518), .Z(n32515) );
  AND U33017 ( .A(b[6]), .B(a[28]), .Z(n32514) );
  XOR U33018 ( .A(n32519), .B(n32323), .Z(n32325) );
  XOR U33019 ( .A(n32520), .B(n32521), .Z(n32323) );
  AND U33020 ( .A(n32522), .B(n32523), .Z(n32520) );
  AND U33021 ( .A(b[5]), .B(a[29]), .Z(n32519) );
  XOR U33022 ( .A(n32524), .B(n32328), .Z(n32330) );
  XOR U33023 ( .A(n32525), .B(n32526), .Z(n32328) );
  AND U33024 ( .A(n32527), .B(n32528), .Z(n32525) );
  AND U33025 ( .A(b[4]), .B(a[30]), .Z(n32524) );
  XNOR U33026 ( .A(n32529), .B(n32530), .Z(n32338) );
  NANDN U33027 ( .A(n32531), .B(n32532), .Z(n32530) );
  XOR U33028 ( .A(n32533), .B(n32333), .Z(n32335) );
  XNOR U33029 ( .A(n32534), .B(n32535), .Z(n32333) );
  AND U33030 ( .A(n32536), .B(n32537), .Z(n32534) );
  AND U33031 ( .A(b[3]), .B(a[31]), .Z(n32533) );
  NANDN U33032 ( .A(n31777), .B(n31775), .Z(n32342) );
  XNOR U33033 ( .A(n32531), .B(n32532), .Z(n31775) );
  XOR U33034 ( .A(n32529), .B(n32538), .Z(n32532) );
  NAND U33035 ( .A(b[1]), .B(a[32]), .Z(n32538) );
  XOR U33036 ( .A(n32537), .B(n32539), .Z(n32531) );
  XOR U33037 ( .A(n32529), .B(n32536), .Z(n32539) );
  XNOR U33038 ( .A(n32540), .B(n32535), .Z(n32536) );
  AND U33039 ( .A(b[2]), .B(a[31]), .Z(n32540) );
  NANDN U33040 ( .A(n31782), .B(n31780), .Z(n32529) );
  XNOR U33041 ( .A(n32541), .B(n32542), .Z(n31780) );
  NAND U33042 ( .A(a[32]), .B(b[0]), .Z(n31782) );
  XOR U33043 ( .A(n32535), .B(n32527), .Z(n32543) );
  XNOR U33044 ( .A(n32526), .B(n32522), .Z(n32544) );
  XNOR U33045 ( .A(n32521), .B(n32517), .Z(n32545) );
  XNOR U33046 ( .A(n32516), .B(n32512), .Z(n32546) );
  XNOR U33047 ( .A(n32511), .B(n32507), .Z(n32547) );
  XNOR U33048 ( .A(n32506), .B(n32502), .Z(n32548) );
  XNOR U33049 ( .A(n32501), .B(n32497), .Z(n32549) );
  XNOR U33050 ( .A(n32496), .B(n32492), .Z(n32550) );
  XNOR U33051 ( .A(n32491), .B(n32487), .Z(n32551) );
  XNOR U33052 ( .A(n32486), .B(n32482), .Z(n32552) );
  XNOR U33053 ( .A(n32481), .B(n32477), .Z(n32553) );
  XNOR U33054 ( .A(n32476), .B(n32472), .Z(n32554) );
  XNOR U33055 ( .A(n32471), .B(n32467), .Z(n32555) );
  XNOR U33056 ( .A(n32466), .B(n32462), .Z(n32556) );
  XNOR U33057 ( .A(n32461), .B(n32457), .Z(n32557) );
  XNOR U33058 ( .A(n32456), .B(n32452), .Z(n32558) );
  XNOR U33059 ( .A(n32451), .B(n32447), .Z(n32559) );
  XNOR U33060 ( .A(n32446), .B(n32442), .Z(n32560) );
  XNOR U33061 ( .A(n32441), .B(n32437), .Z(n32561) );
  XNOR U33062 ( .A(n32436), .B(n32432), .Z(n32562) );
  XNOR U33063 ( .A(n32431), .B(n32427), .Z(n32563) );
  XNOR U33064 ( .A(n32426), .B(n32422), .Z(n32564) );
  XNOR U33065 ( .A(n32421), .B(n32417), .Z(n32565) );
  XNOR U33066 ( .A(n32416), .B(n32412), .Z(n32566) );
  XNOR U33067 ( .A(n32411), .B(n32407), .Z(n32567) );
  XNOR U33068 ( .A(n32406), .B(n32402), .Z(n32568) );
  XNOR U33069 ( .A(n32401), .B(n32397), .Z(n32569) );
  XNOR U33070 ( .A(n32396), .B(n32392), .Z(n32570) );
  XNOR U33071 ( .A(n32391), .B(n32387), .Z(n32571) );
  XNOR U33072 ( .A(n32386), .B(n32382), .Z(n32572) );
  XOR U33073 ( .A(n32573), .B(n32381), .Z(n32382) );
  AND U33074 ( .A(a[0]), .B(b[33]), .Z(n32573) );
  XOR U33075 ( .A(n32574), .B(n32381), .Z(n32383) );
  XNOR U33076 ( .A(n32575), .B(n32576), .Z(n32381) );
  AND U33077 ( .A(n32577), .B(n32578), .Z(n32575) );
  AND U33078 ( .A(a[1]), .B(b[32]), .Z(n32574) );
  XOR U33079 ( .A(n32579), .B(n32386), .Z(n32388) );
  XOR U33080 ( .A(n32580), .B(n32581), .Z(n32386) );
  AND U33081 ( .A(n32582), .B(n32583), .Z(n32580) );
  AND U33082 ( .A(a[2]), .B(b[31]), .Z(n32579) );
  XOR U33083 ( .A(n32584), .B(n32391), .Z(n32393) );
  XOR U33084 ( .A(n32585), .B(n32586), .Z(n32391) );
  AND U33085 ( .A(n32587), .B(n32588), .Z(n32585) );
  AND U33086 ( .A(a[3]), .B(b[30]), .Z(n32584) );
  XOR U33087 ( .A(n32589), .B(n32396), .Z(n32398) );
  XOR U33088 ( .A(n32590), .B(n32591), .Z(n32396) );
  AND U33089 ( .A(n32592), .B(n32593), .Z(n32590) );
  AND U33090 ( .A(a[4]), .B(b[29]), .Z(n32589) );
  XOR U33091 ( .A(n32594), .B(n32401), .Z(n32403) );
  XOR U33092 ( .A(n32595), .B(n32596), .Z(n32401) );
  AND U33093 ( .A(n32597), .B(n32598), .Z(n32595) );
  AND U33094 ( .A(a[5]), .B(b[28]), .Z(n32594) );
  XOR U33095 ( .A(n32599), .B(n32406), .Z(n32408) );
  XOR U33096 ( .A(n32600), .B(n32601), .Z(n32406) );
  AND U33097 ( .A(n32602), .B(n32603), .Z(n32600) );
  AND U33098 ( .A(a[6]), .B(b[27]), .Z(n32599) );
  XOR U33099 ( .A(n32604), .B(n32411), .Z(n32413) );
  XOR U33100 ( .A(n32605), .B(n32606), .Z(n32411) );
  AND U33101 ( .A(n32607), .B(n32608), .Z(n32605) );
  AND U33102 ( .A(a[7]), .B(b[26]), .Z(n32604) );
  XOR U33103 ( .A(n32609), .B(n32416), .Z(n32418) );
  XOR U33104 ( .A(n32610), .B(n32611), .Z(n32416) );
  AND U33105 ( .A(n32612), .B(n32613), .Z(n32610) );
  AND U33106 ( .A(a[8]), .B(b[25]), .Z(n32609) );
  XOR U33107 ( .A(n32614), .B(n32421), .Z(n32423) );
  XOR U33108 ( .A(n32615), .B(n32616), .Z(n32421) );
  AND U33109 ( .A(n32617), .B(n32618), .Z(n32615) );
  AND U33110 ( .A(a[9]), .B(b[24]), .Z(n32614) );
  XOR U33111 ( .A(n32619), .B(n32426), .Z(n32428) );
  XOR U33112 ( .A(n32620), .B(n32621), .Z(n32426) );
  AND U33113 ( .A(n32622), .B(n32623), .Z(n32620) );
  AND U33114 ( .A(a[10]), .B(b[23]), .Z(n32619) );
  XOR U33115 ( .A(n32624), .B(n32431), .Z(n32433) );
  XOR U33116 ( .A(n32625), .B(n32626), .Z(n32431) );
  AND U33117 ( .A(n32627), .B(n32628), .Z(n32625) );
  AND U33118 ( .A(a[11]), .B(b[22]), .Z(n32624) );
  XOR U33119 ( .A(n32629), .B(n32436), .Z(n32438) );
  XOR U33120 ( .A(n32630), .B(n32631), .Z(n32436) );
  AND U33121 ( .A(n32632), .B(n32633), .Z(n32630) );
  AND U33122 ( .A(a[12]), .B(b[21]), .Z(n32629) );
  XOR U33123 ( .A(n32634), .B(n32441), .Z(n32443) );
  XOR U33124 ( .A(n32635), .B(n32636), .Z(n32441) );
  AND U33125 ( .A(n32637), .B(n32638), .Z(n32635) );
  AND U33126 ( .A(a[13]), .B(b[20]), .Z(n32634) );
  XOR U33127 ( .A(n32639), .B(n32446), .Z(n32448) );
  XOR U33128 ( .A(n32640), .B(n32641), .Z(n32446) );
  AND U33129 ( .A(n32642), .B(n32643), .Z(n32640) );
  AND U33130 ( .A(a[14]), .B(b[19]), .Z(n32639) );
  XOR U33131 ( .A(n32644), .B(n32451), .Z(n32453) );
  XOR U33132 ( .A(n32645), .B(n32646), .Z(n32451) );
  AND U33133 ( .A(n32647), .B(n32648), .Z(n32645) );
  AND U33134 ( .A(a[15]), .B(b[18]), .Z(n32644) );
  XOR U33135 ( .A(n32649), .B(n32456), .Z(n32458) );
  XOR U33136 ( .A(n32650), .B(n32651), .Z(n32456) );
  AND U33137 ( .A(n32652), .B(n32653), .Z(n32650) );
  AND U33138 ( .A(a[16]), .B(b[17]), .Z(n32649) );
  XOR U33139 ( .A(n32654), .B(n32461), .Z(n32463) );
  XOR U33140 ( .A(n32655), .B(n32656), .Z(n32461) );
  AND U33141 ( .A(n32657), .B(n32658), .Z(n32655) );
  AND U33142 ( .A(b[16]), .B(a[17]), .Z(n32654) );
  XOR U33143 ( .A(n32659), .B(n32466), .Z(n32468) );
  XOR U33144 ( .A(n32660), .B(n32661), .Z(n32466) );
  AND U33145 ( .A(n32662), .B(n32663), .Z(n32660) );
  AND U33146 ( .A(b[15]), .B(a[18]), .Z(n32659) );
  XOR U33147 ( .A(n32664), .B(n32471), .Z(n32473) );
  XOR U33148 ( .A(n32665), .B(n32666), .Z(n32471) );
  AND U33149 ( .A(n32667), .B(n32668), .Z(n32665) );
  AND U33150 ( .A(b[14]), .B(a[19]), .Z(n32664) );
  XOR U33151 ( .A(n32669), .B(n32476), .Z(n32478) );
  XOR U33152 ( .A(n32670), .B(n32671), .Z(n32476) );
  AND U33153 ( .A(n32672), .B(n32673), .Z(n32670) );
  AND U33154 ( .A(b[13]), .B(a[20]), .Z(n32669) );
  XOR U33155 ( .A(n32674), .B(n32481), .Z(n32483) );
  XOR U33156 ( .A(n32675), .B(n32676), .Z(n32481) );
  AND U33157 ( .A(n32677), .B(n32678), .Z(n32675) );
  AND U33158 ( .A(b[12]), .B(a[21]), .Z(n32674) );
  XOR U33159 ( .A(n32679), .B(n32486), .Z(n32488) );
  XOR U33160 ( .A(n32680), .B(n32681), .Z(n32486) );
  AND U33161 ( .A(n32682), .B(n32683), .Z(n32680) );
  AND U33162 ( .A(b[11]), .B(a[22]), .Z(n32679) );
  XOR U33163 ( .A(n32684), .B(n32491), .Z(n32493) );
  XOR U33164 ( .A(n32685), .B(n32686), .Z(n32491) );
  AND U33165 ( .A(n32687), .B(n32688), .Z(n32685) );
  AND U33166 ( .A(b[10]), .B(a[23]), .Z(n32684) );
  XOR U33167 ( .A(n32689), .B(n32496), .Z(n32498) );
  XOR U33168 ( .A(n32690), .B(n32691), .Z(n32496) );
  AND U33169 ( .A(n32692), .B(n32693), .Z(n32690) );
  AND U33170 ( .A(b[9]), .B(a[24]), .Z(n32689) );
  XOR U33171 ( .A(n32694), .B(n32501), .Z(n32503) );
  XOR U33172 ( .A(n32695), .B(n32696), .Z(n32501) );
  AND U33173 ( .A(n32697), .B(n32698), .Z(n32695) );
  AND U33174 ( .A(b[8]), .B(a[25]), .Z(n32694) );
  XOR U33175 ( .A(n32699), .B(n32506), .Z(n32508) );
  XOR U33176 ( .A(n32700), .B(n32701), .Z(n32506) );
  AND U33177 ( .A(n32702), .B(n32703), .Z(n32700) );
  AND U33178 ( .A(b[7]), .B(a[26]), .Z(n32699) );
  XOR U33179 ( .A(n32704), .B(n32511), .Z(n32513) );
  XOR U33180 ( .A(n32705), .B(n32706), .Z(n32511) );
  AND U33181 ( .A(n32707), .B(n32708), .Z(n32705) );
  AND U33182 ( .A(b[6]), .B(a[27]), .Z(n32704) );
  XOR U33183 ( .A(n32709), .B(n32516), .Z(n32518) );
  XOR U33184 ( .A(n32710), .B(n32711), .Z(n32516) );
  AND U33185 ( .A(n32712), .B(n32713), .Z(n32710) );
  AND U33186 ( .A(b[5]), .B(a[28]), .Z(n32709) );
  XOR U33187 ( .A(n32714), .B(n32521), .Z(n32523) );
  XOR U33188 ( .A(n32715), .B(n32716), .Z(n32521) );
  AND U33189 ( .A(n32717), .B(n32718), .Z(n32715) );
  AND U33190 ( .A(b[4]), .B(a[29]), .Z(n32714) );
  XNOR U33191 ( .A(n32719), .B(n32720), .Z(n32535) );
  NANDN U33192 ( .A(n32541), .B(n32542), .Z(n32720) );
  XOR U33193 ( .A(n32719), .B(n32721), .Z(n32542) );
  NAND U33194 ( .A(b[1]), .B(a[31]), .Z(n32721) );
  XOR U33195 ( .A(n32722), .B(n32723), .Z(n32541) );
  XOR U33196 ( .A(n32719), .B(n32724), .Z(n32723) );
  NANDN U33197 ( .A(n31787), .B(n31785), .Z(n32719) );
  XNOR U33198 ( .A(n32725), .B(n32726), .Z(n31785) );
  NAND U33199 ( .A(a[31]), .B(b[0]), .Z(n31787) );
  XOR U33200 ( .A(n32727), .B(n32526), .Z(n32528) );
  XNOR U33201 ( .A(n32728), .B(n32729), .Z(n32526) );
  AND U33202 ( .A(n32724), .B(n32722), .Z(n32728) );
  XOR U33203 ( .A(n32729), .B(n32717), .Z(n32730) );
  XNOR U33204 ( .A(n32716), .B(n32712), .Z(n32731) );
  XNOR U33205 ( .A(n32711), .B(n32707), .Z(n32732) );
  XNOR U33206 ( .A(n32706), .B(n32702), .Z(n32733) );
  XNOR U33207 ( .A(n32701), .B(n32697), .Z(n32734) );
  XNOR U33208 ( .A(n32696), .B(n32692), .Z(n32735) );
  XNOR U33209 ( .A(n32691), .B(n32687), .Z(n32736) );
  XNOR U33210 ( .A(n32686), .B(n32682), .Z(n32737) );
  XNOR U33211 ( .A(n32681), .B(n32677), .Z(n32738) );
  XNOR U33212 ( .A(n32676), .B(n32672), .Z(n32739) );
  XNOR U33213 ( .A(n32671), .B(n32667), .Z(n32740) );
  XNOR U33214 ( .A(n32666), .B(n32662), .Z(n32741) );
  XNOR U33215 ( .A(n32661), .B(n32657), .Z(n32742) );
  XNOR U33216 ( .A(n32656), .B(n32652), .Z(n32743) );
  XNOR U33217 ( .A(n32651), .B(n32647), .Z(n32744) );
  XNOR U33218 ( .A(n32646), .B(n32642), .Z(n32745) );
  XNOR U33219 ( .A(n32641), .B(n32637), .Z(n32746) );
  XNOR U33220 ( .A(n32636), .B(n32632), .Z(n32747) );
  XNOR U33221 ( .A(n32631), .B(n32627), .Z(n32748) );
  XNOR U33222 ( .A(n32626), .B(n32622), .Z(n32749) );
  XNOR U33223 ( .A(n32621), .B(n32617), .Z(n32750) );
  XNOR U33224 ( .A(n32616), .B(n32612), .Z(n32751) );
  XNOR U33225 ( .A(n32611), .B(n32607), .Z(n32752) );
  XNOR U33226 ( .A(n32606), .B(n32602), .Z(n32753) );
  XNOR U33227 ( .A(n32601), .B(n32597), .Z(n32754) );
  XNOR U33228 ( .A(n32596), .B(n32592), .Z(n32755) );
  XNOR U33229 ( .A(n32591), .B(n32587), .Z(n32756) );
  XNOR U33230 ( .A(n32586), .B(n32582), .Z(n32757) );
  XNOR U33231 ( .A(n32581), .B(n32577), .Z(n32758) );
  XNOR U33232 ( .A(n32759), .B(n32576), .Z(n32577) );
  AND U33233 ( .A(a[0]), .B(b[32]), .Z(n32759) );
  XNOR U33234 ( .A(n32760), .B(n32576), .Z(n32578) );
  XNOR U33235 ( .A(n32761), .B(n32762), .Z(n32576) );
  AND U33236 ( .A(n32763), .B(n32764), .Z(n32761) );
  AND U33237 ( .A(a[1]), .B(b[31]), .Z(n32760) );
  XOR U33238 ( .A(n32765), .B(n32581), .Z(n32583) );
  XOR U33239 ( .A(n32766), .B(n32767), .Z(n32581) );
  AND U33240 ( .A(n32768), .B(n32769), .Z(n32766) );
  AND U33241 ( .A(a[2]), .B(b[30]), .Z(n32765) );
  XOR U33242 ( .A(n32770), .B(n32586), .Z(n32588) );
  XOR U33243 ( .A(n32771), .B(n32772), .Z(n32586) );
  AND U33244 ( .A(n32773), .B(n32774), .Z(n32771) );
  AND U33245 ( .A(a[3]), .B(b[29]), .Z(n32770) );
  XOR U33246 ( .A(n32775), .B(n32591), .Z(n32593) );
  XOR U33247 ( .A(n32776), .B(n32777), .Z(n32591) );
  AND U33248 ( .A(n32778), .B(n32779), .Z(n32776) );
  AND U33249 ( .A(a[4]), .B(b[28]), .Z(n32775) );
  XOR U33250 ( .A(n32780), .B(n32596), .Z(n32598) );
  XOR U33251 ( .A(n32781), .B(n32782), .Z(n32596) );
  AND U33252 ( .A(n32783), .B(n32784), .Z(n32781) );
  AND U33253 ( .A(a[5]), .B(b[27]), .Z(n32780) );
  XOR U33254 ( .A(n32785), .B(n32601), .Z(n32603) );
  XOR U33255 ( .A(n32786), .B(n32787), .Z(n32601) );
  AND U33256 ( .A(n32788), .B(n32789), .Z(n32786) );
  AND U33257 ( .A(a[6]), .B(b[26]), .Z(n32785) );
  XOR U33258 ( .A(n32790), .B(n32606), .Z(n32608) );
  XOR U33259 ( .A(n32791), .B(n32792), .Z(n32606) );
  AND U33260 ( .A(n32793), .B(n32794), .Z(n32791) );
  AND U33261 ( .A(a[7]), .B(b[25]), .Z(n32790) );
  XOR U33262 ( .A(n32795), .B(n32611), .Z(n32613) );
  XOR U33263 ( .A(n32796), .B(n32797), .Z(n32611) );
  AND U33264 ( .A(n32798), .B(n32799), .Z(n32796) );
  AND U33265 ( .A(a[8]), .B(b[24]), .Z(n32795) );
  XOR U33266 ( .A(n32800), .B(n32616), .Z(n32618) );
  XOR U33267 ( .A(n32801), .B(n32802), .Z(n32616) );
  AND U33268 ( .A(n32803), .B(n32804), .Z(n32801) );
  AND U33269 ( .A(a[9]), .B(b[23]), .Z(n32800) );
  XOR U33270 ( .A(n32805), .B(n32621), .Z(n32623) );
  XOR U33271 ( .A(n32806), .B(n32807), .Z(n32621) );
  AND U33272 ( .A(n32808), .B(n32809), .Z(n32806) );
  AND U33273 ( .A(a[10]), .B(b[22]), .Z(n32805) );
  XOR U33274 ( .A(n32810), .B(n32626), .Z(n32628) );
  XOR U33275 ( .A(n32811), .B(n32812), .Z(n32626) );
  AND U33276 ( .A(n32813), .B(n32814), .Z(n32811) );
  AND U33277 ( .A(a[11]), .B(b[21]), .Z(n32810) );
  XOR U33278 ( .A(n32815), .B(n32631), .Z(n32633) );
  XOR U33279 ( .A(n32816), .B(n32817), .Z(n32631) );
  AND U33280 ( .A(n32818), .B(n32819), .Z(n32816) );
  AND U33281 ( .A(a[12]), .B(b[20]), .Z(n32815) );
  XOR U33282 ( .A(n32820), .B(n32636), .Z(n32638) );
  XOR U33283 ( .A(n32821), .B(n32822), .Z(n32636) );
  AND U33284 ( .A(n32823), .B(n32824), .Z(n32821) );
  AND U33285 ( .A(a[13]), .B(b[19]), .Z(n32820) );
  XOR U33286 ( .A(n32825), .B(n32641), .Z(n32643) );
  XOR U33287 ( .A(n32826), .B(n32827), .Z(n32641) );
  AND U33288 ( .A(n32828), .B(n32829), .Z(n32826) );
  AND U33289 ( .A(a[14]), .B(b[18]), .Z(n32825) );
  XOR U33290 ( .A(n32830), .B(n32646), .Z(n32648) );
  XOR U33291 ( .A(n32831), .B(n32832), .Z(n32646) );
  AND U33292 ( .A(n32833), .B(n32834), .Z(n32831) );
  AND U33293 ( .A(a[15]), .B(b[17]), .Z(n32830) );
  XOR U33294 ( .A(n32835), .B(n32651), .Z(n32653) );
  XOR U33295 ( .A(n32836), .B(n32837), .Z(n32651) );
  AND U33296 ( .A(n32838), .B(n32839), .Z(n32836) );
  AND U33297 ( .A(a[16]), .B(b[16]), .Z(n32835) );
  XOR U33298 ( .A(n32840), .B(n32656), .Z(n32658) );
  XOR U33299 ( .A(n32841), .B(n32842), .Z(n32656) );
  AND U33300 ( .A(n32843), .B(n32844), .Z(n32841) );
  AND U33301 ( .A(b[15]), .B(a[17]), .Z(n32840) );
  XOR U33302 ( .A(n32845), .B(n32661), .Z(n32663) );
  XOR U33303 ( .A(n32846), .B(n32847), .Z(n32661) );
  AND U33304 ( .A(n32848), .B(n32849), .Z(n32846) );
  AND U33305 ( .A(b[14]), .B(a[18]), .Z(n32845) );
  XOR U33306 ( .A(n32850), .B(n32666), .Z(n32668) );
  XOR U33307 ( .A(n32851), .B(n32852), .Z(n32666) );
  AND U33308 ( .A(n32853), .B(n32854), .Z(n32851) );
  AND U33309 ( .A(b[13]), .B(a[19]), .Z(n32850) );
  XOR U33310 ( .A(n32855), .B(n32671), .Z(n32673) );
  XOR U33311 ( .A(n32856), .B(n32857), .Z(n32671) );
  AND U33312 ( .A(n32858), .B(n32859), .Z(n32856) );
  AND U33313 ( .A(b[12]), .B(a[20]), .Z(n32855) );
  XOR U33314 ( .A(n32860), .B(n32676), .Z(n32678) );
  XOR U33315 ( .A(n32861), .B(n32862), .Z(n32676) );
  AND U33316 ( .A(n32863), .B(n32864), .Z(n32861) );
  AND U33317 ( .A(b[11]), .B(a[21]), .Z(n32860) );
  XOR U33318 ( .A(n32865), .B(n32681), .Z(n32683) );
  XOR U33319 ( .A(n32866), .B(n32867), .Z(n32681) );
  AND U33320 ( .A(n32868), .B(n32869), .Z(n32866) );
  AND U33321 ( .A(b[10]), .B(a[22]), .Z(n32865) );
  XOR U33322 ( .A(n32870), .B(n32686), .Z(n32688) );
  XOR U33323 ( .A(n32871), .B(n32872), .Z(n32686) );
  AND U33324 ( .A(n32873), .B(n32874), .Z(n32871) );
  AND U33325 ( .A(b[9]), .B(a[23]), .Z(n32870) );
  XOR U33326 ( .A(n32875), .B(n32691), .Z(n32693) );
  XOR U33327 ( .A(n32876), .B(n32877), .Z(n32691) );
  AND U33328 ( .A(n32878), .B(n32879), .Z(n32876) );
  AND U33329 ( .A(b[8]), .B(a[24]), .Z(n32875) );
  XOR U33330 ( .A(n32880), .B(n32696), .Z(n32698) );
  XOR U33331 ( .A(n32881), .B(n32882), .Z(n32696) );
  AND U33332 ( .A(n32883), .B(n32884), .Z(n32881) );
  AND U33333 ( .A(b[7]), .B(a[25]), .Z(n32880) );
  XOR U33334 ( .A(n32885), .B(n32701), .Z(n32703) );
  XOR U33335 ( .A(n32886), .B(n32887), .Z(n32701) );
  AND U33336 ( .A(n32888), .B(n32889), .Z(n32886) );
  AND U33337 ( .A(b[6]), .B(a[26]), .Z(n32885) );
  XOR U33338 ( .A(n32890), .B(n32706), .Z(n32708) );
  XOR U33339 ( .A(n32891), .B(n32892), .Z(n32706) );
  AND U33340 ( .A(n32893), .B(n32894), .Z(n32891) );
  AND U33341 ( .A(b[5]), .B(a[27]), .Z(n32890) );
  XOR U33342 ( .A(n32895), .B(n32711), .Z(n32713) );
  XOR U33343 ( .A(n32896), .B(n32897), .Z(n32711) );
  AND U33344 ( .A(n32898), .B(n32899), .Z(n32896) );
  AND U33345 ( .A(b[4]), .B(a[28]), .Z(n32895) );
  XOR U33346 ( .A(n32900), .B(n32716), .Z(n32718) );
  XNOR U33347 ( .A(n32901), .B(n32902), .Z(n32716) );
  AND U33348 ( .A(n32903), .B(n32904), .Z(n32901) );
  AND U33349 ( .A(b[3]), .B(a[29]), .Z(n32900) );
  XNOR U33350 ( .A(n32905), .B(n32729), .Z(n32724) );
  XNOR U33351 ( .A(n32906), .B(n32907), .Z(n32729) );
  NANDN U33352 ( .A(n32725), .B(n32726), .Z(n32907) );
  XOR U33353 ( .A(n32906), .B(n32908), .Z(n32726) );
  NAND U33354 ( .A(b[1]), .B(a[30]), .Z(n32908) );
  XOR U33355 ( .A(n32904), .B(n32909), .Z(n32725) );
  XOR U33356 ( .A(n32906), .B(n32903), .Z(n32909) );
  XNOR U33357 ( .A(n32910), .B(n32902), .Z(n32903) );
  AND U33358 ( .A(b[2]), .B(a[29]), .Z(n32910) );
  XOR U33359 ( .A(n32902), .B(n32898), .Z(n32911) );
  XNOR U33360 ( .A(n32897), .B(n32893), .Z(n32912) );
  XNOR U33361 ( .A(n32892), .B(n32888), .Z(n32913) );
  XNOR U33362 ( .A(n32887), .B(n32883), .Z(n32914) );
  XNOR U33363 ( .A(n32882), .B(n32878), .Z(n32915) );
  XNOR U33364 ( .A(n32877), .B(n32873), .Z(n32916) );
  XNOR U33365 ( .A(n32872), .B(n32868), .Z(n32917) );
  XNOR U33366 ( .A(n32867), .B(n32863), .Z(n32918) );
  XNOR U33367 ( .A(n32862), .B(n32858), .Z(n32919) );
  XNOR U33368 ( .A(n32857), .B(n32853), .Z(n32920) );
  XNOR U33369 ( .A(n32852), .B(n32848), .Z(n32921) );
  XNOR U33370 ( .A(n32847), .B(n32843), .Z(n32922) );
  XNOR U33371 ( .A(n32842), .B(n32838), .Z(n32923) );
  XNOR U33372 ( .A(n32837), .B(n32833), .Z(n32924) );
  XNOR U33373 ( .A(n32832), .B(n32828), .Z(n32925) );
  XNOR U33374 ( .A(n32827), .B(n32823), .Z(n32926) );
  XNOR U33375 ( .A(n32822), .B(n32818), .Z(n32927) );
  XNOR U33376 ( .A(n32817), .B(n32813), .Z(n32928) );
  XNOR U33377 ( .A(n32812), .B(n32808), .Z(n32929) );
  XNOR U33378 ( .A(n32807), .B(n32803), .Z(n32930) );
  XNOR U33379 ( .A(n32802), .B(n32798), .Z(n32931) );
  XNOR U33380 ( .A(n32797), .B(n32793), .Z(n32932) );
  XNOR U33381 ( .A(n32792), .B(n32788), .Z(n32933) );
  XNOR U33382 ( .A(n32787), .B(n32783), .Z(n32934) );
  XNOR U33383 ( .A(n32782), .B(n32778), .Z(n32935) );
  XNOR U33384 ( .A(n32777), .B(n32773), .Z(n32936) );
  XNOR U33385 ( .A(n32772), .B(n32768), .Z(n32937) );
  XNOR U33386 ( .A(n32767), .B(n32763), .Z(n32938) );
  XOR U33387 ( .A(n32939), .B(n32762), .Z(n32763) );
  AND U33388 ( .A(a[0]), .B(b[31]), .Z(n32939) );
  XOR U33389 ( .A(n32940), .B(n32762), .Z(n32764) );
  XNOR U33390 ( .A(n32941), .B(n32942), .Z(n32762) );
  AND U33391 ( .A(n32943), .B(n32944), .Z(n32941) );
  AND U33392 ( .A(a[1]), .B(b[30]), .Z(n32940) );
  XOR U33393 ( .A(n32945), .B(n32767), .Z(n32769) );
  XOR U33394 ( .A(n32946), .B(n32947), .Z(n32767) );
  AND U33395 ( .A(n32948), .B(n32949), .Z(n32946) );
  AND U33396 ( .A(a[2]), .B(b[29]), .Z(n32945) );
  XOR U33397 ( .A(n32950), .B(n32772), .Z(n32774) );
  XOR U33398 ( .A(n32951), .B(n32952), .Z(n32772) );
  AND U33399 ( .A(n32953), .B(n32954), .Z(n32951) );
  AND U33400 ( .A(a[3]), .B(b[28]), .Z(n32950) );
  XOR U33401 ( .A(n32955), .B(n32777), .Z(n32779) );
  XOR U33402 ( .A(n32956), .B(n32957), .Z(n32777) );
  AND U33403 ( .A(n32958), .B(n32959), .Z(n32956) );
  AND U33404 ( .A(a[4]), .B(b[27]), .Z(n32955) );
  XOR U33405 ( .A(n32960), .B(n32782), .Z(n32784) );
  XOR U33406 ( .A(n32961), .B(n32962), .Z(n32782) );
  AND U33407 ( .A(n32963), .B(n32964), .Z(n32961) );
  AND U33408 ( .A(a[5]), .B(b[26]), .Z(n32960) );
  XOR U33409 ( .A(n32965), .B(n32787), .Z(n32789) );
  XOR U33410 ( .A(n32966), .B(n32967), .Z(n32787) );
  AND U33411 ( .A(n32968), .B(n32969), .Z(n32966) );
  AND U33412 ( .A(a[6]), .B(b[25]), .Z(n32965) );
  XOR U33413 ( .A(n32970), .B(n32792), .Z(n32794) );
  XOR U33414 ( .A(n32971), .B(n32972), .Z(n32792) );
  AND U33415 ( .A(n32973), .B(n32974), .Z(n32971) );
  AND U33416 ( .A(a[7]), .B(b[24]), .Z(n32970) );
  XOR U33417 ( .A(n32975), .B(n32797), .Z(n32799) );
  XOR U33418 ( .A(n32976), .B(n32977), .Z(n32797) );
  AND U33419 ( .A(n32978), .B(n32979), .Z(n32976) );
  AND U33420 ( .A(a[8]), .B(b[23]), .Z(n32975) );
  XOR U33421 ( .A(n32980), .B(n32802), .Z(n32804) );
  XOR U33422 ( .A(n32981), .B(n32982), .Z(n32802) );
  AND U33423 ( .A(n32983), .B(n32984), .Z(n32981) );
  AND U33424 ( .A(a[9]), .B(b[22]), .Z(n32980) );
  XOR U33425 ( .A(n32985), .B(n32807), .Z(n32809) );
  XOR U33426 ( .A(n32986), .B(n32987), .Z(n32807) );
  AND U33427 ( .A(n32988), .B(n32989), .Z(n32986) );
  AND U33428 ( .A(a[10]), .B(b[21]), .Z(n32985) );
  XOR U33429 ( .A(n32990), .B(n32812), .Z(n32814) );
  XOR U33430 ( .A(n32991), .B(n32992), .Z(n32812) );
  AND U33431 ( .A(n32993), .B(n32994), .Z(n32991) );
  AND U33432 ( .A(a[11]), .B(b[20]), .Z(n32990) );
  XOR U33433 ( .A(n32995), .B(n32817), .Z(n32819) );
  XOR U33434 ( .A(n32996), .B(n32997), .Z(n32817) );
  AND U33435 ( .A(n32998), .B(n32999), .Z(n32996) );
  AND U33436 ( .A(a[12]), .B(b[19]), .Z(n32995) );
  XOR U33437 ( .A(n33000), .B(n32822), .Z(n32824) );
  XOR U33438 ( .A(n33001), .B(n33002), .Z(n32822) );
  AND U33439 ( .A(n33003), .B(n33004), .Z(n33001) );
  AND U33440 ( .A(a[13]), .B(b[18]), .Z(n33000) );
  XOR U33441 ( .A(n33005), .B(n32827), .Z(n32829) );
  XOR U33442 ( .A(n33006), .B(n33007), .Z(n32827) );
  AND U33443 ( .A(n33008), .B(n33009), .Z(n33006) );
  AND U33444 ( .A(a[14]), .B(b[17]), .Z(n33005) );
  XOR U33445 ( .A(n33010), .B(n32832), .Z(n32834) );
  XOR U33446 ( .A(n33011), .B(n33012), .Z(n32832) );
  AND U33447 ( .A(n33013), .B(n33014), .Z(n33011) );
  AND U33448 ( .A(a[15]), .B(b[16]), .Z(n33010) );
  XOR U33449 ( .A(n33015), .B(n32837), .Z(n32839) );
  XOR U33450 ( .A(n33016), .B(n33017), .Z(n32837) );
  AND U33451 ( .A(n33018), .B(n33019), .Z(n33016) );
  AND U33452 ( .A(b[15]), .B(a[16]), .Z(n33015) );
  XOR U33453 ( .A(n33020), .B(n32842), .Z(n32844) );
  XOR U33454 ( .A(n33021), .B(n33022), .Z(n32842) );
  AND U33455 ( .A(n33023), .B(n33024), .Z(n33021) );
  AND U33456 ( .A(b[14]), .B(a[17]), .Z(n33020) );
  XOR U33457 ( .A(n33025), .B(n32847), .Z(n32849) );
  XOR U33458 ( .A(n33026), .B(n33027), .Z(n32847) );
  AND U33459 ( .A(n33028), .B(n33029), .Z(n33026) );
  AND U33460 ( .A(b[13]), .B(a[18]), .Z(n33025) );
  XOR U33461 ( .A(n33030), .B(n32852), .Z(n32854) );
  XOR U33462 ( .A(n33031), .B(n33032), .Z(n32852) );
  AND U33463 ( .A(n33033), .B(n33034), .Z(n33031) );
  AND U33464 ( .A(b[12]), .B(a[19]), .Z(n33030) );
  XOR U33465 ( .A(n33035), .B(n32857), .Z(n32859) );
  XOR U33466 ( .A(n33036), .B(n33037), .Z(n32857) );
  AND U33467 ( .A(n33038), .B(n33039), .Z(n33036) );
  AND U33468 ( .A(b[11]), .B(a[20]), .Z(n33035) );
  XOR U33469 ( .A(n33040), .B(n32862), .Z(n32864) );
  XOR U33470 ( .A(n33041), .B(n33042), .Z(n32862) );
  AND U33471 ( .A(n33043), .B(n33044), .Z(n33041) );
  AND U33472 ( .A(b[10]), .B(a[21]), .Z(n33040) );
  XOR U33473 ( .A(n33045), .B(n32867), .Z(n32869) );
  XOR U33474 ( .A(n33046), .B(n33047), .Z(n32867) );
  AND U33475 ( .A(n33048), .B(n33049), .Z(n33046) );
  AND U33476 ( .A(b[9]), .B(a[22]), .Z(n33045) );
  XOR U33477 ( .A(n33050), .B(n32872), .Z(n32874) );
  XOR U33478 ( .A(n33051), .B(n33052), .Z(n32872) );
  AND U33479 ( .A(n33053), .B(n33054), .Z(n33051) );
  AND U33480 ( .A(b[8]), .B(a[23]), .Z(n33050) );
  XOR U33481 ( .A(n33055), .B(n32877), .Z(n32879) );
  XOR U33482 ( .A(n33056), .B(n33057), .Z(n32877) );
  AND U33483 ( .A(n33058), .B(n33059), .Z(n33056) );
  AND U33484 ( .A(b[7]), .B(a[24]), .Z(n33055) );
  XOR U33485 ( .A(n33060), .B(n32882), .Z(n32884) );
  XOR U33486 ( .A(n33061), .B(n33062), .Z(n32882) );
  AND U33487 ( .A(n33063), .B(n33064), .Z(n33061) );
  AND U33488 ( .A(b[6]), .B(a[25]), .Z(n33060) );
  XOR U33489 ( .A(n33065), .B(n32887), .Z(n32889) );
  XOR U33490 ( .A(n33066), .B(n33067), .Z(n32887) );
  AND U33491 ( .A(n33068), .B(n33069), .Z(n33066) );
  AND U33492 ( .A(b[5]), .B(a[26]), .Z(n33065) );
  XOR U33493 ( .A(n33070), .B(n32892), .Z(n32894) );
  XOR U33494 ( .A(n33071), .B(n33072), .Z(n32892) );
  AND U33495 ( .A(n33073), .B(n33074), .Z(n33071) );
  AND U33496 ( .A(b[4]), .B(a[27]), .Z(n33070) );
  XNOR U33497 ( .A(n33075), .B(n33076), .Z(n32902) );
  NANDN U33498 ( .A(n33077), .B(n33078), .Z(n33076) );
  XOR U33499 ( .A(n33079), .B(n32897), .Z(n32899) );
  XNOR U33500 ( .A(n33080), .B(n33081), .Z(n32897) );
  AND U33501 ( .A(n33082), .B(n33083), .Z(n33080) );
  AND U33502 ( .A(b[3]), .B(a[28]), .Z(n33079) );
  NANDN U33503 ( .A(n31792), .B(n31790), .Z(n32906) );
  XNOR U33504 ( .A(n33077), .B(n33078), .Z(n31790) );
  XOR U33505 ( .A(n33075), .B(n33084), .Z(n33078) );
  NAND U33506 ( .A(b[1]), .B(a[29]), .Z(n33084) );
  XOR U33507 ( .A(n33083), .B(n33085), .Z(n33077) );
  XOR U33508 ( .A(n33075), .B(n33082), .Z(n33085) );
  XNOR U33509 ( .A(n33086), .B(n33081), .Z(n33082) );
  AND U33510 ( .A(b[2]), .B(a[28]), .Z(n33086) );
  NANDN U33511 ( .A(n31797), .B(n31795), .Z(n33075) );
  XNOR U33512 ( .A(n33087), .B(n33088), .Z(n31795) );
  NAND U33513 ( .A(a[29]), .B(b[0]), .Z(n31797) );
  XOR U33514 ( .A(n33081), .B(n33073), .Z(n33089) );
  XNOR U33515 ( .A(n33072), .B(n33068), .Z(n33090) );
  XNOR U33516 ( .A(n33067), .B(n33063), .Z(n33091) );
  XNOR U33517 ( .A(n33062), .B(n33058), .Z(n33092) );
  XNOR U33518 ( .A(n33057), .B(n33053), .Z(n33093) );
  XNOR U33519 ( .A(n33052), .B(n33048), .Z(n33094) );
  XNOR U33520 ( .A(n33047), .B(n33043), .Z(n33095) );
  XNOR U33521 ( .A(n33042), .B(n33038), .Z(n33096) );
  XNOR U33522 ( .A(n33037), .B(n33033), .Z(n33097) );
  XNOR U33523 ( .A(n33032), .B(n33028), .Z(n33098) );
  XNOR U33524 ( .A(n33027), .B(n33023), .Z(n33099) );
  XNOR U33525 ( .A(n33022), .B(n33018), .Z(n33100) );
  XNOR U33526 ( .A(n33017), .B(n33013), .Z(n33101) );
  XNOR U33527 ( .A(n33012), .B(n33008), .Z(n33102) );
  XNOR U33528 ( .A(n33007), .B(n33003), .Z(n33103) );
  XNOR U33529 ( .A(n33002), .B(n32998), .Z(n33104) );
  XNOR U33530 ( .A(n32997), .B(n32993), .Z(n33105) );
  XNOR U33531 ( .A(n32992), .B(n32988), .Z(n33106) );
  XNOR U33532 ( .A(n32987), .B(n32983), .Z(n33107) );
  XNOR U33533 ( .A(n32982), .B(n32978), .Z(n33108) );
  XNOR U33534 ( .A(n32977), .B(n32973), .Z(n33109) );
  XNOR U33535 ( .A(n32972), .B(n32968), .Z(n33110) );
  XNOR U33536 ( .A(n32967), .B(n32963), .Z(n33111) );
  XNOR U33537 ( .A(n32962), .B(n32958), .Z(n33112) );
  XNOR U33538 ( .A(n32957), .B(n32953), .Z(n33113) );
  XNOR U33539 ( .A(n32952), .B(n32948), .Z(n33114) );
  XNOR U33540 ( .A(n32947), .B(n32943), .Z(n33115) );
  XNOR U33541 ( .A(n33116), .B(n32942), .Z(n32943) );
  AND U33542 ( .A(a[0]), .B(b[30]), .Z(n33116) );
  XNOR U33543 ( .A(n33117), .B(n32942), .Z(n32944) );
  XNOR U33544 ( .A(n33118), .B(n33119), .Z(n32942) );
  AND U33545 ( .A(n33120), .B(n33121), .Z(n33118) );
  AND U33546 ( .A(a[1]), .B(b[29]), .Z(n33117) );
  XOR U33547 ( .A(n33122), .B(n32947), .Z(n32949) );
  XOR U33548 ( .A(n33123), .B(n33124), .Z(n32947) );
  AND U33549 ( .A(n33125), .B(n33126), .Z(n33123) );
  AND U33550 ( .A(a[2]), .B(b[28]), .Z(n33122) );
  XOR U33551 ( .A(n33127), .B(n32952), .Z(n32954) );
  XOR U33552 ( .A(n33128), .B(n33129), .Z(n32952) );
  AND U33553 ( .A(n33130), .B(n33131), .Z(n33128) );
  AND U33554 ( .A(a[3]), .B(b[27]), .Z(n33127) );
  XOR U33555 ( .A(n33132), .B(n32957), .Z(n32959) );
  XOR U33556 ( .A(n33133), .B(n33134), .Z(n32957) );
  AND U33557 ( .A(n33135), .B(n33136), .Z(n33133) );
  AND U33558 ( .A(a[4]), .B(b[26]), .Z(n33132) );
  XOR U33559 ( .A(n33137), .B(n32962), .Z(n32964) );
  XOR U33560 ( .A(n33138), .B(n33139), .Z(n32962) );
  AND U33561 ( .A(n33140), .B(n33141), .Z(n33138) );
  AND U33562 ( .A(a[5]), .B(b[25]), .Z(n33137) );
  XOR U33563 ( .A(n33142), .B(n32967), .Z(n32969) );
  XOR U33564 ( .A(n33143), .B(n33144), .Z(n32967) );
  AND U33565 ( .A(n33145), .B(n33146), .Z(n33143) );
  AND U33566 ( .A(a[6]), .B(b[24]), .Z(n33142) );
  XOR U33567 ( .A(n33147), .B(n32972), .Z(n32974) );
  XOR U33568 ( .A(n33148), .B(n33149), .Z(n32972) );
  AND U33569 ( .A(n33150), .B(n33151), .Z(n33148) );
  AND U33570 ( .A(a[7]), .B(b[23]), .Z(n33147) );
  XOR U33571 ( .A(n33152), .B(n32977), .Z(n32979) );
  XOR U33572 ( .A(n33153), .B(n33154), .Z(n32977) );
  AND U33573 ( .A(n33155), .B(n33156), .Z(n33153) );
  AND U33574 ( .A(a[8]), .B(b[22]), .Z(n33152) );
  XOR U33575 ( .A(n33157), .B(n32982), .Z(n32984) );
  XOR U33576 ( .A(n33158), .B(n33159), .Z(n32982) );
  AND U33577 ( .A(n33160), .B(n33161), .Z(n33158) );
  AND U33578 ( .A(a[9]), .B(b[21]), .Z(n33157) );
  XOR U33579 ( .A(n33162), .B(n32987), .Z(n32989) );
  XOR U33580 ( .A(n33163), .B(n33164), .Z(n32987) );
  AND U33581 ( .A(n33165), .B(n33166), .Z(n33163) );
  AND U33582 ( .A(a[10]), .B(b[20]), .Z(n33162) );
  XOR U33583 ( .A(n33167), .B(n32992), .Z(n32994) );
  XOR U33584 ( .A(n33168), .B(n33169), .Z(n32992) );
  AND U33585 ( .A(n33170), .B(n33171), .Z(n33168) );
  AND U33586 ( .A(a[11]), .B(b[19]), .Z(n33167) );
  XOR U33587 ( .A(n33172), .B(n32997), .Z(n32999) );
  XOR U33588 ( .A(n33173), .B(n33174), .Z(n32997) );
  AND U33589 ( .A(n33175), .B(n33176), .Z(n33173) );
  AND U33590 ( .A(a[12]), .B(b[18]), .Z(n33172) );
  XOR U33591 ( .A(n33177), .B(n33002), .Z(n33004) );
  XOR U33592 ( .A(n33178), .B(n33179), .Z(n33002) );
  AND U33593 ( .A(n33180), .B(n33181), .Z(n33178) );
  AND U33594 ( .A(a[13]), .B(b[17]), .Z(n33177) );
  XOR U33595 ( .A(n33182), .B(n33007), .Z(n33009) );
  XOR U33596 ( .A(n33183), .B(n33184), .Z(n33007) );
  AND U33597 ( .A(n33185), .B(n33186), .Z(n33183) );
  AND U33598 ( .A(a[14]), .B(b[16]), .Z(n33182) );
  XOR U33599 ( .A(n33187), .B(n33012), .Z(n33014) );
  XOR U33600 ( .A(n33188), .B(n33189), .Z(n33012) );
  AND U33601 ( .A(n33190), .B(n33191), .Z(n33188) );
  AND U33602 ( .A(a[15]), .B(b[15]), .Z(n33187) );
  XOR U33603 ( .A(n33192), .B(n33017), .Z(n33019) );
  XOR U33604 ( .A(n33193), .B(n33194), .Z(n33017) );
  AND U33605 ( .A(n33195), .B(n33196), .Z(n33193) );
  AND U33606 ( .A(b[14]), .B(a[16]), .Z(n33192) );
  XOR U33607 ( .A(n33197), .B(n33022), .Z(n33024) );
  XOR U33608 ( .A(n33198), .B(n33199), .Z(n33022) );
  AND U33609 ( .A(n33200), .B(n33201), .Z(n33198) );
  AND U33610 ( .A(b[13]), .B(a[17]), .Z(n33197) );
  XOR U33611 ( .A(n33202), .B(n33027), .Z(n33029) );
  XOR U33612 ( .A(n33203), .B(n33204), .Z(n33027) );
  AND U33613 ( .A(n33205), .B(n33206), .Z(n33203) );
  AND U33614 ( .A(b[12]), .B(a[18]), .Z(n33202) );
  XOR U33615 ( .A(n33207), .B(n33032), .Z(n33034) );
  XOR U33616 ( .A(n33208), .B(n33209), .Z(n33032) );
  AND U33617 ( .A(n33210), .B(n33211), .Z(n33208) );
  AND U33618 ( .A(b[11]), .B(a[19]), .Z(n33207) );
  XOR U33619 ( .A(n33212), .B(n33037), .Z(n33039) );
  XOR U33620 ( .A(n33213), .B(n33214), .Z(n33037) );
  AND U33621 ( .A(n33215), .B(n33216), .Z(n33213) );
  AND U33622 ( .A(b[10]), .B(a[20]), .Z(n33212) );
  XOR U33623 ( .A(n33217), .B(n33042), .Z(n33044) );
  XOR U33624 ( .A(n33218), .B(n33219), .Z(n33042) );
  AND U33625 ( .A(n33220), .B(n33221), .Z(n33218) );
  AND U33626 ( .A(b[9]), .B(a[21]), .Z(n33217) );
  XOR U33627 ( .A(n33222), .B(n33047), .Z(n33049) );
  XOR U33628 ( .A(n33223), .B(n33224), .Z(n33047) );
  AND U33629 ( .A(n33225), .B(n33226), .Z(n33223) );
  AND U33630 ( .A(b[8]), .B(a[22]), .Z(n33222) );
  XOR U33631 ( .A(n33227), .B(n33052), .Z(n33054) );
  XOR U33632 ( .A(n33228), .B(n33229), .Z(n33052) );
  AND U33633 ( .A(n33230), .B(n33231), .Z(n33228) );
  AND U33634 ( .A(b[7]), .B(a[23]), .Z(n33227) );
  XOR U33635 ( .A(n33232), .B(n33057), .Z(n33059) );
  XOR U33636 ( .A(n33233), .B(n33234), .Z(n33057) );
  AND U33637 ( .A(n33235), .B(n33236), .Z(n33233) );
  AND U33638 ( .A(b[6]), .B(a[24]), .Z(n33232) );
  XOR U33639 ( .A(n33237), .B(n33062), .Z(n33064) );
  XOR U33640 ( .A(n33238), .B(n33239), .Z(n33062) );
  AND U33641 ( .A(n33240), .B(n33241), .Z(n33238) );
  AND U33642 ( .A(b[5]), .B(a[25]), .Z(n33237) );
  XOR U33643 ( .A(n33242), .B(n33067), .Z(n33069) );
  XOR U33644 ( .A(n33243), .B(n33244), .Z(n33067) );
  AND U33645 ( .A(n33245), .B(n33246), .Z(n33243) );
  AND U33646 ( .A(b[4]), .B(a[26]), .Z(n33242) );
  XNOR U33647 ( .A(n33247), .B(n33248), .Z(n33081) );
  NANDN U33648 ( .A(n33087), .B(n33088), .Z(n33248) );
  XOR U33649 ( .A(n33247), .B(n33249), .Z(n33088) );
  NAND U33650 ( .A(b[1]), .B(a[28]), .Z(n33249) );
  XOR U33651 ( .A(n33250), .B(n33251), .Z(n33087) );
  XOR U33652 ( .A(n33247), .B(n33252), .Z(n33251) );
  NANDN U33653 ( .A(n31802), .B(n31800), .Z(n33247) );
  XNOR U33654 ( .A(n33253), .B(n33254), .Z(n31800) );
  NAND U33655 ( .A(a[28]), .B(b[0]), .Z(n31802) );
  XOR U33656 ( .A(n33255), .B(n33072), .Z(n33074) );
  XNOR U33657 ( .A(n33256), .B(n33257), .Z(n33072) );
  AND U33658 ( .A(n33252), .B(n33250), .Z(n33256) );
  XOR U33659 ( .A(n33257), .B(n33245), .Z(n33258) );
  XNOR U33660 ( .A(n33244), .B(n33240), .Z(n33259) );
  XNOR U33661 ( .A(n33239), .B(n33235), .Z(n33260) );
  XNOR U33662 ( .A(n33234), .B(n33230), .Z(n33261) );
  XNOR U33663 ( .A(n33229), .B(n33225), .Z(n33262) );
  XNOR U33664 ( .A(n33224), .B(n33220), .Z(n33263) );
  XNOR U33665 ( .A(n33219), .B(n33215), .Z(n33264) );
  XNOR U33666 ( .A(n33214), .B(n33210), .Z(n33265) );
  XNOR U33667 ( .A(n33209), .B(n33205), .Z(n33266) );
  XNOR U33668 ( .A(n33204), .B(n33200), .Z(n33267) );
  XNOR U33669 ( .A(n33199), .B(n33195), .Z(n33268) );
  XNOR U33670 ( .A(n33194), .B(n33190), .Z(n33269) );
  XNOR U33671 ( .A(n33189), .B(n33185), .Z(n33270) );
  XNOR U33672 ( .A(n33184), .B(n33180), .Z(n33271) );
  XNOR U33673 ( .A(n33179), .B(n33175), .Z(n33272) );
  XNOR U33674 ( .A(n33174), .B(n33170), .Z(n33273) );
  XNOR U33675 ( .A(n33169), .B(n33165), .Z(n33274) );
  XNOR U33676 ( .A(n33164), .B(n33160), .Z(n33275) );
  XNOR U33677 ( .A(n33159), .B(n33155), .Z(n33276) );
  XNOR U33678 ( .A(n33154), .B(n33150), .Z(n33277) );
  XNOR U33679 ( .A(n33149), .B(n33145), .Z(n33278) );
  XNOR U33680 ( .A(n33144), .B(n33140), .Z(n33279) );
  XNOR U33681 ( .A(n33139), .B(n33135), .Z(n33280) );
  XNOR U33682 ( .A(n33134), .B(n33130), .Z(n33281) );
  XNOR U33683 ( .A(n33129), .B(n33125), .Z(n33282) );
  XNOR U33684 ( .A(n33124), .B(n33120), .Z(n33283) );
  XOR U33685 ( .A(n33284), .B(n33119), .Z(n33120) );
  AND U33686 ( .A(a[0]), .B(b[29]), .Z(n33284) );
  XOR U33687 ( .A(n33285), .B(n33119), .Z(n33121) );
  XNOR U33688 ( .A(n33286), .B(n33287), .Z(n33119) );
  AND U33689 ( .A(n33288), .B(n33289), .Z(n33286) );
  AND U33690 ( .A(a[1]), .B(b[28]), .Z(n33285) );
  XOR U33691 ( .A(n33290), .B(n33124), .Z(n33126) );
  XOR U33692 ( .A(n33291), .B(n33292), .Z(n33124) );
  AND U33693 ( .A(n33293), .B(n33294), .Z(n33291) );
  AND U33694 ( .A(a[2]), .B(b[27]), .Z(n33290) );
  XOR U33695 ( .A(n33295), .B(n33129), .Z(n33131) );
  XOR U33696 ( .A(n33296), .B(n33297), .Z(n33129) );
  AND U33697 ( .A(n33298), .B(n33299), .Z(n33296) );
  AND U33698 ( .A(a[3]), .B(b[26]), .Z(n33295) );
  XOR U33699 ( .A(n33300), .B(n33134), .Z(n33136) );
  XOR U33700 ( .A(n33301), .B(n33302), .Z(n33134) );
  AND U33701 ( .A(n33303), .B(n33304), .Z(n33301) );
  AND U33702 ( .A(a[4]), .B(b[25]), .Z(n33300) );
  XOR U33703 ( .A(n33305), .B(n33139), .Z(n33141) );
  XOR U33704 ( .A(n33306), .B(n33307), .Z(n33139) );
  AND U33705 ( .A(n33308), .B(n33309), .Z(n33306) );
  AND U33706 ( .A(a[5]), .B(b[24]), .Z(n33305) );
  XOR U33707 ( .A(n33310), .B(n33144), .Z(n33146) );
  XOR U33708 ( .A(n33311), .B(n33312), .Z(n33144) );
  AND U33709 ( .A(n33313), .B(n33314), .Z(n33311) );
  AND U33710 ( .A(a[6]), .B(b[23]), .Z(n33310) );
  XOR U33711 ( .A(n33315), .B(n33149), .Z(n33151) );
  XOR U33712 ( .A(n33316), .B(n33317), .Z(n33149) );
  AND U33713 ( .A(n33318), .B(n33319), .Z(n33316) );
  AND U33714 ( .A(a[7]), .B(b[22]), .Z(n33315) );
  XOR U33715 ( .A(n33320), .B(n33154), .Z(n33156) );
  XOR U33716 ( .A(n33321), .B(n33322), .Z(n33154) );
  AND U33717 ( .A(n33323), .B(n33324), .Z(n33321) );
  AND U33718 ( .A(a[8]), .B(b[21]), .Z(n33320) );
  XOR U33719 ( .A(n33325), .B(n33159), .Z(n33161) );
  XOR U33720 ( .A(n33326), .B(n33327), .Z(n33159) );
  AND U33721 ( .A(n33328), .B(n33329), .Z(n33326) );
  AND U33722 ( .A(a[9]), .B(b[20]), .Z(n33325) );
  XOR U33723 ( .A(n33330), .B(n33164), .Z(n33166) );
  XOR U33724 ( .A(n33331), .B(n33332), .Z(n33164) );
  AND U33725 ( .A(n33333), .B(n33334), .Z(n33331) );
  AND U33726 ( .A(a[10]), .B(b[19]), .Z(n33330) );
  XOR U33727 ( .A(n33335), .B(n33169), .Z(n33171) );
  XOR U33728 ( .A(n33336), .B(n33337), .Z(n33169) );
  AND U33729 ( .A(n33338), .B(n33339), .Z(n33336) );
  AND U33730 ( .A(a[11]), .B(b[18]), .Z(n33335) );
  XOR U33731 ( .A(n33340), .B(n33174), .Z(n33176) );
  XOR U33732 ( .A(n33341), .B(n33342), .Z(n33174) );
  AND U33733 ( .A(n33343), .B(n33344), .Z(n33341) );
  AND U33734 ( .A(a[12]), .B(b[17]), .Z(n33340) );
  XOR U33735 ( .A(n33345), .B(n33179), .Z(n33181) );
  XOR U33736 ( .A(n33346), .B(n33347), .Z(n33179) );
  AND U33737 ( .A(n33348), .B(n33349), .Z(n33346) );
  AND U33738 ( .A(a[13]), .B(b[16]), .Z(n33345) );
  XOR U33739 ( .A(n33350), .B(n33184), .Z(n33186) );
  XOR U33740 ( .A(n33351), .B(n33352), .Z(n33184) );
  AND U33741 ( .A(n33353), .B(n33354), .Z(n33351) );
  AND U33742 ( .A(a[14]), .B(b[15]), .Z(n33350) );
  XOR U33743 ( .A(n33355), .B(n33189), .Z(n33191) );
  XOR U33744 ( .A(n33356), .B(n33357), .Z(n33189) );
  AND U33745 ( .A(n33358), .B(n33359), .Z(n33356) );
  AND U33746 ( .A(b[14]), .B(a[15]), .Z(n33355) );
  XOR U33747 ( .A(n33360), .B(n33194), .Z(n33196) );
  XOR U33748 ( .A(n33361), .B(n33362), .Z(n33194) );
  AND U33749 ( .A(n33363), .B(n33364), .Z(n33361) );
  AND U33750 ( .A(b[13]), .B(a[16]), .Z(n33360) );
  XOR U33751 ( .A(n33365), .B(n33199), .Z(n33201) );
  XOR U33752 ( .A(n33366), .B(n33367), .Z(n33199) );
  AND U33753 ( .A(n33368), .B(n33369), .Z(n33366) );
  AND U33754 ( .A(b[12]), .B(a[17]), .Z(n33365) );
  XOR U33755 ( .A(n33370), .B(n33204), .Z(n33206) );
  XOR U33756 ( .A(n33371), .B(n33372), .Z(n33204) );
  AND U33757 ( .A(n33373), .B(n33374), .Z(n33371) );
  AND U33758 ( .A(b[11]), .B(a[18]), .Z(n33370) );
  XOR U33759 ( .A(n33375), .B(n33209), .Z(n33211) );
  XOR U33760 ( .A(n33376), .B(n33377), .Z(n33209) );
  AND U33761 ( .A(n33378), .B(n33379), .Z(n33376) );
  AND U33762 ( .A(b[10]), .B(a[19]), .Z(n33375) );
  XOR U33763 ( .A(n33380), .B(n33214), .Z(n33216) );
  XOR U33764 ( .A(n33381), .B(n33382), .Z(n33214) );
  AND U33765 ( .A(n33383), .B(n33384), .Z(n33381) );
  AND U33766 ( .A(b[9]), .B(a[20]), .Z(n33380) );
  XOR U33767 ( .A(n33385), .B(n33219), .Z(n33221) );
  XOR U33768 ( .A(n33386), .B(n33387), .Z(n33219) );
  AND U33769 ( .A(n33388), .B(n33389), .Z(n33386) );
  AND U33770 ( .A(b[8]), .B(a[21]), .Z(n33385) );
  XOR U33771 ( .A(n33390), .B(n33224), .Z(n33226) );
  XOR U33772 ( .A(n33391), .B(n33392), .Z(n33224) );
  AND U33773 ( .A(n33393), .B(n33394), .Z(n33391) );
  AND U33774 ( .A(b[7]), .B(a[22]), .Z(n33390) );
  XOR U33775 ( .A(n33395), .B(n33229), .Z(n33231) );
  XOR U33776 ( .A(n33396), .B(n33397), .Z(n33229) );
  AND U33777 ( .A(n33398), .B(n33399), .Z(n33396) );
  AND U33778 ( .A(b[6]), .B(a[23]), .Z(n33395) );
  XOR U33779 ( .A(n33400), .B(n33234), .Z(n33236) );
  XOR U33780 ( .A(n33401), .B(n33402), .Z(n33234) );
  AND U33781 ( .A(n33403), .B(n33404), .Z(n33401) );
  AND U33782 ( .A(b[5]), .B(a[24]), .Z(n33400) );
  XOR U33783 ( .A(n33405), .B(n33239), .Z(n33241) );
  XOR U33784 ( .A(n33406), .B(n33407), .Z(n33239) );
  AND U33785 ( .A(n33408), .B(n33409), .Z(n33406) );
  AND U33786 ( .A(b[4]), .B(a[25]), .Z(n33405) );
  XOR U33787 ( .A(n33410), .B(n33244), .Z(n33246) );
  XNOR U33788 ( .A(n33411), .B(n33412), .Z(n33244) );
  AND U33789 ( .A(n33413), .B(n33414), .Z(n33411) );
  AND U33790 ( .A(b[3]), .B(a[26]), .Z(n33410) );
  XNOR U33791 ( .A(n33415), .B(n33257), .Z(n33252) );
  XNOR U33792 ( .A(n33416), .B(n33417), .Z(n33257) );
  NANDN U33793 ( .A(n33253), .B(n33254), .Z(n33417) );
  XOR U33794 ( .A(n33416), .B(n33418), .Z(n33254) );
  NAND U33795 ( .A(b[1]), .B(a[27]), .Z(n33418) );
  XOR U33796 ( .A(n33414), .B(n33419), .Z(n33253) );
  XOR U33797 ( .A(n33416), .B(n33413), .Z(n33419) );
  XNOR U33798 ( .A(n33420), .B(n33412), .Z(n33413) );
  AND U33799 ( .A(b[2]), .B(a[26]), .Z(n33420) );
  XOR U33800 ( .A(n33412), .B(n33408), .Z(n33421) );
  XNOR U33801 ( .A(n33407), .B(n33403), .Z(n33422) );
  XNOR U33802 ( .A(n33402), .B(n33398), .Z(n33423) );
  XNOR U33803 ( .A(n33397), .B(n33393), .Z(n33424) );
  XNOR U33804 ( .A(n33392), .B(n33388), .Z(n33425) );
  XNOR U33805 ( .A(n33387), .B(n33383), .Z(n33426) );
  XNOR U33806 ( .A(n33382), .B(n33378), .Z(n33427) );
  XNOR U33807 ( .A(n33377), .B(n33373), .Z(n33428) );
  XNOR U33808 ( .A(n33372), .B(n33368), .Z(n33429) );
  XNOR U33809 ( .A(n33367), .B(n33363), .Z(n33430) );
  XNOR U33810 ( .A(n33362), .B(n33358), .Z(n33431) );
  XNOR U33811 ( .A(n33357), .B(n33353), .Z(n33432) );
  XNOR U33812 ( .A(n33352), .B(n33348), .Z(n33433) );
  XNOR U33813 ( .A(n33347), .B(n33343), .Z(n33434) );
  XNOR U33814 ( .A(n33342), .B(n33338), .Z(n33435) );
  XNOR U33815 ( .A(n33337), .B(n33333), .Z(n33436) );
  XNOR U33816 ( .A(n33332), .B(n33328), .Z(n33437) );
  XNOR U33817 ( .A(n33327), .B(n33323), .Z(n33438) );
  XNOR U33818 ( .A(n33322), .B(n33318), .Z(n33439) );
  XNOR U33819 ( .A(n33317), .B(n33313), .Z(n33440) );
  XNOR U33820 ( .A(n33312), .B(n33308), .Z(n33441) );
  XNOR U33821 ( .A(n33307), .B(n33303), .Z(n33442) );
  XNOR U33822 ( .A(n33302), .B(n33298), .Z(n33443) );
  XNOR U33823 ( .A(n33297), .B(n33293), .Z(n33444) );
  XNOR U33824 ( .A(n33292), .B(n33288), .Z(n33445) );
  XNOR U33825 ( .A(n33446), .B(n33287), .Z(n33288) );
  AND U33826 ( .A(a[0]), .B(b[28]), .Z(n33446) );
  XNOR U33827 ( .A(n33447), .B(n33287), .Z(n33289) );
  XNOR U33828 ( .A(n33448), .B(n33449), .Z(n33287) );
  AND U33829 ( .A(n33450), .B(n33451), .Z(n33448) );
  AND U33830 ( .A(a[1]), .B(b[27]), .Z(n33447) );
  XOR U33831 ( .A(n33452), .B(n33292), .Z(n33294) );
  XOR U33832 ( .A(n33453), .B(n33454), .Z(n33292) );
  AND U33833 ( .A(n33455), .B(n33456), .Z(n33453) );
  AND U33834 ( .A(a[2]), .B(b[26]), .Z(n33452) );
  XOR U33835 ( .A(n33457), .B(n33297), .Z(n33299) );
  XOR U33836 ( .A(n33458), .B(n33459), .Z(n33297) );
  AND U33837 ( .A(n33460), .B(n33461), .Z(n33458) );
  AND U33838 ( .A(a[3]), .B(b[25]), .Z(n33457) );
  XOR U33839 ( .A(n33462), .B(n33302), .Z(n33304) );
  XOR U33840 ( .A(n33463), .B(n33464), .Z(n33302) );
  AND U33841 ( .A(n33465), .B(n33466), .Z(n33463) );
  AND U33842 ( .A(a[4]), .B(b[24]), .Z(n33462) );
  XOR U33843 ( .A(n33467), .B(n33307), .Z(n33309) );
  XOR U33844 ( .A(n33468), .B(n33469), .Z(n33307) );
  AND U33845 ( .A(n33470), .B(n33471), .Z(n33468) );
  AND U33846 ( .A(a[5]), .B(b[23]), .Z(n33467) );
  XOR U33847 ( .A(n33472), .B(n33312), .Z(n33314) );
  XOR U33848 ( .A(n33473), .B(n33474), .Z(n33312) );
  AND U33849 ( .A(n33475), .B(n33476), .Z(n33473) );
  AND U33850 ( .A(a[6]), .B(b[22]), .Z(n33472) );
  XOR U33851 ( .A(n33477), .B(n33317), .Z(n33319) );
  XOR U33852 ( .A(n33478), .B(n33479), .Z(n33317) );
  AND U33853 ( .A(n33480), .B(n33481), .Z(n33478) );
  AND U33854 ( .A(a[7]), .B(b[21]), .Z(n33477) );
  XOR U33855 ( .A(n33482), .B(n33322), .Z(n33324) );
  XOR U33856 ( .A(n33483), .B(n33484), .Z(n33322) );
  AND U33857 ( .A(n33485), .B(n33486), .Z(n33483) );
  AND U33858 ( .A(a[8]), .B(b[20]), .Z(n33482) );
  XOR U33859 ( .A(n33487), .B(n33327), .Z(n33329) );
  XOR U33860 ( .A(n33488), .B(n33489), .Z(n33327) );
  AND U33861 ( .A(n33490), .B(n33491), .Z(n33488) );
  AND U33862 ( .A(a[9]), .B(b[19]), .Z(n33487) );
  XOR U33863 ( .A(n33492), .B(n33332), .Z(n33334) );
  XOR U33864 ( .A(n33493), .B(n33494), .Z(n33332) );
  AND U33865 ( .A(n33495), .B(n33496), .Z(n33493) );
  AND U33866 ( .A(a[10]), .B(b[18]), .Z(n33492) );
  XOR U33867 ( .A(n33497), .B(n33337), .Z(n33339) );
  XOR U33868 ( .A(n33498), .B(n33499), .Z(n33337) );
  AND U33869 ( .A(n33500), .B(n33501), .Z(n33498) );
  AND U33870 ( .A(a[11]), .B(b[17]), .Z(n33497) );
  XOR U33871 ( .A(n33502), .B(n33342), .Z(n33344) );
  XOR U33872 ( .A(n33503), .B(n33504), .Z(n33342) );
  AND U33873 ( .A(n33505), .B(n33506), .Z(n33503) );
  AND U33874 ( .A(a[12]), .B(b[16]), .Z(n33502) );
  XOR U33875 ( .A(n33507), .B(n33347), .Z(n33349) );
  XOR U33876 ( .A(n33508), .B(n33509), .Z(n33347) );
  AND U33877 ( .A(n33510), .B(n33511), .Z(n33508) );
  AND U33878 ( .A(a[13]), .B(b[15]), .Z(n33507) );
  XOR U33879 ( .A(n33512), .B(n33352), .Z(n33354) );
  XOR U33880 ( .A(n33513), .B(n33514), .Z(n33352) );
  AND U33881 ( .A(n33515), .B(n33516), .Z(n33513) );
  AND U33882 ( .A(a[14]), .B(b[14]), .Z(n33512) );
  XOR U33883 ( .A(n33517), .B(n33357), .Z(n33359) );
  XOR U33884 ( .A(n33518), .B(n33519), .Z(n33357) );
  AND U33885 ( .A(n33520), .B(n33521), .Z(n33518) );
  AND U33886 ( .A(b[13]), .B(a[15]), .Z(n33517) );
  XOR U33887 ( .A(n33522), .B(n33362), .Z(n33364) );
  XOR U33888 ( .A(n33523), .B(n33524), .Z(n33362) );
  AND U33889 ( .A(n33525), .B(n33526), .Z(n33523) );
  AND U33890 ( .A(b[12]), .B(a[16]), .Z(n33522) );
  XOR U33891 ( .A(n33527), .B(n33367), .Z(n33369) );
  XOR U33892 ( .A(n33528), .B(n33529), .Z(n33367) );
  AND U33893 ( .A(n33530), .B(n33531), .Z(n33528) );
  AND U33894 ( .A(b[11]), .B(a[17]), .Z(n33527) );
  XOR U33895 ( .A(n33532), .B(n33372), .Z(n33374) );
  XOR U33896 ( .A(n33533), .B(n33534), .Z(n33372) );
  AND U33897 ( .A(n33535), .B(n33536), .Z(n33533) );
  AND U33898 ( .A(b[10]), .B(a[18]), .Z(n33532) );
  XOR U33899 ( .A(n33537), .B(n33377), .Z(n33379) );
  XOR U33900 ( .A(n33538), .B(n33539), .Z(n33377) );
  AND U33901 ( .A(n33540), .B(n33541), .Z(n33538) );
  AND U33902 ( .A(b[9]), .B(a[19]), .Z(n33537) );
  XOR U33903 ( .A(n33542), .B(n33382), .Z(n33384) );
  XOR U33904 ( .A(n33543), .B(n33544), .Z(n33382) );
  AND U33905 ( .A(n33545), .B(n33546), .Z(n33543) );
  AND U33906 ( .A(b[8]), .B(a[20]), .Z(n33542) );
  XOR U33907 ( .A(n33547), .B(n33387), .Z(n33389) );
  XOR U33908 ( .A(n33548), .B(n33549), .Z(n33387) );
  AND U33909 ( .A(n33550), .B(n33551), .Z(n33548) );
  AND U33910 ( .A(b[7]), .B(a[21]), .Z(n33547) );
  XOR U33911 ( .A(n33552), .B(n33392), .Z(n33394) );
  XOR U33912 ( .A(n33553), .B(n33554), .Z(n33392) );
  AND U33913 ( .A(n33555), .B(n33556), .Z(n33553) );
  AND U33914 ( .A(b[6]), .B(a[22]), .Z(n33552) );
  XOR U33915 ( .A(n33557), .B(n33397), .Z(n33399) );
  XOR U33916 ( .A(n33558), .B(n33559), .Z(n33397) );
  AND U33917 ( .A(n33560), .B(n33561), .Z(n33558) );
  AND U33918 ( .A(b[5]), .B(a[23]), .Z(n33557) );
  XOR U33919 ( .A(n33562), .B(n33402), .Z(n33404) );
  XOR U33920 ( .A(n33563), .B(n33564), .Z(n33402) );
  AND U33921 ( .A(n33565), .B(n33566), .Z(n33563) );
  AND U33922 ( .A(b[4]), .B(a[24]), .Z(n33562) );
  XNOR U33923 ( .A(n33567), .B(n33568), .Z(n33412) );
  NANDN U33924 ( .A(n33569), .B(n33570), .Z(n33568) );
  XOR U33925 ( .A(n33571), .B(n33407), .Z(n33409) );
  XNOR U33926 ( .A(n33572), .B(n33573), .Z(n33407) );
  AND U33927 ( .A(n33574), .B(n33575), .Z(n33572) );
  AND U33928 ( .A(b[3]), .B(a[25]), .Z(n33571) );
  NANDN U33929 ( .A(n31807), .B(n31805), .Z(n33416) );
  XNOR U33930 ( .A(n33569), .B(n33570), .Z(n31805) );
  XOR U33931 ( .A(n33567), .B(n33576), .Z(n33570) );
  NAND U33932 ( .A(b[1]), .B(a[26]), .Z(n33576) );
  XOR U33933 ( .A(n33575), .B(n33577), .Z(n33569) );
  XOR U33934 ( .A(n33567), .B(n33574), .Z(n33577) );
  XNOR U33935 ( .A(n33578), .B(n33573), .Z(n33574) );
  AND U33936 ( .A(b[2]), .B(a[25]), .Z(n33578) );
  NANDN U33937 ( .A(n31812), .B(n31810), .Z(n33567) );
  XNOR U33938 ( .A(n33579), .B(n33580), .Z(n31810) );
  NAND U33939 ( .A(a[26]), .B(b[0]), .Z(n31812) );
  XOR U33940 ( .A(n33573), .B(n33565), .Z(n33581) );
  XNOR U33941 ( .A(n33564), .B(n33560), .Z(n33582) );
  XNOR U33942 ( .A(n33559), .B(n33555), .Z(n33583) );
  XNOR U33943 ( .A(n33554), .B(n33550), .Z(n33584) );
  XNOR U33944 ( .A(n33549), .B(n33545), .Z(n33585) );
  XNOR U33945 ( .A(n33544), .B(n33540), .Z(n33586) );
  XNOR U33946 ( .A(n33539), .B(n33535), .Z(n33587) );
  XNOR U33947 ( .A(n33534), .B(n33530), .Z(n33588) );
  XNOR U33948 ( .A(n33529), .B(n33525), .Z(n33589) );
  XNOR U33949 ( .A(n33524), .B(n33520), .Z(n33590) );
  XNOR U33950 ( .A(n33519), .B(n33515), .Z(n33591) );
  XNOR U33951 ( .A(n33514), .B(n33510), .Z(n33592) );
  XNOR U33952 ( .A(n33509), .B(n33505), .Z(n33593) );
  XNOR U33953 ( .A(n33504), .B(n33500), .Z(n33594) );
  XNOR U33954 ( .A(n33499), .B(n33495), .Z(n33595) );
  XNOR U33955 ( .A(n33494), .B(n33490), .Z(n33596) );
  XNOR U33956 ( .A(n33489), .B(n33485), .Z(n33597) );
  XNOR U33957 ( .A(n33484), .B(n33480), .Z(n33598) );
  XNOR U33958 ( .A(n33479), .B(n33475), .Z(n33599) );
  XNOR U33959 ( .A(n33474), .B(n33470), .Z(n33600) );
  XNOR U33960 ( .A(n33469), .B(n33465), .Z(n33601) );
  XNOR U33961 ( .A(n33464), .B(n33460), .Z(n33602) );
  XNOR U33962 ( .A(n33459), .B(n33455), .Z(n33603) );
  XNOR U33963 ( .A(n33454), .B(n33450), .Z(n33604) );
  XOR U33964 ( .A(n33605), .B(n33449), .Z(n33450) );
  AND U33965 ( .A(a[0]), .B(b[27]), .Z(n33605) );
  XOR U33966 ( .A(n33606), .B(n33449), .Z(n33451) );
  XNOR U33967 ( .A(n33607), .B(n33608), .Z(n33449) );
  AND U33968 ( .A(n33609), .B(n33610), .Z(n33607) );
  AND U33969 ( .A(a[1]), .B(b[26]), .Z(n33606) );
  XOR U33970 ( .A(n33611), .B(n33454), .Z(n33456) );
  XOR U33971 ( .A(n33612), .B(n33613), .Z(n33454) );
  AND U33972 ( .A(n33614), .B(n33615), .Z(n33612) );
  AND U33973 ( .A(a[2]), .B(b[25]), .Z(n33611) );
  XOR U33974 ( .A(n33616), .B(n33459), .Z(n33461) );
  XOR U33975 ( .A(n33617), .B(n33618), .Z(n33459) );
  AND U33976 ( .A(n33619), .B(n33620), .Z(n33617) );
  AND U33977 ( .A(a[3]), .B(b[24]), .Z(n33616) );
  XOR U33978 ( .A(n33621), .B(n33464), .Z(n33466) );
  XOR U33979 ( .A(n33622), .B(n33623), .Z(n33464) );
  AND U33980 ( .A(n33624), .B(n33625), .Z(n33622) );
  AND U33981 ( .A(a[4]), .B(b[23]), .Z(n33621) );
  XOR U33982 ( .A(n33626), .B(n33469), .Z(n33471) );
  XOR U33983 ( .A(n33627), .B(n33628), .Z(n33469) );
  AND U33984 ( .A(n33629), .B(n33630), .Z(n33627) );
  AND U33985 ( .A(a[5]), .B(b[22]), .Z(n33626) );
  XOR U33986 ( .A(n33631), .B(n33474), .Z(n33476) );
  XOR U33987 ( .A(n33632), .B(n33633), .Z(n33474) );
  AND U33988 ( .A(n33634), .B(n33635), .Z(n33632) );
  AND U33989 ( .A(a[6]), .B(b[21]), .Z(n33631) );
  XOR U33990 ( .A(n33636), .B(n33479), .Z(n33481) );
  XOR U33991 ( .A(n33637), .B(n33638), .Z(n33479) );
  AND U33992 ( .A(n33639), .B(n33640), .Z(n33637) );
  AND U33993 ( .A(a[7]), .B(b[20]), .Z(n33636) );
  XOR U33994 ( .A(n33641), .B(n33484), .Z(n33486) );
  XOR U33995 ( .A(n33642), .B(n33643), .Z(n33484) );
  AND U33996 ( .A(n33644), .B(n33645), .Z(n33642) );
  AND U33997 ( .A(a[8]), .B(b[19]), .Z(n33641) );
  XOR U33998 ( .A(n33646), .B(n33489), .Z(n33491) );
  XOR U33999 ( .A(n33647), .B(n33648), .Z(n33489) );
  AND U34000 ( .A(n33649), .B(n33650), .Z(n33647) );
  AND U34001 ( .A(a[9]), .B(b[18]), .Z(n33646) );
  XOR U34002 ( .A(n33651), .B(n33494), .Z(n33496) );
  XOR U34003 ( .A(n33652), .B(n33653), .Z(n33494) );
  AND U34004 ( .A(n33654), .B(n33655), .Z(n33652) );
  AND U34005 ( .A(a[10]), .B(b[17]), .Z(n33651) );
  XOR U34006 ( .A(n33656), .B(n33499), .Z(n33501) );
  XOR U34007 ( .A(n33657), .B(n33658), .Z(n33499) );
  AND U34008 ( .A(n33659), .B(n33660), .Z(n33657) );
  AND U34009 ( .A(a[11]), .B(b[16]), .Z(n33656) );
  XOR U34010 ( .A(n33661), .B(n33504), .Z(n33506) );
  XOR U34011 ( .A(n33662), .B(n33663), .Z(n33504) );
  AND U34012 ( .A(n33664), .B(n33665), .Z(n33662) );
  AND U34013 ( .A(a[12]), .B(b[15]), .Z(n33661) );
  XOR U34014 ( .A(n33666), .B(n33509), .Z(n33511) );
  XOR U34015 ( .A(n33667), .B(n33668), .Z(n33509) );
  AND U34016 ( .A(n33669), .B(n33670), .Z(n33667) );
  AND U34017 ( .A(a[13]), .B(b[14]), .Z(n33666) );
  XOR U34018 ( .A(n33671), .B(n33514), .Z(n33516) );
  XOR U34019 ( .A(n33672), .B(n33673), .Z(n33514) );
  AND U34020 ( .A(n33674), .B(n33675), .Z(n33672) );
  AND U34021 ( .A(b[13]), .B(a[14]), .Z(n33671) );
  XOR U34022 ( .A(n33676), .B(n33519), .Z(n33521) );
  XOR U34023 ( .A(n33677), .B(n33678), .Z(n33519) );
  AND U34024 ( .A(n33679), .B(n33680), .Z(n33677) );
  AND U34025 ( .A(b[12]), .B(a[15]), .Z(n33676) );
  XOR U34026 ( .A(n33681), .B(n33524), .Z(n33526) );
  XOR U34027 ( .A(n33682), .B(n33683), .Z(n33524) );
  AND U34028 ( .A(n33684), .B(n33685), .Z(n33682) );
  AND U34029 ( .A(b[11]), .B(a[16]), .Z(n33681) );
  XOR U34030 ( .A(n33686), .B(n33529), .Z(n33531) );
  XOR U34031 ( .A(n33687), .B(n33688), .Z(n33529) );
  AND U34032 ( .A(n33689), .B(n33690), .Z(n33687) );
  AND U34033 ( .A(b[10]), .B(a[17]), .Z(n33686) );
  XOR U34034 ( .A(n33691), .B(n33534), .Z(n33536) );
  XOR U34035 ( .A(n33692), .B(n33693), .Z(n33534) );
  AND U34036 ( .A(n33694), .B(n33695), .Z(n33692) );
  AND U34037 ( .A(b[9]), .B(a[18]), .Z(n33691) );
  XOR U34038 ( .A(n33696), .B(n33539), .Z(n33541) );
  XOR U34039 ( .A(n33697), .B(n33698), .Z(n33539) );
  AND U34040 ( .A(n33699), .B(n33700), .Z(n33697) );
  AND U34041 ( .A(b[8]), .B(a[19]), .Z(n33696) );
  XOR U34042 ( .A(n33701), .B(n33544), .Z(n33546) );
  XOR U34043 ( .A(n33702), .B(n33703), .Z(n33544) );
  AND U34044 ( .A(n33704), .B(n33705), .Z(n33702) );
  AND U34045 ( .A(b[7]), .B(a[20]), .Z(n33701) );
  XOR U34046 ( .A(n33706), .B(n33549), .Z(n33551) );
  XOR U34047 ( .A(n33707), .B(n33708), .Z(n33549) );
  AND U34048 ( .A(n33709), .B(n33710), .Z(n33707) );
  AND U34049 ( .A(b[6]), .B(a[21]), .Z(n33706) );
  XOR U34050 ( .A(n33711), .B(n33554), .Z(n33556) );
  XOR U34051 ( .A(n33712), .B(n33713), .Z(n33554) );
  AND U34052 ( .A(n33714), .B(n33715), .Z(n33712) );
  AND U34053 ( .A(b[5]), .B(a[22]), .Z(n33711) );
  XOR U34054 ( .A(n33716), .B(n33559), .Z(n33561) );
  XOR U34055 ( .A(n33717), .B(n33718), .Z(n33559) );
  AND U34056 ( .A(n33719), .B(n33720), .Z(n33717) );
  AND U34057 ( .A(b[4]), .B(a[23]), .Z(n33716) );
  XNOR U34058 ( .A(n33721), .B(n33722), .Z(n33573) );
  NANDN U34059 ( .A(n33579), .B(n33580), .Z(n33722) );
  XOR U34060 ( .A(n33721), .B(n33723), .Z(n33580) );
  NAND U34061 ( .A(b[1]), .B(a[25]), .Z(n33723) );
  XOR U34062 ( .A(n33724), .B(n33725), .Z(n33579) );
  XOR U34063 ( .A(n33721), .B(n33726), .Z(n33725) );
  NANDN U34064 ( .A(n31817), .B(n31815), .Z(n33721) );
  XNOR U34065 ( .A(n33727), .B(n33728), .Z(n31815) );
  NAND U34066 ( .A(a[25]), .B(b[0]), .Z(n31817) );
  XOR U34067 ( .A(n33729), .B(n33564), .Z(n33566) );
  XNOR U34068 ( .A(n33730), .B(n33731), .Z(n33564) );
  AND U34069 ( .A(n33726), .B(n33724), .Z(n33730) );
  XOR U34070 ( .A(n33731), .B(n33719), .Z(n33732) );
  XNOR U34071 ( .A(n33718), .B(n33714), .Z(n33733) );
  XNOR U34072 ( .A(n33713), .B(n33709), .Z(n33734) );
  XNOR U34073 ( .A(n33708), .B(n33704), .Z(n33735) );
  XNOR U34074 ( .A(n33703), .B(n33699), .Z(n33736) );
  XNOR U34075 ( .A(n33698), .B(n33694), .Z(n33737) );
  XNOR U34076 ( .A(n33693), .B(n33689), .Z(n33738) );
  XNOR U34077 ( .A(n33688), .B(n33684), .Z(n33739) );
  XNOR U34078 ( .A(n33683), .B(n33679), .Z(n33740) );
  XNOR U34079 ( .A(n33678), .B(n33674), .Z(n33741) );
  XNOR U34080 ( .A(n33673), .B(n33669), .Z(n33742) );
  XNOR U34081 ( .A(n33668), .B(n33664), .Z(n33743) );
  XNOR U34082 ( .A(n33663), .B(n33659), .Z(n33744) );
  XNOR U34083 ( .A(n33658), .B(n33654), .Z(n33745) );
  XNOR U34084 ( .A(n33653), .B(n33649), .Z(n33746) );
  XNOR U34085 ( .A(n33648), .B(n33644), .Z(n33747) );
  XNOR U34086 ( .A(n33643), .B(n33639), .Z(n33748) );
  XNOR U34087 ( .A(n33638), .B(n33634), .Z(n33749) );
  XNOR U34088 ( .A(n33633), .B(n33629), .Z(n33750) );
  XNOR U34089 ( .A(n33628), .B(n33624), .Z(n33751) );
  XNOR U34090 ( .A(n33623), .B(n33619), .Z(n33752) );
  XNOR U34091 ( .A(n33618), .B(n33614), .Z(n33753) );
  XNOR U34092 ( .A(n33613), .B(n33609), .Z(n33754) );
  XNOR U34093 ( .A(n33755), .B(n33608), .Z(n33609) );
  AND U34094 ( .A(a[0]), .B(b[26]), .Z(n33755) );
  XNOR U34095 ( .A(n33756), .B(n33608), .Z(n33610) );
  XNOR U34096 ( .A(n33757), .B(n33758), .Z(n33608) );
  AND U34097 ( .A(n33759), .B(n33760), .Z(n33757) );
  AND U34098 ( .A(a[1]), .B(b[25]), .Z(n33756) );
  XOR U34099 ( .A(n33761), .B(n33613), .Z(n33615) );
  XOR U34100 ( .A(n33762), .B(n33763), .Z(n33613) );
  AND U34101 ( .A(n33764), .B(n33765), .Z(n33762) );
  AND U34102 ( .A(a[2]), .B(b[24]), .Z(n33761) );
  XOR U34103 ( .A(n33766), .B(n33618), .Z(n33620) );
  XOR U34104 ( .A(n33767), .B(n33768), .Z(n33618) );
  AND U34105 ( .A(n33769), .B(n33770), .Z(n33767) );
  AND U34106 ( .A(a[3]), .B(b[23]), .Z(n33766) );
  XOR U34107 ( .A(n33771), .B(n33623), .Z(n33625) );
  XOR U34108 ( .A(n33772), .B(n33773), .Z(n33623) );
  AND U34109 ( .A(n33774), .B(n33775), .Z(n33772) );
  AND U34110 ( .A(a[4]), .B(b[22]), .Z(n33771) );
  XOR U34111 ( .A(n33776), .B(n33628), .Z(n33630) );
  XOR U34112 ( .A(n33777), .B(n33778), .Z(n33628) );
  AND U34113 ( .A(n33779), .B(n33780), .Z(n33777) );
  AND U34114 ( .A(a[5]), .B(b[21]), .Z(n33776) );
  XOR U34115 ( .A(n33781), .B(n33633), .Z(n33635) );
  XOR U34116 ( .A(n33782), .B(n33783), .Z(n33633) );
  AND U34117 ( .A(n33784), .B(n33785), .Z(n33782) );
  AND U34118 ( .A(a[6]), .B(b[20]), .Z(n33781) );
  XOR U34119 ( .A(n33786), .B(n33638), .Z(n33640) );
  XOR U34120 ( .A(n33787), .B(n33788), .Z(n33638) );
  AND U34121 ( .A(n33789), .B(n33790), .Z(n33787) );
  AND U34122 ( .A(a[7]), .B(b[19]), .Z(n33786) );
  XOR U34123 ( .A(n33791), .B(n33643), .Z(n33645) );
  XOR U34124 ( .A(n33792), .B(n33793), .Z(n33643) );
  AND U34125 ( .A(n33794), .B(n33795), .Z(n33792) );
  AND U34126 ( .A(a[8]), .B(b[18]), .Z(n33791) );
  XOR U34127 ( .A(n33796), .B(n33648), .Z(n33650) );
  XOR U34128 ( .A(n33797), .B(n33798), .Z(n33648) );
  AND U34129 ( .A(n33799), .B(n33800), .Z(n33797) );
  AND U34130 ( .A(a[9]), .B(b[17]), .Z(n33796) );
  XOR U34131 ( .A(n33801), .B(n33653), .Z(n33655) );
  XOR U34132 ( .A(n33802), .B(n33803), .Z(n33653) );
  AND U34133 ( .A(n33804), .B(n33805), .Z(n33802) );
  AND U34134 ( .A(a[10]), .B(b[16]), .Z(n33801) );
  XOR U34135 ( .A(n33806), .B(n33658), .Z(n33660) );
  XOR U34136 ( .A(n33807), .B(n33808), .Z(n33658) );
  AND U34137 ( .A(n33809), .B(n33810), .Z(n33807) );
  AND U34138 ( .A(a[11]), .B(b[15]), .Z(n33806) );
  XOR U34139 ( .A(n33811), .B(n33663), .Z(n33665) );
  XOR U34140 ( .A(n33812), .B(n33813), .Z(n33663) );
  AND U34141 ( .A(n33814), .B(n33815), .Z(n33812) );
  AND U34142 ( .A(a[12]), .B(b[14]), .Z(n33811) );
  XOR U34143 ( .A(n33816), .B(n33668), .Z(n33670) );
  XOR U34144 ( .A(n33817), .B(n33818), .Z(n33668) );
  AND U34145 ( .A(n33819), .B(n33820), .Z(n33817) );
  AND U34146 ( .A(a[13]), .B(b[13]), .Z(n33816) );
  XOR U34147 ( .A(n33821), .B(n33673), .Z(n33675) );
  XOR U34148 ( .A(n33822), .B(n33823), .Z(n33673) );
  AND U34149 ( .A(n33824), .B(n33825), .Z(n33822) );
  AND U34150 ( .A(b[12]), .B(a[14]), .Z(n33821) );
  XOR U34151 ( .A(n33826), .B(n33678), .Z(n33680) );
  XOR U34152 ( .A(n33827), .B(n33828), .Z(n33678) );
  AND U34153 ( .A(n33829), .B(n33830), .Z(n33827) );
  AND U34154 ( .A(b[11]), .B(a[15]), .Z(n33826) );
  XOR U34155 ( .A(n33831), .B(n33683), .Z(n33685) );
  XOR U34156 ( .A(n33832), .B(n33833), .Z(n33683) );
  AND U34157 ( .A(n33834), .B(n33835), .Z(n33832) );
  AND U34158 ( .A(b[10]), .B(a[16]), .Z(n33831) );
  XOR U34159 ( .A(n33836), .B(n33688), .Z(n33690) );
  XOR U34160 ( .A(n33837), .B(n33838), .Z(n33688) );
  AND U34161 ( .A(n33839), .B(n33840), .Z(n33837) );
  AND U34162 ( .A(b[9]), .B(a[17]), .Z(n33836) );
  XOR U34163 ( .A(n33841), .B(n33693), .Z(n33695) );
  XOR U34164 ( .A(n33842), .B(n33843), .Z(n33693) );
  AND U34165 ( .A(n33844), .B(n33845), .Z(n33842) );
  AND U34166 ( .A(b[8]), .B(a[18]), .Z(n33841) );
  XOR U34167 ( .A(n33846), .B(n33698), .Z(n33700) );
  XOR U34168 ( .A(n33847), .B(n33848), .Z(n33698) );
  AND U34169 ( .A(n33849), .B(n33850), .Z(n33847) );
  AND U34170 ( .A(b[7]), .B(a[19]), .Z(n33846) );
  XOR U34171 ( .A(n33851), .B(n33703), .Z(n33705) );
  XOR U34172 ( .A(n33852), .B(n33853), .Z(n33703) );
  AND U34173 ( .A(n33854), .B(n33855), .Z(n33852) );
  AND U34174 ( .A(b[6]), .B(a[20]), .Z(n33851) );
  XOR U34175 ( .A(n33856), .B(n33708), .Z(n33710) );
  XOR U34176 ( .A(n33857), .B(n33858), .Z(n33708) );
  AND U34177 ( .A(n33859), .B(n33860), .Z(n33857) );
  AND U34178 ( .A(b[5]), .B(a[21]), .Z(n33856) );
  XOR U34179 ( .A(n33861), .B(n33713), .Z(n33715) );
  XOR U34180 ( .A(n33862), .B(n33863), .Z(n33713) );
  AND U34181 ( .A(n33864), .B(n33865), .Z(n33862) );
  AND U34182 ( .A(b[4]), .B(a[22]), .Z(n33861) );
  XOR U34183 ( .A(n33866), .B(n33718), .Z(n33720) );
  XNOR U34184 ( .A(n33867), .B(n33868), .Z(n33718) );
  AND U34185 ( .A(n33869), .B(n33870), .Z(n33867) );
  AND U34186 ( .A(b[3]), .B(a[23]), .Z(n33866) );
  XNOR U34187 ( .A(n33871), .B(n33731), .Z(n33726) );
  XNOR U34188 ( .A(n33872), .B(n33873), .Z(n33731) );
  NANDN U34189 ( .A(n33727), .B(n33728), .Z(n33873) );
  XOR U34190 ( .A(n33872), .B(n33874), .Z(n33728) );
  NAND U34191 ( .A(b[1]), .B(a[24]), .Z(n33874) );
  XOR U34192 ( .A(n33870), .B(n33875), .Z(n33727) );
  XOR U34193 ( .A(n33872), .B(n33869), .Z(n33875) );
  XNOR U34194 ( .A(n33876), .B(n33868), .Z(n33869) );
  AND U34195 ( .A(b[2]), .B(a[23]), .Z(n33876) );
  XOR U34196 ( .A(n33868), .B(n33864), .Z(n33877) );
  XNOR U34197 ( .A(n33863), .B(n33859), .Z(n33878) );
  XNOR U34198 ( .A(n33858), .B(n33854), .Z(n33879) );
  XNOR U34199 ( .A(n33853), .B(n33849), .Z(n33880) );
  XNOR U34200 ( .A(n33848), .B(n33844), .Z(n33881) );
  XNOR U34201 ( .A(n33843), .B(n33839), .Z(n33882) );
  XNOR U34202 ( .A(n33838), .B(n33834), .Z(n33883) );
  XNOR U34203 ( .A(n33833), .B(n33829), .Z(n33884) );
  XNOR U34204 ( .A(n33828), .B(n33824), .Z(n33885) );
  XNOR U34205 ( .A(n33823), .B(n33819), .Z(n33886) );
  XNOR U34206 ( .A(n33818), .B(n33814), .Z(n33887) );
  XNOR U34207 ( .A(n33813), .B(n33809), .Z(n33888) );
  XNOR U34208 ( .A(n33808), .B(n33804), .Z(n33889) );
  XNOR U34209 ( .A(n33803), .B(n33799), .Z(n33890) );
  XNOR U34210 ( .A(n33798), .B(n33794), .Z(n33891) );
  XNOR U34211 ( .A(n33793), .B(n33789), .Z(n33892) );
  XNOR U34212 ( .A(n33788), .B(n33784), .Z(n33893) );
  XNOR U34213 ( .A(n33783), .B(n33779), .Z(n33894) );
  XNOR U34214 ( .A(n33778), .B(n33774), .Z(n33895) );
  XNOR U34215 ( .A(n33773), .B(n33769), .Z(n33896) );
  XNOR U34216 ( .A(n33768), .B(n33764), .Z(n33897) );
  XNOR U34217 ( .A(n33763), .B(n33759), .Z(n33898) );
  XOR U34218 ( .A(n33899), .B(n33758), .Z(n33759) );
  AND U34219 ( .A(a[0]), .B(b[25]), .Z(n33899) );
  XOR U34220 ( .A(n33900), .B(n33758), .Z(n33760) );
  XNOR U34221 ( .A(n33901), .B(n33902), .Z(n33758) );
  AND U34222 ( .A(n33903), .B(n33904), .Z(n33901) );
  AND U34223 ( .A(a[1]), .B(b[24]), .Z(n33900) );
  XOR U34224 ( .A(n33905), .B(n33763), .Z(n33765) );
  XOR U34225 ( .A(n33906), .B(n33907), .Z(n33763) );
  AND U34226 ( .A(n33908), .B(n33909), .Z(n33906) );
  AND U34227 ( .A(a[2]), .B(b[23]), .Z(n33905) );
  XOR U34228 ( .A(n33910), .B(n33768), .Z(n33770) );
  XOR U34229 ( .A(n33911), .B(n33912), .Z(n33768) );
  AND U34230 ( .A(n33913), .B(n33914), .Z(n33911) );
  AND U34231 ( .A(a[3]), .B(b[22]), .Z(n33910) );
  XOR U34232 ( .A(n33915), .B(n33773), .Z(n33775) );
  XOR U34233 ( .A(n33916), .B(n33917), .Z(n33773) );
  AND U34234 ( .A(n33918), .B(n33919), .Z(n33916) );
  AND U34235 ( .A(a[4]), .B(b[21]), .Z(n33915) );
  XOR U34236 ( .A(n33920), .B(n33778), .Z(n33780) );
  XOR U34237 ( .A(n33921), .B(n33922), .Z(n33778) );
  AND U34238 ( .A(n33923), .B(n33924), .Z(n33921) );
  AND U34239 ( .A(a[5]), .B(b[20]), .Z(n33920) );
  XOR U34240 ( .A(n33925), .B(n33783), .Z(n33785) );
  XOR U34241 ( .A(n33926), .B(n33927), .Z(n33783) );
  AND U34242 ( .A(n33928), .B(n33929), .Z(n33926) );
  AND U34243 ( .A(a[6]), .B(b[19]), .Z(n33925) );
  XOR U34244 ( .A(n33930), .B(n33788), .Z(n33790) );
  XOR U34245 ( .A(n33931), .B(n33932), .Z(n33788) );
  AND U34246 ( .A(n33933), .B(n33934), .Z(n33931) );
  AND U34247 ( .A(a[7]), .B(b[18]), .Z(n33930) );
  XOR U34248 ( .A(n33935), .B(n33793), .Z(n33795) );
  XOR U34249 ( .A(n33936), .B(n33937), .Z(n33793) );
  AND U34250 ( .A(n33938), .B(n33939), .Z(n33936) );
  AND U34251 ( .A(a[8]), .B(b[17]), .Z(n33935) );
  XOR U34252 ( .A(n33940), .B(n33798), .Z(n33800) );
  XOR U34253 ( .A(n33941), .B(n33942), .Z(n33798) );
  AND U34254 ( .A(n33943), .B(n33944), .Z(n33941) );
  AND U34255 ( .A(a[9]), .B(b[16]), .Z(n33940) );
  XOR U34256 ( .A(n33945), .B(n33803), .Z(n33805) );
  XOR U34257 ( .A(n33946), .B(n33947), .Z(n33803) );
  AND U34258 ( .A(n33948), .B(n33949), .Z(n33946) );
  AND U34259 ( .A(a[10]), .B(b[15]), .Z(n33945) );
  XOR U34260 ( .A(n33950), .B(n33808), .Z(n33810) );
  XOR U34261 ( .A(n33951), .B(n33952), .Z(n33808) );
  AND U34262 ( .A(n33953), .B(n33954), .Z(n33951) );
  AND U34263 ( .A(a[11]), .B(b[14]), .Z(n33950) );
  XOR U34264 ( .A(n33955), .B(n33813), .Z(n33815) );
  XOR U34265 ( .A(n33956), .B(n33957), .Z(n33813) );
  AND U34266 ( .A(n33958), .B(n33959), .Z(n33956) );
  AND U34267 ( .A(a[12]), .B(b[13]), .Z(n33955) );
  XOR U34268 ( .A(n33960), .B(n33818), .Z(n33820) );
  XOR U34269 ( .A(n33961), .B(n33962), .Z(n33818) );
  AND U34270 ( .A(n33963), .B(n33964), .Z(n33961) );
  AND U34271 ( .A(b[12]), .B(a[13]), .Z(n33960) );
  XOR U34272 ( .A(n33965), .B(n33823), .Z(n33825) );
  XOR U34273 ( .A(n33966), .B(n33967), .Z(n33823) );
  AND U34274 ( .A(n33968), .B(n33969), .Z(n33966) );
  AND U34275 ( .A(b[11]), .B(a[14]), .Z(n33965) );
  XOR U34276 ( .A(n33970), .B(n33828), .Z(n33830) );
  XOR U34277 ( .A(n33971), .B(n33972), .Z(n33828) );
  AND U34278 ( .A(n33973), .B(n33974), .Z(n33971) );
  AND U34279 ( .A(b[10]), .B(a[15]), .Z(n33970) );
  XOR U34280 ( .A(n33975), .B(n33833), .Z(n33835) );
  XOR U34281 ( .A(n33976), .B(n33977), .Z(n33833) );
  AND U34282 ( .A(n33978), .B(n33979), .Z(n33976) );
  AND U34283 ( .A(b[9]), .B(a[16]), .Z(n33975) );
  XOR U34284 ( .A(n33980), .B(n33838), .Z(n33840) );
  XOR U34285 ( .A(n33981), .B(n33982), .Z(n33838) );
  AND U34286 ( .A(n33983), .B(n33984), .Z(n33981) );
  AND U34287 ( .A(b[8]), .B(a[17]), .Z(n33980) );
  XOR U34288 ( .A(n33985), .B(n33843), .Z(n33845) );
  XOR U34289 ( .A(n33986), .B(n33987), .Z(n33843) );
  AND U34290 ( .A(n33988), .B(n33989), .Z(n33986) );
  AND U34291 ( .A(b[7]), .B(a[18]), .Z(n33985) );
  XOR U34292 ( .A(n33990), .B(n33848), .Z(n33850) );
  XOR U34293 ( .A(n33991), .B(n33992), .Z(n33848) );
  AND U34294 ( .A(n33993), .B(n33994), .Z(n33991) );
  AND U34295 ( .A(b[6]), .B(a[19]), .Z(n33990) );
  XOR U34296 ( .A(n33995), .B(n33853), .Z(n33855) );
  XOR U34297 ( .A(n33996), .B(n33997), .Z(n33853) );
  AND U34298 ( .A(n33998), .B(n33999), .Z(n33996) );
  AND U34299 ( .A(b[5]), .B(a[20]), .Z(n33995) );
  XOR U34300 ( .A(n34000), .B(n33858), .Z(n33860) );
  XOR U34301 ( .A(n34001), .B(n34002), .Z(n33858) );
  AND U34302 ( .A(n34003), .B(n34004), .Z(n34001) );
  AND U34303 ( .A(b[4]), .B(a[21]), .Z(n34000) );
  XNOR U34304 ( .A(n34005), .B(n34006), .Z(n33868) );
  NANDN U34305 ( .A(n34007), .B(n34008), .Z(n34006) );
  XOR U34306 ( .A(n34009), .B(n33863), .Z(n33865) );
  XNOR U34307 ( .A(n34010), .B(n34011), .Z(n33863) );
  AND U34308 ( .A(n34012), .B(n34013), .Z(n34010) );
  AND U34309 ( .A(b[3]), .B(a[22]), .Z(n34009) );
  NANDN U34310 ( .A(n31822), .B(n31820), .Z(n33872) );
  XNOR U34311 ( .A(n34007), .B(n34008), .Z(n31820) );
  XOR U34312 ( .A(n34005), .B(n34014), .Z(n34008) );
  NAND U34313 ( .A(b[1]), .B(a[23]), .Z(n34014) );
  XOR U34314 ( .A(n34013), .B(n34015), .Z(n34007) );
  XOR U34315 ( .A(n34005), .B(n34012), .Z(n34015) );
  XNOR U34316 ( .A(n34016), .B(n34011), .Z(n34012) );
  AND U34317 ( .A(b[2]), .B(a[22]), .Z(n34016) );
  NANDN U34318 ( .A(n31827), .B(n31825), .Z(n34005) );
  XNOR U34319 ( .A(n34017), .B(n34018), .Z(n31825) );
  NAND U34320 ( .A(a[23]), .B(b[0]), .Z(n31827) );
  XOR U34321 ( .A(n34011), .B(n34003), .Z(n34019) );
  XNOR U34322 ( .A(n34002), .B(n33998), .Z(n34020) );
  XNOR U34323 ( .A(n33997), .B(n33993), .Z(n34021) );
  XNOR U34324 ( .A(n33992), .B(n33988), .Z(n34022) );
  XNOR U34325 ( .A(n33987), .B(n33983), .Z(n34023) );
  XNOR U34326 ( .A(n33982), .B(n33978), .Z(n34024) );
  XNOR U34327 ( .A(n33977), .B(n33973), .Z(n34025) );
  XNOR U34328 ( .A(n33972), .B(n33968), .Z(n34026) );
  XNOR U34329 ( .A(n33967), .B(n33963), .Z(n34027) );
  XNOR U34330 ( .A(n33962), .B(n33958), .Z(n34028) );
  XNOR U34331 ( .A(n33957), .B(n33953), .Z(n34029) );
  XNOR U34332 ( .A(n33952), .B(n33948), .Z(n34030) );
  XNOR U34333 ( .A(n33947), .B(n33943), .Z(n34031) );
  XNOR U34334 ( .A(n33942), .B(n33938), .Z(n34032) );
  XNOR U34335 ( .A(n33937), .B(n33933), .Z(n34033) );
  XNOR U34336 ( .A(n33932), .B(n33928), .Z(n34034) );
  XNOR U34337 ( .A(n33927), .B(n33923), .Z(n34035) );
  XNOR U34338 ( .A(n33922), .B(n33918), .Z(n34036) );
  XNOR U34339 ( .A(n33917), .B(n33913), .Z(n34037) );
  XNOR U34340 ( .A(n33912), .B(n33908), .Z(n34038) );
  XNOR U34341 ( .A(n33907), .B(n33903), .Z(n34039) );
  XNOR U34342 ( .A(n34040), .B(n33902), .Z(n33903) );
  AND U34343 ( .A(a[0]), .B(b[24]), .Z(n34040) );
  XNOR U34344 ( .A(n34041), .B(n33902), .Z(n33904) );
  XNOR U34345 ( .A(n34042), .B(n34043), .Z(n33902) );
  AND U34346 ( .A(n34044), .B(n34045), .Z(n34042) );
  AND U34347 ( .A(a[1]), .B(b[23]), .Z(n34041) );
  XOR U34348 ( .A(n34046), .B(n33907), .Z(n33909) );
  XOR U34349 ( .A(n34047), .B(n34048), .Z(n33907) );
  AND U34350 ( .A(n34049), .B(n34050), .Z(n34047) );
  AND U34351 ( .A(a[2]), .B(b[22]), .Z(n34046) );
  XOR U34352 ( .A(n34051), .B(n33912), .Z(n33914) );
  XOR U34353 ( .A(n34052), .B(n34053), .Z(n33912) );
  AND U34354 ( .A(n34054), .B(n34055), .Z(n34052) );
  AND U34355 ( .A(a[3]), .B(b[21]), .Z(n34051) );
  XOR U34356 ( .A(n34056), .B(n33917), .Z(n33919) );
  XOR U34357 ( .A(n34057), .B(n34058), .Z(n33917) );
  AND U34358 ( .A(n34059), .B(n34060), .Z(n34057) );
  AND U34359 ( .A(a[4]), .B(b[20]), .Z(n34056) );
  XOR U34360 ( .A(n34061), .B(n33922), .Z(n33924) );
  XOR U34361 ( .A(n34062), .B(n34063), .Z(n33922) );
  AND U34362 ( .A(n34064), .B(n34065), .Z(n34062) );
  AND U34363 ( .A(a[5]), .B(b[19]), .Z(n34061) );
  XOR U34364 ( .A(n34066), .B(n33927), .Z(n33929) );
  XOR U34365 ( .A(n34067), .B(n34068), .Z(n33927) );
  AND U34366 ( .A(n34069), .B(n34070), .Z(n34067) );
  AND U34367 ( .A(a[6]), .B(b[18]), .Z(n34066) );
  XOR U34368 ( .A(n34071), .B(n33932), .Z(n33934) );
  XOR U34369 ( .A(n34072), .B(n34073), .Z(n33932) );
  AND U34370 ( .A(n34074), .B(n34075), .Z(n34072) );
  AND U34371 ( .A(a[7]), .B(b[17]), .Z(n34071) );
  XOR U34372 ( .A(n34076), .B(n33937), .Z(n33939) );
  XOR U34373 ( .A(n34077), .B(n34078), .Z(n33937) );
  AND U34374 ( .A(n34079), .B(n34080), .Z(n34077) );
  AND U34375 ( .A(a[8]), .B(b[16]), .Z(n34076) );
  XOR U34376 ( .A(n34081), .B(n33942), .Z(n33944) );
  XOR U34377 ( .A(n34082), .B(n34083), .Z(n33942) );
  AND U34378 ( .A(n34084), .B(n34085), .Z(n34082) );
  AND U34379 ( .A(a[9]), .B(b[15]), .Z(n34081) );
  XOR U34380 ( .A(n34086), .B(n33947), .Z(n33949) );
  XOR U34381 ( .A(n34087), .B(n34088), .Z(n33947) );
  AND U34382 ( .A(n34089), .B(n34090), .Z(n34087) );
  AND U34383 ( .A(a[10]), .B(b[14]), .Z(n34086) );
  XOR U34384 ( .A(n34091), .B(n33952), .Z(n33954) );
  XOR U34385 ( .A(n34092), .B(n34093), .Z(n33952) );
  AND U34386 ( .A(n34094), .B(n34095), .Z(n34092) );
  AND U34387 ( .A(a[11]), .B(b[13]), .Z(n34091) );
  XOR U34388 ( .A(n34096), .B(n33957), .Z(n33959) );
  XOR U34389 ( .A(n34097), .B(n34098), .Z(n33957) );
  AND U34390 ( .A(n34099), .B(n34100), .Z(n34097) );
  AND U34391 ( .A(a[12]), .B(b[12]), .Z(n34096) );
  XOR U34392 ( .A(n34101), .B(n33962), .Z(n33964) );
  XOR U34393 ( .A(n34102), .B(n34103), .Z(n33962) );
  AND U34394 ( .A(n34104), .B(n34105), .Z(n34102) );
  AND U34395 ( .A(b[11]), .B(a[13]), .Z(n34101) );
  XOR U34396 ( .A(n34106), .B(n33967), .Z(n33969) );
  XOR U34397 ( .A(n34107), .B(n34108), .Z(n33967) );
  AND U34398 ( .A(n34109), .B(n34110), .Z(n34107) );
  AND U34399 ( .A(b[10]), .B(a[14]), .Z(n34106) );
  XOR U34400 ( .A(n34111), .B(n33972), .Z(n33974) );
  XOR U34401 ( .A(n34112), .B(n34113), .Z(n33972) );
  AND U34402 ( .A(n34114), .B(n34115), .Z(n34112) );
  AND U34403 ( .A(b[9]), .B(a[15]), .Z(n34111) );
  XOR U34404 ( .A(n34116), .B(n33977), .Z(n33979) );
  XOR U34405 ( .A(n34117), .B(n34118), .Z(n33977) );
  AND U34406 ( .A(n34119), .B(n34120), .Z(n34117) );
  AND U34407 ( .A(b[8]), .B(a[16]), .Z(n34116) );
  XOR U34408 ( .A(n34121), .B(n33982), .Z(n33984) );
  XOR U34409 ( .A(n34122), .B(n34123), .Z(n33982) );
  AND U34410 ( .A(n34124), .B(n34125), .Z(n34122) );
  AND U34411 ( .A(b[7]), .B(a[17]), .Z(n34121) );
  XOR U34412 ( .A(n34126), .B(n33987), .Z(n33989) );
  XOR U34413 ( .A(n34127), .B(n34128), .Z(n33987) );
  AND U34414 ( .A(n34129), .B(n34130), .Z(n34127) );
  AND U34415 ( .A(b[6]), .B(a[18]), .Z(n34126) );
  XOR U34416 ( .A(n34131), .B(n33992), .Z(n33994) );
  XOR U34417 ( .A(n34132), .B(n34133), .Z(n33992) );
  AND U34418 ( .A(n34134), .B(n34135), .Z(n34132) );
  AND U34419 ( .A(b[5]), .B(a[19]), .Z(n34131) );
  XOR U34420 ( .A(n34136), .B(n33997), .Z(n33999) );
  XOR U34421 ( .A(n34137), .B(n34138), .Z(n33997) );
  AND U34422 ( .A(n34139), .B(n34140), .Z(n34137) );
  AND U34423 ( .A(b[4]), .B(a[20]), .Z(n34136) );
  XNOR U34424 ( .A(n34141), .B(n34142), .Z(n34011) );
  NANDN U34425 ( .A(n34017), .B(n34018), .Z(n34142) );
  XOR U34426 ( .A(n34141), .B(n34143), .Z(n34018) );
  NAND U34427 ( .A(b[1]), .B(a[22]), .Z(n34143) );
  XOR U34428 ( .A(n34144), .B(n34145), .Z(n34017) );
  XOR U34429 ( .A(n34141), .B(n34146), .Z(n34145) );
  NANDN U34430 ( .A(n31832), .B(n31830), .Z(n34141) );
  XNOR U34431 ( .A(n34147), .B(n34148), .Z(n31830) );
  NAND U34432 ( .A(a[22]), .B(b[0]), .Z(n31832) );
  XOR U34433 ( .A(n34149), .B(n34002), .Z(n34004) );
  XNOR U34434 ( .A(n34150), .B(n34151), .Z(n34002) );
  AND U34435 ( .A(n34146), .B(n34144), .Z(n34150) );
  XOR U34436 ( .A(n34151), .B(n34139), .Z(n34152) );
  XNOR U34437 ( .A(n34138), .B(n34134), .Z(n34153) );
  XNOR U34438 ( .A(n34133), .B(n34129), .Z(n34154) );
  XNOR U34439 ( .A(n34128), .B(n34124), .Z(n34155) );
  XNOR U34440 ( .A(n34123), .B(n34119), .Z(n34156) );
  XNOR U34441 ( .A(n34118), .B(n34114), .Z(n34157) );
  XNOR U34442 ( .A(n34113), .B(n34109), .Z(n34158) );
  XNOR U34443 ( .A(n34108), .B(n34104), .Z(n34159) );
  XNOR U34444 ( .A(n34103), .B(n34099), .Z(n34160) );
  XNOR U34445 ( .A(n34098), .B(n34094), .Z(n34161) );
  XNOR U34446 ( .A(n34093), .B(n34089), .Z(n34162) );
  XNOR U34447 ( .A(n34088), .B(n34084), .Z(n34163) );
  XNOR U34448 ( .A(n34083), .B(n34079), .Z(n34164) );
  XNOR U34449 ( .A(n34078), .B(n34074), .Z(n34165) );
  XNOR U34450 ( .A(n34073), .B(n34069), .Z(n34166) );
  XNOR U34451 ( .A(n34068), .B(n34064), .Z(n34167) );
  XNOR U34452 ( .A(n34063), .B(n34059), .Z(n34168) );
  XNOR U34453 ( .A(n34058), .B(n34054), .Z(n34169) );
  XNOR U34454 ( .A(n34053), .B(n34049), .Z(n34170) );
  XNOR U34455 ( .A(n34048), .B(n34044), .Z(n34171) );
  XOR U34456 ( .A(n34172), .B(n34043), .Z(n34044) );
  AND U34457 ( .A(a[0]), .B(b[23]), .Z(n34172) );
  XOR U34458 ( .A(n34173), .B(n34043), .Z(n34045) );
  XNOR U34459 ( .A(n34174), .B(n34175), .Z(n34043) );
  AND U34460 ( .A(n34176), .B(n34177), .Z(n34174) );
  AND U34461 ( .A(a[1]), .B(b[22]), .Z(n34173) );
  XOR U34462 ( .A(n34178), .B(n34048), .Z(n34050) );
  XOR U34463 ( .A(n34179), .B(n34180), .Z(n34048) );
  AND U34464 ( .A(n34181), .B(n34182), .Z(n34179) );
  AND U34465 ( .A(a[2]), .B(b[21]), .Z(n34178) );
  XOR U34466 ( .A(n34183), .B(n34053), .Z(n34055) );
  XOR U34467 ( .A(n34184), .B(n34185), .Z(n34053) );
  AND U34468 ( .A(n34186), .B(n34187), .Z(n34184) );
  AND U34469 ( .A(a[3]), .B(b[20]), .Z(n34183) );
  XOR U34470 ( .A(n34188), .B(n34058), .Z(n34060) );
  XOR U34471 ( .A(n34189), .B(n34190), .Z(n34058) );
  AND U34472 ( .A(n34191), .B(n34192), .Z(n34189) );
  AND U34473 ( .A(a[4]), .B(b[19]), .Z(n34188) );
  XOR U34474 ( .A(n34193), .B(n34063), .Z(n34065) );
  XOR U34475 ( .A(n34194), .B(n34195), .Z(n34063) );
  AND U34476 ( .A(n34196), .B(n34197), .Z(n34194) );
  AND U34477 ( .A(a[5]), .B(b[18]), .Z(n34193) );
  XOR U34478 ( .A(n34198), .B(n34068), .Z(n34070) );
  XOR U34479 ( .A(n34199), .B(n34200), .Z(n34068) );
  AND U34480 ( .A(n34201), .B(n34202), .Z(n34199) );
  AND U34481 ( .A(a[6]), .B(b[17]), .Z(n34198) );
  XOR U34482 ( .A(n34203), .B(n34073), .Z(n34075) );
  XOR U34483 ( .A(n34204), .B(n34205), .Z(n34073) );
  AND U34484 ( .A(n34206), .B(n34207), .Z(n34204) );
  AND U34485 ( .A(a[7]), .B(b[16]), .Z(n34203) );
  XOR U34486 ( .A(n34208), .B(n34078), .Z(n34080) );
  XOR U34487 ( .A(n34209), .B(n34210), .Z(n34078) );
  AND U34488 ( .A(n34211), .B(n34212), .Z(n34209) );
  AND U34489 ( .A(a[8]), .B(b[15]), .Z(n34208) );
  XOR U34490 ( .A(n34213), .B(n34083), .Z(n34085) );
  XOR U34491 ( .A(n34214), .B(n34215), .Z(n34083) );
  AND U34492 ( .A(n34216), .B(n34217), .Z(n34214) );
  AND U34493 ( .A(a[9]), .B(b[14]), .Z(n34213) );
  XOR U34494 ( .A(n34218), .B(n34088), .Z(n34090) );
  XOR U34495 ( .A(n34219), .B(n34220), .Z(n34088) );
  AND U34496 ( .A(n34221), .B(n34222), .Z(n34219) );
  AND U34497 ( .A(a[10]), .B(b[13]), .Z(n34218) );
  XOR U34498 ( .A(n34223), .B(n34093), .Z(n34095) );
  XOR U34499 ( .A(n34224), .B(n34225), .Z(n34093) );
  AND U34500 ( .A(n34226), .B(n34227), .Z(n34224) );
  AND U34501 ( .A(a[11]), .B(b[12]), .Z(n34223) );
  XOR U34502 ( .A(n34228), .B(n34098), .Z(n34100) );
  XOR U34503 ( .A(n34229), .B(n34230), .Z(n34098) );
  AND U34504 ( .A(n34231), .B(n34232), .Z(n34229) );
  AND U34505 ( .A(b[11]), .B(a[12]), .Z(n34228) );
  XOR U34506 ( .A(n34233), .B(n34103), .Z(n34105) );
  XOR U34507 ( .A(n34234), .B(n34235), .Z(n34103) );
  AND U34508 ( .A(n34236), .B(n34237), .Z(n34234) );
  AND U34509 ( .A(b[10]), .B(a[13]), .Z(n34233) );
  XOR U34510 ( .A(n34238), .B(n34108), .Z(n34110) );
  XOR U34511 ( .A(n34239), .B(n34240), .Z(n34108) );
  AND U34512 ( .A(n34241), .B(n34242), .Z(n34239) );
  AND U34513 ( .A(b[9]), .B(a[14]), .Z(n34238) );
  XOR U34514 ( .A(n34243), .B(n34113), .Z(n34115) );
  XOR U34515 ( .A(n34244), .B(n34245), .Z(n34113) );
  AND U34516 ( .A(n34246), .B(n34247), .Z(n34244) );
  AND U34517 ( .A(b[8]), .B(a[15]), .Z(n34243) );
  XOR U34518 ( .A(n34248), .B(n34118), .Z(n34120) );
  XOR U34519 ( .A(n34249), .B(n34250), .Z(n34118) );
  AND U34520 ( .A(n34251), .B(n34252), .Z(n34249) );
  AND U34521 ( .A(b[7]), .B(a[16]), .Z(n34248) );
  XOR U34522 ( .A(n34253), .B(n34123), .Z(n34125) );
  XOR U34523 ( .A(n34254), .B(n34255), .Z(n34123) );
  AND U34524 ( .A(n34256), .B(n34257), .Z(n34254) );
  AND U34525 ( .A(b[6]), .B(a[17]), .Z(n34253) );
  XOR U34526 ( .A(n34258), .B(n34128), .Z(n34130) );
  XOR U34527 ( .A(n34259), .B(n34260), .Z(n34128) );
  AND U34528 ( .A(n34261), .B(n34262), .Z(n34259) );
  AND U34529 ( .A(b[5]), .B(a[18]), .Z(n34258) );
  XOR U34530 ( .A(n34263), .B(n34133), .Z(n34135) );
  XOR U34531 ( .A(n34264), .B(n34265), .Z(n34133) );
  AND U34532 ( .A(n34266), .B(n34267), .Z(n34264) );
  AND U34533 ( .A(b[4]), .B(a[19]), .Z(n34263) );
  XOR U34534 ( .A(n34268), .B(n34138), .Z(n34140) );
  XNOR U34535 ( .A(n34269), .B(n34270), .Z(n34138) );
  AND U34536 ( .A(n34271), .B(n34272), .Z(n34269) );
  AND U34537 ( .A(b[3]), .B(a[20]), .Z(n34268) );
  XNOR U34538 ( .A(n34273), .B(n34151), .Z(n34146) );
  XNOR U34539 ( .A(n34274), .B(n34275), .Z(n34151) );
  NANDN U34540 ( .A(n34147), .B(n34148), .Z(n34275) );
  XOR U34541 ( .A(n34274), .B(n34276), .Z(n34148) );
  NAND U34542 ( .A(b[1]), .B(a[21]), .Z(n34276) );
  XOR U34543 ( .A(n34272), .B(n34277), .Z(n34147) );
  XOR U34544 ( .A(n34274), .B(n34271), .Z(n34277) );
  XNOR U34545 ( .A(n34278), .B(n34270), .Z(n34271) );
  AND U34546 ( .A(b[2]), .B(a[20]), .Z(n34278) );
  XOR U34547 ( .A(n34270), .B(n34266), .Z(n34279) );
  XNOR U34548 ( .A(n34265), .B(n34261), .Z(n34280) );
  XNOR U34549 ( .A(n34260), .B(n34256), .Z(n34281) );
  XNOR U34550 ( .A(n34255), .B(n34251), .Z(n34282) );
  XNOR U34551 ( .A(n34250), .B(n34246), .Z(n34283) );
  XNOR U34552 ( .A(n34245), .B(n34241), .Z(n34284) );
  XNOR U34553 ( .A(n34240), .B(n34236), .Z(n34285) );
  XNOR U34554 ( .A(n34235), .B(n34231), .Z(n34286) );
  XNOR U34555 ( .A(n34230), .B(n34226), .Z(n34287) );
  XNOR U34556 ( .A(n34225), .B(n34221), .Z(n34288) );
  XNOR U34557 ( .A(n34220), .B(n34216), .Z(n34289) );
  XNOR U34558 ( .A(n34215), .B(n34211), .Z(n34290) );
  XNOR U34559 ( .A(n34210), .B(n34206), .Z(n34291) );
  XNOR U34560 ( .A(n34205), .B(n34201), .Z(n34292) );
  XNOR U34561 ( .A(n34200), .B(n34196), .Z(n34293) );
  XNOR U34562 ( .A(n34195), .B(n34191), .Z(n34294) );
  XNOR U34563 ( .A(n34190), .B(n34186), .Z(n34295) );
  XNOR U34564 ( .A(n34185), .B(n34181), .Z(n34296) );
  XNOR U34565 ( .A(n34180), .B(n34176), .Z(n34297) );
  XNOR U34566 ( .A(n34298), .B(n34175), .Z(n34176) );
  AND U34567 ( .A(a[0]), .B(b[22]), .Z(n34298) );
  XNOR U34568 ( .A(n34299), .B(n34175), .Z(n34177) );
  XNOR U34569 ( .A(n34300), .B(n34301), .Z(n34175) );
  AND U34570 ( .A(n34302), .B(n34303), .Z(n34300) );
  AND U34571 ( .A(a[1]), .B(b[21]), .Z(n34299) );
  XOR U34572 ( .A(n34304), .B(n34180), .Z(n34182) );
  XOR U34573 ( .A(n34305), .B(n34306), .Z(n34180) );
  AND U34574 ( .A(n34307), .B(n34308), .Z(n34305) );
  AND U34575 ( .A(a[2]), .B(b[20]), .Z(n34304) );
  XOR U34576 ( .A(n34309), .B(n34185), .Z(n34187) );
  XOR U34577 ( .A(n34310), .B(n34311), .Z(n34185) );
  AND U34578 ( .A(n34312), .B(n34313), .Z(n34310) );
  AND U34579 ( .A(a[3]), .B(b[19]), .Z(n34309) );
  XOR U34580 ( .A(n34314), .B(n34190), .Z(n34192) );
  XOR U34581 ( .A(n34315), .B(n34316), .Z(n34190) );
  AND U34582 ( .A(n34317), .B(n34318), .Z(n34315) );
  AND U34583 ( .A(a[4]), .B(b[18]), .Z(n34314) );
  XOR U34584 ( .A(n34319), .B(n34195), .Z(n34197) );
  XOR U34585 ( .A(n34320), .B(n34321), .Z(n34195) );
  AND U34586 ( .A(n34322), .B(n34323), .Z(n34320) );
  AND U34587 ( .A(a[5]), .B(b[17]), .Z(n34319) );
  XOR U34588 ( .A(n34324), .B(n34200), .Z(n34202) );
  XOR U34589 ( .A(n34325), .B(n34326), .Z(n34200) );
  AND U34590 ( .A(n34327), .B(n34328), .Z(n34325) );
  AND U34591 ( .A(a[6]), .B(b[16]), .Z(n34324) );
  XOR U34592 ( .A(n34329), .B(n34205), .Z(n34207) );
  XOR U34593 ( .A(n34330), .B(n34331), .Z(n34205) );
  AND U34594 ( .A(n34332), .B(n34333), .Z(n34330) );
  AND U34595 ( .A(a[7]), .B(b[15]), .Z(n34329) );
  XOR U34596 ( .A(n34334), .B(n34210), .Z(n34212) );
  XOR U34597 ( .A(n34335), .B(n34336), .Z(n34210) );
  AND U34598 ( .A(n34337), .B(n34338), .Z(n34335) );
  AND U34599 ( .A(a[8]), .B(b[14]), .Z(n34334) );
  XOR U34600 ( .A(n34339), .B(n34215), .Z(n34217) );
  XOR U34601 ( .A(n34340), .B(n34341), .Z(n34215) );
  AND U34602 ( .A(n34342), .B(n34343), .Z(n34340) );
  AND U34603 ( .A(a[9]), .B(b[13]), .Z(n34339) );
  XOR U34604 ( .A(n34344), .B(n34220), .Z(n34222) );
  XOR U34605 ( .A(n34345), .B(n34346), .Z(n34220) );
  AND U34606 ( .A(n34347), .B(n34348), .Z(n34345) );
  AND U34607 ( .A(a[10]), .B(b[12]), .Z(n34344) );
  XOR U34608 ( .A(n34349), .B(n34225), .Z(n34227) );
  XOR U34609 ( .A(n34350), .B(n34351), .Z(n34225) );
  AND U34610 ( .A(n34352), .B(n34353), .Z(n34350) );
  AND U34611 ( .A(a[11]), .B(b[11]), .Z(n34349) );
  XOR U34612 ( .A(n34354), .B(n34230), .Z(n34232) );
  XOR U34613 ( .A(n34355), .B(n34356), .Z(n34230) );
  AND U34614 ( .A(n34357), .B(n34358), .Z(n34355) );
  AND U34615 ( .A(b[10]), .B(a[12]), .Z(n34354) );
  XOR U34616 ( .A(n34359), .B(n34235), .Z(n34237) );
  XOR U34617 ( .A(n34360), .B(n34361), .Z(n34235) );
  AND U34618 ( .A(n34362), .B(n34363), .Z(n34360) );
  AND U34619 ( .A(b[9]), .B(a[13]), .Z(n34359) );
  XOR U34620 ( .A(n34364), .B(n34240), .Z(n34242) );
  XOR U34621 ( .A(n34365), .B(n34366), .Z(n34240) );
  AND U34622 ( .A(n34367), .B(n34368), .Z(n34365) );
  AND U34623 ( .A(b[8]), .B(a[14]), .Z(n34364) );
  XOR U34624 ( .A(n34369), .B(n34245), .Z(n34247) );
  XOR U34625 ( .A(n34370), .B(n34371), .Z(n34245) );
  AND U34626 ( .A(n34372), .B(n34373), .Z(n34370) );
  AND U34627 ( .A(b[7]), .B(a[15]), .Z(n34369) );
  XOR U34628 ( .A(n34374), .B(n34250), .Z(n34252) );
  XOR U34629 ( .A(n34375), .B(n34376), .Z(n34250) );
  AND U34630 ( .A(n34377), .B(n34378), .Z(n34375) );
  AND U34631 ( .A(b[6]), .B(a[16]), .Z(n34374) );
  XOR U34632 ( .A(n34379), .B(n34255), .Z(n34257) );
  XOR U34633 ( .A(n34380), .B(n34381), .Z(n34255) );
  AND U34634 ( .A(n34382), .B(n34383), .Z(n34380) );
  AND U34635 ( .A(b[5]), .B(a[17]), .Z(n34379) );
  XOR U34636 ( .A(n34384), .B(n34260), .Z(n34262) );
  XOR U34637 ( .A(n34385), .B(n34386), .Z(n34260) );
  AND U34638 ( .A(n34387), .B(n34388), .Z(n34385) );
  AND U34639 ( .A(b[4]), .B(a[18]), .Z(n34384) );
  XNOR U34640 ( .A(n34389), .B(n34390), .Z(n34270) );
  NANDN U34641 ( .A(n34391), .B(n34392), .Z(n34390) );
  XOR U34642 ( .A(n34393), .B(n34265), .Z(n34267) );
  XNOR U34643 ( .A(n34394), .B(n34395), .Z(n34265) );
  AND U34644 ( .A(n34396), .B(n34397), .Z(n34394) );
  AND U34645 ( .A(b[3]), .B(a[19]), .Z(n34393) );
  NANDN U34646 ( .A(n31837), .B(n31835), .Z(n34274) );
  XNOR U34647 ( .A(n34391), .B(n34392), .Z(n31835) );
  XOR U34648 ( .A(n34389), .B(n34398), .Z(n34392) );
  NAND U34649 ( .A(b[1]), .B(a[20]), .Z(n34398) );
  XOR U34650 ( .A(n34397), .B(n34399), .Z(n34391) );
  XOR U34651 ( .A(n34389), .B(n34396), .Z(n34399) );
  XNOR U34652 ( .A(n34400), .B(n34395), .Z(n34396) );
  AND U34653 ( .A(b[2]), .B(a[19]), .Z(n34400) );
  NANDN U34654 ( .A(n31842), .B(n31840), .Z(n34389) );
  XNOR U34655 ( .A(n34401), .B(n34402), .Z(n31840) );
  NAND U34656 ( .A(a[20]), .B(b[0]), .Z(n31842) );
  XOR U34657 ( .A(n34395), .B(n34387), .Z(n34403) );
  XNOR U34658 ( .A(n34386), .B(n34382), .Z(n34404) );
  XNOR U34659 ( .A(n34381), .B(n34377), .Z(n34405) );
  XNOR U34660 ( .A(n34376), .B(n34372), .Z(n34406) );
  XNOR U34661 ( .A(n34371), .B(n34367), .Z(n34407) );
  XNOR U34662 ( .A(n34366), .B(n34362), .Z(n34408) );
  XNOR U34663 ( .A(n34361), .B(n34357), .Z(n34409) );
  XNOR U34664 ( .A(n34356), .B(n34352), .Z(n34410) );
  XNOR U34665 ( .A(n34351), .B(n34347), .Z(n34411) );
  XNOR U34666 ( .A(n34346), .B(n34342), .Z(n34412) );
  XNOR U34667 ( .A(n34341), .B(n34337), .Z(n34413) );
  XNOR U34668 ( .A(n34336), .B(n34332), .Z(n34414) );
  XNOR U34669 ( .A(n34331), .B(n34327), .Z(n34415) );
  XNOR U34670 ( .A(n34326), .B(n34322), .Z(n34416) );
  XNOR U34671 ( .A(n34321), .B(n34317), .Z(n34417) );
  XNOR U34672 ( .A(n34316), .B(n34312), .Z(n34418) );
  XNOR U34673 ( .A(n34311), .B(n34307), .Z(n34419) );
  XNOR U34674 ( .A(n34306), .B(n34302), .Z(n34420) );
  XOR U34675 ( .A(n34421), .B(n34301), .Z(n34302) );
  AND U34676 ( .A(a[0]), .B(b[21]), .Z(n34421) );
  XOR U34677 ( .A(n34422), .B(n34301), .Z(n34303) );
  XNOR U34678 ( .A(n34423), .B(n34424), .Z(n34301) );
  AND U34679 ( .A(n34425), .B(n34426), .Z(n34423) );
  AND U34680 ( .A(a[1]), .B(b[20]), .Z(n34422) );
  XOR U34681 ( .A(n34427), .B(n34306), .Z(n34308) );
  XOR U34682 ( .A(n34428), .B(n34429), .Z(n34306) );
  AND U34683 ( .A(n34430), .B(n34431), .Z(n34428) );
  AND U34684 ( .A(a[2]), .B(b[19]), .Z(n34427) );
  XOR U34685 ( .A(n34432), .B(n34311), .Z(n34313) );
  XOR U34686 ( .A(n34433), .B(n34434), .Z(n34311) );
  AND U34687 ( .A(n34435), .B(n34436), .Z(n34433) );
  AND U34688 ( .A(a[3]), .B(b[18]), .Z(n34432) );
  XOR U34689 ( .A(n34437), .B(n34316), .Z(n34318) );
  XOR U34690 ( .A(n34438), .B(n34439), .Z(n34316) );
  AND U34691 ( .A(n34440), .B(n34441), .Z(n34438) );
  AND U34692 ( .A(a[4]), .B(b[17]), .Z(n34437) );
  XOR U34693 ( .A(n34442), .B(n34321), .Z(n34323) );
  XOR U34694 ( .A(n34443), .B(n34444), .Z(n34321) );
  AND U34695 ( .A(n34445), .B(n34446), .Z(n34443) );
  AND U34696 ( .A(a[5]), .B(b[16]), .Z(n34442) );
  XOR U34697 ( .A(n34447), .B(n34326), .Z(n34328) );
  XOR U34698 ( .A(n34448), .B(n34449), .Z(n34326) );
  AND U34699 ( .A(n34450), .B(n34451), .Z(n34448) );
  AND U34700 ( .A(a[6]), .B(b[15]), .Z(n34447) );
  XOR U34701 ( .A(n34452), .B(n34331), .Z(n34333) );
  XOR U34702 ( .A(n34453), .B(n34454), .Z(n34331) );
  AND U34703 ( .A(n34455), .B(n34456), .Z(n34453) );
  AND U34704 ( .A(a[7]), .B(b[14]), .Z(n34452) );
  XOR U34705 ( .A(n34457), .B(n34336), .Z(n34338) );
  XOR U34706 ( .A(n34458), .B(n34459), .Z(n34336) );
  AND U34707 ( .A(n34460), .B(n34461), .Z(n34458) );
  AND U34708 ( .A(a[8]), .B(b[13]), .Z(n34457) );
  XOR U34709 ( .A(n34462), .B(n34341), .Z(n34343) );
  XOR U34710 ( .A(n34463), .B(n34464), .Z(n34341) );
  AND U34711 ( .A(n34465), .B(n34466), .Z(n34463) );
  AND U34712 ( .A(a[9]), .B(b[12]), .Z(n34462) );
  XOR U34713 ( .A(n34467), .B(n34346), .Z(n34348) );
  XOR U34714 ( .A(n34468), .B(n34469), .Z(n34346) );
  AND U34715 ( .A(n34470), .B(n34471), .Z(n34468) );
  AND U34716 ( .A(a[10]), .B(b[11]), .Z(n34467) );
  XOR U34717 ( .A(n34472), .B(n34351), .Z(n34353) );
  XOR U34718 ( .A(n34473), .B(n34474), .Z(n34351) );
  AND U34719 ( .A(n34475), .B(n34476), .Z(n34473) );
  AND U34720 ( .A(b[10]), .B(a[11]), .Z(n34472) );
  XOR U34721 ( .A(n34477), .B(n34356), .Z(n34358) );
  XOR U34722 ( .A(n34478), .B(n34479), .Z(n34356) );
  AND U34723 ( .A(n34480), .B(n34481), .Z(n34478) );
  AND U34724 ( .A(b[9]), .B(a[12]), .Z(n34477) );
  XOR U34725 ( .A(n34482), .B(n34361), .Z(n34363) );
  XOR U34726 ( .A(n34483), .B(n34484), .Z(n34361) );
  AND U34727 ( .A(n34485), .B(n34486), .Z(n34483) );
  AND U34728 ( .A(b[8]), .B(a[13]), .Z(n34482) );
  XOR U34729 ( .A(n34487), .B(n34366), .Z(n34368) );
  XOR U34730 ( .A(n34488), .B(n34489), .Z(n34366) );
  AND U34731 ( .A(n34490), .B(n34491), .Z(n34488) );
  AND U34732 ( .A(b[7]), .B(a[14]), .Z(n34487) );
  XOR U34733 ( .A(n34492), .B(n34371), .Z(n34373) );
  XOR U34734 ( .A(n34493), .B(n34494), .Z(n34371) );
  AND U34735 ( .A(n34495), .B(n34496), .Z(n34493) );
  AND U34736 ( .A(b[6]), .B(a[15]), .Z(n34492) );
  XOR U34737 ( .A(n34497), .B(n34376), .Z(n34378) );
  XOR U34738 ( .A(n34498), .B(n34499), .Z(n34376) );
  AND U34739 ( .A(n34500), .B(n34501), .Z(n34498) );
  AND U34740 ( .A(b[5]), .B(a[16]), .Z(n34497) );
  XOR U34741 ( .A(n34502), .B(n34381), .Z(n34383) );
  XOR U34742 ( .A(n34503), .B(n34504), .Z(n34381) );
  AND U34743 ( .A(n34505), .B(n34506), .Z(n34503) );
  AND U34744 ( .A(b[4]), .B(a[17]), .Z(n34502) );
  XNOR U34745 ( .A(n34507), .B(n34508), .Z(n34395) );
  NANDN U34746 ( .A(n34401), .B(n34402), .Z(n34508) );
  XOR U34747 ( .A(n34507), .B(n34509), .Z(n34402) );
  NAND U34748 ( .A(b[1]), .B(a[19]), .Z(n34509) );
  XOR U34749 ( .A(n34510), .B(n34511), .Z(n34401) );
  XOR U34750 ( .A(n34507), .B(n34512), .Z(n34511) );
  NANDN U34751 ( .A(n31847), .B(n31845), .Z(n34507) );
  XNOR U34752 ( .A(n34513), .B(n34514), .Z(n31845) );
  NAND U34753 ( .A(a[19]), .B(b[0]), .Z(n31847) );
  XOR U34754 ( .A(n34515), .B(n34386), .Z(n34388) );
  XNOR U34755 ( .A(n34516), .B(n34517), .Z(n34386) );
  AND U34756 ( .A(n34512), .B(n34510), .Z(n34516) );
  XOR U34757 ( .A(n34517), .B(n34505), .Z(n34518) );
  XNOR U34758 ( .A(n34504), .B(n34500), .Z(n34519) );
  XNOR U34759 ( .A(n34499), .B(n34495), .Z(n34520) );
  XNOR U34760 ( .A(n34494), .B(n34490), .Z(n34521) );
  XNOR U34761 ( .A(n34489), .B(n34485), .Z(n34522) );
  XNOR U34762 ( .A(n34484), .B(n34480), .Z(n34523) );
  XNOR U34763 ( .A(n34479), .B(n34475), .Z(n34524) );
  XNOR U34764 ( .A(n34474), .B(n34470), .Z(n34525) );
  XNOR U34765 ( .A(n34469), .B(n34465), .Z(n34526) );
  XNOR U34766 ( .A(n34464), .B(n34460), .Z(n34527) );
  XNOR U34767 ( .A(n34459), .B(n34455), .Z(n34528) );
  XNOR U34768 ( .A(n34454), .B(n34450), .Z(n34529) );
  XNOR U34769 ( .A(n34449), .B(n34445), .Z(n34530) );
  XNOR U34770 ( .A(n34444), .B(n34440), .Z(n34531) );
  XNOR U34771 ( .A(n34439), .B(n34435), .Z(n34532) );
  XNOR U34772 ( .A(n34434), .B(n34430), .Z(n34533) );
  XNOR U34773 ( .A(n34429), .B(n34425), .Z(n34534) );
  XNOR U34774 ( .A(n34535), .B(n34424), .Z(n34425) );
  AND U34775 ( .A(a[0]), .B(b[20]), .Z(n34535) );
  XNOR U34776 ( .A(n34536), .B(n34424), .Z(n34426) );
  XNOR U34777 ( .A(n34537), .B(n34538), .Z(n34424) );
  AND U34778 ( .A(n34539), .B(n34540), .Z(n34537) );
  AND U34779 ( .A(a[1]), .B(b[19]), .Z(n34536) );
  XOR U34780 ( .A(n34541), .B(n34429), .Z(n34431) );
  XOR U34781 ( .A(n34542), .B(n34543), .Z(n34429) );
  AND U34782 ( .A(n34544), .B(n34545), .Z(n34542) );
  AND U34783 ( .A(a[2]), .B(b[18]), .Z(n34541) );
  XOR U34784 ( .A(n34546), .B(n34434), .Z(n34436) );
  XOR U34785 ( .A(n34547), .B(n34548), .Z(n34434) );
  AND U34786 ( .A(n34549), .B(n34550), .Z(n34547) );
  AND U34787 ( .A(a[3]), .B(b[17]), .Z(n34546) );
  XOR U34788 ( .A(n34551), .B(n34439), .Z(n34441) );
  XOR U34789 ( .A(n34552), .B(n34553), .Z(n34439) );
  AND U34790 ( .A(n34554), .B(n34555), .Z(n34552) );
  AND U34791 ( .A(a[4]), .B(b[16]), .Z(n34551) );
  XOR U34792 ( .A(n34556), .B(n34444), .Z(n34446) );
  XOR U34793 ( .A(n34557), .B(n34558), .Z(n34444) );
  AND U34794 ( .A(n34559), .B(n34560), .Z(n34557) );
  AND U34795 ( .A(a[5]), .B(b[15]), .Z(n34556) );
  XOR U34796 ( .A(n34561), .B(n34449), .Z(n34451) );
  XOR U34797 ( .A(n34562), .B(n34563), .Z(n34449) );
  AND U34798 ( .A(n34564), .B(n34565), .Z(n34562) );
  AND U34799 ( .A(a[6]), .B(b[14]), .Z(n34561) );
  XOR U34800 ( .A(n34566), .B(n34454), .Z(n34456) );
  XOR U34801 ( .A(n34567), .B(n34568), .Z(n34454) );
  AND U34802 ( .A(n34569), .B(n34570), .Z(n34567) );
  AND U34803 ( .A(a[7]), .B(b[13]), .Z(n34566) );
  XOR U34804 ( .A(n34571), .B(n34459), .Z(n34461) );
  XOR U34805 ( .A(n34572), .B(n34573), .Z(n34459) );
  AND U34806 ( .A(n34574), .B(n34575), .Z(n34572) );
  AND U34807 ( .A(a[8]), .B(b[12]), .Z(n34571) );
  XOR U34808 ( .A(n34576), .B(n34464), .Z(n34466) );
  XOR U34809 ( .A(n34577), .B(n34578), .Z(n34464) );
  AND U34810 ( .A(n34579), .B(n34580), .Z(n34577) );
  AND U34811 ( .A(a[9]), .B(b[11]), .Z(n34576) );
  XOR U34812 ( .A(n34581), .B(n34469), .Z(n34471) );
  XOR U34813 ( .A(n34582), .B(n34583), .Z(n34469) );
  AND U34814 ( .A(n34584), .B(n34585), .Z(n34582) );
  AND U34815 ( .A(a[10]), .B(b[10]), .Z(n34581) );
  XOR U34816 ( .A(n34586), .B(n34474), .Z(n34476) );
  XOR U34817 ( .A(n34587), .B(n34588), .Z(n34474) );
  AND U34818 ( .A(n34589), .B(n34590), .Z(n34587) );
  AND U34819 ( .A(b[9]), .B(a[11]), .Z(n34586) );
  XOR U34820 ( .A(n34591), .B(n34479), .Z(n34481) );
  XOR U34821 ( .A(n34592), .B(n34593), .Z(n34479) );
  AND U34822 ( .A(n34594), .B(n34595), .Z(n34592) );
  AND U34823 ( .A(b[8]), .B(a[12]), .Z(n34591) );
  XOR U34824 ( .A(n34596), .B(n34484), .Z(n34486) );
  XOR U34825 ( .A(n34597), .B(n34598), .Z(n34484) );
  AND U34826 ( .A(n34599), .B(n34600), .Z(n34597) );
  AND U34827 ( .A(b[7]), .B(a[13]), .Z(n34596) );
  XOR U34828 ( .A(n34601), .B(n34489), .Z(n34491) );
  XOR U34829 ( .A(n34602), .B(n34603), .Z(n34489) );
  AND U34830 ( .A(n34604), .B(n34605), .Z(n34602) );
  AND U34831 ( .A(b[6]), .B(a[14]), .Z(n34601) );
  XOR U34832 ( .A(n34606), .B(n34494), .Z(n34496) );
  XOR U34833 ( .A(n34607), .B(n34608), .Z(n34494) );
  AND U34834 ( .A(n34609), .B(n34610), .Z(n34607) );
  AND U34835 ( .A(b[5]), .B(a[15]), .Z(n34606) );
  XOR U34836 ( .A(n34611), .B(n34499), .Z(n34501) );
  XOR U34837 ( .A(n34612), .B(n34613), .Z(n34499) );
  AND U34838 ( .A(n34614), .B(n34615), .Z(n34612) );
  AND U34839 ( .A(b[4]), .B(a[16]), .Z(n34611) );
  XOR U34840 ( .A(n34616), .B(n34504), .Z(n34506) );
  XNOR U34841 ( .A(n34617), .B(n34618), .Z(n34504) );
  AND U34842 ( .A(n34619), .B(n34620), .Z(n34617) );
  AND U34843 ( .A(b[3]), .B(a[17]), .Z(n34616) );
  XNOR U34844 ( .A(n34621), .B(n34517), .Z(n34512) );
  XNOR U34845 ( .A(n34622), .B(n34623), .Z(n34517) );
  NANDN U34846 ( .A(n34513), .B(n34514), .Z(n34623) );
  XOR U34847 ( .A(n34622), .B(n34624), .Z(n34514) );
  NAND U34848 ( .A(b[1]), .B(a[18]), .Z(n34624) );
  XOR U34849 ( .A(n34620), .B(n34625), .Z(n34513) );
  XOR U34850 ( .A(n34622), .B(n34619), .Z(n34625) );
  XNOR U34851 ( .A(n34626), .B(n34618), .Z(n34619) );
  AND U34852 ( .A(b[2]), .B(a[17]), .Z(n34626) );
  XOR U34853 ( .A(n34618), .B(n34614), .Z(n34627) );
  XNOR U34854 ( .A(n34613), .B(n34609), .Z(n34628) );
  XNOR U34855 ( .A(n34608), .B(n34604), .Z(n34629) );
  XNOR U34856 ( .A(n34603), .B(n34599), .Z(n34630) );
  XNOR U34857 ( .A(n34598), .B(n34594), .Z(n34631) );
  XNOR U34858 ( .A(n34593), .B(n34589), .Z(n34632) );
  XNOR U34859 ( .A(n34588), .B(n34584), .Z(n34633) );
  XNOR U34860 ( .A(n34583), .B(n34579), .Z(n34634) );
  XNOR U34861 ( .A(n34578), .B(n34574), .Z(n34635) );
  XNOR U34862 ( .A(n34573), .B(n34569), .Z(n34636) );
  XNOR U34863 ( .A(n34568), .B(n34564), .Z(n34637) );
  XNOR U34864 ( .A(n34563), .B(n34559), .Z(n34638) );
  XNOR U34865 ( .A(n34558), .B(n34554), .Z(n34639) );
  XNOR U34866 ( .A(n34553), .B(n34549), .Z(n34640) );
  XNOR U34867 ( .A(n34548), .B(n34544), .Z(n34641) );
  XNOR U34868 ( .A(n34543), .B(n34539), .Z(n34642) );
  XOR U34869 ( .A(n34643), .B(n34538), .Z(n34539) );
  AND U34870 ( .A(a[0]), .B(b[19]), .Z(n34643) );
  XOR U34871 ( .A(n34644), .B(n34538), .Z(n34540) );
  XNOR U34872 ( .A(n34645), .B(n34646), .Z(n34538) );
  AND U34873 ( .A(n34647), .B(n34648), .Z(n34645) );
  AND U34874 ( .A(a[1]), .B(b[18]), .Z(n34644) );
  XOR U34875 ( .A(n34649), .B(n34543), .Z(n34545) );
  XOR U34876 ( .A(n34650), .B(n34651), .Z(n34543) );
  AND U34877 ( .A(n34652), .B(n34653), .Z(n34650) );
  AND U34878 ( .A(a[2]), .B(b[17]), .Z(n34649) );
  XOR U34879 ( .A(n34654), .B(n34548), .Z(n34550) );
  XOR U34880 ( .A(n34655), .B(n34656), .Z(n34548) );
  AND U34881 ( .A(n34657), .B(n34658), .Z(n34655) );
  AND U34882 ( .A(a[3]), .B(b[16]), .Z(n34654) );
  XOR U34883 ( .A(n34659), .B(n34553), .Z(n34555) );
  XOR U34884 ( .A(n34660), .B(n34661), .Z(n34553) );
  AND U34885 ( .A(n34662), .B(n34663), .Z(n34660) );
  AND U34886 ( .A(a[4]), .B(b[15]), .Z(n34659) );
  XOR U34887 ( .A(n34664), .B(n34558), .Z(n34560) );
  XOR U34888 ( .A(n34665), .B(n34666), .Z(n34558) );
  AND U34889 ( .A(n34667), .B(n34668), .Z(n34665) );
  AND U34890 ( .A(a[5]), .B(b[14]), .Z(n34664) );
  XOR U34891 ( .A(n34669), .B(n34563), .Z(n34565) );
  XOR U34892 ( .A(n34670), .B(n34671), .Z(n34563) );
  AND U34893 ( .A(n34672), .B(n34673), .Z(n34670) );
  AND U34894 ( .A(a[6]), .B(b[13]), .Z(n34669) );
  XOR U34895 ( .A(n34674), .B(n34568), .Z(n34570) );
  XOR U34896 ( .A(n34675), .B(n34676), .Z(n34568) );
  AND U34897 ( .A(n34677), .B(n34678), .Z(n34675) );
  AND U34898 ( .A(a[7]), .B(b[12]), .Z(n34674) );
  XOR U34899 ( .A(n34679), .B(n34573), .Z(n34575) );
  XOR U34900 ( .A(n34680), .B(n34681), .Z(n34573) );
  AND U34901 ( .A(n34682), .B(n34683), .Z(n34680) );
  AND U34902 ( .A(a[8]), .B(b[11]), .Z(n34679) );
  XOR U34903 ( .A(n34684), .B(n34578), .Z(n34580) );
  XOR U34904 ( .A(n34685), .B(n34686), .Z(n34578) );
  AND U34905 ( .A(n34687), .B(n34688), .Z(n34685) );
  AND U34906 ( .A(a[9]), .B(b[10]), .Z(n34684) );
  XOR U34907 ( .A(n34689), .B(n34583), .Z(n34585) );
  XOR U34908 ( .A(n34690), .B(n34691), .Z(n34583) );
  AND U34909 ( .A(n34692), .B(n34693), .Z(n34690) );
  AND U34910 ( .A(b[9]), .B(a[10]), .Z(n34689) );
  XOR U34911 ( .A(n34694), .B(n34588), .Z(n34590) );
  XOR U34912 ( .A(n34695), .B(n34696), .Z(n34588) );
  AND U34913 ( .A(n34697), .B(n34698), .Z(n34695) );
  AND U34914 ( .A(b[8]), .B(a[11]), .Z(n34694) );
  XOR U34915 ( .A(n34699), .B(n34593), .Z(n34595) );
  XOR U34916 ( .A(n34700), .B(n34701), .Z(n34593) );
  AND U34917 ( .A(n34702), .B(n34703), .Z(n34700) );
  AND U34918 ( .A(b[7]), .B(a[12]), .Z(n34699) );
  XOR U34919 ( .A(n34704), .B(n34598), .Z(n34600) );
  XOR U34920 ( .A(n34705), .B(n34706), .Z(n34598) );
  AND U34921 ( .A(n34707), .B(n34708), .Z(n34705) );
  AND U34922 ( .A(b[6]), .B(a[13]), .Z(n34704) );
  XOR U34923 ( .A(n34709), .B(n34603), .Z(n34605) );
  XOR U34924 ( .A(n34710), .B(n34711), .Z(n34603) );
  AND U34925 ( .A(n34712), .B(n34713), .Z(n34710) );
  AND U34926 ( .A(b[5]), .B(a[14]), .Z(n34709) );
  XOR U34927 ( .A(n34714), .B(n34608), .Z(n34610) );
  XOR U34928 ( .A(n34715), .B(n34716), .Z(n34608) );
  AND U34929 ( .A(n34717), .B(n34718), .Z(n34715) );
  AND U34930 ( .A(b[4]), .B(a[15]), .Z(n34714) );
  XNOR U34931 ( .A(n34719), .B(n34720), .Z(n34618) );
  NANDN U34932 ( .A(n34721), .B(n34722), .Z(n34720) );
  XOR U34933 ( .A(n34723), .B(n34613), .Z(n34615) );
  XNOR U34934 ( .A(n34724), .B(n34725), .Z(n34613) );
  AND U34935 ( .A(n34726), .B(n34727), .Z(n34724) );
  AND U34936 ( .A(b[3]), .B(a[16]), .Z(n34723) );
  NANDN U34937 ( .A(n31852), .B(n31850), .Z(n34622) );
  XNOR U34938 ( .A(n34721), .B(n34722), .Z(n31850) );
  XOR U34939 ( .A(n34719), .B(n34728), .Z(n34722) );
  NAND U34940 ( .A(b[1]), .B(a[17]), .Z(n34728) );
  XOR U34941 ( .A(n34727), .B(n34729), .Z(n34721) );
  XOR U34942 ( .A(n34719), .B(n34726), .Z(n34729) );
  XNOR U34943 ( .A(n34730), .B(n34725), .Z(n34726) );
  AND U34944 ( .A(b[2]), .B(a[16]), .Z(n34730) );
  NANDN U34945 ( .A(n31857), .B(n31855), .Z(n34719) );
  XNOR U34946 ( .A(n34731), .B(n34732), .Z(n31855) );
  NAND U34947 ( .A(a[17]), .B(b[0]), .Z(n31857) );
  XOR U34948 ( .A(n34725), .B(n34717), .Z(n34733) );
  XNOR U34949 ( .A(n34716), .B(n34712), .Z(n34734) );
  XNOR U34950 ( .A(n34711), .B(n34707), .Z(n34735) );
  XNOR U34951 ( .A(n34706), .B(n34702), .Z(n34736) );
  XNOR U34952 ( .A(n34701), .B(n34697), .Z(n34737) );
  XNOR U34953 ( .A(n34696), .B(n34692), .Z(n34738) );
  XNOR U34954 ( .A(n34691), .B(n34687), .Z(n34739) );
  XNOR U34955 ( .A(n34686), .B(n34682), .Z(n34740) );
  XNOR U34956 ( .A(n34681), .B(n34677), .Z(n34741) );
  XNOR U34957 ( .A(n34676), .B(n34672), .Z(n34742) );
  XNOR U34958 ( .A(n34671), .B(n34667), .Z(n34743) );
  XNOR U34959 ( .A(n34666), .B(n34662), .Z(n34744) );
  XNOR U34960 ( .A(n34661), .B(n34657), .Z(n34745) );
  XNOR U34961 ( .A(n34656), .B(n34652), .Z(n34746) );
  XNOR U34962 ( .A(n34651), .B(n34647), .Z(n34747) );
  XNOR U34963 ( .A(n34748), .B(n34646), .Z(n34647) );
  AND U34964 ( .A(a[0]), .B(b[18]), .Z(n34748) );
  XNOR U34965 ( .A(n34749), .B(n34646), .Z(n34648) );
  XNOR U34966 ( .A(n34750), .B(n34751), .Z(n34646) );
  AND U34967 ( .A(n34752), .B(n34753), .Z(n34750) );
  AND U34968 ( .A(a[1]), .B(b[17]), .Z(n34749) );
  XOR U34969 ( .A(n34754), .B(n34651), .Z(n34653) );
  XOR U34970 ( .A(n34755), .B(n34756), .Z(n34651) );
  AND U34971 ( .A(n34757), .B(n34758), .Z(n34755) );
  AND U34972 ( .A(a[2]), .B(b[16]), .Z(n34754) );
  XOR U34973 ( .A(n34759), .B(n34656), .Z(n34658) );
  XOR U34974 ( .A(n34760), .B(n34761), .Z(n34656) );
  AND U34975 ( .A(n34762), .B(n34763), .Z(n34760) );
  AND U34976 ( .A(a[3]), .B(b[15]), .Z(n34759) );
  XOR U34977 ( .A(n34764), .B(n34661), .Z(n34663) );
  XOR U34978 ( .A(n34765), .B(n34766), .Z(n34661) );
  AND U34979 ( .A(n34767), .B(n34768), .Z(n34765) );
  AND U34980 ( .A(a[4]), .B(b[14]), .Z(n34764) );
  XOR U34981 ( .A(n34769), .B(n34666), .Z(n34668) );
  XOR U34982 ( .A(n34770), .B(n34771), .Z(n34666) );
  AND U34983 ( .A(n34772), .B(n34773), .Z(n34770) );
  AND U34984 ( .A(a[5]), .B(b[13]), .Z(n34769) );
  XOR U34985 ( .A(n34774), .B(n34671), .Z(n34673) );
  XOR U34986 ( .A(n34775), .B(n34776), .Z(n34671) );
  AND U34987 ( .A(n34777), .B(n34778), .Z(n34775) );
  AND U34988 ( .A(a[6]), .B(b[12]), .Z(n34774) );
  XOR U34989 ( .A(n34779), .B(n34676), .Z(n34678) );
  XOR U34990 ( .A(n34780), .B(n34781), .Z(n34676) );
  AND U34991 ( .A(n34782), .B(n34783), .Z(n34780) );
  AND U34992 ( .A(a[7]), .B(b[11]), .Z(n34779) );
  XOR U34993 ( .A(n34784), .B(n34681), .Z(n34683) );
  XOR U34994 ( .A(n34785), .B(n34786), .Z(n34681) );
  AND U34995 ( .A(n34787), .B(n34788), .Z(n34785) );
  AND U34996 ( .A(a[8]), .B(b[10]), .Z(n34784) );
  XOR U34997 ( .A(n34789), .B(n34686), .Z(n34688) );
  XOR U34998 ( .A(n34790), .B(n34791), .Z(n34686) );
  AND U34999 ( .A(n34792), .B(n34793), .Z(n34790) );
  AND U35000 ( .A(a[9]), .B(b[9]), .Z(n34789) );
  XOR U35001 ( .A(n34794), .B(n34691), .Z(n34693) );
  XOR U35002 ( .A(n34795), .B(n34796), .Z(n34691) );
  AND U35003 ( .A(n34797), .B(n34798), .Z(n34795) );
  AND U35004 ( .A(b[8]), .B(a[10]), .Z(n34794) );
  XOR U35005 ( .A(n34799), .B(n34696), .Z(n34698) );
  XOR U35006 ( .A(n34800), .B(n34801), .Z(n34696) );
  AND U35007 ( .A(n34802), .B(n34803), .Z(n34800) );
  AND U35008 ( .A(b[7]), .B(a[11]), .Z(n34799) );
  XOR U35009 ( .A(n34804), .B(n34701), .Z(n34703) );
  XOR U35010 ( .A(n34805), .B(n34806), .Z(n34701) );
  AND U35011 ( .A(n34807), .B(n34808), .Z(n34805) );
  AND U35012 ( .A(b[6]), .B(a[12]), .Z(n34804) );
  XOR U35013 ( .A(n34809), .B(n34706), .Z(n34708) );
  XOR U35014 ( .A(n34810), .B(n34811), .Z(n34706) );
  AND U35015 ( .A(n34812), .B(n34813), .Z(n34810) );
  AND U35016 ( .A(b[5]), .B(a[13]), .Z(n34809) );
  XOR U35017 ( .A(n34814), .B(n34711), .Z(n34713) );
  XOR U35018 ( .A(n34815), .B(n34816), .Z(n34711) );
  AND U35019 ( .A(n34817), .B(n34818), .Z(n34815) );
  AND U35020 ( .A(b[4]), .B(a[14]), .Z(n34814) );
  XNOR U35021 ( .A(n34819), .B(n34820), .Z(n34725) );
  NANDN U35022 ( .A(n34731), .B(n34732), .Z(n34820) );
  XOR U35023 ( .A(n34819), .B(n34821), .Z(n34732) );
  NAND U35024 ( .A(b[1]), .B(a[16]), .Z(n34821) );
  XOR U35025 ( .A(n34822), .B(n34823), .Z(n34731) );
  XOR U35026 ( .A(n34819), .B(n34824), .Z(n34823) );
  NANDN U35027 ( .A(n31862), .B(n31860), .Z(n34819) );
  XNOR U35028 ( .A(n34825), .B(n34826), .Z(n31860) );
  NAND U35029 ( .A(a[16]), .B(b[0]), .Z(n31862) );
  XOR U35030 ( .A(n34827), .B(n34716), .Z(n34718) );
  XNOR U35031 ( .A(n34828), .B(n34829), .Z(n34716) );
  AND U35032 ( .A(n34824), .B(n34822), .Z(n34828) );
  XOR U35033 ( .A(n34829), .B(n34817), .Z(n34830) );
  XNOR U35034 ( .A(n34816), .B(n34812), .Z(n34831) );
  XNOR U35035 ( .A(n34811), .B(n34807), .Z(n34832) );
  XNOR U35036 ( .A(n34806), .B(n34802), .Z(n34833) );
  XNOR U35037 ( .A(n34801), .B(n34797), .Z(n34834) );
  XNOR U35038 ( .A(n34796), .B(n34792), .Z(n34835) );
  XNOR U35039 ( .A(n34791), .B(n34787), .Z(n34836) );
  XNOR U35040 ( .A(n34786), .B(n34782), .Z(n34837) );
  XNOR U35041 ( .A(n34781), .B(n34777), .Z(n34838) );
  XNOR U35042 ( .A(n34776), .B(n34772), .Z(n34839) );
  XNOR U35043 ( .A(n34771), .B(n34767), .Z(n34840) );
  XNOR U35044 ( .A(n34766), .B(n34762), .Z(n34841) );
  XNOR U35045 ( .A(n34761), .B(n34757), .Z(n34842) );
  XNOR U35046 ( .A(n34756), .B(n34752), .Z(n34843) );
  XOR U35047 ( .A(n34844), .B(n34751), .Z(n34752) );
  AND U35048 ( .A(a[0]), .B(b[17]), .Z(n34844) );
  XOR U35049 ( .A(n34845), .B(n34751), .Z(n34753) );
  XNOR U35050 ( .A(n34846), .B(n34847), .Z(n34751) );
  AND U35051 ( .A(n34848), .B(n34849), .Z(n34846) );
  AND U35052 ( .A(a[1]), .B(b[16]), .Z(n34845) );
  XOR U35053 ( .A(n34850), .B(n34756), .Z(n34758) );
  XOR U35054 ( .A(n34851), .B(n34852), .Z(n34756) );
  AND U35055 ( .A(n34853), .B(n34854), .Z(n34851) );
  AND U35056 ( .A(a[2]), .B(b[15]), .Z(n34850) );
  XOR U35057 ( .A(n34855), .B(n34761), .Z(n34763) );
  XOR U35058 ( .A(n34856), .B(n34857), .Z(n34761) );
  AND U35059 ( .A(n34858), .B(n34859), .Z(n34856) );
  AND U35060 ( .A(a[3]), .B(b[14]), .Z(n34855) );
  XOR U35061 ( .A(n34860), .B(n34766), .Z(n34768) );
  XOR U35062 ( .A(n34861), .B(n34862), .Z(n34766) );
  AND U35063 ( .A(n34863), .B(n34864), .Z(n34861) );
  AND U35064 ( .A(a[4]), .B(b[13]), .Z(n34860) );
  XOR U35065 ( .A(n34865), .B(n34771), .Z(n34773) );
  XOR U35066 ( .A(n34866), .B(n34867), .Z(n34771) );
  AND U35067 ( .A(n34868), .B(n34869), .Z(n34866) );
  AND U35068 ( .A(a[5]), .B(b[12]), .Z(n34865) );
  XOR U35069 ( .A(n34870), .B(n34776), .Z(n34778) );
  XOR U35070 ( .A(n34871), .B(n34872), .Z(n34776) );
  AND U35071 ( .A(n34873), .B(n34874), .Z(n34871) );
  AND U35072 ( .A(a[6]), .B(b[11]), .Z(n34870) );
  XOR U35073 ( .A(n34875), .B(n34781), .Z(n34783) );
  XOR U35074 ( .A(n34876), .B(n34877), .Z(n34781) );
  AND U35075 ( .A(n34878), .B(n34879), .Z(n34876) );
  AND U35076 ( .A(a[7]), .B(b[10]), .Z(n34875) );
  XOR U35077 ( .A(n34880), .B(n34786), .Z(n34788) );
  XOR U35078 ( .A(n34881), .B(n34882), .Z(n34786) );
  AND U35079 ( .A(n34883), .B(n34884), .Z(n34881) );
  AND U35080 ( .A(a[8]), .B(b[9]), .Z(n34880) );
  XOR U35081 ( .A(n34885), .B(n34791), .Z(n34793) );
  XOR U35082 ( .A(n34886), .B(n34887), .Z(n34791) );
  AND U35083 ( .A(n34888), .B(n34889), .Z(n34886) );
  AND U35084 ( .A(b[8]), .B(a[9]), .Z(n34885) );
  XOR U35085 ( .A(n34890), .B(n34796), .Z(n34798) );
  XOR U35086 ( .A(n34891), .B(n34892), .Z(n34796) );
  AND U35087 ( .A(n34893), .B(n34894), .Z(n34891) );
  AND U35088 ( .A(b[7]), .B(a[10]), .Z(n34890) );
  XOR U35089 ( .A(n34895), .B(n34801), .Z(n34803) );
  XOR U35090 ( .A(n34896), .B(n34897), .Z(n34801) );
  AND U35091 ( .A(n34898), .B(n34899), .Z(n34896) );
  AND U35092 ( .A(b[6]), .B(a[11]), .Z(n34895) );
  XOR U35093 ( .A(n34900), .B(n34806), .Z(n34808) );
  XOR U35094 ( .A(n34901), .B(n34902), .Z(n34806) );
  AND U35095 ( .A(n34903), .B(n34904), .Z(n34901) );
  AND U35096 ( .A(b[5]), .B(a[12]), .Z(n34900) );
  XOR U35097 ( .A(n34905), .B(n34811), .Z(n34813) );
  XOR U35098 ( .A(n34906), .B(n34907), .Z(n34811) );
  AND U35099 ( .A(n34908), .B(n34909), .Z(n34906) );
  AND U35100 ( .A(b[4]), .B(a[13]), .Z(n34905) );
  XOR U35101 ( .A(n34910), .B(n34816), .Z(n34818) );
  XNOR U35102 ( .A(n34911), .B(n34912), .Z(n34816) );
  AND U35103 ( .A(n34913), .B(n34914), .Z(n34911) );
  AND U35104 ( .A(b[3]), .B(a[14]), .Z(n34910) );
  XNOR U35105 ( .A(n34915), .B(n34829), .Z(n34824) );
  XNOR U35106 ( .A(n34916), .B(n34917), .Z(n34829) );
  NANDN U35107 ( .A(n34825), .B(n34826), .Z(n34917) );
  XOR U35108 ( .A(n34916), .B(n34918), .Z(n34826) );
  NAND U35109 ( .A(b[1]), .B(a[15]), .Z(n34918) );
  XOR U35110 ( .A(n34914), .B(n34919), .Z(n34825) );
  XOR U35111 ( .A(n34916), .B(n34913), .Z(n34919) );
  XNOR U35112 ( .A(n34920), .B(n34912), .Z(n34913) );
  AND U35113 ( .A(b[2]), .B(a[14]), .Z(n34920) );
  XOR U35114 ( .A(n34912), .B(n34908), .Z(n34921) );
  XNOR U35115 ( .A(n34907), .B(n34903), .Z(n34922) );
  XNOR U35116 ( .A(n34902), .B(n34898), .Z(n34923) );
  XNOR U35117 ( .A(n34897), .B(n34893), .Z(n34924) );
  XNOR U35118 ( .A(n34892), .B(n34888), .Z(n34925) );
  XNOR U35119 ( .A(n34887), .B(n34883), .Z(n34926) );
  XNOR U35120 ( .A(n34882), .B(n34878), .Z(n34927) );
  XNOR U35121 ( .A(n34877), .B(n34873), .Z(n34928) );
  XNOR U35122 ( .A(n34872), .B(n34868), .Z(n34929) );
  XNOR U35123 ( .A(n34867), .B(n34863), .Z(n34930) );
  XNOR U35124 ( .A(n34862), .B(n34858), .Z(n34931) );
  XNOR U35125 ( .A(n34857), .B(n34853), .Z(n34932) );
  XNOR U35126 ( .A(n34852), .B(n34848), .Z(n34933) );
  XNOR U35127 ( .A(n34934), .B(n34847), .Z(n34848) );
  AND U35128 ( .A(a[0]), .B(b[16]), .Z(n34934) );
  XNOR U35129 ( .A(n34935), .B(n34847), .Z(n34849) );
  XNOR U35130 ( .A(n34936), .B(n34937), .Z(n34847) );
  AND U35131 ( .A(n34938), .B(n34939), .Z(n34936) );
  AND U35132 ( .A(a[1]), .B(b[15]), .Z(n34935) );
  XOR U35133 ( .A(n34940), .B(n34852), .Z(n34854) );
  XOR U35134 ( .A(n34941), .B(n34942), .Z(n34852) );
  AND U35135 ( .A(n34943), .B(n34944), .Z(n34941) );
  AND U35136 ( .A(a[2]), .B(b[14]), .Z(n34940) );
  XOR U35137 ( .A(n34945), .B(n34857), .Z(n34859) );
  XOR U35138 ( .A(n34946), .B(n34947), .Z(n34857) );
  AND U35139 ( .A(n34948), .B(n34949), .Z(n34946) );
  AND U35140 ( .A(a[3]), .B(b[13]), .Z(n34945) );
  XOR U35141 ( .A(n34950), .B(n34862), .Z(n34864) );
  XOR U35142 ( .A(n34951), .B(n34952), .Z(n34862) );
  AND U35143 ( .A(n34953), .B(n34954), .Z(n34951) );
  AND U35144 ( .A(a[4]), .B(b[12]), .Z(n34950) );
  XOR U35145 ( .A(n34955), .B(n34867), .Z(n34869) );
  XOR U35146 ( .A(n34956), .B(n34957), .Z(n34867) );
  AND U35147 ( .A(n34958), .B(n34959), .Z(n34956) );
  AND U35148 ( .A(a[5]), .B(b[11]), .Z(n34955) );
  XOR U35149 ( .A(n34960), .B(n34872), .Z(n34874) );
  XOR U35150 ( .A(n34961), .B(n34962), .Z(n34872) );
  AND U35151 ( .A(n34963), .B(n34964), .Z(n34961) );
  AND U35152 ( .A(a[6]), .B(b[10]), .Z(n34960) );
  XOR U35153 ( .A(n34965), .B(n34877), .Z(n34879) );
  XOR U35154 ( .A(n34966), .B(n34967), .Z(n34877) );
  AND U35155 ( .A(n34968), .B(n34969), .Z(n34966) );
  AND U35156 ( .A(a[7]), .B(b[9]), .Z(n34965) );
  XOR U35157 ( .A(n34970), .B(n34882), .Z(n34884) );
  XOR U35158 ( .A(n34971), .B(n34972), .Z(n34882) );
  AND U35159 ( .A(n34973), .B(n34974), .Z(n34971) );
  AND U35160 ( .A(a[8]), .B(b[8]), .Z(n34970) );
  XOR U35161 ( .A(n34975), .B(n34887), .Z(n34889) );
  XOR U35162 ( .A(n34976), .B(n34977), .Z(n34887) );
  AND U35163 ( .A(n34978), .B(n34979), .Z(n34976) );
  AND U35164 ( .A(b[7]), .B(a[9]), .Z(n34975) );
  XOR U35165 ( .A(n34980), .B(n34892), .Z(n34894) );
  XOR U35166 ( .A(n34981), .B(n34982), .Z(n34892) );
  AND U35167 ( .A(n34983), .B(n34984), .Z(n34981) );
  AND U35168 ( .A(b[6]), .B(a[10]), .Z(n34980) );
  XOR U35169 ( .A(n34985), .B(n34897), .Z(n34899) );
  XOR U35170 ( .A(n34986), .B(n34987), .Z(n34897) );
  AND U35171 ( .A(n34988), .B(n34989), .Z(n34986) );
  AND U35172 ( .A(b[5]), .B(a[11]), .Z(n34985) );
  XOR U35173 ( .A(n34990), .B(n34902), .Z(n34904) );
  XOR U35174 ( .A(n34991), .B(n34992), .Z(n34902) );
  AND U35175 ( .A(n34993), .B(n34994), .Z(n34991) );
  AND U35176 ( .A(b[4]), .B(a[12]), .Z(n34990) );
  XNOR U35177 ( .A(n34995), .B(n34996), .Z(n34912) );
  NANDN U35178 ( .A(n34997), .B(n34998), .Z(n34996) );
  XOR U35179 ( .A(n34999), .B(n34907), .Z(n34909) );
  XNOR U35180 ( .A(n35000), .B(n35001), .Z(n34907) );
  AND U35181 ( .A(n35002), .B(n35003), .Z(n35000) );
  AND U35182 ( .A(b[3]), .B(a[13]), .Z(n34999) );
  NANDN U35183 ( .A(n31867), .B(n31865), .Z(n34916) );
  XNOR U35184 ( .A(n34997), .B(n34998), .Z(n31865) );
  XOR U35185 ( .A(n34995), .B(n35004), .Z(n34998) );
  NAND U35186 ( .A(b[1]), .B(a[14]), .Z(n35004) );
  XOR U35187 ( .A(n35003), .B(n35005), .Z(n34997) );
  XOR U35188 ( .A(n34995), .B(n35002), .Z(n35005) );
  XNOR U35189 ( .A(n35006), .B(n35001), .Z(n35002) );
  AND U35190 ( .A(b[2]), .B(a[13]), .Z(n35006) );
  NANDN U35191 ( .A(n31872), .B(n31870), .Z(n34995) );
  XNOR U35192 ( .A(n35007), .B(n35008), .Z(n31870) );
  NAND U35193 ( .A(a[14]), .B(b[0]), .Z(n31872) );
  XOR U35194 ( .A(n35001), .B(n34993), .Z(n35009) );
  XNOR U35195 ( .A(n34992), .B(n34988), .Z(n35010) );
  XNOR U35196 ( .A(n34987), .B(n34983), .Z(n35011) );
  XNOR U35197 ( .A(n34982), .B(n34978), .Z(n35012) );
  XNOR U35198 ( .A(n34977), .B(n34973), .Z(n35013) );
  XNOR U35199 ( .A(n34972), .B(n34968), .Z(n35014) );
  XNOR U35200 ( .A(n34967), .B(n34963), .Z(n35015) );
  XNOR U35201 ( .A(n34962), .B(n34958), .Z(n35016) );
  XNOR U35202 ( .A(n34957), .B(n34953), .Z(n35017) );
  XNOR U35203 ( .A(n34952), .B(n34948), .Z(n35018) );
  XNOR U35204 ( .A(n34947), .B(n34943), .Z(n35019) );
  XNOR U35205 ( .A(n34942), .B(n34938), .Z(n35020) );
  XOR U35206 ( .A(n35021), .B(n34937), .Z(n34938) );
  AND U35207 ( .A(a[0]), .B(b[15]), .Z(n35021) );
  XOR U35208 ( .A(n35022), .B(n34937), .Z(n34939) );
  XNOR U35209 ( .A(n35023), .B(n35024), .Z(n34937) );
  AND U35210 ( .A(n35025), .B(n35026), .Z(n35023) );
  AND U35211 ( .A(a[1]), .B(b[14]), .Z(n35022) );
  XOR U35212 ( .A(n35027), .B(n34942), .Z(n34944) );
  XOR U35213 ( .A(n35028), .B(n35029), .Z(n34942) );
  AND U35214 ( .A(n35030), .B(n35031), .Z(n35028) );
  AND U35215 ( .A(a[2]), .B(b[13]), .Z(n35027) );
  XOR U35216 ( .A(n35032), .B(n34947), .Z(n34949) );
  XOR U35217 ( .A(n35033), .B(n35034), .Z(n34947) );
  AND U35218 ( .A(n35035), .B(n35036), .Z(n35033) );
  AND U35219 ( .A(a[3]), .B(b[12]), .Z(n35032) );
  XOR U35220 ( .A(n35037), .B(n34952), .Z(n34954) );
  XOR U35221 ( .A(n35038), .B(n35039), .Z(n34952) );
  AND U35222 ( .A(n35040), .B(n35041), .Z(n35038) );
  AND U35223 ( .A(a[4]), .B(b[11]), .Z(n35037) );
  XOR U35224 ( .A(n35042), .B(n34957), .Z(n34959) );
  XOR U35225 ( .A(n35043), .B(n35044), .Z(n34957) );
  AND U35226 ( .A(n35045), .B(n35046), .Z(n35043) );
  AND U35227 ( .A(a[5]), .B(b[10]), .Z(n35042) );
  XOR U35228 ( .A(n35047), .B(n34962), .Z(n34964) );
  XOR U35229 ( .A(n35048), .B(n35049), .Z(n34962) );
  AND U35230 ( .A(n35050), .B(n35051), .Z(n35048) );
  AND U35231 ( .A(a[6]), .B(b[9]), .Z(n35047) );
  XOR U35232 ( .A(n35052), .B(n34967), .Z(n34969) );
  XOR U35233 ( .A(n35053), .B(n35054), .Z(n34967) );
  AND U35234 ( .A(n35055), .B(n35056), .Z(n35053) );
  AND U35235 ( .A(a[7]), .B(b[8]), .Z(n35052) );
  XOR U35236 ( .A(n35057), .B(n34972), .Z(n34974) );
  XOR U35237 ( .A(n35058), .B(n35059), .Z(n34972) );
  AND U35238 ( .A(n35060), .B(n35061), .Z(n35058) );
  AND U35239 ( .A(b[7]), .B(a[8]), .Z(n35057) );
  XOR U35240 ( .A(n35062), .B(n34977), .Z(n34979) );
  XOR U35241 ( .A(n35063), .B(n35064), .Z(n34977) );
  AND U35242 ( .A(n35065), .B(n35066), .Z(n35063) );
  AND U35243 ( .A(b[6]), .B(a[9]), .Z(n35062) );
  XOR U35244 ( .A(n35067), .B(n34982), .Z(n34984) );
  XOR U35245 ( .A(n35068), .B(n35069), .Z(n34982) );
  AND U35246 ( .A(n35070), .B(n35071), .Z(n35068) );
  AND U35247 ( .A(b[5]), .B(a[10]), .Z(n35067) );
  XOR U35248 ( .A(n35072), .B(n34987), .Z(n34989) );
  XOR U35249 ( .A(n35073), .B(n35074), .Z(n34987) );
  AND U35250 ( .A(n35075), .B(n35076), .Z(n35073) );
  AND U35251 ( .A(b[4]), .B(a[11]), .Z(n35072) );
  XNOR U35252 ( .A(n35077), .B(n35078), .Z(n35001) );
  NANDN U35253 ( .A(n35007), .B(n35008), .Z(n35078) );
  XOR U35254 ( .A(n35077), .B(n35079), .Z(n35008) );
  NAND U35255 ( .A(b[1]), .B(a[13]), .Z(n35079) );
  XOR U35256 ( .A(n35080), .B(n35081), .Z(n35007) );
  XOR U35257 ( .A(n35077), .B(n35082), .Z(n35081) );
  NANDN U35258 ( .A(n31877), .B(n31875), .Z(n35077) );
  XNOR U35259 ( .A(n35083), .B(n35084), .Z(n31875) );
  NAND U35260 ( .A(a[13]), .B(b[0]), .Z(n31877) );
  XOR U35261 ( .A(n35085), .B(n34992), .Z(n34994) );
  XNOR U35262 ( .A(n35086), .B(n35087), .Z(n34992) );
  AND U35263 ( .A(n35082), .B(n35080), .Z(n35086) );
  XOR U35264 ( .A(n35087), .B(n35075), .Z(n35088) );
  XNOR U35265 ( .A(n35074), .B(n35070), .Z(n35089) );
  XNOR U35266 ( .A(n35069), .B(n35065), .Z(n35090) );
  XNOR U35267 ( .A(n35064), .B(n35060), .Z(n35091) );
  XNOR U35268 ( .A(n35059), .B(n35055), .Z(n35092) );
  XNOR U35269 ( .A(n35054), .B(n35050), .Z(n35093) );
  XNOR U35270 ( .A(n35049), .B(n35045), .Z(n35094) );
  XNOR U35271 ( .A(n35044), .B(n35040), .Z(n35095) );
  XNOR U35272 ( .A(n35039), .B(n35035), .Z(n35096) );
  XNOR U35273 ( .A(n35034), .B(n35030), .Z(n35097) );
  XNOR U35274 ( .A(n35029), .B(n35025), .Z(n35098) );
  XNOR U35275 ( .A(n35099), .B(n35024), .Z(n35025) );
  AND U35276 ( .A(a[0]), .B(b[14]), .Z(n35099) );
  XNOR U35277 ( .A(n35100), .B(n35024), .Z(n35026) );
  XNOR U35278 ( .A(n35101), .B(n35102), .Z(n35024) );
  AND U35279 ( .A(n35103), .B(n35104), .Z(n35101) );
  AND U35280 ( .A(a[1]), .B(b[13]), .Z(n35100) );
  XOR U35281 ( .A(n35105), .B(n35029), .Z(n35031) );
  XOR U35282 ( .A(n35106), .B(n35107), .Z(n35029) );
  AND U35283 ( .A(n35108), .B(n35109), .Z(n35106) );
  AND U35284 ( .A(a[2]), .B(b[12]), .Z(n35105) );
  XOR U35285 ( .A(n35110), .B(n35034), .Z(n35036) );
  XOR U35286 ( .A(n35111), .B(n35112), .Z(n35034) );
  AND U35287 ( .A(n35113), .B(n35114), .Z(n35111) );
  AND U35288 ( .A(a[3]), .B(b[11]), .Z(n35110) );
  XOR U35289 ( .A(n35115), .B(n35039), .Z(n35041) );
  XOR U35290 ( .A(n35116), .B(n35117), .Z(n35039) );
  AND U35291 ( .A(n35118), .B(n35119), .Z(n35116) );
  AND U35292 ( .A(a[4]), .B(b[10]), .Z(n35115) );
  XOR U35293 ( .A(n35120), .B(n35044), .Z(n35046) );
  XOR U35294 ( .A(n35121), .B(n35122), .Z(n35044) );
  AND U35295 ( .A(n35123), .B(n35124), .Z(n35121) );
  AND U35296 ( .A(a[5]), .B(b[9]), .Z(n35120) );
  XOR U35297 ( .A(n35125), .B(n35049), .Z(n35051) );
  XOR U35298 ( .A(n35126), .B(n35127), .Z(n35049) );
  AND U35299 ( .A(n35128), .B(n35129), .Z(n35126) );
  AND U35300 ( .A(a[6]), .B(b[8]), .Z(n35125) );
  XOR U35301 ( .A(n35130), .B(n35054), .Z(n35056) );
  XOR U35302 ( .A(n35131), .B(n35132), .Z(n35054) );
  AND U35303 ( .A(n35133), .B(n35134), .Z(n35131) );
  AND U35304 ( .A(a[7]), .B(b[7]), .Z(n35130) );
  XOR U35305 ( .A(n35135), .B(n35059), .Z(n35061) );
  XOR U35306 ( .A(n35136), .B(n35137), .Z(n35059) );
  AND U35307 ( .A(n35138), .B(n35139), .Z(n35136) );
  AND U35308 ( .A(b[6]), .B(a[8]), .Z(n35135) );
  XOR U35309 ( .A(n35140), .B(n35064), .Z(n35066) );
  XOR U35310 ( .A(n35141), .B(n35142), .Z(n35064) );
  AND U35311 ( .A(n35143), .B(n35144), .Z(n35141) );
  AND U35312 ( .A(b[5]), .B(a[9]), .Z(n35140) );
  XOR U35313 ( .A(n35145), .B(n35069), .Z(n35071) );
  XOR U35314 ( .A(n35146), .B(n35147), .Z(n35069) );
  AND U35315 ( .A(n35148), .B(n35149), .Z(n35146) );
  AND U35316 ( .A(b[4]), .B(a[10]), .Z(n35145) );
  XOR U35317 ( .A(n35150), .B(n35074), .Z(n35076) );
  XNOR U35318 ( .A(n35151), .B(n35152), .Z(n35074) );
  AND U35319 ( .A(n35153), .B(n35154), .Z(n35151) );
  AND U35320 ( .A(b[3]), .B(a[11]), .Z(n35150) );
  XNOR U35321 ( .A(n35155), .B(n35087), .Z(n35082) );
  XNOR U35322 ( .A(n35156), .B(n35157), .Z(n35087) );
  NANDN U35323 ( .A(n35083), .B(n35084), .Z(n35157) );
  XOR U35324 ( .A(n35156), .B(n35158), .Z(n35084) );
  NAND U35325 ( .A(b[1]), .B(a[12]), .Z(n35158) );
  XOR U35326 ( .A(n35154), .B(n35159), .Z(n35083) );
  XOR U35327 ( .A(n35156), .B(n35153), .Z(n35159) );
  XNOR U35328 ( .A(n35160), .B(n35152), .Z(n35153) );
  AND U35329 ( .A(b[2]), .B(a[11]), .Z(n35160) );
  XOR U35330 ( .A(n35152), .B(n35148), .Z(n35161) );
  XNOR U35331 ( .A(n35147), .B(n35143), .Z(n35162) );
  XNOR U35332 ( .A(n35142), .B(n35138), .Z(n35163) );
  XNOR U35333 ( .A(n35137), .B(n35133), .Z(n35164) );
  XNOR U35334 ( .A(n35132), .B(n35128), .Z(n35165) );
  XNOR U35335 ( .A(n35127), .B(n35123), .Z(n35166) );
  XNOR U35336 ( .A(n35122), .B(n35118), .Z(n35167) );
  XNOR U35337 ( .A(n35117), .B(n35113), .Z(n35168) );
  XNOR U35338 ( .A(n35112), .B(n35108), .Z(n35169) );
  XNOR U35339 ( .A(n35107), .B(n35103), .Z(n35170) );
  XOR U35340 ( .A(n35171), .B(n35102), .Z(n35103) );
  AND U35341 ( .A(a[0]), .B(b[13]), .Z(n35171) );
  XOR U35342 ( .A(n35172), .B(n35102), .Z(n35104) );
  XNOR U35343 ( .A(n35173), .B(n35174), .Z(n35102) );
  AND U35344 ( .A(n35175), .B(n35176), .Z(n35173) );
  AND U35345 ( .A(a[1]), .B(b[12]), .Z(n35172) );
  XOR U35346 ( .A(n35177), .B(n35107), .Z(n35109) );
  XOR U35347 ( .A(n35178), .B(n35179), .Z(n35107) );
  AND U35348 ( .A(n35180), .B(n35181), .Z(n35178) );
  AND U35349 ( .A(a[2]), .B(b[11]), .Z(n35177) );
  XOR U35350 ( .A(n35182), .B(n35112), .Z(n35114) );
  XOR U35351 ( .A(n35183), .B(n35184), .Z(n35112) );
  AND U35352 ( .A(n35185), .B(n35186), .Z(n35183) );
  AND U35353 ( .A(a[3]), .B(b[10]), .Z(n35182) );
  XOR U35354 ( .A(n35187), .B(n35117), .Z(n35119) );
  XOR U35355 ( .A(n35188), .B(n35189), .Z(n35117) );
  AND U35356 ( .A(n35190), .B(n35191), .Z(n35188) );
  AND U35357 ( .A(a[4]), .B(b[9]), .Z(n35187) );
  XOR U35358 ( .A(n35192), .B(n35122), .Z(n35124) );
  XOR U35359 ( .A(n35193), .B(n35194), .Z(n35122) );
  AND U35360 ( .A(n35195), .B(n35196), .Z(n35193) );
  AND U35361 ( .A(a[5]), .B(b[8]), .Z(n35192) );
  XOR U35362 ( .A(n35197), .B(n35127), .Z(n35129) );
  XOR U35363 ( .A(n35198), .B(n35199), .Z(n35127) );
  AND U35364 ( .A(n35200), .B(n35201), .Z(n35198) );
  AND U35365 ( .A(a[6]), .B(b[7]), .Z(n35197) );
  XOR U35366 ( .A(n35202), .B(n35132), .Z(n35134) );
  XOR U35367 ( .A(n35203), .B(n35204), .Z(n35132) );
  AND U35368 ( .A(n35205), .B(n35206), .Z(n35203) );
  AND U35369 ( .A(b[6]), .B(a[7]), .Z(n35202) );
  XOR U35370 ( .A(n35207), .B(n35137), .Z(n35139) );
  XOR U35371 ( .A(n35208), .B(n35209), .Z(n35137) );
  AND U35372 ( .A(n35210), .B(n35211), .Z(n35208) );
  AND U35373 ( .A(b[5]), .B(a[8]), .Z(n35207) );
  XOR U35374 ( .A(n35212), .B(n35142), .Z(n35144) );
  XOR U35375 ( .A(n35213), .B(n35214), .Z(n35142) );
  AND U35376 ( .A(n35215), .B(n35216), .Z(n35213) );
  AND U35377 ( .A(b[4]), .B(a[9]), .Z(n35212) );
  XNOR U35378 ( .A(n35217), .B(n35218), .Z(n35152) );
  NANDN U35379 ( .A(n35219), .B(n35220), .Z(n35218) );
  XOR U35380 ( .A(n35221), .B(n35147), .Z(n35149) );
  XNOR U35381 ( .A(n35222), .B(n35223), .Z(n35147) );
  AND U35382 ( .A(n35224), .B(n35225), .Z(n35222) );
  AND U35383 ( .A(b[3]), .B(a[10]), .Z(n35221) );
  NANDN U35384 ( .A(n31882), .B(n31880), .Z(n35156) );
  XNOR U35385 ( .A(n35219), .B(n35220), .Z(n31880) );
  XOR U35386 ( .A(n35217), .B(n35226), .Z(n35220) );
  NAND U35387 ( .A(b[1]), .B(a[11]), .Z(n35226) );
  XOR U35388 ( .A(n35225), .B(n35227), .Z(n35219) );
  XOR U35389 ( .A(n35217), .B(n35224), .Z(n35227) );
  XNOR U35390 ( .A(n35228), .B(n35223), .Z(n35224) );
  AND U35391 ( .A(b[2]), .B(a[10]), .Z(n35228) );
  NANDN U35392 ( .A(n31887), .B(n31885), .Z(n35217) );
  XNOR U35393 ( .A(n35229), .B(n35230), .Z(n31885) );
  NAND U35394 ( .A(a[11]), .B(b[0]), .Z(n31887) );
  XOR U35395 ( .A(n35223), .B(n35215), .Z(n35231) );
  XNOR U35396 ( .A(n35214), .B(n35210), .Z(n35232) );
  XNOR U35397 ( .A(n35209), .B(n35205), .Z(n35233) );
  XNOR U35398 ( .A(n35204), .B(n35200), .Z(n35234) );
  XNOR U35399 ( .A(n35199), .B(n35195), .Z(n35235) );
  XNOR U35400 ( .A(n35194), .B(n35190), .Z(n35236) );
  XNOR U35401 ( .A(n35189), .B(n35185), .Z(n35237) );
  XNOR U35402 ( .A(n35184), .B(n35180), .Z(n35238) );
  XNOR U35403 ( .A(n35179), .B(n35175), .Z(n35239) );
  XNOR U35404 ( .A(n35240), .B(n35174), .Z(n35175) );
  AND U35405 ( .A(a[0]), .B(b[12]), .Z(n35240) );
  XNOR U35406 ( .A(n35241), .B(n35174), .Z(n35176) );
  XNOR U35407 ( .A(n35242), .B(n35243), .Z(n35174) );
  AND U35408 ( .A(n35244), .B(n35245), .Z(n35242) );
  AND U35409 ( .A(a[1]), .B(b[11]), .Z(n35241) );
  XOR U35410 ( .A(n35246), .B(n35179), .Z(n35181) );
  XOR U35411 ( .A(n35247), .B(n35248), .Z(n35179) );
  AND U35412 ( .A(n35249), .B(n35250), .Z(n35247) );
  AND U35413 ( .A(a[2]), .B(b[10]), .Z(n35246) );
  XOR U35414 ( .A(n35251), .B(n35184), .Z(n35186) );
  XOR U35415 ( .A(n35252), .B(n35253), .Z(n35184) );
  AND U35416 ( .A(n35254), .B(n35255), .Z(n35252) );
  AND U35417 ( .A(a[3]), .B(b[9]), .Z(n35251) );
  XOR U35418 ( .A(n35256), .B(n35189), .Z(n35191) );
  XOR U35419 ( .A(n35257), .B(n35258), .Z(n35189) );
  AND U35420 ( .A(n35259), .B(n35260), .Z(n35257) );
  AND U35421 ( .A(a[4]), .B(b[8]), .Z(n35256) );
  XOR U35422 ( .A(n35261), .B(n35194), .Z(n35196) );
  XOR U35423 ( .A(n35262), .B(n35263), .Z(n35194) );
  AND U35424 ( .A(n35264), .B(n35265), .Z(n35262) );
  AND U35425 ( .A(a[5]), .B(b[7]), .Z(n35261) );
  XOR U35426 ( .A(n35266), .B(n35199), .Z(n35201) );
  XOR U35427 ( .A(n35267), .B(n35268), .Z(n35199) );
  AND U35428 ( .A(n35269), .B(n35270), .Z(n35267) );
  AND U35429 ( .A(a[6]), .B(b[6]), .Z(n35266) );
  XOR U35430 ( .A(n35271), .B(n35204), .Z(n35206) );
  XOR U35431 ( .A(n35272), .B(n35273), .Z(n35204) );
  AND U35432 ( .A(n35274), .B(n35275), .Z(n35272) );
  AND U35433 ( .A(b[5]), .B(a[7]), .Z(n35271) );
  XOR U35434 ( .A(n35276), .B(n35209), .Z(n35211) );
  XOR U35435 ( .A(n35277), .B(n35278), .Z(n35209) );
  AND U35436 ( .A(n35279), .B(n35280), .Z(n35277) );
  AND U35437 ( .A(b[4]), .B(a[8]), .Z(n35276) );
  XNOR U35438 ( .A(n35281), .B(n35282), .Z(n35223) );
  NANDN U35439 ( .A(n35229), .B(n35230), .Z(n35282) );
  XOR U35440 ( .A(n35281), .B(n35283), .Z(n35230) );
  NAND U35441 ( .A(b[1]), .B(a[10]), .Z(n35283) );
  XOR U35442 ( .A(n35284), .B(n35285), .Z(n35229) );
  XOR U35443 ( .A(n35281), .B(n35286), .Z(n35285) );
  NANDN U35444 ( .A(n31892), .B(n31890), .Z(n35281) );
  XNOR U35445 ( .A(n35287), .B(n35288), .Z(n31890) );
  NAND U35446 ( .A(a[10]), .B(b[0]), .Z(n31892) );
  XOR U35447 ( .A(n35289), .B(n35214), .Z(n35216) );
  XNOR U35448 ( .A(n35290), .B(n35291), .Z(n35214) );
  AND U35449 ( .A(n35286), .B(n35284), .Z(n35290) );
  XOR U35450 ( .A(n35291), .B(n35279), .Z(n35292) );
  XNOR U35451 ( .A(n35278), .B(n35274), .Z(n35293) );
  XNOR U35452 ( .A(n35273), .B(n35269), .Z(n35294) );
  XNOR U35453 ( .A(n35268), .B(n35264), .Z(n35295) );
  XNOR U35454 ( .A(n35263), .B(n35259), .Z(n35296) );
  XNOR U35455 ( .A(n35258), .B(n35254), .Z(n35297) );
  XNOR U35456 ( .A(n35253), .B(n35249), .Z(n35298) );
  XNOR U35457 ( .A(n35248), .B(n35244), .Z(n35299) );
  XOR U35458 ( .A(n35300), .B(n35243), .Z(n35244) );
  AND U35459 ( .A(a[0]), .B(b[11]), .Z(n35300) );
  XOR U35460 ( .A(n35301), .B(n35243), .Z(n35245) );
  XNOR U35461 ( .A(n35302), .B(n35303), .Z(n35243) );
  AND U35462 ( .A(n35304), .B(n35305), .Z(n35302) );
  AND U35463 ( .A(a[1]), .B(b[10]), .Z(n35301) );
  XOR U35464 ( .A(n35306), .B(n35248), .Z(n35250) );
  XOR U35465 ( .A(n35307), .B(n35308), .Z(n35248) );
  AND U35466 ( .A(n35309), .B(n35310), .Z(n35307) );
  AND U35467 ( .A(a[2]), .B(b[9]), .Z(n35306) );
  XOR U35468 ( .A(n35311), .B(n35253), .Z(n35255) );
  XOR U35469 ( .A(n35312), .B(n35313), .Z(n35253) );
  AND U35470 ( .A(n35314), .B(n35315), .Z(n35312) );
  AND U35471 ( .A(a[3]), .B(b[8]), .Z(n35311) );
  XOR U35472 ( .A(n35316), .B(n35258), .Z(n35260) );
  XOR U35473 ( .A(n35317), .B(n35318), .Z(n35258) );
  AND U35474 ( .A(n35319), .B(n35320), .Z(n35317) );
  AND U35475 ( .A(a[4]), .B(b[7]), .Z(n35316) );
  XOR U35476 ( .A(n35321), .B(n35263), .Z(n35265) );
  XOR U35477 ( .A(n35322), .B(n35323), .Z(n35263) );
  AND U35478 ( .A(n35324), .B(n35325), .Z(n35322) );
  AND U35479 ( .A(a[5]), .B(b[6]), .Z(n35321) );
  XOR U35480 ( .A(n35326), .B(n35268), .Z(n35270) );
  XOR U35481 ( .A(n35327), .B(n35328), .Z(n35268) );
  AND U35482 ( .A(n35329), .B(n35330), .Z(n35327) );
  AND U35483 ( .A(b[5]), .B(a[6]), .Z(n35326) );
  XOR U35484 ( .A(n35331), .B(n35273), .Z(n35275) );
  XOR U35485 ( .A(n35332), .B(n35333), .Z(n35273) );
  AND U35486 ( .A(n35334), .B(n35335), .Z(n35332) );
  AND U35487 ( .A(b[4]), .B(a[7]), .Z(n35331) );
  XOR U35488 ( .A(n35336), .B(n35278), .Z(n35280) );
  XNOR U35489 ( .A(n35337), .B(n35338), .Z(n35278) );
  AND U35490 ( .A(n35339), .B(n35340), .Z(n35337) );
  AND U35491 ( .A(b[3]), .B(a[8]), .Z(n35336) );
  XNOR U35492 ( .A(n35341), .B(n35291), .Z(n35286) );
  XNOR U35493 ( .A(n35342), .B(n35343), .Z(n35291) );
  NANDN U35494 ( .A(n35287), .B(n35288), .Z(n35343) );
  XOR U35495 ( .A(n35342), .B(n35344), .Z(n35288) );
  NAND U35496 ( .A(b[1]), .B(a[9]), .Z(n35344) );
  XOR U35497 ( .A(n35340), .B(n35345), .Z(n35287) );
  XOR U35498 ( .A(n35342), .B(n35339), .Z(n35345) );
  XNOR U35499 ( .A(n35346), .B(n35338), .Z(n35339) );
  AND U35500 ( .A(b[2]), .B(a[8]), .Z(n35346) );
  XOR U35501 ( .A(n35338), .B(n35334), .Z(n35347) );
  XNOR U35502 ( .A(n35333), .B(n35329), .Z(n35348) );
  XNOR U35503 ( .A(n35328), .B(n35324), .Z(n35349) );
  XNOR U35504 ( .A(n35323), .B(n35319), .Z(n35350) );
  XNOR U35505 ( .A(n35318), .B(n35314), .Z(n35351) );
  XNOR U35506 ( .A(n35313), .B(n35309), .Z(n35352) );
  XNOR U35507 ( .A(n35308), .B(n35304), .Z(n35353) );
  XNOR U35508 ( .A(n35354), .B(n35303), .Z(n35304) );
  AND U35509 ( .A(a[0]), .B(b[10]), .Z(n35354) );
  XNOR U35510 ( .A(n35355), .B(n35303), .Z(n35305) );
  XNOR U35511 ( .A(n35356), .B(n35357), .Z(n35303) );
  AND U35512 ( .A(n35358), .B(n35359), .Z(n35356) );
  AND U35513 ( .A(a[1]), .B(b[9]), .Z(n35355) );
  XOR U35514 ( .A(n35360), .B(n35308), .Z(n35310) );
  XOR U35515 ( .A(n35361), .B(n35362), .Z(n35308) );
  AND U35516 ( .A(n35363), .B(n35364), .Z(n35361) );
  AND U35517 ( .A(a[2]), .B(b[8]), .Z(n35360) );
  XOR U35518 ( .A(n35365), .B(n35313), .Z(n35315) );
  XOR U35519 ( .A(n35366), .B(n35367), .Z(n35313) );
  AND U35520 ( .A(n35368), .B(n35369), .Z(n35366) );
  AND U35521 ( .A(a[3]), .B(b[7]), .Z(n35365) );
  XOR U35522 ( .A(n35370), .B(n35318), .Z(n35320) );
  XOR U35523 ( .A(n35371), .B(n35372), .Z(n35318) );
  AND U35524 ( .A(n35373), .B(n35374), .Z(n35371) );
  AND U35525 ( .A(a[4]), .B(b[6]), .Z(n35370) );
  XOR U35526 ( .A(n35375), .B(n35323), .Z(n35325) );
  XOR U35527 ( .A(n35376), .B(n35377), .Z(n35323) );
  AND U35528 ( .A(n35378), .B(n35379), .Z(n35376) );
  AND U35529 ( .A(a[5]), .B(b[5]), .Z(n35375) );
  XOR U35530 ( .A(n35380), .B(n35328), .Z(n35330) );
  XOR U35531 ( .A(n35381), .B(n35382), .Z(n35328) );
  AND U35532 ( .A(n35383), .B(n35384), .Z(n35381) );
  AND U35533 ( .A(b[4]), .B(a[6]), .Z(n35380) );
  XNOR U35534 ( .A(n35385), .B(n35386), .Z(n35338) );
  NANDN U35535 ( .A(n35387), .B(n35388), .Z(n35386) );
  XOR U35536 ( .A(n35389), .B(n35333), .Z(n35335) );
  XNOR U35537 ( .A(n35390), .B(n35391), .Z(n35333) );
  AND U35538 ( .A(n35392), .B(n35393), .Z(n35390) );
  AND U35539 ( .A(b[3]), .B(a[7]), .Z(n35389) );
  NANDN U35540 ( .A(n31897), .B(n31895), .Z(n35342) );
  XNOR U35541 ( .A(n35387), .B(n35388), .Z(n31895) );
  XOR U35542 ( .A(n35385), .B(n35394), .Z(n35388) );
  NAND U35543 ( .A(b[1]), .B(a[8]), .Z(n35394) );
  XOR U35544 ( .A(n35393), .B(n35395), .Z(n35387) );
  XOR U35545 ( .A(n35385), .B(n35392), .Z(n35395) );
  XNOR U35546 ( .A(n35396), .B(n35391), .Z(n35392) );
  AND U35547 ( .A(b[2]), .B(a[7]), .Z(n35396) );
  NANDN U35548 ( .A(n31902), .B(n31900), .Z(n35385) );
  XNOR U35549 ( .A(n35397), .B(n35398), .Z(n31900) );
  NAND U35550 ( .A(a[8]), .B(b[0]), .Z(n31902) );
  XOR U35551 ( .A(n35391), .B(n35383), .Z(n35399) );
  XNOR U35552 ( .A(n35382), .B(n35378), .Z(n35400) );
  XNOR U35553 ( .A(n35377), .B(n35373), .Z(n35401) );
  XNOR U35554 ( .A(n35372), .B(n35368), .Z(n35402) );
  XNOR U35555 ( .A(n35367), .B(n35363), .Z(n35403) );
  XNOR U35556 ( .A(n35362), .B(n35358), .Z(n35404) );
  XOR U35557 ( .A(n35405), .B(n35357), .Z(n35358) );
  AND U35558 ( .A(a[0]), .B(b[9]), .Z(n35405) );
  XOR U35559 ( .A(n35406), .B(n35357), .Z(n35359) );
  XNOR U35560 ( .A(n35407), .B(n35408), .Z(n35357) );
  AND U35561 ( .A(n35409), .B(n35410), .Z(n35407) );
  AND U35562 ( .A(a[1]), .B(b[8]), .Z(n35406) );
  XOR U35563 ( .A(n35411), .B(n35362), .Z(n35364) );
  XOR U35564 ( .A(n35412), .B(n35413), .Z(n35362) );
  AND U35565 ( .A(n35414), .B(n35415), .Z(n35412) );
  AND U35566 ( .A(a[2]), .B(b[7]), .Z(n35411) );
  XOR U35567 ( .A(n35416), .B(n35367), .Z(n35369) );
  XOR U35568 ( .A(n35417), .B(n35418), .Z(n35367) );
  AND U35569 ( .A(n35419), .B(n35420), .Z(n35417) );
  AND U35570 ( .A(a[3]), .B(b[6]), .Z(n35416) );
  XOR U35571 ( .A(n35421), .B(n35372), .Z(n35374) );
  XOR U35572 ( .A(n35422), .B(n35423), .Z(n35372) );
  AND U35573 ( .A(n35424), .B(n35425), .Z(n35422) );
  AND U35574 ( .A(a[4]), .B(b[5]), .Z(n35421) );
  XOR U35575 ( .A(n35426), .B(n35377), .Z(n35379) );
  XOR U35576 ( .A(n35427), .B(n35428), .Z(n35377) );
  AND U35577 ( .A(n35429), .B(n35430), .Z(n35427) );
  AND U35578 ( .A(b[4]), .B(a[5]), .Z(n35426) );
  XNOR U35579 ( .A(n35431), .B(n35432), .Z(n35391) );
  NANDN U35580 ( .A(n35397), .B(n35398), .Z(n35432) );
  XOR U35581 ( .A(n35431), .B(n35433), .Z(n35398) );
  NAND U35582 ( .A(b[1]), .B(a[7]), .Z(n35433) );
  XOR U35583 ( .A(n35434), .B(n35435), .Z(n35397) );
  XOR U35584 ( .A(n35431), .B(n35436), .Z(n35435) );
  NANDN U35585 ( .A(n31907), .B(n31905), .Z(n35431) );
  XNOR U35586 ( .A(n35437), .B(n35438), .Z(n31905) );
  NAND U35587 ( .A(a[7]), .B(b[0]), .Z(n31907) );
  XOR U35588 ( .A(n35439), .B(n35382), .Z(n35384) );
  XNOR U35589 ( .A(n35440), .B(n35441), .Z(n35382) );
  AND U35590 ( .A(n35436), .B(n35434), .Z(n35440) );
  XOR U35591 ( .A(n35441), .B(n35429), .Z(n35442) );
  XNOR U35592 ( .A(n35428), .B(n35424), .Z(n35443) );
  XNOR U35593 ( .A(n35423), .B(n35419), .Z(n35444) );
  XNOR U35594 ( .A(n35418), .B(n35414), .Z(n35445) );
  XNOR U35595 ( .A(n35413), .B(n35409), .Z(n35446) );
  XNOR U35596 ( .A(n35447), .B(n35408), .Z(n35409) );
  AND U35597 ( .A(a[0]), .B(b[8]), .Z(n35447) );
  XNOR U35598 ( .A(n35448), .B(n35408), .Z(n35410) );
  XNOR U35599 ( .A(n35449), .B(n35450), .Z(n35408) );
  AND U35600 ( .A(n35451), .B(n35452), .Z(n35449) );
  AND U35601 ( .A(a[1]), .B(b[7]), .Z(n35448) );
  XOR U35602 ( .A(n35453), .B(n35413), .Z(n35415) );
  XOR U35603 ( .A(n35454), .B(n35455), .Z(n35413) );
  AND U35604 ( .A(n35456), .B(n35457), .Z(n35454) );
  AND U35605 ( .A(a[2]), .B(b[6]), .Z(n35453) );
  XOR U35606 ( .A(n35458), .B(n35418), .Z(n35420) );
  XOR U35607 ( .A(n35459), .B(n35460), .Z(n35418) );
  AND U35608 ( .A(n35461), .B(n35462), .Z(n35459) );
  AND U35609 ( .A(a[3]), .B(b[5]), .Z(n35458) );
  XOR U35610 ( .A(n35463), .B(n35423), .Z(n35425) );
  XOR U35611 ( .A(n35464), .B(n35465), .Z(n35423) );
  AND U35612 ( .A(n35466), .B(n35467), .Z(n35464) );
  AND U35613 ( .A(a[4]), .B(b[4]), .Z(n35463) );
  XOR U35614 ( .A(n35468), .B(n35428), .Z(n35430) );
  XNOR U35615 ( .A(n35469), .B(n35470), .Z(n35428) );
  AND U35616 ( .A(n35471), .B(n35472), .Z(n35469) );
  AND U35617 ( .A(b[3]), .B(a[5]), .Z(n35468) );
  XNOR U35618 ( .A(n35473), .B(n35441), .Z(n35436) );
  XNOR U35619 ( .A(n35474), .B(n35475), .Z(n35441) );
  NANDN U35620 ( .A(n35437), .B(n35438), .Z(n35475) );
  XOR U35621 ( .A(n35474), .B(n35476), .Z(n35438) );
  NAND U35622 ( .A(b[1]), .B(a[6]), .Z(n35476) );
  XOR U35623 ( .A(n35472), .B(n35477), .Z(n35437) );
  XOR U35624 ( .A(n35474), .B(n35471), .Z(n35477) );
  XNOR U35625 ( .A(n35478), .B(n35470), .Z(n35471) );
  AND U35626 ( .A(b[2]), .B(a[5]), .Z(n35478) );
  XOR U35627 ( .A(n35470), .B(n35466), .Z(n35479) );
  XNOR U35628 ( .A(n35465), .B(n35461), .Z(n35480) );
  XNOR U35629 ( .A(n35460), .B(n35456), .Z(n35481) );
  XNOR U35630 ( .A(n35455), .B(n35451), .Z(n35482) );
  XOR U35631 ( .A(n35483), .B(n35450), .Z(n35451) );
  AND U35632 ( .A(a[0]), .B(b[7]), .Z(n35483) );
  XOR U35633 ( .A(n35484), .B(n35450), .Z(n35452) );
  XNOR U35634 ( .A(n35485), .B(n35486), .Z(n35450) );
  AND U35635 ( .A(n35487), .B(n35488), .Z(n35485) );
  AND U35636 ( .A(a[1]), .B(b[6]), .Z(n35484) );
  XOR U35637 ( .A(n35489), .B(n35455), .Z(n35457) );
  XOR U35638 ( .A(n35490), .B(n35491), .Z(n35455) );
  AND U35639 ( .A(n35492), .B(n35493), .Z(n35490) );
  AND U35640 ( .A(a[2]), .B(b[5]), .Z(n35489) );
  XOR U35641 ( .A(n35494), .B(n35460), .Z(n35462) );
  XOR U35642 ( .A(n35495), .B(n35496), .Z(n35460) );
  AND U35643 ( .A(n35497), .B(n35498), .Z(n35495) );
  AND U35644 ( .A(a[3]), .B(b[4]), .Z(n35494) );
  XNOR U35645 ( .A(n35499), .B(n35500), .Z(n35470) );
  NANDN U35646 ( .A(n35501), .B(n35502), .Z(n35500) );
  XOR U35647 ( .A(n35503), .B(n35465), .Z(n35467) );
  XNOR U35648 ( .A(n35504), .B(n35505), .Z(n35465) );
  AND U35649 ( .A(n35506), .B(n35507), .Z(n35504) );
  AND U35650 ( .A(b[3]), .B(a[4]), .Z(n35503) );
  NANDN U35651 ( .A(n31912), .B(n31910), .Z(n35474) );
  XNOR U35652 ( .A(n35501), .B(n35502), .Z(n31910) );
  XOR U35653 ( .A(n35499), .B(n35508), .Z(n35502) );
  NAND U35654 ( .A(b[1]), .B(a[5]), .Z(n35508) );
  XOR U35655 ( .A(n35507), .B(n35509), .Z(n35501) );
  XOR U35656 ( .A(n35499), .B(n35506), .Z(n35509) );
  XNOR U35657 ( .A(n35510), .B(n35505), .Z(n35506) );
  AND U35658 ( .A(b[2]), .B(a[4]), .Z(n35510) );
  NANDN U35659 ( .A(n31917), .B(n31915), .Z(n35499) );
  XNOR U35660 ( .A(n35511), .B(n35512), .Z(n31915) );
  NAND U35661 ( .A(a[5]), .B(b[0]), .Z(n31917) );
  XOR U35662 ( .A(n35505), .B(n35497), .Z(n35513) );
  XNOR U35663 ( .A(n35496), .B(n35492), .Z(n35514) );
  XNOR U35664 ( .A(n35491), .B(n35487), .Z(n35515) );
  XNOR U35665 ( .A(n35516), .B(n35486), .Z(n35487) );
  AND U35666 ( .A(a[0]), .B(b[6]), .Z(n35516) );
  XNOR U35667 ( .A(n35517), .B(n35486), .Z(n35488) );
  XNOR U35668 ( .A(n35518), .B(n35519), .Z(n35486) );
  AND U35669 ( .A(n35520), .B(n35521), .Z(n35518) );
  AND U35670 ( .A(a[1]), .B(b[5]), .Z(n35517) );
  XOR U35671 ( .A(n35522), .B(n35491), .Z(n35493) );
  XOR U35672 ( .A(n35523), .B(n35524), .Z(n35491) );
  AND U35673 ( .A(n35525), .B(n35526), .Z(n35523) );
  AND U35674 ( .A(a[2]), .B(b[4]), .Z(n35522) );
  XNOR U35675 ( .A(n35527), .B(n35528), .Z(n35505) );
  NANDN U35676 ( .A(n35511), .B(n35512), .Z(n35528) );
  XOR U35677 ( .A(n35527), .B(n35529), .Z(n35512) );
  NAND U35678 ( .A(b[1]), .B(a[4]), .Z(n35529) );
  XOR U35679 ( .A(n35530), .B(n35531), .Z(n35511) );
  XOR U35680 ( .A(n35527), .B(n35532), .Z(n35531) );
  NANDN U35681 ( .A(n31922), .B(n31920), .Z(n35527) );
  XNOR U35682 ( .A(n35533), .B(n35534), .Z(n31920) );
  NAND U35683 ( .A(a[4]), .B(b[0]), .Z(n31922) );
  XOR U35684 ( .A(n35535), .B(n35496), .Z(n35498) );
  XNOR U35685 ( .A(n35536), .B(n35537), .Z(n35496) );
  AND U35686 ( .A(n35532), .B(n35530), .Z(n35536) );
  XOR U35687 ( .A(n35537), .B(n35525), .Z(n35538) );
  XNOR U35688 ( .A(n35524), .B(n35520), .Z(n35539) );
  XOR U35689 ( .A(n35540), .B(n35519), .Z(n35520) );
  AND U35690 ( .A(a[0]), .B(b[5]), .Z(n35540) );
  XOR U35691 ( .A(n35541), .B(n35519), .Z(n35521) );
  XNOR U35692 ( .A(n35542), .B(n35543), .Z(n35519) );
  AND U35693 ( .A(n35544), .B(n35545), .Z(n35542) );
  AND U35694 ( .A(a[1]), .B(b[4]), .Z(n35541) );
  XOR U35695 ( .A(n35546), .B(n35524), .Z(n35526) );
  XNOR U35696 ( .A(n35547), .B(n35548), .Z(n35524) );
  AND U35697 ( .A(n35549), .B(n35550), .Z(n35547) );
  AND U35698 ( .A(a[2]), .B(b[3]), .Z(n35546) );
  XNOR U35699 ( .A(n35551), .B(n35537), .Z(n35532) );
  XNOR U35700 ( .A(n35552), .B(n35553), .Z(n35537) );
  NANDN U35701 ( .A(n35533), .B(n35534), .Z(n35553) );
  XOR U35702 ( .A(n35552), .B(n35554), .Z(n35534) );
  NAND U35703 ( .A(b[1]), .B(a[3]), .Z(n35554) );
  XOR U35704 ( .A(n35550), .B(n35555), .Z(n35533) );
  XOR U35705 ( .A(n35552), .B(n35549), .Z(n35555) );
  XNOR U35706 ( .A(n35556), .B(n35548), .Z(n35549) );
  AND U35707 ( .A(a[2]), .B(b[2]), .Z(n35556) );
  XOR U35708 ( .A(n35548), .B(n35544), .Z(n35557) );
  XNOR U35709 ( .A(n35558), .B(n35543), .Z(n35544) );
  AND U35710 ( .A(a[0]), .B(b[4]), .Z(n35558) );
  XNOR U35711 ( .A(n35559), .B(n35560), .Z(n35548) );
  NANDN U35712 ( .A(n35561), .B(n35562), .Z(n35560) );
  XNOR U35713 ( .A(n35563), .B(n35543), .Z(n35545) );
  XNOR U35714 ( .A(n35564), .B(n35565), .Z(n35543) );
  AND U35715 ( .A(n35566), .B(n35567), .Z(n35564) );
  AND U35716 ( .A(a[1]), .B(b[3]), .Z(n35563) );
  NANDN U35717 ( .A(n31927), .B(n31925), .Z(n35552) );
  XNOR U35718 ( .A(n35561), .B(n35562), .Z(n31925) );
  XOR U35719 ( .A(n35559), .B(n35568), .Z(n35562) );
  NAND U35720 ( .A(b[1]), .B(a[2]), .Z(n35568) );
  XOR U35721 ( .A(n35567), .B(n35569), .Z(n35561) );
  XOR U35722 ( .A(n35559), .B(n35566), .Z(n35569) );
  XOR U35723 ( .A(n35570), .B(n35565), .Z(n35566) );
  AND U35724 ( .A(a[1]), .B(b[2]), .Z(n35570) );
  NANDN U35725 ( .A(n31932), .B(n31930), .Z(n35559) );
  XNOR U35726 ( .A(n35571), .B(n35572), .Z(n31930) );
  NAND U35727 ( .A(a[2]), .B(b[0]), .Z(n31932) );
  XOR U35728 ( .A(n35573), .B(n35565), .Z(n35567) );
  XOR U35729 ( .A(n35574), .B(n35575), .Z(n35565) );
  NANDN U35730 ( .A(n35571), .B(n35572), .Z(n35575) );
  XOR U35731 ( .A(n35574), .B(n35576), .Z(n35572) );
  NAND U35732 ( .A(a[1]), .B(b[1]), .Z(n35576) );
  XNOR U35733 ( .A(n35574), .B(n35577), .Z(n35571) );
  NAND U35734 ( .A(a[0]), .B(b[2]), .Z(n35577) );
  OR U35735 ( .A(n31937), .B(n31936), .Z(n35574) );
  NAND U35736 ( .A(a[1]), .B(b[0]), .Z(n31936) );
  NAND U35737 ( .A(a[0]), .B(b[1]), .Z(n31937) );
  AND U35738 ( .A(a[0]), .B(b[3]), .Z(n35573) );
  NAND U35739 ( .A(a[3]), .B(b[0]), .Z(n31927) );
  AND U35740 ( .A(b[2]), .B(a[3]), .Z(n35551) );
  AND U35741 ( .A(a[3]), .B(b[3]), .Z(n35535) );
  NAND U35742 ( .A(a[6]), .B(b[0]), .Z(n31912) );
  AND U35743 ( .A(b[2]), .B(a[6]), .Z(n35473) );
  AND U35744 ( .A(b[3]), .B(a[6]), .Z(n35439) );
  NAND U35745 ( .A(a[9]), .B(b[0]), .Z(n31897) );
  AND U35746 ( .A(b[2]), .B(a[9]), .Z(n35341) );
  AND U35747 ( .A(b[3]), .B(a[9]), .Z(n35289) );
  NAND U35748 ( .A(a[12]), .B(b[0]), .Z(n31882) );
  AND U35749 ( .A(b[2]), .B(a[12]), .Z(n35155) );
  AND U35750 ( .A(b[3]), .B(a[12]), .Z(n35085) );
  NAND U35751 ( .A(a[15]), .B(b[0]), .Z(n31867) );
  AND U35752 ( .A(b[2]), .B(a[15]), .Z(n34915) );
  AND U35753 ( .A(b[3]), .B(a[15]), .Z(n34827) );
  NAND U35754 ( .A(a[18]), .B(b[0]), .Z(n31852) );
  AND U35755 ( .A(b[2]), .B(a[18]), .Z(n34621) );
  AND U35756 ( .A(b[3]), .B(a[18]), .Z(n34515) );
  NAND U35757 ( .A(a[21]), .B(b[0]), .Z(n31837) );
  AND U35758 ( .A(b[2]), .B(a[21]), .Z(n34273) );
  AND U35759 ( .A(b[3]), .B(a[21]), .Z(n34149) );
  NAND U35760 ( .A(a[24]), .B(b[0]), .Z(n31822) );
  AND U35761 ( .A(b[2]), .B(a[24]), .Z(n33871) );
  AND U35762 ( .A(b[3]), .B(a[24]), .Z(n33729) );
  NAND U35763 ( .A(a[27]), .B(b[0]), .Z(n31807) );
  AND U35764 ( .A(b[2]), .B(a[27]), .Z(n33415) );
  AND U35765 ( .A(b[3]), .B(a[27]), .Z(n33255) );
  NAND U35766 ( .A(a[30]), .B(b[0]), .Z(n31792) );
  AND U35767 ( .A(b[2]), .B(a[30]), .Z(n32905) );
  AND U35768 ( .A(b[3]), .B(a[30]), .Z(n32727) );
  NAND U35769 ( .A(a[33]), .B(b[0]), .Z(n31777) );
  AND U35770 ( .A(b[2]), .B(a[33]), .Z(n32341) );
  AND U35771 ( .A(b[3]), .B(a[33]), .Z(n32145) );
endmodule

