
module mult_N8_CC2 ( clk, rst, a, b, c );
  input [7:0] a;
  input [3:0] b;
  output [15:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197;
  wire   [15:0] sreg;

  DFF \sreg_reg[11]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(sreg[11]) );
  DFF \sreg_reg[10]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(sreg[10]) );
  DFF \sreg_reg[9]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(sreg[9]) );
  DFF \sreg_reg[8]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(sreg[8]) );
  DFF \sreg_reg[7]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(sreg[7]) );
  DFF \sreg_reg[6]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(sreg[6]) );
  DFF \sreg_reg[5]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(sreg[5]) );
  DFF \sreg_reg[4]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(sreg[4]) );
  DFF \sreg_reg[3]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[0]) );
  AND U7 ( .A(n74), .B(n75), .Z(n98) );
  XOR U8 ( .A(n103), .B(n104), .Z(n1) );
  NANDN U9 ( .A(n105), .B(n1), .Z(n2) );
  NAND U10 ( .A(n103), .B(n104), .Z(n3) );
  AND U11 ( .A(n2), .B(n3), .Z(n128) );
  NAND U12 ( .A(n120), .B(n121), .Z(n4) );
  XOR U13 ( .A(n120), .B(n121), .Z(n5) );
  NANDN U14 ( .A(n119), .B(n5), .Z(n6) );
  NAND U15 ( .A(n4), .B(n6), .Z(n147) );
  XOR U16 ( .A(n134), .B(n135), .Z(n7) );
  NANDN U17 ( .A(n136), .B(n7), .Z(n8) );
  NAND U18 ( .A(n134), .B(n135), .Z(n9) );
  AND U19 ( .A(n8), .B(n9), .Z(n156) );
  XOR U20 ( .A(n164), .B(n165), .Z(n10) );
  NANDN U21 ( .A(n166), .B(n10), .Z(n11) );
  NAND U22 ( .A(n164), .B(n165), .Z(n12) );
  AND U23 ( .A(n11), .B(n12), .Z(n180) );
  NAND U24 ( .A(n80), .B(n81), .Z(n13) );
  XOR U25 ( .A(n80), .B(n81), .Z(n14) );
  NANDN U26 ( .A(n79), .B(n14), .Z(n15) );
  NAND U27 ( .A(n13), .B(n15), .Z(n96) );
  NAND U28 ( .A(n123), .B(n125), .Z(n16) );
  XOR U29 ( .A(n123), .B(n125), .Z(n17) );
  NAND U30 ( .A(n17), .B(n124), .Z(n18) );
  NAND U31 ( .A(n16), .B(n18), .Z(n142) );
  XOR U32 ( .A(sreg[8]), .B(n115), .Z(n19) );
  NANDN U33 ( .A(n116), .B(n19), .Z(n20) );
  NAND U34 ( .A(sreg[8]), .B(n115), .Z(n21) );
  AND U35 ( .A(n20), .B(n21), .Z(n131) );
  AND U36 ( .A(n90), .B(n91), .Z(n105) );
  NANDN U37 ( .A(n97), .B(n120), .Z(n22) );
  ANDN U38 ( .B(n22), .A(n98), .Z(n108) );
  NAND U39 ( .A(n172), .B(n173), .Z(n23) );
  XOR U40 ( .A(n172), .B(n173), .Z(n24) );
  NANDN U41 ( .A(n171), .B(n24), .Z(n25) );
  NAND U42 ( .A(n23), .B(n25), .Z(n184) );
  NAND U43 ( .A(n131), .B(n130), .Z(n26) );
  XOR U44 ( .A(n131), .B(n130), .Z(n27) );
  NANDN U45 ( .A(sreg[9]), .B(n27), .Z(n28) );
  NAND U46 ( .A(n26), .B(n28), .Z(n150) );
  NAND U47 ( .A(n109), .B(n110), .Z(n29) );
  XOR U48 ( .A(n109), .B(n110), .Z(n30) );
  NANDN U49 ( .A(n108), .B(n30), .Z(n31) );
  NAND U50 ( .A(n29), .B(n31), .Z(n125) );
  NAND U51 ( .A(n127), .B(n128), .Z(n32) );
  XOR U52 ( .A(n127), .B(n128), .Z(n33) );
  NANDN U53 ( .A(n126), .B(n33), .Z(n34) );
  NAND U54 ( .A(n32), .B(n34), .Z(n140) );
  NAND U55 ( .A(n155), .B(n156), .Z(n35) );
  XOR U56 ( .A(n155), .B(n156), .Z(n36) );
  NANDN U57 ( .A(n154), .B(n36), .Z(n37) );
  NAND U58 ( .A(n35), .B(n37), .Z(n172) );
  XOR U59 ( .A(n180), .B(n179), .Z(n38) );
  NANDN U60 ( .A(n178), .B(n38), .Z(n39) );
  NAND U61 ( .A(n180), .B(n179), .Z(n40) );
  AND U62 ( .A(n39), .B(n40), .Z(n182) );
  XOR U63 ( .A(sreg[7]), .B(n100), .Z(n41) );
  NANDN U64 ( .A(n101), .B(n41), .Z(n42) );
  NAND U65 ( .A(sreg[7]), .B(n100), .Z(n43) );
  AND U66 ( .A(n42), .B(n43), .Z(n116) );
  NAND U67 ( .A(n153), .B(n152), .Z(n44) );
  XOR U68 ( .A(n153), .B(n152), .Z(n45) );
  NANDN U69 ( .A(sreg[11]), .B(n45), .Z(n46) );
  NAND U70 ( .A(n44), .B(n46), .Z(n169) );
  NAND U71 ( .A(n95), .B(n96), .Z(n47) );
  XOR U72 ( .A(n95), .B(n96), .Z(n48) );
  NANDN U73 ( .A(n94), .B(n48), .Z(n49) );
  NAND U74 ( .A(n47), .B(n49), .Z(n109) );
  NAND U75 ( .A(n112), .B(n113), .Z(n50) );
  XOR U76 ( .A(n112), .B(n113), .Z(n51) );
  NANDN U77 ( .A(n111), .B(n51), .Z(n52) );
  NAND U78 ( .A(n50), .B(n52), .Z(n124) );
  NAND U79 ( .A(n146), .B(n147), .Z(n53) );
  XOR U80 ( .A(n146), .B(n147), .Z(n54) );
  NANDN U81 ( .A(n145), .B(n54), .Z(n55) );
  NAND U82 ( .A(n53), .B(n55), .Z(n159) );
  NAND U83 ( .A(n150), .B(n149), .Z(n56) );
  XOR U84 ( .A(n150), .B(n149), .Z(n57) );
  NANDN U85 ( .A(sreg[10]), .B(n57), .Z(n58) );
  NAND U86 ( .A(n56), .B(n58), .Z(n153) );
  NANDN U87 ( .A(n182), .B(n183), .Z(n59) );
  XNOR U88 ( .A(n182), .B(n183), .Z(n60) );
  NAND U89 ( .A(n184), .B(n60), .Z(n61) );
  AND U90 ( .A(n59), .B(n61), .Z(n62) );
  XNOR U91 ( .A(n193), .B(n62), .Z(n190) );
  AND U92 ( .A(a[0]), .B(b[0]), .Z(n63) );
  XOR U93 ( .A(n63), .B(sreg[4]), .Z(c[4]) );
  NAND U94 ( .A(b[1]), .B(a[0]), .Z(n97) );
  AND U95 ( .A(b[0]), .B(a[1]), .Z(n65) );
  XOR U96 ( .A(n97), .B(n65), .Z(n69) );
  NAND U97 ( .A(n63), .B(sreg[4]), .Z(n68) );
  IV U98 ( .A(n68), .Z(n67) );
  XOR U99 ( .A(sreg[5]), .B(n67), .Z(n64) );
  XNOR U100 ( .A(n69), .B(n64), .Z(c[5]) );
  NAND U101 ( .A(a[0]), .B(b[2]), .Z(n79) );
  ANDN U102 ( .B(n65), .A(n97), .Z(n81) );
  AND U103 ( .A(b[0]), .B(a[2]), .Z(n75) );
  AND U104 ( .A(b[1]), .B(a[1]), .Z(n74) );
  XOR U105 ( .A(n75), .B(n74), .Z(n80) );
  XNOR U106 ( .A(n81), .B(n80), .Z(n66) );
  XOR U107 ( .A(n79), .B(n66), .Z(n85) );
  IV U108 ( .A(n85), .Z(n83) );
  OR U109 ( .A(sreg[5]), .B(n67), .Z(n72) );
  ANDN U110 ( .B(sreg[5]), .A(n68), .Z(n70) );
  NANDN U111 ( .A(n70), .B(n69), .Z(n71) );
  AND U112 ( .A(n72), .B(n71), .Z(n84) );
  XOR U113 ( .A(n83), .B(n84), .Z(n73) );
  XNOR U114 ( .A(sreg[6]), .B(n73), .Z(c[6]) );
  AND U115 ( .A(a[1]), .B(b[2]), .Z(n91) );
  AND U116 ( .A(b[0]), .B(a[3]), .Z(n90) );
  XOR U117 ( .A(n91), .B(n90), .Z(n95) );
  AND U118 ( .A(a[2]), .B(b[1]), .Z(n77) );
  AND U119 ( .A(a[0]), .B(b[3]), .Z(n76) );
  XNOR U120 ( .A(n77), .B(n76), .Z(n78) );
  XOR U121 ( .A(n98), .B(n78), .Z(n94) );
  XNOR U122 ( .A(n94), .B(n96), .Z(n82) );
  XOR U123 ( .A(n95), .B(n82), .Z(n100) );
  NANDN U124 ( .A(n83), .B(n84), .Z(n88) );
  NOR U125 ( .A(n85), .B(n84), .Z(n86) );
  NANDN U126 ( .A(n86), .B(sreg[6]), .Z(n87) );
  AND U127 ( .A(n88), .B(n87), .Z(n101) );
  XNOR U128 ( .A(n101), .B(sreg[7]), .Z(n89) );
  XOR U129 ( .A(n100), .B(n89), .Z(c[7]) );
  NAND U130 ( .A(a[2]), .B(b[2]), .Z(n104) );
  NAND U131 ( .A(b[3]), .B(a[1]), .Z(n103) );
  XOR U132 ( .A(n105), .B(n103), .Z(n92) );
  XOR U133 ( .A(n104), .B(n92), .Z(n112) );
  AND U134 ( .A(b[1]), .B(a[3]), .Z(n113) );
  NAND U135 ( .A(b[0]), .B(a[4]), .Z(n111) );
  XOR U136 ( .A(n113), .B(n111), .Z(n93) );
  XNOR U137 ( .A(n112), .B(n93), .Z(n110) );
  AND U138 ( .A(b[3]), .B(a[2]), .Z(n120) );
  XNOR U139 ( .A(n109), .B(n108), .Z(n99) );
  XOR U140 ( .A(n110), .B(n99), .Z(n115) );
  XNOR U141 ( .A(n116), .B(sreg[8]), .Z(n102) );
  XOR U142 ( .A(n115), .B(n102), .Z(c[8]) );
  NAND U143 ( .A(b[0]), .B(a[5]), .Z(n126) );
  NAND U144 ( .A(b[2]), .B(a[3]), .Z(n119) );
  AND U145 ( .A(b[1]), .B(a[4]), .Z(n121) );
  XNOR U146 ( .A(n120), .B(n121), .Z(n106) );
  XOR U147 ( .A(n119), .B(n106), .Z(n127) );
  XNOR U148 ( .A(n128), .B(n127), .Z(n107) );
  XOR U149 ( .A(n126), .B(n107), .Z(n123) );
  XNOR U150 ( .A(n125), .B(n124), .Z(n114) );
  XOR U151 ( .A(n123), .B(n114), .Z(n130) );
  XNOR U152 ( .A(n131), .B(sreg[9]), .Z(n117) );
  XNOR U153 ( .A(n130), .B(n117), .Z(c[9]) );
  NAND U154 ( .A(b[2]), .B(a[4]), .Z(n135) );
  AND U155 ( .A(b[1]), .B(a[5]), .Z(n136) );
  NAND U156 ( .A(b[3]), .B(a[3]), .Z(n134) );
  XOR U157 ( .A(n136), .B(n134), .Z(n118) );
  XOR U158 ( .A(n135), .B(n118), .Z(n146) );
  NAND U159 ( .A(b[0]), .B(a[6]), .Z(n145) );
  XOR U160 ( .A(n147), .B(n145), .Z(n122) );
  XOR U161 ( .A(n146), .B(n122), .Z(n139) );
  IV U162 ( .A(n139), .Z(n138) );
  XNOR U163 ( .A(n142), .B(n140), .Z(n129) );
  XOR U164 ( .A(n138), .B(n129), .Z(n149) );
  XNOR U165 ( .A(n150), .B(sreg[10]), .Z(n132) );
  XNOR U166 ( .A(n149), .B(n132), .Z(c[10]) );
  NAND U167 ( .A(b[2]), .B(a[5]), .Z(n165) );
  AND U168 ( .A(b[1]), .B(a[6]), .Z(n166) );
  NAND U169 ( .A(b[3]), .B(a[4]), .Z(n164) );
  XOR U170 ( .A(n166), .B(n164), .Z(n133) );
  XOR U171 ( .A(n165), .B(n133), .Z(n155) );
  NAND U172 ( .A(a[7]), .B(b[0]), .Z(n154) );
  XOR U173 ( .A(n156), .B(n154), .Z(n137) );
  XOR U174 ( .A(n155), .B(n137), .Z(n158) );
  IV U175 ( .A(n158), .Z(n157) );
  OR U176 ( .A(n140), .B(n138), .Z(n144) );
  ANDN U177 ( .B(n140), .A(n139), .Z(n141) );
  OR U178 ( .A(n142), .B(n141), .Z(n143) );
  AND U179 ( .A(n144), .B(n143), .Z(n161) );
  XNOR U180 ( .A(n161), .B(n159), .Z(n148) );
  XOR U181 ( .A(n157), .B(n148), .Z(n152) );
  XNOR U182 ( .A(n153), .B(sreg[11]), .Z(n151) );
  XNOR U183 ( .A(n152), .B(n151), .Z(c[11]) );
  OR U184 ( .A(n159), .B(n157), .Z(n163) );
  ANDN U185 ( .B(n159), .A(n158), .Z(n160) );
  OR U186 ( .A(n161), .B(n160), .Z(n162) );
  AND U187 ( .A(n163), .B(n162), .Z(n173) );
  AND U188 ( .A(b[3]), .B(a[5]), .Z(n179) );
  AND U189 ( .A(b[2]), .B(a[6]), .Z(n191) );
  AND U190 ( .A(a[7]), .B(b[1]), .Z(n185) );
  XNOR U191 ( .A(n191), .B(n185), .Z(n178) );
  XOR U192 ( .A(n179), .B(n178), .Z(n167) );
  XOR U193 ( .A(n180), .B(n167), .Z(n171) );
  XOR U194 ( .A(n173), .B(n171), .Z(n168) );
  XNOR U195 ( .A(n172), .B(n168), .Z(n170) );
  XNOR U196 ( .A(n169), .B(n170), .Z(c[12]) );
  ANDN U197 ( .B(n170), .A(n169), .Z(n189) );
  AND U198 ( .A(n191), .B(n185), .Z(n177) );
  AND U199 ( .A(b[2]), .B(a[7]), .Z(n175) );
  NAND U200 ( .A(a[6]), .B(b[3]), .Z(n174) );
  XNOR U201 ( .A(n175), .B(n174), .Z(n176) );
  XOR U202 ( .A(n177), .B(n176), .Z(n183) );
  XOR U203 ( .A(n183), .B(n182), .Z(n181) );
  XNOR U204 ( .A(n184), .B(n181), .Z(n188) );
  XOR U205 ( .A(n189), .B(n188), .Z(c[13]) );
  AND U206 ( .A(b[3]), .B(a[7]), .Z(n193) );
  OR U207 ( .A(n193), .B(n185), .Z(n186) );
  AND U208 ( .A(n191), .B(n186), .Z(n187) );
  XNOR U209 ( .A(n190), .B(n187), .Z(n195) );
  AND U210 ( .A(n189), .B(n188), .Z(n194) );
  XNOR U211 ( .A(n195), .B(n194), .Z(c[14]) );
  NANDN U212 ( .A(n191), .B(n190), .Z(n192) );
  AND U213 ( .A(n193), .B(n192), .Z(n197) );
  NANDN U214 ( .A(n195), .B(n194), .Z(n196) );
  NANDN U215 ( .A(n197), .B(n196), .Z(c[15]) );
endmodule

