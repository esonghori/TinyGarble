
module sum_N1024_CC1 ( clk, rst, a, b, c );
  input [1023:0] a;
  input [1023:0] b;
  output [1023:0] c;
  input clk, rst;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091;

  XOR U2 ( .A(a[0]), .B(b[0]), .Z(c[0]) );
  XOR U3 ( .A(a[1000]), .B(b[1000]), .Z(n2000) );
  NAND U4 ( .A(b[999]), .B(a[999]), .Z(n1999) );
  XNOR U5 ( .A(b[999]), .B(a[999]), .Z(n4087) );
  NAND U6 ( .A(b[998]), .B(a[998]), .Z(n1997) );
  NAND U7 ( .A(b[997]), .B(a[997]), .Z(n1995) );
  NAND U8 ( .A(b[996]), .B(a[996]), .Z(n1993) );
  NAND U9 ( .A(b[995]), .B(a[995]), .Z(n1991) );
  NAND U10 ( .A(b[994]), .B(a[994]), .Z(n1989) );
  NAND U11 ( .A(b[993]), .B(a[993]), .Z(n1987) );
  NAND U12 ( .A(b[992]), .B(a[992]), .Z(n1985) );
  NAND U13 ( .A(b[991]), .B(a[991]), .Z(n1983) );
  NAND U14 ( .A(b[990]), .B(a[990]), .Z(n1981) );
  NAND U15 ( .A(b[989]), .B(a[989]), .Z(n1979) );
  NAND U16 ( .A(b[988]), .B(a[988]), .Z(n1977) );
  NAND U17 ( .A(b[987]), .B(a[987]), .Z(n1975) );
  NAND U18 ( .A(b[986]), .B(a[986]), .Z(n1973) );
  NAND U19 ( .A(b[985]), .B(a[985]), .Z(n1971) );
  NAND U20 ( .A(b[984]), .B(a[984]), .Z(n1969) );
  NAND U21 ( .A(b[983]), .B(a[983]), .Z(n1967) );
  NAND U22 ( .A(b[982]), .B(a[982]), .Z(n1965) );
  NAND U23 ( .A(b[981]), .B(a[981]), .Z(n1963) );
  NAND U24 ( .A(b[980]), .B(a[980]), .Z(n1961) );
  NAND U25 ( .A(b[979]), .B(a[979]), .Z(n1959) );
  NAND U26 ( .A(b[978]), .B(a[978]), .Z(n1957) );
  NAND U27 ( .A(b[977]), .B(a[977]), .Z(n1955) );
  NAND U28 ( .A(b[976]), .B(a[976]), .Z(n1953) );
  NAND U29 ( .A(b[975]), .B(a[975]), .Z(n1951) );
  NAND U30 ( .A(b[974]), .B(a[974]), .Z(n1949) );
  NAND U31 ( .A(b[973]), .B(a[973]), .Z(n1947) );
  NAND U32 ( .A(b[972]), .B(a[972]), .Z(n1945) );
  NAND U33 ( .A(b[971]), .B(a[971]), .Z(n1943) );
  NAND U34 ( .A(b[970]), .B(a[970]), .Z(n1941) );
  NAND U35 ( .A(b[969]), .B(a[969]), .Z(n1939) );
  NAND U36 ( .A(b[968]), .B(a[968]), .Z(n1937) );
  NAND U37 ( .A(b[967]), .B(a[967]), .Z(n1935) );
  NAND U38 ( .A(b[966]), .B(a[966]), .Z(n1933) );
  NAND U39 ( .A(b[965]), .B(a[965]), .Z(n1931) );
  NAND U40 ( .A(b[964]), .B(a[964]), .Z(n1929) );
  NAND U41 ( .A(b[963]), .B(a[963]), .Z(n1927) );
  NAND U42 ( .A(b[962]), .B(a[962]), .Z(n1925) );
  NAND U43 ( .A(b[961]), .B(a[961]), .Z(n1923) );
  NAND U44 ( .A(b[960]), .B(a[960]), .Z(n1921) );
  NAND U45 ( .A(b[959]), .B(a[959]), .Z(n1919) );
  NAND U46 ( .A(b[958]), .B(a[958]), .Z(n1917) );
  NAND U47 ( .A(b[957]), .B(a[957]), .Z(n1915) );
  NAND U48 ( .A(b[956]), .B(a[956]), .Z(n1913) );
  NAND U49 ( .A(b[955]), .B(a[955]), .Z(n1911) );
  NAND U50 ( .A(b[954]), .B(a[954]), .Z(n1909) );
  NAND U51 ( .A(b[953]), .B(a[953]), .Z(n1907) );
  NAND U52 ( .A(b[952]), .B(a[952]), .Z(n1905) );
  NAND U53 ( .A(b[951]), .B(a[951]), .Z(n1903) );
  NAND U54 ( .A(b[950]), .B(a[950]), .Z(n1901) );
  NAND U55 ( .A(b[949]), .B(a[949]), .Z(n1899) );
  NAND U56 ( .A(b[948]), .B(a[948]), .Z(n1897) );
  NAND U57 ( .A(b[947]), .B(a[947]), .Z(n1895) );
  NAND U58 ( .A(b[946]), .B(a[946]), .Z(n1893) );
  NAND U59 ( .A(b[945]), .B(a[945]), .Z(n1891) );
  NAND U60 ( .A(b[944]), .B(a[944]), .Z(n1889) );
  NAND U61 ( .A(b[943]), .B(a[943]), .Z(n1887) );
  NAND U62 ( .A(b[942]), .B(a[942]), .Z(n1885) );
  NAND U63 ( .A(b[941]), .B(a[941]), .Z(n1883) );
  NAND U64 ( .A(b[940]), .B(a[940]), .Z(n1881) );
  NAND U65 ( .A(b[939]), .B(a[939]), .Z(n1879) );
  NAND U66 ( .A(b[938]), .B(a[938]), .Z(n1877) );
  NAND U67 ( .A(b[937]), .B(a[937]), .Z(n1875) );
  NAND U68 ( .A(b[936]), .B(a[936]), .Z(n1873) );
  NAND U69 ( .A(b[935]), .B(a[935]), .Z(n1871) );
  NAND U70 ( .A(b[934]), .B(a[934]), .Z(n1869) );
  NAND U71 ( .A(b[933]), .B(a[933]), .Z(n1867) );
  NAND U72 ( .A(b[932]), .B(a[932]), .Z(n1865) );
  NAND U73 ( .A(b[931]), .B(a[931]), .Z(n1863) );
  NAND U74 ( .A(b[930]), .B(a[930]), .Z(n1861) );
  NAND U75 ( .A(b[929]), .B(a[929]), .Z(n1859) );
  NAND U76 ( .A(b[928]), .B(a[928]), .Z(n1857) );
  NAND U77 ( .A(b[927]), .B(a[927]), .Z(n1855) );
  NAND U78 ( .A(b[926]), .B(a[926]), .Z(n1853) );
  NAND U79 ( .A(b[925]), .B(a[925]), .Z(n1851) );
  NAND U80 ( .A(b[924]), .B(a[924]), .Z(n1849) );
  NAND U81 ( .A(b[923]), .B(a[923]), .Z(n1847) );
  NAND U82 ( .A(b[922]), .B(a[922]), .Z(n1845) );
  NAND U83 ( .A(b[921]), .B(a[921]), .Z(n1843) );
  NAND U84 ( .A(b[920]), .B(a[920]), .Z(n1841) );
  NAND U85 ( .A(b[919]), .B(a[919]), .Z(n1839) );
  NAND U86 ( .A(b[918]), .B(a[918]), .Z(n1837) );
  NAND U87 ( .A(b[917]), .B(a[917]), .Z(n1835) );
  NAND U88 ( .A(b[916]), .B(a[916]), .Z(n1833) );
  NAND U89 ( .A(b[915]), .B(a[915]), .Z(n1831) );
  NAND U90 ( .A(b[914]), .B(a[914]), .Z(n1829) );
  NAND U91 ( .A(b[913]), .B(a[913]), .Z(n1827) );
  NAND U92 ( .A(b[912]), .B(a[912]), .Z(n1825) );
  NAND U93 ( .A(b[911]), .B(a[911]), .Z(n1823) );
  NAND U94 ( .A(b[910]), .B(a[910]), .Z(n1821) );
  NAND U95 ( .A(b[909]), .B(a[909]), .Z(n1819) );
  NAND U96 ( .A(b[908]), .B(a[908]), .Z(n1817) );
  NAND U97 ( .A(b[907]), .B(a[907]), .Z(n1815) );
  NAND U98 ( .A(b[906]), .B(a[906]), .Z(n1813) );
  NAND U99 ( .A(b[905]), .B(a[905]), .Z(n1811) );
  NAND U100 ( .A(b[904]), .B(a[904]), .Z(n1809) );
  NAND U101 ( .A(b[903]), .B(a[903]), .Z(n1807) );
  NAND U102 ( .A(b[902]), .B(a[902]), .Z(n1805) );
  NAND U103 ( .A(b[901]), .B(a[901]), .Z(n1803) );
  NAND U104 ( .A(b[900]), .B(a[900]), .Z(n1801) );
  NAND U105 ( .A(b[899]), .B(a[899]), .Z(n1799) );
  NAND U106 ( .A(b[898]), .B(a[898]), .Z(n1797) );
  NAND U107 ( .A(b[897]), .B(a[897]), .Z(n1795) );
  NAND U108 ( .A(b[896]), .B(a[896]), .Z(n1793) );
  NAND U109 ( .A(b[895]), .B(a[895]), .Z(n1791) );
  NAND U110 ( .A(b[894]), .B(a[894]), .Z(n1789) );
  NAND U111 ( .A(b[893]), .B(a[893]), .Z(n1787) );
  NAND U112 ( .A(b[892]), .B(a[892]), .Z(n1785) );
  NAND U113 ( .A(b[891]), .B(a[891]), .Z(n1783) );
  NAND U114 ( .A(b[890]), .B(a[890]), .Z(n1781) );
  NAND U115 ( .A(b[889]), .B(a[889]), .Z(n1779) );
  NAND U116 ( .A(b[888]), .B(a[888]), .Z(n1777) );
  NAND U117 ( .A(b[887]), .B(a[887]), .Z(n1775) );
  NAND U118 ( .A(b[886]), .B(a[886]), .Z(n1773) );
  NAND U119 ( .A(b[885]), .B(a[885]), .Z(n1771) );
  NAND U120 ( .A(b[884]), .B(a[884]), .Z(n1769) );
  NAND U121 ( .A(b[883]), .B(a[883]), .Z(n1767) );
  NAND U122 ( .A(b[882]), .B(a[882]), .Z(n1765) );
  NAND U123 ( .A(b[881]), .B(a[881]), .Z(n1763) );
  NAND U124 ( .A(b[880]), .B(a[880]), .Z(n1761) );
  NAND U125 ( .A(b[879]), .B(a[879]), .Z(n1759) );
  NAND U126 ( .A(b[878]), .B(a[878]), .Z(n1757) );
  NAND U127 ( .A(b[877]), .B(a[877]), .Z(n1755) );
  NAND U128 ( .A(b[876]), .B(a[876]), .Z(n1753) );
  NAND U129 ( .A(b[875]), .B(a[875]), .Z(n1751) );
  NAND U130 ( .A(b[874]), .B(a[874]), .Z(n1749) );
  NAND U131 ( .A(b[873]), .B(a[873]), .Z(n1747) );
  NAND U132 ( .A(b[872]), .B(a[872]), .Z(n1745) );
  NAND U133 ( .A(b[871]), .B(a[871]), .Z(n1743) );
  NAND U134 ( .A(b[870]), .B(a[870]), .Z(n1741) );
  NAND U135 ( .A(b[869]), .B(a[869]), .Z(n1739) );
  NAND U136 ( .A(b[868]), .B(a[868]), .Z(n1737) );
  NAND U137 ( .A(b[867]), .B(a[867]), .Z(n1735) );
  NAND U138 ( .A(b[866]), .B(a[866]), .Z(n1733) );
  NAND U139 ( .A(b[865]), .B(a[865]), .Z(n1731) );
  NAND U140 ( .A(b[864]), .B(a[864]), .Z(n1729) );
  NAND U141 ( .A(b[863]), .B(a[863]), .Z(n1727) );
  NAND U142 ( .A(b[862]), .B(a[862]), .Z(n1725) );
  NAND U143 ( .A(b[861]), .B(a[861]), .Z(n1723) );
  NAND U144 ( .A(b[860]), .B(a[860]), .Z(n1721) );
  NAND U145 ( .A(b[859]), .B(a[859]), .Z(n1719) );
  NAND U146 ( .A(b[858]), .B(a[858]), .Z(n1717) );
  NAND U147 ( .A(b[857]), .B(a[857]), .Z(n1715) );
  NAND U148 ( .A(b[856]), .B(a[856]), .Z(n1713) );
  NAND U149 ( .A(b[855]), .B(a[855]), .Z(n1711) );
  NAND U150 ( .A(b[854]), .B(a[854]), .Z(n1709) );
  NAND U151 ( .A(b[853]), .B(a[853]), .Z(n1707) );
  NAND U152 ( .A(b[852]), .B(a[852]), .Z(n1705) );
  NAND U153 ( .A(b[851]), .B(a[851]), .Z(n1703) );
  NAND U154 ( .A(b[850]), .B(a[850]), .Z(n1701) );
  NAND U155 ( .A(b[849]), .B(a[849]), .Z(n1699) );
  NAND U156 ( .A(b[848]), .B(a[848]), .Z(n1697) );
  NAND U157 ( .A(b[847]), .B(a[847]), .Z(n1695) );
  NAND U158 ( .A(b[846]), .B(a[846]), .Z(n1693) );
  NAND U159 ( .A(b[845]), .B(a[845]), .Z(n1691) );
  NAND U160 ( .A(b[844]), .B(a[844]), .Z(n1689) );
  NAND U161 ( .A(b[843]), .B(a[843]), .Z(n1687) );
  NAND U162 ( .A(b[842]), .B(a[842]), .Z(n1685) );
  NAND U163 ( .A(b[841]), .B(a[841]), .Z(n1683) );
  NAND U164 ( .A(b[840]), .B(a[840]), .Z(n1681) );
  NAND U165 ( .A(b[839]), .B(a[839]), .Z(n1679) );
  NAND U166 ( .A(b[838]), .B(a[838]), .Z(n1677) );
  NAND U167 ( .A(b[837]), .B(a[837]), .Z(n1675) );
  NAND U168 ( .A(b[836]), .B(a[836]), .Z(n1673) );
  NAND U169 ( .A(b[835]), .B(a[835]), .Z(n1671) );
  NAND U170 ( .A(b[834]), .B(a[834]), .Z(n1669) );
  NAND U171 ( .A(b[833]), .B(a[833]), .Z(n1667) );
  NAND U172 ( .A(b[832]), .B(a[832]), .Z(n1665) );
  NAND U173 ( .A(b[831]), .B(a[831]), .Z(n1663) );
  NAND U174 ( .A(b[830]), .B(a[830]), .Z(n1661) );
  NAND U175 ( .A(b[829]), .B(a[829]), .Z(n1659) );
  NAND U176 ( .A(b[828]), .B(a[828]), .Z(n1657) );
  NAND U177 ( .A(b[827]), .B(a[827]), .Z(n1655) );
  NAND U178 ( .A(b[826]), .B(a[826]), .Z(n1653) );
  NAND U179 ( .A(b[825]), .B(a[825]), .Z(n1651) );
  NAND U180 ( .A(b[824]), .B(a[824]), .Z(n1649) );
  NAND U181 ( .A(b[823]), .B(a[823]), .Z(n1647) );
  NAND U182 ( .A(b[822]), .B(a[822]), .Z(n1645) );
  NAND U183 ( .A(b[821]), .B(a[821]), .Z(n1643) );
  NAND U184 ( .A(b[820]), .B(a[820]), .Z(n1641) );
  NAND U185 ( .A(b[819]), .B(a[819]), .Z(n1639) );
  NAND U186 ( .A(b[818]), .B(a[818]), .Z(n1637) );
  NAND U187 ( .A(b[817]), .B(a[817]), .Z(n1635) );
  NAND U188 ( .A(b[816]), .B(a[816]), .Z(n1633) );
  NAND U189 ( .A(b[815]), .B(a[815]), .Z(n1631) );
  NAND U190 ( .A(b[814]), .B(a[814]), .Z(n1629) );
  NAND U191 ( .A(b[813]), .B(a[813]), .Z(n1627) );
  NAND U192 ( .A(b[812]), .B(a[812]), .Z(n1625) );
  NAND U193 ( .A(b[811]), .B(a[811]), .Z(n1623) );
  NAND U194 ( .A(b[810]), .B(a[810]), .Z(n1621) );
  NAND U195 ( .A(b[809]), .B(a[809]), .Z(n1619) );
  NAND U196 ( .A(b[808]), .B(a[808]), .Z(n1617) );
  NAND U197 ( .A(b[807]), .B(a[807]), .Z(n1615) );
  NAND U198 ( .A(b[806]), .B(a[806]), .Z(n1613) );
  NAND U199 ( .A(b[805]), .B(a[805]), .Z(n1611) );
  NAND U200 ( .A(b[804]), .B(a[804]), .Z(n1609) );
  NAND U201 ( .A(b[803]), .B(a[803]), .Z(n1607) );
  NAND U202 ( .A(b[802]), .B(a[802]), .Z(n1605) );
  NAND U203 ( .A(b[801]), .B(a[801]), .Z(n1603) );
  NAND U204 ( .A(b[800]), .B(a[800]), .Z(n1601) );
  NAND U205 ( .A(b[799]), .B(a[799]), .Z(n1599) );
  NAND U206 ( .A(b[798]), .B(a[798]), .Z(n1597) );
  NAND U207 ( .A(b[797]), .B(a[797]), .Z(n1595) );
  NAND U208 ( .A(b[796]), .B(a[796]), .Z(n1593) );
  NAND U209 ( .A(b[795]), .B(a[795]), .Z(n1591) );
  NAND U210 ( .A(b[794]), .B(a[794]), .Z(n1589) );
  NAND U211 ( .A(b[793]), .B(a[793]), .Z(n1587) );
  NAND U212 ( .A(b[792]), .B(a[792]), .Z(n1585) );
  NAND U213 ( .A(b[791]), .B(a[791]), .Z(n1583) );
  NAND U214 ( .A(b[790]), .B(a[790]), .Z(n1581) );
  NAND U215 ( .A(b[789]), .B(a[789]), .Z(n1579) );
  NAND U216 ( .A(b[788]), .B(a[788]), .Z(n1577) );
  NAND U217 ( .A(b[787]), .B(a[787]), .Z(n1575) );
  NAND U218 ( .A(b[786]), .B(a[786]), .Z(n1573) );
  NAND U219 ( .A(b[785]), .B(a[785]), .Z(n1571) );
  NAND U220 ( .A(b[784]), .B(a[784]), .Z(n1569) );
  NAND U221 ( .A(b[783]), .B(a[783]), .Z(n1567) );
  NAND U222 ( .A(b[782]), .B(a[782]), .Z(n1565) );
  NAND U223 ( .A(b[781]), .B(a[781]), .Z(n1563) );
  NAND U224 ( .A(b[780]), .B(a[780]), .Z(n1561) );
  NAND U225 ( .A(b[779]), .B(a[779]), .Z(n1559) );
  NAND U226 ( .A(b[778]), .B(a[778]), .Z(n1557) );
  NAND U227 ( .A(b[777]), .B(a[777]), .Z(n1555) );
  NAND U228 ( .A(b[776]), .B(a[776]), .Z(n1553) );
  NAND U229 ( .A(b[775]), .B(a[775]), .Z(n1551) );
  NAND U230 ( .A(b[774]), .B(a[774]), .Z(n1549) );
  NAND U231 ( .A(b[773]), .B(a[773]), .Z(n1547) );
  NAND U232 ( .A(b[772]), .B(a[772]), .Z(n1545) );
  NAND U233 ( .A(b[771]), .B(a[771]), .Z(n1543) );
  NAND U234 ( .A(b[770]), .B(a[770]), .Z(n1541) );
  NAND U235 ( .A(b[769]), .B(a[769]), .Z(n1539) );
  NAND U236 ( .A(b[768]), .B(a[768]), .Z(n1537) );
  NAND U237 ( .A(b[767]), .B(a[767]), .Z(n1535) );
  NAND U238 ( .A(b[766]), .B(a[766]), .Z(n1533) );
  NAND U239 ( .A(b[765]), .B(a[765]), .Z(n1531) );
  NAND U240 ( .A(b[764]), .B(a[764]), .Z(n1529) );
  NAND U241 ( .A(b[763]), .B(a[763]), .Z(n1527) );
  NAND U242 ( .A(b[762]), .B(a[762]), .Z(n1525) );
  NAND U243 ( .A(b[761]), .B(a[761]), .Z(n1523) );
  NAND U244 ( .A(b[760]), .B(a[760]), .Z(n1521) );
  NAND U245 ( .A(b[759]), .B(a[759]), .Z(n1519) );
  NAND U246 ( .A(b[758]), .B(a[758]), .Z(n1517) );
  NAND U247 ( .A(b[757]), .B(a[757]), .Z(n1515) );
  NAND U248 ( .A(b[756]), .B(a[756]), .Z(n1513) );
  NAND U249 ( .A(b[755]), .B(a[755]), .Z(n1511) );
  NAND U250 ( .A(b[754]), .B(a[754]), .Z(n1509) );
  NAND U251 ( .A(b[753]), .B(a[753]), .Z(n1507) );
  NAND U252 ( .A(b[752]), .B(a[752]), .Z(n1505) );
  NAND U253 ( .A(b[751]), .B(a[751]), .Z(n1503) );
  NAND U254 ( .A(b[750]), .B(a[750]), .Z(n1501) );
  NAND U255 ( .A(b[749]), .B(a[749]), .Z(n1499) );
  NAND U256 ( .A(b[748]), .B(a[748]), .Z(n1497) );
  NAND U257 ( .A(b[747]), .B(a[747]), .Z(n1495) );
  NAND U258 ( .A(b[746]), .B(a[746]), .Z(n1493) );
  NAND U259 ( .A(b[745]), .B(a[745]), .Z(n1491) );
  NAND U260 ( .A(b[744]), .B(a[744]), .Z(n1489) );
  NAND U261 ( .A(b[743]), .B(a[743]), .Z(n1487) );
  NAND U262 ( .A(b[742]), .B(a[742]), .Z(n1485) );
  NAND U263 ( .A(b[741]), .B(a[741]), .Z(n1483) );
  NAND U264 ( .A(b[740]), .B(a[740]), .Z(n1481) );
  NAND U265 ( .A(b[739]), .B(a[739]), .Z(n1479) );
  NAND U266 ( .A(b[738]), .B(a[738]), .Z(n1477) );
  NAND U267 ( .A(b[737]), .B(a[737]), .Z(n1475) );
  NAND U268 ( .A(b[736]), .B(a[736]), .Z(n1473) );
  NAND U269 ( .A(b[735]), .B(a[735]), .Z(n1471) );
  NAND U270 ( .A(b[734]), .B(a[734]), .Z(n1469) );
  NAND U271 ( .A(b[733]), .B(a[733]), .Z(n1467) );
  NAND U272 ( .A(b[732]), .B(a[732]), .Z(n1465) );
  NAND U273 ( .A(b[731]), .B(a[731]), .Z(n1463) );
  NAND U274 ( .A(b[730]), .B(a[730]), .Z(n1461) );
  NAND U275 ( .A(b[729]), .B(a[729]), .Z(n1459) );
  NAND U276 ( .A(b[728]), .B(a[728]), .Z(n1457) );
  NAND U277 ( .A(b[727]), .B(a[727]), .Z(n1455) );
  NAND U278 ( .A(b[726]), .B(a[726]), .Z(n1453) );
  NAND U279 ( .A(b[725]), .B(a[725]), .Z(n1451) );
  NAND U280 ( .A(b[724]), .B(a[724]), .Z(n1449) );
  NAND U281 ( .A(b[723]), .B(a[723]), .Z(n1447) );
  NAND U282 ( .A(b[722]), .B(a[722]), .Z(n1445) );
  NAND U283 ( .A(b[721]), .B(a[721]), .Z(n1443) );
  NAND U284 ( .A(b[720]), .B(a[720]), .Z(n1441) );
  NAND U285 ( .A(b[719]), .B(a[719]), .Z(n1439) );
  NAND U286 ( .A(b[718]), .B(a[718]), .Z(n1437) );
  NAND U287 ( .A(b[717]), .B(a[717]), .Z(n1435) );
  NAND U288 ( .A(b[716]), .B(a[716]), .Z(n1433) );
  NAND U289 ( .A(b[715]), .B(a[715]), .Z(n1431) );
  NAND U290 ( .A(b[714]), .B(a[714]), .Z(n1429) );
  NAND U291 ( .A(b[713]), .B(a[713]), .Z(n1427) );
  NAND U292 ( .A(b[712]), .B(a[712]), .Z(n1425) );
  NAND U293 ( .A(b[711]), .B(a[711]), .Z(n1423) );
  NAND U294 ( .A(b[710]), .B(a[710]), .Z(n1421) );
  NAND U295 ( .A(b[709]), .B(a[709]), .Z(n1419) );
  NAND U296 ( .A(b[708]), .B(a[708]), .Z(n1417) );
  NAND U297 ( .A(b[707]), .B(a[707]), .Z(n1415) );
  NAND U298 ( .A(b[706]), .B(a[706]), .Z(n1413) );
  NAND U299 ( .A(b[705]), .B(a[705]), .Z(n1411) );
  NAND U300 ( .A(b[704]), .B(a[704]), .Z(n1409) );
  NAND U301 ( .A(b[703]), .B(a[703]), .Z(n1407) );
  NAND U302 ( .A(b[702]), .B(a[702]), .Z(n1405) );
  NAND U303 ( .A(b[701]), .B(a[701]), .Z(n1403) );
  NAND U304 ( .A(b[700]), .B(a[700]), .Z(n1401) );
  NAND U305 ( .A(b[699]), .B(a[699]), .Z(n1399) );
  NAND U306 ( .A(b[698]), .B(a[698]), .Z(n1397) );
  NAND U307 ( .A(b[697]), .B(a[697]), .Z(n1395) );
  NAND U308 ( .A(b[696]), .B(a[696]), .Z(n1393) );
  NAND U309 ( .A(b[695]), .B(a[695]), .Z(n1391) );
  NAND U310 ( .A(b[694]), .B(a[694]), .Z(n1389) );
  NAND U311 ( .A(b[693]), .B(a[693]), .Z(n1387) );
  NAND U312 ( .A(b[692]), .B(a[692]), .Z(n1385) );
  NAND U313 ( .A(b[691]), .B(a[691]), .Z(n1383) );
  NAND U314 ( .A(b[690]), .B(a[690]), .Z(n1381) );
  NAND U315 ( .A(b[689]), .B(a[689]), .Z(n1379) );
  NAND U316 ( .A(b[688]), .B(a[688]), .Z(n1377) );
  NAND U317 ( .A(b[687]), .B(a[687]), .Z(n1375) );
  NAND U318 ( .A(b[686]), .B(a[686]), .Z(n1373) );
  NAND U319 ( .A(b[685]), .B(a[685]), .Z(n1371) );
  NAND U320 ( .A(b[684]), .B(a[684]), .Z(n1369) );
  NAND U321 ( .A(b[683]), .B(a[683]), .Z(n1367) );
  NAND U322 ( .A(b[682]), .B(a[682]), .Z(n1365) );
  NAND U323 ( .A(b[681]), .B(a[681]), .Z(n1363) );
  NAND U324 ( .A(b[680]), .B(a[680]), .Z(n1361) );
  NAND U325 ( .A(b[679]), .B(a[679]), .Z(n1359) );
  NAND U326 ( .A(b[678]), .B(a[678]), .Z(n1357) );
  NAND U327 ( .A(b[677]), .B(a[677]), .Z(n1355) );
  NAND U328 ( .A(b[676]), .B(a[676]), .Z(n1353) );
  NAND U329 ( .A(b[675]), .B(a[675]), .Z(n1351) );
  NAND U330 ( .A(b[674]), .B(a[674]), .Z(n1349) );
  NAND U331 ( .A(b[673]), .B(a[673]), .Z(n1347) );
  NAND U332 ( .A(b[672]), .B(a[672]), .Z(n1345) );
  NAND U333 ( .A(b[671]), .B(a[671]), .Z(n1343) );
  NAND U334 ( .A(b[670]), .B(a[670]), .Z(n1341) );
  NAND U335 ( .A(b[669]), .B(a[669]), .Z(n1339) );
  NAND U336 ( .A(b[668]), .B(a[668]), .Z(n1337) );
  NAND U337 ( .A(b[667]), .B(a[667]), .Z(n1335) );
  NAND U338 ( .A(b[666]), .B(a[666]), .Z(n1333) );
  NAND U339 ( .A(b[665]), .B(a[665]), .Z(n1331) );
  NAND U340 ( .A(b[664]), .B(a[664]), .Z(n1329) );
  NAND U341 ( .A(b[663]), .B(a[663]), .Z(n1327) );
  NAND U342 ( .A(b[662]), .B(a[662]), .Z(n1325) );
  NAND U343 ( .A(b[661]), .B(a[661]), .Z(n1323) );
  NAND U344 ( .A(b[660]), .B(a[660]), .Z(n1321) );
  NAND U345 ( .A(b[659]), .B(a[659]), .Z(n1319) );
  NAND U346 ( .A(b[658]), .B(a[658]), .Z(n1317) );
  NAND U347 ( .A(b[657]), .B(a[657]), .Z(n1315) );
  NAND U348 ( .A(b[656]), .B(a[656]), .Z(n1313) );
  NAND U349 ( .A(b[655]), .B(a[655]), .Z(n1311) );
  NAND U350 ( .A(b[654]), .B(a[654]), .Z(n1309) );
  NAND U351 ( .A(b[653]), .B(a[653]), .Z(n1307) );
  NAND U352 ( .A(b[652]), .B(a[652]), .Z(n1305) );
  NAND U353 ( .A(b[651]), .B(a[651]), .Z(n1303) );
  NAND U354 ( .A(b[650]), .B(a[650]), .Z(n1301) );
  NAND U355 ( .A(b[649]), .B(a[649]), .Z(n1299) );
  NAND U356 ( .A(b[648]), .B(a[648]), .Z(n1297) );
  NAND U357 ( .A(b[647]), .B(a[647]), .Z(n1295) );
  NAND U358 ( .A(b[646]), .B(a[646]), .Z(n1293) );
  NAND U359 ( .A(b[645]), .B(a[645]), .Z(n1291) );
  NAND U360 ( .A(b[644]), .B(a[644]), .Z(n1289) );
  NAND U361 ( .A(b[643]), .B(a[643]), .Z(n1287) );
  NAND U362 ( .A(b[642]), .B(a[642]), .Z(n1285) );
  NAND U363 ( .A(b[641]), .B(a[641]), .Z(n1283) );
  NAND U364 ( .A(b[640]), .B(a[640]), .Z(n1281) );
  NAND U365 ( .A(b[639]), .B(a[639]), .Z(n1279) );
  NAND U366 ( .A(b[638]), .B(a[638]), .Z(n1277) );
  NAND U367 ( .A(b[637]), .B(a[637]), .Z(n1275) );
  NAND U368 ( .A(b[636]), .B(a[636]), .Z(n1273) );
  NAND U369 ( .A(b[635]), .B(a[635]), .Z(n1271) );
  NAND U370 ( .A(b[634]), .B(a[634]), .Z(n1269) );
  NAND U371 ( .A(b[633]), .B(a[633]), .Z(n1267) );
  NAND U372 ( .A(b[632]), .B(a[632]), .Z(n1265) );
  NAND U373 ( .A(b[631]), .B(a[631]), .Z(n1263) );
  NAND U374 ( .A(b[630]), .B(a[630]), .Z(n1261) );
  NAND U375 ( .A(b[629]), .B(a[629]), .Z(n1259) );
  NAND U376 ( .A(b[628]), .B(a[628]), .Z(n1257) );
  NAND U377 ( .A(b[627]), .B(a[627]), .Z(n1255) );
  NAND U378 ( .A(b[626]), .B(a[626]), .Z(n1253) );
  NAND U379 ( .A(b[625]), .B(a[625]), .Z(n1251) );
  NAND U380 ( .A(b[624]), .B(a[624]), .Z(n1249) );
  NAND U381 ( .A(b[623]), .B(a[623]), .Z(n1247) );
  NAND U382 ( .A(b[622]), .B(a[622]), .Z(n1245) );
  NAND U383 ( .A(b[621]), .B(a[621]), .Z(n1243) );
  NAND U384 ( .A(b[620]), .B(a[620]), .Z(n1241) );
  NAND U385 ( .A(b[619]), .B(a[619]), .Z(n1239) );
  NAND U386 ( .A(b[618]), .B(a[618]), .Z(n1237) );
  NAND U387 ( .A(b[617]), .B(a[617]), .Z(n1235) );
  NAND U388 ( .A(b[616]), .B(a[616]), .Z(n1233) );
  NAND U389 ( .A(b[615]), .B(a[615]), .Z(n1231) );
  NAND U390 ( .A(b[614]), .B(a[614]), .Z(n1229) );
  NAND U391 ( .A(b[613]), .B(a[613]), .Z(n1227) );
  NAND U392 ( .A(b[612]), .B(a[612]), .Z(n1225) );
  NAND U393 ( .A(b[611]), .B(a[611]), .Z(n1223) );
  NAND U394 ( .A(b[610]), .B(a[610]), .Z(n1221) );
  NAND U395 ( .A(b[609]), .B(a[609]), .Z(n1219) );
  NAND U396 ( .A(b[608]), .B(a[608]), .Z(n1217) );
  NAND U397 ( .A(b[607]), .B(a[607]), .Z(n1215) );
  NAND U398 ( .A(b[606]), .B(a[606]), .Z(n1213) );
  NAND U399 ( .A(b[605]), .B(a[605]), .Z(n1211) );
  NAND U400 ( .A(b[604]), .B(a[604]), .Z(n1209) );
  NAND U401 ( .A(b[603]), .B(a[603]), .Z(n1207) );
  NAND U402 ( .A(b[602]), .B(a[602]), .Z(n1205) );
  NAND U403 ( .A(b[601]), .B(a[601]), .Z(n1203) );
  NAND U404 ( .A(b[600]), .B(a[600]), .Z(n1201) );
  NAND U405 ( .A(b[599]), .B(a[599]), .Z(n1199) );
  NAND U406 ( .A(b[598]), .B(a[598]), .Z(n1197) );
  NAND U407 ( .A(b[597]), .B(a[597]), .Z(n1195) );
  NAND U408 ( .A(b[596]), .B(a[596]), .Z(n1193) );
  NAND U409 ( .A(b[595]), .B(a[595]), .Z(n1191) );
  NAND U410 ( .A(b[594]), .B(a[594]), .Z(n1189) );
  NAND U411 ( .A(b[593]), .B(a[593]), .Z(n1187) );
  NAND U412 ( .A(b[592]), .B(a[592]), .Z(n1185) );
  NAND U413 ( .A(b[591]), .B(a[591]), .Z(n1183) );
  NAND U414 ( .A(b[590]), .B(a[590]), .Z(n1181) );
  NAND U415 ( .A(b[589]), .B(a[589]), .Z(n1179) );
  NAND U416 ( .A(b[588]), .B(a[588]), .Z(n1177) );
  NAND U417 ( .A(b[587]), .B(a[587]), .Z(n1175) );
  NAND U418 ( .A(b[586]), .B(a[586]), .Z(n1173) );
  NAND U419 ( .A(b[585]), .B(a[585]), .Z(n1171) );
  NAND U420 ( .A(b[584]), .B(a[584]), .Z(n1169) );
  NAND U421 ( .A(b[583]), .B(a[583]), .Z(n1167) );
  NAND U422 ( .A(b[582]), .B(a[582]), .Z(n1165) );
  NAND U423 ( .A(b[581]), .B(a[581]), .Z(n1163) );
  NAND U424 ( .A(b[580]), .B(a[580]), .Z(n1161) );
  NAND U425 ( .A(b[579]), .B(a[579]), .Z(n1159) );
  NAND U426 ( .A(b[578]), .B(a[578]), .Z(n1157) );
  NAND U427 ( .A(b[577]), .B(a[577]), .Z(n1155) );
  NAND U428 ( .A(b[576]), .B(a[576]), .Z(n1153) );
  NAND U429 ( .A(b[575]), .B(a[575]), .Z(n1151) );
  NAND U430 ( .A(b[574]), .B(a[574]), .Z(n1149) );
  NAND U431 ( .A(b[573]), .B(a[573]), .Z(n1147) );
  NAND U432 ( .A(b[572]), .B(a[572]), .Z(n1145) );
  NAND U433 ( .A(b[571]), .B(a[571]), .Z(n1143) );
  NAND U434 ( .A(b[570]), .B(a[570]), .Z(n1141) );
  NAND U435 ( .A(b[569]), .B(a[569]), .Z(n1139) );
  NAND U436 ( .A(b[568]), .B(a[568]), .Z(n1137) );
  NAND U437 ( .A(b[567]), .B(a[567]), .Z(n1135) );
  NAND U438 ( .A(b[566]), .B(a[566]), .Z(n1133) );
  NAND U439 ( .A(b[565]), .B(a[565]), .Z(n1131) );
  NAND U440 ( .A(b[564]), .B(a[564]), .Z(n1129) );
  NAND U441 ( .A(b[563]), .B(a[563]), .Z(n1127) );
  NAND U442 ( .A(b[562]), .B(a[562]), .Z(n1125) );
  NAND U443 ( .A(b[561]), .B(a[561]), .Z(n1123) );
  NAND U444 ( .A(b[560]), .B(a[560]), .Z(n1121) );
  NAND U445 ( .A(b[559]), .B(a[559]), .Z(n1119) );
  NAND U446 ( .A(b[558]), .B(a[558]), .Z(n1117) );
  NAND U447 ( .A(b[557]), .B(a[557]), .Z(n1115) );
  NAND U448 ( .A(b[556]), .B(a[556]), .Z(n1113) );
  NAND U449 ( .A(b[555]), .B(a[555]), .Z(n1111) );
  NAND U450 ( .A(b[554]), .B(a[554]), .Z(n1109) );
  NAND U451 ( .A(b[553]), .B(a[553]), .Z(n1107) );
  NAND U452 ( .A(b[552]), .B(a[552]), .Z(n1105) );
  NAND U453 ( .A(b[551]), .B(a[551]), .Z(n1103) );
  NAND U454 ( .A(b[550]), .B(a[550]), .Z(n1101) );
  NAND U455 ( .A(b[549]), .B(a[549]), .Z(n1099) );
  NAND U456 ( .A(b[548]), .B(a[548]), .Z(n1097) );
  NAND U457 ( .A(b[547]), .B(a[547]), .Z(n1095) );
  NAND U458 ( .A(b[546]), .B(a[546]), .Z(n1093) );
  NAND U459 ( .A(b[545]), .B(a[545]), .Z(n1091) );
  NAND U460 ( .A(b[544]), .B(a[544]), .Z(n1089) );
  NAND U461 ( .A(b[543]), .B(a[543]), .Z(n1087) );
  NAND U462 ( .A(b[542]), .B(a[542]), .Z(n1085) );
  NAND U463 ( .A(b[541]), .B(a[541]), .Z(n1083) );
  NAND U464 ( .A(b[540]), .B(a[540]), .Z(n1081) );
  NAND U465 ( .A(b[539]), .B(a[539]), .Z(n1079) );
  NAND U466 ( .A(b[538]), .B(a[538]), .Z(n1077) );
  NAND U467 ( .A(b[537]), .B(a[537]), .Z(n1075) );
  NAND U468 ( .A(b[536]), .B(a[536]), .Z(n1073) );
  NAND U469 ( .A(b[535]), .B(a[535]), .Z(n1071) );
  NAND U470 ( .A(b[534]), .B(a[534]), .Z(n1069) );
  NAND U471 ( .A(b[533]), .B(a[533]), .Z(n1067) );
  NAND U472 ( .A(b[532]), .B(a[532]), .Z(n1065) );
  NAND U473 ( .A(b[531]), .B(a[531]), .Z(n1063) );
  NAND U474 ( .A(b[530]), .B(a[530]), .Z(n1061) );
  NAND U475 ( .A(b[529]), .B(a[529]), .Z(n1059) );
  NAND U476 ( .A(b[528]), .B(a[528]), .Z(n1057) );
  NAND U477 ( .A(b[527]), .B(a[527]), .Z(n1055) );
  NAND U478 ( .A(b[526]), .B(a[526]), .Z(n1053) );
  NAND U479 ( .A(b[525]), .B(a[525]), .Z(n1051) );
  NAND U480 ( .A(b[524]), .B(a[524]), .Z(n1049) );
  NAND U481 ( .A(b[523]), .B(a[523]), .Z(n1047) );
  NAND U482 ( .A(b[522]), .B(a[522]), .Z(n1045) );
  NAND U483 ( .A(b[521]), .B(a[521]), .Z(n1043) );
  NAND U484 ( .A(b[520]), .B(a[520]), .Z(n1041) );
  NAND U485 ( .A(b[519]), .B(a[519]), .Z(n1039) );
  NAND U486 ( .A(b[518]), .B(a[518]), .Z(n1037) );
  NAND U487 ( .A(b[517]), .B(a[517]), .Z(n1035) );
  NAND U488 ( .A(b[516]), .B(a[516]), .Z(n1033) );
  NAND U489 ( .A(b[515]), .B(a[515]), .Z(n1031) );
  NAND U490 ( .A(b[514]), .B(a[514]), .Z(n1029) );
  NAND U491 ( .A(b[513]), .B(a[513]), .Z(n1027) );
  NAND U492 ( .A(b[512]), .B(a[512]), .Z(n1025) );
  NAND U493 ( .A(b[511]), .B(a[511]), .Z(n1023) );
  NAND U494 ( .A(b[510]), .B(a[510]), .Z(n1021) );
  NAND U495 ( .A(b[509]), .B(a[509]), .Z(n1019) );
  NAND U496 ( .A(b[508]), .B(a[508]), .Z(n1017) );
  NAND U497 ( .A(b[507]), .B(a[507]), .Z(n1015) );
  NAND U498 ( .A(b[506]), .B(a[506]), .Z(n1013) );
  NAND U499 ( .A(b[505]), .B(a[505]), .Z(n1011) );
  NAND U500 ( .A(b[504]), .B(a[504]), .Z(n1009) );
  NAND U501 ( .A(b[503]), .B(a[503]), .Z(n1007) );
  NAND U502 ( .A(b[502]), .B(a[502]), .Z(n1005) );
  NAND U503 ( .A(b[501]), .B(a[501]), .Z(n1003) );
  NAND U504 ( .A(b[500]), .B(a[500]), .Z(n1001) );
  NAND U505 ( .A(b[499]), .B(a[499]), .Z(n999) );
  NAND U506 ( .A(b[498]), .B(a[498]), .Z(n997) );
  NAND U507 ( .A(b[497]), .B(a[497]), .Z(n995) );
  NAND U508 ( .A(b[496]), .B(a[496]), .Z(n993) );
  NAND U509 ( .A(b[495]), .B(a[495]), .Z(n991) );
  NAND U510 ( .A(b[494]), .B(a[494]), .Z(n989) );
  NAND U511 ( .A(b[493]), .B(a[493]), .Z(n987) );
  NAND U512 ( .A(b[492]), .B(a[492]), .Z(n985) );
  NAND U513 ( .A(b[491]), .B(a[491]), .Z(n983) );
  NAND U514 ( .A(b[490]), .B(a[490]), .Z(n981) );
  NAND U515 ( .A(b[489]), .B(a[489]), .Z(n979) );
  NAND U516 ( .A(b[488]), .B(a[488]), .Z(n977) );
  NAND U517 ( .A(b[487]), .B(a[487]), .Z(n975) );
  NAND U518 ( .A(b[486]), .B(a[486]), .Z(n973) );
  NAND U519 ( .A(b[485]), .B(a[485]), .Z(n971) );
  NAND U520 ( .A(b[484]), .B(a[484]), .Z(n969) );
  NAND U521 ( .A(b[483]), .B(a[483]), .Z(n967) );
  NAND U522 ( .A(b[482]), .B(a[482]), .Z(n965) );
  NAND U523 ( .A(b[481]), .B(a[481]), .Z(n963) );
  NAND U524 ( .A(b[480]), .B(a[480]), .Z(n961) );
  NAND U525 ( .A(b[479]), .B(a[479]), .Z(n959) );
  NAND U526 ( .A(b[478]), .B(a[478]), .Z(n957) );
  NAND U527 ( .A(b[477]), .B(a[477]), .Z(n955) );
  NAND U528 ( .A(b[476]), .B(a[476]), .Z(n953) );
  NAND U529 ( .A(b[475]), .B(a[475]), .Z(n951) );
  NAND U530 ( .A(b[474]), .B(a[474]), .Z(n949) );
  NAND U531 ( .A(b[473]), .B(a[473]), .Z(n947) );
  NAND U532 ( .A(b[472]), .B(a[472]), .Z(n945) );
  NAND U533 ( .A(b[471]), .B(a[471]), .Z(n943) );
  NAND U534 ( .A(b[470]), .B(a[470]), .Z(n941) );
  NAND U535 ( .A(b[469]), .B(a[469]), .Z(n939) );
  NAND U536 ( .A(b[468]), .B(a[468]), .Z(n937) );
  NAND U537 ( .A(b[467]), .B(a[467]), .Z(n935) );
  NAND U538 ( .A(b[466]), .B(a[466]), .Z(n933) );
  NAND U539 ( .A(b[465]), .B(a[465]), .Z(n931) );
  NAND U540 ( .A(b[464]), .B(a[464]), .Z(n929) );
  NAND U541 ( .A(b[463]), .B(a[463]), .Z(n927) );
  NAND U542 ( .A(b[462]), .B(a[462]), .Z(n925) );
  NAND U543 ( .A(b[461]), .B(a[461]), .Z(n923) );
  NAND U544 ( .A(b[460]), .B(a[460]), .Z(n921) );
  NAND U545 ( .A(b[459]), .B(a[459]), .Z(n919) );
  NAND U546 ( .A(b[458]), .B(a[458]), .Z(n917) );
  NAND U547 ( .A(b[457]), .B(a[457]), .Z(n915) );
  NAND U548 ( .A(b[456]), .B(a[456]), .Z(n913) );
  NAND U549 ( .A(b[455]), .B(a[455]), .Z(n911) );
  NAND U550 ( .A(b[454]), .B(a[454]), .Z(n909) );
  NAND U551 ( .A(b[453]), .B(a[453]), .Z(n907) );
  NAND U552 ( .A(b[452]), .B(a[452]), .Z(n905) );
  NAND U553 ( .A(b[451]), .B(a[451]), .Z(n903) );
  NAND U554 ( .A(b[450]), .B(a[450]), .Z(n901) );
  NAND U555 ( .A(b[449]), .B(a[449]), .Z(n899) );
  NAND U556 ( .A(b[448]), .B(a[448]), .Z(n897) );
  NAND U557 ( .A(b[447]), .B(a[447]), .Z(n895) );
  NAND U558 ( .A(b[446]), .B(a[446]), .Z(n893) );
  NAND U559 ( .A(b[445]), .B(a[445]), .Z(n891) );
  NAND U560 ( .A(b[444]), .B(a[444]), .Z(n889) );
  NAND U561 ( .A(b[443]), .B(a[443]), .Z(n887) );
  NAND U562 ( .A(b[442]), .B(a[442]), .Z(n885) );
  NAND U563 ( .A(b[441]), .B(a[441]), .Z(n883) );
  NAND U564 ( .A(b[440]), .B(a[440]), .Z(n881) );
  NAND U565 ( .A(b[439]), .B(a[439]), .Z(n879) );
  NAND U566 ( .A(b[438]), .B(a[438]), .Z(n877) );
  NAND U567 ( .A(b[437]), .B(a[437]), .Z(n875) );
  NAND U568 ( .A(b[436]), .B(a[436]), .Z(n873) );
  NAND U569 ( .A(b[435]), .B(a[435]), .Z(n871) );
  NAND U570 ( .A(b[434]), .B(a[434]), .Z(n869) );
  NAND U571 ( .A(b[433]), .B(a[433]), .Z(n867) );
  NAND U572 ( .A(b[432]), .B(a[432]), .Z(n865) );
  NAND U573 ( .A(b[431]), .B(a[431]), .Z(n863) );
  NAND U574 ( .A(b[430]), .B(a[430]), .Z(n861) );
  NAND U575 ( .A(b[429]), .B(a[429]), .Z(n859) );
  NAND U576 ( .A(b[428]), .B(a[428]), .Z(n857) );
  NAND U577 ( .A(b[427]), .B(a[427]), .Z(n855) );
  NAND U578 ( .A(b[426]), .B(a[426]), .Z(n853) );
  NAND U579 ( .A(b[425]), .B(a[425]), .Z(n851) );
  NAND U580 ( .A(b[424]), .B(a[424]), .Z(n849) );
  NAND U581 ( .A(b[423]), .B(a[423]), .Z(n847) );
  NAND U582 ( .A(b[422]), .B(a[422]), .Z(n845) );
  NAND U583 ( .A(b[421]), .B(a[421]), .Z(n843) );
  NAND U584 ( .A(b[420]), .B(a[420]), .Z(n841) );
  NAND U585 ( .A(b[419]), .B(a[419]), .Z(n839) );
  NAND U586 ( .A(b[418]), .B(a[418]), .Z(n837) );
  NAND U587 ( .A(b[417]), .B(a[417]), .Z(n835) );
  NAND U588 ( .A(b[416]), .B(a[416]), .Z(n833) );
  NAND U589 ( .A(b[415]), .B(a[415]), .Z(n831) );
  NAND U590 ( .A(b[414]), .B(a[414]), .Z(n829) );
  NAND U591 ( .A(b[413]), .B(a[413]), .Z(n827) );
  NAND U592 ( .A(b[412]), .B(a[412]), .Z(n825) );
  NAND U593 ( .A(b[411]), .B(a[411]), .Z(n823) );
  NAND U594 ( .A(b[410]), .B(a[410]), .Z(n821) );
  NAND U595 ( .A(b[409]), .B(a[409]), .Z(n819) );
  NAND U596 ( .A(b[408]), .B(a[408]), .Z(n817) );
  NAND U597 ( .A(b[407]), .B(a[407]), .Z(n815) );
  NAND U598 ( .A(b[406]), .B(a[406]), .Z(n813) );
  NAND U599 ( .A(b[405]), .B(a[405]), .Z(n811) );
  NAND U600 ( .A(b[404]), .B(a[404]), .Z(n809) );
  NAND U601 ( .A(b[403]), .B(a[403]), .Z(n807) );
  NAND U602 ( .A(b[402]), .B(a[402]), .Z(n805) );
  NAND U603 ( .A(b[401]), .B(a[401]), .Z(n803) );
  NAND U604 ( .A(b[400]), .B(a[400]), .Z(n801) );
  NAND U605 ( .A(b[399]), .B(a[399]), .Z(n799) );
  NAND U606 ( .A(b[398]), .B(a[398]), .Z(n797) );
  NAND U607 ( .A(b[397]), .B(a[397]), .Z(n795) );
  NAND U608 ( .A(b[396]), .B(a[396]), .Z(n793) );
  NAND U609 ( .A(b[395]), .B(a[395]), .Z(n791) );
  NAND U610 ( .A(b[394]), .B(a[394]), .Z(n789) );
  NAND U611 ( .A(b[393]), .B(a[393]), .Z(n787) );
  NAND U612 ( .A(b[392]), .B(a[392]), .Z(n785) );
  NAND U613 ( .A(b[391]), .B(a[391]), .Z(n783) );
  NAND U614 ( .A(b[390]), .B(a[390]), .Z(n781) );
  NAND U615 ( .A(b[389]), .B(a[389]), .Z(n779) );
  NAND U616 ( .A(b[388]), .B(a[388]), .Z(n777) );
  NAND U617 ( .A(b[387]), .B(a[387]), .Z(n775) );
  NAND U618 ( .A(b[386]), .B(a[386]), .Z(n773) );
  NAND U619 ( .A(b[385]), .B(a[385]), .Z(n771) );
  NAND U620 ( .A(b[384]), .B(a[384]), .Z(n769) );
  NAND U621 ( .A(b[383]), .B(a[383]), .Z(n767) );
  NAND U622 ( .A(b[382]), .B(a[382]), .Z(n765) );
  NAND U623 ( .A(b[381]), .B(a[381]), .Z(n763) );
  NAND U624 ( .A(b[380]), .B(a[380]), .Z(n761) );
  NAND U625 ( .A(b[379]), .B(a[379]), .Z(n759) );
  NAND U626 ( .A(b[378]), .B(a[378]), .Z(n757) );
  NAND U627 ( .A(b[377]), .B(a[377]), .Z(n755) );
  NAND U628 ( .A(b[376]), .B(a[376]), .Z(n753) );
  NAND U629 ( .A(b[375]), .B(a[375]), .Z(n751) );
  NAND U630 ( .A(b[374]), .B(a[374]), .Z(n749) );
  NAND U631 ( .A(b[373]), .B(a[373]), .Z(n747) );
  NAND U632 ( .A(b[372]), .B(a[372]), .Z(n745) );
  NAND U633 ( .A(b[371]), .B(a[371]), .Z(n743) );
  NAND U634 ( .A(b[370]), .B(a[370]), .Z(n741) );
  NAND U635 ( .A(b[369]), .B(a[369]), .Z(n739) );
  NAND U636 ( .A(b[368]), .B(a[368]), .Z(n737) );
  NAND U637 ( .A(b[367]), .B(a[367]), .Z(n735) );
  NAND U638 ( .A(b[366]), .B(a[366]), .Z(n733) );
  NAND U639 ( .A(b[365]), .B(a[365]), .Z(n731) );
  NAND U640 ( .A(b[364]), .B(a[364]), .Z(n729) );
  NAND U641 ( .A(b[363]), .B(a[363]), .Z(n727) );
  NAND U642 ( .A(b[362]), .B(a[362]), .Z(n725) );
  NAND U643 ( .A(b[361]), .B(a[361]), .Z(n723) );
  NAND U644 ( .A(b[360]), .B(a[360]), .Z(n721) );
  NAND U645 ( .A(b[359]), .B(a[359]), .Z(n719) );
  NAND U646 ( .A(b[358]), .B(a[358]), .Z(n717) );
  NAND U647 ( .A(b[357]), .B(a[357]), .Z(n715) );
  NAND U648 ( .A(b[356]), .B(a[356]), .Z(n713) );
  NAND U649 ( .A(b[355]), .B(a[355]), .Z(n711) );
  NAND U650 ( .A(b[354]), .B(a[354]), .Z(n709) );
  NAND U651 ( .A(b[353]), .B(a[353]), .Z(n707) );
  NAND U652 ( .A(b[352]), .B(a[352]), .Z(n705) );
  NAND U653 ( .A(b[351]), .B(a[351]), .Z(n703) );
  NAND U654 ( .A(b[350]), .B(a[350]), .Z(n701) );
  NAND U655 ( .A(b[349]), .B(a[349]), .Z(n699) );
  NAND U656 ( .A(b[348]), .B(a[348]), .Z(n697) );
  NAND U657 ( .A(b[347]), .B(a[347]), .Z(n695) );
  NAND U658 ( .A(b[346]), .B(a[346]), .Z(n693) );
  NAND U659 ( .A(b[345]), .B(a[345]), .Z(n691) );
  NAND U660 ( .A(b[344]), .B(a[344]), .Z(n689) );
  NAND U661 ( .A(b[343]), .B(a[343]), .Z(n687) );
  NAND U662 ( .A(b[342]), .B(a[342]), .Z(n685) );
  NAND U663 ( .A(b[341]), .B(a[341]), .Z(n683) );
  NAND U664 ( .A(b[340]), .B(a[340]), .Z(n681) );
  NAND U665 ( .A(b[339]), .B(a[339]), .Z(n679) );
  NAND U666 ( .A(b[338]), .B(a[338]), .Z(n677) );
  NAND U667 ( .A(b[337]), .B(a[337]), .Z(n675) );
  NAND U668 ( .A(b[336]), .B(a[336]), .Z(n673) );
  NAND U669 ( .A(b[335]), .B(a[335]), .Z(n671) );
  NAND U670 ( .A(b[334]), .B(a[334]), .Z(n669) );
  NAND U671 ( .A(b[333]), .B(a[333]), .Z(n667) );
  NAND U672 ( .A(b[332]), .B(a[332]), .Z(n665) );
  NAND U673 ( .A(b[331]), .B(a[331]), .Z(n663) );
  NAND U674 ( .A(b[330]), .B(a[330]), .Z(n661) );
  NAND U675 ( .A(b[329]), .B(a[329]), .Z(n659) );
  NAND U676 ( .A(b[328]), .B(a[328]), .Z(n657) );
  NAND U677 ( .A(b[327]), .B(a[327]), .Z(n655) );
  NAND U678 ( .A(b[326]), .B(a[326]), .Z(n653) );
  NAND U679 ( .A(b[325]), .B(a[325]), .Z(n651) );
  NAND U680 ( .A(b[324]), .B(a[324]), .Z(n649) );
  NAND U681 ( .A(b[323]), .B(a[323]), .Z(n647) );
  NAND U682 ( .A(b[322]), .B(a[322]), .Z(n645) );
  NAND U683 ( .A(b[321]), .B(a[321]), .Z(n643) );
  NAND U684 ( .A(b[320]), .B(a[320]), .Z(n641) );
  NAND U685 ( .A(b[319]), .B(a[319]), .Z(n639) );
  NAND U686 ( .A(b[318]), .B(a[318]), .Z(n637) );
  NAND U687 ( .A(b[317]), .B(a[317]), .Z(n635) );
  NAND U688 ( .A(b[316]), .B(a[316]), .Z(n633) );
  NAND U689 ( .A(b[315]), .B(a[315]), .Z(n631) );
  NAND U690 ( .A(b[314]), .B(a[314]), .Z(n629) );
  NAND U691 ( .A(b[313]), .B(a[313]), .Z(n627) );
  NAND U692 ( .A(b[312]), .B(a[312]), .Z(n625) );
  NAND U693 ( .A(b[311]), .B(a[311]), .Z(n623) );
  NAND U694 ( .A(b[310]), .B(a[310]), .Z(n621) );
  NAND U695 ( .A(b[309]), .B(a[309]), .Z(n619) );
  NAND U696 ( .A(b[308]), .B(a[308]), .Z(n617) );
  NAND U697 ( .A(b[307]), .B(a[307]), .Z(n615) );
  NAND U698 ( .A(b[306]), .B(a[306]), .Z(n613) );
  NAND U699 ( .A(b[305]), .B(a[305]), .Z(n611) );
  NAND U700 ( .A(b[304]), .B(a[304]), .Z(n609) );
  NAND U701 ( .A(b[303]), .B(a[303]), .Z(n607) );
  NAND U702 ( .A(b[302]), .B(a[302]), .Z(n605) );
  NAND U703 ( .A(b[301]), .B(a[301]), .Z(n603) );
  NAND U704 ( .A(b[300]), .B(a[300]), .Z(n601) );
  NAND U705 ( .A(b[299]), .B(a[299]), .Z(n599) );
  NAND U706 ( .A(b[298]), .B(a[298]), .Z(n597) );
  NAND U707 ( .A(b[297]), .B(a[297]), .Z(n595) );
  NAND U708 ( .A(b[296]), .B(a[296]), .Z(n593) );
  NAND U709 ( .A(b[295]), .B(a[295]), .Z(n591) );
  NAND U710 ( .A(b[294]), .B(a[294]), .Z(n589) );
  NAND U711 ( .A(b[293]), .B(a[293]), .Z(n587) );
  NAND U712 ( .A(b[292]), .B(a[292]), .Z(n585) );
  NAND U713 ( .A(b[291]), .B(a[291]), .Z(n583) );
  NAND U714 ( .A(b[290]), .B(a[290]), .Z(n581) );
  NAND U715 ( .A(b[289]), .B(a[289]), .Z(n579) );
  NAND U716 ( .A(b[288]), .B(a[288]), .Z(n577) );
  NAND U717 ( .A(b[287]), .B(a[287]), .Z(n575) );
  NAND U718 ( .A(b[286]), .B(a[286]), .Z(n573) );
  NAND U719 ( .A(b[285]), .B(a[285]), .Z(n571) );
  NAND U720 ( .A(b[284]), .B(a[284]), .Z(n569) );
  NAND U721 ( .A(b[283]), .B(a[283]), .Z(n567) );
  NAND U722 ( .A(b[282]), .B(a[282]), .Z(n565) );
  NAND U723 ( .A(b[281]), .B(a[281]), .Z(n563) );
  NAND U724 ( .A(b[280]), .B(a[280]), .Z(n561) );
  NAND U725 ( .A(b[279]), .B(a[279]), .Z(n559) );
  NAND U726 ( .A(b[278]), .B(a[278]), .Z(n557) );
  NAND U727 ( .A(b[277]), .B(a[277]), .Z(n555) );
  NAND U728 ( .A(b[276]), .B(a[276]), .Z(n553) );
  NAND U729 ( .A(b[275]), .B(a[275]), .Z(n551) );
  NAND U730 ( .A(b[274]), .B(a[274]), .Z(n549) );
  NAND U731 ( .A(b[273]), .B(a[273]), .Z(n547) );
  NAND U732 ( .A(b[272]), .B(a[272]), .Z(n545) );
  NAND U733 ( .A(b[271]), .B(a[271]), .Z(n543) );
  NAND U734 ( .A(b[270]), .B(a[270]), .Z(n541) );
  NAND U735 ( .A(b[269]), .B(a[269]), .Z(n539) );
  NAND U736 ( .A(b[268]), .B(a[268]), .Z(n537) );
  NAND U737 ( .A(b[267]), .B(a[267]), .Z(n535) );
  NAND U738 ( .A(b[266]), .B(a[266]), .Z(n533) );
  NAND U739 ( .A(b[265]), .B(a[265]), .Z(n531) );
  NAND U740 ( .A(b[264]), .B(a[264]), .Z(n529) );
  NAND U741 ( .A(b[263]), .B(a[263]), .Z(n527) );
  NAND U742 ( .A(b[262]), .B(a[262]), .Z(n525) );
  NAND U743 ( .A(b[261]), .B(a[261]), .Z(n523) );
  NAND U744 ( .A(b[260]), .B(a[260]), .Z(n521) );
  NAND U745 ( .A(b[259]), .B(a[259]), .Z(n519) );
  NAND U746 ( .A(b[258]), .B(a[258]), .Z(n517) );
  NAND U747 ( .A(b[257]), .B(a[257]), .Z(n515) );
  NAND U748 ( .A(b[256]), .B(a[256]), .Z(n513) );
  NAND U749 ( .A(b[255]), .B(a[255]), .Z(n511) );
  NAND U750 ( .A(b[254]), .B(a[254]), .Z(n509) );
  NAND U751 ( .A(b[253]), .B(a[253]), .Z(n507) );
  NAND U752 ( .A(b[252]), .B(a[252]), .Z(n505) );
  NAND U753 ( .A(b[251]), .B(a[251]), .Z(n503) );
  NAND U754 ( .A(b[250]), .B(a[250]), .Z(n501) );
  NAND U755 ( .A(b[249]), .B(a[249]), .Z(n499) );
  NAND U756 ( .A(b[248]), .B(a[248]), .Z(n497) );
  NAND U757 ( .A(b[247]), .B(a[247]), .Z(n495) );
  NAND U758 ( .A(b[246]), .B(a[246]), .Z(n493) );
  NAND U759 ( .A(b[245]), .B(a[245]), .Z(n491) );
  NAND U760 ( .A(b[244]), .B(a[244]), .Z(n489) );
  NAND U761 ( .A(b[243]), .B(a[243]), .Z(n487) );
  NAND U762 ( .A(b[242]), .B(a[242]), .Z(n485) );
  NAND U763 ( .A(b[241]), .B(a[241]), .Z(n483) );
  NAND U764 ( .A(b[240]), .B(a[240]), .Z(n481) );
  NAND U765 ( .A(b[239]), .B(a[239]), .Z(n479) );
  NAND U766 ( .A(b[238]), .B(a[238]), .Z(n477) );
  NAND U767 ( .A(b[237]), .B(a[237]), .Z(n475) );
  NAND U768 ( .A(b[236]), .B(a[236]), .Z(n473) );
  NAND U769 ( .A(b[235]), .B(a[235]), .Z(n471) );
  NAND U770 ( .A(b[234]), .B(a[234]), .Z(n469) );
  NAND U771 ( .A(b[233]), .B(a[233]), .Z(n467) );
  NAND U772 ( .A(b[232]), .B(a[232]), .Z(n465) );
  NAND U773 ( .A(b[231]), .B(a[231]), .Z(n463) );
  NAND U774 ( .A(b[230]), .B(a[230]), .Z(n461) );
  NAND U775 ( .A(b[229]), .B(a[229]), .Z(n459) );
  NAND U776 ( .A(b[228]), .B(a[228]), .Z(n457) );
  NAND U777 ( .A(b[227]), .B(a[227]), .Z(n455) );
  NAND U778 ( .A(b[226]), .B(a[226]), .Z(n453) );
  NAND U779 ( .A(b[225]), .B(a[225]), .Z(n451) );
  NAND U780 ( .A(b[224]), .B(a[224]), .Z(n449) );
  NAND U781 ( .A(b[223]), .B(a[223]), .Z(n447) );
  NAND U782 ( .A(b[222]), .B(a[222]), .Z(n445) );
  NAND U783 ( .A(b[221]), .B(a[221]), .Z(n443) );
  NAND U784 ( .A(b[220]), .B(a[220]), .Z(n441) );
  NAND U785 ( .A(b[219]), .B(a[219]), .Z(n439) );
  NAND U786 ( .A(b[218]), .B(a[218]), .Z(n437) );
  NAND U787 ( .A(b[217]), .B(a[217]), .Z(n435) );
  NAND U788 ( .A(b[216]), .B(a[216]), .Z(n433) );
  NAND U789 ( .A(b[215]), .B(a[215]), .Z(n431) );
  NAND U790 ( .A(b[214]), .B(a[214]), .Z(n429) );
  NAND U791 ( .A(b[213]), .B(a[213]), .Z(n427) );
  NAND U792 ( .A(b[212]), .B(a[212]), .Z(n425) );
  NAND U793 ( .A(b[211]), .B(a[211]), .Z(n423) );
  NAND U794 ( .A(b[210]), .B(a[210]), .Z(n421) );
  NAND U795 ( .A(b[209]), .B(a[209]), .Z(n419) );
  NAND U796 ( .A(b[208]), .B(a[208]), .Z(n417) );
  NAND U797 ( .A(b[207]), .B(a[207]), .Z(n415) );
  NAND U798 ( .A(b[206]), .B(a[206]), .Z(n413) );
  NAND U799 ( .A(b[205]), .B(a[205]), .Z(n411) );
  NAND U800 ( .A(b[204]), .B(a[204]), .Z(n409) );
  NAND U801 ( .A(b[203]), .B(a[203]), .Z(n407) );
  NAND U802 ( .A(b[202]), .B(a[202]), .Z(n405) );
  NAND U803 ( .A(b[201]), .B(a[201]), .Z(n403) );
  NAND U804 ( .A(b[200]), .B(a[200]), .Z(n401) );
  NAND U805 ( .A(b[199]), .B(a[199]), .Z(n399) );
  NAND U806 ( .A(b[198]), .B(a[198]), .Z(n397) );
  NAND U807 ( .A(b[197]), .B(a[197]), .Z(n395) );
  NAND U808 ( .A(b[196]), .B(a[196]), .Z(n393) );
  NAND U809 ( .A(b[195]), .B(a[195]), .Z(n391) );
  NAND U810 ( .A(b[194]), .B(a[194]), .Z(n389) );
  NAND U811 ( .A(b[193]), .B(a[193]), .Z(n387) );
  NAND U812 ( .A(b[192]), .B(a[192]), .Z(n385) );
  NAND U813 ( .A(b[191]), .B(a[191]), .Z(n383) );
  NAND U814 ( .A(b[190]), .B(a[190]), .Z(n381) );
  NAND U815 ( .A(b[189]), .B(a[189]), .Z(n379) );
  NAND U816 ( .A(b[188]), .B(a[188]), .Z(n377) );
  NAND U817 ( .A(b[187]), .B(a[187]), .Z(n375) );
  NAND U818 ( .A(b[186]), .B(a[186]), .Z(n373) );
  NAND U819 ( .A(b[185]), .B(a[185]), .Z(n371) );
  NAND U820 ( .A(b[184]), .B(a[184]), .Z(n369) );
  NAND U821 ( .A(b[183]), .B(a[183]), .Z(n367) );
  NAND U822 ( .A(b[182]), .B(a[182]), .Z(n365) );
  NAND U823 ( .A(b[181]), .B(a[181]), .Z(n363) );
  NAND U824 ( .A(b[180]), .B(a[180]), .Z(n361) );
  NAND U825 ( .A(b[179]), .B(a[179]), .Z(n359) );
  NAND U826 ( .A(b[178]), .B(a[178]), .Z(n357) );
  NAND U827 ( .A(b[177]), .B(a[177]), .Z(n355) );
  NAND U828 ( .A(b[176]), .B(a[176]), .Z(n353) );
  NAND U829 ( .A(b[175]), .B(a[175]), .Z(n351) );
  NAND U830 ( .A(b[174]), .B(a[174]), .Z(n349) );
  NAND U831 ( .A(b[173]), .B(a[173]), .Z(n347) );
  NAND U832 ( .A(b[172]), .B(a[172]), .Z(n345) );
  NAND U833 ( .A(b[171]), .B(a[171]), .Z(n343) );
  NAND U834 ( .A(b[170]), .B(a[170]), .Z(n341) );
  NAND U835 ( .A(b[169]), .B(a[169]), .Z(n339) );
  NAND U836 ( .A(b[168]), .B(a[168]), .Z(n337) );
  NAND U837 ( .A(b[167]), .B(a[167]), .Z(n335) );
  NAND U838 ( .A(b[166]), .B(a[166]), .Z(n333) );
  NAND U839 ( .A(b[165]), .B(a[165]), .Z(n331) );
  NAND U840 ( .A(b[164]), .B(a[164]), .Z(n329) );
  NAND U841 ( .A(b[163]), .B(a[163]), .Z(n327) );
  NAND U842 ( .A(b[162]), .B(a[162]), .Z(n325) );
  NAND U843 ( .A(b[161]), .B(a[161]), .Z(n323) );
  NAND U844 ( .A(b[160]), .B(a[160]), .Z(n321) );
  NAND U845 ( .A(b[159]), .B(a[159]), .Z(n319) );
  NAND U846 ( .A(b[158]), .B(a[158]), .Z(n317) );
  NAND U847 ( .A(b[157]), .B(a[157]), .Z(n315) );
  NAND U848 ( .A(b[156]), .B(a[156]), .Z(n313) );
  NAND U849 ( .A(b[155]), .B(a[155]), .Z(n311) );
  NAND U850 ( .A(b[154]), .B(a[154]), .Z(n309) );
  NAND U851 ( .A(b[153]), .B(a[153]), .Z(n307) );
  NAND U852 ( .A(b[152]), .B(a[152]), .Z(n305) );
  NAND U853 ( .A(b[151]), .B(a[151]), .Z(n303) );
  NAND U854 ( .A(b[150]), .B(a[150]), .Z(n301) );
  NAND U855 ( .A(b[149]), .B(a[149]), .Z(n299) );
  NAND U856 ( .A(b[148]), .B(a[148]), .Z(n297) );
  NAND U857 ( .A(b[147]), .B(a[147]), .Z(n295) );
  NAND U858 ( .A(b[146]), .B(a[146]), .Z(n293) );
  NAND U859 ( .A(b[145]), .B(a[145]), .Z(n291) );
  NAND U860 ( .A(b[144]), .B(a[144]), .Z(n289) );
  NAND U861 ( .A(b[143]), .B(a[143]), .Z(n287) );
  NAND U862 ( .A(b[142]), .B(a[142]), .Z(n285) );
  NAND U863 ( .A(b[141]), .B(a[141]), .Z(n283) );
  NAND U864 ( .A(b[140]), .B(a[140]), .Z(n281) );
  NAND U865 ( .A(b[139]), .B(a[139]), .Z(n279) );
  NAND U866 ( .A(b[138]), .B(a[138]), .Z(n277) );
  NAND U867 ( .A(b[137]), .B(a[137]), .Z(n275) );
  NAND U868 ( .A(b[136]), .B(a[136]), .Z(n273) );
  NAND U869 ( .A(b[135]), .B(a[135]), .Z(n271) );
  NAND U870 ( .A(b[134]), .B(a[134]), .Z(n269) );
  NAND U871 ( .A(b[133]), .B(a[133]), .Z(n267) );
  NAND U872 ( .A(b[132]), .B(a[132]), .Z(n265) );
  NAND U873 ( .A(b[131]), .B(a[131]), .Z(n263) );
  NAND U874 ( .A(b[130]), .B(a[130]), .Z(n261) );
  NAND U875 ( .A(b[129]), .B(a[129]), .Z(n259) );
  NAND U876 ( .A(b[128]), .B(a[128]), .Z(n257) );
  NAND U877 ( .A(b[127]), .B(a[127]), .Z(n255) );
  NAND U878 ( .A(b[126]), .B(a[126]), .Z(n253) );
  NAND U879 ( .A(b[125]), .B(a[125]), .Z(n251) );
  NAND U880 ( .A(b[124]), .B(a[124]), .Z(n249) );
  NAND U881 ( .A(b[123]), .B(a[123]), .Z(n247) );
  NAND U882 ( .A(b[122]), .B(a[122]), .Z(n245) );
  NAND U883 ( .A(b[121]), .B(a[121]), .Z(n243) );
  NAND U884 ( .A(b[120]), .B(a[120]), .Z(n241) );
  NAND U885 ( .A(b[119]), .B(a[119]), .Z(n239) );
  NAND U886 ( .A(b[118]), .B(a[118]), .Z(n237) );
  NAND U887 ( .A(b[117]), .B(a[117]), .Z(n235) );
  NAND U888 ( .A(b[116]), .B(a[116]), .Z(n233) );
  NAND U889 ( .A(b[115]), .B(a[115]), .Z(n231) );
  NAND U890 ( .A(b[114]), .B(a[114]), .Z(n229) );
  NAND U891 ( .A(b[113]), .B(a[113]), .Z(n227) );
  NAND U892 ( .A(b[112]), .B(a[112]), .Z(n225) );
  NAND U893 ( .A(b[111]), .B(a[111]), .Z(n223) );
  NAND U894 ( .A(b[110]), .B(a[110]), .Z(n221) );
  NAND U895 ( .A(b[109]), .B(a[109]), .Z(n219) );
  NAND U896 ( .A(b[108]), .B(a[108]), .Z(n217) );
  NAND U897 ( .A(b[107]), .B(a[107]), .Z(n215) );
  NAND U898 ( .A(b[106]), .B(a[106]), .Z(n213) );
  NAND U899 ( .A(b[105]), .B(a[105]), .Z(n211) );
  NAND U900 ( .A(b[104]), .B(a[104]), .Z(n209) );
  NAND U901 ( .A(b[103]), .B(a[103]), .Z(n207) );
  NAND U902 ( .A(b[102]), .B(a[102]), .Z(n205) );
  NAND U903 ( .A(b[101]), .B(a[101]), .Z(n203) );
  NAND U904 ( .A(b[100]), .B(a[100]), .Z(n201) );
  NAND U905 ( .A(b[99]), .B(a[99]), .Z(n199) );
  XNOR U906 ( .A(b[99]), .B(a[99]), .Z(n4089) );
  NAND U907 ( .A(b[98]), .B(a[98]), .Z(n197) );
  NAND U908 ( .A(b[97]), .B(a[97]), .Z(n195) );
  NAND U909 ( .A(b[96]), .B(a[96]), .Z(n193) );
  NAND U910 ( .A(b[95]), .B(a[95]), .Z(n191) );
  NAND U911 ( .A(b[94]), .B(a[94]), .Z(n189) );
  NAND U912 ( .A(b[93]), .B(a[93]), .Z(n187) );
  NAND U913 ( .A(b[92]), .B(a[92]), .Z(n185) );
  NAND U914 ( .A(b[91]), .B(a[91]), .Z(n183) );
  NAND U915 ( .A(b[90]), .B(a[90]), .Z(n181) );
  NAND U916 ( .A(b[89]), .B(a[89]), .Z(n179) );
  NAND U917 ( .A(b[88]), .B(a[88]), .Z(n177) );
  NAND U918 ( .A(b[87]), .B(a[87]), .Z(n175) );
  NAND U919 ( .A(b[86]), .B(a[86]), .Z(n173) );
  NAND U920 ( .A(b[85]), .B(a[85]), .Z(n171) );
  NAND U921 ( .A(b[84]), .B(a[84]), .Z(n169) );
  NAND U922 ( .A(b[83]), .B(a[83]), .Z(n167) );
  NAND U923 ( .A(b[82]), .B(a[82]), .Z(n165) );
  NAND U924 ( .A(b[81]), .B(a[81]), .Z(n163) );
  NAND U925 ( .A(b[80]), .B(a[80]), .Z(n161) );
  NAND U926 ( .A(b[79]), .B(a[79]), .Z(n159) );
  NAND U927 ( .A(b[78]), .B(a[78]), .Z(n157) );
  NAND U928 ( .A(b[77]), .B(a[77]), .Z(n155) );
  NAND U929 ( .A(b[76]), .B(a[76]), .Z(n153) );
  NAND U930 ( .A(b[75]), .B(a[75]), .Z(n151) );
  NAND U931 ( .A(b[74]), .B(a[74]), .Z(n149) );
  NAND U932 ( .A(b[73]), .B(a[73]), .Z(n147) );
  NAND U933 ( .A(b[72]), .B(a[72]), .Z(n145) );
  NAND U934 ( .A(b[71]), .B(a[71]), .Z(n143) );
  NAND U935 ( .A(b[70]), .B(a[70]), .Z(n141) );
  NAND U936 ( .A(b[69]), .B(a[69]), .Z(n139) );
  NAND U937 ( .A(b[68]), .B(a[68]), .Z(n137) );
  NAND U938 ( .A(b[67]), .B(a[67]), .Z(n135) );
  NAND U939 ( .A(b[66]), .B(a[66]), .Z(n133) );
  NAND U940 ( .A(b[65]), .B(a[65]), .Z(n131) );
  NAND U941 ( .A(b[64]), .B(a[64]), .Z(n129) );
  NAND U942 ( .A(b[63]), .B(a[63]), .Z(n127) );
  NAND U943 ( .A(b[62]), .B(a[62]), .Z(n125) );
  NAND U944 ( .A(b[61]), .B(a[61]), .Z(n123) );
  NAND U945 ( .A(b[60]), .B(a[60]), .Z(n121) );
  NAND U946 ( .A(b[59]), .B(a[59]), .Z(n119) );
  NAND U947 ( .A(b[58]), .B(a[58]), .Z(n117) );
  NAND U948 ( .A(b[57]), .B(a[57]), .Z(n115) );
  NAND U949 ( .A(b[56]), .B(a[56]), .Z(n113) );
  NAND U950 ( .A(b[55]), .B(a[55]), .Z(n111) );
  NAND U951 ( .A(b[54]), .B(a[54]), .Z(n109) );
  NAND U952 ( .A(b[53]), .B(a[53]), .Z(n107) );
  NAND U953 ( .A(b[52]), .B(a[52]), .Z(n105) );
  NAND U954 ( .A(b[51]), .B(a[51]), .Z(n103) );
  NAND U955 ( .A(b[50]), .B(a[50]), .Z(n101) );
  NAND U956 ( .A(b[49]), .B(a[49]), .Z(n99) );
  NAND U957 ( .A(b[48]), .B(a[48]), .Z(n97) );
  NAND U958 ( .A(b[47]), .B(a[47]), .Z(n95) );
  NAND U959 ( .A(b[46]), .B(a[46]), .Z(n93) );
  NAND U960 ( .A(b[45]), .B(a[45]), .Z(n91) );
  NAND U961 ( .A(b[44]), .B(a[44]), .Z(n89) );
  NAND U962 ( .A(b[43]), .B(a[43]), .Z(n87) );
  NAND U963 ( .A(b[42]), .B(a[42]), .Z(n85) );
  NAND U964 ( .A(b[41]), .B(a[41]), .Z(n83) );
  NAND U965 ( .A(b[40]), .B(a[40]), .Z(n81) );
  NAND U966 ( .A(b[39]), .B(a[39]), .Z(n79) );
  NAND U967 ( .A(b[38]), .B(a[38]), .Z(n77) );
  NAND U968 ( .A(b[37]), .B(a[37]), .Z(n75) );
  NAND U969 ( .A(b[36]), .B(a[36]), .Z(n73) );
  NAND U970 ( .A(b[35]), .B(a[35]), .Z(n71) );
  NAND U971 ( .A(b[34]), .B(a[34]), .Z(n69) );
  NAND U972 ( .A(b[33]), .B(a[33]), .Z(n67) );
  NAND U973 ( .A(b[32]), .B(a[32]), .Z(n65) );
  NAND U974 ( .A(b[31]), .B(a[31]), .Z(n63) );
  NAND U975 ( .A(b[30]), .B(a[30]), .Z(n61) );
  NAND U976 ( .A(b[29]), .B(a[29]), .Z(n59) );
  NAND U977 ( .A(b[28]), .B(a[28]), .Z(n57) );
  NAND U978 ( .A(b[27]), .B(a[27]), .Z(n55) );
  NAND U979 ( .A(b[26]), .B(a[26]), .Z(n53) );
  NAND U980 ( .A(b[25]), .B(a[25]), .Z(n51) );
  NAND U981 ( .A(b[24]), .B(a[24]), .Z(n49) );
  NAND U982 ( .A(b[23]), .B(a[23]), .Z(n47) );
  NAND U983 ( .A(b[22]), .B(a[22]), .Z(n45) );
  NAND U984 ( .A(b[21]), .B(a[21]), .Z(n43) );
  NAND U985 ( .A(b[20]), .B(a[20]), .Z(n41) );
  NAND U986 ( .A(b[19]), .B(a[19]), .Z(n39) );
  NAND U987 ( .A(b[18]), .B(a[18]), .Z(n37) );
  NAND U988 ( .A(b[17]), .B(a[17]), .Z(n35) );
  NAND U989 ( .A(b[16]), .B(a[16]), .Z(n33) );
  NAND U990 ( .A(b[15]), .B(a[15]), .Z(n31) );
  NAND U991 ( .A(b[14]), .B(a[14]), .Z(n29) );
  NAND U992 ( .A(b[13]), .B(a[13]), .Z(n27) );
  NAND U993 ( .A(b[12]), .B(a[12]), .Z(n25) );
  NAND U994 ( .A(b[11]), .B(a[11]), .Z(n23) );
  NAND U995 ( .A(b[10]), .B(a[10]), .Z(n21) );
  NAND U996 ( .A(b[9]), .B(a[9]), .Z(n19) );
  XNOR U997 ( .A(b[9]), .B(a[9]), .Z(n4091) );
  NAND U998 ( .A(b[8]), .B(a[8]), .Z(n17) );
  NAND U999 ( .A(b[7]), .B(a[7]), .Z(n15) );
  NAND U1000 ( .A(b[6]), .B(a[6]), .Z(n13) );
  NAND U1001 ( .A(b[5]), .B(a[5]), .Z(n11) );
  NAND U1002 ( .A(b[4]), .B(a[4]), .Z(n9) );
  NAND U1003 ( .A(b[3]), .B(a[3]), .Z(n7) );
  NAND U1004 ( .A(b[2]), .B(a[2]), .Z(n5) );
  NAND U1005 ( .A(b[1]), .B(a[1]), .Z(n3) );
  NAND U1006 ( .A(a[0]), .B(b[0]), .Z(n2314) );
  XOR U1007 ( .A(a[1]), .B(b[1]), .Z(n2315) );
  NANDN U1008 ( .A(n2314), .B(n2315), .Z(n2) );
  AND U1009 ( .A(n3), .B(n2), .Z(n2536) );
  XOR U1010 ( .A(a[2]), .B(b[2]), .Z(n2537) );
  NANDN U1011 ( .A(n2536), .B(n2537), .Z(n4) );
  AND U1012 ( .A(n5), .B(n4), .Z(n2758) );
  XOR U1013 ( .A(a[3]), .B(b[3]), .Z(n2759) );
  NANDN U1014 ( .A(n2758), .B(n2759), .Z(n6) );
  AND U1015 ( .A(n7), .B(n6), .Z(n2980) );
  XOR U1016 ( .A(a[4]), .B(b[4]), .Z(n2981) );
  NANDN U1017 ( .A(n2980), .B(n2981), .Z(n8) );
  AND U1018 ( .A(n9), .B(n8), .Z(n3202) );
  XOR U1019 ( .A(a[5]), .B(b[5]), .Z(n3203) );
  NANDN U1020 ( .A(n3202), .B(n3203), .Z(n10) );
  AND U1021 ( .A(n11), .B(n10), .Z(n3424) );
  XOR U1022 ( .A(a[6]), .B(b[6]), .Z(n3425) );
  NANDN U1023 ( .A(n3424), .B(n3425), .Z(n12) );
  AND U1024 ( .A(n13), .B(n12), .Z(n3646) );
  XOR U1025 ( .A(a[7]), .B(b[7]), .Z(n3647) );
  NANDN U1026 ( .A(n3646), .B(n3647), .Z(n14) );
  AND U1027 ( .A(n15), .B(n14), .Z(n3868) );
  XOR U1028 ( .A(a[8]), .B(b[8]), .Z(n3869) );
  NANDN U1029 ( .A(n3868), .B(n3869), .Z(n16) );
  AND U1030 ( .A(n17), .B(n16), .Z(n4090) );
  OR U1031 ( .A(n4091), .B(n4090), .Z(n18) );
  AND U1032 ( .A(n19), .B(n18), .Z(n2114) );
  XOR U1033 ( .A(a[10]), .B(b[10]), .Z(n2115) );
  NANDN U1034 ( .A(n2114), .B(n2115), .Z(n20) );
  AND U1035 ( .A(n21), .B(n20), .Z(n2136) );
  XOR U1036 ( .A(a[11]), .B(b[11]), .Z(n2137) );
  NANDN U1037 ( .A(n2136), .B(n2137), .Z(n22) );
  AND U1038 ( .A(n23), .B(n22), .Z(n2158) );
  XOR U1039 ( .A(a[12]), .B(b[12]), .Z(n2159) );
  NANDN U1040 ( .A(n2158), .B(n2159), .Z(n24) );
  AND U1041 ( .A(n25), .B(n24), .Z(n2180) );
  XOR U1042 ( .A(a[13]), .B(b[13]), .Z(n2181) );
  NANDN U1043 ( .A(n2180), .B(n2181), .Z(n26) );
  AND U1044 ( .A(n27), .B(n26), .Z(n2202) );
  XOR U1045 ( .A(a[14]), .B(b[14]), .Z(n2203) );
  NANDN U1046 ( .A(n2202), .B(n2203), .Z(n28) );
  AND U1047 ( .A(n29), .B(n28), .Z(n2224) );
  XOR U1048 ( .A(a[15]), .B(b[15]), .Z(n2225) );
  NANDN U1049 ( .A(n2224), .B(n2225), .Z(n30) );
  AND U1050 ( .A(n31), .B(n30), .Z(n2246) );
  XOR U1051 ( .A(a[16]), .B(b[16]), .Z(n2247) );
  NANDN U1052 ( .A(n2246), .B(n2247), .Z(n32) );
  AND U1053 ( .A(n33), .B(n32), .Z(n2268) );
  XOR U1054 ( .A(a[17]), .B(b[17]), .Z(n2269) );
  NANDN U1055 ( .A(n2268), .B(n2269), .Z(n34) );
  AND U1056 ( .A(n35), .B(n34), .Z(n2290) );
  XOR U1057 ( .A(a[18]), .B(b[18]), .Z(n2291) );
  NANDN U1058 ( .A(n2290), .B(n2291), .Z(n36) );
  AND U1059 ( .A(n37), .B(n36), .Z(n2312) );
  XOR U1060 ( .A(a[19]), .B(b[19]), .Z(n2313) );
  NANDN U1061 ( .A(n2312), .B(n2313), .Z(n38) );
  AND U1062 ( .A(n39), .B(n38), .Z(n2336) );
  XOR U1063 ( .A(a[20]), .B(b[20]), .Z(n2337) );
  NANDN U1064 ( .A(n2336), .B(n2337), .Z(n40) );
  AND U1065 ( .A(n41), .B(n40), .Z(n2358) );
  XOR U1066 ( .A(a[21]), .B(b[21]), .Z(n2359) );
  NANDN U1067 ( .A(n2358), .B(n2359), .Z(n42) );
  AND U1068 ( .A(n43), .B(n42), .Z(n2380) );
  XOR U1069 ( .A(a[22]), .B(b[22]), .Z(n2381) );
  NANDN U1070 ( .A(n2380), .B(n2381), .Z(n44) );
  AND U1071 ( .A(n45), .B(n44), .Z(n2402) );
  XOR U1072 ( .A(a[23]), .B(b[23]), .Z(n2403) );
  NANDN U1073 ( .A(n2402), .B(n2403), .Z(n46) );
  AND U1074 ( .A(n47), .B(n46), .Z(n2424) );
  XOR U1075 ( .A(a[24]), .B(b[24]), .Z(n2425) );
  NANDN U1076 ( .A(n2424), .B(n2425), .Z(n48) );
  AND U1077 ( .A(n49), .B(n48), .Z(n2446) );
  XOR U1078 ( .A(a[25]), .B(b[25]), .Z(n2447) );
  NANDN U1079 ( .A(n2446), .B(n2447), .Z(n50) );
  AND U1080 ( .A(n51), .B(n50), .Z(n2468) );
  XOR U1081 ( .A(a[26]), .B(b[26]), .Z(n2469) );
  NANDN U1082 ( .A(n2468), .B(n2469), .Z(n52) );
  AND U1083 ( .A(n53), .B(n52), .Z(n2490) );
  XOR U1084 ( .A(a[27]), .B(b[27]), .Z(n2491) );
  NANDN U1085 ( .A(n2490), .B(n2491), .Z(n54) );
  AND U1086 ( .A(n55), .B(n54), .Z(n2512) );
  XOR U1087 ( .A(a[28]), .B(b[28]), .Z(n2513) );
  NANDN U1088 ( .A(n2512), .B(n2513), .Z(n56) );
  AND U1089 ( .A(n57), .B(n56), .Z(n2534) );
  XOR U1090 ( .A(a[29]), .B(b[29]), .Z(n2535) );
  NANDN U1091 ( .A(n2534), .B(n2535), .Z(n58) );
  AND U1092 ( .A(n59), .B(n58), .Z(n2558) );
  XOR U1093 ( .A(a[30]), .B(b[30]), .Z(n2559) );
  NANDN U1094 ( .A(n2558), .B(n2559), .Z(n60) );
  AND U1095 ( .A(n61), .B(n60), .Z(n2580) );
  XOR U1096 ( .A(a[31]), .B(b[31]), .Z(n2581) );
  NANDN U1097 ( .A(n2580), .B(n2581), .Z(n62) );
  AND U1098 ( .A(n63), .B(n62), .Z(n2602) );
  XOR U1099 ( .A(a[32]), .B(b[32]), .Z(n2603) );
  NANDN U1100 ( .A(n2602), .B(n2603), .Z(n64) );
  AND U1101 ( .A(n65), .B(n64), .Z(n2624) );
  XOR U1102 ( .A(a[33]), .B(b[33]), .Z(n2625) );
  NANDN U1103 ( .A(n2624), .B(n2625), .Z(n66) );
  AND U1104 ( .A(n67), .B(n66), .Z(n2646) );
  XOR U1105 ( .A(a[34]), .B(b[34]), .Z(n2647) );
  NANDN U1106 ( .A(n2646), .B(n2647), .Z(n68) );
  AND U1107 ( .A(n69), .B(n68), .Z(n2668) );
  XOR U1108 ( .A(a[35]), .B(b[35]), .Z(n2669) );
  NANDN U1109 ( .A(n2668), .B(n2669), .Z(n70) );
  AND U1110 ( .A(n71), .B(n70), .Z(n2690) );
  XOR U1111 ( .A(a[36]), .B(b[36]), .Z(n2691) );
  NANDN U1112 ( .A(n2690), .B(n2691), .Z(n72) );
  AND U1113 ( .A(n73), .B(n72), .Z(n2712) );
  XOR U1114 ( .A(a[37]), .B(b[37]), .Z(n2713) );
  NANDN U1115 ( .A(n2712), .B(n2713), .Z(n74) );
  AND U1116 ( .A(n75), .B(n74), .Z(n2734) );
  XOR U1117 ( .A(a[38]), .B(b[38]), .Z(n2735) );
  NANDN U1118 ( .A(n2734), .B(n2735), .Z(n76) );
  AND U1119 ( .A(n77), .B(n76), .Z(n2756) );
  XOR U1120 ( .A(a[39]), .B(b[39]), .Z(n2757) );
  NANDN U1121 ( .A(n2756), .B(n2757), .Z(n78) );
  AND U1122 ( .A(n79), .B(n78), .Z(n2780) );
  XOR U1123 ( .A(a[40]), .B(b[40]), .Z(n2781) );
  NANDN U1124 ( .A(n2780), .B(n2781), .Z(n80) );
  AND U1125 ( .A(n81), .B(n80), .Z(n2802) );
  XOR U1126 ( .A(a[41]), .B(b[41]), .Z(n2803) );
  NANDN U1127 ( .A(n2802), .B(n2803), .Z(n82) );
  AND U1128 ( .A(n83), .B(n82), .Z(n2824) );
  XOR U1129 ( .A(a[42]), .B(b[42]), .Z(n2825) );
  NANDN U1130 ( .A(n2824), .B(n2825), .Z(n84) );
  AND U1131 ( .A(n85), .B(n84), .Z(n2846) );
  XOR U1132 ( .A(a[43]), .B(b[43]), .Z(n2847) );
  NANDN U1133 ( .A(n2846), .B(n2847), .Z(n86) );
  AND U1134 ( .A(n87), .B(n86), .Z(n2868) );
  XOR U1135 ( .A(a[44]), .B(b[44]), .Z(n2869) );
  NANDN U1136 ( .A(n2868), .B(n2869), .Z(n88) );
  AND U1137 ( .A(n89), .B(n88), .Z(n2890) );
  XOR U1138 ( .A(a[45]), .B(b[45]), .Z(n2891) );
  NANDN U1139 ( .A(n2890), .B(n2891), .Z(n90) );
  AND U1140 ( .A(n91), .B(n90), .Z(n2912) );
  XOR U1141 ( .A(a[46]), .B(b[46]), .Z(n2913) );
  NANDN U1142 ( .A(n2912), .B(n2913), .Z(n92) );
  AND U1143 ( .A(n93), .B(n92), .Z(n2934) );
  XOR U1144 ( .A(a[47]), .B(b[47]), .Z(n2935) );
  NANDN U1145 ( .A(n2934), .B(n2935), .Z(n94) );
  AND U1146 ( .A(n95), .B(n94), .Z(n2956) );
  XOR U1147 ( .A(a[48]), .B(b[48]), .Z(n2957) );
  NANDN U1148 ( .A(n2956), .B(n2957), .Z(n96) );
  AND U1149 ( .A(n97), .B(n96), .Z(n2978) );
  XOR U1150 ( .A(a[49]), .B(b[49]), .Z(n2979) );
  NANDN U1151 ( .A(n2978), .B(n2979), .Z(n98) );
  AND U1152 ( .A(n99), .B(n98), .Z(n3002) );
  XOR U1153 ( .A(a[50]), .B(b[50]), .Z(n3003) );
  NANDN U1154 ( .A(n3002), .B(n3003), .Z(n100) );
  AND U1155 ( .A(n101), .B(n100), .Z(n3024) );
  XOR U1156 ( .A(a[51]), .B(b[51]), .Z(n3025) );
  NANDN U1157 ( .A(n3024), .B(n3025), .Z(n102) );
  AND U1158 ( .A(n103), .B(n102), .Z(n3046) );
  XOR U1159 ( .A(a[52]), .B(b[52]), .Z(n3047) );
  NANDN U1160 ( .A(n3046), .B(n3047), .Z(n104) );
  AND U1161 ( .A(n105), .B(n104), .Z(n3068) );
  XOR U1162 ( .A(a[53]), .B(b[53]), .Z(n3069) );
  NANDN U1163 ( .A(n3068), .B(n3069), .Z(n106) );
  AND U1164 ( .A(n107), .B(n106), .Z(n3090) );
  XOR U1165 ( .A(a[54]), .B(b[54]), .Z(n3091) );
  NANDN U1166 ( .A(n3090), .B(n3091), .Z(n108) );
  AND U1167 ( .A(n109), .B(n108), .Z(n3112) );
  XOR U1168 ( .A(a[55]), .B(b[55]), .Z(n3113) );
  NANDN U1169 ( .A(n3112), .B(n3113), .Z(n110) );
  AND U1170 ( .A(n111), .B(n110), .Z(n3134) );
  XOR U1171 ( .A(a[56]), .B(b[56]), .Z(n3135) );
  NANDN U1172 ( .A(n3134), .B(n3135), .Z(n112) );
  AND U1173 ( .A(n113), .B(n112), .Z(n3156) );
  XOR U1174 ( .A(a[57]), .B(b[57]), .Z(n3157) );
  NANDN U1175 ( .A(n3156), .B(n3157), .Z(n114) );
  AND U1176 ( .A(n115), .B(n114), .Z(n3178) );
  XOR U1177 ( .A(a[58]), .B(b[58]), .Z(n3179) );
  NANDN U1178 ( .A(n3178), .B(n3179), .Z(n116) );
  AND U1179 ( .A(n117), .B(n116), .Z(n3200) );
  XOR U1180 ( .A(a[59]), .B(b[59]), .Z(n3201) );
  NANDN U1181 ( .A(n3200), .B(n3201), .Z(n118) );
  AND U1182 ( .A(n119), .B(n118), .Z(n3224) );
  XOR U1183 ( .A(a[60]), .B(b[60]), .Z(n3225) );
  NANDN U1184 ( .A(n3224), .B(n3225), .Z(n120) );
  AND U1185 ( .A(n121), .B(n120), .Z(n3246) );
  XOR U1186 ( .A(a[61]), .B(b[61]), .Z(n3247) );
  NANDN U1187 ( .A(n3246), .B(n3247), .Z(n122) );
  AND U1188 ( .A(n123), .B(n122), .Z(n3268) );
  XOR U1189 ( .A(a[62]), .B(b[62]), .Z(n3269) );
  NANDN U1190 ( .A(n3268), .B(n3269), .Z(n124) );
  AND U1191 ( .A(n125), .B(n124), .Z(n3290) );
  XOR U1192 ( .A(a[63]), .B(b[63]), .Z(n3291) );
  NANDN U1193 ( .A(n3290), .B(n3291), .Z(n126) );
  AND U1194 ( .A(n127), .B(n126), .Z(n3312) );
  XOR U1195 ( .A(a[64]), .B(b[64]), .Z(n3313) );
  NANDN U1196 ( .A(n3312), .B(n3313), .Z(n128) );
  AND U1197 ( .A(n129), .B(n128), .Z(n3334) );
  XOR U1198 ( .A(a[65]), .B(b[65]), .Z(n3335) );
  NANDN U1199 ( .A(n3334), .B(n3335), .Z(n130) );
  AND U1200 ( .A(n131), .B(n130), .Z(n3356) );
  XOR U1201 ( .A(a[66]), .B(b[66]), .Z(n3357) );
  NANDN U1202 ( .A(n3356), .B(n3357), .Z(n132) );
  AND U1203 ( .A(n133), .B(n132), .Z(n3378) );
  XOR U1204 ( .A(a[67]), .B(b[67]), .Z(n3379) );
  NANDN U1205 ( .A(n3378), .B(n3379), .Z(n134) );
  AND U1206 ( .A(n135), .B(n134), .Z(n3400) );
  XOR U1207 ( .A(a[68]), .B(b[68]), .Z(n3401) );
  NANDN U1208 ( .A(n3400), .B(n3401), .Z(n136) );
  AND U1209 ( .A(n137), .B(n136), .Z(n3422) );
  XOR U1210 ( .A(a[69]), .B(b[69]), .Z(n3423) );
  NANDN U1211 ( .A(n3422), .B(n3423), .Z(n138) );
  AND U1212 ( .A(n139), .B(n138), .Z(n3446) );
  XOR U1213 ( .A(a[70]), .B(b[70]), .Z(n3447) );
  NANDN U1214 ( .A(n3446), .B(n3447), .Z(n140) );
  AND U1215 ( .A(n141), .B(n140), .Z(n3468) );
  XOR U1216 ( .A(a[71]), .B(b[71]), .Z(n3469) );
  NANDN U1217 ( .A(n3468), .B(n3469), .Z(n142) );
  AND U1218 ( .A(n143), .B(n142), .Z(n3490) );
  XOR U1219 ( .A(a[72]), .B(b[72]), .Z(n3491) );
  NANDN U1220 ( .A(n3490), .B(n3491), .Z(n144) );
  AND U1221 ( .A(n145), .B(n144), .Z(n3512) );
  XOR U1222 ( .A(a[73]), .B(b[73]), .Z(n3513) );
  NANDN U1223 ( .A(n3512), .B(n3513), .Z(n146) );
  AND U1224 ( .A(n147), .B(n146), .Z(n3534) );
  XOR U1225 ( .A(a[74]), .B(b[74]), .Z(n3535) );
  NANDN U1226 ( .A(n3534), .B(n3535), .Z(n148) );
  AND U1227 ( .A(n149), .B(n148), .Z(n3556) );
  XOR U1228 ( .A(a[75]), .B(b[75]), .Z(n3557) );
  NANDN U1229 ( .A(n3556), .B(n3557), .Z(n150) );
  AND U1230 ( .A(n151), .B(n150), .Z(n3578) );
  XOR U1231 ( .A(a[76]), .B(b[76]), .Z(n3579) );
  NANDN U1232 ( .A(n3578), .B(n3579), .Z(n152) );
  AND U1233 ( .A(n153), .B(n152), .Z(n3600) );
  XOR U1234 ( .A(a[77]), .B(b[77]), .Z(n3601) );
  NANDN U1235 ( .A(n3600), .B(n3601), .Z(n154) );
  AND U1236 ( .A(n155), .B(n154), .Z(n3622) );
  XOR U1237 ( .A(a[78]), .B(b[78]), .Z(n3623) );
  NANDN U1238 ( .A(n3622), .B(n3623), .Z(n156) );
  AND U1239 ( .A(n157), .B(n156), .Z(n3644) );
  XOR U1240 ( .A(a[79]), .B(b[79]), .Z(n3645) );
  NANDN U1241 ( .A(n3644), .B(n3645), .Z(n158) );
  AND U1242 ( .A(n159), .B(n158), .Z(n3668) );
  XOR U1243 ( .A(a[80]), .B(b[80]), .Z(n3669) );
  NANDN U1244 ( .A(n3668), .B(n3669), .Z(n160) );
  AND U1245 ( .A(n161), .B(n160), .Z(n3690) );
  XOR U1246 ( .A(a[81]), .B(b[81]), .Z(n3691) );
  NANDN U1247 ( .A(n3690), .B(n3691), .Z(n162) );
  AND U1248 ( .A(n163), .B(n162), .Z(n3712) );
  XOR U1249 ( .A(a[82]), .B(b[82]), .Z(n3713) );
  NANDN U1250 ( .A(n3712), .B(n3713), .Z(n164) );
  AND U1251 ( .A(n165), .B(n164), .Z(n3734) );
  XOR U1252 ( .A(a[83]), .B(b[83]), .Z(n3735) );
  NANDN U1253 ( .A(n3734), .B(n3735), .Z(n166) );
  AND U1254 ( .A(n167), .B(n166), .Z(n3756) );
  XOR U1255 ( .A(a[84]), .B(b[84]), .Z(n3757) );
  NANDN U1256 ( .A(n3756), .B(n3757), .Z(n168) );
  AND U1257 ( .A(n169), .B(n168), .Z(n3778) );
  XOR U1258 ( .A(a[85]), .B(b[85]), .Z(n3779) );
  NANDN U1259 ( .A(n3778), .B(n3779), .Z(n170) );
  AND U1260 ( .A(n171), .B(n170), .Z(n3800) );
  XOR U1261 ( .A(a[86]), .B(b[86]), .Z(n3801) );
  NANDN U1262 ( .A(n3800), .B(n3801), .Z(n172) );
  AND U1263 ( .A(n173), .B(n172), .Z(n3822) );
  XOR U1264 ( .A(a[87]), .B(b[87]), .Z(n3823) );
  NANDN U1265 ( .A(n3822), .B(n3823), .Z(n174) );
  AND U1266 ( .A(n175), .B(n174), .Z(n3844) );
  XOR U1267 ( .A(a[88]), .B(b[88]), .Z(n3845) );
  NANDN U1268 ( .A(n3844), .B(n3845), .Z(n176) );
  AND U1269 ( .A(n177), .B(n176), .Z(n3866) );
  XOR U1270 ( .A(a[89]), .B(b[89]), .Z(n3867) );
  NANDN U1271 ( .A(n3866), .B(n3867), .Z(n178) );
  AND U1272 ( .A(n179), .B(n178), .Z(n3890) );
  XOR U1273 ( .A(a[90]), .B(b[90]), .Z(n3891) );
  NANDN U1274 ( .A(n3890), .B(n3891), .Z(n180) );
  AND U1275 ( .A(n181), .B(n180), .Z(n3912) );
  XOR U1276 ( .A(a[91]), .B(b[91]), .Z(n3913) );
  NANDN U1277 ( .A(n3912), .B(n3913), .Z(n182) );
  AND U1278 ( .A(n183), .B(n182), .Z(n3934) );
  XOR U1279 ( .A(a[92]), .B(b[92]), .Z(n3935) );
  NANDN U1280 ( .A(n3934), .B(n3935), .Z(n184) );
  AND U1281 ( .A(n185), .B(n184), .Z(n3956) );
  XOR U1282 ( .A(a[93]), .B(b[93]), .Z(n3957) );
  NANDN U1283 ( .A(n3956), .B(n3957), .Z(n186) );
  AND U1284 ( .A(n187), .B(n186), .Z(n3978) );
  XOR U1285 ( .A(a[94]), .B(b[94]), .Z(n3979) );
  NANDN U1286 ( .A(n3978), .B(n3979), .Z(n188) );
  AND U1287 ( .A(n189), .B(n188), .Z(n4000) );
  XOR U1288 ( .A(a[95]), .B(b[95]), .Z(n4001) );
  NANDN U1289 ( .A(n4000), .B(n4001), .Z(n190) );
  AND U1290 ( .A(n191), .B(n190), .Z(n4022) );
  XOR U1291 ( .A(a[96]), .B(b[96]), .Z(n4023) );
  NANDN U1292 ( .A(n4022), .B(n4023), .Z(n192) );
  AND U1293 ( .A(n193), .B(n192), .Z(n4044) );
  XOR U1294 ( .A(a[97]), .B(b[97]), .Z(n4045) );
  NANDN U1295 ( .A(n4044), .B(n4045), .Z(n194) );
  AND U1296 ( .A(n195), .B(n194), .Z(n4066) );
  XOR U1297 ( .A(a[98]), .B(b[98]), .Z(n4067) );
  NANDN U1298 ( .A(n4066), .B(n4067), .Z(n196) );
  AND U1299 ( .A(n197), .B(n196), .Z(n4088) );
  OR U1300 ( .A(n4089), .B(n4088), .Z(n198) );
  AND U1301 ( .A(n199), .B(n198), .Z(n2036) );
  XOR U1302 ( .A(a[100]), .B(b[100]), .Z(n2037) );
  NANDN U1303 ( .A(n2036), .B(n2037), .Z(n200) );
  AND U1304 ( .A(n201), .B(n200), .Z(n2078) );
  XOR U1305 ( .A(a[101]), .B(b[101]), .Z(n2079) );
  NANDN U1306 ( .A(n2078), .B(n2079), .Z(n202) );
  AND U1307 ( .A(n203), .B(n202), .Z(n2098) );
  XOR U1308 ( .A(a[102]), .B(b[102]), .Z(n2099) );
  NANDN U1309 ( .A(n2098), .B(n2099), .Z(n204) );
  AND U1310 ( .A(n205), .B(n204), .Z(n2100) );
  XOR U1311 ( .A(a[103]), .B(b[103]), .Z(n2101) );
  NANDN U1312 ( .A(n2100), .B(n2101), .Z(n206) );
  AND U1313 ( .A(n207), .B(n206), .Z(n2102) );
  XOR U1314 ( .A(a[104]), .B(b[104]), .Z(n2103) );
  NANDN U1315 ( .A(n2102), .B(n2103), .Z(n208) );
  AND U1316 ( .A(n209), .B(n208), .Z(n2104) );
  XOR U1317 ( .A(a[105]), .B(b[105]), .Z(n2105) );
  NANDN U1318 ( .A(n2104), .B(n2105), .Z(n210) );
  AND U1319 ( .A(n211), .B(n210), .Z(n2106) );
  XOR U1320 ( .A(a[106]), .B(b[106]), .Z(n2107) );
  NANDN U1321 ( .A(n2106), .B(n2107), .Z(n212) );
  AND U1322 ( .A(n213), .B(n212), .Z(n2108) );
  XOR U1323 ( .A(a[107]), .B(b[107]), .Z(n2109) );
  NANDN U1324 ( .A(n2108), .B(n2109), .Z(n214) );
  AND U1325 ( .A(n215), .B(n214), .Z(n2110) );
  XOR U1326 ( .A(a[108]), .B(b[108]), .Z(n2111) );
  NANDN U1327 ( .A(n2110), .B(n2111), .Z(n216) );
  AND U1328 ( .A(n217), .B(n216), .Z(n2112) );
  XOR U1329 ( .A(a[109]), .B(b[109]), .Z(n2113) );
  NANDN U1330 ( .A(n2112), .B(n2113), .Z(n218) );
  AND U1331 ( .A(n219), .B(n218), .Z(n2116) );
  XOR U1332 ( .A(a[110]), .B(b[110]), .Z(n2117) );
  NANDN U1333 ( .A(n2116), .B(n2117), .Z(n220) );
  AND U1334 ( .A(n221), .B(n220), .Z(n2118) );
  XOR U1335 ( .A(a[111]), .B(b[111]), .Z(n2119) );
  NANDN U1336 ( .A(n2118), .B(n2119), .Z(n222) );
  AND U1337 ( .A(n223), .B(n222), .Z(n2120) );
  XOR U1338 ( .A(a[112]), .B(b[112]), .Z(n2121) );
  NANDN U1339 ( .A(n2120), .B(n2121), .Z(n224) );
  AND U1340 ( .A(n225), .B(n224), .Z(n2122) );
  XOR U1341 ( .A(a[113]), .B(b[113]), .Z(n2123) );
  NANDN U1342 ( .A(n2122), .B(n2123), .Z(n226) );
  AND U1343 ( .A(n227), .B(n226), .Z(n2124) );
  XOR U1344 ( .A(a[114]), .B(b[114]), .Z(n2125) );
  NANDN U1345 ( .A(n2124), .B(n2125), .Z(n228) );
  AND U1346 ( .A(n229), .B(n228), .Z(n2126) );
  XOR U1347 ( .A(a[115]), .B(b[115]), .Z(n2127) );
  NANDN U1348 ( .A(n2126), .B(n2127), .Z(n230) );
  AND U1349 ( .A(n231), .B(n230), .Z(n2128) );
  XOR U1350 ( .A(a[116]), .B(b[116]), .Z(n2129) );
  NANDN U1351 ( .A(n2128), .B(n2129), .Z(n232) );
  AND U1352 ( .A(n233), .B(n232), .Z(n2130) );
  XOR U1353 ( .A(a[117]), .B(b[117]), .Z(n2131) );
  NANDN U1354 ( .A(n2130), .B(n2131), .Z(n234) );
  AND U1355 ( .A(n235), .B(n234), .Z(n2132) );
  XOR U1356 ( .A(a[118]), .B(b[118]), .Z(n2133) );
  NANDN U1357 ( .A(n2132), .B(n2133), .Z(n236) );
  AND U1358 ( .A(n237), .B(n236), .Z(n2134) );
  XOR U1359 ( .A(a[119]), .B(b[119]), .Z(n2135) );
  NANDN U1360 ( .A(n2134), .B(n2135), .Z(n238) );
  AND U1361 ( .A(n239), .B(n238), .Z(n2138) );
  XOR U1362 ( .A(a[120]), .B(b[120]), .Z(n2139) );
  NANDN U1363 ( .A(n2138), .B(n2139), .Z(n240) );
  AND U1364 ( .A(n241), .B(n240), .Z(n2140) );
  XOR U1365 ( .A(a[121]), .B(b[121]), .Z(n2141) );
  NANDN U1366 ( .A(n2140), .B(n2141), .Z(n242) );
  AND U1367 ( .A(n243), .B(n242), .Z(n2142) );
  XOR U1368 ( .A(a[122]), .B(b[122]), .Z(n2143) );
  NANDN U1369 ( .A(n2142), .B(n2143), .Z(n244) );
  AND U1370 ( .A(n245), .B(n244), .Z(n2144) );
  XOR U1371 ( .A(a[123]), .B(b[123]), .Z(n2145) );
  NANDN U1372 ( .A(n2144), .B(n2145), .Z(n246) );
  AND U1373 ( .A(n247), .B(n246), .Z(n2146) );
  XOR U1374 ( .A(a[124]), .B(b[124]), .Z(n2147) );
  NANDN U1375 ( .A(n2146), .B(n2147), .Z(n248) );
  AND U1376 ( .A(n249), .B(n248), .Z(n2148) );
  XOR U1377 ( .A(a[125]), .B(b[125]), .Z(n2149) );
  NANDN U1378 ( .A(n2148), .B(n2149), .Z(n250) );
  AND U1379 ( .A(n251), .B(n250), .Z(n2150) );
  XOR U1380 ( .A(a[126]), .B(b[126]), .Z(n2151) );
  NANDN U1381 ( .A(n2150), .B(n2151), .Z(n252) );
  AND U1382 ( .A(n253), .B(n252), .Z(n2152) );
  XOR U1383 ( .A(a[127]), .B(b[127]), .Z(n2153) );
  NANDN U1384 ( .A(n2152), .B(n2153), .Z(n254) );
  AND U1385 ( .A(n255), .B(n254), .Z(n2154) );
  XOR U1386 ( .A(a[128]), .B(b[128]), .Z(n2155) );
  NANDN U1387 ( .A(n2154), .B(n2155), .Z(n256) );
  AND U1388 ( .A(n257), .B(n256), .Z(n2156) );
  XOR U1389 ( .A(a[129]), .B(b[129]), .Z(n2157) );
  NANDN U1390 ( .A(n2156), .B(n2157), .Z(n258) );
  AND U1391 ( .A(n259), .B(n258), .Z(n2160) );
  XOR U1392 ( .A(a[130]), .B(b[130]), .Z(n2161) );
  NANDN U1393 ( .A(n2160), .B(n2161), .Z(n260) );
  AND U1394 ( .A(n261), .B(n260), .Z(n2162) );
  XOR U1395 ( .A(a[131]), .B(b[131]), .Z(n2163) );
  NANDN U1396 ( .A(n2162), .B(n2163), .Z(n262) );
  AND U1397 ( .A(n263), .B(n262), .Z(n2164) );
  XOR U1398 ( .A(a[132]), .B(b[132]), .Z(n2165) );
  NANDN U1399 ( .A(n2164), .B(n2165), .Z(n264) );
  AND U1400 ( .A(n265), .B(n264), .Z(n2166) );
  XOR U1401 ( .A(a[133]), .B(b[133]), .Z(n2167) );
  NANDN U1402 ( .A(n2166), .B(n2167), .Z(n266) );
  AND U1403 ( .A(n267), .B(n266), .Z(n2168) );
  XOR U1404 ( .A(a[134]), .B(b[134]), .Z(n2169) );
  NANDN U1405 ( .A(n2168), .B(n2169), .Z(n268) );
  AND U1406 ( .A(n269), .B(n268), .Z(n2170) );
  XOR U1407 ( .A(a[135]), .B(b[135]), .Z(n2171) );
  NANDN U1408 ( .A(n2170), .B(n2171), .Z(n270) );
  AND U1409 ( .A(n271), .B(n270), .Z(n2172) );
  XOR U1410 ( .A(a[136]), .B(b[136]), .Z(n2173) );
  NANDN U1411 ( .A(n2172), .B(n2173), .Z(n272) );
  AND U1412 ( .A(n273), .B(n272), .Z(n2174) );
  XOR U1413 ( .A(a[137]), .B(b[137]), .Z(n2175) );
  NANDN U1414 ( .A(n2174), .B(n2175), .Z(n274) );
  AND U1415 ( .A(n275), .B(n274), .Z(n2176) );
  XOR U1416 ( .A(a[138]), .B(b[138]), .Z(n2177) );
  NANDN U1417 ( .A(n2176), .B(n2177), .Z(n276) );
  AND U1418 ( .A(n277), .B(n276), .Z(n2178) );
  XOR U1419 ( .A(a[139]), .B(b[139]), .Z(n2179) );
  NANDN U1420 ( .A(n2178), .B(n2179), .Z(n278) );
  AND U1421 ( .A(n279), .B(n278), .Z(n2182) );
  XOR U1422 ( .A(a[140]), .B(b[140]), .Z(n2183) );
  NANDN U1423 ( .A(n2182), .B(n2183), .Z(n280) );
  AND U1424 ( .A(n281), .B(n280), .Z(n2184) );
  XOR U1425 ( .A(a[141]), .B(b[141]), .Z(n2185) );
  NANDN U1426 ( .A(n2184), .B(n2185), .Z(n282) );
  AND U1427 ( .A(n283), .B(n282), .Z(n2186) );
  XOR U1428 ( .A(a[142]), .B(b[142]), .Z(n2187) );
  NANDN U1429 ( .A(n2186), .B(n2187), .Z(n284) );
  AND U1430 ( .A(n285), .B(n284), .Z(n2188) );
  XOR U1431 ( .A(a[143]), .B(b[143]), .Z(n2189) );
  NANDN U1432 ( .A(n2188), .B(n2189), .Z(n286) );
  AND U1433 ( .A(n287), .B(n286), .Z(n2190) );
  XOR U1434 ( .A(a[144]), .B(b[144]), .Z(n2191) );
  NANDN U1435 ( .A(n2190), .B(n2191), .Z(n288) );
  AND U1436 ( .A(n289), .B(n288), .Z(n2192) );
  XOR U1437 ( .A(a[145]), .B(b[145]), .Z(n2193) );
  NANDN U1438 ( .A(n2192), .B(n2193), .Z(n290) );
  AND U1439 ( .A(n291), .B(n290), .Z(n2194) );
  XOR U1440 ( .A(a[146]), .B(b[146]), .Z(n2195) );
  NANDN U1441 ( .A(n2194), .B(n2195), .Z(n292) );
  AND U1442 ( .A(n293), .B(n292), .Z(n2196) );
  XOR U1443 ( .A(a[147]), .B(b[147]), .Z(n2197) );
  NANDN U1444 ( .A(n2196), .B(n2197), .Z(n294) );
  AND U1445 ( .A(n295), .B(n294), .Z(n2198) );
  XOR U1446 ( .A(a[148]), .B(b[148]), .Z(n2199) );
  NANDN U1447 ( .A(n2198), .B(n2199), .Z(n296) );
  AND U1448 ( .A(n297), .B(n296), .Z(n2200) );
  XOR U1449 ( .A(a[149]), .B(b[149]), .Z(n2201) );
  NANDN U1450 ( .A(n2200), .B(n2201), .Z(n298) );
  AND U1451 ( .A(n299), .B(n298), .Z(n2204) );
  XOR U1452 ( .A(a[150]), .B(b[150]), .Z(n2205) );
  NANDN U1453 ( .A(n2204), .B(n2205), .Z(n300) );
  AND U1454 ( .A(n301), .B(n300), .Z(n2206) );
  XOR U1455 ( .A(a[151]), .B(b[151]), .Z(n2207) );
  NANDN U1456 ( .A(n2206), .B(n2207), .Z(n302) );
  AND U1457 ( .A(n303), .B(n302), .Z(n2208) );
  XOR U1458 ( .A(a[152]), .B(b[152]), .Z(n2209) );
  NANDN U1459 ( .A(n2208), .B(n2209), .Z(n304) );
  AND U1460 ( .A(n305), .B(n304), .Z(n2210) );
  XOR U1461 ( .A(a[153]), .B(b[153]), .Z(n2211) );
  NANDN U1462 ( .A(n2210), .B(n2211), .Z(n306) );
  AND U1463 ( .A(n307), .B(n306), .Z(n2212) );
  XOR U1464 ( .A(a[154]), .B(b[154]), .Z(n2213) );
  NANDN U1465 ( .A(n2212), .B(n2213), .Z(n308) );
  AND U1466 ( .A(n309), .B(n308), .Z(n2214) );
  XOR U1467 ( .A(a[155]), .B(b[155]), .Z(n2215) );
  NANDN U1468 ( .A(n2214), .B(n2215), .Z(n310) );
  AND U1469 ( .A(n311), .B(n310), .Z(n2216) );
  XOR U1470 ( .A(a[156]), .B(b[156]), .Z(n2217) );
  NANDN U1471 ( .A(n2216), .B(n2217), .Z(n312) );
  AND U1472 ( .A(n313), .B(n312), .Z(n2218) );
  XOR U1473 ( .A(a[157]), .B(b[157]), .Z(n2219) );
  NANDN U1474 ( .A(n2218), .B(n2219), .Z(n314) );
  AND U1475 ( .A(n315), .B(n314), .Z(n2220) );
  XOR U1476 ( .A(a[158]), .B(b[158]), .Z(n2221) );
  NANDN U1477 ( .A(n2220), .B(n2221), .Z(n316) );
  AND U1478 ( .A(n317), .B(n316), .Z(n2222) );
  XOR U1479 ( .A(a[159]), .B(b[159]), .Z(n2223) );
  NANDN U1480 ( .A(n2222), .B(n2223), .Z(n318) );
  AND U1481 ( .A(n319), .B(n318), .Z(n2226) );
  XOR U1482 ( .A(a[160]), .B(b[160]), .Z(n2227) );
  NANDN U1483 ( .A(n2226), .B(n2227), .Z(n320) );
  AND U1484 ( .A(n321), .B(n320), .Z(n2228) );
  XOR U1485 ( .A(a[161]), .B(b[161]), .Z(n2229) );
  NANDN U1486 ( .A(n2228), .B(n2229), .Z(n322) );
  AND U1487 ( .A(n323), .B(n322), .Z(n2230) );
  XOR U1488 ( .A(a[162]), .B(b[162]), .Z(n2231) );
  NANDN U1489 ( .A(n2230), .B(n2231), .Z(n324) );
  AND U1490 ( .A(n325), .B(n324), .Z(n2232) );
  XOR U1491 ( .A(a[163]), .B(b[163]), .Z(n2233) );
  NANDN U1492 ( .A(n2232), .B(n2233), .Z(n326) );
  AND U1493 ( .A(n327), .B(n326), .Z(n2234) );
  XOR U1494 ( .A(a[164]), .B(b[164]), .Z(n2235) );
  NANDN U1495 ( .A(n2234), .B(n2235), .Z(n328) );
  AND U1496 ( .A(n329), .B(n328), .Z(n2236) );
  XOR U1497 ( .A(a[165]), .B(b[165]), .Z(n2237) );
  NANDN U1498 ( .A(n2236), .B(n2237), .Z(n330) );
  AND U1499 ( .A(n331), .B(n330), .Z(n2238) );
  XOR U1500 ( .A(a[166]), .B(b[166]), .Z(n2239) );
  NANDN U1501 ( .A(n2238), .B(n2239), .Z(n332) );
  AND U1502 ( .A(n333), .B(n332), .Z(n2240) );
  XOR U1503 ( .A(a[167]), .B(b[167]), .Z(n2241) );
  NANDN U1504 ( .A(n2240), .B(n2241), .Z(n334) );
  AND U1505 ( .A(n335), .B(n334), .Z(n2242) );
  XOR U1506 ( .A(a[168]), .B(b[168]), .Z(n2243) );
  NANDN U1507 ( .A(n2242), .B(n2243), .Z(n336) );
  AND U1508 ( .A(n337), .B(n336), .Z(n2244) );
  XOR U1509 ( .A(a[169]), .B(b[169]), .Z(n2245) );
  NANDN U1510 ( .A(n2244), .B(n2245), .Z(n338) );
  AND U1511 ( .A(n339), .B(n338), .Z(n2248) );
  XOR U1512 ( .A(a[170]), .B(b[170]), .Z(n2249) );
  NANDN U1513 ( .A(n2248), .B(n2249), .Z(n340) );
  AND U1514 ( .A(n341), .B(n340), .Z(n2250) );
  XOR U1515 ( .A(a[171]), .B(b[171]), .Z(n2251) );
  NANDN U1516 ( .A(n2250), .B(n2251), .Z(n342) );
  AND U1517 ( .A(n343), .B(n342), .Z(n2252) );
  XOR U1518 ( .A(a[172]), .B(b[172]), .Z(n2253) );
  NANDN U1519 ( .A(n2252), .B(n2253), .Z(n344) );
  AND U1520 ( .A(n345), .B(n344), .Z(n2254) );
  XOR U1521 ( .A(a[173]), .B(b[173]), .Z(n2255) );
  NANDN U1522 ( .A(n2254), .B(n2255), .Z(n346) );
  AND U1523 ( .A(n347), .B(n346), .Z(n2256) );
  XOR U1524 ( .A(a[174]), .B(b[174]), .Z(n2257) );
  NANDN U1525 ( .A(n2256), .B(n2257), .Z(n348) );
  AND U1526 ( .A(n349), .B(n348), .Z(n2258) );
  XOR U1527 ( .A(a[175]), .B(b[175]), .Z(n2259) );
  NANDN U1528 ( .A(n2258), .B(n2259), .Z(n350) );
  AND U1529 ( .A(n351), .B(n350), .Z(n2260) );
  XOR U1530 ( .A(a[176]), .B(b[176]), .Z(n2261) );
  NANDN U1531 ( .A(n2260), .B(n2261), .Z(n352) );
  AND U1532 ( .A(n353), .B(n352), .Z(n2262) );
  XOR U1533 ( .A(a[177]), .B(b[177]), .Z(n2263) );
  NANDN U1534 ( .A(n2262), .B(n2263), .Z(n354) );
  AND U1535 ( .A(n355), .B(n354), .Z(n2264) );
  XOR U1536 ( .A(a[178]), .B(b[178]), .Z(n2265) );
  NANDN U1537 ( .A(n2264), .B(n2265), .Z(n356) );
  AND U1538 ( .A(n357), .B(n356), .Z(n2266) );
  XOR U1539 ( .A(a[179]), .B(b[179]), .Z(n2267) );
  NANDN U1540 ( .A(n2266), .B(n2267), .Z(n358) );
  AND U1541 ( .A(n359), .B(n358), .Z(n2270) );
  XOR U1542 ( .A(a[180]), .B(b[180]), .Z(n2271) );
  NANDN U1543 ( .A(n2270), .B(n2271), .Z(n360) );
  AND U1544 ( .A(n361), .B(n360), .Z(n2272) );
  XOR U1545 ( .A(a[181]), .B(b[181]), .Z(n2273) );
  NANDN U1546 ( .A(n2272), .B(n2273), .Z(n362) );
  AND U1547 ( .A(n363), .B(n362), .Z(n2274) );
  XOR U1548 ( .A(a[182]), .B(b[182]), .Z(n2275) );
  NANDN U1549 ( .A(n2274), .B(n2275), .Z(n364) );
  AND U1550 ( .A(n365), .B(n364), .Z(n2276) );
  XOR U1551 ( .A(a[183]), .B(b[183]), .Z(n2277) );
  NANDN U1552 ( .A(n2276), .B(n2277), .Z(n366) );
  AND U1553 ( .A(n367), .B(n366), .Z(n2278) );
  XOR U1554 ( .A(a[184]), .B(b[184]), .Z(n2279) );
  NANDN U1555 ( .A(n2278), .B(n2279), .Z(n368) );
  AND U1556 ( .A(n369), .B(n368), .Z(n2280) );
  XOR U1557 ( .A(a[185]), .B(b[185]), .Z(n2281) );
  NANDN U1558 ( .A(n2280), .B(n2281), .Z(n370) );
  AND U1559 ( .A(n371), .B(n370), .Z(n2282) );
  XOR U1560 ( .A(a[186]), .B(b[186]), .Z(n2283) );
  NANDN U1561 ( .A(n2282), .B(n2283), .Z(n372) );
  AND U1562 ( .A(n373), .B(n372), .Z(n2284) );
  XOR U1563 ( .A(a[187]), .B(b[187]), .Z(n2285) );
  NANDN U1564 ( .A(n2284), .B(n2285), .Z(n374) );
  AND U1565 ( .A(n375), .B(n374), .Z(n2286) );
  XOR U1566 ( .A(a[188]), .B(b[188]), .Z(n2287) );
  NANDN U1567 ( .A(n2286), .B(n2287), .Z(n376) );
  AND U1568 ( .A(n377), .B(n376), .Z(n2288) );
  XOR U1569 ( .A(a[189]), .B(b[189]), .Z(n2289) );
  NANDN U1570 ( .A(n2288), .B(n2289), .Z(n378) );
  AND U1571 ( .A(n379), .B(n378), .Z(n2292) );
  XOR U1572 ( .A(a[190]), .B(b[190]), .Z(n2293) );
  NANDN U1573 ( .A(n2292), .B(n2293), .Z(n380) );
  AND U1574 ( .A(n381), .B(n380), .Z(n2294) );
  XOR U1575 ( .A(a[191]), .B(b[191]), .Z(n2295) );
  NANDN U1576 ( .A(n2294), .B(n2295), .Z(n382) );
  AND U1577 ( .A(n383), .B(n382), .Z(n2296) );
  XOR U1578 ( .A(a[192]), .B(b[192]), .Z(n2297) );
  NANDN U1579 ( .A(n2296), .B(n2297), .Z(n384) );
  AND U1580 ( .A(n385), .B(n384), .Z(n2298) );
  XOR U1581 ( .A(a[193]), .B(b[193]), .Z(n2299) );
  NANDN U1582 ( .A(n2298), .B(n2299), .Z(n386) );
  AND U1583 ( .A(n387), .B(n386), .Z(n2300) );
  XOR U1584 ( .A(a[194]), .B(b[194]), .Z(n2301) );
  NANDN U1585 ( .A(n2300), .B(n2301), .Z(n388) );
  AND U1586 ( .A(n389), .B(n388), .Z(n2302) );
  XOR U1587 ( .A(a[195]), .B(b[195]), .Z(n2303) );
  NANDN U1588 ( .A(n2302), .B(n2303), .Z(n390) );
  AND U1589 ( .A(n391), .B(n390), .Z(n2304) );
  XOR U1590 ( .A(a[196]), .B(b[196]), .Z(n2305) );
  NANDN U1591 ( .A(n2304), .B(n2305), .Z(n392) );
  AND U1592 ( .A(n393), .B(n392), .Z(n2306) );
  XOR U1593 ( .A(a[197]), .B(b[197]), .Z(n2307) );
  NANDN U1594 ( .A(n2306), .B(n2307), .Z(n394) );
  AND U1595 ( .A(n395), .B(n394), .Z(n2308) );
  XOR U1596 ( .A(a[198]), .B(b[198]), .Z(n2309) );
  NANDN U1597 ( .A(n2308), .B(n2309), .Z(n396) );
  AND U1598 ( .A(n397), .B(n396), .Z(n2310) );
  XOR U1599 ( .A(a[199]), .B(b[199]), .Z(n2311) );
  NANDN U1600 ( .A(n2310), .B(n2311), .Z(n398) );
  AND U1601 ( .A(n399), .B(n398), .Z(n2316) );
  XOR U1602 ( .A(a[200]), .B(b[200]), .Z(n2317) );
  NANDN U1603 ( .A(n2316), .B(n2317), .Z(n400) );
  AND U1604 ( .A(n401), .B(n400), .Z(n2318) );
  XOR U1605 ( .A(a[201]), .B(b[201]), .Z(n2319) );
  NANDN U1606 ( .A(n2318), .B(n2319), .Z(n402) );
  AND U1607 ( .A(n403), .B(n402), .Z(n2320) );
  XOR U1608 ( .A(a[202]), .B(b[202]), .Z(n2321) );
  NANDN U1609 ( .A(n2320), .B(n2321), .Z(n404) );
  AND U1610 ( .A(n405), .B(n404), .Z(n2322) );
  XOR U1611 ( .A(a[203]), .B(b[203]), .Z(n2323) );
  NANDN U1612 ( .A(n2322), .B(n2323), .Z(n406) );
  AND U1613 ( .A(n407), .B(n406), .Z(n2324) );
  XOR U1614 ( .A(a[204]), .B(b[204]), .Z(n2325) );
  NANDN U1615 ( .A(n2324), .B(n2325), .Z(n408) );
  AND U1616 ( .A(n409), .B(n408), .Z(n2326) );
  XOR U1617 ( .A(a[205]), .B(b[205]), .Z(n2327) );
  NANDN U1618 ( .A(n2326), .B(n2327), .Z(n410) );
  AND U1619 ( .A(n411), .B(n410), .Z(n2328) );
  XOR U1620 ( .A(a[206]), .B(b[206]), .Z(n2329) );
  NANDN U1621 ( .A(n2328), .B(n2329), .Z(n412) );
  AND U1622 ( .A(n413), .B(n412), .Z(n2330) );
  XOR U1623 ( .A(a[207]), .B(b[207]), .Z(n2331) );
  NANDN U1624 ( .A(n2330), .B(n2331), .Z(n414) );
  AND U1625 ( .A(n415), .B(n414), .Z(n2332) );
  XOR U1626 ( .A(a[208]), .B(b[208]), .Z(n2333) );
  NANDN U1627 ( .A(n2332), .B(n2333), .Z(n416) );
  AND U1628 ( .A(n417), .B(n416), .Z(n2334) );
  XOR U1629 ( .A(a[209]), .B(b[209]), .Z(n2335) );
  NANDN U1630 ( .A(n2334), .B(n2335), .Z(n418) );
  AND U1631 ( .A(n419), .B(n418), .Z(n2338) );
  XOR U1632 ( .A(a[210]), .B(b[210]), .Z(n2339) );
  NANDN U1633 ( .A(n2338), .B(n2339), .Z(n420) );
  AND U1634 ( .A(n421), .B(n420), .Z(n2340) );
  XOR U1635 ( .A(a[211]), .B(b[211]), .Z(n2341) );
  NANDN U1636 ( .A(n2340), .B(n2341), .Z(n422) );
  AND U1637 ( .A(n423), .B(n422), .Z(n2342) );
  XOR U1638 ( .A(a[212]), .B(b[212]), .Z(n2343) );
  NANDN U1639 ( .A(n2342), .B(n2343), .Z(n424) );
  AND U1640 ( .A(n425), .B(n424), .Z(n2344) );
  XOR U1641 ( .A(a[213]), .B(b[213]), .Z(n2345) );
  NANDN U1642 ( .A(n2344), .B(n2345), .Z(n426) );
  AND U1643 ( .A(n427), .B(n426), .Z(n2346) );
  XOR U1644 ( .A(a[214]), .B(b[214]), .Z(n2347) );
  NANDN U1645 ( .A(n2346), .B(n2347), .Z(n428) );
  AND U1646 ( .A(n429), .B(n428), .Z(n2348) );
  XOR U1647 ( .A(a[215]), .B(b[215]), .Z(n2349) );
  NANDN U1648 ( .A(n2348), .B(n2349), .Z(n430) );
  AND U1649 ( .A(n431), .B(n430), .Z(n2350) );
  XOR U1650 ( .A(a[216]), .B(b[216]), .Z(n2351) );
  NANDN U1651 ( .A(n2350), .B(n2351), .Z(n432) );
  AND U1652 ( .A(n433), .B(n432), .Z(n2352) );
  XOR U1653 ( .A(a[217]), .B(b[217]), .Z(n2353) );
  NANDN U1654 ( .A(n2352), .B(n2353), .Z(n434) );
  AND U1655 ( .A(n435), .B(n434), .Z(n2354) );
  XOR U1656 ( .A(a[218]), .B(b[218]), .Z(n2355) );
  NANDN U1657 ( .A(n2354), .B(n2355), .Z(n436) );
  AND U1658 ( .A(n437), .B(n436), .Z(n2356) );
  XOR U1659 ( .A(a[219]), .B(b[219]), .Z(n2357) );
  NANDN U1660 ( .A(n2356), .B(n2357), .Z(n438) );
  AND U1661 ( .A(n439), .B(n438), .Z(n2360) );
  XOR U1662 ( .A(a[220]), .B(b[220]), .Z(n2361) );
  NANDN U1663 ( .A(n2360), .B(n2361), .Z(n440) );
  AND U1664 ( .A(n441), .B(n440), .Z(n2362) );
  XOR U1665 ( .A(a[221]), .B(b[221]), .Z(n2363) );
  NANDN U1666 ( .A(n2362), .B(n2363), .Z(n442) );
  AND U1667 ( .A(n443), .B(n442), .Z(n2364) );
  XOR U1668 ( .A(a[222]), .B(b[222]), .Z(n2365) );
  NANDN U1669 ( .A(n2364), .B(n2365), .Z(n444) );
  AND U1670 ( .A(n445), .B(n444), .Z(n2366) );
  XOR U1671 ( .A(a[223]), .B(b[223]), .Z(n2367) );
  NANDN U1672 ( .A(n2366), .B(n2367), .Z(n446) );
  AND U1673 ( .A(n447), .B(n446), .Z(n2368) );
  XOR U1674 ( .A(a[224]), .B(b[224]), .Z(n2369) );
  NANDN U1675 ( .A(n2368), .B(n2369), .Z(n448) );
  AND U1676 ( .A(n449), .B(n448), .Z(n2370) );
  XOR U1677 ( .A(a[225]), .B(b[225]), .Z(n2371) );
  NANDN U1678 ( .A(n2370), .B(n2371), .Z(n450) );
  AND U1679 ( .A(n451), .B(n450), .Z(n2372) );
  XOR U1680 ( .A(a[226]), .B(b[226]), .Z(n2373) );
  NANDN U1681 ( .A(n2372), .B(n2373), .Z(n452) );
  AND U1682 ( .A(n453), .B(n452), .Z(n2374) );
  XOR U1683 ( .A(a[227]), .B(b[227]), .Z(n2375) );
  NANDN U1684 ( .A(n2374), .B(n2375), .Z(n454) );
  AND U1685 ( .A(n455), .B(n454), .Z(n2376) );
  XOR U1686 ( .A(a[228]), .B(b[228]), .Z(n2377) );
  NANDN U1687 ( .A(n2376), .B(n2377), .Z(n456) );
  AND U1688 ( .A(n457), .B(n456), .Z(n2378) );
  XOR U1689 ( .A(a[229]), .B(b[229]), .Z(n2379) );
  NANDN U1690 ( .A(n2378), .B(n2379), .Z(n458) );
  AND U1691 ( .A(n459), .B(n458), .Z(n2382) );
  XOR U1692 ( .A(a[230]), .B(b[230]), .Z(n2383) );
  NANDN U1693 ( .A(n2382), .B(n2383), .Z(n460) );
  AND U1694 ( .A(n461), .B(n460), .Z(n2384) );
  XOR U1695 ( .A(a[231]), .B(b[231]), .Z(n2385) );
  NANDN U1696 ( .A(n2384), .B(n2385), .Z(n462) );
  AND U1697 ( .A(n463), .B(n462), .Z(n2386) );
  XOR U1698 ( .A(a[232]), .B(b[232]), .Z(n2387) );
  NANDN U1699 ( .A(n2386), .B(n2387), .Z(n464) );
  AND U1700 ( .A(n465), .B(n464), .Z(n2388) );
  XOR U1701 ( .A(a[233]), .B(b[233]), .Z(n2389) );
  NANDN U1702 ( .A(n2388), .B(n2389), .Z(n466) );
  AND U1703 ( .A(n467), .B(n466), .Z(n2390) );
  XOR U1704 ( .A(a[234]), .B(b[234]), .Z(n2391) );
  NANDN U1705 ( .A(n2390), .B(n2391), .Z(n468) );
  AND U1706 ( .A(n469), .B(n468), .Z(n2392) );
  XOR U1707 ( .A(a[235]), .B(b[235]), .Z(n2393) );
  NANDN U1708 ( .A(n2392), .B(n2393), .Z(n470) );
  AND U1709 ( .A(n471), .B(n470), .Z(n2394) );
  XOR U1710 ( .A(a[236]), .B(b[236]), .Z(n2395) );
  NANDN U1711 ( .A(n2394), .B(n2395), .Z(n472) );
  AND U1712 ( .A(n473), .B(n472), .Z(n2396) );
  XOR U1713 ( .A(a[237]), .B(b[237]), .Z(n2397) );
  NANDN U1714 ( .A(n2396), .B(n2397), .Z(n474) );
  AND U1715 ( .A(n475), .B(n474), .Z(n2398) );
  XOR U1716 ( .A(a[238]), .B(b[238]), .Z(n2399) );
  NANDN U1717 ( .A(n2398), .B(n2399), .Z(n476) );
  AND U1718 ( .A(n477), .B(n476), .Z(n2400) );
  XOR U1719 ( .A(a[239]), .B(b[239]), .Z(n2401) );
  NANDN U1720 ( .A(n2400), .B(n2401), .Z(n478) );
  AND U1721 ( .A(n479), .B(n478), .Z(n2404) );
  XOR U1722 ( .A(a[240]), .B(b[240]), .Z(n2405) );
  NANDN U1723 ( .A(n2404), .B(n2405), .Z(n480) );
  AND U1724 ( .A(n481), .B(n480), .Z(n2406) );
  XOR U1725 ( .A(a[241]), .B(b[241]), .Z(n2407) );
  NANDN U1726 ( .A(n2406), .B(n2407), .Z(n482) );
  AND U1727 ( .A(n483), .B(n482), .Z(n2408) );
  XOR U1728 ( .A(a[242]), .B(b[242]), .Z(n2409) );
  NANDN U1729 ( .A(n2408), .B(n2409), .Z(n484) );
  AND U1730 ( .A(n485), .B(n484), .Z(n2410) );
  XOR U1731 ( .A(a[243]), .B(b[243]), .Z(n2411) );
  NANDN U1732 ( .A(n2410), .B(n2411), .Z(n486) );
  AND U1733 ( .A(n487), .B(n486), .Z(n2412) );
  XOR U1734 ( .A(a[244]), .B(b[244]), .Z(n2413) );
  NANDN U1735 ( .A(n2412), .B(n2413), .Z(n488) );
  AND U1736 ( .A(n489), .B(n488), .Z(n2414) );
  XOR U1737 ( .A(a[245]), .B(b[245]), .Z(n2415) );
  NANDN U1738 ( .A(n2414), .B(n2415), .Z(n490) );
  AND U1739 ( .A(n491), .B(n490), .Z(n2416) );
  XOR U1740 ( .A(a[246]), .B(b[246]), .Z(n2417) );
  NANDN U1741 ( .A(n2416), .B(n2417), .Z(n492) );
  AND U1742 ( .A(n493), .B(n492), .Z(n2418) );
  XOR U1743 ( .A(a[247]), .B(b[247]), .Z(n2419) );
  NANDN U1744 ( .A(n2418), .B(n2419), .Z(n494) );
  AND U1745 ( .A(n495), .B(n494), .Z(n2420) );
  XOR U1746 ( .A(a[248]), .B(b[248]), .Z(n2421) );
  NANDN U1747 ( .A(n2420), .B(n2421), .Z(n496) );
  AND U1748 ( .A(n497), .B(n496), .Z(n2422) );
  XOR U1749 ( .A(a[249]), .B(b[249]), .Z(n2423) );
  NANDN U1750 ( .A(n2422), .B(n2423), .Z(n498) );
  AND U1751 ( .A(n499), .B(n498), .Z(n2426) );
  XOR U1752 ( .A(a[250]), .B(b[250]), .Z(n2427) );
  NANDN U1753 ( .A(n2426), .B(n2427), .Z(n500) );
  AND U1754 ( .A(n501), .B(n500), .Z(n2428) );
  XOR U1755 ( .A(a[251]), .B(b[251]), .Z(n2429) );
  NANDN U1756 ( .A(n2428), .B(n2429), .Z(n502) );
  AND U1757 ( .A(n503), .B(n502), .Z(n2430) );
  XOR U1758 ( .A(a[252]), .B(b[252]), .Z(n2431) );
  NANDN U1759 ( .A(n2430), .B(n2431), .Z(n504) );
  AND U1760 ( .A(n505), .B(n504), .Z(n2432) );
  XOR U1761 ( .A(a[253]), .B(b[253]), .Z(n2433) );
  NANDN U1762 ( .A(n2432), .B(n2433), .Z(n506) );
  AND U1763 ( .A(n507), .B(n506), .Z(n2434) );
  XOR U1764 ( .A(a[254]), .B(b[254]), .Z(n2435) );
  NANDN U1765 ( .A(n2434), .B(n2435), .Z(n508) );
  AND U1766 ( .A(n509), .B(n508), .Z(n2436) );
  XOR U1767 ( .A(a[255]), .B(b[255]), .Z(n2437) );
  NANDN U1768 ( .A(n2436), .B(n2437), .Z(n510) );
  AND U1769 ( .A(n511), .B(n510), .Z(n2438) );
  XOR U1770 ( .A(a[256]), .B(b[256]), .Z(n2439) );
  NANDN U1771 ( .A(n2438), .B(n2439), .Z(n512) );
  AND U1772 ( .A(n513), .B(n512), .Z(n2440) );
  XOR U1773 ( .A(a[257]), .B(b[257]), .Z(n2441) );
  NANDN U1774 ( .A(n2440), .B(n2441), .Z(n514) );
  AND U1775 ( .A(n515), .B(n514), .Z(n2442) );
  XOR U1776 ( .A(a[258]), .B(b[258]), .Z(n2443) );
  NANDN U1777 ( .A(n2442), .B(n2443), .Z(n516) );
  AND U1778 ( .A(n517), .B(n516), .Z(n2444) );
  XOR U1779 ( .A(a[259]), .B(b[259]), .Z(n2445) );
  NANDN U1780 ( .A(n2444), .B(n2445), .Z(n518) );
  AND U1781 ( .A(n519), .B(n518), .Z(n2448) );
  XOR U1782 ( .A(a[260]), .B(b[260]), .Z(n2449) );
  NANDN U1783 ( .A(n2448), .B(n2449), .Z(n520) );
  AND U1784 ( .A(n521), .B(n520), .Z(n2450) );
  XOR U1785 ( .A(a[261]), .B(b[261]), .Z(n2451) );
  NANDN U1786 ( .A(n2450), .B(n2451), .Z(n522) );
  AND U1787 ( .A(n523), .B(n522), .Z(n2452) );
  XOR U1788 ( .A(a[262]), .B(b[262]), .Z(n2453) );
  NANDN U1789 ( .A(n2452), .B(n2453), .Z(n524) );
  AND U1790 ( .A(n525), .B(n524), .Z(n2454) );
  XOR U1791 ( .A(a[263]), .B(b[263]), .Z(n2455) );
  NANDN U1792 ( .A(n2454), .B(n2455), .Z(n526) );
  AND U1793 ( .A(n527), .B(n526), .Z(n2456) );
  XOR U1794 ( .A(a[264]), .B(b[264]), .Z(n2457) );
  NANDN U1795 ( .A(n2456), .B(n2457), .Z(n528) );
  AND U1796 ( .A(n529), .B(n528), .Z(n2458) );
  XOR U1797 ( .A(a[265]), .B(b[265]), .Z(n2459) );
  NANDN U1798 ( .A(n2458), .B(n2459), .Z(n530) );
  AND U1799 ( .A(n531), .B(n530), .Z(n2460) );
  XOR U1800 ( .A(a[266]), .B(b[266]), .Z(n2461) );
  NANDN U1801 ( .A(n2460), .B(n2461), .Z(n532) );
  AND U1802 ( .A(n533), .B(n532), .Z(n2462) );
  XOR U1803 ( .A(a[267]), .B(b[267]), .Z(n2463) );
  NANDN U1804 ( .A(n2462), .B(n2463), .Z(n534) );
  AND U1805 ( .A(n535), .B(n534), .Z(n2464) );
  XOR U1806 ( .A(a[268]), .B(b[268]), .Z(n2465) );
  NANDN U1807 ( .A(n2464), .B(n2465), .Z(n536) );
  AND U1808 ( .A(n537), .B(n536), .Z(n2466) );
  XOR U1809 ( .A(a[269]), .B(b[269]), .Z(n2467) );
  NANDN U1810 ( .A(n2466), .B(n2467), .Z(n538) );
  AND U1811 ( .A(n539), .B(n538), .Z(n2470) );
  XOR U1812 ( .A(a[270]), .B(b[270]), .Z(n2471) );
  NANDN U1813 ( .A(n2470), .B(n2471), .Z(n540) );
  AND U1814 ( .A(n541), .B(n540), .Z(n2472) );
  XOR U1815 ( .A(a[271]), .B(b[271]), .Z(n2473) );
  NANDN U1816 ( .A(n2472), .B(n2473), .Z(n542) );
  AND U1817 ( .A(n543), .B(n542), .Z(n2474) );
  XOR U1818 ( .A(a[272]), .B(b[272]), .Z(n2475) );
  NANDN U1819 ( .A(n2474), .B(n2475), .Z(n544) );
  AND U1820 ( .A(n545), .B(n544), .Z(n2476) );
  XOR U1821 ( .A(a[273]), .B(b[273]), .Z(n2477) );
  NANDN U1822 ( .A(n2476), .B(n2477), .Z(n546) );
  AND U1823 ( .A(n547), .B(n546), .Z(n2478) );
  XOR U1824 ( .A(a[274]), .B(b[274]), .Z(n2479) );
  NANDN U1825 ( .A(n2478), .B(n2479), .Z(n548) );
  AND U1826 ( .A(n549), .B(n548), .Z(n2480) );
  XOR U1827 ( .A(a[275]), .B(b[275]), .Z(n2481) );
  NANDN U1828 ( .A(n2480), .B(n2481), .Z(n550) );
  AND U1829 ( .A(n551), .B(n550), .Z(n2482) );
  XOR U1830 ( .A(a[276]), .B(b[276]), .Z(n2483) );
  NANDN U1831 ( .A(n2482), .B(n2483), .Z(n552) );
  AND U1832 ( .A(n553), .B(n552), .Z(n2484) );
  XOR U1833 ( .A(a[277]), .B(b[277]), .Z(n2485) );
  NANDN U1834 ( .A(n2484), .B(n2485), .Z(n554) );
  AND U1835 ( .A(n555), .B(n554), .Z(n2486) );
  XOR U1836 ( .A(a[278]), .B(b[278]), .Z(n2487) );
  NANDN U1837 ( .A(n2486), .B(n2487), .Z(n556) );
  AND U1838 ( .A(n557), .B(n556), .Z(n2488) );
  XOR U1839 ( .A(a[279]), .B(b[279]), .Z(n2489) );
  NANDN U1840 ( .A(n2488), .B(n2489), .Z(n558) );
  AND U1841 ( .A(n559), .B(n558), .Z(n2492) );
  XOR U1842 ( .A(a[280]), .B(b[280]), .Z(n2493) );
  NANDN U1843 ( .A(n2492), .B(n2493), .Z(n560) );
  AND U1844 ( .A(n561), .B(n560), .Z(n2494) );
  XOR U1845 ( .A(a[281]), .B(b[281]), .Z(n2495) );
  NANDN U1846 ( .A(n2494), .B(n2495), .Z(n562) );
  AND U1847 ( .A(n563), .B(n562), .Z(n2496) );
  XOR U1848 ( .A(a[282]), .B(b[282]), .Z(n2497) );
  NANDN U1849 ( .A(n2496), .B(n2497), .Z(n564) );
  AND U1850 ( .A(n565), .B(n564), .Z(n2498) );
  XOR U1851 ( .A(a[283]), .B(b[283]), .Z(n2499) );
  NANDN U1852 ( .A(n2498), .B(n2499), .Z(n566) );
  AND U1853 ( .A(n567), .B(n566), .Z(n2500) );
  XOR U1854 ( .A(a[284]), .B(b[284]), .Z(n2501) );
  NANDN U1855 ( .A(n2500), .B(n2501), .Z(n568) );
  AND U1856 ( .A(n569), .B(n568), .Z(n2502) );
  XOR U1857 ( .A(a[285]), .B(b[285]), .Z(n2503) );
  NANDN U1858 ( .A(n2502), .B(n2503), .Z(n570) );
  AND U1859 ( .A(n571), .B(n570), .Z(n2504) );
  XOR U1860 ( .A(a[286]), .B(b[286]), .Z(n2505) );
  NANDN U1861 ( .A(n2504), .B(n2505), .Z(n572) );
  AND U1862 ( .A(n573), .B(n572), .Z(n2506) );
  XOR U1863 ( .A(a[287]), .B(b[287]), .Z(n2507) );
  NANDN U1864 ( .A(n2506), .B(n2507), .Z(n574) );
  AND U1865 ( .A(n575), .B(n574), .Z(n2508) );
  XOR U1866 ( .A(a[288]), .B(b[288]), .Z(n2509) );
  NANDN U1867 ( .A(n2508), .B(n2509), .Z(n576) );
  AND U1868 ( .A(n577), .B(n576), .Z(n2510) );
  XOR U1869 ( .A(a[289]), .B(b[289]), .Z(n2511) );
  NANDN U1870 ( .A(n2510), .B(n2511), .Z(n578) );
  AND U1871 ( .A(n579), .B(n578), .Z(n2514) );
  XOR U1872 ( .A(a[290]), .B(b[290]), .Z(n2515) );
  NANDN U1873 ( .A(n2514), .B(n2515), .Z(n580) );
  AND U1874 ( .A(n581), .B(n580), .Z(n2516) );
  XOR U1875 ( .A(a[291]), .B(b[291]), .Z(n2517) );
  NANDN U1876 ( .A(n2516), .B(n2517), .Z(n582) );
  AND U1877 ( .A(n583), .B(n582), .Z(n2518) );
  XOR U1878 ( .A(a[292]), .B(b[292]), .Z(n2519) );
  NANDN U1879 ( .A(n2518), .B(n2519), .Z(n584) );
  AND U1880 ( .A(n585), .B(n584), .Z(n2520) );
  XOR U1881 ( .A(a[293]), .B(b[293]), .Z(n2521) );
  NANDN U1882 ( .A(n2520), .B(n2521), .Z(n586) );
  AND U1883 ( .A(n587), .B(n586), .Z(n2522) );
  XOR U1884 ( .A(a[294]), .B(b[294]), .Z(n2523) );
  NANDN U1885 ( .A(n2522), .B(n2523), .Z(n588) );
  AND U1886 ( .A(n589), .B(n588), .Z(n2524) );
  XOR U1887 ( .A(a[295]), .B(b[295]), .Z(n2525) );
  NANDN U1888 ( .A(n2524), .B(n2525), .Z(n590) );
  AND U1889 ( .A(n591), .B(n590), .Z(n2526) );
  XOR U1890 ( .A(a[296]), .B(b[296]), .Z(n2527) );
  NANDN U1891 ( .A(n2526), .B(n2527), .Z(n592) );
  AND U1892 ( .A(n593), .B(n592), .Z(n2528) );
  XOR U1893 ( .A(a[297]), .B(b[297]), .Z(n2529) );
  NANDN U1894 ( .A(n2528), .B(n2529), .Z(n594) );
  AND U1895 ( .A(n595), .B(n594), .Z(n2530) );
  XOR U1896 ( .A(a[298]), .B(b[298]), .Z(n2531) );
  NANDN U1897 ( .A(n2530), .B(n2531), .Z(n596) );
  AND U1898 ( .A(n597), .B(n596), .Z(n2532) );
  XOR U1899 ( .A(a[299]), .B(b[299]), .Z(n2533) );
  NANDN U1900 ( .A(n2532), .B(n2533), .Z(n598) );
  AND U1901 ( .A(n599), .B(n598), .Z(n2538) );
  XOR U1902 ( .A(a[300]), .B(b[300]), .Z(n2539) );
  NANDN U1903 ( .A(n2538), .B(n2539), .Z(n600) );
  AND U1904 ( .A(n601), .B(n600), .Z(n2540) );
  XOR U1905 ( .A(a[301]), .B(b[301]), .Z(n2541) );
  NANDN U1906 ( .A(n2540), .B(n2541), .Z(n602) );
  AND U1907 ( .A(n603), .B(n602), .Z(n2542) );
  XOR U1908 ( .A(a[302]), .B(b[302]), .Z(n2543) );
  NANDN U1909 ( .A(n2542), .B(n2543), .Z(n604) );
  AND U1910 ( .A(n605), .B(n604), .Z(n2544) );
  XOR U1911 ( .A(a[303]), .B(b[303]), .Z(n2545) );
  NANDN U1912 ( .A(n2544), .B(n2545), .Z(n606) );
  AND U1913 ( .A(n607), .B(n606), .Z(n2546) );
  XOR U1914 ( .A(a[304]), .B(b[304]), .Z(n2547) );
  NANDN U1915 ( .A(n2546), .B(n2547), .Z(n608) );
  AND U1916 ( .A(n609), .B(n608), .Z(n2548) );
  XOR U1917 ( .A(a[305]), .B(b[305]), .Z(n2549) );
  NANDN U1918 ( .A(n2548), .B(n2549), .Z(n610) );
  AND U1919 ( .A(n611), .B(n610), .Z(n2550) );
  XOR U1920 ( .A(a[306]), .B(b[306]), .Z(n2551) );
  NANDN U1921 ( .A(n2550), .B(n2551), .Z(n612) );
  AND U1922 ( .A(n613), .B(n612), .Z(n2552) );
  XOR U1923 ( .A(a[307]), .B(b[307]), .Z(n2553) );
  NANDN U1924 ( .A(n2552), .B(n2553), .Z(n614) );
  AND U1925 ( .A(n615), .B(n614), .Z(n2554) );
  XOR U1926 ( .A(a[308]), .B(b[308]), .Z(n2555) );
  NANDN U1927 ( .A(n2554), .B(n2555), .Z(n616) );
  AND U1928 ( .A(n617), .B(n616), .Z(n2556) );
  XOR U1929 ( .A(a[309]), .B(b[309]), .Z(n2557) );
  NANDN U1930 ( .A(n2556), .B(n2557), .Z(n618) );
  AND U1931 ( .A(n619), .B(n618), .Z(n2560) );
  XOR U1932 ( .A(a[310]), .B(b[310]), .Z(n2561) );
  NANDN U1933 ( .A(n2560), .B(n2561), .Z(n620) );
  AND U1934 ( .A(n621), .B(n620), .Z(n2562) );
  XOR U1935 ( .A(a[311]), .B(b[311]), .Z(n2563) );
  NANDN U1936 ( .A(n2562), .B(n2563), .Z(n622) );
  AND U1937 ( .A(n623), .B(n622), .Z(n2564) );
  XOR U1938 ( .A(a[312]), .B(b[312]), .Z(n2565) );
  NANDN U1939 ( .A(n2564), .B(n2565), .Z(n624) );
  AND U1940 ( .A(n625), .B(n624), .Z(n2566) );
  XOR U1941 ( .A(a[313]), .B(b[313]), .Z(n2567) );
  NANDN U1942 ( .A(n2566), .B(n2567), .Z(n626) );
  AND U1943 ( .A(n627), .B(n626), .Z(n2568) );
  XOR U1944 ( .A(a[314]), .B(b[314]), .Z(n2569) );
  NANDN U1945 ( .A(n2568), .B(n2569), .Z(n628) );
  AND U1946 ( .A(n629), .B(n628), .Z(n2570) );
  XOR U1947 ( .A(a[315]), .B(b[315]), .Z(n2571) );
  NANDN U1948 ( .A(n2570), .B(n2571), .Z(n630) );
  AND U1949 ( .A(n631), .B(n630), .Z(n2572) );
  XOR U1950 ( .A(a[316]), .B(b[316]), .Z(n2573) );
  NANDN U1951 ( .A(n2572), .B(n2573), .Z(n632) );
  AND U1952 ( .A(n633), .B(n632), .Z(n2574) );
  XOR U1953 ( .A(a[317]), .B(b[317]), .Z(n2575) );
  NANDN U1954 ( .A(n2574), .B(n2575), .Z(n634) );
  AND U1955 ( .A(n635), .B(n634), .Z(n2576) );
  XOR U1956 ( .A(a[318]), .B(b[318]), .Z(n2577) );
  NANDN U1957 ( .A(n2576), .B(n2577), .Z(n636) );
  AND U1958 ( .A(n637), .B(n636), .Z(n2578) );
  XOR U1959 ( .A(a[319]), .B(b[319]), .Z(n2579) );
  NANDN U1960 ( .A(n2578), .B(n2579), .Z(n638) );
  AND U1961 ( .A(n639), .B(n638), .Z(n2582) );
  XOR U1962 ( .A(a[320]), .B(b[320]), .Z(n2583) );
  NANDN U1963 ( .A(n2582), .B(n2583), .Z(n640) );
  AND U1964 ( .A(n641), .B(n640), .Z(n2584) );
  XOR U1965 ( .A(a[321]), .B(b[321]), .Z(n2585) );
  NANDN U1966 ( .A(n2584), .B(n2585), .Z(n642) );
  AND U1967 ( .A(n643), .B(n642), .Z(n2586) );
  XOR U1968 ( .A(a[322]), .B(b[322]), .Z(n2587) );
  NANDN U1969 ( .A(n2586), .B(n2587), .Z(n644) );
  AND U1970 ( .A(n645), .B(n644), .Z(n2588) );
  XOR U1971 ( .A(a[323]), .B(b[323]), .Z(n2589) );
  NANDN U1972 ( .A(n2588), .B(n2589), .Z(n646) );
  AND U1973 ( .A(n647), .B(n646), .Z(n2590) );
  XOR U1974 ( .A(a[324]), .B(b[324]), .Z(n2591) );
  NANDN U1975 ( .A(n2590), .B(n2591), .Z(n648) );
  AND U1976 ( .A(n649), .B(n648), .Z(n2592) );
  XOR U1977 ( .A(a[325]), .B(b[325]), .Z(n2593) );
  NANDN U1978 ( .A(n2592), .B(n2593), .Z(n650) );
  AND U1979 ( .A(n651), .B(n650), .Z(n2594) );
  XOR U1980 ( .A(a[326]), .B(b[326]), .Z(n2595) );
  NANDN U1981 ( .A(n2594), .B(n2595), .Z(n652) );
  AND U1982 ( .A(n653), .B(n652), .Z(n2596) );
  XOR U1983 ( .A(a[327]), .B(b[327]), .Z(n2597) );
  NANDN U1984 ( .A(n2596), .B(n2597), .Z(n654) );
  AND U1985 ( .A(n655), .B(n654), .Z(n2598) );
  XOR U1986 ( .A(a[328]), .B(b[328]), .Z(n2599) );
  NANDN U1987 ( .A(n2598), .B(n2599), .Z(n656) );
  AND U1988 ( .A(n657), .B(n656), .Z(n2600) );
  XOR U1989 ( .A(a[329]), .B(b[329]), .Z(n2601) );
  NANDN U1990 ( .A(n2600), .B(n2601), .Z(n658) );
  AND U1991 ( .A(n659), .B(n658), .Z(n2604) );
  XOR U1992 ( .A(a[330]), .B(b[330]), .Z(n2605) );
  NANDN U1993 ( .A(n2604), .B(n2605), .Z(n660) );
  AND U1994 ( .A(n661), .B(n660), .Z(n2606) );
  XOR U1995 ( .A(a[331]), .B(b[331]), .Z(n2607) );
  NANDN U1996 ( .A(n2606), .B(n2607), .Z(n662) );
  AND U1997 ( .A(n663), .B(n662), .Z(n2608) );
  XOR U1998 ( .A(a[332]), .B(b[332]), .Z(n2609) );
  NANDN U1999 ( .A(n2608), .B(n2609), .Z(n664) );
  AND U2000 ( .A(n665), .B(n664), .Z(n2610) );
  XOR U2001 ( .A(a[333]), .B(b[333]), .Z(n2611) );
  NANDN U2002 ( .A(n2610), .B(n2611), .Z(n666) );
  AND U2003 ( .A(n667), .B(n666), .Z(n2612) );
  XOR U2004 ( .A(a[334]), .B(b[334]), .Z(n2613) );
  NANDN U2005 ( .A(n2612), .B(n2613), .Z(n668) );
  AND U2006 ( .A(n669), .B(n668), .Z(n2614) );
  XOR U2007 ( .A(a[335]), .B(b[335]), .Z(n2615) );
  NANDN U2008 ( .A(n2614), .B(n2615), .Z(n670) );
  AND U2009 ( .A(n671), .B(n670), .Z(n2616) );
  XOR U2010 ( .A(a[336]), .B(b[336]), .Z(n2617) );
  NANDN U2011 ( .A(n2616), .B(n2617), .Z(n672) );
  AND U2012 ( .A(n673), .B(n672), .Z(n2618) );
  XOR U2013 ( .A(a[337]), .B(b[337]), .Z(n2619) );
  NANDN U2014 ( .A(n2618), .B(n2619), .Z(n674) );
  AND U2015 ( .A(n675), .B(n674), .Z(n2620) );
  XOR U2016 ( .A(a[338]), .B(b[338]), .Z(n2621) );
  NANDN U2017 ( .A(n2620), .B(n2621), .Z(n676) );
  AND U2018 ( .A(n677), .B(n676), .Z(n2622) );
  XOR U2019 ( .A(a[339]), .B(b[339]), .Z(n2623) );
  NANDN U2020 ( .A(n2622), .B(n2623), .Z(n678) );
  AND U2021 ( .A(n679), .B(n678), .Z(n2626) );
  XOR U2022 ( .A(a[340]), .B(b[340]), .Z(n2627) );
  NANDN U2023 ( .A(n2626), .B(n2627), .Z(n680) );
  AND U2024 ( .A(n681), .B(n680), .Z(n2628) );
  XOR U2025 ( .A(a[341]), .B(b[341]), .Z(n2629) );
  NANDN U2026 ( .A(n2628), .B(n2629), .Z(n682) );
  AND U2027 ( .A(n683), .B(n682), .Z(n2630) );
  XOR U2028 ( .A(a[342]), .B(b[342]), .Z(n2631) );
  NANDN U2029 ( .A(n2630), .B(n2631), .Z(n684) );
  AND U2030 ( .A(n685), .B(n684), .Z(n2632) );
  XOR U2031 ( .A(a[343]), .B(b[343]), .Z(n2633) );
  NANDN U2032 ( .A(n2632), .B(n2633), .Z(n686) );
  AND U2033 ( .A(n687), .B(n686), .Z(n2634) );
  XOR U2034 ( .A(a[344]), .B(b[344]), .Z(n2635) );
  NANDN U2035 ( .A(n2634), .B(n2635), .Z(n688) );
  AND U2036 ( .A(n689), .B(n688), .Z(n2636) );
  XOR U2037 ( .A(a[345]), .B(b[345]), .Z(n2637) );
  NANDN U2038 ( .A(n2636), .B(n2637), .Z(n690) );
  AND U2039 ( .A(n691), .B(n690), .Z(n2638) );
  XOR U2040 ( .A(a[346]), .B(b[346]), .Z(n2639) );
  NANDN U2041 ( .A(n2638), .B(n2639), .Z(n692) );
  AND U2042 ( .A(n693), .B(n692), .Z(n2640) );
  XOR U2043 ( .A(a[347]), .B(b[347]), .Z(n2641) );
  NANDN U2044 ( .A(n2640), .B(n2641), .Z(n694) );
  AND U2045 ( .A(n695), .B(n694), .Z(n2642) );
  XOR U2046 ( .A(a[348]), .B(b[348]), .Z(n2643) );
  NANDN U2047 ( .A(n2642), .B(n2643), .Z(n696) );
  AND U2048 ( .A(n697), .B(n696), .Z(n2644) );
  XOR U2049 ( .A(a[349]), .B(b[349]), .Z(n2645) );
  NANDN U2050 ( .A(n2644), .B(n2645), .Z(n698) );
  AND U2051 ( .A(n699), .B(n698), .Z(n2648) );
  XOR U2052 ( .A(a[350]), .B(b[350]), .Z(n2649) );
  NANDN U2053 ( .A(n2648), .B(n2649), .Z(n700) );
  AND U2054 ( .A(n701), .B(n700), .Z(n2650) );
  XOR U2055 ( .A(a[351]), .B(b[351]), .Z(n2651) );
  NANDN U2056 ( .A(n2650), .B(n2651), .Z(n702) );
  AND U2057 ( .A(n703), .B(n702), .Z(n2652) );
  XOR U2058 ( .A(a[352]), .B(b[352]), .Z(n2653) );
  NANDN U2059 ( .A(n2652), .B(n2653), .Z(n704) );
  AND U2060 ( .A(n705), .B(n704), .Z(n2654) );
  XOR U2061 ( .A(a[353]), .B(b[353]), .Z(n2655) );
  NANDN U2062 ( .A(n2654), .B(n2655), .Z(n706) );
  AND U2063 ( .A(n707), .B(n706), .Z(n2656) );
  XOR U2064 ( .A(a[354]), .B(b[354]), .Z(n2657) );
  NANDN U2065 ( .A(n2656), .B(n2657), .Z(n708) );
  AND U2066 ( .A(n709), .B(n708), .Z(n2658) );
  XOR U2067 ( .A(a[355]), .B(b[355]), .Z(n2659) );
  NANDN U2068 ( .A(n2658), .B(n2659), .Z(n710) );
  AND U2069 ( .A(n711), .B(n710), .Z(n2660) );
  XOR U2070 ( .A(a[356]), .B(b[356]), .Z(n2661) );
  NANDN U2071 ( .A(n2660), .B(n2661), .Z(n712) );
  AND U2072 ( .A(n713), .B(n712), .Z(n2662) );
  XOR U2073 ( .A(a[357]), .B(b[357]), .Z(n2663) );
  NANDN U2074 ( .A(n2662), .B(n2663), .Z(n714) );
  AND U2075 ( .A(n715), .B(n714), .Z(n2664) );
  XOR U2076 ( .A(a[358]), .B(b[358]), .Z(n2665) );
  NANDN U2077 ( .A(n2664), .B(n2665), .Z(n716) );
  AND U2078 ( .A(n717), .B(n716), .Z(n2666) );
  XOR U2079 ( .A(a[359]), .B(b[359]), .Z(n2667) );
  NANDN U2080 ( .A(n2666), .B(n2667), .Z(n718) );
  AND U2081 ( .A(n719), .B(n718), .Z(n2670) );
  XOR U2082 ( .A(a[360]), .B(b[360]), .Z(n2671) );
  NANDN U2083 ( .A(n2670), .B(n2671), .Z(n720) );
  AND U2084 ( .A(n721), .B(n720), .Z(n2672) );
  XOR U2085 ( .A(a[361]), .B(b[361]), .Z(n2673) );
  NANDN U2086 ( .A(n2672), .B(n2673), .Z(n722) );
  AND U2087 ( .A(n723), .B(n722), .Z(n2674) );
  XOR U2088 ( .A(a[362]), .B(b[362]), .Z(n2675) );
  NANDN U2089 ( .A(n2674), .B(n2675), .Z(n724) );
  AND U2090 ( .A(n725), .B(n724), .Z(n2676) );
  XOR U2091 ( .A(a[363]), .B(b[363]), .Z(n2677) );
  NANDN U2092 ( .A(n2676), .B(n2677), .Z(n726) );
  AND U2093 ( .A(n727), .B(n726), .Z(n2678) );
  XOR U2094 ( .A(a[364]), .B(b[364]), .Z(n2679) );
  NANDN U2095 ( .A(n2678), .B(n2679), .Z(n728) );
  AND U2096 ( .A(n729), .B(n728), .Z(n2680) );
  XOR U2097 ( .A(a[365]), .B(b[365]), .Z(n2681) );
  NANDN U2098 ( .A(n2680), .B(n2681), .Z(n730) );
  AND U2099 ( .A(n731), .B(n730), .Z(n2682) );
  XOR U2100 ( .A(a[366]), .B(b[366]), .Z(n2683) );
  NANDN U2101 ( .A(n2682), .B(n2683), .Z(n732) );
  AND U2102 ( .A(n733), .B(n732), .Z(n2684) );
  XOR U2103 ( .A(a[367]), .B(b[367]), .Z(n2685) );
  NANDN U2104 ( .A(n2684), .B(n2685), .Z(n734) );
  AND U2105 ( .A(n735), .B(n734), .Z(n2686) );
  XOR U2106 ( .A(a[368]), .B(b[368]), .Z(n2687) );
  NANDN U2107 ( .A(n2686), .B(n2687), .Z(n736) );
  AND U2108 ( .A(n737), .B(n736), .Z(n2688) );
  XOR U2109 ( .A(a[369]), .B(b[369]), .Z(n2689) );
  NANDN U2110 ( .A(n2688), .B(n2689), .Z(n738) );
  AND U2111 ( .A(n739), .B(n738), .Z(n2692) );
  XOR U2112 ( .A(a[370]), .B(b[370]), .Z(n2693) );
  NANDN U2113 ( .A(n2692), .B(n2693), .Z(n740) );
  AND U2114 ( .A(n741), .B(n740), .Z(n2694) );
  XOR U2115 ( .A(a[371]), .B(b[371]), .Z(n2695) );
  NANDN U2116 ( .A(n2694), .B(n2695), .Z(n742) );
  AND U2117 ( .A(n743), .B(n742), .Z(n2696) );
  XOR U2118 ( .A(a[372]), .B(b[372]), .Z(n2697) );
  NANDN U2119 ( .A(n2696), .B(n2697), .Z(n744) );
  AND U2120 ( .A(n745), .B(n744), .Z(n2698) );
  XOR U2121 ( .A(a[373]), .B(b[373]), .Z(n2699) );
  NANDN U2122 ( .A(n2698), .B(n2699), .Z(n746) );
  AND U2123 ( .A(n747), .B(n746), .Z(n2700) );
  XOR U2124 ( .A(a[374]), .B(b[374]), .Z(n2701) );
  NANDN U2125 ( .A(n2700), .B(n2701), .Z(n748) );
  AND U2126 ( .A(n749), .B(n748), .Z(n2702) );
  XOR U2127 ( .A(a[375]), .B(b[375]), .Z(n2703) );
  NANDN U2128 ( .A(n2702), .B(n2703), .Z(n750) );
  AND U2129 ( .A(n751), .B(n750), .Z(n2704) );
  XOR U2130 ( .A(a[376]), .B(b[376]), .Z(n2705) );
  NANDN U2131 ( .A(n2704), .B(n2705), .Z(n752) );
  AND U2132 ( .A(n753), .B(n752), .Z(n2706) );
  XOR U2133 ( .A(a[377]), .B(b[377]), .Z(n2707) );
  NANDN U2134 ( .A(n2706), .B(n2707), .Z(n754) );
  AND U2135 ( .A(n755), .B(n754), .Z(n2708) );
  XOR U2136 ( .A(a[378]), .B(b[378]), .Z(n2709) );
  NANDN U2137 ( .A(n2708), .B(n2709), .Z(n756) );
  AND U2138 ( .A(n757), .B(n756), .Z(n2710) );
  XOR U2139 ( .A(a[379]), .B(b[379]), .Z(n2711) );
  NANDN U2140 ( .A(n2710), .B(n2711), .Z(n758) );
  AND U2141 ( .A(n759), .B(n758), .Z(n2714) );
  XOR U2142 ( .A(a[380]), .B(b[380]), .Z(n2715) );
  NANDN U2143 ( .A(n2714), .B(n2715), .Z(n760) );
  AND U2144 ( .A(n761), .B(n760), .Z(n2716) );
  XOR U2145 ( .A(a[381]), .B(b[381]), .Z(n2717) );
  NANDN U2146 ( .A(n2716), .B(n2717), .Z(n762) );
  AND U2147 ( .A(n763), .B(n762), .Z(n2718) );
  XOR U2148 ( .A(a[382]), .B(b[382]), .Z(n2719) );
  NANDN U2149 ( .A(n2718), .B(n2719), .Z(n764) );
  AND U2150 ( .A(n765), .B(n764), .Z(n2720) );
  XOR U2151 ( .A(a[383]), .B(b[383]), .Z(n2721) );
  NANDN U2152 ( .A(n2720), .B(n2721), .Z(n766) );
  AND U2153 ( .A(n767), .B(n766), .Z(n2722) );
  XOR U2154 ( .A(a[384]), .B(b[384]), .Z(n2723) );
  NANDN U2155 ( .A(n2722), .B(n2723), .Z(n768) );
  AND U2156 ( .A(n769), .B(n768), .Z(n2724) );
  XOR U2157 ( .A(a[385]), .B(b[385]), .Z(n2725) );
  NANDN U2158 ( .A(n2724), .B(n2725), .Z(n770) );
  AND U2159 ( .A(n771), .B(n770), .Z(n2726) );
  XOR U2160 ( .A(a[386]), .B(b[386]), .Z(n2727) );
  NANDN U2161 ( .A(n2726), .B(n2727), .Z(n772) );
  AND U2162 ( .A(n773), .B(n772), .Z(n2728) );
  XOR U2163 ( .A(a[387]), .B(b[387]), .Z(n2729) );
  NANDN U2164 ( .A(n2728), .B(n2729), .Z(n774) );
  AND U2165 ( .A(n775), .B(n774), .Z(n2730) );
  XOR U2166 ( .A(a[388]), .B(b[388]), .Z(n2731) );
  NANDN U2167 ( .A(n2730), .B(n2731), .Z(n776) );
  AND U2168 ( .A(n777), .B(n776), .Z(n2732) );
  XOR U2169 ( .A(a[389]), .B(b[389]), .Z(n2733) );
  NANDN U2170 ( .A(n2732), .B(n2733), .Z(n778) );
  AND U2171 ( .A(n779), .B(n778), .Z(n2736) );
  XOR U2172 ( .A(a[390]), .B(b[390]), .Z(n2737) );
  NANDN U2173 ( .A(n2736), .B(n2737), .Z(n780) );
  AND U2174 ( .A(n781), .B(n780), .Z(n2738) );
  XOR U2175 ( .A(a[391]), .B(b[391]), .Z(n2739) );
  NANDN U2176 ( .A(n2738), .B(n2739), .Z(n782) );
  AND U2177 ( .A(n783), .B(n782), .Z(n2740) );
  XOR U2178 ( .A(a[392]), .B(b[392]), .Z(n2741) );
  NANDN U2179 ( .A(n2740), .B(n2741), .Z(n784) );
  AND U2180 ( .A(n785), .B(n784), .Z(n2742) );
  XOR U2181 ( .A(a[393]), .B(b[393]), .Z(n2743) );
  NANDN U2182 ( .A(n2742), .B(n2743), .Z(n786) );
  AND U2183 ( .A(n787), .B(n786), .Z(n2744) );
  XOR U2184 ( .A(a[394]), .B(b[394]), .Z(n2745) );
  NANDN U2185 ( .A(n2744), .B(n2745), .Z(n788) );
  AND U2186 ( .A(n789), .B(n788), .Z(n2746) );
  XOR U2187 ( .A(a[395]), .B(b[395]), .Z(n2747) );
  NANDN U2188 ( .A(n2746), .B(n2747), .Z(n790) );
  AND U2189 ( .A(n791), .B(n790), .Z(n2748) );
  XOR U2190 ( .A(a[396]), .B(b[396]), .Z(n2749) );
  NANDN U2191 ( .A(n2748), .B(n2749), .Z(n792) );
  AND U2192 ( .A(n793), .B(n792), .Z(n2750) );
  XOR U2193 ( .A(a[397]), .B(b[397]), .Z(n2751) );
  NANDN U2194 ( .A(n2750), .B(n2751), .Z(n794) );
  AND U2195 ( .A(n795), .B(n794), .Z(n2752) );
  XOR U2196 ( .A(a[398]), .B(b[398]), .Z(n2753) );
  NANDN U2197 ( .A(n2752), .B(n2753), .Z(n796) );
  AND U2198 ( .A(n797), .B(n796), .Z(n2754) );
  XOR U2199 ( .A(a[399]), .B(b[399]), .Z(n2755) );
  NANDN U2200 ( .A(n2754), .B(n2755), .Z(n798) );
  AND U2201 ( .A(n799), .B(n798), .Z(n2760) );
  XOR U2202 ( .A(a[400]), .B(b[400]), .Z(n2761) );
  NANDN U2203 ( .A(n2760), .B(n2761), .Z(n800) );
  AND U2204 ( .A(n801), .B(n800), .Z(n2762) );
  XOR U2205 ( .A(a[401]), .B(b[401]), .Z(n2763) );
  NANDN U2206 ( .A(n2762), .B(n2763), .Z(n802) );
  AND U2207 ( .A(n803), .B(n802), .Z(n2764) );
  XOR U2208 ( .A(a[402]), .B(b[402]), .Z(n2765) );
  NANDN U2209 ( .A(n2764), .B(n2765), .Z(n804) );
  AND U2210 ( .A(n805), .B(n804), .Z(n2766) );
  XOR U2211 ( .A(a[403]), .B(b[403]), .Z(n2767) );
  NANDN U2212 ( .A(n2766), .B(n2767), .Z(n806) );
  AND U2213 ( .A(n807), .B(n806), .Z(n2768) );
  XOR U2214 ( .A(a[404]), .B(b[404]), .Z(n2769) );
  NANDN U2215 ( .A(n2768), .B(n2769), .Z(n808) );
  AND U2216 ( .A(n809), .B(n808), .Z(n2770) );
  XOR U2217 ( .A(a[405]), .B(b[405]), .Z(n2771) );
  NANDN U2218 ( .A(n2770), .B(n2771), .Z(n810) );
  AND U2219 ( .A(n811), .B(n810), .Z(n2772) );
  XOR U2220 ( .A(a[406]), .B(b[406]), .Z(n2773) );
  NANDN U2221 ( .A(n2772), .B(n2773), .Z(n812) );
  AND U2222 ( .A(n813), .B(n812), .Z(n2774) );
  XOR U2223 ( .A(a[407]), .B(b[407]), .Z(n2775) );
  NANDN U2224 ( .A(n2774), .B(n2775), .Z(n814) );
  AND U2225 ( .A(n815), .B(n814), .Z(n2776) );
  XOR U2226 ( .A(a[408]), .B(b[408]), .Z(n2777) );
  NANDN U2227 ( .A(n2776), .B(n2777), .Z(n816) );
  AND U2228 ( .A(n817), .B(n816), .Z(n2778) );
  XOR U2229 ( .A(a[409]), .B(b[409]), .Z(n2779) );
  NANDN U2230 ( .A(n2778), .B(n2779), .Z(n818) );
  AND U2231 ( .A(n819), .B(n818), .Z(n2782) );
  XOR U2232 ( .A(a[410]), .B(b[410]), .Z(n2783) );
  NANDN U2233 ( .A(n2782), .B(n2783), .Z(n820) );
  AND U2234 ( .A(n821), .B(n820), .Z(n2784) );
  XOR U2235 ( .A(a[411]), .B(b[411]), .Z(n2785) );
  NANDN U2236 ( .A(n2784), .B(n2785), .Z(n822) );
  AND U2237 ( .A(n823), .B(n822), .Z(n2786) );
  XOR U2238 ( .A(a[412]), .B(b[412]), .Z(n2787) );
  NANDN U2239 ( .A(n2786), .B(n2787), .Z(n824) );
  AND U2240 ( .A(n825), .B(n824), .Z(n2788) );
  XOR U2241 ( .A(a[413]), .B(b[413]), .Z(n2789) );
  NANDN U2242 ( .A(n2788), .B(n2789), .Z(n826) );
  AND U2243 ( .A(n827), .B(n826), .Z(n2790) );
  XOR U2244 ( .A(a[414]), .B(b[414]), .Z(n2791) );
  NANDN U2245 ( .A(n2790), .B(n2791), .Z(n828) );
  AND U2246 ( .A(n829), .B(n828), .Z(n2792) );
  XOR U2247 ( .A(a[415]), .B(b[415]), .Z(n2793) );
  NANDN U2248 ( .A(n2792), .B(n2793), .Z(n830) );
  AND U2249 ( .A(n831), .B(n830), .Z(n2794) );
  XOR U2250 ( .A(a[416]), .B(b[416]), .Z(n2795) );
  NANDN U2251 ( .A(n2794), .B(n2795), .Z(n832) );
  AND U2252 ( .A(n833), .B(n832), .Z(n2796) );
  XOR U2253 ( .A(a[417]), .B(b[417]), .Z(n2797) );
  NANDN U2254 ( .A(n2796), .B(n2797), .Z(n834) );
  AND U2255 ( .A(n835), .B(n834), .Z(n2798) );
  XOR U2256 ( .A(a[418]), .B(b[418]), .Z(n2799) );
  NANDN U2257 ( .A(n2798), .B(n2799), .Z(n836) );
  AND U2258 ( .A(n837), .B(n836), .Z(n2800) );
  XOR U2259 ( .A(a[419]), .B(b[419]), .Z(n2801) );
  NANDN U2260 ( .A(n2800), .B(n2801), .Z(n838) );
  AND U2261 ( .A(n839), .B(n838), .Z(n2804) );
  XOR U2262 ( .A(a[420]), .B(b[420]), .Z(n2805) );
  NANDN U2263 ( .A(n2804), .B(n2805), .Z(n840) );
  AND U2264 ( .A(n841), .B(n840), .Z(n2806) );
  XOR U2265 ( .A(a[421]), .B(b[421]), .Z(n2807) );
  NANDN U2266 ( .A(n2806), .B(n2807), .Z(n842) );
  AND U2267 ( .A(n843), .B(n842), .Z(n2808) );
  XOR U2268 ( .A(a[422]), .B(b[422]), .Z(n2809) );
  NANDN U2269 ( .A(n2808), .B(n2809), .Z(n844) );
  AND U2270 ( .A(n845), .B(n844), .Z(n2810) );
  XOR U2271 ( .A(a[423]), .B(b[423]), .Z(n2811) );
  NANDN U2272 ( .A(n2810), .B(n2811), .Z(n846) );
  AND U2273 ( .A(n847), .B(n846), .Z(n2812) );
  XOR U2274 ( .A(a[424]), .B(b[424]), .Z(n2813) );
  NANDN U2275 ( .A(n2812), .B(n2813), .Z(n848) );
  AND U2276 ( .A(n849), .B(n848), .Z(n2814) );
  XOR U2277 ( .A(a[425]), .B(b[425]), .Z(n2815) );
  NANDN U2278 ( .A(n2814), .B(n2815), .Z(n850) );
  AND U2279 ( .A(n851), .B(n850), .Z(n2816) );
  XOR U2280 ( .A(a[426]), .B(b[426]), .Z(n2817) );
  NANDN U2281 ( .A(n2816), .B(n2817), .Z(n852) );
  AND U2282 ( .A(n853), .B(n852), .Z(n2818) );
  XOR U2283 ( .A(a[427]), .B(b[427]), .Z(n2819) );
  NANDN U2284 ( .A(n2818), .B(n2819), .Z(n854) );
  AND U2285 ( .A(n855), .B(n854), .Z(n2820) );
  XOR U2286 ( .A(a[428]), .B(b[428]), .Z(n2821) );
  NANDN U2287 ( .A(n2820), .B(n2821), .Z(n856) );
  AND U2288 ( .A(n857), .B(n856), .Z(n2822) );
  XOR U2289 ( .A(a[429]), .B(b[429]), .Z(n2823) );
  NANDN U2290 ( .A(n2822), .B(n2823), .Z(n858) );
  AND U2291 ( .A(n859), .B(n858), .Z(n2826) );
  XOR U2292 ( .A(a[430]), .B(b[430]), .Z(n2827) );
  NANDN U2293 ( .A(n2826), .B(n2827), .Z(n860) );
  AND U2294 ( .A(n861), .B(n860), .Z(n2828) );
  XOR U2295 ( .A(a[431]), .B(b[431]), .Z(n2829) );
  NANDN U2296 ( .A(n2828), .B(n2829), .Z(n862) );
  AND U2297 ( .A(n863), .B(n862), .Z(n2830) );
  XOR U2298 ( .A(a[432]), .B(b[432]), .Z(n2831) );
  NANDN U2299 ( .A(n2830), .B(n2831), .Z(n864) );
  AND U2300 ( .A(n865), .B(n864), .Z(n2832) );
  XOR U2301 ( .A(a[433]), .B(b[433]), .Z(n2833) );
  NANDN U2302 ( .A(n2832), .B(n2833), .Z(n866) );
  AND U2303 ( .A(n867), .B(n866), .Z(n2834) );
  XOR U2304 ( .A(a[434]), .B(b[434]), .Z(n2835) );
  NANDN U2305 ( .A(n2834), .B(n2835), .Z(n868) );
  AND U2306 ( .A(n869), .B(n868), .Z(n2836) );
  XOR U2307 ( .A(a[435]), .B(b[435]), .Z(n2837) );
  NANDN U2308 ( .A(n2836), .B(n2837), .Z(n870) );
  AND U2309 ( .A(n871), .B(n870), .Z(n2838) );
  XOR U2310 ( .A(a[436]), .B(b[436]), .Z(n2839) );
  NANDN U2311 ( .A(n2838), .B(n2839), .Z(n872) );
  AND U2312 ( .A(n873), .B(n872), .Z(n2840) );
  XOR U2313 ( .A(a[437]), .B(b[437]), .Z(n2841) );
  NANDN U2314 ( .A(n2840), .B(n2841), .Z(n874) );
  AND U2315 ( .A(n875), .B(n874), .Z(n2842) );
  XOR U2316 ( .A(a[438]), .B(b[438]), .Z(n2843) );
  NANDN U2317 ( .A(n2842), .B(n2843), .Z(n876) );
  AND U2318 ( .A(n877), .B(n876), .Z(n2844) );
  XOR U2319 ( .A(a[439]), .B(b[439]), .Z(n2845) );
  NANDN U2320 ( .A(n2844), .B(n2845), .Z(n878) );
  AND U2321 ( .A(n879), .B(n878), .Z(n2848) );
  XOR U2322 ( .A(a[440]), .B(b[440]), .Z(n2849) );
  NANDN U2323 ( .A(n2848), .B(n2849), .Z(n880) );
  AND U2324 ( .A(n881), .B(n880), .Z(n2850) );
  XOR U2325 ( .A(a[441]), .B(b[441]), .Z(n2851) );
  NANDN U2326 ( .A(n2850), .B(n2851), .Z(n882) );
  AND U2327 ( .A(n883), .B(n882), .Z(n2852) );
  XOR U2328 ( .A(a[442]), .B(b[442]), .Z(n2853) );
  NANDN U2329 ( .A(n2852), .B(n2853), .Z(n884) );
  AND U2330 ( .A(n885), .B(n884), .Z(n2854) );
  XOR U2331 ( .A(a[443]), .B(b[443]), .Z(n2855) );
  NANDN U2332 ( .A(n2854), .B(n2855), .Z(n886) );
  AND U2333 ( .A(n887), .B(n886), .Z(n2856) );
  XOR U2334 ( .A(a[444]), .B(b[444]), .Z(n2857) );
  NANDN U2335 ( .A(n2856), .B(n2857), .Z(n888) );
  AND U2336 ( .A(n889), .B(n888), .Z(n2858) );
  XOR U2337 ( .A(a[445]), .B(b[445]), .Z(n2859) );
  NANDN U2338 ( .A(n2858), .B(n2859), .Z(n890) );
  AND U2339 ( .A(n891), .B(n890), .Z(n2860) );
  XOR U2340 ( .A(a[446]), .B(b[446]), .Z(n2861) );
  NANDN U2341 ( .A(n2860), .B(n2861), .Z(n892) );
  AND U2342 ( .A(n893), .B(n892), .Z(n2862) );
  XOR U2343 ( .A(a[447]), .B(b[447]), .Z(n2863) );
  NANDN U2344 ( .A(n2862), .B(n2863), .Z(n894) );
  AND U2345 ( .A(n895), .B(n894), .Z(n2864) );
  XOR U2346 ( .A(a[448]), .B(b[448]), .Z(n2865) );
  NANDN U2347 ( .A(n2864), .B(n2865), .Z(n896) );
  AND U2348 ( .A(n897), .B(n896), .Z(n2866) );
  XOR U2349 ( .A(a[449]), .B(b[449]), .Z(n2867) );
  NANDN U2350 ( .A(n2866), .B(n2867), .Z(n898) );
  AND U2351 ( .A(n899), .B(n898), .Z(n2870) );
  XOR U2352 ( .A(a[450]), .B(b[450]), .Z(n2871) );
  NANDN U2353 ( .A(n2870), .B(n2871), .Z(n900) );
  AND U2354 ( .A(n901), .B(n900), .Z(n2872) );
  XOR U2355 ( .A(a[451]), .B(b[451]), .Z(n2873) );
  NANDN U2356 ( .A(n2872), .B(n2873), .Z(n902) );
  AND U2357 ( .A(n903), .B(n902), .Z(n2874) );
  XOR U2358 ( .A(a[452]), .B(b[452]), .Z(n2875) );
  NANDN U2359 ( .A(n2874), .B(n2875), .Z(n904) );
  AND U2360 ( .A(n905), .B(n904), .Z(n2876) );
  XOR U2361 ( .A(a[453]), .B(b[453]), .Z(n2877) );
  NANDN U2362 ( .A(n2876), .B(n2877), .Z(n906) );
  AND U2363 ( .A(n907), .B(n906), .Z(n2878) );
  XOR U2364 ( .A(a[454]), .B(b[454]), .Z(n2879) );
  NANDN U2365 ( .A(n2878), .B(n2879), .Z(n908) );
  AND U2366 ( .A(n909), .B(n908), .Z(n2880) );
  XOR U2367 ( .A(a[455]), .B(b[455]), .Z(n2881) );
  NANDN U2368 ( .A(n2880), .B(n2881), .Z(n910) );
  AND U2369 ( .A(n911), .B(n910), .Z(n2882) );
  XOR U2370 ( .A(a[456]), .B(b[456]), .Z(n2883) );
  NANDN U2371 ( .A(n2882), .B(n2883), .Z(n912) );
  AND U2372 ( .A(n913), .B(n912), .Z(n2884) );
  XOR U2373 ( .A(a[457]), .B(b[457]), .Z(n2885) );
  NANDN U2374 ( .A(n2884), .B(n2885), .Z(n914) );
  AND U2375 ( .A(n915), .B(n914), .Z(n2886) );
  XOR U2376 ( .A(a[458]), .B(b[458]), .Z(n2887) );
  NANDN U2377 ( .A(n2886), .B(n2887), .Z(n916) );
  AND U2378 ( .A(n917), .B(n916), .Z(n2888) );
  XOR U2379 ( .A(a[459]), .B(b[459]), .Z(n2889) );
  NANDN U2380 ( .A(n2888), .B(n2889), .Z(n918) );
  AND U2381 ( .A(n919), .B(n918), .Z(n2892) );
  XOR U2382 ( .A(a[460]), .B(b[460]), .Z(n2893) );
  NANDN U2383 ( .A(n2892), .B(n2893), .Z(n920) );
  AND U2384 ( .A(n921), .B(n920), .Z(n2894) );
  XOR U2385 ( .A(a[461]), .B(b[461]), .Z(n2895) );
  NANDN U2386 ( .A(n2894), .B(n2895), .Z(n922) );
  AND U2387 ( .A(n923), .B(n922), .Z(n2896) );
  XOR U2388 ( .A(a[462]), .B(b[462]), .Z(n2897) );
  NANDN U2389 ( .A(n2896), .B(n2897), .Z(n924) );
  AND U2390 ( .A(n925), .B(n924), .Z(n2898) );
  XOR U2391 ( .A(a[463]), .B(b[463]), .Z(n2899) );
  NANDN U2392 ( .A(n2898), .B(n2899), .Z(n926) );
  AND U2393 ( .A(n927), .B(n926), .Z(n2900) );
  XOR U2394 ( .A(a[464]), .B(b[464]), .Z(n2901) );
  NANDN U2395 ( .A(n2900), .B(n2901), .Z(n928) );
  AND U2396 ( .A(n929), .B(n928), .Z(n2902) );
  XOR U2397 ( .A(a[465]), .B(b[465]), .Z(n2903) );
  NANDN U2398 ( .A(n2902), .B(n2903), .Z(n930) );
  AND U2399 ( .A(n931), .B(n930), .Z(n2904) );
  XOR U2400 ( .A(a[466]), .B(b[466]), .Z(n2905) );
  NANDN U2401 ( .A(n2904), .B(n2905), .Z(n932) );
  AND U2402 ( .A(n933), .B(n932), .Z(n2906) );
  XOR U2403 ( .A(a[467]), .B(b[467]), .Z(n2907) );
  NANDN U2404 ( .A(n2906), .B(n2907), .Z(n934) );
  AND U2405 ( .A(n935), .B(n934), .Z(n2908) );
  XOR U2406 ( .A(a[468]), .B(b[468]), .Z(n2909) );
  NANDN U2407 ( .A(n2908), .B(n2909), .Z(n936) );
  AND U2408 ( .A(n937), .B(n936), .Z(n2910) );
  XOR U2409 ( .A(a[469]), .B(b[469]), .Z(n2911) );
  NANDN U2410 ( .A(n2910), .B(n2911), .Z(n938) );
  AND U2411 ( .A(n939), .B(n938), .Z(n2914) );
  XOR U2412 ( .A(a[470]), .B(b[470]), .Z(n2915) );
  NANDN U2413 ( .A(n2914), .B(n2915), .Z(n940) );
  AND U2414 ( .A(n941), .B(n940), .Z(n2916) );
  XOR U2415 ( .A(a[471]), .B(b[471]), .Z(n2917) );
  NANDN U2416 ( .A(n2916), .B(n2917), .Z(n942) );
  AND U2417 ( .A(n943), .B(n942), .Z(n2918) );
  XOR U2418 ( .A(a[472]), .B(b[472]), .Z(n2919) );
  NANDN U2419 ( .A(n2918), .B(n2919), .Z(n944) );
  AND U2420 ( .A(n945), .B(n944), .Z(n2920) );
  XOR U2421 ( .A(a[473]), .B(b[473]), .Z(n2921) );
  NANDN U2422 ( .A(n2920), .B(n2921), .Z(n946) );
  AND U2423 ( .A(n947), .B(n946), .Z(n2922) );
  XOR U2424 ( .A(a[474]), .B(b[474]), .Z(n2923) );
  NANDN U2425 ( .A(n2922), .B(n2923), .Z(n948) );
  AND U2426 ( .A(n949), .B(n948), .Z(n2924) );
  XOR U2427 ( .A(a[475]), .B(b[475]), .Z(n2925) );
  NANDN U2428 ( .A(n2924), .B(n2925), .Z(n950) );
  AND U2429 ( .A(n951), .B(n950), .Z(n2926) );
  XOR U2430 ( .A(a[476]), .B(b[476]), .Z(n2927) );
  NANDN U2431 ( .A(n2926), .B(n2927), .Z(n952) );
  AND U2432 ( .A(n953), .B(n952), .Z(n2928) );
  XOR U2433 ( .A(a[477]), .B(b[477]), .Z(n2929) );
  NANDN U2434 ( .A(n2928), .B(n2929), .Z(n954) );
  AND U2435 ( .A(n955), .B(n954), .Z(n2930) );
  XOR U2436 ( .A(a[478]), .B(b[478]), .Z(n2931) );
  NANDN U2437 ( .A(n2930), .B(n2931), .Z(n956) );
  AND U2438 ( .A(n957), .B(n956), .Z(n2932) );
  XOR U2439 ( .A(a[479]), .B(b[479]), .Z(n2933) );
  NANDN U2440 ( .A(n2932), .B(n2933), .Z(n958) );
  AND U2441 ( .A(n959), .B(n958), .Z(n2936) );
  XOR U2442 ( .A(a[480]), .B(b[480]), .Z(n2937) );
  NANDN U2443 ( .A(n2936), .B(n2937), .Z(n960) );
  AND U2444 ( .A(n961), .B(n960), .Z(n2938) );
  XOR U2445 ( .A(a[481]), .B(b[481]), .Z(n2939) );
  NANDN U2446 ( .A(n2938), .B(n2939), .Z(n962) );
  AND U2447 ( .A(n963), .B(n962), .Z(n2940) );
  XOR U2448 ( .A(a[482]), .B(b[482]), .Z(n2941) );
  NANDN U2449 ( .A(n2940), .B(n2941), .Z(n964) );
  AND U2450 ( .A(n965), .B(n964), .Z(n2942) );
  XOR U2451 ( .A(a[483]), .B(b[483]), .Z(n2943) );
  NANDN U2452 ( .A(n2942), .B(n2943), .Z(n966) );
  AND U2453 ( .A(n967), .B(n966), .Z(n2944) );
  XOR U2454 ( .A(a[484]), .B(b[484]), .Z(n2945) );
  NANDN U2455 ( .A(n2944), .B(n2945), .Z(n968) );
  AND U2456 ( .A(n969), .B(n968), .Z(n2946) );
  XOR U2457 ( .A(a[485]), .B(b[485]), .Z(n2947) );
  NANDN U2458 ( .A(n2946), .B(n2947), .Z(n970) );
  AND U2459 ( .A(n971), .B(n970), .Z(n2948) );
  XOR U2460 ( .A(a[486]), .B(b[486]), .Z(n2949) );
  NANDN U2461 ( .A(n2948), .B(n2949), .Z(n972) );
  AND U2462 ( .A(n973), .B(n972), .Z(n2950) );
  XOR U2463 ( .A(a[487]), .B(b[487]), .Z(n2951) );
  NANDN U2464 ( .A(n2950), .B(n2951), .Z(n974) );
  AND U2465 ( .A(n975), .B(n974), .Z(n2952) );
  XOR U2466 ( .A(a[488]), .B(b[488]), .Z(n2953) );
  NANDN U2467 ( .A(n2952), .B(n2953), .Z(n976) );
  AND U2468 ( .A(n977), .B(n976), .Z(n2954) );
  XOR U2469 ( .A(a[489]), .B(b[489]), .Z(n2955) );
  NANDN U2470 ( .A(n2954), .B(n2955), .Z(n978) );
  AND U2471 ( .A(n979), .B(n978), .Z(n2958) );
  XOR U2472 ( .A(a[490]), .B(b[490]), .Z(n2959) );
  NANDN U2473 ( .A(n2958), .B(n2959), .Z(n980) );
  AND U2474 ( .A(n981), .B(n980), .Z(n2960) );
  XOR U2475 ( .A(a[491]), .B(b[491]), .Z(n2961) );
  NANDN U2476 ( .A(n2960), .B(n2961), .Z(n982) );
  AND U2477 ( .A(n983), .B(n982), .Z(n2962) );
  XOR U2478 ( .A(a[492]), .B(b[492]), .Z(n2963) );
  NANDN U2479 ( .A(n2962), .B(n2963), .Z(n984) );
  AND U2480 ( .A(n985), .B(n984), .Z(n2964) );
  XOR U2481 ( .A(a[493]), .B(b[493]), .Z(n2965) );
  NANDN U2482 ( .A(n2964), .B(n2965), .Z(n986) );
  AND U2483 ( .A(n987), .B(n986), .Z(n2966) );
  XOR U2484 ( .A(a[494]), .B(b[494]), .Z(n2967) );
  NANDN U2485 ( .A(n2966), .B(n2967), .Z(n988) );
  AND U2486 ( .A(n989), .B(n988), .Z(n2968) );
  XOR U2487 ( .A(a[495]), .B(b[495]), .Z(n2969) );
  NANDN U2488 ( .A(n2968), .B(n2969), .Z(n990) );
  AND U2489 ( .A(n991), .B(n990), .Z(n2970) );
  XOR U2490 ( .A(a[496]), .B(b[496]), .Z(n2971) );
  NANDN U2491 ( .A(n2970), .B(n2971), .Z(n992) );
  AND U2492 ( .A(n993), .B(n992), .Z(n2972) );
  XOR U2493 ( .A(a[497]), .B(b[497]), .Z(n2973) );
  NANDN U2494 ( .A(n2972), .B(n2973), .Z(n994) );
  AND U2495 ( .A(n995), .B(n994), .Z(n2974) );
  XOR U2496 ( .A(a[498]), .B(b[498]), .Z(n2975) );
  NANDN U2497 ( .A(n2974), .B(n2975), .Z(n996) );
  AND U2498 ( .A(n997), .B(n996), .Z(n2976) );
  XOR U2499 ( .A(a[499]), .B(b[499]), .Z(n2977) );
  NANDN U2500 ( .A(n2976), .B(n2977), .Z(n998) );
  AND U2501 ( .A(n999), .B(n998), .Z(n2982) );
  XOR U2502 ( .A(a[500]), .B(b[500]), .Z(n2983) );
  NANDN U2503 ( .A(n2982), .B(n2983), .Z(n1000) );
  AND U2504 ( .A(n1001), .B(n1000), .Z(n2984) );
  XOR U2505 ( .A(a[501]), .B(b[501]), .Z(n2985) );
  NANDN U2506 ( .A(n2984), .B(n2985), .Z(n1002) );
  AND U2507 ( .A(n1003), .B(n1002), .Z(n2986) );
  XOR U2508 ( .A(a[502]), .B(b[502]), .Z(n2987) );
  NANDN U2509 ( .A(n2986), .B(n2987), .Z(n1004) );
  AND U2510 ( .A(n1005), .B(n1004), .Z(n2988) );
  XOR U2511 ( .A(a[503]), .B(b[503]), .Z(n2989) );
  NANDN U2512 ( .A(n2988), .B(n2989), .Z(n1006) );
  AND U2513 ( .A(n1007), .B(n1006), .Z(n2990) );
  XOR U2514 ( .A(a[504]), .B(b[504]), .Z(n2991) );
  NANDN U2515 ( .A(n2990), .B(n2991), .Z(n1008) );
  AND U2516 ( .A(n1009), .B(n1008), .Z(n2992) );
  XOR U2517 ( .A(a[505]), .B(b[505]), .Z(n2993) );
  NANDN U2518 ( .A(n2992), .B(n2993), .Z(n1010) );
  AND U2519 ( .A(n1011), .B(n1010), .Z(n2994) );
  XOR U2520 ( .A(a[506]), .B(b[506]), .Z(n2995) );
  NANDN U2521 ( .A(n2994), .B(n2995), .Z(n1012) );
  AND U2522 ( .A(n1013), .B(n1012), .Z(n2996) );
  XOR U2523 ( .A(a[507]), .B(b[507]), .Z(n2997) );
  NANDN U2524 ( .A(n2996), .B(n2997), .Z(n1014) );
  AND U2525 ( .A(n1015), .B(n1014), .Z(n2998) );
  XOR U2526 ( .A(a[508]), .B(b[508]), .Z(n2999) );
  NANDN U2527 ( .A(n2998), .B(n2999), .Z(n1016) );
  AND U2528 ( .A(n1017), .B(n1016), .Z(n3000) );
  XOR U2529 ( .A(a[509]), .B(b[509]), .Z(n3001) );
  NANDN U2530 ( .A(n3000), .B(n3001), .Z(n1018) );
  AND U2531 ( .A(n1019), .B(n1018), .Z(n3004) );
  XOR U2532 ( .A(a[510]), .B(b[510]), .Z(n3005) );
  NANDN U2533 ( .A(n3004), .B(n3005), .Z(n1020) );
  AND U2534 ( .A(n1021), .B(n1020), .Z(n3006) );
  XOR U2535 ( .A(a[511]), .B(b[511]), .Z(n3007) );
  NANDN U2536 ( .A(n3006), .B(n3007), .Z(n1022) );
  AND U2537 ( .A(n1023), .B(n1022), .Z(n3008) );
  XOR U2538 ( .A(a[512]), .B(b[512]), .Z(n3009) );
  NANDN U2539 ( .A(n3008), .B(n3009), .Z(n1024) );
  AND U2540 ( .A(n1025), .B(n1024), .Z(n3010) );
  XOR U2541 ( .A(a[513]), .B(b[513]), .Z(n3011) );
  NANDN U2542 ( .A(n3010), .B(n3011), .Z(n1026) );
  AND U2543 ( .A(n1027), .B(n1026), .Z(n3012) );
  XOR U2544 ( .A(a[514]), .B(b[514]), .Z(n3013) );
  NANDN U2545 ( .A(n3012), .B(n3013), .Z(n1028) );
  AND U2546 ( .A(n1029), .B(n1028), .Z(n3014) );
  XOR U2547 ( .A(a[515]), .B(b[515]), .Z(n3015) );
  NANDN U2548 ( .A(n3014), .B(n3015), .Z(n1030) );
  AND U2549 ( .A(n1031), .B(n1030), .Z(n3016) );
  XOR U2550 ( .A(a[516]), .B(b[516]), .Z(n3017) );
  NANDN U2551 ( .A(n3016), .B(n3017), .Z(n1032) );
  AND U2552 ( .A(n1033), .B(n1032), .Z(n3018) );
  XOR U2553 ( .A(a[517]), .B(b[517]), .Z(n3019) );
  NANDN U2554 ( .A(n3018), .B(n3019), .Z(n1034) );
  AND U2555 ( .A(n1035), .B(n1034), .Z(n3020) );
  XOR U2556 ( .A(a[518]), .B(b[518]), .Z(n3021) );
  NANDN U2557 ( .A(n3020), .B(n3021), .Z(n1036) );
  AND U2558 ( .A(n1037), .B(n1036), .Z(n3022) );
  XOR U2559 ( .A(a[519]), .B(b[519]), .Z(n3023) );
  NANDN U2560 ( .A(n3022), .B(n3023), .Z(n1038) );
  AND U2561 ( .A(n1039), .B(n1038), .Z(n3026) );
  XOR U2562 ( .A(a[520]), .B(b[520]), .Z(n3027) );
  NANDN U2563 ( .A(n3026), .B(n3027), .Z(n1040) );
  AND U2564 ( .A(n1041), .B(n1040), .Z(n3028) );
  XOR U2565 ( .A(a[521]), .B(b[521]), .Z(n3029) );
  NANDN U2566 ( .A(n3028), .B(n3029), .Z(n1042) );
  AND U2567 ( .A(n1043), .B(n1042), .Z(n3030) );
  XOR U2568 ( .A(a[522]), .B(b[522]), .Z(n3031) );
  NANDN U2569 ( .A(n3030), .B(n3031), .Z(n1044) );
  AND U2570 ( .A(n1045), .B(n1044), .Z(n3032) );
  XOR U2571 ( .A(a[523]), .B(b[523]), .Z(n3033) );
  NANDN U2572 ( .A(n3032), .B(n3033), .Z(n1046) );
  AND U2573 ( .A(n1047), .B(n1046), .Z(n3034) );
  XOR U2574 ( .A(a[524]), .B(b[524]), .Z(n3035) );
  NANDN U2575 ( .A(n3034), .B(n3035), .Z(n1048) );
  AND U2576 ( .A(n1049), .B(n1048), .Z(n3036) );
  XOR U2577 ( .A(a[525]), .B(b[525]), .Z(n3037) );
  NANDN U2578 ( .A(n3036), .B(n3037), .Z(n1050) );
  AND U2579 ( .A(n1051), .B(n1050), .Z(n3038) );
  XOR U2580 ( .A(a[526]), .B(b[526]), .Z(n3039) );
  NANDN U2581 ( .A(n3038), .B(n3039), .Z(n1052) );
  AND U2582 ( .A(n1053), .B(n1052), .Z(n3040) );
  XOR U2583 ( .A(a[527]), .B(b[527]), .Z(n3041) );
  NANDN U2584 ( .A(n3040), .B(n3041), .Z(n1054) );
  AND U2585 ( .A(n1055), .B(n1054), .Z(n3042) );
  XOR U2586 ( .A(a[528]), .B(b[528]), .Z(n3043) );
  NANDN U2587 ( .A(n3042), .B(n3043), .Z(n1056) );
  AND U2588 ( .A(n1057), .B(n1056), .Z(n3044) );
  XOR U2589 ( .A(a[529]), .B(b[529]), .Z(n3045) );
  NANDN U2590 ( .A(n3044), .B(n3045), .Z(n1058) );
  AND U2591 ( .A(n1059), .B(n1058), .Z(n3048) );
  XOR U2592 ( .A(a[530]), .B(b[530]), .Z(n3049) );
  NANDN U2593 ( .A(n3048), .B(n3049), .Z(n1060) );
  AND U2594 ( .A(n1061), .B(n1060), .Z(n3050) );
  XOR U2595 ( .A(a[531]), .B(b[531]), .Z(n3051) );
  NANDN U2596 ( .A(n3050), .B(n3051), .Z(n1062) );
  AND U2597 ( .A(n1063), .B(n1062), .Z(n3052) );
  XOR U2598 ( .A(a[532]), .B(b[532]), .Z(n3053) );
  NANDN U2599 ( .A(n3052), .B(n3053), .Z(n1064) );
  AND U2600 ( .A(n1065), .B(n1064), .Z(n3054) );
  XOR U2601 ( .A(a[533]), .B(b[533]), .Z(n3055) );
  NANDN U2602 ( .A(n3054), .B(n3055), .Z(n1066) );
  AND U2603 ( .A(n1067), .B(n1066), .Z(n3056) );
  XOR U2604 ( .A(a[534]), .B(b[534]), .Z(n3057) );
  NANDN U2605 ( .A(n3056), .B(n3057), .Z(n1068) );
  AND U2606 ( .A(n1069), .B(n1068), .Z(n3058) );
  XOR U2607 ( .A(a[535]), .B(b[535]), .Z(n3059) );
  NANDN U2608 ( .A(n3058), .B(n3059), .Z(n1070) );
  AND U2609 ( .A(n1071), .B(n1070), .Z(n3060) );
  XOR U2610 ( .A(a[536]), .B(b[536]), .Z(n3061) );
  NANDN U2611 ( .A(n3060), .B(n3061), .Z(n1072) );
  AND U2612 ( .A(n1073), .B(n1072), .Z(n3062) );
  XOR U2613 ( .A(a[537]), .B(b[537]), .Z(n3063) );
  NANDN U2614 ( .A(n3062), .B(n3063), .Z(n1074) );
  AND U2615 ( .A(n1075), .B(n1074), .Z(n3064) );
  XOR U2616 ( .A(a[538]), .B(b[538]), .Z(n3065) );
  NANDN U2617 ( .A(n3064), .B(n3065), .Z(n1076) );
  AND U2618 ( .A(n1077), .B(n1076), .Z(n3066) );
  XOR U2619 ( .A(a[539]), .B(b[539]), .Z(n3067) );
  NANDN U2620 ( .A(n3066), .B(n3067), .Z(n1078) );
  AND U2621 ( .A(n1079), .B(n1078), .Z(n3070) );
  XOR U2622 ( .A(a[540]), .B(b[540]), .Z(n3071) );
  NANDN U2623 ( .A(n3070), .B(n3071), .Z(n1080) );
  AND U2624 ( .A(n1081), .B(n1080), .Z(n3072) );
  XOR U2625 ( .A(a[541]), .B(b[541]), .Z(n3073) );
  NANDN U2626 ( .A(n3072), .B(n3073), .Z(n1082) );
  AND U2627 ( .A(n1083), .B(n1082), .Z(n3074) );
  XOR U2628 ( .A(a[542]), .B(b[542]), .Z(n3075) );
  NANDN U2629 ( .A(n3074), .B(n3075), .Z(n1084) );
  AND U2630 ( .A(n1085), .B(n1084), .Z(n3076) );
  XOR U2631 ( .A(a[543]), .B(b[543]), .Z(n3077) );
  NANDN U2632 ( .A(n3076), .B(n3077), .Z(n1086) );
  AND U2633 ( .A(n1087), .B(n1086), .Z(n3078) );
  XOR U2634 ( .A(a[544]), .B(b[544]), .Z(n3079) );
  NANDN U2635 ( .A(n3078), .B(n3079), .Z(n1088) );
  AND U2636 ( .A(n1089), .B(n1088), .Z(n3080) );
  XOR U2637 ( .A(a[545]), .B(b[545]), .Z(n3081) );
  NANDN U2638 ( .A(n3080), .B(n3081), .Z(n1090) );
  AND U2639 ( .A(n1091), .B(n1090), .Z(n3082) );
  XOR U2640 ( .A(a[546]), .B(b[546]), .Z(n3083) );
  NANDN U2641 ( .A(n3082), .B(n3083), .Z(n1092) );
  AND U2642 ( .A(n1093), .B(n1092), .Z(n3084) );
  XOR U2643 ( .A(a[547]), .B(b[547]), .Z(n3085) );
  NANDN U2644 ( .A(n3084), .B(n3085), .Z(n1094) );
  AND U2645 ( .A(n1095), .B(n1094), .Z(n3086) );
  XOR U2646 ( .A(a[548]), .B(b[548]), .Z(n3087) );
  NANDN U2647 ( .A(n3086), .B(n3087), .Z(n1096) );
  AND U2648 ( .A(n1097), .B(n1096), .Z(n3088) );
  XOR U2649 ( .A(a[549]), .B(b[549]), .Z(n3089) );
  NANDN U2650 ( .A(n3088), .B(n3089), .Z(n1098) );
  AND U2651 ( .A(n1099), .B(n1098), .Z(n3092) );
  XOR U2652 ( .A(a[550]), .B(b[550]), .Z(n3093) );
  NANDN U2653 ( .A(n3092), .B(n3093), .Z(n1100) );
  AND U2654 ( .A(n1101), .B(n1100), .Z(n3094) );
  XOR U2655 ( .A(a[551]), .B(b[551]), .Z(n3095) );
  NANDN U2656 ( .A(n3094), .B(n3095), .Z(n1102) );
  AND U2657 ( .A(n1103), .B(n1102), .Z(n3096) );
  XOR U2658 ( .A(a[552]), .B(b[552]), .Z(n3097) );
  NANDN U2659 ( .A(n3096), .B(n3097), .Z(n1104) );
  AND U2660 ( .A(n1105), .B(n1104), .Z(n3098) );
  XOR U2661 ( .A(a[553]), .B(b[553]), .Z(n3099) );
  NANDN U2662 ( .A(n3098), .B(n3099), .Z(n1106) );
  AND U2663 ( .A(n1107), .B(n1106), .Z(n3100) );
  XOR U2664 ( .A(a[554]), .B(b[554]), .Z(n3101) );
  NANDN U2665 ( .A(n3100), .B(n3101), .Z(n1108) );
  AND U2666 ( .A(n1109), .B(n1108), .Z(n3102) );
  XOR U2667 ( .A(a[555]), .B(b[555]), .Z(n3103) );
  NANDN U2668 ( .A(n3102), .B(n3103), .Z(n1110) );
  AND U2669 ( .A(n1111), .B(n1110), .Z(n3104) );
  XOR U2670 ( .A(a[556]), .B(b[556]), .Z(n3105) );
  NANDN U2671 ( .A(n3104), .B(n3105), .Z(n1112) );
  AND U2672 ( .A(n1113), .B(n1112), .Z(n3106) );
  XOR U2673 ( .A(a[557]), .B(b[557]), .Z(n3107) );
  NANDN U2674 ( .A(n3106), .B(n3107), .Z(n1114) );
  AND U2675 ( .A(n1115), .B(n1114), .Z(n3108) );
  XOR U2676 ( .A(a[558]), .B(b[558]), .Z(n3109) );
  NANDN U2677 ( .A(n3108), .B(n3109), .Z(n1116) );
  AND U2678 ( .A(n1117), .B(n1116), .Z(n3110) );
  XOR U2679 ( .A(a[559]), .B(b[559]), .Z(n3111) );
  NANDN U2680 ( .A(n3110), .B(n3111), .Z(n1118) );
  AND U2681 ( .A(n1119), .B(n1118), .Z(n3114) );
  XOR U2682 ( .A(a[560]), .B(b[560]), .Z(n3115) );
  NANDN U2683 ( .A(n3114), .B(n3115), .Z(n1120) );
  AND U2684 ( .A(n1121), .B(n1120), .Z(n3116) );
  XOR U2685 ( .A(a[561]), .B(b[561]), .Z(n3117) );
  NANDN U2686 ( .A(n3116), .B(n3117), .Z(n1122) );
  AND U2687 ( .A(n1123), .B(n1122), .Z(n3118) );
  XOR U2688 ( .A(a[562]), .B(b[562]), .Z(n3119) );
  NANDN U2689 ( .A(n3118), .B(n3119), .Z(n1124) );
  AND U2690 ( .A(n1125), .B(n1124), .Z(n3120) );
  XOR U2691 ( .A(a[563]), .B(b[563]), .Z(n3121) );
  NANDN U2692 ( .A(n3120), .B(n3121), .Z(n1126) );
  AND U2693 ( .A(n1127), .B(n1126), .Z(n3122) );
  XOR U2694 ( .A(a[564]), .B(b[564]), .Z(n3123) );
  NANDN U2695 ( .A(n3122), .B(n3123), .Z(n1128) );
  AND U2696 ( .A(n1129), .B(n1128), .Z(n3124) );
  XOR U2697 ( .A(a[565]), .B(b[565]), .Z(n3125) );
  NANDN U2698 ( .A(n3124), .B(n3125), .Z(n1130) );
  AND U2699 ( .A(n1131), .B(n1130), .Z(n3126) );
  XOR U2700 ( .A(a[566]), .B(b[566]), .Z(n3127) );
  NANDN U2701 ( .A(n3126), .B(n3127), .Z(n1132) );
  AND U2702 ( .A(n1133), .B(n1132), .Z(n3128) );
  XOR U2703 ( .A(a[567]), .B(b[567]), .Z(n3129) );
  NANDN U2704 ( .A(n3128), .B(n3129), .Z(n1134) );
  AND U2705 ( .A(n1135), .B(n1134), .Z(n3130) );
  XOR U2706 ( .A(a[568]), .B(b[568]), .Z(n3131) );
  NANDN U2707 ( .A(n3130), .B(n3131), .Z(n1136) );
  AND U2708 ( .A(n1137), .B(n1136), .Z(n3132) );
  XOR U2709 ( .A(a[569]), .B(b[569]), .Z(n3133) );
  NANDN U2710 ( .A(n3132), .B(n3133), .Z(n1138) );
  AND U2711 ( .A(n1139), .B(n1138), .Z(n3136) );
  XOR U2712 ( .A(a[570]), .B(b[570]), .Z(n3137) );
  NANDN U2713 ( .A(n3136), .B(n3137), .Z(n1140) );
  AND U2714 ( .A(n1141), .B(n1140), .Z(n3138) );
  XOR U2715 ( .A(a[571]), .B(b[571]), .Z(n3139) );
  NANDN U2716 ( .A(n3138), .B(n3139), .Z(n1142) );
  AND U2717 ( .A(n1143), .B(n1142), .Z(n3140) );
  XOR U2718 ( .A(a[572]), .B(b[572]), .Z(n3141) );
  NANDN U2719 ( .A(n3140), .B(n3141), .Z(n1144) );
  AND U2720 ( .A(n1145), .B(n1144), .Z(n3142) );
  XOR U2721 ( .A(a[573]), .B(b[573]), .Z(n3143) );
  NANDN U2722 ( .A(n3142), .B(n3143), .Z(n1146) );
  AND U2723 ( .A(n1147), .B(n1146), .Z(n3144) );
  XOR U2724 ( .A(a[574]), .B(b[574]), .Z(n3145) );
  NANDN U2725 ( .A(n3144), .B(n3145), .Z(n1148) );
  AND U2726 ( .A(n1149), .B(n1148), .Z(n3146) );
  XOR U2727 ( .A(a[575]), .B(b[575]), .Z(n3147) );
  NANDN U2728 ( .A(n3146), .B(n3147), .Z(n1150) );
  AND U2729 ( .A(n1151), .B(n1150), .Z(n3148) );
  XOR U2730 ( .A(a[576]), .B(b[576]), .Z(n3149) );
  NANDN U2731 ( .A(n3148), .B(n3149), .Z(n1152) );
  AND U2732 ( .A(n1153), .B(n1152), .Z(n3150) );
  XOR U2733 ( .A(a[577]), .B(b[577]), .Z(n3151) );
  NANDN U2734 ( .A(n3150), .B(n3151), .Z(n1154) );
  AND U2735 ( .A(n1155), .B(n1154), .Z(n3152) );
  XOR U2736 ( .A(a[578]), .B(b[578]), .Z(n3153) );
  NANDN U2737 ( .A(n3152), .B(n3153), .Z(n1156) );
  AND U2738 ( .A(n1157), .B(n1156), .Z(n3154) );
  XOR U2739 ( .A(a[579]), .B(b[579]), .Z(n3155) );
  NANDN U2740 ( .A(n3154), .B(n3155), .Z(n1158) );
  AND U2741 ( .A(n1159), .B(n1158), .Z(n3158) );
  XOR U2742 ( .A(a[580]), .B(b[580]), .Z(n3159) );
  NANDN U2743 ( .A(n3158), .B(n3159), .Z(n1160) );
  AND U2744 ( .A(n1161), .B(n1160), .Z(n3160) );
  XOR U2745 ( .A(a[581]), .B(b[581]), .Z(n3161) );
  NANDN U2746 ( .A(n3160), .B(n3161), .Z(n1162) );
  AND U2747 ( .A(n1163), .B(n1162), .Z(n3162) );
  XOR U2748 ( .A(a[582]), .B(b[582]), .Z(n3163) );
  NANDN U2749 ( .A(n3162), .B(n3163), .Z(n1164) );
  AND U2750 ( .A(n1165), .B(n1164), .Z(n3164) );
  XOR U2751 ( .A(a[583]), .B(b[583]), .Z(n3165) );
  NANDN U2752 ( .A(n3164), .B(n3165), .Z(n1166) );
  AND U2753 ( .A(n1167), .B(n1166), .Z(n3166) );
  XOR U2754 ( .A(a[584]), .B(b[584]), .Z(n3167) );
  NANDN U2755 ( .A(n3166), .B(n3167), .Z(n1168) );
  AND U2756 ( .A(n1169), .B(n1168), .Z(n3168) );
  XOR U2757 ( .A(a[585]), .B(b[585]), .Z(n3169) );
  NANDN U2758 ( .A(n3168), .B(n3169), .Z(n1170) );
  AND U2759 ( .A(n1171), .B(n1170), .Z(n3170) );
  XOR U2760 ( .A(a[586]), .B(b[586]), .Z(n3171) );
  NANDN U2761 ( .A(n3170), .B(n3171), .Z(n1172) );
  AND U2762 ( .A(n1173), .B(n1172), .Z(n3172) );
  XOR U2763 ( .A(a[587]), .B(b[587]), .Z(n3173) );
  NANDN U2764 ( .A(n3172), .B(n3173), .Z(n1174) );
  AND U2765 ( .A(n1175), .B(n1174), .Z(n3174) );
  XOR U2766 ( .A(a[588]), .B(b[588]), .Z(n3175) );
  NANDN U2767 ( .A(n3174), .B(n3175), .Z(n1176) );
  AND U2768 ( .A(n1177), .B(n1176), .Z(n3176) );
  XOR U2769 ( .A(a[589]), .B(b[589]), .Z(n3177) );
  NANDN U2770 ( .A(n3176), .B(n3177), .Z(n1178) );
  AND U2771 ( .A(n1179), .B(n1178), .Z(n3180) );
  XOR U2772 ( .A(a[590]), .B(b[590]), .Z(n3181) );
  NANDN U2773 ( .A(n3180), .B(n3181), .Z(n1180) );
  AND U2774 ( .A(n1181), .B(n1180), .Z(n3182) );
  XOR U2775 ( .A(a[591]), .B(b[591]), .Z(n3183) );
  NANDN U2776 ( .A(n3182), .B(n3183), .Z(n1182) );
  AND U2777 ( .A(n1183), .B(n1182), .Z(n3184) );
  XOR U2778 ( .A(a[592]), .B(b[592]), .Z(n3185) );
  NANDN U2779 ( .A(n3184), .B(n3185), .Z(n1184) );
  AND U2780 ( .A(n1185), .B(n1184), .Z(n3186) );
  XOR U2781 ( .A(a[593]), .B(b[593]), .Z(n3187) );
  NANDN U2782 ( .A(n3186), .B(n3187), .Z(n1186) );
  AND U2783 ( .A(n1187), .B(n1186), .Z(n3188) );
  XOR U2784 ( .A(a[594]), .B(b[594]), .Z(n3189) );
  NANDN U2785 ( .A(n3188), .B(n3189), .Z(n1188) );
  AND U2786 ( .A(n1189), .B(n1188), .Z(n3190) );
  XOR U2787 ( .A(a[595]), .B(b[595]), .Z(n3191) );
  NANDN U2788 ( .A(n3190), .B(n3191), .Z(n1190) );
  AND U2789 ( .A(n1191), .B(n1190), .Z(n3192) );
  XOR U2790 ( .A(a[596]), .B(b[596]), .Z(n3193) );
  NANDN U2791 ( .A(n3192), .B(n3193), .Z(n1192) );
  AND U2792 ( .A(n1193), .B(n1192), .Z(n3194) );
  XOR U2793 ( .A(a[597]), .B(b[597]), .Z(n3195) );
  NANDN U2794 ( .A(n3194), .B(n3195), .Z(n1194) );
  AND U2795 ( .A(n1195), .B(n1194), .Z(n3196) );
  XOR U2796 ( .A(a[598]), .B(b[598]), .Z(n3197) );
  NANDN U2797 ( .A(n3196), .B(n3197), .Z(n1196) );
  AND U2798 ( .A(n1197), .B(n1196), .Z(n3198) );
  XOR U2799 ( .A(a[599]), .B(b[599]), .Z(n3199) );
  NANDN U2800 ( .A(n3198), .B(n3199), .Z(n1198) );
  AND U2801 ( .A(n1199), .B(n1198), .Z(n3204) );
  XOR U2802 ( .A(a[600]), .B(b[600]), .Z(n3205) );
  NANDN U2803 ( .A(n3204), .B(n3205), .Z(n1200) );
  AND U2804 ( .A(n1201), .B(n1200), .Z(n3206) );
  XOR U2805 ( .A(a[601]), .B(b[601]), .Z(n3207) );
  NANDN U2806 ( .A(n3206), .B(n3207), .Z(n1202) );
  AND U2807 ( .A(n1203), .B(n1202), .Z(n3208) );
  XOR U2808 ( .A(a[602]), .B(b[602]), .Z(n3209) );
  NANDN U2809 ( .A(n3208), .B(n3209), .Z(n1204) );
  AND U2810 ( .A(n1205), .B(n1204), .Z(n3210) );
  XOR U2811 ( .A(a[603]), .B(b[603]), .Z(n3211) );
  NANDN U2812 ( .A(n3210), .B(n3211), .Z(n1206) );
  AND U2813 ( .A(n1207), .B(n1206), .Z(n3212) );
  XOR U2814 ( .A(a[604]), .B(b[604]), .Z(n3213) );
  NANDN U2815 ( .A(n3212), .B(n3213), .Z(n1208) );
  AND U2816 ( .A(n1209), .B(n1208), .Z(n3214) );
  XOR U2817 ( .A(a[605]), .B(b[605]), .Z(n3215) );
  NANDN U2818 ( .A(n3214), .B(n3215), .Z(n1210) );
  AND U2819 ( .A(n1211), .B(n1210), .Z(n3216) );
  XOR U2820 ( .A(a[606]), .B(b[606]), .Z(n3217) );
  NANDN U2821 ( .A(n3216), .B(n3217), .Z(n1212) );
  AND U2822 ( .A(n1213), .B(n1212), .Z(n3218) );
  XOR U2823 ( .A(a[607]), .B(b[607]), .Z(n3219) );
  NANDN U2824 ( .A(n3218), .B(n3219), .Z(n1214) );
  AND U2825 ( .A(n1215), .B(n1214), .Z(n3220) );
  XOR U2826 ( .A(a[608]), .B(b[608]), .Z(n3221) );
  NANDN U2827 ( .A(n3220), .B(n3221), .Z(n1216) );
  AND U2828 ( .A(n1217), .B(n1216), .Z(n3222) );
  XOR U2829 ( .A(a[609]), .B(b[609]), .Z(n3223) );
  NANDN U2830 ( .A(n3222), .B(n3223), .Z(n1218) );
  AND U2831 ( .A(n1219), .B(n1218), .Z(n3226) );
  XOR U2832 ( .A(a[610]), .B(b[610]), .Z(n3227) );
  NANDN U2833 ( .A(n3226), .B(n3227), .Z(n1220) );
  AND U2834 ( .A(n1221), .B(n1220), .Z(n3228) );
  XOR U2835 ( .A(a[611]), .B(b[611]), .Z(n3229) );
  NANDN U2836 ( .A(n3228), .B(n3229), .Z(n1222) );
  AND U2837 ( .A(n1223), .B(n1222), .Z(n3230) );
  XOR U2838 ( .A(a[612]), .B(b[612]), .Z(n3231) );
  NANDN U2839 ( .A(n3230), .B(n3231), .Z(n1224) );
  AND U2840 ( .A(n1225), .B(n1224), .Z(n3232) );
  XOR U2841 ( .A(a[613]), .B(b[613]), .Z(n3233) );
  NANDN U2842 ( .A(n3232), .B(n3233), .Z(n1226) );
  AND U2843 ( .A(n1227), .B(n1226), .Z(n3234) );
  XOR U2844 ( .A(a[614]), .B(b[614]), .Z(n3235) );
  NANDN U2845 ( .A(n3234), .B(n3235), .Z(n1228) );
  AND U2846 ( .A(n1229), .B(n1228), .Z(n3236) );
  XOR U2847 ( .A(a[615]), .B(b[615]), .Z(n3237) );
  NANDN U2848 ( .A(n3236), .B(n3237), .Z(n1230) );
  AND U2849 ( .A(n1231), .B(n1230), .Z(n3238) );
  XOR U2850 ( .A(a[616]), .B(b[616]), .Z(n3239) );
  NANDN U2851 ( .A(n3238), .B(n3239), .Z(n1232) );
  AND U2852 ( .A(n1233), .B(n1232), .Z(n3240) );
  XOR U2853 ( .A(a[617]), .B(b[617]), .Z(n3241) );
  NANDN U2854 ( .A(n3240), .B(n3241), .Z(n1234) );
  AND U2855 ( .A(n1235), .B(n1234), .Z(n3242) );
  XOR U2856 ( .A(a[618]), .B(b[618]), .Z(n3243) );
  NANDN U2857 ( .A(n3242), .B(n3243), .Z(n1236) );
  AND U2858 ( .A(n1237), .B(n1236), .Z(n3244) );
  XOR U2859 ( .A(a[619]), .B(b[619]), .Z(n3245) );
  NANDN U2860 ( .A(n3244), .B(n3245), .Z(n1238) );
  AND U2861 ( .A(n1239), .B(n1238), .Z(n3248) );
  XOR U2862 ( .A(a[620]), .B(b[620]), .Z(n3249) );
  NANDN U2863 ( .A(n3248), .B(n3249), .Z(n1240) );
  AND U2864 ( .A(n1241), .B(n1240), .Z(n3250) );
  XOR U2865 ( .A(a[621]), .B(b[621]), .Z(n3251) );
  NANDN U2866 ( .A(n3250), .B(n3251), .Z(n1242) );
  AND U2867 ( .A(n1243), .B(n1242), .Z(n3252) );
  XOR U2868 ( .A(a[622]), .B(b[622]), .Z(n3253) );
  NANDN U2869 ( .A(n3252), .B(n3253), .Z(n1244) );
  AND U2870 ( .A(n1245), .B(n1244), .Z(n3254) );
  XOR U2871 ( .A(a[623]), .B(b[623]), .Z(n3255) );
  NANDN U2872 ( .A(n3254), .B(n3255), .Z(n1246) );
  AND U2873 ( .A(n1247), .B(n1246), .Z(n3256) );
  XOR U2874 ( .A(a[624]), .B(b[624]), .Z(n3257) );
  NANDN U2875 ( .A(n3256), .B(n3257), .Z(n1248) );
  AND U2876 ( .A(n1249), .B(n1248), .Z(n3258) );
  XOR U2877 ( .A(a[625]), .B(b[625]), .Z(n3259) );
  NANDN U2878 ( .A(n3258), .B(n3259), .Z(n1250) );
  AND U2879 ( .A(n1251), .B(n1250), .Z(n3260) );
  XOR U2880 ( .A(a[626]), .B(b[626]), .Z(n3261) );
  NANDN U2881 ( .A(n3260), .B(n3261), .Z(n1252) );
  AND U2882 ( .A(n1253), .B(n1252), .Z(n3262) );
  XOR U2883 ( .A(a[627]), .B(b[627]), .Z(n3263) );
  NANDN U2884 ( .A(n3262), .B(n3263), .Z(n1254) );
  AND U2885 ( .A(n1255), .B(n1254), .Z(n3264) );
  XOR U2886 ( .A(a[628]), .B(b[628]), .Z(n3265) );
  NANDN U2887 ( .A(n3264), .B(n3265), .Z(n1256) );
  AND U2888 ( .A(n1257), .B(n1256), .Z(n3266) );
  XOR U2889 ( .A(a[629]), .B(b[629]), .Z(n3267) );
  NANDN U2890 ( .A(n3266), .B(n3267), .Z(n1258) );
  AND U2891 ( .A(n1259), .B(n1258), .Z(n3270) );
  XOR U2892 ( .A(a[630]), .B(b[630]), .Z(n3271) );
  NANDN U2893 ( .A(n3270), .B(n3271), .Z(n1260) );
  AND U2894 ( .A(n1261), .B(n1260), .Z(n3272) );
  XOR U2895 ( .A(a[631]), .B(b[631]), .Z(n3273) );
  NANDN U2896 ( .A(n3272), .B(n3273), .Z(n1262) );
  AND U2897 ( .A(n1263), .B(n1262), .Z(n3274) );
  XOR U2898 ( .A(a[632]), .B(b[632]), .Z(n3275) );
  NANDN U2899 ( .A(n3274), .B(n3275), .Z(n1264) );
  AND U2900 ( .A(n1265), .B(n1264), .Z(n3276) );
  XOR U2901 ( .A(a[633]), .B(b[633]), .Z(n3277) );
  NANDN U2902 ( .A(n3276), .B(n3277), .Z(n1266) );
  AND U2903 ( .A(n1267), .B(n1266), .Z(n3278) );
  XOR U2904 ( .A(a[634]), .B(b[634]), .Z(n3279) );
  NANDN U2905 ( .A(n3278), .B(n3279), .Z(n1268) );
  AND U2906 ( .A(n1269), .B(n1268), .Z(n3280) );
  XOR U2907 ( .A(a[635]), .B(b[635]), .Z(n3281) );
  NANDN U2908 ( .A(n3280), .B(n3281), .Z(n1270) );
  AND U2909 ( .A(n1271), .B(n1270), .Z(n3282) );
  XOR U2910 ( .A(a[636]), .B(b[636]), .Z(n3283) );
  NANDN U2911 ( .A(n3282), .B(n3283), .Z(n1272) );
  AND U2912 ( .A(n1273), .B(n1272), .Z(n3284) );
  XOR U2913 ( .A(a[637]), .B(b[637]), .Z(n3285) );
  NANDN U2914 ( .A(n3284), .B(n3285), .Z(n1274) );
  AND U2915 ( .A(n1275), .B(n1274), .Z(n3286) );
  XOR U2916 ( .A(a[638]), .B(b[638]), .Z(n3287) );
  NANDN U2917 ( .A(n3286), .B(n3287), .Z(n1276) );
  AND U2918 ( .A(n1277), .B(n1276), .Z(n3288) );
  XOR U2919 ( .A(a[639]), .B(b[639]), .Z(n3289) );
  NANDN U2920 ( .A(n3288), .B(n3289), .Z(n1278) );
  AND U2921 ( .A(n1279), .B(n1278), .Z(n3292) );
  XOR U2922 ( .A(a[640]), .B(b[640]), .Z(n3293) );
  NANDN U2923 ( .A(n3292), .B(n3293), .Z(n1280) );
  AND U2924 ( .A(n1281), .B(n1280), .Z(n3294) );
  XOR U2925 ( .A(a[641]), .B(b[641]), .Z(n3295) );
  NANDN U2926 ( .A(n3294), .B(n3295), .Z(n1282) );
  AND U2927 ( .A(n1283), .B(n1282), .Z(n3296) );
  XOR U2928 ( .A(a[642]), .B(b[642]), .Z(n3297) );
  NANDN U2929 ( .A(n3296), .B(n3297), .Z(n1284) );
  AND U2930 ( .A(n1285), .B(n1284), .Z(n3298) );
  XOR U2931 ( .A(a[643]), .B(b[643]), .Z(n3299) );
  NANDN U2932 ( .A(n3298), .B(n3299), .Z(n1286) );
  AND U2933 ( .A(n1287), .B(n1286), .Z(n3300) );
  XOR U2934 ( .A(a[644]), .B(b[644]), .Z(n3301) );
  NANDN U2935 ( .A(n3300), .B(n3301), .Z(n1288) );
  AND U2936 ( .A(n1289), .B(n1288), .Z(n3302) );
  XOR U2937 ( .A(a[645]), .B(b[645]), .Z(n3303) );
  NANDN U2938 ( .A(n3302), .B(n3303), .Z(n1290) );
  AND U2939 ( .A(n1291), .B(n1290), .Z(n3304) );
  XOR U2940 ( .A(a[646]), .B(b[646]), .Z(n3305) );
  NANDN U2941 ( .A(n3304), .B(n3305), .Z(n1292) );
  AND U2942 ( .A(n1293), .B(n1292), .Z(n3306) );
  XOR U2943 ( .A(a[647]), .B(b[647]), .Z(n3307) );
  NANDN U2944 ( .A(n3306), .B(n3307), .Z(n1294) );
  AND U2945 ( .A(n1295), .B(n1294), .Z(n3308) );
  XOR U2946 ( .A(a[648]), .B(b[648]), .Z(n3309) );
  NANDN U2947 ( .A(n3308), .B(n3309), .Z(n1296) );
  AND U2948 ( .A(n1297), .B(n1296), .Z(n3310) );
  XOR U2949 ( .A(a[649]), .B(b[649]), .Z(n3311) );
  NANDN U2950 ( .A(n3310), .B(n3311), .Z(n1298) );
  AND U2951 ( .A(n1299), .B(n1298), .Z(n3314) );
  XOR U2952 ( .A(a[650]), .B(b[650]), .Z(n3315) );
  NANDN U2953 ( .A(n3314), .B(n3315), .Z(n1300) );
  AND U2954 ( .A(n1301), .B(n1300), .Z(n3316) );
  XOR U2955 ( .A(a[651]), .B(b[651]), .Z(n3317) );
  NANDN U2956 ( .A(n3316), .B(n3317), .Z(n1302) );
  AND U2957 ( .A(n1303), .B(n1302), .Z(n3318) );
  XOR U2958 ( .A(a[652]), .B(b[652]), .Z(n3319) );
  NANDN U2959 ( .A(n3318), .B(n3319), .Z(n1304) );
  AND U2960 ( .A(n1305), .B(n1304), .Z(n3320) );
  XOR U2961 ( .A(a[653]), .B(b[653]), .Z(n3321) );
  NANDN U2962 ( .A(n3320), .B(n3321), .Z(n1306) );
  AND U2963 ( .A(n1307), .B(n1306), .Z(n3322) );
  XOR U2964 ( .A(a[654]), .B(b[654]), .Z(n3323) );
  NANDN U2965 ( .A(n3322), .B(n3323), .Z(n1308) );
  AND U2966 ( .A(n1309), .B(n1308), .Z(n3324) );
  XOR U2967 ( .A(a[655]), .B(b[655]), .Z(n3325) );
  NANDN U2968 ( .A(n3324), .B(n3325), .Z(n1310) );
  AND U2969 ( .A(n1311), .B(n1310), .Z(n3326) );
  XOR U2970 ( .A(a[656]), .B(b[656]), .Z(n3327) );
  NANDN U2971 ( .A(n3326), .B(n3327), .Z(n1312) );
  AND U2972 ( .A(n1313), .B(n1312), .Z(n3328) );
  XOR U2973 ( .A(a[657]), .B(b[657]), .Z(n3329) );
  NANDN U2974 ( .A(n3328), .B(n3329), .Z(n1314) );
  AND U2975 ( .A(n1315), .B(n1314), .Z(n3330) );
  XOR U2976 ( .A(a[658]), .B(b[658]), .Z(n3331) );
  NANDN U2977 ( .A(n3330), .B(n3331), .Z(n1316) );
  AND U2978 ( .A(n1317), .B(n1316), .Z(n3332) );
  XOR U2979 ( .A(a[659]), .B(b[659]), .Z(n3333) );
  NANDN U2980 ( .A(n3332), .B(n3333), .Z(n1318) );
  AND U2981 ( .A(n1319), .B(n1318), .Z(n3336) );
  XOR U2982 ( .A(a[660]), .B(b[660]), .Z(n3337) );
  NANDN U2983 ( .A(n3336), .B(n3337), .Z(n1320) );
  AND U2984 ( .A(n1321), .B(n1320), .Z(n3338) );
  XOR U2985 ( .A(a[661]), .B(b[661]), .Z(n3339) );
  NANDN U2986 ( .A(n3338), .B(n3339), .Z(n1322) );
  AND U2987 ( .A(n1323), .B(n1322), .Z(n3340) );
  XOR U2988 ( .A(a[662]), .B(b[662]), .Z(n3341) );
  NANDN U2989 ( .A(n3340), .B(n3341), .Z(n1324) );
  AND U2990 ( .A(n1325), .B(n1324), .Z(n3342) );
  XOR U2991 ( .A(a[663]), .B(b[663]), .Z(n3343) );
  NANDN U2992 ( .A(n3342), .B(n3343), .Z(n1326) );
  AND U2993 ( .A(n1327), .B(n1326), .Z(n3344) );
  XOR U2994 ( .A(a[664]), .B(b[664]), .Z(n3345) );
  NANDN U2995 ( .A(n3344), .B(n3345), .Z(n1328) );
  AND U2996 ( .A(n1329), .B(n1328), .Z(n3346) );
  XOR U2997 ( .A(a[665]), .B(b[665]), .Z(n3347) );
  NANDN U2998 ( .A(n3346), .B(n3347), .Z(n1330) );
  AND U2999 ( .A(n1331), .B(n1330), .Z(n3348) );
  XOR U3000 ( .A(a[666]), .B(b[666]), .Z(n3349) );
  NANDN U3001 ( .A(n3348), .B(n3349), .Z(n1332) );
  AND U3002 ( .A(n1333), .B(n1332), .Z(n3350) );
  XOR U3003 ( .A(a[667]), .B(b[667]), .Z(n3351) );
  NANDN U3004 ( .A(n3350), .B(n3351), .Z(n1334) );
  AND U3005 ( .A(n1335), .B(n1334), .Z(n3352) );
  XOR U3006 ( .A(a[668]), .B(b[668]), .Z(n3353) );
  NANDN U3007 ( .A(n3352), .B(n3353), .Z(n1336) );
  AND U3008 ( .A(n1337), .B(n1336), .Z(n3354) );
  XOR U3009 ( .A(a[669]), .B(b[669]), .Z(n3355) );
  NANDN U3010 ( .A(n3354), .B(n3355), .Z(n1338) );
  AND U3011 ( .A(n1339), .B(n1338), .Z(n3358) );
  XOR U3012 ( .A(a[670]), .B(b[670]), .Z(n3359) );
  NANDN U3013 ( .A(n3358), .B(n3359), .Z(n1340) );
  AND U3014 ( .A(n1341), .B(n1340), .Z(n3360) );
  XOR U3015 ( .A(a[671]), .B(b[671]), .Z(n3361) );
  NANDN U3016 ( .A(n3360), .B(n3361), .Z(n1342) );
  AND U3017 ( .A(n1343), .B(n1342), .Z(n3362) );
  XOR U3018 ( .A(a[672]), .B(b[672]), .Z(n3363) );
  NANDN U3019 ( .A(n3362), .B(n3363), .Z(n1344) );
  AND U3020 ( .A(n1345), .B(n1344), .Z(n3364) );
  XOR U3021 ( .A(a[673]), .B(b[673]), .Z(n3365) );
  NANDN U3022 ( .A(n3364), .B(n3365), .Z(n1346) );
  AND U3023 ( .A(n1347), .B(n1346), .Z(n3366) );
  XOR U3024 ( .A(a[674]), .B(b[674]), .Z(n3367) );
  NANDN U3025 ( .A(n3366), .B(n3367), .Z(n1348) );
  AND U3026 ( .A(n1349), .B(n1348), .Z(n3368) );
  XOR U3027 ( .A(a[675]), .B(b[675]), .Z(n3369) );
  NANDN U3028 ( .A(n3368), .B(n3369), .Z(n1350) );
  AND U3029 ( .A(n1351), .B(n1350), .Z(n3370) );
  XOR U3030 ( .A(a[676]), .B(b[676]), .Z(n3371) );
  NANDN U3031 ( .A(n3370), .B(n3371), .Z(n1352) );
  AND U3032 ( .A(n1353), .B(n1352), .Z(n3372) );
  XOR U3033 ( .A(a[677]), .B(b[677]), .Z(n3373) );
  NANDN U3034 ( .A(n3372), .B(n3373), .Z(n1354) );
  AND U3035 ( .A(n1355), .B(n1354), .Z(n3374) );
  XOR U3036 ( .A(a[678]), .B(b[678]), .Z(n3375) );
  NANDN U3037 ( .A(n3374), .B(n3375), .Z(n1356) );
  AND U3038 ( .A(n1357), .B(n1356), .Z(n3376) );
  XOR U3039 ( .A(a[679]), .B(b[679]), .Z(n3377) );
  NANDN U3040 ( .A(n3376), .B(n3377), .Z(n1358) );
  AND U3041 ( .A(n1359), .B(n1358), .Z(n3380) );
  XOR U3042 ( .A(a[680]), .B(b[680]), .Z(n3381) );
  NANDN U3043 ( .A(n3380), .B(n3381), .Z(n1360) );
  AND U3044 ( .A(n1361), .B(n1360), .Z(n3382) );
  XOR U3045 ( .A(a[681]), .B(b[681]), .Z(n3383) );
  NANDN U3046 ( .A(n3382), .B(n3383), .Z(n1362) );
  AND U3047 ( .A(n1363), .B(n1362), .Z(n3384) );
  XOR U3048 ( .A(a[682]), .B(b[682]), .Z(n3385) );
  NANDN U3049 ( .A(n3384), .B(n3385), .Z(n1364) );
  AND U3050 ( .A(n1365), .B(n1364), .Z(n3386) );
  XOR U3051 ( .A(a[683]), .B(b[683]), .Z(n3387) );
  NANDN U3052 ( .A(n3386), .B(n3387), .Z(n1366) );
  AND U3053 ( .A(n1367), .B(n1366), .Z(n3388) );
  XOR U3054 ( .A(a[684]), .B(b[684]), .Z(n3389) );
  NANDN U3055 ( .A(n3388), .B(n3389), .Z(n1368) );
  AND U3056 ( .A(n1369), .B(n1368), .Z(n3390) );
  XOR U3057 ( .A(a[685]), .B(b[685]), .Z(n3391) );
  NANDN U3058 ( .A(n3390), .B(n3391), .Z(n1370) );
  AND U3059 ( .A(n1371), .B(n1370), .Z(n3392) );
  XOR U3060 ( .A(a[686]), .B(b[686]), .Z(n3393) );
  NANDN U3061 ( .A(n3392), .B(n3393), .Z(n1372) );
  AND U3062 ( .A(n1373), .B(n1372), .Z(n3394) );
  XOR U3063 ( .A(a[687]), .B(b[687]), .Z(n3395) );
  NANDN U3064 ( .A(n3394), .B(n3395), .Z(n1374) );
  AND U3065 ( .A(n1375), .B(n1374), .Z(n3396) );
  XOR U3066 ( .A(a[688]), .B(b[688]), .Z(n3397) );
  NANDN U3067 ( .A(n3396), .B(n3397), .Z(n1376) );
  AND U3068 ( .A(n1377), .B(n1376), .Z(n3398) );
  XOR U3069 ( .A(a[689]), .B(b[689]), .Z(n3399) );
  NANDN U3070 ( .A(n3398), .B(n3399), .Z(n1378) );
  AND U3071 ( .A(n1379), .B(n1378), .Z(n3402) );
  XOR U3072 ( .A(a[690]), .B(b[690]), .Z(n3403) );
  NANDN U3073 ( .A(n3402), .B(n3403), .Z(n1380) );
  AND U3074 ( .A(n1381), .B(n1380), .Z(n3404) );
  XOR U3075 ( .A(a[691]), .B(b[691]), .Z(n3405) );
  NANDN U3076 ( .A(n3404), .B(n3405), .Z(n1382) );
  AND U3077 ( .A(n1383), .B(n1382), .Z(n3406) );
  XOR U3078 ( .A(a[692]), .B(b[692]), .Z(n3407) );
  NANDN U3079 ( .A(n3406), .B(n3407), .Z(n1384) );
  AND U3080 ( .A(n1385), .B(n1384), .Z(n3408) );
  XOR U3081 ( .A(a[693]), .B(b[693]), .Z(n3409) );
  NANDN U3082 ( .A(n3408), .B(n3409), .Z(n1386) );
  AND U3083 ( .A(n1387), .B(n1386), .Z(n3410) );
  XOR U3084 ( .A(a[694]), .B(b[694]), .Z(n3411) );
  NANDN U3085 ( .A(n3410), .B(n3411), .Z(n1388) );
  AND U3086 ( .A(n1389), .B(n1388), .Z(n3412) );
  XOR U3087 ( .A(a[695]), .B(b[695]), .Z(n3413) );
  NANDN U3088 ( .A(n3412), .B(n3413), .Z(n1390) );
  AND U3089 ( .A(n1391), .B(n1390), .Z(n3414) );
  XOR U3090 ( .A(a[696]), .B(b[696]), .Z(n3415) );
  NANDN U3091 ( .A(n3414), .B(n3415), .Z(n1392) );
  AND U3092 ( .A(n1393), .B(n1392), .Z(n3416) );
  XOR U3093 ( .A(a[697]), .B(b[697]), .Z(n3417) );
  NANDN U3094 ( .A(n3416), .B(n3417), .Z(n1394) );
  AND U3095 ( .A(n1395), .B(n1394), .Z(n3418) );
  XOR U3096 ( .A(a[698]), .B(b[698]), .Z(n3419) );
  NANDN U3097 ( .A(n3418), .B(n3419), .Z(n1396) );
  AND U3098 ( .A(n1397), .B(n1396), .Z(n3420) );
  XOR U3099 ( .A(a[699]), .B(b[699]), .Z(n3421) );
  NANDN U3100 ( .A(n3420), .B(n3421), .Z(n1398) );
  AND U3101 ( .A(n1399), .B(n1398), .Z(n3426) );
  XOR U3102 ( .A(a[700]), .B(b[700]), .Z(n3427) );
  NANDN U3103 ( .A(n3426), .B(n3427), .Z(n1400) );
  AND U3104 ( .A(n1401), .B(n1400), .Z(n3428) );
  XOR U3105 ( .A(a[701]), .B(b[701]), .Z(n3429) );
  NANDN U3106 ( .A(n3428), .B(n3429), .Z(n1402) );
  AND U3107 ( .A(n1403), .B(n1402), .Z(n3430) );
  XOR U3108 ( .A(a[702]), .B(b[702]), .Z(n3431) );
  NANDN U3109 ( .A(n3430), .B(n3431), .Z(n1404) );
  AND U3110 ( .A(n1405), .B(n1404), .Z(n3432) );
  XOR U3111 ( .A(a[703]), .B(b[703]), .Z(n3433) );
  NANDN U3112 ( .A(n3432), .B(n3433), .Z(n1406) );
  AND U3113 ( .A(n1407), .B(n1406), .Z(n3434) );
  XOR U3114 ( .A(a[704]), .B(b[704]), .Z(n3435) );
  NANDN U3115 ( .A(n3434), .B(n3435), .Z(n1408) );
  AND U3116 ( .A(n1409), .B(n1408), .Z(n3436) );
  XOR U3117 ( .A(a[705]), .B(b[705]), .Z(n3437) );
  NANDN U3118 ( .A(n3436), .B(n3437), .Z(n1410) );
  AND U3119 ( .A(n1411), .B(n1410), .Z(n3438) );
  XOR U3120 ( .A(a[706]), .B(b[706]), .Z(n3439) );
  NANDN U3121 ( .A(n3438), .B(n3439), .Z(n1412) );
  AND U3122 ( .A(n1413), .B(n1412), .Z(n3440) );
  XOR U3123 ( .A(a[707]), .B(b[707]), .Z(n3441) );
  NANDN U3124 ( .A(n3440), .B(n3441), .Z(n1414) );
  AND U3125 ( .A(n1415), .B(n1414), .Z(n3442) );
  XOR U3126 ( .A(a[708]), .B(b[708]), .Z(n3443) );
  NANDN U3127 ( .A(n3442), .B(n3443), .Z(n1416) );
  AND U3128 ( .A(n1417), .B(n1416), .Z(n3444) );
  XOR U3129 ( .A(a[709]), .B(b[709]), .Z(n3445) );
  NANDN U3130 ( .A(n3444), .B(n3445), .Z(n1418) );
  AND U3131 ( .A(n1419), .B(n1418), .Z(n3448) );
  XOR U3132 ( .A(a[710]), .B(b[710]), .Z(n3449) );
  NANDN U3133 ( .A(n3448), .B(n3449), .Z(n1420) );
  AND U3134 ( .A(n1421), .B(n1420), .Z(n3450) );
  XOR U3135 ( .A(a[711]), .B(b[711]), .Z(n3451) );
  NANDN U3136 ( .A(n3450), .B(n3451), .Z(n1422) );
  AND U3137 ( .A(n1423), .B(n1422), .Z(n3452) );
  XOR U3138 ( .A(a[712]), .B(b[712]), .Z(n3453) );
  NANDN U3139 ( .A(n3452), .B(n3453), .Z(n1424) );
  AND U3140 ( .A(n1425), .B(n1424), .Z(n3454) );
  XOR U3141 ( .A(a[713]), .B(b[713]), .Z(n3455) );
  NANDN U3142 ( .A(n3454), .B(n3455), .Z(n1426) );
  AND U3143 ( .A(n1427), .B(n1426), .Z(n3456) );
  XOR U3144 ( .A(a[714]), .B(b[714]), .Z(n3457) );
  NANDN U3145 ( .A(n3456), .B(n3457), .Z(n1428) );
  AND U3146 ( .A(n1429), .B(n1428), .Z(n3458) );
  XOR U3147 ( .A(a[715]), .B(b[715]), .Z(n3459) );
  NANDN U3148 ( .A(n3458), .B(n3459), .Z(n1430) );
  AND U3149 ( .A(n1431), .B(n1430), .Z(n3460) );
  XOR U3150 ( .A(a[716]), .B(b[716]), .Z(n3461) );
  NANDN U3151 ( .A(n3460), .B(n3461), .Z(n1432) );
  AND U3152 ( .A(n1433), .B(n1432), .Z(n3462) );
  XOR U3153 ( .A(a[717]), .B(b[717]), .Z(n3463) );
  NANDN U3154 ( .A(n3462), .B(n3463), .Z(n1434) );
  AND U3155 ( .A(n1435), .B(n1434), .Z(n3464) );
  XOR U3156 ( .A(a[718]), .B(b[718]), .Z(n3465) );
  NANDN U3157 ( .A(n3464), .B(n3465), .Z(n1436) );
  AND U3158 ( .A(n1437), .B(n1436), .Z(n3466) );
  XOR U3159 ( .A(a[719]), .B(b[719]), .Z(n3467) );
  NANDN U3160 ( .A(n3466), .B(n3467), .Z(n1438) );
  AND U3161 ( .A(n1439), .B(n1438), .Z(n3470) );
  XOR U3162 ( .A(a[720]), .B(b[720]), .Z(n3471) );
  NANDN U3163 ( .A(n3470), .B(n3471), .Z(n1440) );
  AND U3164 ( .A(n1441), .B(n1440), .Z(n3472) );
  XOR U3165 ( .A(a[721]), .B(b[721]), .Z(n3473) );
  NANDN U3166 ( .A(n3472), .B(n3473), .Z(n1442) );
  AND U3167 ( .A(n1443), .B(n1442), .Z(n3474) );
  XOR U3168 ( .A(a[722]), .B(b[722]), .Z(n3475) );
  NANDN U3169 ( .A(n3474), .B(n3475), .Z(n1444) );
  AND U3170 ( .A(n1445), .B(n1444), .Z(n3476) );
  XOR U3171 ( .A(a[723]), .B(b[723]), .Z(n3477) );
  NANDN U3172 ( .A(n3476), .B(n3477), .Z(n1446) );
  AND U3173 ( .A(n1447), .B(n1446), .Z(n3478) );
  XOR U3174 ( .A(a[724]), .B(b[724]), .Z(n3479) );
  NANDN U3175 ( .A(n3478), .B(n3479), .Z(n1448) );
  AND U3176 ( .A(n1449), .B(n1448), .Z(n3480) );
  XOR U3177 ( .A(a[725]), .B(b[725]), .Z(n3481) );
  NANDN U3178 ( .A(n3480), .B(n3481), .Z(n1450) );
  AND U3179 ( .A(n1451), .B(n1450), .Z(n3482) );
  XOR U3180 ( .A(a[726]), .B(b[726]), .Z(n3483) );
  NANDN U3181 ( .A(n3482), .B(n3483), .Z(n1452) );
  AND U3182 ( .A(n1453), .B(n1452), .Z(n3484) );
  XOR U3183 ( .A(a[727]), .B(b[727]), .Z(n3485) );
  NANDN U3184 ( .A(n3484), .B(n3485), .Z(n1454) );
  AND U3185 ( .A(n1455), .B(n1454), .Z(n3486) );
  XOR U3186 ( .A(a[728]), .B(b[728]), .Z(n3487) );
  NANDN U3187 ( .A(n3486), .B(n3487), .Z(n1456) );
  AND U3188 ( .A(n1457), .B(n1456), .Z(n3488) );
  XOR U3189 ( .A(a[729]), .B(b[729]), .Z(n3489) );
  NANDN U3190 ( .A(n3488), .B(n3489), .Z(n1458) );
  AND U3191 ( .A(n1459), .B(n1458), .Z(n3492) );
  XOR U3192 ( .A(a[730]), .B(b[730]), .Z(n3493) );
  NANDN U3193 ( .A(n3492), .B(n3493), .Z(n1460) );
  AND U3194 ( .A(n1461), .B(n1460), .Z(n3494) );
  XOR U3195 ( .A(a[731]), .B(b[731]), .Z(n3495) );
  NANDN U3196 ( .A(n3494), .B(n3495), .Z(n1462) );
  AND U3197 ( .A(n1463), .B(n1462), .Z(n3496) );
  XOR U3198 ( .A(a[732]), .B(b[732]), .Z(n3497) );
  NANDN U3199 ( .A(n3496), .B(n3497), .Z(n1464) );
  AND U3200 ( .A(n1465), .B(n1464), .Z(n3498) );
  XOR U3201 ( .A(a[733]), .B(b[733]), .Z(n3499) );
  NANDN U3202 ( .A(n3498), .B(n3499), .Z(n1466) );
  AND U3203 ( .A(n1467), .B(n1466), .Z(n3500) );
  XOR U3204 ( .A(a[734]), .B(b[734]), .Z(n3501) );
  NANDN U3205 ( .A(n3500), .B(n3501), .Z(n1468) );
  AND U3206 ( .A(n1469), .B(n1468), .Z(n3502) );
  XOR U3207 ( .A(a[735]), .B(b[735]), .Z(n3503) );
  NANDN U3208 ( .A(n3502), .B(n3503), .Z(n1470) );
  AND U3209 ( .A(n1471), .B(n1470), .Z(n3504) );
  XOR U3210 ( .A(a[736]), .B(b[736]), .Z(n3505) );
  NANDN U3211 ( .A(n3504), .B(n3505), .Z(n1472) );
  AND U3212 ( .A(n1473), .B(n1472), .Z(n3506) );
  XOR U3213 ( .A(a[737]), .B(b[737]), .Z(n3507) );
  NANDN U3214 ( .A(n3506), .B(n3507), .Z(n1474) );
  AND U3215 ( .A(n1475), .B(n1474), .Z(n3508) );
  XOR U3216 ( .A(a[738]), .B(b[738]), .Z(n3509) );
  NANDN U3217 ( .A(n3508), .B(n3509), .Z(n1476) );
  AND U3218 ( .A(n1477), .B(n1476), .Z(n3510) );
  XOR U3219 ( .A(a[739]), .B(b[739]), .Z(n3511) );
  NANDN U3220 ( .A(n3510), .B(n3511), .Z(n1478) );
  AND U3221 ( .A(n1479), .B(n1478), .Z(n3514) );
  XOR U3222 ( .A(a[740]), .B(b[740]), .Z(n3515) );
  NANDN U3223 ( .A(n3514), .B(n3515), .Z(n1480) );
  AND U3224 ( .A(n1481), .B(n1480), .Z(n3516) );
  XOR U3225 ( .A(a[741]), .B(b[741]), .Z(n3517) );
  NANDN U3226 ( .A(n3516), .B(n3517), .Z(n1482) );
  AND U3227 ( .A(n1483), .B(n1482), .Z(n3518) );
  XOR U3228 ( .A(a[742]), .B(b[742]), .Z(n3519) );
  NANDN U3229 ( .A(n3518), .B(n3519), .Z(n1484) );
  AND U3230 ( .A(n1485), .B(n1484), .Z(n3520) );
  XOR U3231 ( .A(a[743]), .B(b[743]), .Z(n3521) );
  NANDN U3232 ( .A(n3520), .B(n3521), .Z(n1486) );
  AND U3233 ( .A(n1487), .B(n1486), .Z(n3522) );
  XOR U3234 ( .A(a[744]), .B(b[744]), .Z(n3523) );
  NANDN U3235 ( .A(n3522), .B(n3523), .Z(n1488) );
  AND U3236 ( .A(n1489), .B(n1488), .Z(n3524) );
  XOR U3237 ( .A(a[745]), .B(b[745]), .Z(n3525) );
  NANDN U3238 ( .A(n3524), .B(n3525), .Z(n1490) );
  AND U3239 ( .A(n1491), .B(n1490), .Z(n3526) );
  XOR U3240 ( .A(a[746]), .B(b[746]), .Z(n3527) );
  NANDN U3241 ( .A(n3526), .B(n3527), .Z(n1492) );
  AND U3242 ( .A(n1493), .B(n1492), .Z(n3528) );
  XOR U3243 ( .A(a[747]), .B(b[747]), .Z(n3529) );
  NANDN U3244 ( .A(n3528), .B(n3529), .Z(n1494) );
  AND U3245 ( .A(n1495), .B(n1494), .Z(n3530) );
  XOR U3246 ( .A(a[748]), .B(b[748]), .Z(n3531) );
  NANDN U3247 ( .A(n3530), .B(n3531), .Z(n1496) );
  AND U3248 ( .A(n1497), .B(n1496), .Z(n3532) );
  XOR U3249 ( .A(a[749]), .B(b[749]), .Z(n3533) );
  NANDN U3250 ( .A(n3532), .B(n3533), .Z(n1498) );
  AND U3251 ( .A(n1499), .B(n1498), .Z(n3536) );
  XOR U3252 ( .A(a[750]), .B(b[750]), .Z(n3537) );
  NANDN U3253 ( .A(n3536), .B(n3537), .Z(n1500) );
  AND U3254 ( .A(n1501), .B(n1500), .Z(n3538) );
  XOR U3255 ( .A(a[751]), .B(b[751]), .Z(n3539) );
  NANDN U3256 ( .A(n3538), .B(n3539), .Z(n1502) );
  AND U3257 ( .A(n1503), .B(n1502), .Z(n3540) );
  XOR U3258 ( .A(a[752]), .B(b[752]), .Z(n3541) );
  NANDN U3259 ( .A(n3540), .B(n3541), .Z(n1504) );
  AND U3260 ( .A(n1505), .B(n1504), .Z(n3542) );
  XOR U3261 ( .A(a[753]), .B(b[753]), .Z(n3543) );
  NANDN U3262 ( .A(n3542), .B(n3543), .Z(n1506) );
  AND U3263 ( .A(n1507), .B(n1506), .Z(n3544) );
  XOR U3264 ( .A(a[754]), .B(b[754]), .Z(n3545) );
  NANDN U3265 ( .A(n3544), .B(n3545), .Z(n1508) );
  AND U3266 ( .A(n1509), .B(n1508), .Z(n3546) );
  XOR U3267 ( .A(a[755]), .B(b[755]), .Z(n3547) );
  NANDN U3268 ( .A(n3546), .B(n3547), .Z(n1510) );
  AND U3269 ( .A(n1511), .B(n1510), .Z(n3548) );
  XOR U3270 ( .A(a[756]), .B(b[756]), .Z(n3549) );
  NANDN U3271 ( .A(n3548), .B(n3549), .Z(n1512) );
  AND U3272 ( .A(n1513), .B(n1512), .Z(n3550) );
  XOR U3273 ( .A(a[757]), .B(b[757]), .Z(n3551) );
  NANDN U3274 ( .A(n3550), .B(n3551), .Z(n1514) );
  AND U3275 ( .A(n1515), .B(n1514), .Z(n3552) );
  XOR U3276 ( .A(a[758]), .B(b[758]), .Z(n3553) );
  NANDN U3277 ( .A(n3552), .B(n3553), .Z(n1516) );
  AND U3278 ( .A(n1517), .B(n1516), .Z(n3554) );
  XOR U3279 ( .A(a[759]), .B(b[759]), .Z(n3555) );
  NANDN U3280 ( .A(n3554), .B(n3555), .Z(n1518) );
  AND U3281 ( .A(n1519), .B(n1518), .Z(n3558) );
  XOR U3282 ( .A(a[760]), .B(b[760]), .Z(n3559) );
  NANDN U3283 ( .A(n3558), .B(n3559), .Z(n1520) );
  AND U3284 ( .A(n1521), .B(n1520), .Z(n3560) );
  XOR U3285 ( .A(a[761]), .B(b[761]), .Z(n3561) );
  NANDN U3286 ( .A(n3560), .B(n3561), .Z(n1522) );
  AND U3287 ( .A(n1523), .B(n1522), .Z(n3562) );
  XOR U3288 ( .A(a[762]), .B(b[762]), .Z(n3563) );
  NANDN U3289 ( .A(n3562), .B(n3563), .Z(n1524) );
  AND U3290 ( .A(n1525), .B(n1524), .Z(n3564) );
  XOR U3291 ( .A(a[763]), .B(b[763]), .Z(n3565) );
  NANDN U3292 ( .A(n3564), .B(n3565), .Z(n1526) );
  AND U3293 ( .A(n1527), .B(n1526), .Z(n3566) );
  XOR U3294 ( .A(a[764]), .B(b[764]), .Z(n3567) );
  NANDN U3295 ( .A(n3566), .B(n3567), .Z(n1528) );
  AND U3296 ( .A(n1529), .B(n1528), .Z(n3568) );
  XOR U3297 ( .A(a[765]), .B(b[765]), .Z(n3569) );
  NANDN U3298 ( .A(n3568), .B(n3569), .Z(n1530) );
  AND U3299 ( .A(n1531), .B(n1530), .Z(n3570) );
  XOR U3300 ( .A(a[766]), .B(b[766]), .Z(n3571) );
  NANDN U3301 ( .A(n3570), .B(n3571), .Z(n1532) );
  AND U3302 ( .A(n1533), .B(n1532), .Z(n3572) );
  XOR U3303 ( .A(a[767]), .B(b[767]), .Z(n3573) );
  NANDN U3304 ( .A(n3572), .B(n3573), .Z(n1534) );
  AND U3305 ( .A(n1535), .B(n1534), .Z(n3574) );
  XOR U3306 ( .A(a[768]), .B(b[768]), .Z(n3575) );
  NANDN U3307 ( .A(n3574), .B(n3575), .Z(n1536) );
  AND U3308 ( .A(n1537), .B(n1536), .Z(n3576) );
  XOR U3309 ( .A(a[769]), .B(b[769]), .Z(n3577) );
  NANDN U3310 ( .A(n3576), .B(n3577), .Z(n1538) );
  AND U3311 ( .A(n1539), .B(n1538), .Z(n3580) );
  XOR U3312 ( .A(a[770]), .B(b[770]), .Z(n3581) );
  NANDN U3313 ( .A(n3580), .B(n3581), .Z(n1540) );
  AND U3314 ( .A(n1541), .B(n1540), .Z(n3582) );
  XOR U3315 ( .A(a[771]), .B(b[771]), .Z(n3583) );
  NANDN U3316 ( .A(n3582), .B(n3583), .Z(n1542) );
  AND U3317 ( .A(n1543), .B(n1542), .Z(n3584) );
  XOR U3318 ( .A(a[772]), .B(b[772]), .Z(n3585) );
  NANDN U3319 ( .A(n3584), .B(n3585), .Z(n1544) );
  AND U3320 ( .A(n1545), .B(n1544), .Z(n3586) );
  XOR U3321 ( .A(a[773]), .B(b[773]), .Z(n3587) );
  NANDN U3322 ( .A(n3586), .B(n3587), .Z(n1546) );
  AND U3323 ( .A(n1547), .B(n1546), .Z(n3588) );
  XOR U3324 ( .A(a[774]), .B(b[774]), .Z(n3589) );
  NANDN U3325 ( .A(n3588), .B(n3589), .Z(n1548) );
  AND U3326 ( .A(n1549), .B(n1548), .Z(n3590) );
  XOR U3327 ( .A(a[775]), .B(b[775]), .Z(n3591) );
  NANDN U3328 ( .A(n3590), .B(n3591), .Z(n1550) );
  AND U3329 ( .A(n1551), .B(n1550), .Z(n3592) );
  XOR U3330 ( .A(a[776]), .B(b[776]), .Z(n3593) );
  NANDN U3331 ( .A(n3592), .B(n3593), .Z(n1552) );
  AND U3332 ( .A(n1553), .B(n1552), .Z(n3594) );
  XOR U3333 ( .A(a[777]), .B(b[777]), .Z(n3595) );
  NANDN U3334 ( .A(n3594), .B(n3595), .Z(n1554) );
  AND U3335 ( .A(n1555), .B(n1554), .Z(n3596) );
  XOR U3336 ( .A(a[778]), .B(b[778]), .Z(n3597) );
  NANDN U3337 ( .A(n3596), .B(n3597), .Z(n1556) );
  AND U3338 ( .A(n1557), .B(n1556), .Z(n3598) );
  XOR U3339 ( .A(a[779]), .B(b[779]), .Z(n3599) );
  NANDN U3340 ( .A(n3598), .B(n3599), .Z(n1558) );
  AND U3341 ( .A(n1559), .B(n1558), .Z(n3602) );
  XOR U3342 ( .A(a[780]), .B(b[780]), .Z(n3603) );
  NANDN U3343 ( .A(n3602), .B(n3603), .Z(n1560) );
  AND U3344 ( .A(n1561), .B(n1560), .Z(n3604) );
  XOR U3345 ( .A(a[781]), .B(b[781]), .Z(n3605) );
  NANDN U3346 ( .A(n3604), .B(n3605), .Z(n1562) );
  AND U3347 ( .A(n1563), .B(n1562), .Z(n3606) );
  XOR U3348 ( .A(a[782]), .B(b[782]), .Z(n3607) );
  NANDN U3349 ( .A(n3606), .B(n3607), .Z(n1564) );
  AND U3350 ( .A(n1565), .B(n1564), .Z(n3608) );
  XOR U3351 ( .A(a[783]), .B(b[783]), .Z(n3609) );
  NANDN U3352 ( .A(n3608), .B(n3609), .Z(n1566) );
  AND U3353 ( .A(n1567), .B(n1566), .Z(n3610) );
  XOR U3354 ( .A(a[784]), .B(b[784]), .Z(n3611) );
  NANDN U3355 ( .A(n3610), .B(n3611), .Z(n1568) );
  AND U3356 ( .A(n1569), .B(n1568), .Z(n3612) );
  XOR U3357 ( .A(a[785]), .B(b[785]), .Z(n3613) );
  NANDN U3358 ( .A(n3612), .B(n3613), .Z(n1570) );
  AND U3359 ( .A(n1571), .B(n1570), .Z(n3614) );
  XOR U3360 ( .A(a[786]), .B(b[786]), .Z(n3615) );
  NANDN U3361 ( .A(n3614), .B(n3615), .Z(n1572) );
  AND U3362 ( .A(n1573), .B(n1572), .Z(n3616) );
  XOR U3363 ( .A(a[787]), .B(b[787]), .Z(n3617) );
  NANDN U3364 ( .A(n3616), .B(n3617), .Z(n1574) );
  AND U3365 ( .A(n1575), .B(n1574), .Z(n3618) );
  XOR U3366 ( .A(a[788]), .B(b[788]), .Z(n3619) );
  NANDN U3367 ( .A(n3618), .B(n3619), .Z(n1576) );
  AND U3368 ( .A(n1577), .B(n1576), .Z(n3620) );
  XOR U3369 ( .A(a[789]), .B(b[789]), .Z(n3621) );
  NANDN U3370 ( .A(n3620), .B(n3621), .Z(n1578) );
  AND U3371 ( .A(n1579), .B(n1578), .Z(n3624) );
  XOR U3372 ( .A(a[790]), .B(b[790]), .Z(n3625) );
  NANDN U3373 ( .A(n3624), .B(n3625), .Z(n1580) );
  AND U3374 ( .A(n1581), .B(n1580), .Z(n3626) );
  XOR U3375 ( .A(a[791]), .B(b[791]), .Z(n3627) );
  NANDN U3376 ( .A(n3626), .B(n3627), .Z(n1582) );
  AND U3377 ( .A(n1583), .B(n1582), .Z(n3628) );
  XOR U3378 ( .A(a[792]), .B(b[792]), .Z(n3629) );
  NANDN U3379 ( .A(n3628), .B(n3629), .Z(n1584) );
  AND U3380 ( .A(n1585), .B(n1584), .Z(n3630) );
  XOR U3381 ( .A(a[793]), .B(b[793]), .Z(n3631) );
  NANDN U3382 ( .A(n3630), .B(n3631), .Z(n1586) );
  AND U3383 ( .A(n1587), .B(n1586), .Z(n3632) );
  XOR U3384 ( .A(a[794]), .B(b[794]), .Z(n3633) );
  NANDN U3385 ( .A(n3632), .B(n3633), .Z(n1588) );
  AND U3386 ( .A(n1589), .B(n1588), .Z(n3634) );
  XOR U3387 ( .A(a[795]), .B(b[795]), .Z(n3635) );
  NANDN U3388 ( .A(n3634), .B(n3635), .Z(n1590) );
  AND U3389 ( .A(n1591), .B(n1590), .Z(n3636) );
  XOR U3390 ( .A(a[796]), .B(b[796]), .Z(n3637) );
  NANDN U3391 ( .A(n3636), .B(n3637), .Z(n1592) );
  AND U3392 ( .A(n1593), .B(n1592), .Z(n3638) );
  XOR U3393 ( .A(a[797]), .B(b[797]), .Z(n3639) );
  NANDN U3394 ( .A(n3638), .B(n3639), .Z(n1594) );
  AND U3395 ( .A(n1595), .B(n1594), .Z(n3640) );
  XOR U3396 ( .A(a[798]), .B(b[798]), .Z(n3641) );
  NANDN U3397 ( .A(n3640), .B(n3641), .Z(n1596) );
  AND U3398 ( .A(n1597), .B(n1596), .Z(n3642) );
  XOR U3399 ( .A(a[799]), .B(b[799]), .Z(n3643) );
  NANDN U3400 ( .A(n3642), .B(n3643), .Z(n1598) );
  AND U3401 ( .A(n1599), .B(n1598), .Z(n3648) );
  XOR U3402 ( .A(a[800]), .B(b[800]), .Z(n3649) );
  NANDN U3403 ( .A(n3648), .B(n3649), .Z(n1600) );
  AND U3404 ( .A(n1601), .B(n1600), .Z(n3650) );
  XOR U3405 ( .A(a[801]), .B(b[801]), .Z(n3651) );
  NANDN U3406 ( .A(n3650), .B(n3651), .Z(n1602) );
  AND U3407 ( .A(n1603), .B(n1602), .Z(n3652) );
  XOR U3408 ( .A(a[802]), .B(b[802]), .Z(n3653) );
  NANDN U3409 ( .A(n3652), .B(n3653), .Z(n1604) );
  AND U3410 ( .A(n1605), .B(n1604), .Z(n3654) );
  XOR U3411 ( .A(a[803]), .B(b[803]), .Z(n3655) );
  NANDN U3412 ( .A(n3654), .B(n3655), .Z(n1606) );
  AND U3413 ( .A(n1607), .B(n1606), .Z(n3656) );
  XOR U3414 ( .A(a[804]), .B(b[804]), .Z(n3657) );
  NANDN U3415 ( .A(n3656), .B(n3657), .Z(n1608) );
  AND U3416 ( .A(n1609), .B(n1608), .Z(n3658) );
  XOR U3417 ( .A(a[805]), .B(b[805]), .Z(n3659) );
  NANDN U3418 ( .A(n3658), .B(n3659), .Z(n1610) );
  AND U3419 ( .A(n1611), .B(n1610), .Z(n3660) );
  XOR U3420 ( .A(a[806]), .B(b[806]), .Z(n3661) );
  NANDN U3421 ( .A(n3660), .B(n3661), .Z(n1612) );
  AND U3422 ( .A(n1613), .B(n1612), .Z(n3662) );
  XOR U3423 ( .A(a[807]), .B(b[807]), .Z(n3663) );
  NANDN U3424 ( .A(n3662), .B(n3663), .Z(n1614) );
  AND U3425 ( .A(n1615), .B(n1614), .Z(n3664) );
  XOR U3426 ( .A(a[808]), .B(b[808]), .Z(n3665) );
  NANDN U3427 ( .A(n3664), .B(n3665), .Z(n1616) );
  AND U3428 ( .A(n1617), .B(n1616), .Z(n3666) );
  XOR U3429 ( .A(a[809]), .B(b[809]), .Z(n3667) );
  NANDN U3430 ( .A(n3666), .B(n3667), .Z(n1618) );
  AND U3431 ( .A(n1619), .B(n1618), .Z(n3670) );
  XOR U3432 ( .A(a[810]), .B(b[810]), .Z(n3671) );
  NANDN U3433 ( .A(n3670), .B(n3671), .Z(n1620) );
  AND U3434 ( .A(n1621), .B(n1620), .Z(n3672) );
  XOR U3435 ( .A(a[811]), .B(b[811]), .Z(n3673) );
  NANDN U3436 ( .A(n3672), .B(n3673), .Z(n1622) );
  AND U3437 ( .A(n1623), .B(n1622), .Z(n3674) );
  XOR U3438 ( .A(a[812]), .B(b[812]), .Z(n3675) );
  NANDN U3439 ( .A(n3674), .B(n3675), .Z(n1624) );
  AND U3440 ( .A(n1625), .B(n1624), .Z(n3676) );
  XOR U3441 ( .A(a[813]), .B(b[813]), .Z(n3677) );
  NANDN U3442 ( .A(n3676), .B(n3677), .Z(n1626) );
  AND U3443 ( .A(n1627), .B(n1626), .Z(n3678) );
  XOR U3444 ( .A(a[814]), .B(b[814]), .Z(n3679) );
  NANDN U3445 ( .A(n3678), .B(n3679), .Z(n1628) );
  AND U3446 ( .A(n1629), .B(n1628), .Z(n3680) );
  XOR U3447 ( .A(a[815]), .B(b[815]), .Z(n3681) );
  NANDN U3448 ( .A(n3680), .B(n3681), .Z(n1630) );
  AND U3449 ( .A(n1631), .B(n1630), .Z(n3682) );
  XOR U3450 ( .A(a[816]), .B(b[816]), .Z(n3683) );
  NANDN U3451 ( .A(n3682), .B(n3683), .Z(n1632) );
  AND U3452 ( .A(n1633), .B(n1632), .Z(n3684) );
  XOR U3453 ( .A(a[817]), .B(b[817]), .Z(n3685) );
  NANDN U3454 ( .A(n3684), .B(n3685), .Z(n1634) );
  AND U3455 ( .A(n1635), .B(n1634), .Z(n3686) );
  XOR U3456 ( .A(a[818]), .B(b[818]), .Z(n3687) );
  NANDN U3457 ( .A(n3686), .B(n3687), .Z(n1636) );
  AND U3458 ( .A(n1637), .B(n1636), .Z(n3688) );
  XOR U3459 ( .A(a[819]), .B(b[819]), .Z(n3689) );
  NANDN U3460 ( .A(n3688), .B(n3689), .Z(n1638) );
  AND U3461 ( .A(n1639), .B(n1638), .Z(n3692) );
  XOR U3462 ( .A(a[820]), .B(b[820]), .Z(n3693) );
  NANDN U3463 ( .A(n3692), .B(n3693), .Z(n1640) );
  AND U3464 ( .A(n1641), .B(n1640), .Z(n3694) );
  XOR U3465 ( .A(a[821]), .B(b[821]), .Z(n3695) );
  NANDN U3466 ( .A(n3694), .B(n3695), .Z(n1642) );
  AND U3467 ( .A(n1643), .B(n1642), .Z(n3696) );
  XOR U3468 ( .A(a[822]), .B(b[822]), .Z(n3697) );
  NANDN U3469 ( .A(n3696), .B(n3697), .Z(n1644) );
  AND U3470 ( .A(n1645), .B(n1644), .Z(n3698) );
  XOR U3471 ( .A(a[823]), .B(b[823]), .Z(n3699) );
  NANDN U3472 ( .A(n3698), .B(n3699), .Z(n1646) );
  AND U3473 ( .A(n1647), .B(n1646), .Z(n3700) );
  XOR U3474 ( .A(a[824]), .B(b[824]), .Z(n3701) );
  NANDN U3475 ( .A(n3700), .B(n3701), .Z(n1648) );
  AND U3476 ( .A(n1649), .B(n1648), .Z(n3702) );
  XOR U3477 ( .A(a[825]), .B(b[825]), .Z(n3703) );
  NANDN U3478 ( .A(n3702), .B(n3703), .Z(n1650) );
  AND U3479 ( .A(n1651), .B(n1650), .Z(n3704) );
  XOR U3480 ( .A(a[826]), .B(b[826]), .Z(n3705) );
  NANDN U3481 ( .A(n3704), .B(n3705), .Z(n1652) );
  AND U3482 ( .A(n1653), .B(n1652), .Z(n3706) );
  XOR U3483 ( .A(a[827]), .B(b[827]), .Z(n3707) );
  NANDN U3484 ( .A(n3706), .B(n3707), .Z(n1654) );
  AND U3485 ( .A(n1655), .B(n1654), .Z(n3708) );
  XOR U3486 ( .A(a[828]), .B(b[828]), .Z(n3709) );
  NANDN U3487 ( .A(n3708), .B(n3709), .Z(n1656) );
  AND U3488 ( .A(n1657), .B(n1656), .Z(n3710) );
  XOR U3489 ( .A(a[829]), .B(b[829]), .Z(n3711) );
  NANDN U3490 ( .A(n3710), .B(n3711), .Z(n1658) );
  AND U3491 ( .A(n1659), .B(n1658), .Z(n3714) );
  XOR U3492 ( .A(a[830]), .B(b[830]), .Z(n3715) );
  NANDN U3493 ( .A(n3714), .B(n3715), .Z(n1660) );
  AND U3494 ( .A(n1661), .B(n1660), .Z(n3716) );
  XOR U3495 ( .A(a[831]), .B(b[831]), .Z(n3717) );
  NANDN U3496 ( .A(n3716), .B(n3717), .Z(n1662) );
  AND U3497 ( .A(n1663), .B(n1662), .Z(n3718) );
  XOR U3498 ( .A(a[832]), .B(b[832]), .Z(n3719) );
  NANDN U3499 ( .A(n3718), .B(n3719), .Z(n1664) );
  AND U3500 ( .A(n1665), .B(n1664), .Z(n3720) );
  XOR U3501 ( .A(a[833]), .B(b[833]), .Z(n3721) );
  NANDN U3502 ( .A(n3720), .B(n3721), .Z(n1666) );
  AND U3503 ( .A(n1667), .B(n1666), .Z(n3722) );
  XOR U3504 ( .A(a[834]), .B(b[834]), .Z(n3723) );
  NANDN U3505 ( .A(n3722), .B(n3723), .Z(n1668) );
  AND U3506 ( .A(n1669), .B(n1668), .Z(n3724) );
  XOR U3507 ( .A(a[835]), .B(b[835]), .Z(n3725) );
  NANDN U3508 ( .A(n3724), .B(n3725), .Z(n1670) );
  AND U3509 ( .A(n1671), .B(n1670), .Z(n3726) );
  XOR U3510 ( .A(a[836]), .B(b[836]), .Z(n3727) );
  NANDN U3511 ( .A(n3726), .B(n3727), .Z(n1672) );
  AND U3512 ( .A(n1673), .B(n1672), .Z(n3728) );
  XOR U3513 ( .A(a[837]), .B(b[837]), .Z(n3729) );
  NANDN U3514 ( .A(n3728), .B(n3729), .Z(n1674) );
  AND U3515 ( .A(n1675), .B(n1674), .Z(n3730) );
  XOR U3516 ( .A(a[838]), .B(b[838]), .Z(n3731) );
  NANDN U3517 ( .A(n3730), .B(n3731), .Z(n1676) );
  AND U3518 ( .A(n1677), .B(n1676), .Z(n3732) );
  XOR U3519 ( .A(a[839]), .B(b[839]), .Z(n3733) );
  NANDN U3520 ( .A(n3732), .B(n3733), .Z(n1678) );
  AND U3521 ( .A(n1679), .B(n1678), .Z(n3736) );
  XOR U3522 ( .A(a[840]), .B(b[840]), .Z(n3737) );
  NANDN U3523 ( .A(n3736), .B(n3737), .Z(n1680) );
  AND U3524 ( .A(n1681), .B(n1680), .Z(n3738) );
  XOR U3525 ( .A(a[841]), .B(b[841]), .Z(n3739) );
  NANDN U3526 ( .A(n3738), .B(n3739), .Z(n1682) );
  AND U3527 ( .A(n1683), .B(n1682), .Z(n3740) );
  XOR U3528 ( .A(a[842]), .B(b[842]), .Z(n3741) );
  NANDN U3529 ( .A(n3740), .B(n3741), .Z(n1684) );
  AND U3530 ( .A(n1685), .B(n1684), .Z(n3742) );
  XOR U3531 ( .A(a[843]), .B(b[843]), .Z(n3743) );
  NANDN U3532 ( .A(n3742), .B(n3743), .Z(n1686) );
  AND U3533 ( .A(n1687), .B(n1686), .Z(n3744) );
  XOR U3534 ( .A(a[844]), .B(b[844]), .Z(n3745) );
  NANDN U3535 ( .A(n3744), .B(n3745), .Z(n1688) );
  AND U3536 ( .A(n1689), .B(n1688), .Z(n3746) );
  XOR U3537 ( .A(a[845]), .B(b[845]), .Z(n3747) );
  NANDN U3538 ( .A(n3746), .B(n3747), .Z(n1690) );
  AND U3539 ( .A(n1691), .B(n1690), .Z(n3748) );
  XOR U3540 ( .A(a[846]), .B(b[846]), .Z(n3749) );
  NANDN U3541 ( .A(n3748), .B(n3749), .Z(n1692) );
  AND U3542 ( .A(n1693), .B(n1692), .Z(n3750) );
  XOR U3543 ( .A(a[847]), .B(b[847]), .Z(n3751) );
  NANDN U3544 ( .A(n3750), .B(n3751), .Z(n1694) );
  AND U3545 ( .A(n1695), .B(n1694), .Z(n3752) );
  XOR U3546 ( .A(a[848]), .B(b[848]), .Z(n3753) );
  NANDN U3547 ( .A(n3752), .B(n3753), .Z(n1696) );
  AND U3548 ( .A(n1697), .B(n1696), .Z(n3754) );
  XOR U3549 ( .A(a[849]), .B(b[849]), .Z(n3755) );
  NANDN U3550 ( .A(n3754), .B(n3755), .Z(n1698) );
  AND U3551 ( .A(n1699), .B(n1698), .Z(n3758) );
  XOR U3552 ( .A(a[850]), .B(b[850]), .Z(n3759) );
  NANDN U3553 ( .A(n3758), .B(n3759), .Z(n1700) );
  AND U3554 ( .A(n1701), .B(n1700), .Z(n3760) );
  XOR U3555 ( .A(a[851]), .B(b[851]), .Z(n3761) );
  NANDN U3556 ( .A(n3760), .B(n3761), .Z(n1702) );
  AND U3557 ( .A(n1703), .B(n1702), .Z(n3762) );
  XOR U3558 ( .A(a[852]), .B(b[852]), .Z(n3763) );
  NANDN U3559 ( .A(n3762), .B(n3763), .Z(n1704) );
  AND U3560 ( .A(n1705), .B(n1704), .Z(n3764) );
  XOR U3561 ( .A(a[853]), .B(b[853]), .Z(n3765) );
  NANDN U3562 ( .A(n3764), .B(n3765), .Z(n1706) );
  AND U3563 ( .A(n1707), .B(n1706), .Z(n3766) );
  XOR U3564 ( .A(a[854]), .B(b[854]), .Z(n3767) );
  NANDN U3565 ( .A(n3766), .B(n3767), .Z(n1708) );
  AND U3566 ( .A(n1709), .B(n1708), .Z(n3768) );
  XOR U3567 ( .A(a[855]), .B(b[855]), .Z(n3769) );
  NANDN U3568 ( .A(n3768), .B(n3769), .Z(n1710) );
  AND U3569 ( .A(n1711), .B(n1710), .Z(n3770) );
  XOR U3570 ( .A(a[856]), .B(b[856]), .Z(n3771) );
  NANDN U3571 ( .A(n3770), .B(n3771), .Z(n1712) );
  AND U3572 ( .A(n1713), .B(n1712), .Z(n3772) );
  XOR U3573 ( .A(a[857]), .B(b[857]), .Z(n3773) );
  NANDN U3574 ( .A(n3772), .B(n3773), .Z(n1714) );
  AND U3575 ( .A(n1715), .B(n1714), .Z(n3774) );
  XOR U3576 ( .A(a[858]), .B(b[858]), .Z(n3775) );
  NANDN U3577 ( .A(n3774), .B(n3775), .Z(n1716) );
  AND U3578 ( .A(n1717), .B(n1716), .Z(n3776) );
  XOR U3579 ( .A(a[859]), .B(b[859]), .Z(n3777) );
  NANDN U3580 ( .A(n3776), .B(n3777), .Z(n1718) );
  AND U3581 ( .A(n1719), .B(n1718), .Z(n3780) );
  XOR U3582 ( .A(a[860]), .B(b[860]), .Z(n3781) );
  NANDN U3583 ( .A(n3780), .B(n3781), .Z(n1720) );
  AND U3584 ( .A(n1721), .B(n1720), .Z(n3782) );
  XOR U3585 ( .A(a[861]), .B(b[861]), .Z(n3783) );
  NANDN U3586 ( .A(n3782), .B(n3783), .Z(n1722) );
  AND U3587 ( .A(n1723), .B(n1722), .Z(n3784) );
  XOR U3588 ( .A(a[862]), .B(b[862]), .Z(n3785) );
  NANDN U3589 ( .A(n3784), .B(n3785), .Z(n1724) );
  AND U3590 ( .A(n1725), .B(n1724), .Z(n3786) );
  XOR U3591 ( .A(a[863]), .B(b[863]), .Z(n3787) );
  NANDN U3592 ( .A(n3786), .B(n3787), .Z(n1726) );
  AND U3593 ( .A(n1727), .B(n1726), .Z(n3788) );
  XOR U3594 ( .A(a[864]), .B(b[864]), .Z(n3789) );
  NANDN U3595 ( .A(n3788), .B(n3789), .Z(n1728) );
  AND U3596 ( .A(n1729), .B(n1728), .Z(n3790) );
  XOR U3597 ( .A(a[865]), .B(b[865]), .Z(n3791) );
  NANDN U3598 ( .A(n3790), .B(n3791), .Z(n1730) );
  AND U3599 ( .A(n1731), .B(n1730), .Z(n3792) );
  XOR U3600 ( .A(a[866]), .B(b[866]), .Z(n3793) );
  NANDN U3601 ( .A(n3792), .B(n3793), .Z(n1732) );
  AND U3602 ( .A(n1733), .B(n1732), .Z(n3794) );
  XOR U3603 ( .A(a[867]), .B(b[867]), .Z(n3795) );
  NANDN U3604 ( .A(n3794), .B(n3795), .Z(n1734) );
  AND U3605 ( .A(n1735), .B(n1734), .Z(n3796) );
  XOR U3606 ( .A(a[868]), .B(b[868]), .Z(n3797) );
  NANDN U3607 ( .A(n3796), .B(n3797), .Z(n1736) );
  AND U3608 ( .A(n1737), .B(n1736), .Z(n3798) );
  XOR U3609 ( .A(a[869]), .B(b[869]), .Z(n3799) );
  NANDN U3610 ( .A(n3798), .B(n3799), .Z(n1738) );
  AND U3611 ( .A(n1739), .B(n1738), .Z(n3802) );
  XOR U3612 ( .A(a[870]), .B(b[870]), .Z(n3803) );
  NANDN U3613 ( .A(n3802), .B(n3803), .Z(n1740) );
  AND U3614 ( .A(n1741), .B(n1740), .Z(n3804) );
  XOR U3615 ( .A(a[871]), .B(b[871]), .Z(n3805) );
  NANDN U3616 ( .A(n3804), .B(n3805), .Z(n1742) );
  AND U3617 ( .A(n1743), .B(n1742), .Z(n3806) );
  XOR U3618 ( .A(a[872]), .B(b[872]), .Z(n3807) );
  NANDN U3619 ( .A(n3806), .B(n3807), .Z(n1744) );
  AND U3620 ( .A(n1745), .B(n1744), .Z(n3808) );
  XOR U3621 ( .A(a[873]), .B(b[873]), .Z(n3809) );
  NANDN U3622 ( .A(n3808), .B(n3809), .Z(n1746) );
  AND U3623 ( .A(n1747), .B(n1746), .Z(n3810) );
  XOR U3624 ( .A(a[874]), .B(b[874]), .Z(n3811) );
  NANDN U3625 ( .A(n3810), .B(n3811), .Z(n1748) );
  AND U3626 ( .A(n1749), .B(n1748), .Z(n3812) );
  XOR U3627 ( .A(a[875]), .B(b[875]), .Z(n3813) );
  NANDN U3628 ( .A(n3812), .B(n3813), .Z(n1750) );
  AND U3629 ( .A(n1751), .B(n1750), .Z(n3814) );
  XOR U3630 ( .A(a[876]), .B(b[876]), .Z(n3815) );
  NANDN U3631 ( .A(n3814), .B(n3815), .Z(n1752) );
  AND U3632 ( .A(n1753), .B(n1752), .Z(n3816) );
  XOR U3633 ( .A(a[877]), .B(b[877]), .Z(n3817) );
  NANDN U3634 ( .A(n3816), .B(n3817), .Z(n1754) );
  AND U3635 ( .A(n1755), .B(n1754), .Z(n3818) );
  XOR U3636 ( .A(a[878]), .B(b[878]), .Z(n3819) );
  NANDN U3637 ( .A(n3818), .B(n3819), .Z(n1756) );
  AND U3638 ( .A(n1757), .B(n1756), .Z(n3820) );
  XOR U3639 ( .A(a[879]), .B(b[879]), .Z(n3821) );
  NANDN U3640 ( .A(n3820), .B(n3821), .Z(n1758) );
  AND U3641 ( .A(n1759), .B(n1758), .Z(n3824) );
  XOR U3642 ( .A(a[880]), .B(b[880]), .Z(n3825) );
  NANDN U3643 ( .A(n3824), .B(n3825), .Z(n1760) );
  AND U3644 ( .A(n1761), .B(n1760), .Z(n3826) );
  XOR U3645 ( .A(a[881]), .B(b[881]), .Z(n3827) );
  NANDN U3646 ( .A(n3826), .B(n3827), .Z(n1762) );
  AND U3647 ( .A(n1763), .B(n1762), .Z(n3828) );
  XOR U3648 ( .A(a[882]), .B(b[882]), .Z(n3829) );
  NANDN U3649 ( .A(n3828), .B(n3829), .Z(n1764) );
  AND U3650 ( .A(n1765), .B(n1764), .Z(n3830) );
  XOR U3651 ( .A(a[883]), .B(b[883]), .Z(n3831) );
  NANDN U3652 ( .A(n3830), .B(n3831), .Z(n1766) );
  AND U3653 ( .A(n1767), .B(n1766), .Z(n3832) );
  XOR U3654 ( .A(a[884]), .B(b[884]), .Z(n3833) );
  NANDN U3655 ( .A(n3832), .B(n3833), .Z(n1768) );
  AND U3656 ( .A(n1769), .B(n1768), .Z(n3834) );
  XOR U3657 ( .A(a[885]), .B(b[885]), .Z(n3835) );
  NANDN U3658 ( .A(n3834), .B(n3835), .Z(n1770) );
  AND U3659 ( .A(n1771), .B(n1770), .Z(n3836) );
  XOR U3660 ( .A(a[886]), .B(b[886]), .Z(n3837) );
  NANDN U3661 ( .A(n3836), .B(n3837), .Z(n1772) );
  AND U3662 ( .A(n1773), .B(n1772), .Z(n3838) );
  XOR U3663 ( .A(a[887]), .B(b[887]), .Z(n3839) );
  NANDN U3664 ( .A(n3838), .B(n3839), .Z(n1774) );
  AND U3665 ( .A(n1775), .B(n1774), .Z(n3840) );
  XOR U3666 ( .A(a[888]), .B(b[888]), .Z(n3841) );
  NANDN U3667 ( .A(n3840), .B(n3841), .Z(n1776) );
  AND U3668 ( .A(n1777), .B(n1776), .Z(n3842) );
  XOR U3669 ( .A(a[889]), .B(b[889]), .Z(n3843) );
  NANDN U3670 ( .A(n3842), .B(n3843), .Z(n1778) );
  AND U3671 ( .A(n1779), .B(n1778), .Z(n3846) );
  XOR U3672 ( .A(a[890]), .B(b[890]), .Z(n3847) );
  NANDN U3673 ( .A(n3846), .B(n3847), .Z(n1780) );
  AND U3674 ( .A(n1781), .B(n1780), .Z(n3848) );
  XOR U3675 ( .A(a[891]), .B(b[891]), .Z(n3849) );
  NANDN U3676 ( .A(n3848), .B(n3849), .Z(n1782) );
  AND U3677 ( .A(n1783), .B(n1782), .Z(n3850) );
  XOR U3678 ( .A(a[892]), .B(b[892]), .Z(n3851) );
  NANDN U3679 ( .A(n3850), .B(n3851), .Z(n1784) );
  AND U3680 ( .A(n1785), .B(n1784), .Z(n3852) );
  XOR U3681 ( .A(a[893]), .B(b[893]), .Z(n3853) );
  NANDN U3682 ( .A(n3852), .B(n3853), .Z(n1786) );
  AND U3683 ( .A(n1787), .B(n1786), .Z(n3854) );
  XOR U3684 ( .A(a[894]), .B(b[894]), .Z(n3855) );
  NANDN U3685 ( .A(n3854), .B(n3855), .Z(n1788) );
  AND U3686 ( .A(n1789), .B(n1788), .Z(n3856) );
  XOR U3687 ( .A(a[895]), .B(b[895]), .Z(n3857) );
  NANDN U3688 ( .A(n3856), .B(n3857), .Z(n1790) );
  AND U3689 ( .A(n1791), .B(n1790), .Z(n3858) );
  XOR U3690 ( .A(a[896]), .B(b[896]), .Z(n3859) );
  NANDN U3691 ( .A(n3858), .B(n3859), .Z(n1792) );
  AND U3692 ( .A(n1793), .B(n1792), .Z(n3860) );
  XOR U3693 ( .A(a[897]), .B(b[897]), .Z(n3861) );
  NANDN U3694 ( .A(n3860), .B(n3861), .Z(n1794) );
  AND U3695 ( .A(n1795), .B(n1794), .Z(n3862) );
  XOR U3696 ( .A(a[898]), .B(b[898]), .Z(n3863) );
  NANDN U3697 ( .A(n3862), .B(n3863), .Z(n1796) );
  AND U3698 ( .A(n1797), .B(n1796), .Z(n3864) );
  XOR U3699 ( .A(a[899]), .B(b[899]), .Z(n3865) );
  NANDN U3700 ( .A(n3864), .B(n3865), .Z(n1798) );
  AND U3701 ( .A(n1799), .B(n1798), .Z(n3870) );
  XOR U3702 ( .A(a[900]), .B(b[900]), .Z(n3871) );
  NANDN U3703 ( .A(n3870), .B(n3871), .Z(n1800) );
  AND U3704 ( .A(n1801), .B(n1800), .Z(n3872) );
  XOR U3705 ( .A(a[901]), .B(b[901]), .Z(n3873) );
  NANDN U3706 ( .A(n3872), .B(n3873), .Z(n1802) );
  AND U3707 ( .A(n1803), .B(n1802), .Z(n3874) );
  XOR U3708 ( .A(a[902]), .B(b[902]), .Z(n3875) );
  NANDN U3709 ( .A(n3874), .B(n3875), .Z(n1804) );
  AND U3710 ( .A(n1805), .B(n1804), .Z(n3876) );
  XOR U3711 ( .A(a[903]), .B(b[903]), .Z(n3877) );
  NANDN U3712 ( .A(n3876), .B(n3877), .Z(n1806) );
  AND U3713 ( .A(n1807), .B(n1806), .Z(n3878) );
  XOR U3714 ( .A(a[904]), .B(b[904]), .Z(n3879) );
  NANDN U3715 ( .A(n3878), .B(n3879), .Z(n1808) );
  AND U3716 ( .A(n1809), .B(n1808), .Z(n3880) );
  XOR U3717 ( .A(a[905]), .B(b[905]), .Z(n3881) );
  NANDN U3718 ( .A(n3880), .B(n3881), .Z(n1810) );
  AND U3719 ( .A(n1811), .B(n1810), .Z(n3882) );
  XOR U3720 ( .A(a[906]), .B(b[906]), .Z(n3883) );
  NANDN U3721 ( .A(n3882), .B(n3883), .Z(n1812) );
  AND U3722 ( .A(n1813), .B(n1812), .Z(n3884) );
  XOR U3723 ( .A(a[907]), .B(b[907]), .Z(n3885) );
  NANDN U3724 ( .A(n3884), .B(n3885), .Z(n1814) );
  AND U3725 ( .A(n1815), .B(n1814), .Z(n3886) );
  XOR U3726 ( .A(a[908]), .B(b[908]), .Z(n3887) );
  NANDN U3727 ( .A(n3886), .B(n3887), .Z(n1816) );
  AND U3728 ( .A(n1817), .B(n1816), .Z(n3888) );
  XOR U3729 ( .A(a[909]), .B(b[909]), .Z(n3889) );
  NANDN U3730 ( .A(n3888), .B(n3889), .Z(n1818) );
  AND U3731 ( .A(n1819), .B(n1818), .Z(n3892) );
  XOR U3732 ( .A(a[910]), .B(b[910]), .Z(n3893) );
  NANDN U3733 ( .A(n3892), .B(n3893), .Z(n1820) );
  AND U3734 ( .A(n1821), .B(n1820), .Z(n3894) );
  XOR U3735 ( .A(a[911]), .B(b[911]), .Z(n3895) );
  NANDN U3736 ( .A(n3894), .B(n3895), .Z(n1822) );
  AND U3737 ( .A(n1823), .B(n1822), .Z(n3896) );
  XOR U3738 ( .A(a[912]), .B(b[912]), .Z(n3897) );
  NANDN U3739 ( .A(n3896), .B(n3897), .Z(n1824) );
  AND U3740 ( .A(n1825), .B(n1824), .Z(n3898) );
  XOR U3741 ( .A(a[913]), .B(b[913]), .Z(n3899) );
  NANDN U3742 ( .A(n3898), .B(n3899), .Z(n1826) );
  AND U3743 ( .A(n1827), .B(n1826), .Z(n3900) );
  XOR U3744 ( .A(a[914]), .B(b[914]), .Z(n3901) );
  NANDN U3745 ( .A(n3900), .B(n3901), .Z(n1828) );
  AND U3746 ( .A(n1829), .B(n1828), .Z(n3902) );
  XOR U3747 ( .A(a[915]), .B(b[915]), .Z(n3903) );
  NANDN U3748 ( .A(n3902), .B(n3903), .Z(n1830) );
  AND U3749 ( .A(n1831), .B(n1830), .Z(n3904) );
  XOR U3750 ( .A(a[916]), .B(b[916]), .Z(n3905) );
  NANDN U3751 ( .A(n3904), .B(n3905), .Z(n1832) );
  AND U3752 ( .A(n1833), .B(n1832), .Z(n3906) );
  XOR U3753 ( .A(a[917]), .B(b[917]), .Z(n3907) );
  NANDN U3754 ( .A(n3906), .B(n3907), .Z(n1834) );
  AND U3755 ( .A(n1835), .B(n1834), .Z(n3908) );
  XOR U3756 ( .A(a[918]), .B(b[918]), .Z(n3909) );
  NANDN U3757 ( .A(n3908), .B(n3909), .Z(n1836) );
  AND U3758 ( .A(n1837), .B(n1836), .Z(n3910) );
  XOR U3759 ( .A(a[919]), .B(b[919]), .Z(n3911) );
  NANDN U3760 ( .A(n3910), .B(n3911), .Z(n1838) );
  AND U3761 ( .A(n1839), .B(n1838), .Z(n3914) );
  XOR U3762 ( .A(a[920]), .B(b[920]), .Z(n3915) );
  NANDN U3763 ( .A(n3914), .B(n3915), .Z(n1840) );
  AND U3764 ( .A(n1841), .B(n1840), .Z(n3916) );
  XOR U3765 ( .A(a[921]), .B(b[921]), .Z(n3917) );
  NANDN U3766 ( .A(n3916), .B(n3917), .Z(n1842) );
  AND U3767 ( .A(n1843), .B(n1842), .Z(n3918) );
  XOR U3768 ( .A(a[922]), .B(b[922]), .Z(n3919) );
  NANDN U3769 ( .A(n3918), .B(n3919), .Z(n1844) );
  AND U3770 ( .A(n1845), .B(n1844), .Z(n3920) );
  XOR U3771 ( .A(a[923]), .B(b[923]), .Z(n3921) );
  NANDN U3772 ( .A(n3920), .B(n3921), .Z(n1846) );
  AND U3773 ( .A(n1847), .B(n1846), .Z(n3922) );
  XOR U3774 ( .A(a[924]), .B(b[924]), .Z(n3923) );
  NANDN U3775 ( .A(n3922), .B(n3923), .Z(n1848) );
  AND U3776 ( .A(n1849), .B(n1848), .Z(n3924) );
  XOR U3777 ( .A(a[925]), .B(b[925]), .Z(n3925) );
  NANDN U3778 ( .A(n3924), .B(n3925), .Z(n1850) );
  AND U3779 ( .A(n1851), .B(n1850), .Z(n3926) );
  XOR U3780 ( .A(a[926]), .B(b[926]), .Z(n3927) );
  NANDN U3781 ( .A(n3926), .B(n3927), .Z(n1852) );
  AND U3782 ( .A(n1853), .B(n1852), .Z(n3928) );
  XOR U3783 ( .A(a[927]), .B(b[927]), .Z(n3929) );
  NANDN U3784 ( .A(n3928), .B(n3929), .Z(n1854) );
  AND U3785 ( .A(n1855), .B(n1854), .Z(n3930) );
  XOR U3786 ( .A(a[928]), .B(b[928]), .Z(n3931) );
  NANDN U3787 ( .A(n3930), .B(n3931), .Z(n1856) );
  AND U3788 ( .A(n1857), .B(n1856), .Z(n3932) );
  XOR U3789 ( .A(a[929]), .B(b[929]), .Z(n3933) );
  NANDN U3790 ( .A(n3932), .B(n3933), .Z(n1858) );
  AND U3791 ( .A(n1859), .B(n1858), .Z(n3936) );
  XOR U3792 ( .A(a[930]), .B(b[930]), .Z(n3937) );
  NANDN U3793 ( .A(n3936), .B(n3937), .Z(n1860) );
  AND U3794 ( .A(n1861), .B(n1860), .Z(n3938) );
  XOR U3795 ( .A(a[931]), .B(b[931]), .Z(n3939) );
  NANDN U3796 ( .A(n3938), .B(n3939), .Z(n1862) );
  AND U3797 ( .A(n1863), .B(n1862), .Z(n3940) );
  XOR U3798 ( .A(a[932]), .B(b[932]), .Z(n3941) );
  NANDN U3799 ( .A(n3940), .B(n3941), .Z(n1864) );
  AND U3800 ( .A(n1865), .B(n1864), .Z(n3942) );
  XOR U3801 ( .A(a[933]), .B(b[933]), .Z(n3943) );
  NANDN U3802 ( .A(n3942), .B(n3943), .Z(n1866) );
  AND U3803 ( .A(n1867), .B(n1866), .Z(n3944) );
  XOR U3804 ( .A(a[934]), .B(b[934]), .Z(n3945) );
  NANDN U3805 ( .A(n3944), .B(n3945), .Z(n1868) );
  AND U3806 ( .A(n1869), .B(n1868), .Z(n3946) );
  XOR U3807 ( .A(a[935]), .B(b[935]), .Z(n3947) );
  NANDN U3808 ( .A(n3946), .B(n3947), .Z(n1870) );
  AND U3809 ( .A(n1871), .B(n1870), .Z(n3948) );
  XOR U3810 ( .A(a[936]), .B(b[936]), .Z(n3949) );
  NANDN U3811 ( .A(n3948), .B(n3949), .Z(n1872) );
  AND U3812 ( .A(n1873), .B(n1872), .Z(n3950) );
  XOR U3813 ( .A(a[937]), .B(b[937]), .Z(n3951) );
  NANDN U3814 ( .A(n3950), .B(n3951), .Z(n1874) );
  AND U3815 ( .A(n1875), .B(n1874), .Z(n3952) );
  XOR U3816 ( .A(a[938]), .B(b[938]), .Z(n3953) );
  NANDN U3817 ( .A(n3952), .B(n3953), .Z(n1876) );
  AND U3818 ( .A(n1877), .B(n1876), .Z(n3954) );
  XOR U3819 ( .A(a[939]), .B(b[939]), .Z(n3955) );
  NANDN U3820 ( .A(n3954), .B(n3955), .Z(n1878) );
  AND U3821 ( .A(n1879), .B(n1878), .Z(n3958) );
  XOR U3822 ( .A(a[940]), .B(b[940]), .Z(n3959) );
  NANDN U3823 ( .A(n3958), .B(n3959), .Z(n1880) );
  AND U3824 ( .A(n1881), .B(n1880), .Z(n3960) );
  XOR U3825 ( .A(a[941]), .B(b[941]), .Z(n3961) );
  NANDN U3826 ( .A(n3960), .B(n3961), .Z(n1882) );
  AND U3827 ( .A(n1883), .B(n1882), .Z(n3962) );
  XOR U3828 ( .A(a[942]), .B(b[942]), .Z(n3963) );
  NANDN U3829 ( .A(n3962), .B(n3963), .Z(n1884) );
  AND U3830 ( .A(n1885), .B(n1884), .Z(n3964) );
  XOR U3831 ( .A(a[943]), .B(b[943]), .Z(n3965) );
  NANDN U3832 ( .A(n3964), .B(n3965), .Z(n1886) );
  AND U3833 ( .A(n1887), .B(n1886), .Z(n3966) );
  XOR U3834 ( .A(a[944]), .B(b[944]), .Z(n3967) );
  NANDN U3835 ( .A(n3966), .B(n3967), .Z(n1888) );
  AND U3836 ( .A(n1889), .B(n1888), .Z(n3968) );
  XOR U3837 ( .A(a[945]), .B(b[945]), .Z(n3969) );
  NANDN U3838 ( .A(n3968), .B(n3969), .Z(n1890) );
  AND U3839 ( .A(n1891), .B(n1890), .Z(n3970) );
  XOR U3840 ( .A(a[946]), .B(b[946]), .Z(n3971) );
  NANDN U3841 ( .A(n3970), .B(n3971), .Z(n1892) );
  AND U3842 ( .A(n1893), .B(n1892), .Z(n3972) );
  XOR U3843 ( .A(a[947]), .B(b[947]), .Z(n3973) );
  NANDN U3844 ( .A(n3972), .B(n3973), .Z(n1894) );
  AND U3845 ( .A(n1895), .B(n1894), .Z(n3974) );
  XOR U3846 ( .A(a[948]), .B(b[948]), .Z(n3975) );
  NANDN U3847 ( .A(n3974), .B(n3975), .Z(n1896) );
  AND U3848 ( .A(n1897), .B(n1896), .Z(n3976) );
  XOR U3849 ( .A(a[949]), .B(b[949]), .Z(n3977) );
  NANDN U3850 ( .A(n3976), .B(n3977), .Z(n1898) );
  AND U3851 ( .A(n1899), .B(n1898), .Z(n3980) );
  XOR U3852 ( .A(a[950]), .B(b[950]), .Z(n3981) );
  NANDN U3853 ( .A(n3980), .B(n3981), .Z(n1900) );
  AND U3854 ( .A(n1901), .B(n1900), .Z(n3982) );
  XOR U3855 ( .A(a[951]), .B(b[951]), .Z(n3983) );
  NANDN U3856 ( .A(n3982), .B(n3983), .Z(n1902) );
  AND U3857 ( .A(n1903), .B(n1902), .Z(n3984) );
  XOR U3858 ( .A(a[952]), .B(b[952]), .Z(n3985) );
  NANDN U3859 ( .A(n3984), .B(n3985), .Z(n1904) );
  AND U3860 ( .A(n1905), .B(n1904), .Z(n3986) );
  XOR U3861 ( .A(a[953]), .B(b[953]), .Z(n3987) );
  NANDN U3862 ( .A(n3986), .B(n3987), .Z(n1906) );
  AND U3863 ( .A(n1907), .B(n1906), .Z(n3988) );
  XOR U3864 ( .A(a[954]), .B(b[954]), .Z(n3989) );
  NANDN U3865 ( .A(n3988), .B(n3989), .Z(n1908) );
  AND U3866 ( .A(n1909), .B(n1908), .Z(n3990) );
  XOR U3867 ( .A(a[955]), .B(b[955]), .Z(n3991) );
  NANDN U3868 ( .A(n3990), .B(n3991), .Z(n1910) );
  AND U3869 ( .A(n1911), .B(n1910), .Z(n3992) );
  XOR U3870 ( .A(a[956]), .B(b[956]), .Z(n3993) );
  NANDN U3871 ( .A(n3992), .B(n3993), .Z(n1912) );
  AND U3872 ( .A(n1913), .B(n1912), .Z(n3994) );
  XOR U3873 ( .A(a[957]), .B(b[957]), .Z(n3995) );
  NANDN U3874 ( .A(n3994), .B(n3995), .Z(n1914) );
  AND U3875 ( .A(n1915), .B(n1914), .Z(n3996) );
  XOR U3876 ( .A(a[958]), .B(b[958]), .Z(n3997) );
  NANDN U3877 ( .A(n3996), .B(n3997), .Z(n1916) );
  AND U3878 ( .A(n1917), .B(n1916), .Z(n3998) );
  XOR U3879 ( .A(a[959]), .B(b[959]), .Z(n3999) );
  NANDN U3880 ( .A(n3998), .B(n3999), .Z(n1918) );
  AND U3881 ( .A(n1919), .B(n1918), .Z(n4002) );
  XOR U3882 ( .A(a[960]), .B(b[960]), .Z(n4003) );
  NANDN U3883 ( .A(n4002), .B(n4003), .Z(n1920) );
  AND U3884 ( .A(n1921), .B(n1920), .Z(n4004) );
  XOR U3885 ( .A(a[961]), .B(b[961]), .Z(n4005) );
  NANDN U3886 ( .A(n4004), .B(n4005), .Z(n1922) );
  AND U3887 ( .A(n1923), .B(n1922), .Z(n4006) );
  XOR U3888 ( .A(a[962]), .B(b[962]), .Z(n4007) );
  NANDN U3889 ( .A(n4006), .B(n4007), .Z(n1924) );
  AND U3890 ( .A(n1925), .B(n1924), .Z(n4008) );
  XOR U3891 ( .A(a[963]), .B(b[963]), .Z(n4009) );
  NANDN U3892 ( .A(n4008), .B(n4009), .Z(n1926) );
  AND U3893 ( .A(n1927), .B(n1926), .Z(n4010) );
  XOR U3894 ( .A(a[964]), .B(b[964]), .Z(n4011) );
  NANDN U3895 ( .A(n4010), .B(n4011), .Z(n1928) );
  AND U3896 ( .A(n1929), .B(n1928), .Z(n4012) );
  XOR U3897 ( .A(a[965]), .B(b[965]), .Z(n4013) );
  NANDN U3898 ( .A(n4012), .B(n4013), .Z(n1930) );
  AND U3899 ( .A(n1931), .B(n1930), .Z(n4014) );
  XOR U3900 ( .A(a[966]), .B(b[966]), .Z(n4015) );
  NANDN U3901 ( .A(n4014), .B(n4015), .Z(n1932) );
  AND U3902 ( .A(n1933), .B(n1932), .Z(n4016) );
  XOR U3903 ( .A(a[967]), .B(b[967]), .Z(n4017) );
  NANDN U3904 ( .A(n4016), .B(n4017), .Z(n1934) );
  AND U3905 ( .A(n1935), .B(n1934), .Z(n4018) );
  XOR U3906 ( .A(a[968]), .B(b[968]), .Z(n4019) );
  NANDN U3907 ( .A(n4018), .B(n4019), .Z(n1936) );
  AND U3908 ( .A(n1937), .B(n1936), .Z(n4020) );
  XOR U3909 ( .A(a[969]), .B(b[969]), .Z(n4021) );
  NANDN U3910 ( .A(n4020), .B(n4021), .Z(n1938) );
  AND U3911 ( .A(n1939), .B(n1938), .Z(n4024) );
  XOR U3912 ( .A(a[970]), .B(b[970]), .Z(n4025) );
  NANDN U3913 ( .A(n4024), .B(n4025), .Z(n1940) );
  AND U3914 ( .A(n1941), .B(n1940), .Z(n4026) );
  XOR U3915 ( .A(a[971]), .B(b[971]), .Z(n4027) );
  NANDN U3916 ( .A(n4026), .B(n4027), .Z(n1942) );
  AND U3917 ( .A(n1943), .B(n1942), .Z(n4028) );
  XOR U3918 ( .A(a[972]), .B(b[972]), .Z(n4029) );
  NANDN U3919 ( .A(n4028), .B(n4029), .Z(n1944) );
  AND U3920 ( .A(n1945), .B(n1944), .Z(n4030) );
  XOR U3921 ( .A(a[973]), .B(b[973]), .Z(n4031) );
  NANDN U3922 ( .A(n4030), .B(n4031), .Z(n1946) );
  AND U3923 ( .A(n1947), .B(n1946), .Z(n4032) );
  XOR U3924 ( .A(a[974]), .B(b[974]), .Z(n4033) );
  NANDN U3925 ( .A(n4032), .B(n4033), .Z(n1948) );
  AND U3926 ( .A(n1949), .B(n1948), .Z(n4034) );
  XOR U3927 ( .A(a[975]), .B(b[975]), .Z(n4035) );
  NANDN U3928 ( .A(n4034), .B(n4035), .Z(n1950) );
  AND U3929 ( .A(n1951), .B(n1950), .Z(n4036) );
  XOR U3930 ( .A(a[976]), .B(b[976]), .Z(n4037) );
  NANDN U3931 ( .A(n4036), .B(n4037), .Z(n1952) );
  AND U3932 ( .A(n1953), .B(n1952), .Z(n4038) );
  XOR U3933 ( .A(a[977]), .B(b[977]), .Z(n4039) );
  NANDN U3934 ( .A(n4038), .B(n4039), .Z(n1954) );
  AND U3935 ( .A(n1955), .B(n1954), .Z(n4040) );
  XOR U3936 ( .A(a[978]), .B(b[978]), .Z(n4041) );
  NANDN U3937 ( .A(n4040), .B(n4041), .Z(n1956) );
  AND U3938 ( .A(n1957), .B(n1956), .Z(n4042) );
  XOR U3939 ( .A(a[979]), .B(b[979]), .Z(n4043) );
  NANDN U3940 ( .A(n4042), .B(n4043), .Z(n1958) );
  AND U3941 ( .A(n1959), .B(n1958), .Z(n4046) );
  XOR U3942 ( .A(a[980]), .B(b[980]), .Z(n4047) );
  NANDN U3943 ( .A(n4046), .B(n4047), .Z(n1960) );
  AND U3944 ( .A(n1961), .B(n1960), .Z(n4048) );
  XOR U3945 ( .A(a[981]), .B(b[981]), .Z(n4049) );
  NANDN U3946 ( .A(n4048), .B(n4049), .Z(n1962) );
  AND U3947 ( .A(n1963), .B(n1962), .Z(n4050) );
  XOR U3948 ( .A(a[982]), .B(b[982]), .Z(n4051) );
  NANDN U3949 ( .A(n4050), .B(n4051), .Z(n1964) );
  AND U3950 ( .A(n1965), .B(n1964), .Z(n4052) );
  XOR U3951 ( .A(a[983]), .B(b[983]), .Z(n4053) );
  NANDN U3952 ( .A(n4052), .B(n4053), .Z(n1966) );
  AND U3953 ( .A(n1967), .B(n1966), .Z(n4054) );
  XOR U3954 ( .A(a[984]), .B(b[984]), .Z(n4055) );
  NANDN U3955 ( .A(n4054), .B(n4055), .Z(n1968) );
  AND U3956 ( .A(n1969), .B(n1968), .Z(n4056) );
  XOR U3957 ( .A(a[985]), .B(b[985]), .Z(n4057) );
  NANDN U3958 ( .A(n4056), .B(n4057), .Z(n1970) );
  AND U3959 ( .A(n1971), .B(n1970), .Z(n4058) );
  XOR U3960 ( .A(a[986]), .B(b[986]), .Z(n4059) );
  NANDN U3961 ( .A(n4058), .B(n4059), .Z(n1972) );
  AND U3962 ( .A(n1973), .B(n1972), .Z(n4060) );
  XOR U3963 ( .A(a[987]), .B(b[987]), .Z(n4061) );
  NANDN U3964 ( .A(n4060), .B(n4061), .Z(n1974) );
  AND U3965 ( .A(n1975), .B(n1974), .Z(n4062) );
  XOR U3966 ( .A(a[988]), .B(b[988]), .Z(n4063) );
  NANDN U3967 ( .A(n4062), .B(n4063), .Z(n1976) );
  AND U3968 ( .A(n1977), .B(n1976), .Z(n4064) );
  XOR U3969 ( .A(a[989]), .B(b[989]), .Z(n4065) );
  NANDN U3970 ( .A(n4064), .B(n4065), .Z(n1978) );
  AND U3971 ( .A(n1979), .B(n1978), .Z(n4068) );
  XOR U3972 ( .A(a[990]), .B(b[990]), .Z(n4069) );
  NANDN U3973 ( .A(n4068), .B(n4069), .Z(n1980) );
  AND U3974 ( .A(n1981), .B(n1980), .Z(n4070) );
  XOR U3975 ( .A(a[991]), .B(b[991]), .Z(n4071) );
  NANDN U3976 ( .A(n4070), .B(n4071), .Z(n1982) );
  AND U3977 ( .A(n1983), .B(n1982), .Z(n4072) );
  XOR U3978 ( .A(a[992]), .B(b[992]), .Z(n4073) );
  NANDN U3979 ( .A(n4072), .B(n4073), .Z(n1984) );
  AND U3980 ( .A(n1985), .B(n1984), .Z(n4074) );
  XOR U3981 ( .A(a[993]), .B(b[993]), .Z(n4075) );
  NANDN U3982 ( .A(n4074), .B(n4075), .Z(n1986) );
  AND U3983 ( .A(n1987), .B(n1986), .Z(n4076) );
  XOR U3984 ( .A(a[994]), .B(b[994]), .Z(n4077) );
  NANDN U3985 ( .A(n4076), .B(n4077), .Z(n1988) );
  AND U3986 ( .A(n1989), .B(n1988), .Z(n4078) );
  XOR U3987 ( .A(a[995]), .B(b[995]), .Z(n4079) );
  NANDN U3988 ( .A(n4078), .B(n4079), .Z(n1990) );
  AND U3989 ( .A(n1991), .B(n1990), .Z(n4080) );
  XOR U3990 ( .A(a[996]), .B(b[996]), .Z(n4081) );
  NANDN U3991 ( .A(n4080), .B(n4081), .Z(n1992) );
  AND U3992 ( .A(n1993), .B(n1992), .Z(n4082) );
  XOR U3993 ( .A(a[997]), .B(b[997]), .Z(n4083) );
  NANDN U3994 ( .A(n4082), .B(n4083), .Z(n1994) );
  AND U3995 ( .A(n1995), .B(n1994), .Z(n4084) );
  XOR U3996 ( .A(a[998]), .B(b[998]), .Z(n4085) );
  NANDN U3997 ( .A(n4084), .B(n4085), .Z(n1996) );
  AND U3998 ( .A(n1997), .B(n1996), .Z(n4086) );
  OR U3999 ( .A(n4087), .B(n4086), .Z(n1998) );
  AND U4000 ( .A(n1999), .B(n1998), .Z(n2001) );
  XNOR U4001 ( .A(n2000), .B(n2001), .Z(c[1000]) );
  XOR U4002 ( .A(a[1001]), .B(b[1001]), .Z(n2004) );
  NAND U4003 ( .A(b[1000]), .B(a[1000]), .Z(n2003) );
  NANDN U4004 ( .A(n2001), .B(n2000), .Z(n2002) );
  AND U4005 ( .A(n2003), .B(n2002), .Z(n2005) );
  XNOR U4006 ( .A(n2004), .B(n2005), .Z(c[1001]) );
  XOR U4007 ( .A(a[1002]), .B(b[1002]), .Z(n2008) );
  NAND U4008 ( .A(b[1001]), .B(a[1001]), .Z(n2007) );
  NANDN U4009 ( .A(n2005), .B(n2004), .Z(n2006) );
  AND U4010 ( .A(n2007), .B(n2006), .Z(n2009) );
  XNOR U4011 ( .A(n2008), .B(n2009), .Z(c[1002]) );
  XOR U4012 ( .A(a[1003]), .B(b[1003]), .Z(n2012) );
  NAND U4013 ( .A(b[1002]), .B(a[1002]), .Z(n2011) );
  NANDN U4014 ( .A(n2009), .B(n2008), .Z(n2010) );
  AND U4015 ( .A(n2011), .B(n2010), .Z(n2013) );
  XNOR U4016 ( .A(n2012), .B(n2013), .Z(c[1003]) );
  XOR U4017 ( .A(a[1004]), .B(b[1004]), .Z(n2016) );
  NAND U4018 ( .A(b[1003]), .B(a[1003]), .Z(n2015) );
  NANDN U4019 ( .A(n2013), .B(n2012), .Z(n2014) );
  AND U4020 ( .A(n2015), .B(n2014), .Z(n2017) );
  XNOR U4021 ( .A(n2016), .B(n2017), .Z(c[1004]) );
  XOR U4022 ( .A(a[1005]), .B(b[1005]), .Z(n2020) );
  NAND U4023 ( .A(b[1004]), .B(a[1004]), .Z(n2019) );
  NANDN U4024 ( .A(n2017), .B(n2016), .Z(n2018) );
  AND U4025 ( .A(n2019), .B(n2018), .Z(n2021) );
  XNOR U4026 ( .A(n2020), .B(n2021), .Z(c[1005]) );
  XOR U4027 ( .A(a[1006]), .B(b[1006]), .Z(n2024) );
  NAND U4028 ( .A(b[1005]), .B(a[1005]), .Z(n2023) );
  NANDN U4029 ( .A(n2021), .B(n2020), .Z(n2022) );
  AND U4030 ( .A(n2023), .B(n2022), .Z(n2025) );
  XNOR U4031 ( .A(n2024), .B(n2025), .Z(c[1006]) );
  XOR U4032 ( .A(a[1007]), .B(b[1007]), .Z(n2028) );
  NAND U4033 ( .A(b[1006]), .B(a[1006]), .Z(n2027) );
  NANDN U4034 ( .A(n2025), .B(n2024), .Z(n2026) );
  AND U4035 ( .A(n2027), .B(n2026), .Z(n2029) );
  XNOR U4036 ( .A(n2028), .B(n2029), .Z(c[1007]) );
  XOR U4037 ( .A(a[1008]), .B(b[1008]), .Z(n2032) );
  NAND U4038 ( .A(b[1007]), .B(a[1007]), .Z(n2031) );
  NANDN U4039 ( .A(n2029), .B(n2028), .Z(n2030) );
  AND U4040 ( .A(n2031), .B(n2030), .Z(n2033) );
  XNOR U4041 ( .A(n2032), .B(n2033), .Z(c[1008]) );
  XOR U4042 ( .A(a[1009]), .B(b[1009]), .Z(n2038) );
  NAND U4043 ( .A(b[1008]), .B(a[1008]), .Z(n2035) );
  NANDN U4044 ( .A(n2033), .B(n2032), .Z(n2034) );
  AND U4045 ( .A(n2035), .B(n2034), .Z(n2039) );
  XNOR U4046 ( .A(n2038), .B(n2039), .Z(c[1009]) );
  XNOR U4047 ( .A(n2037), .B(n2036), .Z(c[100]) );
  XOR U4048 ( .A(a[1010]), .B(b[1010]), .Z(n2042) );
  NAND U4049 ( .A(b[1009]), .B(a[1009]), .Z(n2041) );
  NANDN U4050 ( .A(n2039), .B(n2038), .Z(n2040) );
  AND U4051 ( .A(n2041), .B(n2040), .Z(n2043) );
  XNOR U4052 ( .A(n2042), .B(n2043), .Z(c[1010]) );
  XOR U4053 ( .A(a[1011]), .B(b[1011]), .Z(n2046) );
  NAND U4054 ( .A(b[1010]), .B(a[1010]), .Z(n2045) );
  NANDN U4055 ( .A(n2043), .B(n2042), .Z(n2044) );
  AND U4056 ( .A(n2045), .B(n2044), .Z(n2047) );
  XNOR U4057 ( .A(n2046), .B(n2047), .Z(c[1011]) );
  XOR U4058 ( .A(a[1012]), .B(b[1012]), .Z(n2050) );
  NAND U4059 ( .A(b[1011]), .B(a[1011]), .Z(n2049) );
  NANDN U4060 ( .A(n2047), .B(n2046), .Z(n2048) );
  AND U4061 ( .A(n2049), .B(n2048), .Z(n2051) );
  XNOR U4062 ( .A(n2050), .B(n2051), .Z(c[1012]) );
  XOR U4063 ( .A(a[1013]), .B(b[1013]), .Z(n2054) );
  NAND U4064 ( .A(b[1012]), .B(a[1012]), .Z(n2053) );
  NANDN U4065 ( .A(n2051), .B(n2050), .Z(n2052) );
  AND U4066 ( .A(n2053), .B(n2052), .Z(n2055) );
  XNOR U4067 ( .A(n2054), .B(n2055), .Z(c[1013]) );
  XOR U4068 ( .A(a[1014]), .B(b[1014]), .Z(n2058) );
  NAND U4069 ( .A(b[1013]), .B(a[1013]), .Z(n2057) );
  NANDN U4070 ( .A(n2055), .B(n2054), .Z(n2056) );
  AND U4071 ( .A(n2057), .B(n2056), .Z(n2059) );
  XNOR U4072 ( .A(n2058), .B(n2059), .Z(c[1014]) );
  XOR U4073 ( .A(a[1015]), .B(b[1015]), .Z(n2062) );
  NAND U4074 ( .A(b[1014]), .B(a[1014]), .Z(n2061) );
  NANDN U4075 ( .A(n2059), .B(n2058), .Z(n2060) );
  AND U4076 ( .A(n2061), .B(n2060), .Z(n2063) );
  XNOR U4077 ( .A(n2062), .B(n2063), .Z(c[1015]) );
  XOR U4078 ( .A(a[1016]), .B(b[1016]), .Z(n2066) );
  NAND U4079 ( .A(b[1015]), .B(a[1015]), .Z(n2065) );
  NANDN U4080 ( .A(n2063), .B(n2062), .Z(n2064) );
  AND U4081 ( .A(n2065), .B(n2064), .Z(n2067) );
  XNOR U4082 ( .A(n2066), .B(n2067), .Z(c[1016]) );
  XOR U4083 ( .A(a[1017]), .B(b[1017]), .Z(n2070) );
  NAND U4084 ( .A(b[1016]), .B(a[1016]), .Z(n2069) );
  NANDN U4085 ( .A(n2067), .B(n2066), .Z(n2068) );
  AND U4086 ( .A(n2069), .B(n2068), .Z(n2071) );
  XNOR U4087 ( .A(n2070), .B(n2071), .Z(c[1017]) );
  XOR U4088 ( .A(a[1018]), .B(b[1018]), .Z(n2074) );
  NAND U4089 ( .A(b[1017]), .B(a[1017]), .Z(n2073) );
  NANDN U4090 ( .A(n2071), .B(n2070), .Z(n2072) );
  AND U4091 ( .A(n2073), .B(n2072), .Z(n2075) );
  XNOR U4092 ( .A(n2074), .B(n2075), .Z(c[1018]) );
  XOR U4093 ( .A(a[1019]), .B(b[1019]), .Z(n2080) );
  NAND U4094 ( .A(b[1018]), .B(a[1018]), .Z(n2077) );
  NANDN U4095 ( .A(n2075), .B(n2074), .Z(n2076) );
  AND U4096 ( .A(n2077), .B(n2076), .Z(n2081) );
  XNOR U4097 ( .A(n2080), .B(n2081), .Z(c[1019]) );
  XNOR U4098 ( .A(n2079), .B(n2078), .Z(c[101]) );
  XOR U4099 ( .A(a[1020]), .B(b[1020]), .Z(n2084) );
  NAND U4100 ( .A(b[1019]), .B(a[1019]), .Z(n2083) );
  NANDN U4101 ( .A(n2081), .B(n2080), .Z(n2082) );
  AND U4102 ( .A(n2083), .B(n2082), .Z(n2085) );
  XNOR U4103 ( .A(n2084), .B(n2085), .Z(c[1020]) );
  XOR U4104 ( .A(a[1021]), .B(b[1021]), .Z(n2088) );
  NAND U4105 ( .A(b[1020]), .B(a[1020]), .Z(n2087) );
  NANDN U4106 ( .A(n2085), .B(n2084), .Z(n2086) );
  AND U4107 ( .A(n2087), .B(n2086), .Z(n2089) );
  XNOR U4108 ( .A(n2088), .B(n2089), .Z(c[1021]) );
  XNOR U4109 ( .A(a[1022]), .B(b[1022]), .Z(n2093) );
  NAND U4110 ( .A(b[1021]), .B(a[1021]), .Z(n2091) );
  NANDN U4111 ( .A(n2089), .B(n2088), .Z(n2090) );
  AND U4112 ( .A(n2091), .B(n2090), .Z(n2092) );
  XOR U4113 ( .A(n2093), .B(n2092), .Z(c[1022]) );
  OR U4114 ( .A(n2093), .B(n2092), .Z(n2095) );
  NAND U4115 ( .A(a[1022]), .B(b[1022]), .Z(n2094) );
  NAND U4116 ( .A(n2095), .B(n2094), .Z(n2096) );
  XNOR U4117 ( .A(a[1023]), .B(n2096), .Z(n2097) );
  XNOR U4118 ( .A(b[1023]), .B(n2097), .Z(c[1023]) );
  XNOR U4119 ( .A(n2099), .B(n2098), .Z(c[102]) );
  XNOR U4120 ( .A(n2101), .B(n2100), .Z(c[103]) );
  XNOR U4121 ( .A(n2103), .B(n2102), .Z(c[104]) );
  XNOR U4122 ( .A(n2105), .B(n2104), .Z(c[105]) );
  XNOR U4123 ( .A(n2107), .B(n2106), .Z(c[106]) );
  XNOR U4124 ( .A(n2109), .B(n2108), .Z(c[107]) );
  XNOR U4125 ( .A(n2111), .B(n2110), .Z(c[108]) );
  XNOR U4126 ( .A(n2113), .B(n2112), .Z(c[109]) );
  XNOR U4127 ( .A(n2115), .B(n2114), .Z(c[10]) );
  XNOR U4128 ( .A(n2117), .B(n2116), .Z(c[110]) );
  XNOR U4129 ( .A(n2119), .B(n2118), .Z(c[111]) );
  XNOR U4130 ( .A(n2121), .B(n2120), .Z(c[112]) );
  XNOR U4131 ( .A(n2123), .B(n2122), .Z(c[113]) );
  XNOR U4132 ( .A(n2125), .B(n2124), .Z(c[114]) );
  XNOR U4133 ( .A(n2127), .B(n2126), .Z(c[115]) );
  XNOR U4134 ( .A(n2129), .B(n2128), .Z(c[116]) );
  XNOR U4135 ( .A(n2131), .B(n2130), .Z(c[117]) );
  XNOR U4136 ( .A(n2133), .B(n2132), .Z(c[118]) );
  XNOR U4137 ( .A(n2135), .B(n2134), .Z(c[119]) );
  XNOR U4138 ( .A(n2137), .B(n2136), .Z(c[11]) );
  XNOR U4139 ( .A(n2139), .B(n2138), .Z(c[120]) );
  XNOR U4140 ( .A(n2141), .B(n2140), .Z(c[121]) );
  XNOR U4141 ( .A(n2143), .B(n2142), .Z(c[122]) );
  XNOR U4142 ( .A(n2145), .B(n2144), .Z(c[123]) );
  XNOR U4143 ( .A(n2147), .B(n2146), .Z(c[124]) );
  XNOR U4144 ( .A(n2149), .B(n2148), .Z(c[125]) );
  XNOR U4145 ( .A(n2151), .B(n2150), .Z(c[126]) );
  XNOR U4146 ( .A(n2153), .B(n2152), .Z(c[127]) );
  XNOR U4147 ( .A(n2155), .B(n2154), .Z(c[128]) );
  XNOR U4148 ( .A(n2157), .B(n2156), .Z(c[129]) );
  XNOR U4149 ( .A(n2159), .B(n2158), .Z(c[12]) );
  XNOR U4150 ( .A(n2161), .B(n2160), .Z(c[130]) );
  XNOR U4151 ( .A(n2163), .B(n2162), .Z(c[131]) );
  XNOR U4152 ( .A(n2165), .B(n2164), .Z(c[132]) );
  XNOR U4153 ( .A(n2167), .B(n2166), .Z(c[133]) );
  XNOR U4154 ( .A(n2169), .B(n2168), .Z(c[134]) );
  XNOR U4155 ( .A(n2171), .B(n2170), .Z(c[135]) );
  XNOR U4156 ( .A(n2173), .B(n2172), .Z(c[136]) );
  XNOR U4157 ( .A(n2175), .B(n2174), .Z(c[137]) );
  XNOR U4158 ( .A(n2177), .B(n2176), .Z(c[138]) );
  XNOR U4159 ( .A(n2179), .B(n2178), .Z(c[139]) );
  XNOR U4160 ( .A(n2181), .B(n2180), .Z(c[13]) );
  XNOR U4161 ( .A(n2183), .B(n2182), .Z(c[140]) );
  XNOR U4162 ( .A(n2185), .B(n2184), .Z(c[141]) );
  XNOR U4163 ( .A(n2187), .B(n2186), .Z(c[142]) );
  XNOR U4164 ( .A(n2189), .B(n2188), .Z(c[143]) );
  XNOR U4165 ( .A(n2191), .B(n2190), .Z(c[144]) );
  XNOR U4166 ( .A(n2193), .B(n2192), .Z(c[145]) );
  XNOR U4167 ( .A(n2195), .B(n2194), .Z(c[146]) );
  XNOR U4168 ( .A(n2197), .B(n2196), .Z(c[147]) );
  XNOR U4169 ( .A(n2199), .B(n2198), .Z(c[148]) );
  XNOR U4170 ( .A(n2201), .B(n2200), .Z(c[149]) );
  XNOR U4171 ( .A(n2203), .B(n2202), .Z(c[14]) );
  XNOR U4172 ( .A(n2205), .B(n2204), .Z(c[150]) );
  XNOR U4173 ( .A(n2207), .B(n2206), .Z(c[151]) );
  XNOR U4174 ( .A(n2209), .B(n2208), .Z(c[152]) );
  XNOR U4175 ( .A(n2211), .B(n2210), .Z(c[153]) );
  XNOR U4176 ( .A(n2213), .B(n2212), .Z(c[154]) );
  XNOR U4177 ( .A(n2215), .B(n2214), .Z(c[155]) );
  XNOR U4178 ( .A(n2217), .B(n2216), .Z(c[156]) );
  XNOR U4179 ( .A(n2219), .B(n2218), .Z(c[157]) );
  XNOR U4180 ( .A(n2221), .B(n2220), .Z(c[158]) );
  XNOR U4181 ( .A(n2223), .B(n2222), .Z(c[159]) );
  XNOR U4182 ( .A(n2225), .B(n2224), .Z(c[15]) );
  XNOR U4183 ( .A(n2227), .B(n2226), .Z(c[160]) );
  XNOR U4184 ( .A(n2229), .B(n2228), .Z(c[161]) );
  XNOR U4185 ( .A(n2231), .B(n2230), .Z(c[162]) );
  XNOR U4186 ( .A(n2233), .B(n2232), .Z(c[163]) );
  XNOR U4187 ( .A(n2235), .B(n2234), .Z(c[164]) );
  XNOR U4188 ( .A(n2237), .B(n2236), .Z(c[165]) );
  XNOR U4189 ( .A(n2239), .B(n2238), .Z(c[166]) );
  XNOR U4190 ( .A(n2241), .B(n2240), .Z(c[167]) );
  XNOR U4191 ( .A(n2243), .B(n2242), .Z(c[168]) );
  XNOR U4192 ( .A(n2245), .B(n2244), .Z(c[169]) );
  XNOR U4193 ( .A(n2247), .B(n2246), .Z(c[16]) );
  XNOR U4194 ( .A(n2249), .B(n2248), .Z(c[170]) );
  XNOR U4195 ( .A(n2251), .B(n2250), .Z(c[171]) );
  XNOR U4196 ( .A(n2253), .B(n2252), .Z(c[172]) );
  XNOR U4197 ( .A(n2255), .B(n2254), .Z(c[173]) );
  XNOR U4198 ( .A(n2257), .B(n2256), .Z(c[174]) );
  XNOR U4199 ( .A(n2259), .B(n2258), .Z(c[175]) );
  XNOR U4200 ( .A(n2261), .B(n2260), .Z(c[176]) );
  XNOR U4201 ( .A(n2263), .B(n2262), .Z(c[177]) );
  XNOR U4202 ( .A(n2265), .B(n2264), .Z(c[178]) );
  XNOR U4203 ( .A(n2267), .B(n2266), .Z(c[179]) );
  XNOR U4204 ( .A(n2269), .B(n2268), .Z(c[17]) );
  XNOR U4205 ( .A(n2271), .B(n2270), .Z(c[180]) );
  XNOR U4206 ( .A(n2273), .B(n2272), .Z(c[181]) );
  XNOR U4207 ( .A(n2275), .B(n2274), .Z(c[182]) );
  XNOR U4208 ( .A(n2277), .B(n2276), .Z(c[183]) );
  XNOR U4209 ( .A(n2279), .B(n2278), .Z(c[184]) );
  XNOR U4210 ( .A(n2281), .B(n2280), .Z(c[185]) );
  XNOR U4211 ( .A(n2283), .B(n2282), .Z(c[186]) );
  XNOR U4212 ( .A(n2285), .B(n2284), .Z(c[187]) );
  XNOR U4213 ( .A(n2287), .B(n2286), .Z(c[188]) );
  XNOR U4214 ( .A(n2289), .B(n2288), .Z(c[189]) );
  XNOR U4215 ( .A(n2291), .B(n2290), .Z(c[18]) );
  XNOR U4216 ( .A(n2293), .B(n2292), .Z(c[190]) );
  XNOR U4217 ( .A(n2295), .B(n2294), .Z(c[191]) );
  XNOR U4218 ( .A(n2297), .B(n2296), .Z(c[192]) );
  XNOR U4219 ( .A(n2299), .B(n2298), .Z(c[193]) );
  XNOR U4220 ( .A(n2301), .B(n2300), .Z(c[194]) );
  XNOR U4221 ( .A(n2303), .B(n2302), .Z(c[195]) );
  XNOR U4222 ( .A(n2305), .B(n2304), .Z(c[196]) );
  XNOR U4223 ( .A(n2307), .B(n2306), .Z(c[197]) );
  XNOR U4224 ( .A(n2309), .B(n2308), .Z(c[198]) );
  XNOR U4225 ( .A(n2311), .B(n2310), .Z(c[199]) );
  XNOR U4226 ( .A(n2313), .B(n2312), .Z(c[19]) );
  XNOR U4227 ( .A(n2315), .B(n2314), .Z(c[1]) );
  XNOR U4228 ( .A(n2317), .B(n2316), .Z(c[200]) );
  XNOR U4229 ( .A(n2319), .B(n2318), .Z(c[201]) );
  XNOR U4230 ( .A(n2321), .B(n2320), .Z(c[202]) );
  XNOR U4231 ( .A(n2323), .B(n2322), .Z(c[203]) );
  XNOR U4232 ( .A(n2325), .B(n2324), .Z(c[204]) );
  XNOR U4233 ( .A(n2327), .B(n2326), .Z(c[205]) );
  XNOR U4234 ( .A(n2329), .B(n2328), .Z(c[206]) );
  XNOR U4235 ( .A(n2331), .B(n2330), .Z(c[207]) );
  XNOR U4236 ( .A(n2333), .B(n2332), .Z(c[208]) );
  XNOR U4237 ( .A(n2335), .B(n2334), .Z(c[209]) );
  XNOR U4238 ( .A(n2337), .B(n2336), .Z(c[20]) );
  XNOR U4239 ( .A(n2339), .B(n2338), .Z(c[210]) );
  XNOR U4240 ( .A(n2341), .B(n2340), .Z(c[211]) );
  XNOR U4241 ( .A(n2343), .B(n2342), .Z(c[212]) );
  XNOR U4242 ( .A(n2345), .B(n2344), .Z(c[213]) );
  XNOR U4243 ( .A(n2347), .B(n2346), .Z(c[214]) );
  XNOR U4244 ( .A(n2349), .B(n2348), .Z(c[215]) );
  XNOR U4245 ( .A(n2351), .B(n2350), .Z(c[216]) );
  XNOR U4246 ( .A(n2353), .B(n2352), .Z(c[217]) );
  XNOR U4247 ( .A(n2355), .B(n2354), .Z(c[218]) );
  XNOR U4248 ( .A(n2357), .B(n2356), .Z(c[219]) );
  XNOR U4249 ( .A(n2359), .B(n2358), .Z(c[21]) );
  XNOR U4250 ( .A(n2361), .B(n2360), .Z(c[220]) );
  XNOR U4251 ( .A(n2363), .B(n2362), .Z(c[221]) );
  XNOR U4252 ( .A(n2365), .B(n2364), .Z(c[222]) );
  XNOR U4253 ( .A(n2367), .B(n2366), .Z(c[223]) );
  XNOR U4254 ( .A(n2369), .B(n2368), .Z(c[224]) );
  XNOR U4255 ( .A(n2371), .B(n2370), .Z(c[225]) );
  XNOR U4256 ( .A(n2373), .B(n2372), .Z(c[226]) );
  XNOR U4257 ( .A(n2375), .B(n2374), .Z(c[227]) );
  XNOR U4258 ( .A(n2377), .B(n2376), .Z(c[228]) );
  XNOR U4259 ( .A(n2379), .B(n2378), .Z(c[229]) );
  XNOR U4260 ( .A(n2381), .B(n2380), .Z(c[22]) );
  XNOR U4261 ( .A(n2383), .B(n2382), .Z(c[230]) );
  XNOR U4262 ( .A(n2385), .B(n2384), .Z(c[231]) );
  XNOR U4263 ( .A(n2387), .B(n2386), .Z(c[232]) );
  XNOR U4264 ( .A(n2389), .B(n2388), .Z(c[233]) );
  XNOR U4265 ( .A(n2391), .B(n2390), .Z(c[234]) );
  XNOR U4266 ( .A(n2393), .B(n2392), .Z(c[235]) );
  XNOR U4267 ( .A(n2395), .B(n2394), .Z(c[236]) );
  XNOR U4268 ( .A(n2397), .B(n2396), .Z(c[237]) );
  XNOR U4269 ( .A(n2399), .B(n2398), .Z(c[238]) );
  XNOR U4270 ( .A(n2401), .B(n2400), .Z(c[239]) );
  XNOR U4271 ( .A(n2403), .B(n2402), .Z(c[23]) );
  XNOR U4272 ( .A(n2405), .B(n2404), .Z(c[240]) );
  XNOR U4273 ( .A(n2407), .B(n2406), .Z(c[241]) );
  XNOR U4274 ( .A(n2409), .B(n2408), .Z(c[242]) );
  XNOR U4275 ( .A(n2411), .B(n2410), .Z(c[243]) );
  XNOR U4276 ( .A(n2413), .B(n2412), .Z(c[244]) );
  XNOR U4277 ( .A(n2415), .B(n2414), .Z(c[245]) );
  XNOR U4278 ( .A(n2417), .B(n2416), .Z(c[246]) );
  XNOR U4279 ( .A(n2419), .B(n2418), .Z(c[247]) );
  XNOR U4280 ( .A(n2421), .B(n2420), .Z(c[248]) );
  XNOR U4281 ( .A(n2423), .B(n2422), .Z(c[249]) );
  XNOR U4282 ( .A(n2425), .B(n2424), .Z(c[24]) );
  XNOR U4283 ( .A(n2427), .B(n2426), .Z(c[250]) );
  XNOR U4284 ( .A(n2429), .B(n2428), .Z(c[251]) );
  XNOR U4285 ( .A(n2431), .B(n2430), .Z(c[252]) );
  XNOR U4286 ( .A(n2433), .B(n2432), .Z(c[253]) );
  XNOR U4287 ( .A(n2435), .B(n2434), .Z(c[254]) );
  XNOR U4288 ( .A(n2437), .B(n2436), .Z(c[255]) );
  XNOR U4289 ( .A(n2439), .B(n2438), .Z(c[256]) );
  XNOR U4290 ( .A(n2441), .B(n2440), .Z(c[257]) );
  XNOR U4291 ( .A(n2443), .B(n2442), .Z(c[258]) );
  XNOR U4292 ( .A(n2445), .B(n2444), .Z(c[259]) );
  XNOR U4293 ( .A(n2447), .B(n2446), .Z(c[25]) );
  XNOR U4294 ( .A(n2449), .B(n2448), .Z(c[260]) );
  XNOR U4295 ( .A(n2451), .B(n2450), .Z(c[261]) );
  XNOR U4296 ( .A(n2453), .B(n2452), .Z(c[262]) );
  XNOR U4297 ( .A(n2455), .B(n2454), .Z(c[263]) );
  XNOR U4298 ( .A(n2457), .B(n2456), .Z(c[264]) );
  XNOR U4299 ( .A(n2459), .B(n2458), .Z(c[265]) );
  XNOR U4300 ( .A(n2461), .B(n2460), .Z(c[266]) );
  XNOR U4301 ( .A(n2463), .B(n2462), .Z(c[267]) );
  XNOR U4302 ( .A(n2465), .B(n2464), .Z(c[268]) );
  XNOR U4303 ( .A(n2467), .B(n2466), .Z(c[269]) );
  XNOR U4304 ( .A(n2469), .B(n2468), .Z(c[26]) );
  XNOR U4305 ( .A(n2471), .B(n2470), .Z(c[270]) );
  XNOR U4306 ( .A(n2473), .B(n2472), .Z(c[271]) );
  XNOR U4307 ( .A(n2475), .B(n2474), .Z(c[272]) );
  XNOR U4308 ( .A(n2477), .B(n2476), .Z(c[273]) );
  XNOR U4309 ( .A(n2479), .B(n2478), .Z(c[274]) );
  XNOR U4310 ( .A(n2481), .B(n2480), .Z(c[275]) );
  XNOR U4311 ( .A(n2483), .B(n2482), .Z(c[276]) );
  XNOR U4312 ( .A(n2485), .B(n2484), .Z(c[277]) );
  XNOR U4313 ( .A(n2487), .B(n2486), .Z(c[278]) );
  XNOR U4314 ( .A(n2489), .B(n2488), .Z(c[279]) );
  XNOR U4315 ( .A(n2491), .B(n2490), .Z(c[27]) );
  XNOR U4316 ( .A(n2493), .B(n2492), .Z(c[280]) );
  XNOR U4317 ( .A(n2495), .B(n2494), .Z(c[281]) );
  XNOR U4318 ( .A(n2497), .B(n2496), .Z(c[282]) );
  XNOR U4319 ( .A(n2499), .B(n2498), .Z(c[283]) );
  XNOR U4320 ( .A(n2501), .B(n2500), .Z(c[284]) );
  XNOR U4321 ( .A(n2503), .B(n2502), .Z(c[285]) );
  XNOR U4322 ( .A(n2505), .B(n2504), .Z(c[286]) );
  XNOR U4323 ( .A(n2507), .B(n2506), .Z(c[287]) );
  XNOR U4324 ( .A(n2509), .B(n2508), .Z(c[288]) );
  XNOR U4325 ( .A(n2511), .B(n2510), .Z(c[289]) );
  XNOR U4326 ( .A(n2513), .B(n2512), .Z(c[28]) );
  XNOR U4327 ( .A(n2515), .B(n2514), .Z(c[290]) );
  XNOR U4328 ( .A(n2517), .B(n2516), .Z(c[291]) );
  XNOR U4329 ( .A(n2519), .B(n2518), .Z(c[292]) );
  XNOR U4330 ( .A(n2521), .B(n2520), .Z(c[293]) );
  XNOR U4331 ( .A(n2523), .B(n2522), .Z(c[294]) );
  XNOR U4332 ( .A(n2525), .B(n2524), .Z(c[295]) );
  XNOR U4333 ( .A(n2527), .B(n2526), .Z(c[296]) );
  XNOR U4334 ( .A(n2529), .B(n2528), .Z(c[297]) );
  XNOR U4335 ( .A(n2531), .B(n2530), .Z(c[298]) );
  XNOR U4336 ( .A(n2533), .B(n2532), .Z(c[299]) );
  XNOR U4337 ( .A(n2535), .B(n2534), .Z(c[29]) );
  XNOR U4338 ( .A(n2537), .B(n2536), .Z(c[2]) );
  XNOR U4339 ( .A(n2539), .B(n2538), .Z(c[300]) );
  XNOR U4340 ( .A(n2541), .B(n2540), .Z(c[301]) );
  XNOR U4341 ( .A(n2543), .B(n2542), .Z(c[302]) );
  XNOR U4342 ( .A(n2545), .B(n2544), .Z(c[303]) );
  XNOR U4343 ( .A(n2547), .B(n2546), .Z(c[304]) );
  XNOR U4344 ( .A(n2549), .B(n2548), .Z(c[305]) );
  XNOR U4345 ( .A(n2551), .B(n2550), .Z(c[306]) );
  XNOR U4346 ( .A(n2553), .B(n2552), .Z(c[307]) );
  XNOR U4347 ( .A(n2555), .B(n2554), .Z(c[308]) );
  XNOR U4348 ( .A(n2557), .B(n2556), .Z(c[309]) );
  XNOR U4349 ( .A(n2559), .B(n2558), .Z(c[30]) );
  XNOR U4350 ( .A(n2561), .B(n2560), .Z(c[310]) );
  XNOR U4351 ( .A(n2563), .B(n2562), .Z(c[311]) );
  XNOR U4352 ( .A(n2565), .B(n2564), .Z(c[312]) );
  XNOR U4353 ( .A(n2567), .B(n2566), .Z(c[313]) );
  XNOR U4354 ( .A(n2569), .B(n2568), .Z(c[314]) );
  XNOR U4355 ( .A(n2571), .B(n2570), .Z(c[315]) );
  XNOR U4356 ( .A(n2573), .B(n2572), .Z(c[316]) );
  XNOR U4357 ( .A(n2575), .B(n2574), .Z(c[317]) );
  XNOR U4358 ( .A(n2577), .B(n2576), .Z(c[318]) );
  XNOR U4359 ( .A(n2579), .B(n2578), .Z(c[319]) );
  XNOR U4360 ( .A(n2581), .B(n2580), .Z(c[31]) );
  XNOR U4361 ( .A(n2583), .B(n2582), .Z(c[320]) );
  XNOR U4362 ( .A(n2585), .B(n2584), .Z(c[321]) );
  XNOR U4363 ( .A(n2587), .B(n2586), .Z(c[322]) );
  XNOR U4364 ( .A(n2589), .B(n2588), .Z(c[323]) );
  XNOR U4365 ( .A(n2591), .B(n2590), .Z(c[324]) );
  XNOR U4366 ( .A(n2593), .B(n2592), .Z(c[325]) );
  XNOR U4367 ( .A(n2595), .B(n2594), .Z(c[326]) );
  XNOR U4368 ( .A(n2597), .B(n2596), .Z(c[327]) );
  XNOR U4369 ( .A(n2599), .B(n2598), .Z(c[328]) );
  XNOR U4370 ( .A(n2601), .B(n2600), .Z(c[329]) );
  XNOR U4371 ( .A(n2603), .B(n2602), .Z(c[32]) );
  XNOR U4372 ( .A(n2605), .B(n2604), .Z(c[330]) );
  XNOR U4373 ( .A(n2607), .B(n2606), .Z(c[331]) );
  XNOR U4374 ( .A(n2609), .B(n2608), .Z(c[332]) );
  XNOR U4375 ( .A(n2611), .B(n2610), .Z(c[333]) );
  XNOR U4376 ( .A(n2613), .B(n2612), .Z(c[334]) );
  XNOR U4377 ( .A(n2615), .B(n2614), .Z(c[335]) );
  XNOR U4378 ( .A(n2617), .B(n2616), .Z(c[336]) );
  XNOR U4379 ( .A(n2619), .B(n2618), .Z(c[337]) );
  XNOR U4380 ( .A(n2621), .B(n2620), .Z(c[338]) );
  XNOR U4381 ( .A(n2623), .B(n2622), .Z(c[339]) );
  XNOR U4382 ( .A(n2625), .B(n2624), .Z(c[33]) );
  XNOR U4383 ( .A(n2627), .B(n2626), .Z(c[340]) );
  XNOR U4384 ( .A(n2629), .B(n2628), .Z(c[341]) );
  XNOR U4385 ( .A(n2631), .B(n2630), .Z(c[342]) );
  XNOR U4386 ( .A(n2633), .B(n2632), .Z(c[343]) );
  XNOR U4387 ( .A(n2635), .B(n2634), .Z(c[344]) );
  XNOR U4388 ( .A(n2637), .B(n2636), .Z(c[345]) );
  XNOR U4389 ( .A(n2639), .B(n2638), .Z(c[346]) );
  XNOR U4390 ( .A(n2641), .B(n2640), .Z(c[347]) );
  XNOR U4391 ( .A(n2643), .B(n2642), .Z(c[348]) );
  XNOR U4392 ( .A(n2645), .B(n2644), .Z(c[349]) );
  XNOR U4393 ( .A(n2647), .B(n2646), .Z(c[34]) );
  XNOR U4394 ( .A(n2649), .B(n2648), .Z(c[350]) );
  XNOR U4395 ( .A(n2651), .B(n2650), .Z(c[351]) );
  XNOR U4396 ( .A(n2653), .B(n2652), .Z(c[352]) );
  XNOR U4397 ( .A(n2655), .B(n2654), .Z(c[353]) );
  XNOR U4398 ( .A(n2657), .B(n2656), .Z(c[354]) );
  XNOR U4399 ( .A(n2659), .B(n2658), .Z(c[355]) );
  XNOR U4400 ( .A(n2661), .B(n2660), .Z(c[356]) );
  XNOR U4401 ( .A(n2663), .B(n2662), .Z(c[357]) );
  XNOR U4402 ( .A(n2665), .B(n2664), .Z(c[358]) );
  XNOR U4403 ( .A(n2667), .B(n2666), .Z(c[359]) );
  XNOR U4404 ( .A(n2669), .B(n2668), .Z(c[35]) );
  XNOR U4405 ( .A(n2671), .B(n2670), .Z(c[360]) );
  XNOR U4406 ( .A(n2673), .B(n2672), .Z(c[361]) );
  XNOR U4407 ( .A(n2675), .B(n2674), .Z(c[362]) );
  XNOR U4408 ( .A(n2677), .B(n2676), .Z(c[363]) );
  XNOR U4409 ( .A(n2679), .B(n2678), .Z(c[364]) );
  XNOR U4410 ( .A(n2681), .B(n2680), .Z(c[365]) );
  XNOR U4411 ( .A(n2683), .B(n2682), .Z(c[366]) );
  XNOR U4412 ( .A(n2685), .B(n2684), .Z(c[367]) );
  XNOR U4413 ( .A(n2687), .B(n2686), .Z(c[368]) );
  XNOR U4414 ( .A(n2689), .B(n2688), .Z(c[369]) );
  XNOR U4415 ( .A(n2691), .B(n2690), .Z(c[36]) );
  XNOR U4416 ( .A(n2693), .B(n2692), .Z(c[370]) );
  XNOR U4417 ( .A(n2695), .B(n2694), .Z(c[371]) );
  XNOR U4418 ( .A(n2697), .B(n2696), .Z(c[372]) );
  XNOR U4419 ( .A(n2699), .B(n2698), .Z(c[373]) );
  XNOR U4420 ( .A(n2701), .B(n2700), .Z(c[374]) );
  XNOR U4421 ( .A(n2703), .B(n2702), .Z(c[375]) );
  XNOR U4422 ( .A(n2705), .B(n2704), .Z(c[376]) );
  XNOR U4423 ( .A(n2707), .B(n2706), .Z(c[377]) );
  XNOR U4424 ( .A(n2709), .B(n2708), .Z(c[378]) );
  XNOR U4425 ( .A(n2711), .B(n2710), .Z(c[379]) );
  XNOR U4426 ( .A(n2713), .B(n2712), .Z(c[37]) );
  XNOR U4427 ( .A(n2715), .B(n2714), .Z(c[380]) );
  XNOR U4428 ( .A(n2717), .B(n2716), .Z(c[381]) );
  XNOR U4429 ( .A(n2719), .B(n2718), .Z(c[382]) );
  XNOR U4430 ( .A(n2721), .B(n2720), .Z(c[383]) );
  XNOR U4431 ( .A(n2723), .B(n2722), .Z(c[384]) );
  XNOR U4432 ( .A(n2725), .B(n2724), .Z(c[385]) );
  XNOR U4433 ( .A(n2727), .B(n2726), .Z(c[386]) );
  XNOR U4434 ( .A(n2729), .B(n2728), .Z(c[387]) );
  XNOR U4435 ( .A(n2731), .B(n2730), .Z(c[388]) );
  XNOR U4436 ( .A(n2733), .B(n2732), .Z(c[389]) );
  XNOR U4437 ( .A(n2735), .B(n2734), .Z(c[38]) );
  XNOR U4438 ( .A(n2737), .B(n2736), .Z(c[390]) );
  XNOR U4439 ( .A(n2739), .B(n2738), .Z(c[391]) );
  XNOR U4440 ( .A(n2741), .B(n2740), .Z(c[392]) );
  XNOR U4441 ( .A(n2743), .B(n2742), .Z(c[393]) );
  XNOR U4442 ( .A(n2745), .B(n2744), .Z(c[394]) );
  XNOR U4443 ( .A(n2747), .B(n2746), .Z(c[395]) );
  XNOR U4444 ( .A(n2749), .B(n2748), .Z(c[396]) );
  XNOR U4445 ( .A(n2751), .B(n2750), .Z(c[397]) );
  XNOR U4446 ( .A(n2753), .B(n2752), .Z(c[398]) );
  XNOR U4447 ( .A(n2755), .B(n2754), .Z(c[399]) );
  XNOR U4448 ( .A(n2757), .B(n2756), .Z(c[39]) );
  XNOR U4449 ( .A(n2759), .B(n2758), .Z(c[3]) );
  XNOR U4450 ( .A(n2761), .B(n2760), .Z(c[400]) );
  XNOR U4451 ( .A(n2763), .B(n2762), .Z(c[401]) );
  XNOR U4452 ( .A(n2765), .B(n2764), .Z(c[402]) );
  XNOR U4453 ( .A(n2767), .B(n2766), .Z(c[403]) );
  XNOR U4454 ( .A(n2769), .B(n2768), .Z(c[404]) );
  XNOR U4455 ( .A(n2771), .B(n2770), .Z(c[405]) );
  XNOR U4456 ( .A(n2773), .B(n2772), .Z(c[406]) );
  XNOR U4457 ( .A(n2775), .B(n2774), .Z(c[407]) );
  XNOR U4458 ( .A(n2777), .B(n2776), .Z(c[408]) );
  XNOR U4459 ( .A(n2779), .B(n2778), .Z(c[409]) );
  XNOR U4460 ( .A(n2781), .B(n2780), .Z(c[40]) );
  XNOR U4461 ( .A(n2783), .B(n2782), .Z(c[410]) );
  XNOR U4462 ( .A(n2785), .B(n2784), .Z(c[411]) );
  XNOR U4463 ( .A(n2787), .B(n2786), .Z(c[412]) );
  XNOR U4464 ( .A(n2789), .B(n2788), .Z(c[413]) );
  XNOR U4465 ( .A(n2791), .B(n2790), .Z(c[414]) );
  XNOR U4466 ( .A(n2793), .B(n2792), .Z(c[415]) );
  XNOR U4467 ( .A(n2795), .B(n2794), .Z(c[416]) );
  XNOR U4468 ( .A(n2797), .B(n2796), .Z(c[417]) );
  XNOR U4469 ( .A(n2799), .B(n2798), .Z(c[418]) );
  XNOR U4470 ( .A(n2801), .B(n2800), .Z(c[419]) );
  XNOR U4471 ( .A(n2803), .B(n2802), .Z(c[41]) );
  XNOR U4472 ( .A(n2805), .B(n2804), .Z(c[420]) );
  XNOR U4473 ( .A(n2807), .B(n2806), .Z(c[421]) );
  XNOR U4474 ( .A(n2809), .B(n2808), .Z(c[422]) );
  XNOR U4475 ( .A(n2811), .B(n2810), .Z(c[423]) );
  XNOR U4476 ( .A(n2813), .B(n2812), .Z(c[424]) );
  XNOR U4477 ( .A(n2815), .B(n2814), .Z(c[425]) );
  XNOR U4478 ( .A(n2817), .B(n2816), .Z(c[426]) );
  XNOR U4479 ( .A(n2819), .B(n2818), .Z(c[427]) );
  XNOR U4480 ( .A(n2821), .B(n2820), .Z(c[428]) );
  XNOR U4481 ( .A(n2823), .B(n2822), .Z(c[429]) );
  XNOR U4482 ( .A(n2825), .B(n2824), .Z(c[42]) );
  XNOR U4483 ( .A(n2827), .B(n2826), .Z(c[430]) );
  XNOR U4484 ( .A(n2829), .B(n2828), .Z(c[431]) );
  XNOR U4485 ( .A(n2831), .B(n2830), .Z(c[432]) );
  XNOR U4486 ( .A(n2833), .B(n2832), .Z(c[433]) );
  XNOR U4487 ( .A(n2835), .B(n2834), .Z(c[434]) );
  XNOR U4488 ( .A(n2837), .B(n2836), .Z(c[435]) );
  XNOR U4489 ( .A(n2839), .B(n2838), .Z(c[436]) );
  XNOR U4490 ( .A(n2841), .B(n2840), .Z(c[437]) );
  XNOR U4491 ( .A(n2843), .B(n2842), .Z(c[438]) );
  XNOR U4492 ( .A(n2845), .B(n2844), .Z(c[439]) );
  XNOR U4493 ( .A(n2847), .B(n2846), .Z(c[43]) );
  XNOR U4494 ( .A(n2849), .B(n2848), .Z(c[440]) );
  XNOR U4495 ( .A(n2851), .B(n2850), .Z(c[441]) );
  XNOR U4496 ( .A(n2853), .B(n2852), .Z(c[442]) );
  XNOR U4497 ( .A(n2855), .B(n2854), .Z(c[443]) );
  XNOR U4498 ( .A(n2857), .B(n2856), .Z(c[444]) );
  XNOR U4499 ( .A(n2859), .B(n2858), .Z(c[445]) );
  XNOR U4500 ( .A(n2861), .B(n2860), .Z(c[446]) );
  XNOR U4501 ( .A(n2863), .B(n2862), .Z(c[447]) );
  XNOR U4502 ( .A(n2865), .B(n2864), .Z(c[448]) );
  XNOR U4503 ( .A(n2867), .B(n2866), .Z(c[449]) );
  XNOR U4504 ( .A(n2869), .B(n2868), .Z(c[44]) );
  XNOR U4505 ( .A(n2871), .B(n2870), .Z(c[450]) );
  XNOR U4506 ( .A(n2873), .B(n2872), .Z(c[451]) );
  XNOR U4507 ( .A(n2875), .B(n2874), .Z(c[452]) );
  XNOR U4508 ( .A(n2877), .B(n2876), .Z(c[453]) );
  XNOR U4509 ( .A(n2879), .B(n2878), .Z(c[454]) );
  XNOR U4510 ( .A(n2881), .B(n2880), .Z(c[455]) );
  XNOR U4511 ( .A(n2883), .B(n2882), .Z(c[456]) );
  XNOR U4512 ( .A(n2885), .B(n2884), .Z(c[457]) );
  XNOR U4513 ( .A(n2887), .B(n2886), .Z(c[458]) );
  XNOR U4514 ( .A(n2889), .B(n2888), .Z(c[459]) );
  XNOR U4515 ( .A(n2891), .B(n2890), .Z(c[45]) );
  XNOR U4516 ( .A(n2893), .B(n2892), .Z(c[460]) );
  XNOR U4517 ( .A(n2895), .B(n2894), .Z(c[461]) );
  XNOR U4518 ( .A(n2897), .B(n2896), .Z(c[462]) );
  XNOR U4519 ( .A(n2899), .B(n2898), .Z(c[463]) );
  XNOR U4520 ( .A(n2901), .B(n2900), .Z(c[464]) );
  XNOR U4521 ( .A(n2903), .B(n2902), .Z(c[465]) );
  XNOR U4522 ( .A(n2905), .B(n2904), .Z(c[466]) );
  XNOR U4523 ( .A(n2907), .B(n2906), .Z(c[467]) );
  XNOR U4524 ( .A(n2909), .B(n2908), .Z(c[468]) );
  XNOR U4525 ( .A(n2911), .B(n2910), .Z(c[469]) );
  XNOR U4526 ( .A(n2913), .B(n2912), .Z(c[46]) );
  XNOR U4527 ( .A(n2915), .B(n2914), .Z(c[470]) );
  XNOR U4528 ( .A(n2917), .B(n2916), .Z(c[471]) );
  XNOR U4529 ( .A(n2919), .B(n2918), .Z(c[472]) );
  XNOR U4530 ( .A(n2921), .B(n2920), .Z(c[473]) );
  XNOR U4531 ( .A(n2923), .B(n2922), .Z(c[474]) );
  XNOR U4532 ( .A(n2925), .B(n2924), .Z(c[475]) );
  XNOR U4533 ( .A(n2927), .B(n2926), .Z(c[476]) );
  XNOR U4534 ( .A(n2929), .B(n2928), .Z(c[477]) );
  XNOR U4535 ( .A(n2931), .B(n2930), .Z(c[478]) );
  XNOR U4536 ( .A(n2933), .B(n2932), .Z(c[479]) );
  XNOR U4537 ( .A(n2935), .B(n2934), .Z(c[47]) );
  XNOR U4538 ( .A(n2937), .B(n2936), .Z(c[480]) );
  XNOR U4539 ( .A(n2939), .B(n2938), .Z(c[481]) );
  XNOR U4540 ( .A(n2941), .B(n2940), .Z(c[482]) );
  XNOR U4541 ( .A(n2943), .B(n2942), .Z(c[483]) );
  XNOR U4542 ( .A(n2945), .B(n2944), .Z(c[484]) );
  XNOR U4543 ( .A(n2947), .B(n2946), .Z(c[485]) );
  XNOR U4544 ( .A(n2949), .B(n2948), .Z(c[486]) );
  XNOR U4545 ( .A(n2951), .B(n2950), .Z(c[487]) );
  XNOR U4546 ( .A(n2953), .B(n2952), .Z(c[488]) );
  XNOR U4547 ( .A(n2955), .B(n2954), .Z(c[489]) );
  XNOR U4548 ( .A(n2957), .B(n2956), .Z(c[48]) );
  XNOR U4549 ( .A(n2959), .B(n2958), .Z(c[490]) );
  XNOR U4550 ( .A(n2961), .B(n2960), .Z(c[491]) );
  XNOR U4551 ( .A(n2963), .B(n2962), .Z(c[492]) );
  XNOR U4552 ( .A(n2965), .B(n2964), .Z(c[493]) );
  XNOR U4553 ( .A(n2967), .B(n2966), .Z(c[494]) );
  XNOR U4554 ( .A(n2969), .B(n2968), .Z(c[495]) );
  XNOR U4555 ( .A(n2971), .B(n2970), .Z(c[496]) );
  XNOR U4556 ( .A(n2973), .B(n2972), .Z(c[497]) );
  XNOR U4557 ( .A(n2975), .B(n2974), .Z(c[498]) );
  XNOR U4558 ( .A(n2977), .B(n2976), .Z(c[499]) );
  XNOR U4559 ( .A(n2979), .B(n2978), .Z(c[49]) );
  XNOR U4560 ( .A(n2981), .B(n2980), .Z(c[4]) );
  XNOR U4561 ( .A(n2983), .B(n2982), .Z(c[500]) );
  XNOR U4562 ( .A(n2985), .B(n2984), .Z(c[501]) );
  XNOR U4563 ( .A(n2987), .B(n2986), .Z(c[502]) );
  XNOR U4564 ( .A(n2989), .B(n2988), .Z(c[503]) );
  XNOR U4565 ( .A(n2991), .B(n2990), .Z(c[504]) );
  XNOR U4566 ( .A(n2993), .B(n2992), .Z(c[505]) );
  XNOR U4567 ( .A(n2995), .B(n2994), .Z(c[506]) );
  XNOR U4568 ( .A(n2997), .B(n2996), .Z(c[507]) );
  XNOR U4569 ( .A(n2999), .B(n2998), .Z(c[508]) );
  XNOR U4570 ( .A(n3001), .B(n3000), .Z(c[509]) );
  XNOR U4571 ( .A(n3003), .B(n3002), .Z(c[50]) );
  XNOR U4572 ( .A(n3005), .B(n3004), .Z(c[510]) );
  XNOR U4573 ( .A(n3007), .B(n3006), .Z(c[511]) );
  XNOR U4574 ( .A(n3009), .B(n3008), .Z(c[512]) );
  XNOR U4575 ( .A(n3011), .B(n3010), .Z(c[513]) );
  XNOR U4576 ( .A(n3013), .B(n3012), .Z(c[514]) );
  XNOR U4577 ( .A(n3015), .B(n3014), .Z(c[515]) );
  XNOR U4578 ( .A(n3017), .B(n3016), .Z(c[516]) );
  XNOR U4579 ( .A(n3019), .B(n3018), .Z(c[517]) );
  XNOR U4580 ( .A(n3021), .B(n3020), .Z(c[518]) );
  XNOR U4581 ( .A(n3023), .B(n3022), .Z(c[519]) );
  XNOR U4582 ( .A(n3025), .B(n3024), .Z(c[51]) );
  XNOR U4583 ( .A(n3027), .B(n3026), .Z(c[520]) );
  XNOR U4584 ( .A(n3029), .B(n3028), .Z(c[521]) );
  XNOR U4585 ( .A(n3031), .B(n3030), .Z(c[522]) );
  XNOR U4586 ( .A(n3033), .B(n3032), .Z(c[523]) );
  XNOR U4587 ( .A(n3035), .B(n3034), .Z(c[524]) );
  XNOR U4588 ( .A(n3037), .B(n3036), .Z(c[525]) );
  XNOR U4589 ( .A(n3039), .B(n3038), .Z(c[526]) );
  XNOR U4590 ( .A(n3041), .B(n3040), .Z(c[527]) );
  XNOR U4591 ( .A(n3043), .B(n3042), .Z(c[528]) );
  XNOR U4592 ( .A(n3045), .B(n3044), .Z(c[529]) );
  XNOR U4593 ( .A(n3047), .B(n3046), .Z(c[52]) );
  XNOR U4594 ( .A(n3049), .B(n3048), .Z(c[530]) );
  XNOR U4595 ( .A(n3051), .B(n3050), .Z(c[531]) );
  XNOR U4596 ( .A(n3053), .B(n3052), .Z(c[532]) );
  XNOR U4597 ( .A(n3055), .B(n3054), .Z(c[533]) );
  XNOR U4598 ( .A(n3057), .B(n3056), .Z(c[534]) );
  XNOR U4599 ( .A(n3059), .B(n3058), .Z(c[535]) );
  XNOR U4600 ( .A(n3061), .B(n3060), .Z(c[536]) );
  XNOR U4601 ( .A(n3063), .B(n3062), .Z(c[537]) );
  XNOR U4602 ( .A(n3065), .B(n3064), .Z(c[538]) );
  XNOR U4603 ( .A(n3067), .B(n3066), .Z(c[539]) );
  XNOR U4604 ( .A(n3069), .B(n3068), .Z(c[53]) );
  XNOR U4605 ( .A(n3071), .B(n3070), .Z(c[540]) );
  XNOR U4606 ( .A(n3073), .B(n3072), .Z(c[541]) );
  XNOR U4607 ( .A(n3075), .B(n3074), .Z(c[542]) );
  XNOR U4608 ( .A(n3077), .B(n3076), .Z(c[543]) );
  XNOR U4609 ( .A(n3079), .B(n3078), .Z(c[544]) );
  XNOR U4610 ( .A(n3081), .B(n3080), .Z(c[545]) );
  XNOR U4611 ( .A(n3083), .B(n3082), .Z(c[546]) );
  XNOR U4612 ( .A(n3085), .B(n3084), .Z(c[547]) );
  XNOR U4613 ( .A(n3087), .B(n3086), .Z(c[548]) );
  XNOR U4614 ( .A(n3089), .B(n3088), .Z(c[549]) );
  XNOR U4615 ( .A(n3091), .B(n3090), .Z(c[54]) );
  XNOR U4616 ( .A(n3093), .B(n3092), .Z(c[550]) );
  XNOR U4617 ( .A(n3095), .B(n3094), .Z(c[551]) );
  XNOR U4618 ( .A(n3097), .B(n3096), .Z(c[552]) );
  XNOR U4619 ( .A(n3099), .B(n3098), .Z(c[553]) );
  XNOR U4620 ( .A(n3101), .B(n3100), .Z(c[554]) );
  XNOR U4621 ( .A(n3103), .B(n3102), .Z(c[555]) );
  XNOR U4622 ( .A(n3105), .B(n3104), .Z(c[556]) );
  XNOR U4623 ( .A(n3107), .B(n3106), .Z(c[557]) );
  XNOR U4624 ( .A(n3109), .B(n3108), .Z(c[558]) );
  XNOR U4625 ( .A(n3111), .B(n3110), .Z(c[559]) );
  XNOR U4626 ( .A(n3113), .B(n3112), .Z(c[55]) );
  XNOR U4627 ( .A(n3115), .B(n3114), .Z(c[560]) );
  XNOR U4628 ( .A(n3117), .B(n3116), .Z(c[561]) );
  XNOR U4629 ( .A(n3119), .B(n3118), .Z(c[562]) );
  XNOR U4630 ( .A(n3121), .B(n3120), .Z(c[563]) );
  XNOR U4631 ( .A(n3123), .B(n3122), .Z(c[564]) );
  XNOR U4632 ( .A(n3125), .B(n3124), .Z(c[565]) );
  XNOR U4633 ( .A(n3127), .B(n3126), .Z(c[566]) );
  XNOR U4634 ( .A(n3129), .B(n3128), .Z(c[567]) );
  XNOR U4635 ( .A(n3131), .B(n3130), .Z(c[568]) );
  XNOR U4636 ( .A(n3133), .B(n3132), .Z(c[569]) );
  XNOR U4637 ( .A(n3135), .B(n3134), .Z(c[56]) );
  XNOR U4638 ( .A(n3137), .B(n3136), .Z(c[570]) );
  XNOR U4639 ( .A(n3139), .B(n3138), .Z(c[571]) );
  XNOR U4640 ( .A(n3141), .B(n3140), .Z(c[572]) );
  XNOR U4641 ( .A(n3143), .B(n3142), .Z(c[573]) );
  XNOR U4642 ( .A(n3145), .B(n3144), .Z(c[574]) );
  XNOR U4643 ( .A(n3147), .B(n3146), .Z(c[575]) );
  XNOR U4644 ( .A(n3149), .B(n3148), .Z(c[576]) );
  XNOR U4645 ( .A(n3151), .B(n3150), .Z(c[577]) );
  XNOR U4646 ( .A(n3153), .B(n3152), .Z(c[578]) );
  XNOR U4647 ( .A(n3155), .B(n3154), .Z(c[579]) );
  XNOR U4648 ( .A(n3157), .B(n3156), .Z(c[57]) );
  XNOR U4649 ( .A(n3159), .B(n3158), .Z(c[580]) );
  XNOR U4650 ( .A(n3161), .B(n3160), .Z(c[581]) );
  XNOR U4651 ( .A(n3163), .B(n3162), .Z(c[582]) );
  XNOR U4652 ( .A(n3165), .B(n3164), .Z(c[583]) );
  XNOR U4653 ( .A(n3167), .B(n3166), .Z(c[584]) );
  XNOR U4654 ( .A(n3169), .B(n3168), .Z(c[585]) );
  XNOR U4655 ( .A(n3171), .B(n3170), .Z(c[586]) );
  XNOR U4656 ( .A(n3173), .B(n3172), .Z(c[587]) );
  XNOR U4657 ( .A(n3175), .B(n3174), .Z(c[588]) );
  XNOR U4658 ( .A(n3177), .B(n3176), .Z(c[589]) );
  XNOR U4659 ( .A(n3179), .B(n3178), .Z(c[58]) );
  XNOR U4660 ( .A(n3181), .B(n3180), .Z(c[590]) );
  XNOR U4661 ( .A(n3183), .B(n3182), .Z(c[591]) );
  XNOR U4662 ( .A(n3185), .B(n3184), .Z(c[592]) );
  XNOR U4663 ( .A(n3187), .B(n3186), .Z(c[593]) );
  XNOR U4664 ( .A(n3189), .B(n3188), .Z(c[594]) );
  XNOR U4665 ( .A(n3191), .B(n3190), .Z(c[595]) );
  XNOR U4666 ( .A(n3193), .B(n3192), .Z(c[596]) );
  XNOR U4667 ( .A(n3195), .B(n3194), .Z(c[597]) );
  XNOR U4668 ( .A(n3197), .B(n3196), .Z(c[598]) );
  XNOR U4669 ( .A(n3199), .B(n3198), .Z(c[599]) );
  XNOR U4670 ( .A(n3201), .B(n3200), .Z(c[59]) );
  XNOR U4671 ( .A(n3203), .B(n3202), .Z(c[5]) );
  XNOR U4672 ( .A(n3205), .B(n3204), .Z(c[600]) );
  XNOR U4673 ( .A(n3207), .B(n3206), .Z(c[601]) );
  XNOR U4674 ( .A(n3209), .B(n3208), .Z(c[602]) );
  XNOR U4675 ( .A(n3211), .B(n3210), .Z(c[603]) );
  XNOR U4676 ( .A(n3213), .B(n3212), .Z(c[604]) );
  XNOR U4677 ( .A(n3215), .B(n3214), .Z(c[605]) );
  XNOR U4678 ( .A(n3217), .B(n3216), .Z(c[606]) );
  XNOR U4679 ( .A(n3219), .B(n3218), .Z(c[607]) );
  XNOR U4680 ( .A(n3221), .B(n3220), .Z(c[608]) );
  XNOR U4681 ( .A(n3223), .B(n3222), .Z(c[609]) );
  XNOR U4682 ( .A(n3225), .B(n3224), .Z(c[60]) );
  XNOR U4683 ( .A(n3227), .B(n3226), .Z(c[610]) );
  XNOR U4684 ( .A(n3229), .B(n3228), .Z(c[611]) );
  XNOR U4685 ( .A(n3231), .B(n3230), .Z(c[612]) );
  XNOR U4686 ( .A(n3233), .B(n3232), .Z(c[613]) );
  XNOR U4687 ( .A(n3235), .B(n3234), .Z(c[614]) );
  XNOR U4688 ( .A(n3237), .B(n3236), .Z(c[615]) );
  XNOR U4689 ( .A(n3239), .B(n3238), .Z(c[616]) );
  XNOR U4690 ( .A(n3241), .B(n3240), .Z(c[617]) );
  XNOR U4691 ( .A(n3243), .B(n3242), .Z(c[618]) );
  XNOR U4692 ( .A(n3245), .B(n3244), .Z(c[619]) );
  XNOR U4693 ( .A(n3247), .B(n3246), .Z(c[61]) );
  XNOR U4694 ( .A(n3249), .B(n3248), .Z(c[620]) );
  XNOR U4695 ( .A(n3251), .B(n3250), .Z(c[621]) );
  XNOR U4696 ( .A(n3253), .B(n3252), .Z(c[622]) );
  XNOR U4697 ( .A(n3255), .B(n3254), .Z(c[623]) );
  XNOR U4698 ( .A(n3257), .B(n3256), .Z(c[624]) );
  XNOR U4699 ( .A(n3259), .B(n3258), .Z(c[625]) );
  XNOR U4700 ( .A(n3261), .B(n3260), .Z(c[626]) );
  XNOR U4701 ( .A(n3263), .B(n3262), .Z(c[627]) );
  XNOR U4702 ( .A(n3265), .B(n3264), .Z(c[628]) );
  XNOR U4703 ( .A(n3267), .B(n3266), .Z(c[629]) );
  XNOR U4704 ( .A(n3269), .B(n3268), .Z(c[62]) );
  XNOR U4705 ( .A(n3271), .B(n3270), .Z(c[630]) );
  XNOR U4706 ( .A(n3273), .B(n3272), .Z(c[631]) );
  XNOR U4707 ( .A(n3275), .B(n3274), .Z(c[632]) );
  XNOR U4708 ( .A(n3277), .B(n3276), .Z(c[633]) );
  XNOR U4709 ( .A(n3279), .B(n3278), .Z(c[634]) );
  XNOR U4710 ( .A(n3281), .B(n3280), .Z(c[635]) );
  XNOR U4711 ( .A(n3283), .B(n3282), .Z(c[636]) );
  XNOR U4712 ( .A(n3285), .B(n3284), .Z(c[637]) );
  XNOR U4713 ( .A(n3287), .B(n3286), .Z(c[638]) );
  XNOR U4714 ( .A(n3289), .B(n3288), .Z(c[639]) );
  XNOR U4715 ( .A(n3291), .B(n3290), .Z(c[63]) );
  XNOR U4716 ( .A(n3293), .B(n3292), .Z(c[640]) );
  XNOR U4717 ( .A(n3295), .B(n3294), .Z(c[641]) );
  XNOR U4718 ( .A(n3297), .B(n3296), .Z(c[642]) );
  XNOR U4719 ( .A(n3299), .B(n3298), .Z(c[643]) );
  XNOR U4720 ( .A(n3301), .B(n3300), .Z(c[644]) );
  XNOR U4721 ( .A(n3303), .B(n3302), .Z(c[645]) );
  XNOR U4722 ( .A(n3305), .B(n3304), .Z(c[646]) );
  XNOR U4723 ( .A(n3307), .B(n3306), .Z(c[647]) );
  XNOR U4724 ( .A(n3309), .B(n3308), .Z(c[648]) );
  XNOR U4725 ( .A(n3311), .B(n3310), .Z(c[649]) );
  XNOR U4726 ( .A(n3313), .B(n3312), .Z(c[64]) );
  XNOR U4727 ( .A(n3315), .B(n3314), .Z(c[650]) );
  XNOR U4728 ( .A(n3317), .B(n3316), .Z(c[651]) );
  XNOR U4729 ( .A(n3319), .B(n3318), .Z(c[652]) );
  XNOR U4730 ( .A(n3321), .B(n3320), .Z(c[653]) );
  XNOR U4731 ( .A(n3323), .B(n3322), .Z(c[654]) );
  XNOR U4732 ( .A(n3325), .B(n3324), .Z(c[655]) );
  XNOR U4733 ( .A(n3327), .B(n3326), .Z(c[656]) );
  XNOR U4734 ( .A(n3329), .B(n3328), .Z(c[657]) );
  XNOR U4735 ( .A(n3331), .B(n3330), .Z(c[658]) );
  XNOR U4736 ( .A(n3333), .B(n3332), .Z(c[659]) );
  XNOR U4737 ( .A(n3335), .B(n3334), .Z(c[65]) );
  XNOR U4738 ( .A(n3337), .B(n3336), .Z(c[660]) );
  XNOR U4739 ( .A(n3339), .B(n3338), .Z(c[661]) );
  XNOR U4740 ( .A(n3341), .B(n3340), .Z(c[662]) );
  XNOR U4741 ( .A(n3343), .B(n3342), .Z(c[663]) );
  XNOR U4742 ( .A(n3345), .B(n3344), .Z(c[664]) );
  XNOR U4743 ( .A(n3347), .B(n3346), .Z(c[665]) );
  XNOR U4744 ( .A(n3349), .B(n3348), .Z(c[666]) );
  XNOR U4745 ( .A(n3351), .B(n3350), .Z(c[667]) );
  XNOR U4746 ( .A(n3353), .B(n3352), .Z(c[668]) );
  XNOR U4747 ( .A(n3355), .B(n3354), .Z(c[669]) );
  XNOR U4748 ( .A(n3357), .B(n3356), .Z(c[66]) );
  XNOR U4749 ( .A(n3359), .B(n3358), .Z(c[670]) );
  XNOR U4750 ( .A(n3361), .B(n3360), .Z(c[671]) );
  XNOR U4751 ( .A(n3363), .B(n3362), .Z(c[672]) );
  XNOR U4752 ( .A(n3365), .B(n3364), .Z(c[673]) );
  XNOR U4753 ( .A(n3367), .B(n3366), .Z(c[674]) );
  XNOR U4754 ( .A(n3369), .B(n3368), .Z(c[675]) );
  XNOR U4755 ( .A(n3371), .B(n3370), .Z(c[676]) );
  XNOR U4756 ( .A(n3373), .B(n3372), .Z(c[677]) );
  XNOR U4757 ( .A(n3375), .B(n3374), .Z(c[678]) );
  XNOR U4758 ( .A(n3377), .B(n3376), .Z(c[679]) );
  XNOR U4759 ( .A(n3379), .B(n3378), .Z(c[67]) );
  XNOR U4760 ( .A(n3381), .B(n3380), .Z(c[680]) );
  XNOR U4761 ( .A(n3383), .B(n3382), .Z(c[681]) );
  XNOR U4762 ( .A(n3385), .B(n3384), .Z(c[682]) );
  XNOR U4763 ( .A(n3387), .B(n3386), .Z(c[683]) );
  XNOR U4764 ( .A(n3389), .B(n3388), .Z(c[684]) );
  XNOR U4765 ( .A(n3391), .B(n3390), .Z(c[685]) );
  XNOR U4766 ( .A(n3393), .B(n3392), .Z(c[686]) );
  XNOR U4767 ( .A(n3395), .B(n3394), .Z(c[687]) );
  XNOR U4768 ( .A(n3397), .B(n3396), .Z(c[688]) );
  XNOR U4769 ( .A(n3399), .B(n3398), .Z(c[689]) );
  XNOR U4770 ( .A(n3401), .B(n3400), .Z(c[68]) );
  XNOR U4771 ( .A(n3403), .B(n3402), .Z(c[690]) );
  XNOR U4772 ( .A(n3405), .B(n3404), .Z(c[691]) );
  XNOR U4773 ( .A(n3407), .B(n3406), .Z(c[692]) );
  XNOR U4774 ( .A(n3409), .B(n3408), .Z(c[693]) );
  XNOR U4775 ( .A(n3411), .B(n3410), .Z(c[694]) );
  XNOR U4776 ( .A(n3413), .B(n3412), .Z(c[695]) );
  XNOR U4777 ( .A(n3415), .B(n3414), .Z(c[696]) );
  XNOR U4778 ( .A(n3417), .B(n3416), .Z(c[697]) );
  XNOR U4779 ( .A(n3419), .B(n3418), .Z(c[698]) );
  XNOR U4780 ( .A(n3421), .B(n3420), .Z(c[699]) );
  XNOR U4781 ( .A(n3423), .B(n3422), .Z(c[69]) );
  XNOR U4782 ( .A(n3425), .B(n3424), .Z(c[6]) );
  XNOR U4783 ( .A(n3427), .B(n3426), .Z(c[700]) );
  XNOR U4784 ( .A(n3429), .B(n3428), .Z(c[701]) );
  XNOR U4785 ( .A(n3431), .B(n3430), .Z(c[702]) );
  XNOR U4786 ( .A(n3433), .B(n3432), .Z(c[703]) );
  XNOR U4787 ( .A(n3435), .B(n3434), .Z(c[704]) );
  XNOR U4788 ( .A(n3437), .B(n3436), .Z(c[705]) );
  XNOR U4789 ( .A(n3439), .B(n3438), .Z(c[706]) );
  XNOR U4790 ( .A(n3441), .B(n3440), .Z(c[707]) );
  XNOR U4791 ( .A(n3443), .B(n3442), .Z(c[708]) );
  XNOR U4792 ( .A(n3445), .B(n3444), .Z(c[709]) );
  XNOR U4793 ( .A(n3447), .B(n3446), .Z(c[70]) );
  XNOR U4794 ( .A(n3449), .B(n3448), .Z(c[710]) );
  XNOR U4795 ( .A(n3451), .B(n3450), .Z(c[711]) );
  XNOR U4796 ( .A(n3453), .B(n3452), .Z(c[712]) );
  XNOR U4797 ( .A(n3455), .B(n3454), .Z(c[713]) );
  XNOR U4798 ( .A(n3457), .B(n3456), .Z(c[714]) );
  XNOR U4799 ( .A(n3459), .B(n3458), .Z(c[715]) );
  XNOR U4800 ( .A(n3461), .B(n3460), .Z(c[716]) );
  XNOR U4801 ( .A(n3463), .B(n3462), .Z(c[717]) );
  XNOR U4802 ( .A(n3465), .B(n3464), .Z(c[718]) );
  XNOR U4803 ( .A(n3467), .B(n3466), .Z(c[719]) );
  XNOR U4804 ( .A(n3469), .B(n3468), .Z(c[71]) );
  XNOR U4805 ( .A(n3471), .B(n3470), .Z(c[720]) );
  XNOR U4806 ( .A(n3473), .B(n3472), .Z(c[721]) );
  XNOR U4807 ( .A(n3475), .B(n3474), .Z(c[722]) );
  XNOR U4808 ( .A(n3477), .B(n3476), .Z(c[723]) );
  XNOR U4809 ( .A(n3479), .B(n3478), .Z(c[724]) );
  XNOR U4810 ( .A(n3481), .B(n3480), .Z(c[725]) );
  XNOR U4811 ( .A(n3483), .B(n3482), .Z(c[726]) );
  XNOR U4812 ( .A(n3485), .B(n3484), .Z(c[727]) );
  XNOR U4813 ( .A(n3487), .B(n3486), .Z(c[728]) );
  XNOR U4814 ( .A(n3489), .B(n3488), .Z(c[729]) );
  XNOR U4815 ( .A(n3491), .B(n3490), .Z(c[72]) );
  XNOR U4816 ( .A(n3493), .B(n3492), .Z(c[730]) );
  XNOR U4817 ( .A(n3495), .B(n3494), .Z(c[731]) );
  XNOR U4818 ( .A(n3497), .B(n3496), .Z(c[732]) );
  XNOR U4819 ( .A(n3499), .B(n3498), .Z(c[733]) );
  XNOR U4820 ( .A(n3501), .B(n3500), .Z(c[734]) );
  XNOR U4821 ( .A(n3503), .B(n3502), .Z(c[735]) );
  XNOR U4822 ( .A(n3505), .B(n3504), .Z(c[736]) );
  XNOR U4823 ( .A(n3507), .B(n3506), .Z(c[737]) );
  XNOR U4824 ( .A(n3509), .B(n3508), .Z(c[738]) );
  XNOR U4825 ( .A(n3511), .B(n3510), .Z(c[739]) );
  XNOR U4826 ( .A(n3513), .B(n3512), .Z(c[73]) );
  XNOR U4827 ( .A(n3515), .B(n3514), .Z(c[740]) );
  XNOR U4828 ( .A(n3517), .B(n3516), .Z(c[741]) );
  XNOR U4829 ( .A(n3519), .B(n3518), .Z(c[742]) );
  XNOR U4830 ( .A(n3521), .B(n3520), .Z(c[743]) );
  XNOR U4831 ( .A(n3523), .B(n3522), .Z(c[744]) );
  XNOR U4832 ( .A(n3525), .B(n3524), .Z(c[745]) );
  XNOR U4833 ( .A(n3527), .B(n3526), .Z(c[746]) );
  XNOR U4834 ( .A(n3529), .B(n3528), .Z(c[747]) );
  XNOR U4835 ( .A(n3531), .B(n3530), .Z(c[748]) );
  XNOR U4836 ( .A(n3533), .B(n3532), .Z(c[749]) );
  XNOR U4837 ( .A(n3535), .B(n3534), .Z(c[74]) );
  XNOR U4838 ( .A(n3537), .B(n3536), .Z(c[750]) );
  XNOR U4839 ( .A(n3539), .B(n3538), .Z(c[751]) );
  XNOR U4840 ( .A(n3541), .B(n3540), .Z(c[752]) );
  XNOR U4841 ( .A(n3543), .B(n3542), .Z(c[753]) );
  XNOR U4842 ( .A(n3545), .B(n3544), .Z(c[754]) );
  XNOR U4843 ( .A(n3547), .B(n3546), .Z(c[755]) );
  XNOR U4844 ( .A(n3549), .B(n3548), .Z(c[756]) );
  XNOR U4845 ( .A(n3551), .B(n3550), .Z(c[757]) );
  XNOR U4846 ( .A(n3553), .B(n3552), .Z(c[758]) );
  XNOR U4847 ( .A(n3555), .B(n3554), .Z(c[759]) );
  XNOR U4848 ( .A(n3557), .B(n3556), .Z(c[75]) );
  XNOR U4849 ( .A(n3559), .B(n3558), .Z(c[760]) );
  XNOR U4850 ( .A(n3561), .B(n3560), .Z(c[761]) );
  XNOR U4851 ( .A(n3563), .B(n3562), .Z(c[762]) );
  XNOR U4852 ( .A(n3565), .B(n3564), .Z(c[763]) );
  XNOR U4853 ( .A(n3567), .B(n3566), .Z(c[764]) );
  XNOR U4854 ( .A(n3569), .B(n3568), .Z(c[765]) );
  XNOR U4855 ( .A(n3571), .B(n3570), .Z(c[766]) );
  XNOR U4856 ( .A(n3573), .B(n3572), .Z(c[767]) );
  XNOR U4857 ( .A(n3575), .B(n3574), .Z(c[768]) );
  XNOR U4858 ( .A(n3577), .B(n3576), .Z(c[769]) );
  XNOR U4859 ( .A(n3579), .B(n3578), .Z(c[76]) );
  XNOR U4860 ( .A(n3581), .B(n3580), .Z(c[770]) );
  XNOR U4861 ( .A(n3583), .B(n3582), .Z(c[771]) );
  XNOR U4862 ( .A(n3585), .B(n3584), .Z(c[772]) );
  XNOR U4863 ( .A(n3587), .B(n3586), .Z(c[773]) );
  XNOR U4864 ( .A(n3589), .B(n3588), .Z(c[774]) );
  XNOR U4865 ( .A(n3591), .B(n3590), .Z(c[775]) );
  XNOR U4866 ( .A(n3593), .B(n3592), .Z(c[776]) );
  XNOR U4867 ( .A(n3595), .B(n3594), .Z(c[777]) );
  XNOR U4868 ( .A(n3597), .B(n3596), .Z(c[778]) );
  XNOR U4869 ( .A(n3599), .B(n3598), .Z(c[779]) );
  XNOR U4870 ( .A(n3601), .B(n3600), .Z(c[77]) );
  XNOR U4871 ( .A(n3603), .B(n3602), .Z(c[780]) );
  XNOR U4872 ( .A(n3605), .B(n3604), .Z(c[781]) );
  XNOR U4873 ( .A(n3607), .B(n3606), .Z(c[782]) );
  XNOR U4874 ( .A(n3609), .B(n3608), .Z(c[783]) );
  XNOR U4875 ( .A(n3611), .B(n3610), .Z(c[784]) );
  XNOR U4876 ( .A(n3613), .B(n3612), .Z(c[785]) );
  XNOR U4877 ( .A(n3615), .B(n3614), .Z(c[786]) );
  XNOR U4878 ( .A(n3617), .B(n3616), .Z(c[787]) );
  XNOR U4879 ( .A(n3619), .B(n3618), .Z(c[788]) );
  XNOR U4880 ( .A(n3621), .B(n3620), .Z(c[789]) );
  XNOR U4881 ( .A(n3623), .B(n3622), .Z(c[78]) );
  XNOR U4882 ( .A(n3625), .B(n3624), .Z(c[790]) );
  XNOR U4883 ( .A(n3627), .B(n3626), .Z(c[791]) );
  XNOR U4884 ( .A(n3629), .B(n3628), .Z(c[792]) );
  XNOR U4885 ( .A(n3631), .B(n3630), .Z(c[793]) );
  XNOR U4886 ( .A(n3633), .B(n3632), .Z(c[794]) );
  XNOR U4887 ( .A(n3635), .B(n3634), .Z(c[795]) );
  XNOR U4888 ( .A(n3637), .B(n3636), .Z(c[796]) );
  XNOR U4889 ( .A(n3639), .B(n3638), .Z(c[797]) );
  XNOR U4890 ( .A(n3641), .B(n3640), .Z(c[798]) );
  XNOR U4891 ( .A(n3643), .B(n3642), .Z(c[799]) );
  XNOR U4892 ( .A(n3645), .B(n3644), .Z(c[79]) );
  XNOR U4893 ( .A(n3647), .B(n3646), .Z(c[7]) );
  XNOR U4894 ( .A(n3649), .B(n3648), .Z(c[800]) );
  XNOR U4895 ( .A(n3651), .B(n3650), .Z(c[801]) );
  XNOR U4896 ( .A(n3653), .B(n3652), .Z(c[802]) );
  XNOR U4897 ( .A(n3655), .B(n3654), .Z(c[803]) );
  XNOR U4898 ( .A(n3657), .B(n3656), .Z(c[804]) );
  XNOR U4899 ( .A(n3659), .B(n3658), .Z(c[805]) );
  XNOR U4900 ( .A(n3661), .B(n3660), .Z(c[806]) );
  XNOR U4901 ( .A(n3663), .B(n3662), .Z(c[807]) );
  XNOR U4902 ( .A(n3665), .B(n3664), .Z(c[808]) );
  XNOR U4903 ( .A(n3667), .B(n3666), .Z(c[809]) );
  XNOR U4904 ( .A(n3669), .B(n3668), .Z(c[80]) );
  XNOR U4905 ( .A(n3671), .B(n3670), .Z(c[810]) );
  XNOR U4906 ( .A(n3673), .B(n3672), .Z(c[811]) );
  XNOR U4907 ( .A(n3675), .B(n3674), .Z(c[812]) );
  XNOR U4908 ( .A(n3677), .B(n3676), .Z(c[813]) );
  XNOR U4909 ( .A(n3679), .B(n3678), .Z(c[814]) );
  XNOR U4910 ( .A(n3681), .B(n3680), .Z(c[815]) );
  XNOR U4911 ( .A(n3683), .B(n3682), .Z(c[816]) );
  XNOR U4912 ( .A(n3685), .B(n3684), .Z(c[817]) );
  XNOR U4913 ( .A(n3687), .B(n3686), .Z(c[818]) );
  XNOR U4914 ( .A(n3689), .B(n3688), .Z(c[819]) );
  XNOR U4915 ( .A(n3691), .B(n3690), .Z(c[81]) );
  XNOR U4916 ( .A(n3693), .B(n3692), .Z(c[820]) );
  XNOR U4917 ( .A(n3695), .B(n3694), .Z(c[821]) );
  XNOR U4918 ( .A(n3697), .B(n3696), .Z(c[822]) );
  XNOR U4919 ( .A(n3699), .B(n3698), .Z(c[823]) );
  XNOR U4920 ( .A(n3701), .B(n3700), .Z(c[824]) );
  XNOR U4921 ( .A(n3703), .B(n3702), .Z(c[825]) );
  XNOR U4922 ( .A(n3705), .B(n3704), .Z(c[826]) );
  XNOR U4923 ( .A(n3707), .B(n3706), .Z(c[827]) );
  XNOR U4924 ( .A(n3709), .B(n3708), .Z(c[828]) );
  XNOR U4925 ( .A(n3711), .B(n3710), .Z(c[829]) );
  XNOR U4926 ( .A(n3713), .B(n3712), .Z(c[82]) );
  XNOR U4927 ( .A(n3715), .B(n3714), .Z(c[830]) );
  XNOR U4928 ( .A(n3717), .B(n3716), .Z(c[831]) );
  XNOR U4929 ( .A(n3719), .B(n3718), .Z(c[832]) );
  XNOR U4930 ( .A(n3721), .B(n3720), .Z(c[833]) );
  XNOR U4931 ( .A(n3723), .B(n3722), .Z(c[834]) );
  XNOR U4932 ( .A(n3725), .B(n3724), .Z(c[835]) );
  XNOR U4933 ( .A(n3727), .B(n3726), .Z(c[836]) );
  XNOR U4934 ( .A(n3729), .B(n3728), .Z(c[837]) );
  XNOR U4935 ( .A(n3731), .B(n3730), .Z(c[838]) );
  XNOR U4936 ( .A(n3733), .B(n3732), .Z(c[839]) );
  XNOR U4937 ( .A(n3735), .B(n3734), .Z(c[83]) );
  XNOR U4938 ( .A(n3737), .B(n3736), .Z(c[840]) );
  XNOR U4939 ( .A(n3739), .B(n3738), .Z(c[841]) );
  XNOR U4940 ( .A(n3741), .B(n3740), .Z(c[842]) );
  XNOR U4941 ( .A(n3743), .B(n3742), .Z(c[843]) );
  XNOR U4942 ( .A(n3745), .B(n3744), .Z(c[844]) );
  XNOR U4943 ( .A(n3747), .B(n3746), .Z(c[845]) );
  XNOR U4944 ( .A(n3749), .B(n3748), .Z(c[846]) );
  XNOR U4945 ( .A(n3751), .B(n3750), .Z(c[847]) );
  XNOR U4946 ( .A(n3753), .B(n3752), .Z(c[848]) );
  XNOR U4947 ( .A(n3755), .B(n3754), .Z(c[849]) );
  XNOR U4948 ( .A(n3757), .B(n3756), .Z(c[84]) );
  XNOR U4949 ( .A(n3759), .B(n3758), .Z(c[850]) );
  XNOR U4950 ( .A(n3761), .B(n3760), .Z(c[851]) );
  XNOR U4951 ( .A(n3763), .B(n3762), .Z(c[852]) );
  XNOR U4952 ( .A(n3765), .B(n3764), .Z(c[853]) );
  XNOR U4953 ( .A(n3767), .B(n3766), .Z(c[854]) );
  XNOR U4954 ( .A(n3769), .B(n3768), .Z(c[855]) );
  XNOR U4955 ( .A(n3771), .B(n3770), .Z(c[856]) );
  XNOR U4956 ( .A(n3773), .B(n3772), .Z(c[857]) );
  XNOR U4957 ( .A(n3775), .B(n3774), .Z(c[858]) );
  XNOR U4958 ( .A(n3777), .B(n3776), .Z(c[859]) );
  XNOR U4959 ( .A(n3779), .B(n3778), .Z(c[85]) );
  XNOR U4960 ( .A(n3781), .B(n3780), .Z(c[860]) );
  XNOR U4961 ( .A(n3783), .B(n3782), .Z(c[861]) );
  XNOR U4962 ( .A(n3785), .B(n3784), .Z(c[862]) );
  XNOR U4963 ( .A(n3787), .B(n3786), .Z(c[863]) );
  XNOR U4964 ( .A(n3789), .B(n3788), .Z(c[864]) );
  XNOR U4965 ( .A(n3791), .B(n3790), .Z(c[865]) );
  XNOR U4966 ( .A(n3793), .B(n3792), .Z(c[866]) );
  XNOR U4967 ( .A(n3795), .B(n3794), .Z(c[867]) );
  XNOR U4968 ( .A(n3797), .B(n3796), .Z(c[868]) );
  XNOR U4969 ( .A(n3799), .B(n3798), .Z(c[869]) );
  XNOR U4970 ( .A(n3801), .B(n3800), .Z(c[86]) );
  XNOR U4971 ( .A(n3803), .B(n3802), .Z(c[870]) );
  XNOR U4972 ( .A(n3805), .B(n3804), .Z(c[871]) );
  XNOR U4973 ( .A(n3807), .B(n3806), .Z(c[872]) );
  XNOR U4974 ( .A(n3809), .B(n3808), .Z(c[873]) );
  XNOR U4975 ( .A(n3811), .B(n3810), .Z(c[874]) );
  XNOR U4976 ( .A(n3813), .B(n3812), .Z(c[875]) );
  XNOR U4977 ( .A(n3815), .B(n3814), .Z(c[876]) );
  XNOR U4978 ( .A(n3817), .B(n3816), .Z(c[877]) );
  XNOR U4979 ( .A(n3819), .B(n3818), .Z(c[878]) );
  XNOR U4980 ( .A(n3821), .B(n3820), .Z(c[879]) );
  XNOR U4981 ( .A(n3823), .B(n3822), .Z(c[87]) );
  XNOR U4982 ( .A(n3825), .B(n3824), .Z(c[880]) );
  XNOR U4983 ( .A(n3827), .B(n3826), .Z(c[881]) );
  XNOR U4984 ( .A(n3829), .B(n3828), .Z(c[882]) );
  XNOR U4985 ( .A(n3831), .B(n3830), .Z(c[883]) );
  XNOR U4986 ( .A(n3833), .B(n3832), .Z(c[884]) );
  XNOR U4987 ( .A(n3835), .B(n3834), .Z(c[885]) );
  XNOR U4988 ( .A(n3837), .B(n3836), .Z(c[886]) );
  XNOR U4989 ( .A(n3839), .B(n3838), .Z(c[887]) );
  XNOR U4990 ( .A(n3841), .B(n3840), .Z(c[888]) );
  XNOR U4991 ( .A(n3843), .B(n3842), .Z(c[889]) );
  XNOR U4992 ( .A(n3845), .B(n3844), .Z(c[88]) );
  XNOR U4993 ( .A(n3847), .B(n3846), .Z(c[890]) );
  XNOR U4994 ( .A(n3849), .B(n3848), .Z(c[891]) );
  XNOR U4995 ( .A(n3851), .B(n3850), .Z(c[892]) );
  XNOR U4996 ( .A(n3853), .B(n3852), .Z(c[893]) );
  XNOR U4997 ( .A(n3855), .B(n3854), .Z(c[894]) );
  XNOR U4998 ( .A(n3857), .B(n3856), .Z(c[895]) );
  XNOR U4999 ( .A(n3859), .B(n3858), .Z(c[896]) );
  XNOR U5000 ( .A(n3861), .B(n3860), .Z(c[897]) );
  XNOR U5001 ( .A(n3863), .B(n3862), .Z(c[898]) );
  XNOR U5002 ( .A(n3865), .B(n3864), .Z(c[899]) );
  XNOR U5003 ( .A(n3867), .B(n3866), .Z(c[89]) );
  XNOR U5004 ( .A(n3869), .B(n3868), .Z(c[8]) );
  XNOR U5005 ( .A(n3871), .B(n3870), .Z(c[900]) );
  XNOR U5006 ( .A(n3873), .B(n3872), .Z(c[901]) );
  XNOR U5007 ( .A(n3875), .B(n3874), .Z(c[902]) );
  XNOR U5008 ( .A(n3877), .B(n3876), .Z(c[903]) );
  XNOR U5009 ( .A(n3879), .B(n3878), .Z(c[904]) );
  XNOR U5010 ( .A(n3881), .B(n3880), .Z(c[905]) );
  XNOR U5011 ( .A(n3883), .B(n3882), .Z(c[906]) );
  XNOR U5012 ( .A(n3885), .B(n3884), .Z(c[907]) );
  XNOR U5013 ( .A(n3887), .B(n3886), .Z(c[908]) );
  XNOR U5014 ( .A(n3889), .B(n3888), .Z(c[909]) );
  XNOR U5015 ( .A(n3891), .B(n3890), .Z(c[90]) );
  XNOR U5016 ( .A(n3893), .B(n3892), .Z(c[910]) );
  XNOR U5017 ( .A(n3895), .B(n3894), .Z(c[911]) );
  XNOR U5018 ( .A(n3897), .B(n3896), .Z(c[912]) );
  XNOR U5019 ( .A(n3899), .B(n3898), .Z(c[913]) );
  XNOR U5020 ( .A(n3901), .B(n3900), .Z(c[914]) );
  XNOR U5021 ( .A(n3903), .B(n3902), .Z(c[915]) );
  XNOR U5022 ( .A(n3905), .B(n3904), .Z(c[916]) );
  XNOR U5023 ( .A(n3907), .B(n3906), .Z(c[917]) );
  XNOR U5024 ( .A(n3909), .B(n3908), .Z(c[918]) );
  XNOR U5025 ( .A(n3911), .B(n3910), .Z(c[919]) );
  XNOR U5026 ( .A(n3913), .B(n3912), .Z(c[91]) );
  XNOR U5027 ( .A(n3915), .B(n3914), .Z(c[920]) );
  XNOR U5028 ( .A(n3917), .B(n3916), .Z(c[921]) );
  XNOR U5029 ( .A(n3919), .B(n3918), .Z(c[922]) );
  XNOR U5030 ( .A(n3921), .B(n3920), .Z(c[923]) );
  XNOR U5031 ( .A(n3923), .B(n3922), .Z(c[924]) );
  XNOR U5032 ( .A(n3925), .B(n3924), .Z(c[925]) );
  XNOR U5033 ( .A(n3927), .B(n3926), .Z(c[926]) );
  XNOR U5034 ( .A(n3929), .B(n3928), .Z(c[927]) );
  XNOR U5035 ( .A(n3931), .B(n3930), .Z(c[928]) );
  XNOR U5036 ( .A(n3933), .B(n3932), .Z(c[929]) );
  XNOR U5037 ( .A(n3935), .B(n3934), .Z(c[92]) );
  XNOR U5038 ( .A(n3937), .B(n3936), .Z(c[930]) );
  XNOR U5039 ( .A(n3939), .B(n3938), .Z(c[931]) );
  XNOR U5040 ( .A(n3941), .B(n3940), .Z(c[932]) );
  XNOR U5041 ( .A(n3943), .B(n3942), .Z(c[933]) );
  XNOR U5042 ( .A(n3945), .B(n3944), .Z(c[934]) );
  XNOR U5043 ( .A(n3947), .B(n3946), .Z(c[935]) );
  XNOR U5044 ( .A(n3949), .B(n3948), .Z(c[936]) );
  XNOR U5045 ( .A(n3951), .B(n3950), .Z(c[937]) );
  XNOR U5046 ( .A(n3953), .B(n3952), .Z(c[938]) );
  XNOR U5047 ( .A(n3955), .B(n3954), .Z(c[939]) );
  XNOR U5048 ( .A(n3957), .B(n3956), .Z(c[93]) );
  XNOR U5049 ( .A(n3959), .B(n3958), .Z(c[940]) );
  XNOR U5050 ( .A(n3961), .B(n3960), .Z(c[941]) );
  XNOR U5051 ( .A(n3963), .B(n3962), .Z(c[942]) );
  XNOR U5052 ( .A(n3965), .B(n3964), .Z(c[943]) );
  XNOR U5053 ( .A(n3967), .B(n3966), .Z(c[944]) );
  XNOR U5054 ( .A(n3969), .B(n3968), .Z(c[945]) );
  XNOR U5055 ( .A(n3971), .B(n3970), .Z(c[946]) );
  XNOR U5056 ( .A(n3973), .B(n3972), .Z(c[947]) );
  XNOR U5057 ( .A(n3975), .B(n3974), .Z(c[948]) );
  XNOR U5058 ( .A(n3977), .B(n3976), .Z(c[949]) );
  XNOR U5059 ( .A(n3979), .B(n3978), .Z(c[94]) );
  XNOR U5060 ( .A(n3981), .B(n3980), .Z(c[950]) );
  XNOR U5061 ( .A(n3983), .B(n3982), .Z(c[951]) );
  XNOR U5062 ( .A(n3985), .B(n3984), .Z(c[952]) );
  XNOR U5063 ( .A(n3987), .B(n3986), .Z(c[953]) );
  XNOR U5064 ( .A(n3989), .B(n3988), .Z(c[954]) );
  XNOR U5065 ( .A(n3991), .B(n3990), .Z(c[955]) );
  XNOR U5066 ( .A(n3993), .B(n3992), .Z(c[956]) );
  XNOR U5067 ( .A(n3995), .B(n3994), .Z(c[957]) );
  XNOR U5068 ( .A(n3997), .B(n3996), .Z(c[958]) );
  XNOR U5069 ( .A(n3999), .B(n3998), .Z(c[959]) );
  XNOR U5070 ( .A(n4001), .B(n4000), .Z(c[95]) );
  XNOR U5071 ( .A(n4003), .B(n4002), .Z(c[960]) );
  XNOR U5072 ( .A(n4005), .B(n4004), .Z(c[961]) );
  XNOR U5073 ( .A(n4007), .B(n4006), .Z(c[962]) );
  XNOR U5074 ( .A(n4009), .B(n4008), .Z(c[963]) );
  XNOR U5075 ( .A(n4011), .B(n4010), .Z(c[964]) );
  XNOR U5076 ( .A(n4013), .B(n4012), .Z(c[965]) );
  XNOR U5077 ( .A(n4015), .B(n4014), .Z(c[966]) );
  XNOR U5078 ( .A(n4017), .B(n4016), .Z(c[967]) );
  XNOR U5079 ( .A(n4019), .B(n4018), .Z(c[968]) );
  XNOR U5080 ( .A(n4021), .B(n4020), .Z(c[969]) );
  XNOR U5081 ( .A(n4023), .B(n4022), .Z(c[96]) );
  XNOR U5082 ( .A(n4025), .B(n4024), .Z(c[970]) );
  XNOR U5083 ( .A(n4027), .B(n4026), .Z(c[971]) );
  XNOR U5084 ( .A(n4029), .B(n4028), .Z(c[972]) );
  XNOR U5085 ( .A(n4031), .B(n4030), .Z(c[973]) );
  XNOR U5086 ( .A(n4033), .B(n4032), .Z(c[974]) );
  XNOR U5087 ( .A(n4035), .B(n4034), .Z(c[975]) );
  XNOR U5088 ( .A(n4037), .B(n4036), .Z(c[976]) );
  XNOR U5089 ( .A(n4039), .B(n4038), .Z(c[977]) );
  XNOR U5090 ( .A(n4041), .B(n4040), .Z(c[978]) );
  XNOR U5091 ( .A(n4043), .B(n4042), .Z(c[979]) );
  XNOR U5092 ( .A(n4045), .B(n4044), .Z(c[97]) );
  XNOR U5093 ( .A(n4047), .B(n4046), .Z(c[980]) );
  XNOR U5094 ( .A(n4049), .B(n4048), .Z(c[981]) );
  XNOR U5095 ( .A(n4051), .B(n4050), .Z(c[982]) );
  XNOR U5096 ( .A(n4053), .B(n4052), .Z(c[983]) );
  XNOR U5097 ( .A(n4055), .B(n4054), .Z(c[984]) );
  XNOR U5098 ( .A(n4057), .B(n4056), .Z(c[985]) );
  XNOR U5099 ( .A(n4059), .B(n4058), .Z(c[986]) );
  XNOR U5100 ( .A(n4061), .B(n4060), .Z(c[987]) );
  XNOR U5101 ( .A(n4063), .B(n4062), .Z(c[988]) );
  XNOR U5102 ( .A(n4065), .B(n4064), .Z(c[989]) );
  XNOR U5103 ( .A(n4067), .B(n4066), .Z(c[98]) );
  XNOR U5104 ( .A(n4069), .B(n4068), .Z(c[990]) );
  XNOR U5105 ( .A(n4071), .B(n4070), .Z(c[991]) );
  XNOR U5106 ( .A(n4073), .B(n4072), .Z(c[992]) );
  XNOR U5107 ( .A(n4075), .B(n4074), .Z(c[993]) );
  XNOR U5108 ( .A(n4077), .B(n4076), .Z(c[994]) );
  XNOR U5109 ( .A(n4079), .B(n4078), .Z(c[995]) );
  XNOR U5110 ( .A(n4081), .B(n4080), .Z(c[996]) );
  XNOR U5111 ( .A(n4083), .B(n4082), .Z(c[997]) );
  XNOR U5112 ( .A(n4085), .B(n4084), .Z(c[998]) );
  XOR U5113 ( .A(n4087), .B(n4086), .Z(c[999]) );
  XOR U5114 ( .A(n4089), .B(n4088), .Z(c[99]) );
  XOR U5115 ( .A(n4091), .B(n4090), .Z(c[9]) );
endmodule

