
module hamming_N16000_CC32_DW01_add_0 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45;

  XNOR U1 ( .A(A[9]), .B(n1), .Z(SUM[9]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[8]) );
  XNOR U3 ( .A(B[8]), .B(A[8]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[7]) );
  XNOR U5 ( .A(B[7]), .B(A[7]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[6]) );
  XNOR U7 ( .A(B[6]), .B(A[6]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[5]) );
  XNOR U9 ( .A(B[5]), .B(A[5]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U11 ( .A(B[4]), .B(A[4]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[3]) );
  XNOR U13 ( .A(B[3]), .B(A[3]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[2]) );
  XNOR U15 ( .A(B[2]), .B(A[2]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[1]) );
  XOR U17 ( .A(B[1]), .B(A[1]), .Z(n17) );
  XOR U18 ( .A(A[13]), .B(n18), .Z(SUM[13]) );
  ANDN U19 ( .B(A[12]), .A(n19), .Z(n18) );
  XNOR U20 ( .A(A[12]), .B(n19), .Z(SUM[12]) );
  NANDN U21 ( .A(n20), .B(A[11]), .Z(n19) );
  XNOR U22 ( .A(A[11]), .B(n20), .Z(SUM[11]) );
  NAND U23 ( .A(n21), .B(A[10]), .Z(n20) );
  XOR U24 ( .A(A[10]), .B(n21), .Z(SUM[10]) );
  ANDN U25 ( .B(A[9]), .A(n1), .Z(n21) );
  AND U26 ( .A(n22), .B(n23), .Z(n1) );
  NAND U27 ( .A(n24), .B(B[8]), .Z(n23) );
  NANDN U28 ( .A(A[8]), .B(n2), .Z(n24) );
  NANDN U29 ( .A(n2), .B(A[8]), .Z(n22) );
  AND U30 ( .A(n25), .B(n26), .Z(n2) );
  NAND U31 ( .A(n27), .B(B[7]), .Z(n26) );
  NANDN U32 ( .A(A[7]), .B(n4), .Z(n27) );
  NANDN U33 ( .A(n4), .B(A[7]), .Z(n25) );
  AND U34 ( .A(n28), .B(n29), .Z(n4) );
  NAND U35 ( .A(n30), .B(B[6]), .Z(n29) );
  NANDN U36 ( .A(A[6]), .B(n6), .Z(n30) );
  NANDN U37 ( .A(n6), .B(A[6]), .Z(n28) );
  AND U38 ( .A(n31), .B(n32), .Z(n6) );
  NAND U39 ( .A(n33), .B(B[5]), .Z(n32) );
  NANDN U40 ( .A(A[5]), .B(n8), .Z(n33) );
  NANDN U41 ( .A(n8), .B(A[5]), .Z(n31) );
  AND U42 ( .A(n34), .B(n35), .Z(n8) );
  NAND U43 ( .A(n36), .B(B[4]), .Z(n35) );
  NANDN U44 ( .A(A[4]), .B(n10), .Z(n36) );
  NANDN U45 ( .A(n10), .B(A[4]), .Z(n34) );
  AND U46 ( .A(n37), .B(n38), .Z(n10) );
  NAND U47 ( .A(n39), .B(B[3]), .Z(n38) );
  NANDN U48 ( .A(A[3]), .B(n12), .Z(n39) );
  NANDN U49 ( .A(n12), .B(A[3]), .Z(n37) );
  AND U50 ( .A(n40), .B(n41), .Z(n12) );
  NAND U51 ( .A(n42), .B(B[2]), .Z(n41) );
  NANDN U52 ( .A(A[2]), .B(n14), .Z(n42) );
  NANDN U53 ( .A(n14), .B(A[2]), .Z(n40) );
  AND U54 ( .A(n43), .B(n44), .Z(n14) );
  NAND U55 ( .A(n45), .B(B[1]), .Z(n44) );
  OR U56 ( .A(n16), .B(A[1]), .Z(n45) );
  NAND U57 ( .A(n16), .B(A[1]), .Z(n43) );
  AND U58 ( .A(B[0]), .B(A[0]), .Z(n16) );
  XOR U59 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC32_DW01_add_1 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37;

  IV U1 ( .A(B[8]), .Z(n1) );
  XOR U2 ( .A(n2), .B(n1), .Z(SUM[8]) );
  AND U3 ( .A(n3), .B(n4), .Z(n2) );
  NAND U4 ( .A(n5), .B(B[7]), .Z(n4) );
  NANDN U5 ( .A(A[7]), .B(n6), .Z(n5) );
  NANDN U6 ( .A(n6), .B(A[7]), .Z(n3) );
  XOR U7 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U8 ( .A(B[7]), .B(A[7]), .Z(n7) );
  AND U9 ( .A(n8), .B(n9), .Z(n6) );
  NAND U10 ( .A(n10), .B(B[6]), .Z(n9) );
  NANDN U11 ( .A(A[6]), .B(n11), .Z(n10) );
  NANDN U12 ( .A(n11), .B(A[6]), .Z(n8) );
  XOR U13 ( .A(n11), .B(n12), .Z(SUM[6]) );
  XNOR U14 ( .A(B[6]), .B(A[6]), .Z(n12) );
  AND U15 ( .A(n13), .B(n14), .Z(n11) );
  NAND U16 ( .A(n15), .B(B[5]), .Z(n14) );
  NANDN U17 ( .A(A[5]), .B(n16), .Z(n15) );
  NANDN U18 ( .A(n16), .B(A[5]), .Z(n13) );
  XOR U19 ( .A(n16), .B(n17), .Z(SUM[5]) );
  XNOR U20 ( .A(B[5]), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n18), .B(n19), .Z(n16) );
  NAND U22 ( .A(n20), .B(B[4]), .Z(n19) );
  NANDN U23 ( .A(A[4]), .B(n21), .Z(n20) );
  NANDN U24 ( .A(n21), .B(A[4]), .Z(n18) );
  XOR U25 ( .A(n21), .B(n22), .Z(SUM[4]) );
  XNOR U26 ( .A(B[4]), .B(A[4]), .Z(n22) );
  AND U27 ( .A(n23), .B(n24), .Z(n21) );
  NAND U28 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U29 ( .A(A[3]), .B(n26), .Z(n25) );
  NANDN U30 ( .A(n26), .B(A[3]), .Z(n23) );
  XOR U31 ( .A(n26), .B(n27), .Z(SUM[3]) );
  XNOR U32 ( .A(B[3]), .B(A[3]), .Z(n27) );
  AND U33 ( .A(n28), .B(n29), .Z(n26) );
  NAND U34 ( .A(n30), .B(B[2]), .Z(n29) );
  NANDN U35 ( .A(A[2]), .B(n31), .Z(n30) );
  NANDN U36 ( .A(n31), .B(A[2]), .Z(n28) );
  XOR U37 ( .A(n31), .B(n32), .Z(SUM[2]) );
  XNOR U38 ( .A(B[2]), .B(A[2]), .Z(n32) );
  AND U39 ( .A(n33), .B(n34), .Z(n31) );
  NAND U40 ( .A(n35), .B(B[1]), .Z(n34) );
  OR U41 ( .A(n36), .B(A[1]), .Z(n35) );
  NAND U42 ( .A(n36), .B(A[1]), .Z(n33) );
  XOR U43 ( .A(n36), .B(n37), .Z(SUM[1]) );
  XOR U44 ( .A(B[1]), .B(A[1]), .Z(n37) );
  AND U45 ( .A(B[0]), .B(A[0]), .Z(n36) );
  XOR U46 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC32_DW01_add_2 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[8]) );
  NAND U2 ( .A(n4), .B(B[7]), .Z(n3) );
  NANDN U3 ( .A(A[7]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[7]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[6]), .Z(n8) );
  NANDN U9 ( .A(A[6]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[6]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[6]) );
  XNOR U12 ( .A(B[6]), .B(A[6]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U15 ( .A(A[5]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[5]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[5]) );
  XNOR U18 ( .A(B[5]), .B(A[5]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[4]), .Z(n18) );
  NANDN U21 ( .A(A[4]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[4]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[4]) );
  XNOR U24 ( .A(B[4]), .B(A[4]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[3]), .Z(n23) );
  NANDN U27 ( .A(A[3]), .B(n25), .Z(n24) );
  NANDN U28 ( .A(n25), .B(A[3]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[3]) );
  XNOR U30 ( .A(B[3]), .B(A[3]), .Z(n26) );
  AND U31 ( .A(n27), .B(n28), .Z(n25) );
  NAND U32 ( .A(n29), .B(B[2]), .Z(n28) );
  NANDN U33 ( .A(A[2]), .B(n30), .Z(n29) );
  NANDN U34 ( .A(n30), .B(A[2]), .Z(n27) );
  XOR U35 ( .A(n30), .B(n31), .Z(SUM[2]) );
  XNOR U36 ( .A(B[2]), .B(A[2]), .Z(n31) );
  AND U37 ( .A(n32), .B(n33), .Z(n30) );
  NAND U38 ( .A(n34), .B(B[1]), .Z(n33) );
  OR U39 ( .A(n35), .B(A[1]), .Z(n34) );
  NAND U40 ( .A(n35), .B(A[1]), .Z(n32) );
  XOR U41 ( .A(n35), .B(n36), .Z(SUM[1]) );
  XOR U42 ( .A(B[1]), .B(A[1]), .Z(n36) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n35) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC32_DW01_add_3 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[7]) );
  NAND U2 ( .A(n4), .B(B[6]), .Z(n3) );
  NANDN U3 ( .A(A[6]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[6]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[5]), .Z(n8) );
  NANDN U9 ( .A(A[5]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[5]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U12 ( .A(B[5]), .B(A[5]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[4]), .Z(n13) );
  NANDN U15 ( .A(A[4]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[4]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[4]) );
  XNOR U18 ( .A(B[4]), .B(A[4]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[3]), .Z(n18) );
  NANDN U21 ( .A(A[3]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[3]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[3]) );
  XNOR U24 ( .A(B[3]), .B(A[3]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[2]), .Z(n23) );
  NANDN U27 ( .A(A[2]), .B(n25), .Z(n24) );
  NANDN U28 ( .A(n25), .B(A[2]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[2]) );
  XNOR U30 ( .A(B[2]), .B(A[2]), .Z(n26) );
  AND U31 ( .A(n27), .B(n28), .Z(n25) );
  NAND U32 ( .A(n29), .B(B[1]), .Z(n28) );
  OR U33 ( .A(n30), .B(A[1]), .Z(n29) );
  NAND U34 ( .A(n30), .B(A[1]), .Z(n27) );
  XOR U35 ( .A(n30), .B(n31), .Z(SUM[1]) );
  XOR U36 ( .A(B[1]), .B(A[1]), .Z(n31) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n30) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC32_DW01_add_4 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[7]) );
  NAND U2 ( .A(n4), .B(B[6]), .Z(n3) );
  NANDN U3 ( .A(A[6]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[6]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[5]), .Z(n8) );
  NANDN U9 ( .A(A[5]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[5]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U12 ( .A(B[5]), .B(A[5]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[4]), .Z(n13) );
  NANDN U15 ( .A(A[4]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[4]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[4]) );
  XNOR U18 ( .A(B[4]), .B(A[4]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[3]), .Z(n18) );
  NANDN U21 ( .A(A[3]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[3]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[3]) );
  XNOR U24 ( .A(B[3]), .B(A[3]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[2]), .Z(n23) );
  NANDN U27 ( .A(A[2]), .B(n25), .Z(n24) );
  NANDN U28 ( .A(n25), .B(A[2]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[2]) );
  XNOR U30 ( .A(B[2]), .B(A[2]), .Z(n26) );
  AND U31 ( .A(n27), .B(n28), .Z(n25) );
  NAND U32 ( .A(n29), .B(B[1]), .Z(n28) );
  OR U33 ( .A(n30), .B(A[1]), .Z(n29) );
  NAND U34 ( .A(n30), .B(A[1]), .Z(n27) );
  XOR U35 ( .A(n30), .B(n31), .Z(SUM[1]) );
  XOR U36 ( .A(B[1]), .B(A[1]), .Z(n31) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n30) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC32_DW01_add_5 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29;

  AND U1 ( .A(n2), .B(B[6]), .Z(SUM[7]) );
  IV U2 ( .A(n4), .Z(n2) );
  IV U3 ( .A(B[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n3), .Z(SUM[6]) );
  AND U5 ( .A(n5), .B(n6), .Z(n4) );
  NAND U6 ( .A(n7), .B(B[5]), .Z(n6) );
  NANDN U7 ( .A(A[5]), .B(n8), .Z(n7) );
  NANDN U8 ( .A(n8), .B(A[5]), .Z(n5) );
  XOR U9 ( .A(n8), .B(n9), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n9) );
  AND U11 ( .A(n10), .B(n11), .Z(n8) );
  NAND U12 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U13 ( .A(A[4]), .B(n13), .Z(n12) );
  NANDN U14 ( .A(n13), .B(A[4]), .Z(n10) );
  XOR U15 ( .A(n13), .B(n14), .Z(SUM[4]) );
  XNOR U16 ( .A(B[4]), .B(A[4]), .Z(n14) );
  AND U17 ( .A(n15), .B(n16), .Z(n13) );
  NAND U18 ( .A(n17), .B(B[3]), .Z(n16) );
  NANDN U19 ( .A(A[3]), .B(n18), .Z(n17) );
  NANDN U20 ( .A(n18), .B(A[3]), .Z(n15) );
  XOR U21 ( .A(n18), .B(n19), .Z(SUM[3]) );
  XNOR U22 ( .A(B[3]), .B(A[3]), .Z(n19) );
  AND U23 ( .A(n20), .B(n21), .Z(n18) );
  NAND U24 ( .A(n22), .B(B[2]), .Z(n21) );
  NANDN U25 ( .A(A[2]), .B(n23), .Z(n22) );
  NANDN U26 ( .A(n23), .B(A[2]), .Z(n20) );
  XOR U27 ( .A(n23), .B(n24), .Z(SUM[2]) );
  XNOR U28 ( .A(B[2]), .B(A[2]), .Z(n24) );
  AND U29 ( .A(n25), .B(n26), .Z(n23) );
  NAND U30 ( .A(n27), .B(B[1]), .Z(n26) );
  OR U31 ( .A(n28), .B(A[1]), .Z(n27) );
  NAND U32 ( .A(n28), .B(A[1]), .Z(n25) );
  XOR U33 ( .A(n28), .B(n29), .Z(SUM[1]) );
  XOR U34 ( .A(B[1]), .B(A[1]), .Z(n29) );
  AND U35 ( .A(B[0]), .B(A[0]), .Z(n28) );
  XOR U36 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC32_DW01_add_6 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[6]) );
  NAND U2 ( .A(n4), .B(B[5]), .Z(n3) );
  NANDN U3 ( .A(A[5]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[5]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[5]) );
  XNOR U6 ( .A(B[5]), .B(A[5]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[4]), .Z(n8) );
  NANDN U9 ( .A(A[4]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[4]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[3]), .Z(n13) );
  NANDN U15 ( .A(A[3]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[3]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[3]) );
  XNOR U18 ( .A(B[3]), .B(A[3]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[2]), .Z(n18) );
  NANDN U21 ( .A(A[2]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[2]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[2]) );
  XNOR U24 ( .A(B[2]), .B(A[2]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[1]), .Z(n23) );
  OR U27 ( .A(n25), .B(A[1]), .Z(n24) );
  NAND U28 ( .A(n25), .B(A[1]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[1]) );
  XOR U30 ( .A(B[1]), .B(A[1]), .Z(n26) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n25) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC32_DW01_add_7 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[6]) );
  NAND U2 ( .A(n4), .B(B[5]), .Z(n3) );
  NANDN U3 ( .A(A[5]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[5]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[5]) );
  XNOR U6 ( .A(B[5]), .B(A[5]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[4]), .Z(n8) );
  NANDN U9 ( .A(A[4]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[4]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[3]), .Z(n13) );
  NANDN U15 ( .A(A[3]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[3]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[3]) );
  XNOR U18 ( .A(B[3]), .B(A[3]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[2]), .Z(n18) );
  NANDN U21 ( .A(A[2]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[2]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[2]) );
  XNOR U24 ( .A(B[2]), .B(A[2]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[1]), .Z(n23) );
  OR U27 ( .A(n25), .B(A[1]), .Z(n24) );
  NAND U28 ( .A(n25), .B(A[1]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[1]) );
  XOR U30 ( .A(B[1]), .B(A[1]), .Z(n26) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n25) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC32_DW01_add_8 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[6]) );
  NAND U2 ( .A(n4), .B(B[5]), .Z(n3) );
  NANDN U3 ( .A(A[5]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[5]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[5]) );
  XNOR U6 ( .A(B[5]), .B(A[5]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[4]), .Z(n8) );
  NANDN U9 ( .A(A[4]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[4]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[3]), .Z(n13) );
  NANDN U15 ( .A(A[3]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[3]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[3]) );
  XNOR U18 ( .A(B[3]), .B(A[3]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[2]), .Z(n18) );
  NANDN U21 ( .A(A[2]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[2]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[2]) );
  XNOR U24 ( .A(B[2]), .B(A[2]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[1]), .Z(n23) );
  OR U27 ( .A(n25), .B(A[1]), .Z(n24) );
  NAND U28 ( .A(n25), .B(A[1]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[1]) );
  XOR U30 ( .A(B[1]), .B(A[1]), .Z(n26) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n25) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC32_DW01_add_9 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[6]) );
  NAND U2 ( .A(n4), .B(B[5]), .Z(n3) );
  NANDN U3 ( .A(A[5]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[5]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[5]) );
  XNOR U6 ( .A(B[5]), .B(A[5]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[4]), .Z(n8) );
  NANDN U9 ( .A(A[4]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[4]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[3]), .Z(n13) );
  NANDN U15 ( .A(A[3]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[3]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[3]) );
  XNOR U18 ( .A(B[3]), .B(A[3]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[2]), .Z(n18) );
  NANDN U21 ( .A(A[2]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[2]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[2]) );
  XNOR U24 ( .A(B[2]), .B(A[2]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[1]), .Z(n23) );
  OR U27 ( .A(n25), .B(A[1]), .Z(n24) );
  NAND U28 ( .A(n25), .B(A[1]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[1]) );
  XOR U30 ( .A(B[1]), .B(A[1]), .Z(n26) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n25) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC32_DW01_add_10 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24;

  AND U1 ( .A(n3), .B(B[5]), .Z(SUM[6]) );
  IV U2 ( .A(B[5]), .Z(n2) );
  IV U3 ( .A(n4), .Z(n3) );
  XOR U4 ( .A(n4), .B(n2), .Z(SUM[5]) );
  AND U5 ( .A(n5), .B(n6), .Z(n4) );
  NAND U6 ( .A(n7), .B(B[4]), .Z(n6) );
  NANDN U7 ( .A(A[4]), .B(n8), .Z(n7) );
  NANDN U8 ( .A(n8), .B(A[4]), .Z(n5) );
  XOR U9 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U10 ( .A(B[4]), .B(A[4]), .Z(n9) );
  AND U11 ( .A(n10), .B(n11), .Z(n8) );
  NAND U12 ( .A(n12), .B(B[3]), .Z(n11) );
  NANDN U13 ( .A(A[3]), .B(n13), .Z(n12) );
  NANDN U14 ( .A(n13), .B(A[3]), .Z(n10) );
  XOR U15 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U16 ( .A(B[3]), .B(A[3]), .Z(n14) );
  AND U17 ( .A(n15), .B(n16), .Z(n13) );
  NAND U18 ( .A(n17), .B(B[2]), .Z(n16) );
  NANDN U19 ( .A(A[2]), .B(n18), .Z(n17) );
  NANDN U20 ( .A(n18), .B(A[2]), .Z(n15) );
  XOR U21 ( .A(n18), .B(n19), .Z(SUM[2]) );
  XNOR U22 ( .A(B[2]), .B(A[2]), .Z(n19) );
  AND U23 ( .A(n20), .B(n21), .Z(n18) );
  NAND U24 ( .A(n22), .B(B[1]), .Z(n21) );
  OR U25 ( .A(n23), .B(A[1]), .Z(n22) );
  NAND U26 ( .A(n23), .B(A[1]), .Z(n20) );
  XOR U27 ( .A(n23), .B(n24), .Z(SUM[1]) );
  XOR U28 ( .A(B[1]), .B(A[1]), .Z(n24) );
  AND U29 ( .A(B[0]), .B(A[0]), .Z(n23) );
  XOR U30 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC32_DW01_add_11 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC32_DW01_add_12 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC32_DW01_add_13 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC32_DW01_add_14 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC32_DW01_add_15 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC32_DW01_add_16 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC32_DW01_add_17 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC32_DW01_add_18 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC32_DW01_add_19 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC32_DW01_add_20 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC32 ( clk, rst, x, y, o );
  input [499:0] x;
  input [499:0] y;
  output [13:0] o;
  input clk, rst;
  wire   N2591, N2592, N2593, N2594, N2595, N2600, N2601, N2602, N2603, N2604,
         N2609, N2610, N2611, N2612, N2613, N2618, N2619, N2620, N2621, N2622,
         N2627, N2628, N2629, N2630, N2631, N2636, N2637, N2638, N2639, N2640,
         N2645, N2646, N2647, N2648, N2649, N2654, N2655, N2656, N2657, N2658,
         N2663, N2664, N2665, N2666, N2667, N2672, N2673, N2674, N2675, N2676,
         N2681, N2682, N2683, N2684, N2685, N2690, N2691, N2692, N2693, N2694,
         N2699, N2700, N2701, N2702, N2703, N2708, N2709, N2710, N2711, N2712,
         N2717, N2718, N2719, N2720, N2721, N2726, N2727, N2728, N2729, N2730,
         N2735, N2736, N2737, N2738, N2739, N2744, N2745, N2746, N2747, N2748,
         N2753, N2754, N2755, N2756, N2757, N2762, N2763, N2764, N2765, N2766,
         N2771, N2772, N2773, N2774, N2775, N2780, N2781, N2782, N2783, N2784,
         N2785, N2789, N2790, N2791, N2792, N2793, N2794, N2798, N2799, N2800,
         N2801, N2802, N2803, N2807, N2808, N2809, N2810, N2811, N2812, N2816,
         N2817, N2818, N2819, N2820, N2821, N2825, N2826, N2827, N2828, N2829,
         N2830, N2834, N2835, N2836, N2837, N2838, N2839, N2843, N2844, N2845,
         N2846, N2847, N2848, N2852, N2853, N2854, N2855, N2856, N2857, N2861,
         N2862, N2863, N2864, N2865, N2866, N2870, N2871, N2872, N2873, N2874,
         N2875, N2876, N2879, N2880, N2881, N2882, N2883, N2884, N2885, N2888,
         N2889, N2890, N2891, N2892, N2893, N2894, N2897, N2898, N2899, N2900,
         N2901, N2902, N2903, N2906, N2907, N2908, N2909, N2910, N2911, N2912,
         N2915, N2916, N2917, N2918, N2919, N2920, N2921, N2922, N2924, N2925,
         N2926, N2927, N2928, N2929, N2930, N2931, N2933, N2934, N2935, N2936,
         N2937, N2938, N2939, N2940, N2942, N2943, N2944, N2945, N2946, N2947,
         N2948, N2949, N2950, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411;
  wire   [8:0] olocal;
  wire   [13:0] oglobal;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42;

  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .Q(oglobal[11]) );
  DFF \oglobal_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .Q(oglobal[12]) );
  DFF \oglobal_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .Q(oglobal[13]) );
  hamming_N16000_CC32_DW01_add_0 add_97 ( .A(oglobal), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, olocal}), .CI(1'b0), .SUM(o) );
  hamming_N16000_CC32_DW01_add_1 add_167_root_add_47_I500 ( .A({1'b0, N2940, 
        N2939, N2938, N2937, N2936, N2935, N2934, N2933}), .B({N2950, N2949, 
        N2948, N2947, N2946, N2945, N2944, N2943, N2942}), .CI(1'b0), .SUM(
        olocal) );
  hamming_N16000_CC32_DW01_add_2 add_168_root_add_47_I500 ( .A({1'b0, N2922, 
        N2921, N2920, N2919, N2918, N2917, N2916, N2915}), .B({1'b0, N2931, 
        N2930, N2929, N2928, N2927, N2926, N2925, N2924}), .CI(1'b0), .SUM({
        N2950, N2949, N2948, N2947, N2946, N2945, N2944, N2943, N2942}) );
  hamming_N16000_CC32_DW01_add_3 add_169_root_add_47_I500 ( .A({1'b0, 1'b0, 
        N2903, N2902, N2901, N2900, N2899, N2898, N2897}), .B({1'b0, 1'b0, 
        N2912, N2911, N2910, N2909, N2908, N2907, N2906}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, N2940, N2939, N2938, N2937, N2936, N2935, 
        N2934, N2933}) );
  hamming_N16000_CC32_DW01_add_4 add_170_root_add_47_I500 ( .A({1'b0, 1'b0, 
        N2885, N2884, N2883, N2882, N2881, N2880, N2879}), .B({1'b0, 1'b0, 
        N2894, N2893, N2892, N2891, N2890, N2889, N2888}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1, N2931, N2930, N2929, N2928, N2927, N2926, 
        N2925, N2924}) );
  hamming_N16000_CC32_DW01_add_5 add_171_root_add_47_I500 ( .A({1'b0, 1'b0, 
        1'b0, N2866, N2865, N2864, N2863, N2862, N2861}), .B({1'b0, 1'b0, 
        N2876, N2875, N2874, N2873, N2872, N2871, N2870}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__2, N2922, N2921, N2920, N2919, N2918, N2917, 
        N2916, N2915}) );
  hamming_N16000_CC32_DW01_add_6 add_172_root_add_47_I500 ( .A({1'b0, 1'b0, 
        1'b0, N2848, N2847, N2846, N2845, N2844, N2843}), .B({1'b0, 1'b0, 1'b0, 
        N2857, N2856, N2855, N2854, N2853, N2852}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, N2912, N2911, N2910, 
        N2909, N2908, N2907, N2906}) );
  hamming_N16000_CC32_DW01_add_7 add_173_root_add_47_I500 ( .A({1'b0, 1'b0, 
        1'b0, N2830, N2829, N2828, N2827, N2826, N2825}), .B({1'b0, 1'b0, 1'b0, 
        N2839, N2838, N2837, N2836, N2835, N2834}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, N2903, N2902, N2901, 
        N2900, N2899, N2898, N2897}) );
  hamming_N16000_CC32_DW01_add_8 add_174_root_add_47_I500 ( .A({1'b0, 1'b0, 
        1'b0, N2812, N2811, N2810, N2809, N2808, N2807}), .B({1'b0, 1'b0, 1'b0, 
        N2821, N2820, N2819, N2818, N2817, N2816}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, N2894, N2893, N2892, 
        N2891, N2890, N2889, N2888}) );
  hamming_N16000_CC32_DW01_add_9 add_175_root_add_47_I500 ( .A({1'b0, 1'b0, 
        1'b0, N2794, N2793, N2792, N2791, N2790, N2789}), .B({1'b0, 1'b0, 1'b0, 
        N2803, N2802, N2801, N2800, N2799, N2798}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, N2885, N2884, N2883, 
        N2882, N2881, N2880, N2879}) );
  hamming_N16000_CC32_DW01_add_10 add_176_root_add_47_I500 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N2775, N2774, N2773, N2772, N2771}), .B({1'b0, 1'b0, 1'b0, 
        N2785, N2784, N2783, N2782, N2781, N2780}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, N2876, N2875, 
        N2874, N2873, N2872, N2871, N2870}) );
  hamming_N16000_CC32_DW01_add_11 add_177_root_add_47_I500 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N2757, N2756, N2755, N2754, N2753}), .B({1'b0, 1'b0, 1'b0, 
        1'b0, N2766, N2765, N2764, N2763, N2762}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N2866, N2865, N2864, N2863, N2862, N2861})
         );
  hamming_N16000_CC32_DW01_add_12 add_178_root_add_47_I500 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N2739, N2738, N2737, N2736, N2735}), .B({1'b0, 1'b0, 1'b0, 
        1'b0, N2748, N2747, N2746, N2745, N2744}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, N2857, N2856, N2855, N2854, N2853, N2852})
         );
  hamming_N16000_CC32_DW01_add_13 add_179_root_add_47_I500 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N2721, N2720, N2719, N2718, N2717}), .B({1'b0, 1'b0, 1'b0, 
        1'b0, N2730, N2729, N2728, N2727, N2726}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, N2848, N2847, N2846, N2845, N2844, N2843})
         );
  hamming_N16000_CC32_DW01_add_14 add_180_root_add_47_I500 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N2703, N2702, N2701, N2700, N2699}), .B({1'b0, 1'b0, 1'b0, 
        1'b0, N2712, N2711, N2710, N2709, N2708}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, N2839, N2838, N2837, N2836, N2835, N2834})
         );
  hamming_N16000_CC32_DW01_add_15 add_181_root_add_47_I500 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N2685, N2684, N2683, N2682, N2681}), .B({1'b0, 1'b0, 1'b0, 
        1'b0, N2694, N2693, N2692, N2691, N2690}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, N2830, N2829, N2828, N2827, N2826, N2825})
         );
  hamming_N16000_CC32_DW01_add_16 add_182_root_add_47_I500 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N2667, N2666, N2665, N2664, N2663}), .B({1'b0, 1'b0, 1'b0, 
        1'b0, N2676, N2675, N2674, N2673, N2672}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, N2821, N2820, N2819, N2818, N2817, N2816})
         );
  hamming_N16000_CC32_DW01_add_17 add_183_root_add_47_I500 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N2649, N2648, N2647, N2646, N2645}), .B({1'b0, 1'b0, 1'b0, 
        1'b0, N2658, N2657, N2656, N2655, N2654}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, N2812, N2811, N2810, N2809, N2808, N2807})
         );
  hamming_N16000_CC32_DW01_add_18 add_184_root_add_47_I500 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N2631, N2630, N2629, N2628, N2627}), .B({1'b0, 1'b0, 1'b0, 
        1'b0, N2640, N2639, N2638, N2637, N2636}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, N2803, N2802, N2801, N2800, N2799, N2798})
         );
  hamming_N16000_CC32_DW01_add_19 add_185_root_add_47_I500 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N2613, N2612, N2611, N2610, N2609}), .B({1'b0, 1'b0, 1'b0, 
        1'b0, N2622, N2621, N2620, N2619, N2618}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, N2794, N2793, N2792, N2791, N2790, N2789})
         );
  hamming_N16000_CC32_DW01_add_20 add_186_root_add_47_I500 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N2595, N2594, N2593, N2592, N2591}), .B({1'b0, 1'b0, 1'b0, 
        1'b0, N2604, N2603, N2602, N2601, N2600}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, N2785, N2784, N2783, N2782, N2781, N2780})
         );
  NAND U853 ( .A(n354), .B(n355), .Z(N2775) );
  NANDN U854 ( .A(n356), .B(n357), .Z(n355) );
  OR U855 ( .A(n358), .B(n359), .Z(n357) );
  NAND U856 ( .A(n358), .B(n359), .Z(n354) );
  XOR U857 ( .A(n358), .B(n360), .Z(N2774) );
  XNOR U858 ( .A(n356), .B(n359), .Z(n360) );
  AND U859 ( .A(n361), .B(n362), .Z(n359) );
  NANDN U860 ( .A(n363), .B(n364), .Z(n362) );
  NANDN U861 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U862 ( .A(n366), .B(n365), .Z(n361) );
  NAND U863 ( .A(n367), .B(n368), .Z(n356) );
  NANDN U864 ( .A(n369), .B(n370), .Z(n368) );
  OR U865 ( .A(n371), .B(n372), .Z(n370) );
  NAND U866 ( .A(n372), .B(n371), .Z(n367) );
  AND U867 ( .A(n373), .B(n374), .Z(n358) );
  NANDN U868 ( .A(n375), .B(n376), .Z(n374) );
  NANDN U869 ( .A(n377), .B(n378), .Z(n376) );
  NANDN U870 ( .A(n378), .B(n377), .Z(n373) );
  XOR U871 ( .A(n372), .B(n379), .Z(N2773) );
  XOR U872 ( .A(n369), .B(n371), .Z(n379) );
  XNOR U873 ( .A(n365), .B(n380), .Z(n371) );
  XNOR U874 ( .A(n363), .B(n366), .Z(n380) );
  NAND U875 ( .A(n381), .B(n382), .Z(n366) );
  NAND U876 ( .A(n383), .B(n384), .Z(n382) );
  OR U877 ( .A(n385), .B(n386), .Z(n383) );
  NANDN U878 ( .A(n387), .B(n385), .Z(n381) );
  IV U879 ( .A(n386), .Z(n387) );
  NAND U880 ( .A(n388), .B(n389), .Z(n363) );
  NAND U881 ( .A(n390), .B(n391), .Z(n389) );
  NANDN U882 ( .A(n392), .B(n393), .Z(n390) );
  NANDN U883 ( .A(n393), .B(n392), .Z(n388) );
  AND U884 ( .A(n394), .B(n395), .Z(n365) );
  NAND U885 ( .A(n396), .B(n397), .Z(n395) );
  OR U886 ( .A(n398), .B(n399), .Z(n396) );
  NANDN U887 ( .A(n400), .B(n398), .Z(n394) );
  NAND U888 ( .A(n401), .B(n402), .Z(n369) );
  NANDN U889 ( .A(n403), .B(n404), .Z(n402) );
  OR U890 ( .A(n405), .B(n406), .Z(n404) );
  NANDN U891 ( .A(n407), .B(n405), .Z(n401) );
  IV U892 ( .A(n406), .Z(n407) );
  XNOR U893 ( .A(n377), .B(n408), .Z(n372) );
  XNOR U894 ( .A(n375), .B(n378), .Z(n408) );
  NAND U895 ( .A(n409), .B(n410), .Z(n378) );
  NAND U896 ( .A(n411), .B(n412), .Z(n410) );
  OR U897 ( .A(n413), .B(n414), .Z(n411) );
  NANDN U898 ( .A(n415), .B(n413), .Z(n409) );
  IV U899 ( .A(n414), .Z(n415) );
  NAND U900 ( .A(n416), .B(n417), .Z(n375) );
  NAND U901 ( .A(n418), .B(n419), .Z(n417) );
  NANDN U902 ( .A(n420), .B(n421), .Z(n418) );
  NANDN U903 ( .A(n421), .B(n420), .Z(n416) );
  AND U904 ( .A(n422), .B(n423), .Z(n377) );
  NAND U905 ( .A(n424), .B(n425), .Z(n423) );
  OR U906 ( .A(n426), .B(n427), .Z(n424) );
  NANDN U907 ( .A(n428), .B(n426), .Z(n422) );
  XNOR U908 ( .A(n403), .B(n429), .Z(N2772) );
  XOR U909 ( .A(n405), .B(n406), .Z(n429) );
  XNOR U910 ( .A(n419), .B(n430), .Z(n406) );
  XOR U911 ( .A(n420), .B(n421), .Z(n430) );
  XOR U912 ( .A(n426), .B(n431), .Z(n421) );
  XOR U913 ( .A(n425), .B(n428), .Z(n431) );
  IV U914 ( .A(n427), .Z(n428) );
  NAND U915 ( .A(n432), .B(n433), .Z(n427) );
  OR U916 ( .A(n434), .B(n435), .Z(n433) );
  OR U917 ( .A(n436), .B(n437), .Z(n432) );
  NAND U918 ( .A(n438), .B(n439), .Z(n425) );
  OR U919 ( .A(n440), .B(n441), .Z(n439) );
  OR U920 ( .A(n442), .B(n443), .Z(n438) );
  NOR U921 ( .A(n444), .B(n445), .Z(n426) );
  ANDN U922 ( .B(n446), .A(n447), .Z(n420) );
  XNOR U923 ( .A(n413), .B(n448), .Z(n419) );
  XNOR U924 ( .A(n412), .B(n414), .Z(n448) );
  NAND U925 ( .A(n449), .B(n450), .Z(n414) );
  OR U926 ( .A(n451), .B(n452), .Z(n450) );
  OR U927 ( .A(n453), .B(n454), .Z(n449) );
  NAND U928 ( .A(n455), .B(n456), .Z(n412) );
  OR U929 ( .A(n457), .B(n458), .Z(n456) );
  OR U930 ( .A(n459), .B(n460), .Z(n455) );
  ANDN U931 ( .B(n461), .A(n462), .Z(n413) );
  IV U932 ( .A(n463), .Z(n461) );
  ANDN U933 ( .B(n464), .A(n465), .Z(n405) );
  XOR U934 ( .A(n391), .B(n466), .Z(n403) );
  XOR U935 ( .A(n392), .B(n393), .Z(n466) );
  XOR U936 ( .A(n398), .B(n467), .Z(n393) );
  XOR U937 ( .A(n397), .B(n400), .Z(n467) );
  IV U938 ( .A(n399), .Z(n400) );
  NAND U939 ( .A(n468), .B(n469), .Z(n399) );
  OR U940 ( .A(n470), .B(n471), .Z(n469) );
  OR U941 ( .A(n472), .B(n473), .Z(n468) );
  NAND U942 ( .A(n474), .B(n475), .Z(n397) );
  OR U943 ( .A(n476), .B(n477), .Z(n475) );
  OR U944 ( .A(n478), .B(n479), .Z(n474) );
  NOR U945 ( .A(n480), .B(n481), .Z(n398) );
  ANDN U946 ( .B(n482), .A(n483), .Z(n392) );
  IV U947 ( .A(n484), .Z(n482) );
  XNOR U948 ( .A(n385), .B(n485), .Z(n391) );
  XNOR U949 ( .A(n384), .B(n386), .Z(n485) );
  NAND U950 ( .A(n486), .B(n487), .Z(n386) );
  OR U951 ( .A(n488), .B(n489), .Z(n487) );
  OR U952 ( .A(n490), .B(n491), .Z(n486) );
  NAND U953 ( .A(n492), .B(n493), .Z(n384) );
  OR U954 ( .A(n494), .B(n495), .Z(n493) );
  OR U955 ( .A(n496), .B(n497), .Z(n492) );
  ANDN U956 ( .B(n498), .A(n499), .Z(n385) );
  IV U957 ( .A(n500), .Z(n498) );
  XNOR U958 ( .A(n465), .B(n464), .Z(N2771) );
  XOR U959 ( .A(n484), .B(n483), .Z(n464) );
  XNOR U960 ( .A(n499), .B(n500), .Z(n483) );
  XNOR U961 ( .A(n494), .B(n495), .Z(n500) );
  XNOR U962 ( .A(n496), .B(n497), .Z(n495) );
  XNOR U963 ( .A(y[493]), .B(x[493]), .Z(n497) );
  XNOR U964 ( .A(y[494]), .B(x[494]), .Z(n496) );
  XNOR U965 ( .A(y[492]), .B(x[492]), .Z(n494) );
  XNOR U966 ( .A(n488), .B(n489), .Z(n499) );
  XNOR U967 ( .A(y[489]), .B(x[489]), .Z(n489) );
  XNOR U968 ( .A(n490), .B(n491), .Z(n488) );
  XNOR U969 ( .A(y[490]), .B(x[490]), .Z(n491) );
  XNOR U970 ( .A(y[491]), .B(x[491]), .Z(n490) );
  XNOR U971 ( .A(n481), .B(n480), .Z(n484) );
  XNOR U972 ( .A(n476), .B(n477), .Z(n480) );
  XNOR U973 ( .A(y[486]), .B(x[486]), .Z(n477) );
  XNOR U974 ( .A(n478), .B(n479), .Z(n476) );
  XNOR U975 ( .A(y[487]), .B(x[487]), .Z(n479) );
  XNOR U976 ( .A(y[488]), .B(x[488]), .Z(n478) );
  XNOR U977 ( .A(n470), .B(n471), .Z(n481) );
  XNOR U978 ( .A(y[483]), .B(x[483]), .Z(n471) );
  XNOR U979 ( .A(n472), .B(n473), .Z(n470) );
  XNOR U980 ( .A(y[484]), .B(x[484]), .Z(n473) );
  XNOR U981 ( .A(y[485]), .B(x[485]), .Z(n472) );
  XOR U982 ( .A(n446), .B(n447), .Z(n465) );
  XNOR U983 ( .A(n462), .B(n463), .Z(n447) );
  XNOR U984 ( .A(n457), .B(n458), .Z(n463) );
  XNOR U985 ( .A(n459), .B(n460), .Z(n458) );
  XNOR U986 ( .A(y[481]), .B(x[481]), .Z(n460) );
  XNOR U987 ( .A(y[482]), .B(x[482]), .Z(n459) );
  XNOR U988 ( .A(y[480]), .B(x[480]), .Z(n457) );
  XNOR U989 ( .A(n451), .B(n452), .Z(n462) );
  XNOR U990 ( .A(y[477]), .B(x[477]), .Z(n452) );
  XNOR U991 ( .A(n453), .B(n454), .Z(n451) );
  XNOR U992 ( .A(y[478]), .B(x[478]), .Z(n454) );
  XNOR U993 ( .A(y[479]), .B(x[479]), .Z(n453) );
  XOR U994 ( .A(n445), .B(n444), .Z(n446) );
  XNOR U995 ( .A(n440), .B(n441), .Z(n444) );
  XNOR U996 ( .A(y[474]), .B(x[474]), .Z(n441) );
  XNOR U997 ( .A(n442), .B(n443), .Z(n440) );
  XNOR U998 ( .A(y[475]), .B(x[475]), .Z(n443) );
  XNOR U999 ( .A(y[476]), .B(x[476]), .Z(n442) );
  XNOR U1000 ( .A(n434), .B(n435), .Z(n445) );
  XNOR U1001 ( .A(y[471]), .B(x[471]), .Z(n435) );
  XNOR U1002 ( .A(n436), .B(n437), .Z(n434) );
  XNOR U1003 ( .A(y[472]), .B(x[472]), .Z(n437) );
  XNOR U1004 ( .A(y[473]), .B(x[473]), .Z(n436) );
  NAND U1005 ( .A(n501), .B(n502), .Z(N2766) );
  NANDN U1006 ( .A(n503), .B(n504), .Z(n502) );
  OR U1007 ( .A(n505), .B(n506), .Z(n504) );
  NAND U1008 ( .A(n505), .B(n506), .Z(n501) );
  XOR U1009 ( .A(n505), .B(n507), .Z(N2765) );
  XNOR U1010 ( .A(n503), .B(n506), .Z(n507) );
  AND U1011 ( .A(n508), .B(n509), .Z(n506) );
  NANDN U1012 ( .A(n510), .B(n511), .Z(n509) );
  NANDN U1013 ( .A(n512), .B(n513), .Z(n511) );
  NANDN U1014 ( .A(n513), .B(n512), .Z(n508) );
  NAND U1015 ( .A(n514), .B(n515), .Z(n503) );
  NANDN U1016 ( .A(n516), .B(n517), .Z(n515) );
  OR U1017 ( .A(n518), .B(n519), .Z(n517) );
  NAND U1018 ( .A(n519), .B(n518), .Z(n514) );
  AND U1019 ( .A(n520), .B(n521), .Z(n505) );
  NANDN U1020 ( .A(n522), .B(n523), .Z(n521) );
  NANDN U1021 ( .A(n524), .B(n525), .Z(n523) );
  NANDN U1022 ( .A(n525), .B(n524), .Z(n520) );
  XOR U1023 ( .A(n519), .B(n526), .Z(N2764) );
  XOR U1024 ( .A(n516), .B(n518), .Z(n526) );
  XNOR U1025 ( .A(n512), .B(n527), .Z(n518) );
  XNOR U1026 ( .A(n510), .B(n513), .Z(n527) );
  NAND U1027 ( .A(n528), .B(n529), .Z(n513) );
  NAND U1028 ( .A(n530), .B(n531), .Z(n529) );
  OR U1029 ( .A(n532), .B(n533), .Z(n530) );
  NANDN U1030 ( .A(n534), .B(n532), .Z(n528) );
  IV U1031 ( .A(n533), .Z(n534) );
  NAND U1032 ( .A(n535), .B(n536), .Z(n510) );
  NAND U1033 ( .A(n537), .B(n538), .Z(n536) );
  NANDN U1034 ( .A(n539), .B(n540), .Z(n537) );
  NANDN U1035 ( .A(n540), .B(n539), .Z(n535) );
  AND U1036 ( .A(n541), .B(n542), .Z(n512) );
  NAND U1037 ( .A(n543), .B(n544), .Z(n542) );
  OR U1038 ( .A(n545), .B(n546), .Z(n543) );
  NANDN U1039 ( .A(n547), .B(n545), .Z(n541) );
  NAND U1040 ( .A(n548), .B(n549), .Z(n516) );
  NANDN U1041 ( .A(n550), .B(n551), .Z(n549) );
  OR U1042 ( .A(n552), .B(n553), .Z(n551) );
  NANDN U1043 ( .A(n554), .B(n552), .Z(n548) );
  IV U1044 ( .A(n553), .Z(n554) );
  XNOR U1045 ( .A(n524), .B(n555), .Z(n519) );
  XNOR U1046 ( .A(n522), .B(n525), .Z(n555) );
  NAND U1047 ( .A(n556), .B(n557), .Z(n525) );
  NAND U1048 ( .A(n558), .B(n559), .Z(n557) );
  OR U1049 ( .A(n560), .B(n561), .Z(n558) );
  NANDN U1050 ( .A(n562), .B(n560), .Z(n556) );
  IV U1051 ( .A(n561), .Z(n562) );
  NAND U1052 ( .A(n563), .B(n564), .Z(n522) );
  NAND U1053 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U1054 ( .A(n567), .B(n568), .Z(n565) );
  NANDN U1055 ( .A(n568), .B(n567), .Z(n563) );
  AND U1056 ( .A(n569), .B(n570), .Z(n524) );
  NAND U1057 ( .A(n571), .B(n572), .Z(n570) );
  OR U1058 ( .A(n573), .B(n574), .Z(n571) );
  NANDN U1059 ( .A(n575), .B(n573), .Z(n569) );
  XNOR U1060 ( .A(n550), .B(n576), .Z(N2763) );
  XOR U1061 ( .A(n552), .B(n553), .Z(n576) );
  XNOR U1062 ( .A(n566), .B(n577), .Z(n553) );
  XOR U1063 ( .A(n567), .B(n568), .Z(n577) );
  XOR U1064 ( .A(n573), .B(n578), .Z(n568) );
  XOR U1065 ( .A(n572), .B(n575), .Z(n578) );
  IV U1066 ( .A(n574), .Z(n575) );
  NAND U1067 ( .A(n579), .B(n580), .Z(n574) );
  OR U1068 ( .A(n581), .B(n582), .Z(n580) );
  OR U1069 ( .A(n583), .B(n584), .Z(n579) );
  NAND U1070 ( .A(n585), .B(n586), .Z(n572) );
  OR U1071 ( .A(n587), .B(n588), .Z(n586) );
  OR U1072 ( .A(n589), .B(n590), .Z(n585) );
  NOR U1073 ( .A(n591), .B(n592), .Z(n573) );
  ANDN U1074 ( .B(n593), .A(n594), .Z(n567) );
  XNOR U1075 ( .A(n560), .B(n595), .Z(n566) );
  XNOR U1076 ( .A(n559), .B(n561), .Z(n595) );
  NAND U1077 ( .A(n596), .B(n597), .Z(n561) );
  OR U1078 ( .A(n598), .B(n599), .Z(n597) );
  OR U1079 ( .A(n600), .B(n601), .Z(n596) );
  NAND U1080 ( .A(n602), .B(n603), .Z(n559) );
  OR U1081 ( .A(n604), .B(n605), .Z(n603) );
  OR U1082 ( .A(n606), .B(n607), .Z(n602) );
  ANDN U1083 ( .B(n608), .A(n609), .Z(n560) );
  IV U1084 ( .A(n610), .Z(n608) );
  ANDN U1085 ( .B(n611), .A(n612), .Z(n552) );
  XOR U1086 ( .A(n538), .B(n613), .Z(n550) );
  XOR U1087 ( .A(n539), .B(n540), .Z(n613) );
  XOR U1088 ( .A(n545), .B(n614), .Z(n540) );
  XOR U1089 ( .A(n544), .B(n547), .Z(n614) );
  IV U1090 ( .A(n546), .Z(n547) );
  NAND U1091 ( .A(n615), .B(n616), .Z(n546) );
  OR U1092 ( .A(n617), .B(n618), .Z(n616) );
  OR U1093 ( .A(n619), .B(n620), .Z(n615) );
  NAND U1094 ( .A(n621), .B(n622), .Z(n544) );
  OR U1095 ( .A(n623), .B(n624), .Z(n622) );
  OR U1096 ( .A(n625), .B(n626), .Z(n621) );
  NOR U1097 ( .A(n627), .B(n628), .Z(n545) );
  ANDN U1098 ( .B(n629), .A(n630), .Z(n539) );
  IV U1099 ( .A(n631), .Z(n629) );
  XNOR U1100 ( .A(n532), .B(n632), .Z(n538) );
  XNOR U1101 ( .A(n531), .B(n533), .Z(n632) );
  NAND U1102 ( .A(n633), .B(n634), .Z(n533) );
  OR U1103 ( .A(n635), .B(n636), .Z(n634) );
  OR U1104 ( .A(n637), .B(n638), .Z(n633) );
  NAND U1105 ( .A(n639), .B(n640), .Z(n531) );
  OR U1106 ( .A(n641), .B(n642), .Z(n640) );
  OR U1107 ( .A(n643), .B(n644), .Z(n639) );
  ANDN U1108 ( .B(n645), .A(n646), .Z(n532) );
  IV U1109 ( .A(n647), .Z(n645) );
  XNOR U1110 ( .A(n612), .B(n611), .Z(N2762) );
  XOR U1111 ( .A(n631), .B(n630), .Z(n611) );
  XNOR U1112 ( .A(n646), .B(n647), .Z(n630) );
  XNOR U1113 ( .A(n641), .B(n642), .Z(n647) );
  XNOR U1114 ( .A(n643), .B(n644), .Z(n642) );
  XNOR U1115 ( .A(y[469]), .B(x[469]), .Z(n644) );
  XNOR U1116 ( .A(y[470]), .B(x[470]), .Z(n643) );
  XNOR U1117 ( .A(y[468]), .B(x[468]), .Z(n641) );
  XNOR U1118 ( .A(n635), .B(n636), .Z(n646) );
  XNOR U1119 ( .A(y[465]), .B(x[465]), .Z(n636) );
  XNOR U1120 ( .A(n637), .B(n638), .Z(n635) );
  XNOR U1121 ( .A(y[466]), .B(x[466]), .Z(n638) );
  XNOR U1122 ( .A(y[467]), .B(x[467]), .Z(n637) );
  XNOR U1123 ( .A(n628), .B(n627), .Z(n631) );
  XNOR U1124 ( .A(n623), .B(n624), .Z(n627) );
  XNOR U1125 ( .A(y[462]), .B(x[462]), .Z(n624) );
  XNOR U1126 ( .A(n625), .B(n626), .Z(n623) );
  XNOR U1127 ( .A(y[463]), .B(x[463]), .Z(n626) );
  XNOR U1128 ( .A(y[464]), .B(x[464]), .Z(n625) );
  XNOR U1129 ( .A(n617), .B(n618), .Z(n628) );
  XNOR U1130 ( .A(y[459]), .B(x[459]), .Z(n618) );
  XNOR U1131 ( .A(n619), .B(n620), .Z(n617) );
  XNOR U1132 ( .A(y[460]), .B(x[460]), .Z(n620) );
  XNOR U1133 ( .A(y[461]), .B(x[461]), .Z(n619) );
  XOR U1134 ( .A(n593), .B(n594), .Z(n612) );
  XNOR U1135 ( .A(n609), .B(n610), .Z(n594) );
  XNOR U1136 ( .A(n604), .B(n605), .Z(n610) );
  XNOR U1137 ( .A(n606), .B(n607), .Z(n605) );
  XNOR U1138 ( .A(y[457]), .B(x[457]), .Z(n607) );
  XNOR U1139 ( .A(y[458]), .B(x[458]), .Z(n606) );
  XNOR U1140 ( .A(y[456]), .B(x[456]), .Z(n604) );
  XNOR U1141 ( .A(n598), .B(n599), .Z(n609) );
  XNOR U1142 ( .A(y[453]), .B(x[453]), .Z(n599) );
  XNOR U1143 ( .A(n600), .B(n601), .Z(n598) );
  XNOR U1144 ( .A(y[454]), .B(x[454]), .Z(n601) );
  XNOR U1145 ( .A(y[455]), .B(x[455]), .Z(n600) );
  XOR U1146 ( .A(n592), .B(n591), .Z(n593) );
  XNOR U1147 ( .A(n587), .B(n588), .Z(n591) );
  XNOR U1148 ( .A(y[450]), .B(x[450]), .Z(n588) );
  XNOR U1149 ( .A(n589), .B(n590), .Z(n587) );
  XNOR U1150 ( .A(y[451]), .B(x[451]), .Z(n590) );
  XNOR U1151 ( .A(y[452]), .B(x[452]), .Z(n589) );
  XNOR U1152 ( .A(n581), .B(n582), .Z(n592) );
  XNOR U1153 ( .A(y[447]), .B(x[447]), .Z(n582) );
  XNOR U1154 ( .A(n583), .B(n584), .Z(n581) );
  XNOR U1155 ( .A(y[448]), .B(x[448]), .Z(n584) );
  XNOR U1156 ( .A(y[449]), .B(x[449]), .Z(n583) );
  NAND U1157 ( .A(n648), .B(n649), .Z(N2757) );
  NANDN U1158 ( .A(n650), .B(n651), .Z(n649) );
  OR U1159 ( .A(n652), .B(n653), .Z(n651) );
  NAND U1160 ( .A(n652), .B(n653), .Z(n648) );
  XOR U1161 ( .A(n652), .B(n654), .Z(N2756) );
  XNOR U1162 ( .A(n650), .B(n653), .Z(n654) );
  AND U1163 ( .A(n655), .B(n656), .Z(n653) );
  NANDN U1164 ( .A(n657), .B(n658), .Z(n656) );
  NANDN U1165 ( .A(n659), .B(n660), .Z(n658) );
  NANDN U1166 ( .A(n660), .B(n659), .Z(n655) );
  NAND U1167 ( .A(n661), .B(n662), .Z(n650) );
  NANDN U1168 ( .A(n663), .B(n664), .Z(n662) );
  OR U1169 ( .A(n665), .B(n666), .Z(n664) );
  NAND U1170 ( .A(n666), .B(n665), .Z(n661) );
  AND U1171 ( .A(n667), .B(n668), .Z(n652) );
  NANDN U1172 ( .A(n669), .B(n670), .Z(n668) );
  NANDN U1173 ( .A(n671), .B(n672), .Z(n670) );
  NANDN U1174 ( .A(n672), .B(n671), .Z(n667) );
  XOR U1175 ( .A(n666), .B(n673), .Z(N2755) );
  XOR U1176 ( .A(n663), .B(n665), .Z(n673) );
  XNOR U1177 ( .A(n659), .B(n674), .Z(n665) );
  XNOR U1178 ( .A(n657), .B(n660), .Z(n674) );
  NAND U1179 ( .A(n675), .B(n676), .Z(n660) );
  NAND U1180 ( .A(n677), .B(n678), .Z(n676) );
  OR U1181 ( .A(n679), .B(n680), .Z(n677) );
  NANDN U1182 ( .A(n681), .B(n679), .Z(n675) );
  IV U1183 ( .A(n680), .Z(n681) );
  NAND U1184 ( .A(n682), .B(n683), .Z(n657) );
  NAND U1185 ( .A(n684), .B(n685), .Z(n683) );
  NANDN U1186 ( .A(n686), .B(n687), .Z(n684) );
  NANDN U1187 ( .A(n687), .B(n686), .Z(n682) );
  AND U1188 ( .A(n688), .B(n689), .Z(n659) );
  NAND U1189 ( .A(n690), .B(n691), .Z(n689) );
  OR U1190 ( .A(n692), .B(n693), .Z(n690) );
  NANDN U1191 ( .A(n694), .B(n692), .Z(n688) );
  NAND U1192 ( .A(n695), .B(n696), .Z(n663) );
  NANDN U1193 ( .A(n697), .B(n698), .Z(n696) );
  OR U1194 ( .A(n699), .B(n700), .Z(n698) );
  NANDN U1195 ( .A(n701), .B(n699), .Z(n695) );
  IV U1196 ( .A(n700), .Z(n701) );
  XNOR U1197 ( .A(n671), .B(n702), .Z(n666) );
  XNOR U1198 ( .A(n669), .B(n672), .Z(n702) );
  NAND U1199 ( .A(n703), .B(n704), .Z(n672) );
  NAND U1200 ( .A(n705), .B(n706), .Z(n704) );
  OR U1201 ( .A(n707), .B(n708), .Z(n705) );
  NANDN U1202 ( .A(n709), .B(n707), .Z(n703) );
  IV U1203 ( .A(n708), .Z(n709) );
  NAND U1204 ( .A(n710), .B(n711), .Z(n669) );
  NAND U1205 ( .A(n712), .B(n713), .Z(n711) );
  NANDN U1206 ( .A(n714), .B(n715), .Z(n712) );
  NANDN U1207 ( .A(n715), .B(n714), .Z(n710) );
  AND U1208 ( .A(n716), .B(n717), .Z(n671) );
  NAND U1209 ( .A(n718), .B(n719), .Z(n717) );
  OR U1210 ( .A(n720), .B(n721), .Z(n718) );
  NANDN U1211 ( .A(n722), .B(n720), .Z(n716) );
  XNOR U1212 ( .A(n697), .B(n723), .Z(N2754) );
  XOR U1213 ( .A(n699), .B(n700), .Z(n723) );
  XNOR U1214 ( .A(n713), .B(n724), .Z(n700) );
  XOR U1215 ( .A(n714), .B(n715), .Z(n724) );
  XOR U1216 ( .A(n720), .B(n725), .Z(n715) );
  XOR U1217 ( .A(n719), .B(n722), .Z(n725) );
  IV U1218 ( .A(n721), .Z(n722) );
  NAND U1219 ( .A(n726), .B(n727), .Z(n721) );
  OR U1220 ( .A(n728), .B(n729), .Z(n727) );
  OR U1221 ( .A(n730), .B(n731), .Z(n726) );
  NAND U1222 ( .A(n732), .B(n733), .Z(n719) );
  OR U1223 ( .A(n734), .B(n735), .Z(n733) );
  OR U1224 ( .A(n736), .B(n737), .Z(n732) );
  NOR U1225 ( .A(n738), .B(n739), .Z(n720) );
  ANDN U1226 ( .B(n740), .A(n741), .Z(n714) );
  XNOR U1227 ( .A(n707), .B(n742), .Z(n713) );
  XNOR U1228 ( .A(n706), .B(n708), .Z(n742) );
  NAND U1229 ( .A(n743), .B(n744), .Z(n708) );
  OR U1230 ( .A(n745), .B(n746), .Z(n744) );
  OR U1231 ( .A(n747), .B(n748), .Z(n743) );
  NAND U1232 ( .A(n749), .B(n750), .Z(n706) );
  OR U1233 ( .A(n751), .B(n752), .Z(n750) );
  OR U1234 ( .A(n753), .B(n754), .Z(n749) );
  ANDN U1235 ( .B(n755), .A(n756), .Z(n707) );
  IV U1236 ( .A(n757), .Z(n755) );
  ANDN U1237 ( .B(n758), .A(n759), .Z(n699) );
  XOR U1238 ( .A(n685), .B(n760), .Z(n697) );
  XOR U1239 ( .A(n686), .B(n687), .Z(n760) );
  XOR U1240 ( .A(n692), .B(n761), .Z(n687) );
  XOR U1241 ( .A(n691), .B(n694), .Z(n761) );
  IV U1242 ( .A(n693), .Z(n694) );
  NAND U1243 ( .A(n762), .B(n763), .Z(n693) );
  OR U1244 ( .A(n764), .B(n765), .Z(n763) );
  OR U1245 ( .A(n766), .B(n767), .Z(n762) );
  NAND U1246 ( .A(n768), .B(n769), .Z(n691) );
  OR U1247 ( .A(n770), .B(n771), .Z(n769) );
  OR U1248 ( .A(n772), .B(n773), .Z(n768) );
  NOR U1249 ( .A(n774), .B(n775), .Z(n692) );
  ANDN U1250 ( .B(n776), .A(n777), .Z(n686) );
  IV U1251 ( .A(n778), .Z(n776) );
  XNOR U1252 ( .A(n679), .B(n779), .Z(n685) );
  XNOR U1253 ( .A(n678), .B(n680), .Z(n779) );
  NAND U1254 ( .A(n780), .B(n781), .Z(n680) );
  OR U1255 ( .A(n782), .B(n783), .Z(n781) );
  OR U1256 ( .A(n784), .B(n785), .Z(n780) );
  NAND U1257 ( .A(n786), .B(n787), .Z(n678) );
  OR U1258 ( .A(n788), .B(n789), .Z(n787) );
  OR U1259 ( .A(n790), .B(n791), .Z(n786) );
  ANDN U1260 ( .B(n792), .A(n793), .Z(n679) );
  IV U1261 ( .A(n794), .Z(n792) );
  XNOR U1262 ( .A(n759), .B(n758), .Z(N2753) );
  XOR U1263 ( .A(n778), .B(n777), .Z(n758) );
  XNOR U1264 ( .A(n793), .B(n794), .Z(n777) );
  XNOR U1265 ( .A(n788), .B(n789), .Z(n794) );
  XNOR U1266 ( .A(n790), .B(n791), .Z(n789) );
  XNOR U1267 ( .A(y[445]), .B(x[445]), .Z(n791) );
  XNOR U1268 ( .A(y[446]), .B(x[446]), .Z(n790) );
  XNOR U1269 ( .A(y[444]), .B(x[444]), .Z(n788) );
  XNOR U1270 ( .A(n782), .B(n783), .Z(n793) );
  XNOR U1271 ( .A(y[441]), .B(x[441]), .Z(n783) );
  XNOR U1272 ( .A(n784), .B(n785), .Z(n782) );
  XNOR U1273 ( .A(y[442]), .B(x[442]), .Z(n785) );
  XNOR U1274 ( .A(y[443]), .B(x[443]), .Z(n784) );
  XNOR U1275 ( .A(n775), .B(n774), .Z(n778) );
  XNOR U1276 ( .A(n770), .B(n771), .Z(n774) );
  XNOR U1277 ( .A(y[438]), .B(x[438]), .Z(n771) );
  XNOR U1278 ( .A(n772), .B(n773), .Z(n770) );
  XNOR U1279 ( .A(y[439]), .B(x[439]), .Z(n773) );
  XNOR U1280 ( .A(y[440]), .B(x[440]), .Z(n772) );
  XNOR U1281 ( .A(n764), .B(n765), .Z(n775) );
  XNOR U1282 ( .A(y[435]), .B(x[435]), .Z(n765) );
  XNOR U1283 ( .A(n766), .B(n767), .Z(n764) );
  XNOR U1284 ( .A(y[436]), .B(x[436]), .Z(n767) );
  XNOR U1285 ( .A(y[437]), .B(x[437]), .Z(n766) );
  XOR U1286 ( .A(n740), .B(n741), .Z(n759) );
  XNOR U1287 ( .A(n756), .B(n757), .Z(n741) );
  XNOR U1288 ( .A(n751), .B(n752), .Z(n757) );
  XNOR U1289 ( .A(n753), .B(n754), .Z(n752) );
  XNOR U1290 ( .A(y[433]), .B(x[433]), .Z(n754) );
  XNOR U1291 ( .A(y[434]), .B(x[434]), .Z(n753) );
  XNOR U1292 ( .A(y[432]), .B(x[432]), .Z(n751) );
  XNOR U1293 ( .A(n745), .B(n746), .Z(n756) );
  XNOR U1294 ( .A(y[429]), .B(x[429]), .Z(n746) );
  XNOR U1295 ( .A(n747), .B(n748), .Z(n745) );
  XNOR U1296 ( .A(y[430]), .B(x[430]), .Z(n748) );
  XNOR U1297 ( .A(y[431]), .B(x[431]), .Z(n747) );
  XOR U1298 ( .A(n739), .B(n738), .Z(n740) );
  XNOR U1299 ( .A(n734), .B(n735), .Z(n738) );
  XNOR U1300 ( .A(y[426]), .B(x[426]), .Z(n735) );
  XNOR U1301 ( .A(n736), .B(n737), .Z(n734) );
  XNOR U1302 ( .A(y[427]), .B(x[427]), .Z(n737) );
  XNOR U1303 ( .A(y[428]), .B(x[428]), .Z(n736) );
  XNOR U1304 ( .A(n728), .B(n729), .Z(n739) );
  XNOR U1305 ( .A(y[423]), .B(x[423]), .Z(n729) );
  XNOR U1306 ( .A(n730), .B(n731), .Z(n728) );
  XNOR U1307 ( .A(y[424]), .B(x[424]), .Z(n731) );
  XNOR U1308 ( .A(y[425]), .B(x[425]), .Z(n730) );
  NAND U1309 ( .A(n795), .B(n796), .Z(N2748) );
  NANDN U1310 ( .A(n797), .B(n798), .Z(n796) );
  OR U1311 ( .A(n799), .B(n800), .Z(n798) );
  NAND U1312 ( .A(n799), .B(n800), .Z(n795) );
  XOR U1313 ( .A(n799), .B(n801), .Z(N2747) );
  XNOR U1314 ( .A(n797), .B(n800), .Z(n801) );
  AND U1315 ( .A(n802), .B(n803), .Z(n800) );
  NANDN U1316 ( .A(n804), .B(n805), .Z(n803) );
  NANDN U1317 ( .A(n806), .B(n807), .Z(n805) );
  NANDN U1318 ( .A(n807), .B(n806), .Z(n802) );
  NAND U1319 ( .A(n808), .B(n809), .Z(n797) );
  NANDN U1320 ( .A(n810), .B(n811), .Z(n809) );
  OR U1321 ( .A(n812), .B(n813), .Z(n811) );
  NAND U1322 ( .A(n813), .B(n812), .Z(n808) );
  AND U1323 ( .A(n814), .B(n815), .Z(n799) );
  NANDN U1324 ( .A(n816), .B(n817), .Z(n815) );
  NANDN U1325 ( .A(n818), .B(n819), .Z(n817) );
  NANDN U1326 ( .A(n819), .B(n818), .Z(n814) );
  XOR U1327 ( .A(n813), .B(n820), .Z(N2746) );
  XOR U1328 ( .A(n810), .B(n812), .Z(n820) );
  XNOR U1329 ( .A(n806), .B(n821), .Z(n812) );
  XNOR U1330 ( .A(n804), .B(n807), .Z(n821) );
  NAND U1331 ( .A(n822), .B(n823), .Z(n807) );
  NAND U1332 ( .A(n824), .B(n825), .Z(n823) );
  OR U1333 ( .A(n826), .B(n827), .Z(n824) );
  NANDN U1334 ( .A(n828), .B(n826), .Z(n822) );
  IV U1335 ( .A(n827), .Z(n828) );
  NAND U1336 ( .A(n829), .B(n830), .Z(n804) );
  NAND U1337 ( .A(n831), .B(n832), .Z(n830) );
  NANDN U1338 ( .A(n833), .B(n834), .Z(n831) );
  NANDN U1339 ( .A(n834), .B(n833), .Z(n829) );
  AND U1340 ( .A(n835), .B(n836), .Z(n806) );
  NAND U1341 ( .A(n837), .B(n838), .Z(n836) );
  OR U1342 ( .A(n839), .B(n840), .Z(n837) );
  NANDN U1343 ( .A(n841), .B(n839), .Z(n835) );
  NAND U1344 ( .A(n842), .B(n843), .Z(n810) );
  NANDN U1345 ( .A(n844), .B(n845), .Z(n843) );
  OR U1346 ( .A(n846), .B(n847), .Z(n845) );
  NANDN U1347 ( .A(n848), .B(n846), .Z(n842) );
  IV U1348 ( .A(n847), .Z(n848) );
  XNOR U1349 ( .A(n818), .B(n849), .Z(n813) );
  XNOR U1350 ( .A(n816), .B(n819), .Z(n849) );
  NAND U1351 ( .A(n850), .B(n851), .Z(n819) );
  NAND U1352 ( .A(n852), .B(n853), .Z(n851) );
  OR U1353 ( .A(n854), .B(n855), .Z(n852) );
  NANDN U1354 ( .A(n856), .B(n854), .Z(n850) );
  IV U1355 ( .A(n855), .Z(n856) );
  NAND U1356 ( .A(n857), .B(n858), .Z(n816) );
  NAND U1357 ( .A(n859), .B(n860), .Z(n858) );
  NANDN U1358 ( .A(n861), .B(n862), .Z(n859) );
  NANDN U1359 ( .A(n862), .B(n861), .Z(n857) );
  AND U1360 ( .A(n863), .B(n864), .Z(n818) );
  NAND U1361 ( .A(n865), .B(n866), .Z(n864) );
  OR U1362 ( .A(n867), .B(n868), .Z(n865) );
  NANDN U1363 ( .A(n869), .B(n867), .Z(n863) );
  XNOR U1364 ( .A(n844), .B(n870), .Z(N2745) );
  XOR U1365 ( .A(n846), .B(n847), .Z(n870) );
  XNOR U1366 ( .A(n860), .B(n871), .Z(n847) );
  XOR U1367 ( .A(n861), .B(n862), .Z(n871) );
  XOR U1368 ( .A(n867), .B(n872), .Z(n862) );
  XOR U1369 ( .A(n866), .B(n869), .Z(n872) );
  IV U1370 ( .A(n868), .Z(n869) );
  NAND U1371 ( .A(n873), .B(n874), .Z(n868) );
  OR U1372 ( .A(n875), .B(n876), .Z(n874) );
  OR U1373 ( .A(n877), .B(n878), .Z(n873) );
  NAND U1374 ( .A(n879), .B(n880), .Z(n866) );
  OR U1375 ( .A(n881), .B(n882), .Z(n880) );
  OR U1376 ( .A(n883), .B(n884), .Z(n879) );
  NOR U1377 ( .A(n885), .B(n886), .Z(n867) );
  ANDN U1378 ( .B(n887), .A(n888), .Z(n861) );
  XNOR U1379 ( .A(n854), .B(n889), .Z(n860) );
  XNOR U1380 ( .A(n853), .B(n855), .Z(n889) );
  NAND U1381 ( .A(n890), .B(n891), .Z(n855) );
  OR U1382 ( .A(n892), .B(n893), .Z(n891) );
  OR U1383 ( .A(n894), .B(n895), .Z(n890) );
  NAND U1384 ( .A(n896), .B(n897), .Z(n853) );
  OR U1385 ( .A(n898), .B(n899), .Z(n897) );
  OR U1386 ( .A(n900), .B(n901), .Z(n896) );
  ANDN U1387 ( .B(n902), .A(n903), .Z(n854) );
  IV U1388 ( .A(n904), .Z(n902) );
  ANDN U1389 ( .B(n905), .A(n906), .Z(n846) );
  XOR U1390 ( .A(n832), .B(n907), .Z(n844) );
  XOR U1391 ( .A(n833), .B(n834), .Z(n907) );
  XOR U1392 ( .A(n839), .B(n908), .Z(n834) );
  XOR U1393 ( .A(n838), .B(n841), .Z(n908) );
  IV U1394 ( .A(n840), .Z(n841) );
  NAND U1395 ( .A(n909), .B(n910), .Z(n840) );
  OR U1396 ( .A(n911), .B(n912), .Z(n910) );
  OR U1397 ( .A(n913), .B(n914), .Z(n909) );
  NAND U1398 ( .A(n915), .B(n916), .Z(n838) );
  OR U1399 ( .A(n917), .B(n918), .Z(n916) );
  OR U1400 ( .A(n919), .B(n920), .Z(n915) );
  NOR U1401 ( .A(n921), .B(n922), .Z(n839) );
  ANDN U1402 ( .B(n923), .A(n924), .Z(n833) );
  IV U1403 ( .A(n925), .Z(n923) );
  XNOR U1404 ( .A(n826), .B(n926), .Z(n832) );
  XNOR U1405 ( .A(n825), .B(n827), .Z(n926) );
  NAND U1406 ( .A(n927), .B(n928), .Z(n827) );
  OR U1407 ( .A(n929), .B(n930), .Z(n928) );
  OR U1408 ( .A(n931), .B(n932), .Z(n927) );
  NAND U1409 ( .A(n933), .B(n934), .Z(n825) );
  OR U1410 ( .A(n935), .B(n936), .Z(n934) );
  OR U1411 ( .A(n937), .B(n938), .Z(n933) );
  ANDN U1412 ( .B(n939), .A(n940), .Z(n826) );
  IV U1413 ( .A(n941), .Z(n939) );
  XNOR U1414 ( .A(n906), .B(n905), .Z(N2744) );
  XOR U1415 ( .A(n925), .B(n924), .Z(n905) );
  XNOR U1416 ( .A(n940), .B(n941), .Z(n924) );
  XNOR U1417 ( .A(n935), .B(n936), .Z(n941) );
  XNOR U1418 ( .A(n937), .B(n938), .Z(n936) );
  XNOR U1419 ( .A(y[421]), .B(x[421]), .Z(n938) );
  XNOR U1420 ( .A(y[422]), .B(x[422]), .Z(n937) );
  XNOR U1421 ( .A(y[420]), .B(x[420]), .Z(n935) );
  XNOR U1422 ( .A(n929), .B(n930), .Z(n940) );
  XNOR U1423 ( .A(y[417]), .B(x[417]), .Z(n930) );
  XNOR U1424 ( .A(n931), .B(n932), .Z(n929) );
  XNOR U1425 ( .A(y[418]), .B(x[418]), .Z(n932) );
  XNOR U1426 ( .A(y[419]), .B(x[419]), .Z(n931) );
  XNOR U1427 ( .A(n922), .B(n921), .Z(n925) );
  XNOR U1428 ( .A(n917), .B(n918), .Z(n921) );
  XNOR U1429 ( .A(y[414]), .B(x[414]), .Z(n918) );
  XNOR U1430 ( .A(n919), .B(n920), .Z(n917) );
  XNOR U1431 ( .A(y[415]), .B(x[415]), .Z(n920) );
  XNOR U1432 ( .A(y[416]), .B(x[416]), .Z(n919) );
  XNOR U1433 ( .A(n911), .B(n912), .Z(n922) );
  XNOR U1434 ( .A(y[411]), .B(x[411]), .Z(n912) );
  XNOR U1435 ( .A(n913), .B(n914), .Z(n911) );
  XNOR U1436 ( .A(y[412]), .B(x[412]), .Z(n914) );
  XNOR U1437 ( .A(y[413]), .B(x[413]), .Z(n913) );
  XOR U1438 ( .A(n887), .B(n888), .Z(n906) );
  XNOR U1439 ( .A(n903), .B(n904), .Z(n888) );
  XNOR U1440 ( .A(n898), .B(n899), .Z(n904) );
  XNOR U1441 ( .A(n900), .B(n901), .Z(n899) );
  XNOR U1442 ( .A(y[409]), .B(x[409]), .Z(n901) );
  XNOR U1443 ( .A(y[410]), .B(x[410]), .Z(n900) );
  XNOR U1444 ( .A(y[408]), .B(x[408]), .Z(n898) );
  XNOR U1445 ( .A(n892), .B(n893), .Z(n903) );
  XNOR U1446 ( .A(y[405]), .B(x[405]), .Z(n893) );
  XNOR U1447 ( .A(n894), .B(n895), .Z(n892) );
  XNOR U1448 ( .A(y[406]), .B(x[406]), .Z(n895) );
  XNOR U1449 ( .A(y[407]), .B(x[407]), .Z(n894) );
  XOR U1450 ( .A(n886), .B(n885), .Z(n887) );
  XNOR U1451 ( .A(n881), .B(n882), .Z(n885) );
  XNOR U1452 ( .A(y[402]), .B(x[402]), .Z(n882) );
  XNOR U1453 ( .A(n883), .B(n884), .Z(n881) );
  XNOR U1454 ( .A(y[403]), .B(x[403]), .Z(n884) );
  XNOR U1455 ( .A(y[404]), .B(x[404]), .Z(n883) );
  XNOR U1456 ( .A(n875), .B(n876), .Z(n886) );
  XNOR U1457 ( .A(y[399]), .B(x[399]), .Z(n876) );
  XNOR U1458 ( .A(n877), .B(n878), .Z(n875) );
  XNOR U1459 ( .A(y[400]), .B(x[400]), .Z(n878) );
  XNOR U1460 ( .A(y[401]), .B(x[401]), .Z(n877) );
  NAND U1461 ( .A(n942), .B(n943), .Z(N2739) );
  NANDN U1462 ( .A(n944), .B(n945), .Z(n943) );
  OR U1463 ( .A(n946), .B(n947), .Z(n945) );
  NAND U1464 ( .A(n946), .B(n947), .Z(n942) );
  XOR U1465 ( .A(n946), .B(n948), .Z(N2738) );
  XNOR U1466 ( .A(n944), .B(n947), .Z(n948) );
  AND U1467 ( .A(n949), .B(n950), .Z(n947) );
  NANDN U1468 ( .A(n951), .B(n952), .Z(n950) );
  NANDN U1469 ( .A(n953), .B(n954), .Z(n952) );
  NANDN U1470 ( .A(n954), .B(n953), .Z(n949) );
  NAND U1471 ( .A(n955), .B(n956), .Z(n944) );
  NANDN U1472 ( .A(n957), .B(n958), .Z(n956) );
  OR U1473 ( .A(n959), .B(n960), .Z(n958) );
  NAND U1474 ( .A(n960), .B(n959), .Z(n955) );
  AND U1475 ( .A(n961), .B(n962), .Z(n946) );
  NANDN U1476 ( .A(n963), .B(n964), .Z(n962) );
  NANDN U1477 ( .A(n965), .B(n966), .Z(n964) );
  NANDN U1478 ( .A(n966), .B(n965), .Z(n961) );
  XOR U1479 ( .A(n960), .B(n967), .Z(N2737) );
  XOR U1480 ( .A(n957), .B(n959), .Z(n967) );
  XNOR U1481 ( .A(n953), .B(n968), .Z(n959) );
  XNOR U1482 ( .A(n951), .B(n954), .Z(n968) );
  NAND U1483 ( .A(n969), .B(n970), .Z(n954) );
  NAND U1484 ( .A(n971), .B(n972), .Z(n970) );
  OR U1485 ( .A(n973), .B(n974), .Z(n971) );
  NANDN U1486 ( .A(n975), .B(n973), .Z(n969) );
  IV U1487 ( .A(n974), .Z(n975) );
  NAND U1488 ( .A(n976), .B(n977), .Z(n951) );
  NAND U1489 ( .A(n978), .B(n979), .Z(n977) );
  NANDN U1490 ( .A(n980), .B(n981), .Z(n978) );
  NANDN U1491 ( .A(n981), .B(n980), .Z(n976) );
  AND U1492 ( .A(n982), .B(n983), .Z(n953) );
  NAND U1493 ( .A(n984), .B(n985), .Z(n983) );
  OR U1494 ( .A(n986), .B(n987), .Z(n984) );
  NANDN U1495 ( .A(n988), .B(n986), .Z(n982) );
  NAND U1496 ( .A(n989), .B(n990), .Z(n957) );
  NANDN U1497 ( .A(n991), .B(n992), .Z(n990) );
  OR U1498 ( .A(n993), .B(n994), .Z(n992) );
  NANDN U1499 ( .A(n995), .B(n993), .Z(n989) );
  IV U1500 ( .A(n994), .Z(n995) );
  XNOR U1501 ( .A(n965), .B(n996), .Z(n960) );
  XNOR U1502 ( .A(n963), .B(n966), .Z(n996) );
  NAND U1503 ( .A(n997), .B(n998), .Z(n966) );
  NAND U1504 ( .A(n999), .B(n1000), .Z(n998) );
  OR U1505 ( .A(n1001), .B(n1002), .Z(n999) );
  NANDN U1506 ( .A(n1003), .B(n1001), .Z(n997) );
  IV U1507 ( .A(n1002), .Z(n1003) );
  NAND U1508 ( .A(n1004), .B(n1005), .Z(n963) );
  NAND U1509 ( .A(n1006), .B(n1007), .Z(n1005) );
  NANDN U1510 ( .A(n1008), .B(n1009), .Z(n1006) );
  NANDN U1511 ( .A(n1009), .B(n1008), .Z(n1004) );
  AND U1512 ( .A(n1010), .B(n1011), .Z(n965) );
  NAND U1513 ( .A(n1012), .B(n1013), .Z(n1011) );
  OR U1514 ( .A(n1014), .B(n1015), .Z(n1012) );
  NANDN U1515 ( .A(n1016), .B(n1014), .Z(n1010) );
  XNOR U1516 ( .A(n991), .B(n1017), .Z(N2736) );
  XOR U1517 ( .A(n993), .B(n994), .Z(n1017) );
  XNOR U1518 ( .A(n1007), .B(n1018), .Z(n994) );
  XOR U1519 ( .A(n1008), .B(n1009), .Z(n1018) );
  XOR U1520 ( .A(n1014), .B(n1019), .Z(n1009) );
  XOR U1521 ( .A(n1013), .B(n1016), .Z(n1019) );
  IV U1522 ( .A(n1015), .Z(n1016) );
  NAND U1523 ( .A(n1020), .B(n1021), .Z(n1015) );
  OR U1524 ( .A(n1022), .B(n1023), .Z(n1021) );
  OR U1525 ( .A(n1024), .B(n1025), .Z(n1020) );
  NAND U1526 ( .A(n1026), .B(n1027), .Z(n1013) );
  OR U1527 ( .A(n1028), .B(n1029), .Z(n1027) );
  OR U1528 ( .A(n1030), .B(n1031), .Z(n1026) );
  NOR U1529 ( .A(n1032), .B(n1033), .Z(n1014) );
  ANDN U1530 ( .B(n1034), .A(n1035), .Z(n1008) );
  XNOR U1531 ( .A(n1001), .B(n1036), .Z(n1007) );
  XNOR U1532 ( .A(n1000), .B(n1002), .Z(n1036) );
  NAND U1533 ( .A(n1037), .B(n1038), .Z(n1002) );
  OR U1534 ( .A(n1039), .B(n1040), .Z(n1038) );
  OR U1535 ( .A(n1041), .B(n1042), .Z(n1037) );
  NAND U1536 ( .A(n1043), .B(n1044), .Z(n1000) );
  OR U1537 ( .A(n1045), .B(n1046), .Z(n1044) );
  OR U1538 ( .A(n1047), .B(n1048), .Z(n1043) );
  ANDN U1539 ( .B(n1049), .A(n1050), .Z(n1001) );
  IV U1540 ( .A(n1051), .Z(n1049) );
  ANDN U1541 ( .B(n1052), .A(n1053), .Z(n993) );
  XOR U1542 ( .A(n979), .B(n1054), .Z(n991) );
  XOR U1543 ( .A(n980), .B(n981), .Z(n1054) );
  XOR U1544 ( .A(n986), .B(n1055), .Z(n981) );
  XOR U1545 ( .A(n985), .B(n988), .Z(n1055) );
  IV U1546 ( .A(n987), .Z(n988) );
  NAND U1547 ( .A(n1056), .B(n1057), .Z(n987) );
  OR U1548 ( .A(n1058), .B(n1059), .Z(n1057) );
  OR U1549 ( .A(n1060), .B(n1061), .Z(n1056) );
  NAND U1550 ( .A(n1062), .B(n1063), .Z(n985) );
  OR U1551 ( .A(n1064), .B(n1065), .Z(n1063) );
  OR U1552 ( .A(n1066), .B(n1067), .Z(n1062) );
  NOR U1553 ( .A(n1068), .B(n1069), .Z(n986) );
  ANDN U1554 ( .B(n1070), .A(n1071), .Z(n980) );
  IV U1555 ( .A(n1072), .Z(n1070) );
  XNOR U1556 ( .A(n973), .B(n1073), .Z(n979) );
  XNOR U1557 ( .A(n972), .B(n974), .Z(n1073) );
  NAND U1558 ( .A(n1074), .B(n1075), .Z(n974) );
  OR U1559 ( .A(n1076), .B(n1077), .Z(n1075) );
  OR U1560 ( .A(n1078), .B(n1079), .Z(n1074) );
  NAND U1561 ( .A(n1080), .B(n1081), .Z(n972) );
  OR U1562 ( .A(n1082), .B(n1083), .Z(n1081) );
  OR U1563 ( .A(n1084), .B(n1085), .Z(n1080) );
  ANDN U1564 ( .B(n1086), .A(n1087), .Z(n973) );
  IV U1565 ( .A(n1088), .Z(n1086) );
  XNOR U1566 ( .A(n1053), .B(n1052), .Z(N2735) );
  XOR U1567 ( .A(n1072), .B(n1071), .Z(n1052) );
  XNOR U1568 ( .A(n1087), .B(n1088), .Z(n1071) );
  XNOR U1569 ( .A(n1082), .B(n1083), .Z(n1088) );
  XNOR U1570 ( .A(n1084), .B(n1085), .Z(n1083) );
  XNOR U1571 ( .A(y[397]), .B(x[397]), .Z(n1085) );
  XNOR U1572 ( .A(y[398]), .B(x[398]), .Z(n1084) );
  XNOR U1573 ( .A(y[396]), .B(x[396]), .Z(n1082) );
  XNOR U1574 ( .A(n1076), .B(n1077), .Z(n1087) );
  XNOR U1575 ( .A(y[393]), .B(x[393]), .Z(n1077) );
  XNOR U1576 ( .A(n1078), .B(n1079), .Z(n1076) );
  XNOR U1577 ( .A(y[394]), .B(x[394]), .Z(n1079) );
  XNOR U1578 ( .A(y[395]), .B(x[395]), .Z(n1078) );
  XNOR U1579 ( .A(n1069), .B(n1068), .Z(n1072) );
  XNOR U1580 ( .A(n1064), .B(n1065), .Z(n1068) );
  XNOR U1581 ( .A(y[390]), .B(x[390]), .Z(n1065) );
  XNOR U1582 ( .A(n1066), .B(n1067), .Z(n1064) );
  XNOR U1583 ( .A(y[391]), .B(x[391]), .Z(n1067) );
  XNOR U1584 ( .A(y[392]), .B(x[392]), .Z(n1066) );
  XNOR U1585 ( .A(n1058), .B(n1059), .Z(n1069) );
  XNOR U1586 ( .A(y[387]), .B(x[387]), .Z(n1059) );
  XNOR U1587 ( .A(n1060), .B(n1061), .Z(n1058) );
  XNOR U1588 ( .A(y[388]), .B(x[388]), .Z(n1061) );
  XNOR U1589 ( .A(y[389]), .B(x[389]), .Z(n1060) );
  XOR U1590 ( .A(n1034), .B(n1035), .Z(n1053) );
  XNOR U1591 ( .A(n1050), .B(n1051), .Z(n1035) );
  XNOR U1592 ( .A(n1045), .B(n1046), .Z(n1051) );
  XNOR U1593 ( .A(n1047), .B(n1048), .Z(n1046) );
  XNOR U1594 ( .A(y[385]), .B(x[385]), .Z(n1048) );
  XNOR U1595 ( .A(y[386]), .B(x[386]), .Z(n1047) );
  XNOR U1596 ( .A(y[384]), .B(x[384]), .Z(n1045) );
  XNOR U1597 ( .A(n1039), .B(n1040), .Z(n1050) );
  XNOR U1598 ( .A(y[381]), .B(x[381]), .Z(n1040) );
  XNOR U1599 ( .A(n1041), .B(n1042), .Z(n1039) );
  XNOR U1600 ( .A(y[382]), .B(x[382]), .Z(n1042) );
  XNOR U1601 ( .A(y[383]), .B(x[383]), .Z(n1041) );
  XOR U1602 ( .A(n1033), .B(n1032), .Z(n1034) );
  XNOR U1603 ( .A(n1028), .B(n1029), .Z(n1032) );
  XNOR U1604 ( .A(y[378]), .B(x[378]), .Z(n1029) );
  XNOR U1605 ( .A(n1030), .B(n1031), .Z(n1028) );
  XNOR U1606 ( .A(y[379]), .B(x[379]), .Z(n1031) );
  XNOR U1607 ( .A(y[380]), .B(x[380]), .Z(n1030) );
  XNOR U1608 ( .A(n1022), .B(n1023), .Z(n1033) );
  XNOR U1609 ( .A(y[375]), .B(x[375]), .Z(n1023) );
  XNOR U1610 ( .A(n1024), .B(n1025), .Z(n1022) );
  XNOR U1611 ( .A(y[376]), .B(x[376]), .Z(n1025) );
  XNOR U1612 ( .A(y[377]), .B(x[377]), .Z(n1024) );
  NAND U1613 ( .A(n1089), .B(n1090), .Z(N2730) );
  NANDN U1614 ( .A(n1091), .B(n1092), .Z(n1090) );
  OR U1615 ( .A(n1093), .B(n1094), .Z(n1092) );
  NAND U1616 ( .A(n1093), .B(n1094), .Z(n1089) );
  XOR U1617 ( .A(n1093), .B(n1095), .Z(N2729) );
  XNOR U1618 ( .A(n1091), .B(n1094), .Z(n1095) );
  AND U1619 ( .A(n1096), .B(n1097), .Z(n1094) );
  NANDN U1620 ( .A(n1098), .B(n1099), .Z(n1097) );
  NANDN U1621 ( .A(n1100), .B(n1101), .Z(n1099) );
  NANDN U1622 ( .A(n1101), .B(n1100), .Z(n1096) );
  NAND U1623 ( .A(n1102), .B(n1103), .Z(n1091) );
  NANDN U1624 ( .A(n1104), .B(n1105), .Z(n1103) );
  OR U1625 ( .A(n1106), .B(n1107), .Z(n1105) );
  NAND U1626 ( .A(n1107), .B(n1106), .Z(n1102) );
  AND U1627 ( .A(n1108), .B(n1109), .Z(n1093) );
  NANDN U1628 ( .A(n1110), .B(n1111), .Z(n1109) );
  NANDN U1629 ( .A(n1112), .B(n1113), .Z(n1111) );
  NANDN U1630 ( .A(n1113), .B(n1112), .Z(n1108) );
  XOR U1631 ( .A(n1107), .B(n1114), .Z(N2728) );
  XOR U1632 ( .A(n1104), .B(n1106), .Z(n1114) );
  XNOR U1633 ( .A(n1100), .B(n1115), .Z(n1106) );
  XNOR U1634 ( .A(n1098), .B(n1101), .Z(n1115) );
  NAND U1635 ( .A(n1116), .B(n1117), .Z(n1101) );
  NAND U1636 ( .A(n1118), .B(n1119), .Z(n1117) );
  OR U1637 ( .A(n1120), .B(n1121), .Z(n1118) );
  NANDN U1638 ( .A(n1122), .B(n1120), .Z(n1116) );
  IV U1639 ( .A(n1121), .Z(n1122) );
  NAND U1640 ( .A(n1123), .B(n1124), .Z(n1098) );
  NAND U1641 ( .A(n1125), .B(n1126), .Z(n1124) );
  NANDN U1642 ( .A(n1127), .B(n1128), .Z(n1125) );
  NANDN U1643 ( .A(n1128), .B(n1127), .Z(n1123) );
  AND U1644 ( .A(n1129), .B(n1130), .Z(n1100) );
  NAND U1645 ( .A(n1131), .B(n1132), .Z(n1130) );
  OR U1646 ( .A(n1133), .B(n1134), .Z(n1131) );
  NANDN U1647 ( .A(n1135), .B(n1133), .Z(n1129) );
  NAND U1648 ( .A(n1136), .B(n1137), .Z(n1104) );
  NANDN U1649 ( .A(n1138), .B(n1139), .Z(n1137) );
  OR U1650 ( .A(n1140), .B(n1141), .Z(n1139) );
  NANDN U1651 ( .A(n1142), .B(n1140), .Z(n1136) );
  IV U1652 ( .A(n1141), .Z(n1142) );
  XNOR U1653 ( .A(n1112), .B(n1143), .Z(n1107) );
  XNOR U1654 ( .A(n1110), .B(n1113), .Z(n1143) );
  NAND U1655 ( .A(n1144), .B(n1145), .Z(n1113) );
  NAND U1656 ( .A(n1146), .B(n1147), .Z(n1145) );
  OR U1657 ( .A(n1148), .B(n1149), .Z(n1146) );
  NANDN U1658 ( .A(n1150), .B(n1148), .Z(n1144) );
  IV U1659 ( .A(n1149), .Z(n1150) );
  NAND U1660 ( .A(n1151), .B(n1152), .Z(n1110) );
  NAND U1661 ( .A(n1153), .B(n1154), .Z(n1152) );
  NANDN U1662 ( .A(n1155), .B(n1156), .Z(n1153) );
  NANDN U1663 ( .A(n1156), .B(n1155), .Z(n1151) );
  AND U1664 ( .A(n1157), .B(n1158), .Z(n1112) );
  NAND U1665 ( .A(n1159), .B(n1160), .Z(n1158) );
  OR U1666 ( .A(n1161), .B(n1162), .Z(n1159) );
  NANDN U1667 ( .A(n1163), .B(n1161), .Z(n1157) );
  XNOR U1668 ( .A(n1138), .B(n1164), .Z(N2727) );
  XOR U1669 ( .A(n1140), .B(n1141), .Z(n1164) );
  XNOR U1670 ( .A(n1154), .B(n1165), .Z(n1141) );
  XOR U1671 ( .A(n1155), .B(n1156), .Z(n1165) );
  XOR U1672 ( .A(n1161), .B(n1166), .Z(n1156) );
  XOR U1673 ( .A(n1160), .B(n1163), .Z(n1166) );
  IV U1674 ( .A(n1162), .Z(n1163) );
  NAND U1675 ( .A(n1167), .B(n1168), .Z(n1162) );
  OR U1676 ( .A(n1169), .B(n1170), .Z(n1168) );
  OR U1677 ( .A(n1171), .B(n1172), .Z(n1167) );
  NAND U1678 ( .A(n1173), .B(n1174), .Z(n1160) );
  OR U1679 ( .A(n1175), .B(n1176), .Z(n1174) );
  OR U1680 ( .A(n1177), .B(n1178), .Z(n1173) );
  NOR U1681 ( .A(n1179), .B(n1180), .Z(n1161) );
  ANDN U1682 ( .B(n1181), .A(n1182), .Z(n1155) );
  XNOR U1683 ( .A(n1148), .B(n1183), .Z(n1154) );
  XNOR U1684 ( .A(n1147), .B(n1149), .Z(n1183) );
  NAND U1685 ( .A(n1184), .B(n1185), .Z(n1149) );
  OR U1686 ( .A(n1186), .B(n1187), .Z(n1185) );
  OR U1687 ( .A(n1188), .B(n1189), .Z(n1184) );
  NAND U1688 ( .A(n1190), .B(n1191), .Z(n1147) );
  OR U1689 ( .A(n1192), .B(n1193), .Z(n1191) );
  OR U1690 ( .A(n1194), .B(n1195), .Z(n1190) );
  ANDN U1691 ( .B(n1196), .A(n1197), .Z(n1148) );
  IV U1692 ( .A(n1198), .Z(n1196) );
  ANDN U1693 ( .B(n1199), .A(n1200), .Z(n1140) );
  XOR U1694 ( .A(n1126), .B(n1201), .Z(n1138) );
  XOR U1695 ( .A(n1127), .B(n1128), .Z(n1201) );
  XOR U1696 ( .A(n1133), .B(n1202), .Z(n1128) );
  XOR U1697 ( .A(n1132), .B(n1135), .Z(n1202) );
  IV U1698 ( .A(n1134), .Z(n1135) );
  NAND U1699 ( .A(n1203), .B(n1204), .Z(n1134) );
  OR U1700 ( .A(n1205), .B(n1206), .Z(n1204) );
  OR U1701 ( .A(n1207), .B(n1208), .Z(n1203) );
  NAND U1702 ( .A(n1209), .B(n1210), .Z(n1132) );
  OR U1703 ( .A(n1211), .B(n1212), .Z(n1210) );
  OR U1704 ( .A(n1213), .B(n1214), .Z(n1209) );
  NOR U1705 ( .A(n1215), .B(n1216), .Z(n1133) );
  ANDN U1706 ( .B(n1217), .A(n1218), .Z(n1127) );
  IV U1707 ( .A(n1219), .Z(n1217) );
  XNOR U1708 ( .A(n1120), .B(n1220), .Z(n1126) );
  XNOR U1709 ( .A(n1119), .B(n1121), .Z(n1220) );
  NAND U1710 ( .A(n1221), .B(n1222), .Z(n1121) );
  OR U1711 ( .A(n1223), .B(n1224), .Z(n1222) );
  OR U1712 ( .A(n1225), .B(n1226), .Z(n1221) );
  NAND U1713 ( .A(n1227), .B(n1228), .Z(n1119) );
  OR U1714 ( .A(n1229), .B(n1230), .Z(n1228) );
  OR U1715 ( .A(n1231), .B(n1232), .Z(n1227) );
  ANDN U1716 ( .B(n1233), .A(n1234), .Z(n1120) );
  IV U1717 ( .A(n1235), .Z(n1233) );
  XNOR U1718 ( .A(n1200), .B(n1199), .Z(N2726) );
  XOR U1719 ( .A(n1219), .B(n1218), .Z(n1199) );
  XNOR U1720 ( .A(n1234), .B(n1235), .Z(n1218) );
  XNOR U1721 ( .A(n1229), .B(n1230), .Z(n1235) );
  XNOR U1722 ( .A(n1231), .B(n1232), .Z(n1230) );
  XNOR U1723 ( .A(y[373]), .B(x[373]), .Z(n1232) );
  XNOR U1724 ( .A(y[374]), .B(x[374]), .Z(n1231) );
  XNOR U1725 ( .A(y[372]), .B(x[372]), .Z(n1229) );
  XNOR U1726 ( .A(n1223), .B(n1224), .Z(n1234) );
  XNOR U1727 ( .A(y[369]), .B(x[369]), .Z(n1224) );
  XNOR U1728 ( .A(n1225), .B(n1226), .Z(n1223) );
  XNOR U1729 ( .A(y[370]), .B(x[370]), .Z(n1226) );
  XNOR U1730 ( .A(y[371]), .B(x[371]), .Z(n1225) );
  XNOR U1731 ( .A(n1216), .B(n1215), .Z(n1219) );
  XNOR U1732 ( .A(n1211), .B(n1212), .Z(n1215) );
  XNOR U1733 ( .A(y[366]), .B(x[366]), .Z(n1212) );
  XNOR U1734 ( .A(n1213), .B(n1214), .Z(n1211) );
  XNOR U1735 ( .A(y[367]), .B(x[367]), .Z(n1214) );
  XNOR U1736 ( .A(y[368]), .B(x[368]), .Z(n1213) );
  XNOR U1737 ( .A(n1205), .B(n1206), .Z(n1216) );
  XNOR U1738 ( .A(y[363]), .B(x[363]), .Z(n1206) );
  XNOR U1739 ( .A(n1207), .B(n1208), .Z(n1205) );
  XNOR U1740 ( .A(y[364]), .B(x[364]), .Z(n1208) );
  XNOR U1741 ( .A(y[365]), .B(x[365]), .Z(n1207) );
  XOR U1742 ( .A(n1181), .B(n1182), .Z(n1200) );
  XNOR U1743 ( .A(n1197), .B(n1198), .Z(n1182) );
  XNOR U1744 ( .A(n1192), .B(n1193), .Z(n1198) );
  XNOR U1745 ( .A(n1194), .B(n1195), .Z(n1193) );
  XNOR U1746 ( .A(y[361]), .B(x[361]), .Z(n1195) );
  XNOR U1747 ( .A(y[362]), .B(x[362]), .Z(n1194) );
  XNOR U1748 ( .A(y[360]), .B(x[360]), .Z(n1192) );
  XNOR U1749 ( .A(n1186), .B(n1187), .Z(n1197) );
  XNOR U1750 ( .A(y[357]), .B(x[357]), .Z(n1187) );
  XNOR U1751 ( .A(n1188), .B(n1189), .Z(n1186) );
  XNOR U1752 ( .A(y[358]), .B(x[358]), .Z(n1189) );
  XNOR U1753 ( .A(y[359]), .B(x[359]), .Z(n1188) );
  XOR U1754 ( .A(n1180), .B(n1179), .Z(n1181) );
  XNOR U1755 ( .A(n1175), .B(n1176), .Z(n1179) );
  XNOR U1756 ( .A(y[354]), .B(x[354]), .Z(n1176) );
  XNOR U1757 ( .A(n1177), .B(n1178), .Z(n1175) );
  XNOR U1758 ( .A(y[355]), .B(x[355]), .Z(n1178) );
  XNOR U1759 ( .A(y[356]), .B(x[356]), .Z(n1177) );
  XNOR U1760 ( .A(n1169), .B(n1170), .Z(n1180) );
  XNOR U1761 ( .A(y[351]), .B(x[351]), .Z(n1170) );
  XNOR U1762 ( .A(n1171), .B(n1172), .Z(n1169) );
  XNOR U1763 ( .A(y[352]), .B(x[352]), .Z(n1172) );
  XNOR U1764 ( .A(y[353]), .B(x[353]), .Z(n1171) );
  NAND U1765 ( .A(n1236), .B(n1237), .Z(N2721) );
  NANDN U1766 ( .A(n1238), .B(n1239), .Z(n1237) );
  OR U1767 ( .A(n1240), .B(n1241), .Z(n1239) );
  NAND U1768 ( .A(n1240), .B(n1241), .Z(n1236) );
  XOR U1769 ( .A(n1240), .B(n1242), .Z(N2720) );
  XNOR U1770 ( .A(n1238), .B(n1241), .Z(n1242) );
  AND U1771 ( .A(n1243), .B(n1244), .Z(n1241) );
  NANDN U1772 ( .A(n1245), .B(n1246), .Z(n1244) );
  NANDN U1773 ( .A(n1247), .B(n1248), .Z(n1246) );
  NANDN U1774 ( .A(n1248), .B(n1247), .Z(n1243) );
  NAND U1775 ( .A(n1249), .B(n1250), .Z(n1238) );
  NANDN U1776 ( .A(n1251), .B(n1252), .Z(n1250) );
  OR U1777 ( .A(n1253), .B(n1254), .Z(n1252) );
  NAND U1778 ( .A(n1254), .B(n1253), .Z(n1249) );
  AND U1779 ( .A(n1255), .B(n1256), .Z(n1240) );
  NANDN U1780 ( .A(n1257), .B(n1258), .Z(n1256) );
  NANDN U1781 ( .A(n1259), .B(n1260), .Z(n1258) );
  NANDN U1782 ( .A(n1260), .B(n1259), .Z(n1255) );
  XOR U1783 ( .A(n1254), .B(n1261), .Z(N2719) );
  XOR U1784 ( .A(n1251), .B(n1253), .Z(n1261) );
  XNOR U1785 ( .A(n1247), .B(n1262), .Z(n1253) );
  XNOR U1786 ( .A(n1245), .B(n1248), .Z(n1262) );
  NAND U1787 ( .A(n1263), .B(n1264), .Z(n1248) );
  NAND U1788 ( .A(n1265), .B(n1266), .Z(n1264) );
  OR U1789 ( .A(n1267), .B(n1268), .Z(n1265) );
  NANDN U1790 ( .A(n1269), .B(n1267), .Z(n1263) );
  IV U1791 ( .A(n1268), .Z(n1269) );
  NAND U1792 ( .A(n1270), .B(n1271), .Z(n1245) );
  NAND U1793 ( .A(n1272), .B(n1273), .Z(n1271) );
  NANDN U1794 ( .A(n1274), .B(n1275), .Z(n1272) );
  NANDN U1795 ( .A(n1275), .B(n1274), .Z(n1270) );
  AND U1796 ( .A(n1276), .B(n1277), .Z(n1247) );
  NAND U1797 ( .A(n1278), .B(n1279), .Z(n1277) );
  OR U1798 ( .A(n1280), .B(n1281), .Z(n1278) );
  NANDN U1799 ( .A(n1282), .B(n1280), .Z(n1276) );
  NAND U1800 ( .A(n1283), .B(n1284), .Z(n1251) );
  NANDN U1801 ( .A(n1285), .B(n1286), .Z(n1284) );
  OR U1802 ( .A(n1287), .B(n1288), .Z(n1286) );
  NANDN U1803 ( .A(n1289), .B(n1287), .Z(n1283) );
  IV U1804 ( .A(n1288), .Z(n1289) );
  XNOR U1805 ( .A(n1259), .B(n1290), .Z(n1254) );
  XNOR U1806 ( .A(n1257), .B(n1260), .Z(n1290) );
  NAND U1807 ( .A(n1291), .B(n1292), .Z(n1260) );
  NAND U1808 ( .A(n1293), .B(n1294), .Z(n1292) );
  OR U1809 ( .A(n1295), .B(n1296), .Z(n1293) );
  NANDN U1810 ( .A(n1297), .B(n1295), .Z(n1291) );
  IV U1811 ( .A(n1296), .Z(n1297) );
  NAND U1812 ( .A(n1298), .B(n1299), .Z(n1257) );
  NAND U1813 ( .A(n1300), .B(n1301), .Z(n1299) );
  NANDN U1814 ( .A(n1302), .B(n1303), .Z(n1300) );
  NANDN U1815 ( .A(n1303), .B(n1302), .Z(n1298) );
  AND U1816 ( .A(n1304), .B(n1305), .Z(n1259) );
  NAND U1817 ( .A(n1306), .B(n1307), .Z(n1305) );
  OR U1818 ( .A(n1308), .B(n1309), .Z(n1306) );
  NANDN U1819 ( .A(n1310), .B(n1308), .Z(n1304) );
  XNOR U1820 ( .A(n1285), .B(n1311), .Z(N2718) );
  XOR U1821 ( .A(n1287), .B(n1288), .Z(n1311) );
  XNOR U1822 ( .A(n1301), .B(n1312), .Z(n1288) );
  XOR U1823 ( .A(n1302), .B(n1303), .Z(n1312) );
  XOR U1824 ( .A(n1308), .B(n1313), .Z(n1303) );
  XOR U1825 ( .A(n1307), .B(n1310), .Z(n1313) );
  IV U1826 ( .A(n1309), .Z(n1310) );
  NAND U1827 ( .A(n1314), .B(n1315), .Z(n1309) );
  OR U1828 ( .A(n1316), .B(n1317), .Z(n1315) );
  OR U1829 ( .A(n1318), .B(n1319), .Z(n1314) );
  NAND U1830 ( .A(n1320), .B(n1321), .Z(n1307) );
  OR U1831 ( .A(n1322), .B(n1323), .Z(n1321) );
  OR U1832 ( .A(n1324), .B(n1325), .Z(n1320) );
  NOR U1833 ( .A(n1326), .B(n1327), .Z(n1308) );
  ANDN U1834 ( .B(n1328), .A(n1329), .Z(n1302) );
  XNOR U1835 ( .A(n1295), .B(n1330), .Z(n1301) );
  XNOR U1836 ( .A(n1294), .B(n1296), .Z(n1330) );
  NAND U1837 ( .A(n1331), .B(n1332), .Z(n1296) );
  OR U1838 ( .A(n1333), .B(n1334), .Z(n1332) );
  OR U1839 ( .A(n1335), .B(n1336), .Z(n1331) );
  NAND U1840 ( .A(n1337), .B(n1338), .Z(n1294) );
  OR U1841 ( .A(n1339), .B(n1340), .Z(n1338) );
  OR U1842 ( .A(n1341), .B(n1342), .Z(n1337) );
  ANDN U1843 ( .B(n1343), .A(n1344), .Z(n1295) );
  IV U1844 ( .A(n1345), .Z(n1343) );
  ANDN U1845 ( .B(n1346), .A(n1347), .Z(n1287) );
  XOR U1846 ( .A(n1273), .B(n1348), .Z(n1285) );
  XOR U1847 ( .A(n1274), .B(n1275), .Z(n1348) );
  XOR U1848 ( .A(n1280), .B(n1349), .Z(n1275) );
  XOR U1849 ( .A(n1279), .B(n1282), .Z(n1349) );
  IV U1850 ( .A(n1281), .Z(n1282) );
  NAND U1851 ( .A(n1350), .B(n1351), .Z(n1281) );
  OR U1852 ( .A(n1352), .B(n1353), .Z(n1351) );
  OR U1853 ( .A(n1354), .B(n1355), .Z(n1350) );
  NAND U1854 ( .A(n1356), .B(n1357), .Z(n1279) );
  OR U1855 ( .A(n1358), .B(n1359), .Z(n1357) );
  OR U1856 ( .A(n1360), .B(n1361), .Z(n1356) );
  NOR U1857 ( .A(n1362), .B(n1363), .Z(n1280) );
  ANDN U1858 ( .B(n1364), .A(n1365), .Z(n1274) );
  IV U1859 ( .A(n1366), .Z(n1364) );
  XNOR U1860 ( .A(n1267), .B(n1367), .Z(n1273) );
  XNOR U1861 ( .A(n1266), .B(n1268), .Z(n1367) );
  NAND U1862 ( .A(n1368), .B(n1369), .Z(n1268) );
  OR U1863 ( .A(n1370), .B(n1371), .Z(n1369) );
  OR U1864 ( .A(n1372), .B(n1373), .Z(n1368) );
  NAND U1865 ( .A(n1374), .B(n1375), .Z(n1266) );
  OR U1866 ( .A(n1376), .B(n1377), .Z(n1375) );
  OR U1867 ( .A(n1378), .B(n1379), .Z(n1374) );
  ANDN U1868 ( .B(n1380), .A(n1381), .Z(n1267) );
  IV U1869 ( .A(n1382), .Z(n1380) );
  XNOR U1870 ( .A(n1347), .B(n1346), .Z(N2717) );
  XOR U1871 ( .A(n1366), .B(n1365), .Z(n1346) );
  XNOR U1872 ( .A(n1381), .B(n1382), .Z(n1365) );
  XNOR U1873 ( .A(n1376), .B(n1377), .Z(n1382) );
  XNOR U1874 ( .A(n1378), .B(n1379), .Z(n1377) );
  XNOR U1875 ( .A(y[349]), .B(x[349]), .Z(n1379) );
  XNOR U1876 ( .A(y[350]), .B(x[350]), .Z(n1378) );
  XNOR U1877 ( .A(y[348]), .B(x[348]), .Z(n1376) );
  XNOR U1878 ( .A(n1370), .B(n1371), .Z(n1381) );
  XNOR U1879 ( .A(y[345]), .B(x[345]), .Z(n1371) );
  XNOR U1880 ( .A(n1372), .B(n1373), .Z(n1370) );
  XNOR U1881 ( .A(y[346]), .B(x[346]), .Z(n1373) );
  XNOR U1882 ( .A(y[347]), .B(x[347]), .Z(n1372) );
  XNOR U1883 ( .A(n1363), .B(n1362), .Z(n1366) );
  XNOR U1884 ( .A(n1358), .B(n1359), .Z(n1362) );
  XNOR U1885 ( .A(y[342]), .B(x[342]), .Z(n1359) );
  XNOR U1886 ( .A(n1360), .B(n1361), .Z(n1358) );
  XNOR U1887 ( .A(y[343]), .B(x[343]), .Z(n1361) );
  XNOR U1888 ( .A(y[344]), .B(x[344]), .Z(n1360) );
  XNOR U1889 ( .A(n1352), .B(n1353), .Z(n1363) );
  XNOR U1890 ( .A(y[339]), .B(x[339]), .Z(n1353) );
  XNOR U1891 ( .A(n1354), .B(n1355), .Z(n1352) );
  XNOR U1892 ( .A(y[340]), .B(x[340]), .Z(n1355) );
  XNOR U1893 ( .A(y[341]), .B(x[341]), .Z(n1354) );
  XOR U1894 ( .A(n1328), .B(n1329), .Z(n1347) );
  XNOR U1895 ( .A(n1344), .B(n1345), .Z(n1329) );
  XNOR U1896 ( .A(n1339), .B(n1340), .Z(n1345) );
  XNOR U1897 ( .A(n1341), .B(n1342), .Z(n1340) );
  XNOR U1898 ( .A(y[337]), .B(x[337]), .Z(n1342) );
  XNOR U1899 ( .A(y[338]), .B(x[338]), .Z(n1341) );
  XNOR U1900 ( .A(y[336]), .B(x[336]), .Z(n1339) );
  XNOR U1901 ( .A(n1333), .B(n1334), .Z(n1344) );
  XNOR U1902 ( .A(y[333]), .B(x[333]), .Z(n1334) );
  XNOR U1903 ( .A(n1335), .B(n1336), .Z(n1333) );
  XNOR U1904 ( .A(y[334]), .B(x[334]), .Z(n1336) );
  XNOR U1905 ( .A(y[335]), .B(x[335]), .Z(n1335) );
  XOR U1906 ( .A(n1327), .B(n1326), .Z(n1328) );
  XNOR U1907 ( .A(n1322), .B(n1323), .Z(n1326) );
  XNOR U1908 ( .A(y[330]), .B(x[330]), .Z(n1323) );
  XNOR U1909 ( .A(n1324), .B(n1325), .Z(n1322) );
  XNOR U1910 ( .A(y[331]), .B(x[331]), .Z(n1325) );
  XNOR U1911 ( .A(y[332]), .B(x[332]), .Z(n1324) );
  XNOR U1912 ( .A(n1316), .B(n1317), .Z(n1327) );
  XNOR U1913 ( .A(y[327]), .B(x[327]), .Z(n1317) );
  XNOR U1914 ( .A(n1318), .B(n1319), .Z(n1316) );
  XNOR U1915 ( .A(y[328]), .B(x[328]), .Z(n1319) );
  XNOR U1916 ( .A(y[329]), .B(x[329]), .Z(n1318) );
  NAND U1917 ( .A(n1383), .B(n1384), .Z(N2712) );
  NANDN U1918 ( .A(n1385), .B(n1386), .Z(n1384) );
  OR U1919 ( .A(n1387), .B(n1388), .Z(n1386) );
  NAND U1920 ( .A(n1387), .B(n1388), .Z(n1383) );
  XOR U1921 ( .A(n1387), .B(n1389), .Z(N2711) );
  XNOR U1922 ( .A(n1385), .B(n1388), .Z(n1389) );
  AND U1923 ( .A(n1390), .B(n1391), .Z(n1388) );
  NANDN U1924 ( .A(n1392), .B(n1393), .Z(n1391) );
  NANDN U1925 ( .A(n1394), .B(n1395), .Z(n1393) );
  NANDN U1926 ( .A(n1395), .B(n1394), .Z(n1390) );
  NAND U1927 ( .A(n1396), .B(n1397), .Z(n1385) );
  NANDN U1928 ( .A(n1398), .B(n1399), .Z(n1397) );
  OR U1929 ( .A(n1400), .B(n1401), .Z(n1399) );
  NAND U1930 ( .A(n1401), .B(n1400), .Z(n1396) );
  AND U1931 ( .A(n1402), .B(n1403), .Z(n1387) );
  NANDN U1932 ( .A(n1404), .B(n1405), .Z(n1403) );
  NANDN U1933 ( .A(n1406), .B(n1407), .Z(n1405) );
  NANDN U1934 ( .A(n1407), .B(n1406), .Z(n1402) );
  XOR U1935 ( .A(n1401), .B(n1408), .Z(N2710) );
  XOR U1936 ( .A(n1398), .B(n1400), .Z(n1408) );
  XNOR U1937 ( .A(n1394), .B(n1409), .Z(n1400) );
  XNOR U1938 ( .A(n1392), .B(n1395), .Z(n1409) );
  NAND U1939 ( .A(n1410), .B(n1411), .Z(n1395) );
  NAND U1940 ( .A(n1412), .B(n1413), .Z(n1411) );
  OR U1941 ( .A(n1414), .B(n1415), .Z(n1412) );
  NANDN U1942 ( .A(n1416), .B(n1414), .Z(n1410) );
  IV U1943 ( .A(n1415), .Z(n1416) );
  NAND U1944 ( .A(n1417), .B(n1418), .Z(n1392) );
  NAND U1945 ( .A(n1419), .B(n1420), .Z(n1418) );
  NANDN U1946 ( .A(n1421), .B(n1422), .Z(n1419) );
  NANDN U1947 ( .A(n1422), .B(n1421), .Z(n1417) );
  AND U1948 ( .A(n1423), .B(n1424), .Z(n1394) );
  NAND U1949 ( .A(n1425), .B(n1426), .Z(n1424) );
  OR U1950 ( .A(n1427), .B(n1428), .Z(n1425) );
  NANDN U1951 ( .A(n1429), .B(n1427), .Z(n1423) );
  NAND U1952 ( .A(n1430), .B(n1431), .Z(n1398) );
  NANDN U1953 ( .A(n1432), .B(n1433), .Z(n1431) );
  OR U1954 ( .A(n1434), .B(n1435), .Z(n1433) );
  NANDN U1955 ( .A(n1436), .B(n1434), .Z(n1430) );
  IV U1956 ( .A(n1435), .Z(n1436) );
  XNOR U1957 ( .A(n1406), .B(n1437), .Z(n1401) );
  XNOR U1958 ( .A(n1404), .B(n1407), .Z(n1437) );
  NAND U1959 ( .A(n1438), .B(n1439), .Z(n1407) );
  NAND U1960 ( .A(n1440), .B(n1441), .Z(n1439) );
  OR U1961 ( .A(n1442), .B(n1443), .Z(n1440) );
  NANDN U1962 ( .A(n1444), .B(n1442), .Z(n1438) );
  IV U1963 ( .A(n1443), .Z(n1444) );
  NAND U1964 ( .A(n1445), .B(n1446), .Z(n1404) );
  NAND U1965 ( .A(n1447), .B(n1448), .Z(n1446) );
  NANDN U1966 ( .A(n1449), .B(n1450), .Z(n1447) );
  NANDN U1967 ( .A(n1450), .B(n1449), .Z(n1445) );
  AND U1968 ( .A(n1451), .B(n1452), .Z(n1406) );
  NAND U1969 ( .A(n1453), .B(n1454), .Z(n1452) );
  OR U1970 ( .A(n1455), .B(n1456), .Z(n1453) );
  NANDN U1971 ( .A(n1457), .B(n1455), .Z(n1451) );
  XNOR U1972 ( .A(n1432), .B(n1458), .Z(N2709) );
  XOR U1973 ( .A(n1434), .B(n1435), .Z(n1458) );
  XNOR U1974 ( .A(n1448), .B(n1459), .Z(n1435) );
  XOR U1975 ( .A(n1449), .B(n1450), .Z(n1459) );
  XOR U1976 ( .A(n1455), .B(n1460), .Z(n1450) );
  XOR U1977 ( .A(n1454), .B(n1457), .Z(n1460) );
  IV U1978 ( .A(n1456), .Z(n1457) );
  NAND U1979 ( .A(n1461), .B(n1462), .Z(n1456) );
  OR U1980 ( .A(n1463), .B(n1464), .Z(n1462) );
  OR U1981 ( .A(n1465), .B(n1466), .Z(n1461) );
  NAND U1982 ( .A(n1467), .B(n1468), .Z(n1454) );
  OR U1983 ( .A(n1469), .B(n1470), .Z(n1468) );
  OR U1984 ( .A(n1471), .B(n1472), .Z(n1467) );
  NOR U1985 ( .A(n1473), .B(n1474), .Z(n1455) );
  ANDN U1986 ( .B(n1475), .A(n1476), .Z(n1449) );
  XNOR U1987 ( .A(n1442), .B(n1477), .Z(n1448) );
  XNOR U1988 ( .A(n1441), .B(n1443), .Z(n1477) );
  NAND U1989 ( .A(n1478), .B(n1479), .Z(n1443) );
  OR U1990 ( .A(n1480), .B(n1481), .Z(n1479) );
  OR U1991 ( .A(n1482), .B(n1483), .Z(n1478) );
  NAND U1992 ( .A(n1484), .B(n1485), .Z(n1441) );
  OR U1993 ( .A(n1486), .B(n1487), .Z(n1485) );
  OR U1994 ( .A(n1488), .B(n1489), .Z(n1484) );
  ANDN U1995 ( .B(n1490), .A(n1491), .Z(n1442) );
  IV U1996 ( .A(n1492), .Z(n1490) );
  ANDN U1997 ( .B(n1493), .A(n1494), .Z(n1434) );
  XOR U1998 ( .A(n1420), .B(n1495), .Z(n1432) );
  XOR U1999 ( .A(n1421), .B(n1422), .Z(n1495) );
  XOR U2000 ( .A(n1427), .B(n1496), .Z(n1422) );
  XOR U2001 ( .A(n1426), .B(n1429), .Z(n1496) );
  IV U2002 ( .A(n1428), .Z(n1429) );
  NAND U2003 ( .A(n1497), .B(n1498), .Z(n1428) );
  OR U2004 ( .A(n1499), .B(n1500), .Z(n1498) );
  OR U2005 ( .A(n1501), .B(n1502), .Z(n1497) );
  NAND U2006 ( .A(n1503), .B(n1504), .Z(n1426) );
  OR U2007 ( .A(n1505), .B(n1506), .Z(n1504) );
  OR U2008 ( .A(n1507), .B(n1508), .Z(n1503) );
  NOR U2009 ( .A(n1509), .B(n1510), .Z(n1427) );
  ANDN U2010 ( .B(n1511), .A(n1512), .Z(n1421) );
  IV U2011 ( .A(n1513), .Z(n1511) );
  XNOR U2012 ( .A(n1414), .B(n1514), .Z(n1420) );
  XNOR U2013 ( .A(n1413), .B(n1415), .Z(n1514) );
  NAND U2014 ( .A(n1515), .B(n1516), .Z(n1415) );
  OR U2015 ( .A(n1517), .B(n1518), .Z(n1516) );
  OR U2016 ( .A(n1519), .B(n1520), .Z(n1515) );
  NAND U2017 ( .A(n1521), .B(n1522), .Z(n1413) );
  OR U2018 ( .A(n1523), .B(n1524), .Z(n1522) );
  OR U2019 ( .A(n1525), .B(n1526), .Z(n1521) );
  ANDN U2020 ( .B(n1527), .A(n1528), .Z(n1414) );
  IV U2021 ( .A(n1529), .Z(n1527) );
  XNOR U2022 ( .A(n1494), .B(n1493), .Z(N2708) );
  XOR U2023 ( .A(n1513), .B(n1512), .Z(n1493) );
  XNOR U2024 ( .A(n1528), .B(n1529), .Z(n1512) );
  XNOR U2025 ( .A(n1523), .B(n1524), .Z(n1529) );
  XNOR U2026 ( .A(n1525), .B(n1526), .Z(n1524) );
  XNOR U2027 ( .A(y[325]), .B(x[325]), .Z(n1526) );
  XNOR U2028 ( .A(y[326]), .B(x[326]), .Z(n1525) );
  XNOR U2029 ( .A(y[324]), .B(x[324]), .Z(n1523) );
  XNOR U2030 ( .A(n1517), .B(n1518), .Z(n1528) );
  XNOR U2031 ( .A(y[321]), .B(x[321]), .Z(n1518) );
  XNOR U2032 ( .A(n1519), .B(n1520), .Z(n1517) );
  XNOR U2033 ( .A(y[322]), .B(x[322]), .Z(n1520) );
  XNOR U2034 ( .A(y[323]), .B(x[323]), .Z(n1519) );
  XNOR U2035 ( .A(n1510), .B(n1509), .Z(n1513) );
  XNOR U2036 ( .A(n1505), .B(n1506), .Z(n1509) );
  XNOR U2037 ( .A(y[318]), .B(x[318]), .Z(n1506) );
  XNOR U2038 ( .A(n1507), .B(n1508), .Z(n1505) );
  XNOR U2039 ( .A(y[319]), .B(x[319]), .Z(n1508) );
  XNOR U2040 ( .A(y[320]), .B(x[320]), .Z(n1507) );
  XNOR U2041 ( .A(n1499), .B(n1500), .Z(n1510) );
  XNOR U2042 ( .A(y[315]), .B(x[315]), .Z(n1500) );
  XNOR U2043 ( .A(n1501), .B(n1502), .Z(n1499) );
  XNOR U2044 ( .A(y[316]), .B(x[316]), .Z(n1502) );
  XNOR U2045 ( .A(y[317]), .B(x[317]), .Z(n1501) );
  XOR U2046 ( .A(n1475), .B(n1476), .Z(n1494) );
  XNOR U2047 ( .A(n1491), .B(n1492), .Z(n1476) );
  XNOR U2048 ( .A(n1486), .B(n1487), .Z(n1492) );
  XNOR U2049 ( .A(n1488), .B(n1489), .Z(n1487) );
  XNOR U2050 ( .A(y[313]), .B(x[313]), .Z(n1489) );
  XNOR U2051 ( .A(y[314]), .B(x[314]), .Z(n1488) );
  XNOR U2052 ( .A(y[312]), .B(x[312]), .Z(n1486) );
  XNOR U2053 ( .A(n1480), .B(n1481), .Z(n1491) );
  XNOR U2054 ( .A(y[309]), .B(x[309]), .Z(n1481) );
  XNOR U2055 ( .A(n1482), .B(n1483), .Z(n1480) );
  XNOR U2056 ( .A(y[310]), .B(x[310]), .Z(n1483) );
  XNOR U2057 ( .A(y[311]), .B(x[311]), .Z(n1482) );
  XOR U2058 ( .A(n1474), .B(n1473), .Z(n1475) );
  XNOR U2059 ( .A(n1469), .B(n1470), .Z(n1473) );
  XNOR U2060 ( .A(y[306]), .B(x[306]), .Z(n1470) );
  XNOR U2061 ( .A(n1471), .B(n1472), .Z(n1469) );
  XNOR U2062 ( .A(y[307]), .B(x[307]), .Z(n1472) );
  XNOR U2063 ( .A(y[308]), .B(x[308]), .Z(n1471) );
  XNOR U2064 ( .A(n1463), .B(n1464), .Z(n1474) );
  XNOR U2065 ( .A(y[303]), .B(x[303]), .Z(n1464) );
  XNOR U2066 ( .A(n1465), .B(n1466), .Z(n1463) );
  XNOR U2067 ( .A(y[304]), .B(x[304]), .Z(n1466) );
  XNOR U2068 ( .A(y[305]), .B(x[305]), .Z(n1465) );
  NAND U2069 ( .A(n1530), .B(n1531), .Z(N2703) );
  NANDN U2070 ( .A(n1532), .B(n1533), .Z(n1531) );
  OR U2071 ( .A(n1534), .B(n1535), .Z(n1533) );
  NAND U2072 ( .A(n1534), .B(n1535), .Z(n1530) );
  XOR U2073 ( .A(n1534), .B(n1536), .Z(N2702) );
  XNOR U2074 ( .A(n1532), .B(n1535), .Z(n1536) );
  AND U2075 ( .A(n1537), .B(n1538), .Z(n1535) );
  NANDN U2076 ( .A(n1539), .B(n1540), .Z(n1538) );
  NANDN U2077 ( .A(n1541), .B(n1542), .Z(n1540) );
  NANDN U2078 ( .A(n1542), .B(n1541), .Z(n1537) );
  NAND U2079 ( .A(n1543), .B(n1544), .Z(n1532) );
  NANDN U2080 ( .A(n1545), .B(n1546), .Z(n1544) );
  OR U2081 ( .A(n1547), .B(n1548), .Z(n1546) );
  NAND U2082 ( .A(n1548), .B(n1547), .Z(n1543) );
  AND U2083 ( .A(n1549), .B(n1550), .Z(n1534) );
  NANDN U2084 ( .A(n1551), .B(n1552), .Z(n1550) );
  NANDN U2085 ( .A(n1553), .B(n1554), .Z(n1552) );
  NANDN U2086 ( .A(n1554), .B(n1553), .Z(n1549) );
  XOR U2087 ( .A(n1548), .B(n1555), .Z(N2701) );
  XOR U2088 ( .A(n1545), .B(n1547), .Z(n1555) );
  XNOR U2089 ( .A(n1541), .B(n1556), .Z(n1547) );
  XNOR U2090 ( .A(n1539), .B(n1542), .Z(n1556) );
  NAND U2091 ( .A(n1557), .B(n1558), .Z(n1542) );
  NAND U2092 ( .A(n1559), .B(n1560), .Z(n1558) );
  OR U2093 ( .A(n1561), .B(n1562), .Z(n1559) );
  NANDN U2094 ( .A(n1563), .B(n1561), .Z(n1557) );
  IV U2095 ( .A(n1562), .Z(n1563) );
  NAND U2096 ( .A(n1564), .B(n1565), .Z(n1539) );
  NAND U2097 ( .A(n1566), .B(n1567), .Z(n1565) );
  NANDN U2098 ( .A(n1568), .B(n1569), .Z(n1566) );
  NANDN U2099 ( .A(n1569), .B(n1568), .Z(n1564) );
  AND U2100 ( .A(n1570), .B(n1571), .Z(n1541) );
  NAND U2101 ( .A(n1572), .B(n1573), .Z(n1571) );
  OR U2102 ( .A(n1574), .B(n1575), .Z(n1572) );
  NANDN U2103 ( .A(n1576), .B(n1574), .Z(n1570) );
  NAND U2104 ( .A(n1577), .B(n1578), .Z(n1545) );
  NANDN U2105 ( .A(n1579), .B(n1580), .Z(n1578) );
  OR U2106 ( .A(n1581), .B(n1582), .Z(n1580) );
  NANDN U2107 ( .A(n1583), .B(n1581), .Z(n1577) );
  IV U2108 ( .A(n1582), .Z(n1583) );
  XNOR U2109 ( .A(n1553), .B(n1584), .Z(n1548) );
  XNOR U2110 ( .A(n1551), .B(n1554), .Z(n1584) );
  NAND U2111 ( .A(n1585), .B(n1586), .Z(n1554) );
  NAND U2112 ( .A(n1587), .B(n1588), .Z(n1586) );
  OR U2113 ( .A(n1589), .B(n1590), .Z(n1587) );
  NANDN U2114 ( .A(n1591), .B(n1589), .Z(n1585) );
  IV U2115 ( .A(n1590), .Z(n1591) );
  NAND U2116 ( .A(n1592), .B(n1593), .Z(n1551) );
  NAND U2117 ( .A(n1594), .B(n1595), .Z(n1593) );
  NANDN U2118 ( .A(n1596), .B(n1597), .Z(n1594) );
  NANDN U2119 ( .A(n1597), .B(n1596), .Z(n1592) );
  AND U2120 ( .A(n1598), .B(n1599), .Z(n1553) );
  NAND U2121 ( .A(n1600), .B(n1601), .Z(n1599) );
  OR U2122 ( .A(n1602), .B(n1603), .Z(n1600) );
  NANDN U2123 ( .A(n1604), .B(n1602), .Z(n1598) );
  XNOR U2124 ( .A(n1579), .B(n1605), .Z(N2700) );
  XOR U2125 ( .A(n1581), .B(n1582), .Z(n1605) );
  XNOR U2126 ( .A(n1595), .B(n1606), .Z(n1582) );
  XOR U2127 ( .A(n1596), .B(n1597), .Z(n1606) );
  XOR U2128 ( .A(n1602), .B(n1607), .Z(n1597) );
  XOR U2129 ( .A(n1601), .B(n1604), .Z(n1607) );
  IV U2130 ( .A(n1603), .Z(n1604) );
  NAND U2131 ( .A(n1608), .B(n1609), .Z(n1603) );
  OR U2132 ( .A(n1610), .B(n1611), .Z(n1609) );
  OR U2133 ( .A(n1612), .B(n1613), .Z(n1608) );
  NAND U2134 ( .A(n1614), .B(n1615), .Z(n1601) );
  OR U2135 ( .A(n1616), .B(n1617), .Z(n1615) );
  OR U2136 ( .A(n1618), .B(n1619), .Z(n1614) );
  NOR U2137 ( .A(n1620), .B(n1621), .Z(n1602) );
  ANDN U2138 ( .B(n1622), .A(n1623), .Z(n1596) );
  XNOR U2139 ( .A(n1589), .B(n1624), .Z(n1595) );
  XNOR U2140 ( .A(n1588), .B(n1590), .Z(n1624) );
  NAND U2141 ( .A(n1625), .B(n1626), .Z(n1590) );
  OR U2142 ( .A(n1627), .B(n1628), .Z(n1626) );
  OR U2143 ( .A(n1629), .B(n1630), .Z(n1625) );
  NAND U2144 ( .A(n1631), .B(n1632), .Z(n1588) );
  OR U2145 ( .A(n1633), .B(n1634), .Z(n1632) );
  OR U2146 ( .A(n1635), .B(n1636), .Z(n1631) );
  ANDN U2147 ( .B(n1637), .A(n1638), .Z(n1589) );
  IV U2148 ( .A(n1639), .Z(n1637) );
  ANDN U2149 ( .B(n1640), .A(n1641), .Z(n1581) );
  XOR U2150 ( .A(n1567), .B(n1642), .Z(n1579) );
  XOR U2151 ( .A(n1568), .B(n1569), .Z(n1642) );
  XOR U2152 ( .A(n1574), .B(n1643), .Z(n1569) );
  XOR U2153 ( .A(n1573), .B(n1576), .Z(n1643) );
  IV U2154 ( .A(n1575), .Z(n1576) );
  NAND U2155 ( .A(n1644), .B(n1645), .Z(n1575) );
  OR U2156 ( .A(n1646), .B(n1647), .Z(n1645) );
  OR U2157 ( .A(n1648), .B(n1649), .Z(n1644) );
  NAND U2158 ( .A(n1650), .B(n1651), .Z(n1573) );
  OR U2159 ( .A(n1652), .B(n1653), .Z(n1651) );
  OR U2160 ( .A(n1654), .B(n1655), .Z(n1650) );
  NOR U2161 ( .A(n1656), .B(n1657), .Z(n1574) );
  ANDN U2162 ( .B(n1658), .A(n1659), .Z(n1568) );
  IV U2163 ( .A(n1660), .Z(n1658) );
  XNOR U2164 ( .A(n1561), .B(n1661), .Z(n1567) );
  XNOR U2165 ( .A(n1560), .B(n1562), .Z(n1661) );
  NAND U2166 ( .A(n1662), .B(n1663), .Z(n1562) );
  OR U2167 ( .A(n1664), .B(n1665), .Z(n1663) );
  OR U2168 ( .A(n1666), .B(n1667), .Z(n1662) );
  NAND U2169 ( .A(n1668), .B(n1669), .Z(n1560) );
  OR U2170 ( .A(n1670), .B(n1671), .Z(n1669) );
  OR U2171 ( .A(n1672), .B(n1673), .Z(n1668) );
  ANDN U2172 ( .B(n1674), .A(n1675), .Z(n1561) );
  IV U2173 ( .A(n1676), .Z(n1674) );
  XNOR U2174 ( .A(n1641), .B(n1640), .Z(N2699) );
  XOR U2175 ( .A(n1660), .B(n1659), .Z(n1640) );
  XNOR U2176 ( .A(n1675), .B(n1676), .Z(n1659) );
  XNOR U2177 ( .A(n1670), .B(n1671), .Z(n1676) );
  XNOR U2178 ( .A(n1672), .B(n1673), .Z(n1671) );
  XNOR U2179 ( .A(y[301]), .B(x[301]), .Z(n1673) );
  XNOR U2180 ( .A(y[302]), .B(x[302]), .Z(n1672) );
  XNOR U2181 ( .A(y[300]), .B(x[300]), .Z(n1670) );
  XNOR U2182 ( .A(n1664), .B(n1665), .Z(n1675) );
  XNOR U2183 ( .A(y[297]), .B(x[297]), .Z(n1665) );
  XNOR U2184 ( .A(n1666), .B(n1667), .Z(n1664) );
  XNOR U2185 ( .A(y[298]), .B(x[298]), .Z(n1667) );
  XNOR U2186 ( .A(y[299]), .B(x[299]), .Z(n1666) );
  XNOR U2187 ( .A(n1657), .B(n1656), .Z(n1660) );
  XNOR U2188 ( .A(n1652), .B(n1653), .Z(n1656) );
  XNOR U2189 ( .A(y[294]), .B(x[294]), .Z(n1653) );
  XNOR U2190 ( .A(n1654), .B(n1655), .Z(n1652) );
  XNOR U2191 ( .A(y[295]), .B(x[295]), .Z(n1655) );
  XNOR U2192 ( .A(y[296]), .B(x[296]), .Z(n1654) );
  XNOR U2193 ( .A(n1646), .B(n1647), .Z(n1657) );
  XNOR U2194 ( .A(y[291]), .B(x[291]), .Z(n1647) );
  XNOR U2195 ( .A(n1648), .B(n1649), .Z(n1646) );
  XNOR U2196 ( .A(y[292]), .B(x[292]), .Z(n1649) );
  XNOR U2197 ( .A(y[293]), .B(x[293]), .Z(n1648) );
  XOR U2198 ( .A(n1622), .B(n1623), .Z(n1641) );
  XNOR U2199 ( .A(n1638), .B(n1639), .Z(n1623) );
  XNOR U2200 ( .A(n1633), .B(n1634), .Z(n1639) );
  XNOR U2201 ( .A(n1635), .B(n1636), .Z(n1634) );
  XNOR U2202 ( .A(y[289]), .B(x[289]), .Z(n1636) );
  XNOR U2203 ( .A(y[290]), .B(x[290]), .Z(n1635) );
  XNOR U2204 ( .A(y[288]), .B(x[288]), .Z(n1633) );
  XNOR U2205 ( .A(n1627), .B(n1628), .Z(n1638) );
  XNOR U2206 ( .A(y[285]), .B(x[285]), .Z(n1628) );
  XNOR U2207 ( .A(n1629), .B(n1630), .Z(n1627) );
  XNOR U2208 ( .A(y[286]), .B(x[286]), .Z(n1630) );
  XNOR U2209 ( .A(y[287]), .B(x[287]), .Z(n1629) );
  XOR U2210 ( .A(n1621), .B(n1620), .Z(n1622) );
  XNOR U2211 ( .A(n1616), .B(n1617), .Z(n1620) );
  XNOR U2212 ( .A(y[282]), .B(x[282]), .Z(n1617) );
  XNOR U2213 ( .A(n1618), .B(n1619), .Z(n1616) );
  XNOR U2214 ( .A(y[283]), .B(x[283]), .Z(n1619) );
  XNOR U2215 ( .A(y[284]), .B(x[284]), .Z(n1618) );
  XNOR U2216 ( .A(n1610), .B(n1611), .Z(n1621) );
  XNOR U2217 ( .A(y[279]), .B(x[279]), .Z(n1611) );
  XNOR U2218 ( .A(n1612), .B(n1613), .Z(n1610) );
  XNOR U2219 ( .A(y[280]), .B(x[280]), .Z(n1613) );
  XNOR U2220 ( .A(y[281]), .B(x[281]), .Z(n1612) );
  NAND U2221 ( .A(n1677), .B(n1678), .Z(N2694) );
  NANDN U2222 ( .A(n1679), .B(n1680), .Z(n1678) );
  OR U2223 ( .A(n1681), .B(n1682), .Z(n1680) );
  NAND U2224 ( .A(n1681), .B(n1682), .Z(n1677) );
  XOR U2225 ( .A(n1681), .B(n1683), .Z(N2693) );
  XNOR U2226 ( .A(n1679), .B(n1682), .Z(n1683) );
  AND U2227 ( .A(n1684), .B(n1685), .Z(n1682) );
  NANDN U2228 ( .A(n1686), .B(n1687), .Z(n1685) );
  NANDN U2229 ( .A(n1688), .B(n1689), .Z(n1687) );
  NANDN U2230 ( .A(n1689), .B(n1688), .Z(n1684) );
  NAND U2231 ( .A(n1690), .B(n1691), .Z(n1679) );
  NANDN U2232 ( .A(n1692), .B(n1693), .Z(n1691) );
  OR U2233 ( .A(n1694), .B(n1695), .Z(n1693) );
  NAND U2234 ( .A(n1695), .B(n1694), .Z(n1690) );
  AND U2235 ( .A(n1696), .B(n1697), .Z(n1681) );
  NANDN U2236 ( .A(n1698), .B(n1699), .Z(n1697) );
  NANDN U2237 ( .A(n1700), .B(n1701), .Z(n1699) );
  NANDN U2238 ( .A(n1701), .B(n1700), .Z(n1696) );
  XOR U2239 ( .A(n1695), .B(n1702), .Z(N2692) );
  XOR U2240 ( .A(n1692), .B(n1694), .Z(n1702) );
  XNOR U2241 ( .A(n1688), .B(n1703), .Z(n1694) );
  XNOR U2242 ( .A(n1686), .B(n1689), .Z(n1703) );
  NAND U2243 ( .A(n1704), .B(n1705), .Z(n1689) );
  NAND U2244 ( .A(n1706), .B(n1707), .Z(n1705) );
  OR U2245 ( .A(n1708), .B(n1709), .Z(n1706) );
  NANDN U2246 ( .A(n1710), .B(n1708), .Z(n1704) );
  IV U2247 ( .A(n1709), .Z(n1710) );
  NAND U2248 ( .A(n1711), .B(n1712), .Z(n1686) );
  NAND U2249 ( .A(n1713), .B(n1714), .Z(n1712) );
  NANDN U2250 ( .A(n1715), .B(n1716), .Z(n1713) );
  NANDN U2251 ( .A(n1716), .B(n1715), .Z(n1711) );
  AND U2252 ( .A(n1717), .B(n1718), .Z(n1688) );
  NAND U2253 ( .A(n1719), .B(n1720), .Z(n1718) );
  OR U2254 ( .A(n1721), .B(n1722), .Z(n1719) );
  NANDN U2255 ( .A(n1723), .B(n1721), .Z(n1717) );
  NAND U2256 ( .A(n1724), .B(n1725), .Z(n1692) );
  NANDN U2257 ( .A(n1726), .B(n1727), .Z(n1725) );
  OR U2258 ( .A(n1728), .B(n1729), .Z(n1727) );
  NANDN U2259 ( .A(n1730), .B(n1728), .Z(n1724) );
  IV U2260 ( .A(n1729), .Z(n1730) );
  XNOR U2261 ( .A(n1700), .B(n1731), .Z(n1695) );
  XNOR U2262 ( .A(n1698), .B(n1701), .Z(n1731) );
  NAND U2263 ( .A(n1732), .B(n1733), .Z(n1701) );
  NAND U2264 ( .A(n1734), .B(n1735), .Z(n1733) );
  OR U2265 ( .A(n1736), .B(n1737), .Z(n1734) );
  NANDN U2266 ( .A(n1738), .B(n1736), .Z(n1732) );
  IV U2267 ( .A(n1737), .Z(n1738) );
  NAND U2268 ( .A(n1739), .B(n1740), .Z(n1698) );
  NAND U2269 ( .A(n1741), .B(n1742), .Z(n1740) );
  NANDN U2270 ( .A(n1743), .B(n1744), .Z(n1741) );
  NANDN U2271 ( .A(n1744), .B(n1743), .Z(n1739) );
  AND U2272 ( .A(n1745), .B(n1746), .Z(n1700) );
  NAND U2273 ( .A(n1747), .B(n1748), .Z(n1746) );
  OR U2274 ( .A(n1749), .B(n1750), .Z(n1747) );
  NANDN U2275 ( .A(n1751), .B(n1749), .Z(n1745) );
  XNOR U2276 ( .A(n1726), .B(n1752), .Z(N2691) );
  XOR U2277 ( .A(n1728), .B(n1729), .Z(n1752) );
  XNOR U2278 ( .A(n1742), .B(n1753), .Z(n1729) );
  XOR U2279 ( .A(n1743), .B(n1744), .Z(n1753) );
  XOR U2280 ( .A(n1749), .B(n1754), .Z(n1744) );
  XOR U2281 ( .A(n1748), .B(n1751), .Z(n1754) );
  IV U2282 ( .A(n1750), .Z(n1751) );
  NAND U2283 ( .A(n1755), .B(n1756), .Z(n1750) );
  OR U2284 ( .A(n1757), .B(n1758), .Z(n1756) );
  OR U2285 ( .A(n1759), .B(n1760), .Z(n1755) );
  NAND U2286 ( .A(n1761), .B(n1762), .Z(n1748) );
  OR U2287 ( .A(n1763), .B(n1764), .Z(n1762) );
  OR U2288 ( .A(n1765), .B(n1766), .Z(n1761) );
  NOR U2289 ( .A(n1767), .B(n1768), .Z(n1749) );
  ANDN U2290 ( .B(n1769), .A(n1770), .Z(n1743) );
  XNOR U2291 ( .A(n1736), .B(n1771), .Z(n1742) );
  XNOR U2292 ( .A(n1735), .B(n1737), .Z(n1771) );
  NAND U2293 ( .A(n1772), .B(n1773), .Z(n1737) );
  OR U2294 ( .A(n1774), .B(n1775), .Z(n1773) );
  OR U2295 ( .A(n1776), .B(n1777), .Z(n1772) );
  NAND U2296 ( .A(n1778), .B(n1779), .Z(n1735) );
  OR U2297 ( .A(n1780), .B(n1781), .Z(n1779) );
  OR U2298 ( .A(n1782), .B(n1783), .Z(n1778) );
  ANDN U2299 ( .B(n1784), .A(n1785), .Z(n1736) );
  IV U2300 ( .A(n1786), .Z(n1784) );
  ANDN U2301 ( .B(n1787), .A(n1788), .Z(n1728) );
  XOR U2302 ( .A(n1714), .B(n1789), .Z(n1726) );
  XOR U2303 ( .A(n1715), .B(n1716), .Z(n1789) );
  XOR U2304 ( .A(n1721), .B(n1790), .Z(n1716) );
  XOR U2305 ( .A(n1720), .B(n1723), .Z(n1790) );
  IV U2306 ( .A(n1722), .Z(n1723) );
  NAND U2307 ( .A(n1791), .B(n1792), .Z(n1722) );
  OR U2308 ( .A(n1793), .B(n1794), .Z(n1792) );
  OR U2309 ( .A(n1795), .B(n1796), .Z(n1791) );
  NAND U2310 ( .A(n1797), .B(n1798), .Z(n1720) );
  OR U2311 ( .A(n1799), .B(n1800), .Z(n1798) );
  OR U2312 ( .A(n1801), .B(n1802), .Z(n1797) );
  NOR U2313 ( .A(n1803), .B(n1804), .Z(n1721) );
  ANDN U2314 ( .B(n1805), .A(n1806), .Z(n1715) );
  IV U2315 ( .A(n1807), .Z(n1805) );
  XNOR U2316 ( .A(n1708), .B(n1808), .Z(n1714) );
  XNOR U2317 ( .A(n1707), .B(n1709), .Z(n1808) );
  NAND U2318 ( .A(n1809), .B(n1810), .Z(n1709) );
  OR U2319 ( .A(n1811), .B(n1812), .Z(n1810) );
  OR U2320 ( .A(n1813), .B(n1814), .Z(n1809) );
  NAND U2321 ( .A(n1815), .B(n1816), .Z(n1707) );
  OR U2322 ( .A(n1817), .B(n1818), .Z(n1816) );
  OR U2323 ( .A(n1819), .B(n1820), .Z(n1815) );
  ANDN U2324 ( .B(n1821), .A(n1822), .Z(n1708) );
  IV U2325 ( .A(n1823), .Z(n1821) );
  XNOR U2326 ( .A(n1788), .B(n1787), .Z(N2690) );
  XOR U2327 ( .A(n1807), .B(n1806), .Z(n1787) );
  XNOR U2328 ( .A(n1822), .B(n1823), .Z(n1806) );
  XNOR U2329 ( .A(n1817), .B(n1818), .Z(n1823) );
  XNOR U2330 ( .A(n1819), .B(n1820), .Z(n1818) );
  XNOR U2331 ( .A(y[277]), .B(x[277]), .Z(n1820) );
  XNOR U2332 ( .A(y[278]), .B(x[278]), .Z(n1819) );
  XNOR U2333 ( .A(y[276]), .B(x[276]), .Z(n1817) );
  XNOR U2334 ( .A(n1811), .B(n1812), .Z(n1822) );
  XNOR U2335 ( .A(y[273]), .B(x[273]), .Z(n1812) );
  XNOR U2336 ( .A(n1813), .B(n1814), .Z(n1811) );
  XNOR U2337 ( .A(y[274]), .B(x[274]), .Z(n1814) );
  XNOR U2338 ( .A(y[275]), .B(x[275]), .Z(n1813) );
  XNOR U2339 ( .A(n1804), .B(n1803), .Z(n1807) );
  XNOR U2340 ( .A(n1799), .B(n1800), .Z(n1803) );
  XNOR U2341 ( .A(y[270]), .B(x[270]), .Z(n1800) );
  XNOR U2342 ( .A(n1801), .B(n1802), .Z(n1799) );
  XNOR U2343 ( .A(y[271]), .B(x[271]), .Z(n1802) );
  XNOR U2344 ( .A(y[272]), .B(x[272]), .Z(n1801) );
  XNOR U2345 ( .A(n1793), .B(n1794), .Z(n1804) );
  XNOR U2346 ( .A(y[267]), .B(x[267]), .Z(n1794) );
  XNOR U2347 ( .A(n1795), .B(n1796), .Z(n1793) );
  XNOR U2348 ( .A(y[268]), .B(x[268]), .Z(n1796) );
  XNOR U2349 ( .A(y[269]), .B(x[269]), .Z(n1795) );
  XOR U2350 ( .A(n1769), .B(n1770), .Z(n1788) );
  XNOR U2351 ( .A(n1785), .B(n1786), .Z(n1770) );
  XNOR U2352 ( .A(n1780), .B(n1781), .Z(n1786) );
  XNOR U2353 ( .A(n1782), .B(n1783), .Z(n1781) );
  XNOR U2354 ( .A(y[265]), .B(x[265]), .Z(n1783) );
  XNOR U2355 ( .A(y[266]), .B(x[266]), .Z(n1782) );
  XNOR U2356 ( .A(y[264]), .B(x[264]), .Z(n1780) );
  XNOR U2357 ( .A(n1774), .B(n1775), .Z(n1785) );
  XNOR U2358 ( .A(y[261]), .B(x[261]), .Z(n1775) );
  XNOR U2359 ( .A(n1776), .B(n1777), .Z(n1774) );
  XNOR U2360 ( .A(y[262]), .B(x[262]), .Z(n1777) );
  XNOR U2361 ( .A(y[263]), .B(x[263]), .Z(n1776) );
  XOR U2362 ( .A(n1768), .B(n1767), .Z(n1769) );
  XNOR U2363 ( .A(n1763), .B(n1764), .Z(n1767) );
  XNOR U2364 ( .A(y[258]), .B(x[258]), .Z(n1764) );
  XNOR U2365 ( .A(n1765), .B(n1766), .Z(n1763) );
  XNOR U2366 ( .A(y[259]), .B(x[259]), .Z(n1766) );
  XNOR U2367 ( .A(y[260]), .B(x[260]), .Z(n1765) );
  XNOR U2368 ( .A(n1757), .B(n1758), .Z(n1768) );
  XNOR U2369 ( .A(y[255]), .B(x[255]), .Z(n1758) );
  XNOR U2370 ( .A(n1759), .B(n1760), .Z(n1757) );
  XNOR U2371 ( .A(y[256]), .B(x[256]), .Z(n1760) );
  XNOR U2372 ( .A(y[257]), .B(x[257]), .Z(n1759) );
  NAND U2373 ( .A(n1824), .B(n1825), .Z(N2685) );
  NANDN U2374 ( .A(n1826), .B(n1827), .Z(n1825) );
  OR U2375 ( .A(n1828), .B(n1829), .Z(n1827) );
  NAND U2376 ( .A(n1828), .B(n1829), .Z(n1824) );
  XOR U2377 ( .A(n1828), .B(n1830), .Z(N2684) );
  XNOR U2378 ( .A(n1826), .B(n1829), .Z(n1830) );
  AND U2379 ( .A(n1831), .B(n1832), .Z(n1829) );
  NANDN U2380 ( .A(n1833), .B(n1834), .Z(n1832) );
  NANDN U2381 ( .A(n1835), .B(n1836), .Z(n1834) );
  NANDN U2382 ( .A(n1836), .B(n1835), .Z(n1831) );
  NAND U2383 ( .A(n1837), .B(n1838), .Z(n1826) );
  NANDN U2384 ( .A(n1839), .B(n1840), .Z(n1838) );
  OR U2385 ( .A(n1841), .B(n1842), .Z(n1840) );
  NAND U2386 ( .A(n1842), .B(n1841), .Z(n1837) );
  AND U2387 ( .A(n1843), .B(n1844), .Z(n1828) );
  NANDN U2388 ( .A(n1845), .B(n1846), .Z(n1844) );
  NANDN U2389 ( .A(n1847), .B(n1848), .Z(n1846) );
  NANDN U2390 ( .A(n1848), .B(n1847), .Z(n1843) );
  XOR U2391 ( .A(n1842), .B(n1849), .Z(N2683) );
  XOR U2392 ( .A(n1839), .B(n1841), .Z(n1849) );
  XNOR U2393 ( .A(n1835), .B(n1850), .Z(n1841) );
  XNOR U2394 ( .A(n1833), .B(n1836), .Z(n1850) );
  NAND U2395 ( .A(n1851), .B(n1852), .Z(n1836) );
  NAND U2396 ( .A(n1853), .B(n1854), .Z(n1852) );
  OR U2397 ( .A(n1855), .B(n1856), .Z(n1853) );
  NANDN U2398 ( .A(n1857), .B(n1855), .Z(n1851) );
  IV U2399 ( .A(n1856), .Z(n1857) );
  NAND U2400 ( .A(n1858), .B(n1859), .Z(n1833) );
  NAND U2401 ( .A(n1860), .B(n1861), .Z(n1859) );
  NANDN U2402 ( .A(n1862), .B(n1863), .Z(n1860) );
  NANDN U2403 ( .A(n1863), .B(n1862), .Z(n1858) );
  AND U2404 ( .A(n1864), .B(n1865), .Z(n1835) );
  NAND U2405 ( .A(n1866), .B(n1867), .Z(n1865) );
  OR U2406 ( .A(n1868), .B(n1869), .Z(n1866) );
  NANDN U2407 ( .A(n1870), .B(n1868), .Z(n1864) );
  NAND U2408 ( .A(n1871), .B(n1872), .Z(n1839) );
  NANDN U2409 ( .A(n1873), .B(n1874), .Z(n1872) );
  OR U2410 ( .A(n1875), .B(n1876), .Z(n1874) );
  NANDN U2411 ( .A(n1877), .B(n1875), .Z(n1871) );
  IV U2412 ( .A(n1876), .Z(n1877) );
  XNOR U2413 ( .A(n1847), .B(n1878), .Z(n1842) );
  XNOR U2414 ( .A(n1845), .B(n1848), .Z(n1878) );
  NAND U2415 ( .A(n1879), .B(n1880), .Z(n1848) );
  NAND U2416 ( .A(n1881), .B(n1882), .Z(n1880) );
  OR U2417 ( .A(n1883), .B(n1884), .Z(n1881) );
  NANDN U2418 ( .A(n1885), .B(n1883), .Z(n1879) );
  IV U2419 ( .A(n1884), .Z(n1885) );
  NAND U2420 ( .A(n1886), .B(n1887), .Z(n1845) );
  NAND U2421 ( .A(n1888), .B(n1889), .Z(n1887) );
  NANDN U2422 ( .A(n1890), .B(n1891), .Z(n1888) );
  NANDN U2423 ( .A(n1891), .B(n1890), .Z(n1886) );
  AND U2424 ( .A(n1892), .B(n1893), .Z(n1847) );
  NAND U2425 ( .A(n1894), .B(n1895), .Z(n1893) );
  OR U2426 ( .A(n1896), .B(n1897), .Z(n1894) );
  NANDN U2427 ( .A(n1898), .B(n1896), .Z(n1892) );
  XNOR U2428 ( .A(n1873), .B(n1899), .Z(N2682) );
  XOR U2429 ( .A(n1875), .B(n1876), .Z(n1899) );
  XNOR U2430 ( .A(n1889), .B(n1900), .Z(n1876) );
  XOR U2431 ( .A(n1890), .B(n1891), .Z(n1900) );
  XOR U2432 ( .A(n1896), .B(n1901), .Z(n1891) );
  XOR U2433 ( .A(n1895), .B(n1898), .Z(n1901) );
  IV U2434 ( .A(n1897), .Z(n1898) );
  NAND U2435 ( .A(n1902), .B(n1903), .Z(n1897) );
  OR U2436 ( .A(n1904), .B(n1905), .Z(n1903) );
  OR U2437 ( .A(n1906), .B(n1907), .Z(n1902) );
  NAND U2438 ( .A(n1908), .B(n1909), .Z(n1895) );
  OR U2439 ( .A(n1910), .B(n1911), .Z(n1909) );
  OR U2440 ( .A(n1912), .B(n1913), .Z(n1908) );
  NOR U2441 ( .A(n1914), .B(n1915), .Z(n1896) );
  ANDN U2442 ( .B(n1916), .A(n1917), .Z(n1890) );
  XNOR U2443 ( .A(n1883), .B(n1918), .Z(n1889) );
  XNOR U2444 ( .A(n1882), .B(n1884), .Z(n1918) );
  NAND U2445 ( .A(n1919), .B(n1920), .Z(n1884) );
  OR U2446 ( .A(n1921), .B(n1922), .Z(n1920) );
  OR U2447 ( .A(n1923), .B(n1924), .Z(n1919) );
  NAND U2448 ( .A(n1925), .B(n1926), .Z(n1882) );
  OR U2449 ( .A(n1927), .B(n1928), .Z(n1926) );
  OR U2450 ( .A(n1929), .B(n1930), .Z(n1925) );
  ANDN U2451 ( .B(n1931), .A(n1932), .Z(n1883) );
  IV U2452 ( .A(n1933), .Z(n1931) );
  ANDN U2453 ( .B(n1934), .A(n1935), .Z(n1875) );
  XOR U2454 ( .A(n1861), .B(n1936), .Z(n1873) );
  XOR U2455 ( .A(n1862), .B(n1863), .Z(n1936) );
  XOR U2456 ( .A(n1868), .B(n1937), .Z(n1863) );
  XOR U2457 ( .A(n1867), .B(n1870), .Z(n1937) );
  IV U2458 ( .A(n1869), .Z(n1870) );
  NAND U2459 ( .A(n1938), .B(n1939), .Z(n1869) );
  OR U2460 ( .A(n1940), .B(n1941), .Z(n1939) );
  OR U2461 ( .A(n1942), .B(n1943), .Z(n1938) );
  NAND U2462 ( .A(n1944), .B(n1945), .Z(n1867) );
  OR U2463 ( .A(n1946), .B(n1947), .Z(n1945) );
  OR U2464 ( .A(n1948), .B(n1949), .Z(n1944) );
  NOR U2465 ( .A(n1950), .B(n1951), .Z(n1868) );
  ANDN U2466 ( .B(n1952), .A(n1953), .Z(n1862) );
  IV U2467 ( .A(n1954), .Z(n1952) );
  XNOR U2468 ( .A(n1855), .B(n1955), .Z(n1861) );
  XNOR U2469 ( .A(n1854), .B(n1856), .Z(n1955) );
  NAND U2470 ( .A(n1956), .B(n1957), .Z(n1856) );
  OR U2471 ( .A(n1958), .B(n1959), .Z(n1957) );
  OR U2472 ( .A(n1960), .B(n1961), .Z(n1956) );
  NAND U2473 ( .A(n1962), .B(n1963), .Z(n1854) );
  OR U2474 ( .A(n1964), .B(n1965), .Z(n1963) );
  OR U2475 ( .A(n1966), .B(n1967), .Z(n1962) );
  ANDN U2476 ( .B(n1968), .A(n1969), .Z(n1855) );
  IV U2477 ( .A(n1970), .Z(n1968) );
  XNOR U2478 ( .A(n1935), .B(n1934), .Z(N2681) );
  XOR U2479 ( .A(n1954), .B(n1953), .Z(n1934) );
  XNOR U2480 ( .A(n1969), .B(n1970), .Z(n1953) );
  XNOR U2481 ( .A(n1964), .B(n1965), .Z(n1970) );
  XNOR U2482 ( .A(n1966), .B(n1967), .Z(n1965) );
  XNOR U2483 ( .A(y[253]), .B(x[253]), .Z(n1967) );
  XNOR U2484 ( .A(y[254]), .B(x[254]), .Z(n1966) );
  XNOR U2485 ( .A(y[252]), .B(x[252]), .Z(n1964) );
  XNOR U2486 ( .A(n1958), .B(n1959), .Z(n1969) );
  XNOR U2487 ( .A(y[249]), .B(x[249]), .Z(n1959) );
  XNOR U2488 ( .A(n1960), .B(n1961), .Z(n1958) );
  XNOR U2489 ( .A(y[250]), .B(x[250]), .Z(n1961) );
  XNOR U2490 ( .A(y[251]), .B(x[251]), .Z(n1960) );
  XNOR U2491 ( .A(n1951), .B(n1950), .Z(n1954) );
  XNOR U2492 ( .A(n1946), .B(n1947), .Z(n1950) );
  XNOR U2493 ( .A(y[246]), .B(x[246]), .Z(n1947) );
  XNOR U2494 ( .A(n1948), .B(n1949), .Z(n1946) );
  XNOR U2495 ( .A(y[247]), .B(x[247]), .Z(n1949) );
  XNOR U2496 ( .A(y[248]), .B(x[248]), .Z(n1948) );
  XNOR U2497 ( .A(n1940), .B(n1941), .Z(n1951) );
  XNOR U2498 ( .A(y[243]), .B(x[243]), .Z(n1941) );
  XNOR U2499 ( .A(n1942), .B(n1943), .Z(n1940) );
  XNOR U2500 ( .A(y[244]), .B(x[244]), .Z(n1943) );
  XNOR U2501 ( .A(y[245]), .B(x[245]), .Z(n1942) );
  XOR U2502 ( .A(n1916), .B(n1917), .Z(n1935) );
  XNOR U2503 ( .A(n1932), .B(n1933), .Z(n1917) );
  XNOR U2504 ( .A(n1927), .B(n1928), .Z(n1933) );
  XNOR U2505 ( .A(n1929), .B(n1930), .Z(n1928) );
  XNOR U2506 ( .A(y[241]), .B(x[241]), .Z(n1930) );
  XNOR U2507 ( .A(y[242]), .B(x[242]), .Z(n1929) );
  XNOR U2508 ( .A(y[240]), .B(x[240]), .Z(n1927) );
  XNOR U2509 ( .A(n1921), .B(n1922), .Z(n1932) );
  XNOR U2510 ( .A(y[237]), .B(x[237]), .Z(n1922) );
  XNOR U2511 ( .A(n1923), .B(n1924), .Z(n1921) );
  XNOR U2512 ( .A(y[238]), .B(x[238]), .Z(n1924) );
  XNOR U2513 ( .A(y[239]), .B(x[239]), .Z(n1923) );
  XOR U2514 ( .A(n1915), .B(n1914), .Z(n1916) );
  XNOR U2515 ( .A(n1910), .B(n1911), .Z(n1914) );
  XNOR U2516 ( .A(y[234]), .B(x[234]), .Z(n1911) );
  XNOR U2517 ( .A(n1912), .B(n1913), .Z(n1910) );
  XNOR U2518 ( .A(y[235]), .B(x[235]), .Z(n1913) );
  XNOR U2519 ( .A(y[236]), .B(x[236]), .Z(n1912) );
  XNOR U2520 ( .A(n1904), .B(n1905), .Z(n1915) );
  XNOR U2521 ( .A(y[231]), .B(x[231]), .Z(n1905) );
  XNOR U2522 ( .A(n1906), .B(n1907), .Z(n1904) );
  XNOR U2523 ( .A(y[232]), .B(x[232]), .Z(n1907) );
  XNOR U2524 ( .A(y[233]), .B(x[233]), .Z(n1906) );
  NAND U2525 ( .A(n1971), .B(n1972), .Z(N2676) );
  NANDN U2526 ( .A(n1973), .B(n1974), .Z(n1972) );
  OR U2527 ( .A(n1975), .B(n1976), .Z(n1974) );
  NAND U2528 ( .A(n1975), .B(n1976), .Z(n1971) );
  XOR U2529 ( .A(n1975), .B(n1977), .Z(N2675) );
  XNOR U2530 ( .A(n1973), .B(n1976), .Z(n1977) );
  AND U2531 ( .A(n1978), .B(n1979), .Z(n1976) );
  NANDN U2532 ( .A(n1980), .B(n1981), .Z(n1979) );
  NANDN U2533 ( .A(n1982), .B(n1983), .Z(n1981) );
  NANDN U2534 ( .A(n1983), .B(n1982), .Z(n1978) );
  NAND U2535 ( .A(n1984), .B(n1985), .Z(n1973) );
  NANDN U2536 ( .A(n1986), .B(n1987), .Z(n1985) );
  OR U2537 ( .A(n1988), .B(n1989), .Z(n1987) );
  NAND U2538 ( .A(n1989), .B(n1988), .Z(n1984) );
  AND U2539 ( .A(n1990), .B(n1991), .Z(n1975) );
  NANDN U2540 ( .A(n1992), .B(n1993), .Z(n1991) );
  NANDN U2541 ( .A(n1994), .B(n1995), .Z(n1993) );
  NANDN U2542 ( .A(n1995), .B(n1994), .Z(n1990) );
  XOR U2543 ( .A(n1989), .B(n1996), .Z(N2674) );
  XOR U2544 ( .A(n1986), .B(n1988), .Z(n1996) );
  XNOR U2545 ( .A(n1982), .B(n1997), .Z(n1988) );
  XNOR U2546 ( .A(n1980), .B(n1983), .Z(n1997) );
  NAND U2547 ( .A(n1998), .B(n1999), .Z(n1983) );
  NAND U2548 ( .A(n2000), .B(n2001), .Z(n1999) );
  OR U2549 ( .A(n2002), .B(n2003), .Z(n2000) );
  NANDN U2550 ( .A(n2004), .B(n2002), .Z(n1998) );
  IV U2551 ( .A(n2003), .Z(n2004) );
  NAND U2552 ( .A(n2005), .B(n2006), .Z(n1980) );
  NAND U2553 ( .A(n2007), .B(n2008), .Z(n2006) );
  NANDN U2554 ( .A(n2009), .B(n2010), .Z(n2007) );
  NANDN U2555 ( .A(n2010), .B(n2009), .Z(n2005) );
  AND U2556 ( .A(n2011), .B(n2012), .Z(n1982) );
  NAND U2557 ( .A(n2013), .B(n2014), .Z(n2012) );
  OR U2558 ( .A(n2015), .B(n2016), .Z(n2013) );
  NANDN U2559 ( .A(n2017), .B(n2015), .Z(n2011) );
  NAND U2560 ( .A(n2018), .B(n2019), .Z(n1986) );
  NANDN U2561 ( .A(n2020), .B(n2021), .Z(n2019) );
  OR U2562 ( .A(n2022), .B(n2023), .Z(n2021) );
  NANDN U2563 ( .A(n2024), .B(n2022), .Z(n2018) );
  IV U2564 ( .A(n2023), .Z(n2024) );
  XNOR U2565 ( .A(n1994), .B(n2025), .Z(n1989) );
  XNOR U2566 ( .A(n1992), .B(n1995), .Z(n2025) );
  NAND U2567 ( .A(n2026), .B(n2027), .Z(n1995) );
  NAND U2568 ( .A(n2028), .B(n2029), .Z(n2027) );
  OR U2569 ( .A(n2030), .B(n2031), .Z(n2028) );
  NANDN U2570 ( .A(n2032), .B(n2030), .Z(n2026) );
  IV U2571 ( .A(n2031), .Z(n2032) );
  NAND U2572 ( .A(n2033), .B(n2034), .Z(n1992) );
  NAND U2573 ( .A(n2035), .B(n2036), .Z(n2034) );
  NANDN U2574 ( .A(n2037), .B(n2038), .Z(n2035) );
  NANDN U2575 ( .A(n2038), .B(n2037), .Z(n2033) );
  AND U2576 ( .A(n2039), .B(n2040), .Z(n1994) );
  NAND U2577 ( .A(n2041), .B(n2042), .Z(n2040) );
  OR U2578 ( .A(n2043), .B(n2044), .Z(n2041) );
  NANDN U2579 ( .A(n2045), .B(n2043), .Z(n2039) );
  XNOR U2580 ( .A(n2020), .B(n2046), .Z(N2673) );
  XOR U2581 ( .A(n2022), .B(n2023), .Z(n2046) );
  XNOR U2582 ( .A(n2036), .B(n2047), .Z(n2023) );
  XOR U2583 ( .A(n2037), .B(n2038), .Z(n2047) );
  XOR U2584 ( .A(n2043), .B(n2048), .Z(n2038) );
  XOR U2585 ( .A(n2042), .B(n2045), .Z(n2048) );
  IV U2586 ( .A(n2044), .Z(n2045) );
  NAND U2587 ( .A(n2049), .B(n2050), .Z(n2044) );
  OR U2588 ( .A(n2051), .B(n2052), .Z(n2050) );
  OR U2589 ( .A(n2053), .B(n2054), .Z(n2049) );
  NAND U2590 ( .A(n2055), .B(n2056), .Z(n2042) );
  OR U2591 ( .A(n2057), .B(n2058), .Z(n2056) );
  OR U2592 ( .A(n2059), .B(n2060), .Z(n2055) );
  NOR U2593 ( .A(n2061), .B(n2062), .Z(n2043) );
  ANDN U2594 ( .B(n2063), .A(n2064), .Z(n2037) );
  XNOR U2595 ( .A(n2030), .B(n2065), .Z(n2036) );
  XNOR U2596 ( .A(n2029), .B(n2031), .Z(n2065) );
  NAND U2597 ( .A(n2066), .B(n2067), .Z(n2031) );
  OR U2598 ( .A(n2068), .B(n2069), .Z(n2067) );
  OR U2599 ( .A(n2070), .B(n2071), .Z(n2066) );
  NAND U2600 ( .A(n2072), .B(n2073), .Z(n2029) );
  OR U2601 ( .A(n2074), .B(n2075), .Z(n2073) );
  OR U2602 ( .A(n2076), .B(n2077), .Z(n2072) );
  ANDN U2603 ( .B(n2078), .A(n2079), .Z(n2030) );
  IV U2604 ( .A(n2080), .Z(n2078) );
  ANDN U2605 ( .B(n2081), .A(n2082), .Z(n2022) );
  XOR U2606 ( .A(n2008), .B(n2083), .Z(n2020) );
  XOR U2607 ( .A(n2009), .B(n2010), .Z(n2083) );
  XOR U2608 ( .A(n2015), .B(n2084), .Z(n2010) );
  XOR U2609 ( .A(n2014), .B(n2017), .Z(n2084) );
  IV U2610 ( .A(n2016), .Z(n2017) );
  NAND U2611 ( .A(n2085), .B(n2086), .Z(n2016) );
  OR U2612 ( .A(n2087), .B(n2088), .Z(n2086) );
  OR U2613 ( .A(n2089), .B(n2090), .Z(n2085) );
  NAND U2614 ( .A(n2091), .B(n2092), .Z(n2014) );
  OR U2615 ( .A(n2093), .B(n2094), .Z(n2092) );
  OR U2616 ( .A(n2095), .B(n2096), .Z(n2091) );
  NOR U2617 ( .A(n2097), .B(n2098), .Z(n2015) );
  ANDN U2618 ( .B(n2099), .A(n2100), .Z(n2009) );
  IV U2619 ( .A(n2101), .Z(n2099) );
  XNOR U2620 ( .A(n2002), .B(n2102), .Z(n2008) );
  XNOR U2621 ( .A(n2001), .B(n2003), .Z(n2102) );
  NAND U2622 ( .A(n2103), .B(n2104), .Z(n2003) );
  OR U2623 ( .A(n2105), .B(n2106), .Z(n2104) );
  OR U2624 ( .A(n2107), .B(n2108), .Z(n2103) );
  NAND U2625 ( .A(n2109), .B(n2110), .Z(n2001) );
  OR U2626 ( .A(n2111), .B(n2112), .Z(n2110) );
  OR U2627 ( .A(n2113), .B(n2114), .Z(n2109) );
  ANDN U2628 ( .B(n2115), .A(n2116), .Z(n2002) );
  IV U2629 ( .A(n2117), .Z(n2115) );
  XNOR U2630 ( .A(n2082), .B(n2081), .Z(N2672) );
  XOR U2631 ( .A(n2101), .B(n2100), .Z(n2081) );
  XNOR U2632 ( .A(n2116), .B(n2117), .Z(n2100) );
  XNOR U2633 ( .A(n2111), .B(n2112), .Z(n2117) );
  XNOR U2634 ( .A(n2113), .B(n2114), .Z(n2112) );
  XNOR U2635 ( .A(y[229]), .B(x[229]), .Z(n2114) );
  XNOR U2636 ( .A(y[230]), .B(x[230]), .Z(n2113) );
  XNOR U2637 ( .A(y[228]), .B(x[228]), .Z(n2111) );
  XNOR U2638 ( .A(n2105), .B(n2106), .Z(n2116) );
  XNOR U2639 ( .A(y[225]), .B(x[225]), .Z(n2106) );
  XNOR U2640 ( .A(n2107), .B(n2108), .Z(n2105) );
  XNOR U2641 ( .A(y[226]), .B(x[226]), .Z(n2108) );
  XNOR U2642 ( .A(y[227]), .B(x[227]), .Z(n2107) );
  XNOR U2643 ( .A(n2098), .B(n2097), .Z(n2101) );
  XNOR U2644 ( .A(n2093), .B(n2094), .Z(n2097) );
  XNOR U2645 ( .A(y[222]), .B(x[222]), .Z(n2094) );
  XNOR U2646 ( .A(n2095), .B(n2096), .Z(n2093) );
  XNOR U2647 ( .A(y[223]), .B(x[223]), .Z(n2096) );
  XNOR U2648 ( .A(y[224]), .B(x[224]), .Z(n2095) );
  XNOR U2649 ( .A(n2087), .B(n2088), .Z(n2098) );
  XNOR U2650 ( .A(y[219]), .B(x[219]), .Z(n2088) );
  XNOR U2651 ( .A(n2089), .B(n2090), .Z(n2087) );
  XNOR U2652 ( .A(y[220]), .B(x[220]), .Z(n2090) );
  XNOR U2653 ( .A(y[221]), .B(x[221]), .Z(n2089) );
  XOR U2654 ( .A(n2063), .B(n2064), .Z(n2082) );
  XNOR U2655 ( .A(n2079), .B(n2080), .Z(n2064) );
  XNOR U2656 ( .A(n2074), .B(n2075), .Z(n2080) );
  XNOR U2657 ( .A(n2076), .B(n2077), .Z(n2075) );
  XNOR U2658 ( .A(y[217]), .B(x[217]), .Z(n2077) );
  XNOR U2659 ( .A(y[218]), .B(x[218]), .Z(n2076) );
  XNOR U2660 ( .A(y[216]), .B(x[216]), .Z(n2074) );
  XNOR U2661 ( .A(n2068), .B(n2069), .Z(n2079) );
  XNOR U2662 ( .A(y[213]), .B(x[213]), .Z(n2069) );
  XNOR U2663 ( .A(n2070), .B(n2071), .Z(n2068) );
  XNOR U2664 ( .A(y[214]), .B(x[214]), .Z(n2071) );
  XNOR U2665 ( .A(y[215]), .B(x[215]), .Z(n2070) );
  XOR U2666 ( .A(n2062), .B(n2061), .Z(n2063) );
  XNOR U2667 ( .A(n2057), .B(n2058), .Z(n2061) );
  XNOR U2668 ( .A(y[210]), .B(x[210]), .Z(n2058) );
  XNOR U2669 ( .A(n2059), .B(n2060), .Z(n2057) );
  XNOR U2670 ( .A(y[211]), .B(x[211]), .Z(n2060) );
  XNOR U2671 ( .A(y[212]), .B(x[212]), .Z(n2059) );
  XNOR U2672 ( .A(n2051), .B(n2052), .Z(n2062) );
  XNOR U2673 ( .A(y[207]), .B(x[207]), .Z(n2052) );
  XNOR U2674 ( .A(n2053), .B(n2054), .Z(n2051) );
  XNOR U2675 ( .A(y[208]), .B(x[208]), .Z(n2054) );
  XNOR U2676 ( .A(y[209]), .B(x[209]), .Z(n2053) );
  NAND U2677 ( .A(n2118), .B(n2119), .Z(N2667) );
  NANDN U2678 ( .A(n2120), .B(n2121), .Z(n2119) );
  OR U2679 ( .A(n2122), .B(n2123), .Z(n2121) );
  NAND U2680 ( .A(n2122), .B(n2123), .Z(n2118) );
  XOR U2681 ( .A(n2122), .B(n2124), .Z(N2666) );
  XNOR U2682 ( .A(n2120), .B(n2123), .Z(n2124) );
  AND U2683 ( .A(n2125), .B(n2126), .Z(n2123) );
  NANDN U2684 ( .A(n2127), .B(n2128), .Z(n2126) );
  NANDN U2685 ( .A(n2129), .B(n2130), .Z(n2128) );
  NANDN U2686 ( .A(n2130), .B(n2129), .Z(n2125) );
  NAND U2687 ( .A(n2131), .B(n2132), .Z(n2120) );
  NANDN U2688 ( .A(n2133), .B(n2134), .Z(n2132) );
  OR U2689 ( .A(n2135), .B(n2136), .Z(n2134) );
  NAND U2690 ( .A(n2136), .B(n2135), .Z(n2131) );
  AND U2691 ( .A(n2137), .B(n2138), .Z(n2122) );
  NANDN U2692 ( .A(n2139), .B(n2140), .Z(n2138) );
  NANDN U2693 ( .A(n2141), .B(n2142), .Z(n2140) );
  NANDN U2694 ( .A(n2142), .B(n2141), .Z(n2137) );
  XOR U2695 ( .A(n2136), .B(n2143), .Z(N2665) );
  XOR U2696 ( .A(n2133), .B(n2135), .Z(n2143) );
  XNOR U2697 ( .A(n2129), .B(n2144), .Z(n2135) );
  XNOR U2698 ( .A(n2127), .B(n2130), .Z(n2144) );
  NAND U2699 ( .A(n2145), .B(n2146), .Z(n2130) );
  NAND U2700 ( .A(n2147), .B(n2148), .Z(n2146) );
  OR U2701 ( .A(n2149), .B(n2150), .Z(n2147) );
  NANDN U2702 ( .A(n2151), .B(n2149), .Z(n2145) );
  IV U2703 ( .A(n2150), .Z(n2151) );
  NAND U2704 ( .A(n2152), .B(n2153), .Z(n2127) );
  NAND U2705 ( .A(n2154), .B(n2155), .Z(n2153) );
  NANDN U2706 ( .A(n2156), .B(n2157), .Z(n2154) );
  NANDN U2707 ( .A(n2157), .B(n2156), .Z(n2152) );
  AND U2708 ( .A(n2158), .B(n2159), .Z(n2129) );
  NAND U2709 ( .A(n2160), .B(n2161), .Z(n2159) );
  OR U2710 ( .A(n2162), .B(n2163), .Z(n2160) );
  NANDN U2711 ( .A(n2164), .B(n2162), .Z(n2158) );
  NAND U2712 ( .A(n2165), .B(n2166), .Z(n2133) );
  NANDN U2713 ( .A(n2167), .B(n2168), .Z(n2166) );
  OR U2714 ( .A(n2169), .B(n2170), .Z(n2168) );
  NANDN U2715 ( .A(n2171), .B(n2169), .Z(n2165) );
  IV U2716 ( .A(n2170), .Z(n2171) );
  XNOR U2717 ( .A(n2141), .B(n2172), .Z(n2136) );
  XNOR U2718 ( .A(n2139), .B(n2142), .Z(n2172) );
  NAND U2719 ( .A(n2173), .B(n2174), .Z(n2142) );
  NAND U2720 ( .A(n2175), .B(n2176), .Z(n2174) );
  OR U2721 ( .A(n2177), .B(n2178), .Z(n2175) );
  NANDN U2722 ( .A(n2179), .B(n2177), .Z(n2173) );
  IV U2723 ( .A(n2178), .Z(n2179) );
  NAND U2724 ( .A(n2180), .B(n2181), .Z(n2139) );
  NAND U2725 ( .A(n2182), .B(n2183), .Z(n2181) );
  NANDN U2726 ( .A(n2184), .B(n2185), .Z(n2182) );
  NANDN U2727 ( .A(n2185), .B(n2184), .Z(n2180) );
  AND U2728 ( .A(n2186), .B(n2187), .Z(n2141) );
  NAND U2729 ( .A(n2188), .B(n2189), .Z(n2187) );
  OR U2730 ( .A(n2190), .B(n2191), .Z(n2188) );
  NANDN U2731 ( .A(n2192), .B(n2190), .Z(n2186) );
  XNOR U2732 ( .A(n2167), .B(n2193), .Z(N2664) );
  XOR U2733 ( .A(n2169), .B(n2170), .Z(n2193) );
  XNOR U2734 ( .A(n2183), .B(n2194), .Z(n2170) );
  XOR U2735 ( .A(n2184), .B(n2185), .Z(n2194) );
  XOR U2736 ( .A(n2190), .B(n2195), .Z(n2185) );
  XOR U2737 ( .A(n2189), .B(n2192), .Z(n2195) );
  IV U2738 ( .A(n2191), .Z(n2192) );
  NAND U2739 ( .A(n2196), .B(n2197), .Z(n2191) );
  OR U2740 ( .A(n2198), .B(n2199), .Z(n2197) );
  OR U2741 ( .A(n2200), .B(n2201), .Z(n2196) );
  NAND U2742 ( .A(n2202), .B(n2203), .Z(n2189) );
  OR U2743 ( .A(n2204), .B(n2205), .Z(n2203) );
  OR U2744 ( .A(n2206), .B(n2207), .Z(n2202) );
  NOR U2745 ( .A(n2208), .B(n2209), .Z(n2190) );
  ANDN U2746 ( .B(n2210), .A(n2211), .Z(n2184) );
  XNOR U2747 ( .A(n2177), .B(n2212), .Z(n2183) );
  XNOR U2748 ( .A(n2176), .B(n2178), .Z(n2212) );
  NAND U2749 ( .A(n2213), .B(n2214), .Z(n2178) );
  OR U2750 ( .A(n2215), .B(n2216), .Z(n2214) );
  OR U2751 ( .A(n2217), .B(n2218), .Z(n2213) );
  NAND U2752 ( .A(n2219), .B(n2220), .Z(n2176) );
  OR U2753 ( .A(n2221), .B(n2222), .Z(n2220) );
  OR U2754 ( .A(n2223), .B(n2224), .Z(n2219) );
  ANDN U2755 ( .B(n2225), .A(n2226), .Z(n2177) );
  IV U2756 ( .A(n2227), .Z(n2225) );
  ANDN U2757 ( .B(n2228), .A(n2229), .Z(n2169) );
  XOR U2758 ( .A(n2155), .B(n2230), .Z(n2167) );
  XOR U2759 ( .A(n2156), .B(n2157), .Z(n2230) );
  XOR U2760 ( .A(n2162), .B(n2231), .Z(n2157) );
  XOR U2761 ( .A(n2161), .B(n2164), .Z(n2231) );
  IV U2762 ( .A(n2163), .Z(n2164) );
  NAND U2763 ( .A(n2232), .B(n2233), .Z(n2163) );
  OR U2764 ( .A(n2234), .B(n2235), .Z(n2233) );
  OR U2765 ( .A(n2236), .B(n2237), .Z(n2232) );
  NAND U2766 ( .A(n2238), .B(n2239), .Z(n2161) );
  OR U2767 ( .A(n2240), .B(n2241), .Z(n2239) );
  OR U2768 ( .A(n2242), .B(n2243), .Z(n2238) );
  NOR U2769 ( .A(n2244), .B(n2245), .Z(n2162) );
  ANDN U2770 ( .B(n2246), .A(n2247), .Z(n2156) );
  IV U2771 ( .A(n2248), .Z(n2246) );
  XNOR U2772 ( .A(n2149), .B(n2249), .Z(n2155) );
  XNOR U2773 ( .A(n2148), .B(n2150), .Z(n2249) );
  NAND U2774 ( .A(n2250), .B(n2251), .Z(n2150) );
  OR U2775 ( .A(n2252), .B(n2253), .Z(n2251) );
  OR U2776 ( .A(n2254), .B(n2255), .Z(n2250) );
  NAND U2777 ( .A(n2256), .B(n2257), .Z(n2148) );
  OR U2778 ( .A(n2258), .B(n2259), .Z(n2257) );
  OR U2779 ( .A(n2260), .B(n2261), .Z(n2256) );
  ANDN U2780 ( .B(n2262), .A(n2263), .Z(n2149) );
  IV U2781 ( .A(n2264), .Z(n2262) );
  XNOR U2782 ( .A(n2229), .B(n2228), .Z(N2663) );
  XOR U2783 ( .A(n2248), .B(n2247), .Z(n2228) );
  XNOR U2784 ( .A(n2263), .B(n2264), .Z(n2247) );
  XNOR U2785 ( .A(n2258), .B(n2259), .Z(n2264) );
  XNOR U2786 ( .A(n2260), .B(n2261), .Z(n2259) );
  XNOR U2787 ( .A(y[205]), .B(x[205]), .Z(n2261) );
  XNOR U2788 ( .A(y[206]), .B(x[206]), .Z(n2260) );
  XNOR U2789 ( .A(y[204]), .B(x[204]), .Z(n2258) );
  XNOR U2790 ( .A(n2252), .B(n2253), .Z(n2263) );
  XNOR U2791 ( .A(y[201]), .B(x[201]), .Z(n2253) );
  XNOR U2792 ( .A(n2254), .B(n2255), .Z(n2252) );
  XNOR U2793 ( .A(y[202]), .B(x[202]), .Z(n2255) );
  XNOR U2794 ( .A(y[203]), .B(x[203]), .Z(n2254) );
  XNOR U2795 ( .A(n2245), .B(n2244), .Z(n2248) );
  XNOR U2796 ( .A(n2240), .B(n2241), .Z(n2244) );
  XNOR U2797 ( .A(y[198]), .B(x[198]), .Z(n2241) );
  XNOR U2798 ( .A(n2242), .B(n2243), .Z(n2240) );
  XNOR U2799 ( .A(y[199]), .B(x[199]), .Z(n2243) );
  XNOR U2800 ( .A(y[200]), .B(x[200]), .Z(n2242) );
  XNOR U2801 ( .A(n2234), .B(n2235), .Z(n2245) );
  XNOR U2802 ( .A(y[195]), .B(x[195]), .Z(n2235) );
  XNOR U2803 ( .A(n2236), .B(n2237), .Z(n2234) );
  XNOR U2804 ( .A(y[196]), .B(x[196]), .Z(n2237) );
  XNOR U2805 ( .A(y[197]), .B(x[197]), .Z(n2236) );
  XOR U2806 ( .A(n2210), .B(n2211), .Z(n2229) );
  XNOR U2807 ( .A(n2226), .B(n2227), .Z(n2211) );
  XNOR U2808 ( .A(n2221), .B(n2222), .Z(n2227) );
  XNOR U2809 ( .A(n2223), .B(n2224), .Z(n2222) );
  XNOR U2810 ( .A(y[193]), .B(x[193]), .Z(n2224) );
  XNOR U2811 ( .A(y[194]), .B(x[194]), .Z(n2223) );
  XNOR U2812 ( .A(y[192]), .B(x[192]), .Z(n2221) );
  XNOR U2813 ( .A(n2215), .B(n2216), .Z(n2226) );
  XNOR U2814 ( .A(y[189]), .B(x[189]), .Z(n2216) );
  XNOR U2815 ( .A(n2217), .B(n2218), .Z(n2215) );
  XNOR U2816 ( .A(y[190]), .B(x[190]), .Z(n2218) );
  XNOR U2817 ( .A(y[191]), .B(x[191]), .Z(n2217) );
  XOR U2818 ( .A(n2209), .B(n2208), .Z(n2210) );
  XNOR U2819 ( .A(n2204), .B(n2205), .Z(n2208) );
  XNOR U2820 ( .A(y[186]), .B(x[186]), .Z(n2205) );
  XNOR U2821 ( .A(n2206), .B(n2207), .Z(n2204) );
  XNOR U2822 ( .A(y[187]), .B(x[187]), .Z(n2207) );
  XNOR U2823 ( .A(y[188]), .B(x[188]), .Z(n2206) );
  XNOR U2824 ( .A(n2198), .B(n2199), .Z(n2209) );
  XNOR U2825 ( .A(y[183]), .B(x[183]), .Z(n2199) );
  XNOR U2826 ( .A(n2200), .B(n2201), .Z(n2198) );
  XNOR U2827 ( .A(y[184]), .B(x[184]), .Z(n2201) );
  XNOR U2828 ( .A(y[185]), .B(x[185]), .Z(n2200) );
  NAND U2829 ( .A(n2265), .B(n2266), .Z(N2658) );
  NANDN U2830 ( .A(n2267), .B(n2268), .Z(n2266) );
  OR U2831 ( .A(n2269), .B(n2270), .Z(n2268) );
  NAND U2832 ( .A(n2269), .B(n2270), .Z(n2265) );
  XOR U2833 ( .A(n2269), .B(n2271), .Z(N2657) );
  XNOR U2834 ( .A(n2267), .B(n2270), .Z(n2271) );
  AND U2835 ( .A(n2272), .B(n2273), .Z(n2270) );
  NANDN U2836 ( .A(n2274), .B(n2275), .Z(n2273) );
  NANDN U2837 ( .A(n2276), .B(n2277), .Z(n2275) );
  NANDN U2838 ( .A(n2277), .B(n2276), .Z(n2272) );
  NAND U2839 ( .A(n2278), .B(n2279), .Z(n2267) );
  NANDN U2840 ( .A(n2280), .B(n2281), .Z(n2279) );
  OR U2841 ( .A(n2282), .B(n2283), .Z(n2281) );
  NAND U2842 ( .A(n2283), .B(n2282), .Z(n2278) );
  AND U2843 ( .A(n2284), .B(n2285), .Z(n2269) );
  NANDN U2844 ( .A(n2286), .B(n2287), .Z(n2285) );
  NANDN U2845 ( .A(n2288), .B(n2289), .Z(n2287) );
  NANDN U2846 ( .A(n2289), .B(n2288), .Z(n2284) );
  XOR U2847 ( .A(n2283), .B(n2290), .Z(N2656) );
  XOR U2848 ( .A(n2280), .B(n2282), .Z(n2290) );
  XNOR U2849 ( .A(n2276), .B(n2291), .Z(n2282) );
  XNOR U2850 ( .A(n2274), .B(n2277), .Z(n2291) );
  NAND U2851 ( .A(n2292), .B(n2293), .Z(n2277) );
  NAND U2852 ( .A(n2294), .B(n2295), .Z(n2293) );
  OR U2853 ( .A(n2296), .B(n2297), .Z(n2294) );
  NANDN U2854 ( .A(n2298), .B(n2296), .Z(n2292) );
  IV U2855 ( .A(n2297), .Z(n2298) );
  NAND U2856 ( .A(n2299), .B(n2300), .Z(n2274) );
  NAND U2857 ( .A(n2301), .B(n2302), .Z(n2300) );
  NANDN U2858 ( .A(n2303), .B(n2304), .Z(n2301) );
  NANDN U2859 ( .A(n2304), .B(n2303), .Z(n2299) );
  AND U2860 ( .A(n2305), .B(n2306), .Z(n2276) );
  NAND U2861 ( .A(n2307), .B(n2308), .Z(n2306) );
  OR U2862 ( .A(n2309), .B(n2310), .Z(n2307) );
  NANDN U2863 ( .A(n2311), .B(n2309), .Z(n2305) );
  NAND U2864 ( .A(n2312), .B(n2313), .Z(n2280) );
  NANDN U2865 ( .A(n2314), .B(n2315), .Z(n2313) );
  OR U2866 ( .A(n2316), .B(n2317), .Z(n2315) );
  NANDN U2867 ( .A(n2318), .B(n2316), .Z(n2312) );
  IV U2868 ( .A(n2317), .Z(n2318) );
  XNOR U2869 ( .A(n2288), .B(n2319), .Z(n2283) );
  XNOR U2870 ( .A(n2286), .B(n2289), .Z(n2319) );
  NAND U2871 ( .A(n2320), .B(n2321), .Z(n2289) );
  NAND U2872 ( .A(n2322), .B(n2323), .Z(n2321) );
  OR U2873 ( .A(n2324), .B(n2325), .Z(n2322) );
  NANDN U2874 ( .A(n2326), .B(n2324), .Z(n2320) );
  IV U2875 ( .A(n2325), .Z(n2326) );
  NAND U2876 ( .A(n2327), .B(n2328), .Z(n2286) );
  NAND U2877 ( .A(n2329), .B(n2330), .Z(n2328) );
  NANDN U2878 ( .A(n2331), .B(n2332), .Z(n2329) );
  NANDN U2879 ( .A(n2332), .B(n2331), .Z(n2327) );
  AND U2880 ( .A(n2333), .B(n2334), .Z(n2288) );
  NAND U2881 ( .A(n2335), .B(n2336), .Z(n2334) );
  OR U2882 ( .A(n2337), .B(n2338), .Z(n2335) );
  NANDN U2883 ( .A(n2339), .B(n2337), .Z(n2333) );
  XNOR U2884 ( .A(n2314), .B(n2340), .Z(N2655) );
  XOR U2885 ( .A(n2316), .B(n2317), .Z(n2340) );
  XNOR U2886 ( .A(n2330), .B(n2341), .Z(n2317) );
  XOR U2887 ( .A(n2331), .B(n2332), .Z(n2341) );
  XOR U2888 ( .A(n2337), .B(n2342), .Z(n2332) );
  XOR U2889 ( .A(n2336), .B(n2339), .Z(n2342) );
  IV U2890 ( .A(n2338), .Z(n2339) );
  NAND U2891 ( .A(n2343), .B(n2344), .Z(n2338) );
  OR U2892 ( .A(n2345), .B(n2346), .Z(n2344) );
  OR U2893 ( .A(n2347), .B(n2348), .Z(n2343) );
  NAND U2894 ( .A(n2349), .B(n2350), .Z(n2336) );
  OR U2895 ( .A(n2351), .B(n2352), .Z(n2350) );
  OR U2896 ( .A(n2353), .B(n2354), .Z(n2349) );
  NOR U2897 ( .A(n2355), .B(n2356), .Z(n2337) );
  ANDN U2898 ( .B(n2357), .A(n2358), .Z(n2331) );
  XNOR U2899 ( .A(n2324), .B(n2359), .Z(n2330) );
  XNOR U2900 ( .A(n2323), .B(n2325), .Z(n2359) );
  NAND U2901 ( .A(n2360), .B(n2361), .Z(n2325) );
  OR U2902 ( .A(n2362), .B(n2363), .Z(n2361) );
  OR U2903 ( .A(n2364), .B(n2365), .Z(n2360) );
  NAND U2904 ( .A(n2366), .B(n2367), .Z(n2323) );
  OR U2905 ( .A(n2368), .B(n2369), .Z(n2367) );
  OR U2906 ( .A(n2370), .B(n2371), .Z(n2366) );
  ANDN U2907 ( .B(n2372), .A(n2373), .Z(n2324) );
  IV U2908 ( .A(n2374), .Z(n2372) );
  ANDN U2909 ( .B(n2375), .A(n2376), .Z(n2316) );
  XOR U2910 ( .A(n2302), .B(n2377), .Z(n2314) );
  XOR U2911 ( .A(n2303), .B(n2304), .Z(n2377) );
  XOR U2912 ( .A(n2309), .B(n2378), .Z(n2304) );
  XOR U2913 ( .A(n2308), .B(n2311), .Z(n2378) );
  IV U2914 ( .A(n2310), .Z(n2311) );
  NAND U2915 ( .A(n2379), .B(n2380), .Z(n2310) );
  OR U2916 ( .A(n2381), .B(n2382), .Z(n2380) );
  OR U2917 ( .A(n2383), .B(n2384), .Z(n2379) );
  NAND U2918 ( .A(n2385), .B(n2386), .Z(n2308) );
  OR U2919 ( .A(n2387), .B(n2388), .Z(n2386) );
  OR U2920 ( .A(n2389), .B(n2390), .Z(n2385) );
  NOR U2921 ( .A(n2391), .B(n2392), .Z(n2309) );
  ANDN U2922 ( .B(n2393), .A(n2394), .Z(n2303) );
  IV U2923 ( .A(n2395), .Z(n2393) );
  XNOR U2924 ( .A(n2296), .B(n2396), .Z(n2302) );
  XNOR U2925 ( .A(n2295), .B(n2297), .Z(n2396) );
  NAND U2926 ( .A(n2397), .B(n2398), .Z(n2297) );
  OR U2927 ( .A(n2399), .B(n2400), .Z(n2398) );
  OR U2928 ( .A(n2401), .B(n2402), .Z(n2397) );
  NAND U2929 ( .A(n2403), .B(n2404), .Z(n2295) );
  OR U2930 ( .A(n2405), .B(n2406), .Z(n2404) );
  OR U2931 ( .A(n2407), .B(n2408), .Z(n2403) );
  ANDN U2932 ( .B(n2409), .A(n2410), .Z(n2296) );
  IV U2933 ( .A(n2411), .Z(n2409) );
  XNOR U2934 ( .A(n2376), .B(n2375), .Z(N2654) );
  XOR U2935 ( .A(n2395), .B(n2394), .Z(n2375) );
  XNOR U2936 ( .A(n2410), .B(n2411), .Z(n2394) );
  XNOR U2937 ( .A(n2405), .B(n2406), .Z(n2411) );
  XNOR U2938 ( .A(n2407), .B(n2408), .Z(n2406) );
  XNOR U2939 ( .A(y[181]), .B(x[181]), .Z(n2408) );
  XNOR U2940 ( .A(y[182]), .B(x[182]), .Z(n2407) );
  XNOR U2941 ( .A(y[180]), .B(x[180]), .Z(n2405) );
  XNOR U2942 ( .A(n2399), .B(n2400), .Z(n2410) );
  XNOR U2943 ( .A(y[177]), .B(x[177]), .Z(n2400) );
  XNOR U2944 ( .A(n2401), .B(n2402), .Z(n2399) );
  XNOR U2945 ( .A(y[178]), .B(x[178]), .Z(n2402) );
  XNOR U2946 ( .A(y[179]), .B(x[179]), .Z(n2401) );
  XNOR U2947 ( .A(n2392), .B(n2391), .Z(n2395) );
  XNOR U2948 ( .A(n2387), .B(n2388), .Z(n2391) );
  XNOR U2949 ( .A(y[174]), .B(x[174]), .Z(n2388) );
  XNOR U2950 ( .A(n2389), .B(n2390), .Z(n2387) );
  XNOR U2951 ( .A(y[175]), .B(x[175]), .Z(n2390) );
  XNOR U2952 ( .A(y[176]), .B(x[176]), .Z(n2389) );
  XNOR U2953 ( .A(n2381), .B(n2382), .Z(n2392) );
  XNOR U2954 ( .A(y[171]), .B(x[171]), .Z(n2382) );
  XNOR U2955 ( .A(n2383), .B(n2384), .Z(n2381) );
  XNOR U2956 ( .A(y[172]), .B(x[172]), .Z(n2384) );
  XNOR U2957 ( .A(y[173]), .B(x[173]), .Z(n2383) );
  XOR U2958 ( .A(n2357), .B(n2358), .Z(n2376) );
  XNOR U2959 ( .A(n2373), .B(n2374), .Z(n2358) );
  XNOR U2960 ( .A(n2368), .B(n2369), .Z(n2374) );
  XNOR U2961 ( .A(n2370), .B(n2371), .Z(n2369) );
  XNOR U2962 ( .A(y[169]), .B(x[169]), .Z(n2371) );
  XNOR U2963 ( .A(y[170]), .B(x[170]), .Z(n2370) );
  XNOR U2964 ( .A(y[168]), .B(x[168]), .Z(n2368) );
  XNOR U2965 ( .A(n2362), .B(n2363), .Z(n2373) );
  XNOR U2966 ( .A(y[165]), .B(x[165]), .Z(n2363) );
  XNOR U2967 ( .A(n2364), .B(n2365), .Z(n2362) );
  XNOR U2968 ( .A(y[166]), .B(x[166]), .Z(n2365) );
  XNOR U2969 ( .A(y[167]), .B(x[167]), .Z(n2364) );
  XOR U2970 ( .A(n2356), .B(n2355), .Z(n2357) );
  XNOR U2971 ( .A(n2351), .B(n2352), .Z(n2355) );
  XNOR U2972 ( .A(y[162]), .B(x[162]), .Z(n2352) );
  XNOR U2973 ( .A(n2353), .B(n2354), .Z(n2351) );
  XNOR U2974 ( .A(y[163]), .B(x[163]), .Z(n2354) );
  XNOR U2975 ( .A(y[164]), .B(x[164]), .Z(n2353) );
  XNOR U2976 ( .A(n2345), .B(n2346), .Z(n2356) );
  XNOR U2977 ( .A(y[159]), .B(x[159]), .Z(n2346) );
  XNOR U2978 ( .A(n2347), .B(n2348), .Z(n2345) );
  XNOR U2979 ( .A(y[160]), .B(x[160]), .Z(n2348) );
  XNOR U2980 ( .A(y[161]), .B(x[161]), .Z(n2347) );
  NAND U2981 ( .A(n2412), .B(n2413), .Z(N2649) );
  NANDN U2982 ( .A(n2414), .B(n2415), .Z(n2413) );
  OR U2983 ( .A(n2416), .B(n2417), .Z(n2415) );
  NAND U2984 ( .A(n2416), .B(n2417), .Z(n2412) );
  XOR U2985 ( .A(n2416), .B(n2418), .Z(N2648) );
  XNOR U2986 ( .A(n2414), .B(n2417), .Z(n2418) );
  AND U2987 ( .A(n2419), .B(n2420), .Z(n2417) );
  NANDN U2988 ( .A(n2421), .B(n2422), .Z(n2420) );
  NANDN U2989 ( .A(n2423), .B(n2424), .Z(n2422) );
  NANDN U2990 ( .A(n2424), .B(n2423), .Z(n2419) );
  NAND U2991 ( .A(n2425), .B(n2426), .Z(n2414) );
  NANDN U2992 ( .A(n2427), .B(n2428), .Z(n2426) );
  OR U2993 ( .A(n2429), .B(n2430), .Z(n2428) );
  NAND U2994 ( .A(n2430), .B(n2429), .Z(n2425) );
  AND U2995 ( .A(n2431), .B(n2432), .Z(n2416) );
  NANDN U2996 ( .A(n2433), .B(n2434), .Z(n2432) );
  NANDN U2997 ( .A(n2435), .B(n2436), .Z(n2434) );
  NANDN U2998 ( .A(n2436), .B(n2435), .Z(n2431) );
  XOR U2999 ( .A(n2430), .B(n2437), .Z(N2647) );
  XOR U3000 ( .A(n2427), .B(n2429), .Z(n2437) );
  XNOR U3001 ( .A(n2423), .B(n2438), .Z(n2429) );
  XNOR U3002 ( .A(n2421), .B(n2424), .Z(n2438) );
  NAND U3003 ( .A(n2439), .B(n2440), .Z(n2424) );
  NAND U3004 ( .A(n2441), .B(n2442), .Z(n2440) );
  OR U3005 ( .A(n2443), .B(n2444), .Z(n2441) );
  NANDN U3006 ( .A(n2445), .B(n2443), .Z(n2439) );
  IV U3007 ( .A(n2444), .Z(n2445) );
  NAND U3008 ( .A(n2446), .B(n2447), .Z(n2421) );
  NAND U3009 ( .A(n2448), .B(n2449), .Z(n2447) );
  NANDN U3010 ( .A(n2450), .B(n2451), .Z(n2448) );
  NANDN U3011 ( .A(n2451), .B(n2450), .Z(n2446) );
  AND U3012 ( .A(n2452), .B(n2453), .Z(n2423) );
  NAND U3013 ( .A(n2454), .B(n2455), .Z(n2453) );
  OR U3014 ( .A(n2456), .B(n2457), .Z(n2454) );
  NANDN U3015 ( .A(n2458), .B(n2456), .Z(n2452) );
  NAND U3016 ( .A(n2459), .B(n2460), .Z(n2427) );
  NANDN U3017 ( .A(n2461), .B(n2462), .Z(n2460) );
  OR U3018 ( .A(n2463), .B(n2464), .Z(n2462) );
  NANDN U3019 ( .A(n2465), .B(n2463), .Z(n2459) );
  IV U3020 ( .A(n2464), .Z(n2465) );
  XNOR U3021 ( .A(n2435), .B(n2466), .Z(n2430) );
  XNOR U3022 ( .A(n2433), .B(n2436), .Z(n2466) );
  NAND U3023 ( .A(n2467), .B(n2468), .Z(n2436) );
  NAND U3024 ( .A(n2469), .B(n2470), .Z(n2468) );
  OR U3025 ( .A(n2471), .B(n2472), .Z(n2469) );
  NANDN U3026 ( .A(n2473), .B(n2471), .Z(n2467) );
  IV U3027 ( .A(n2472), .Z(n2473) );
  NAND U3028 ( .A(n2474), .B(n2475), .Z(n2433) );
  NAND U3029 ( .A(n2476), .B(n2477), .Z(n2475) );
  NANDN U3030 ( .A(n2478), .B(n2479), .Z(n2476) );
  NANDN U3031 ( .A(n2479), .B(n2478), .Z(n2474) );
  AND U3032 ( .A(n2480), .B(n2481), .Z(n2435) );
  NAND U3033 ( .A(n2482), .B(n2483), .Z(n2481) );
  OR U3034 ( .A(n2484), .B(n2485), .Z(n2482) );
  NANDN U3035 ( .A(n2486), .B(n2484), .Z(n2480) );
  XNOR U3036 ( .A(n2461), .B(n2487), .Z(N2646) );
  XOR U3037 ( .A(n2463), .B(n2464), .Z(n2487) );
  XNOR U3038 ( .A(n2477), .B(n2488), .Z(n2464) );
  XOR U3039 ( .A(n2478), .B(n2479), .Z(n2488) );
  XOR U3040 ( .A(n2484), .B(n2489), .Z(n2479) );
  XOR U3041 ( .A(n2483), .B(n2486), .Z(n2489) );
  IV U3042 ( .A(n2485), .Z(n2486) );
  NAND U3043 ( .A(n2490), .B(n2491), .Z(n2485) );
  OR U3044 ( .A(n2492), .B(n2493), .Z(n2491) );
  OR U3045 ( .A(n2494), .B(n2495), .Z(n2490) );
  NAND U3046 ( .A(n2496), .B(n2497), .Z(n2483) );
  OR U3047 ( .A(n2498), .B(n2499), .Z(n2497) );
  OR U3048 ( .A(n2500), .B(n2501), .Z(n2496) );
  NOR U3049 ( .A(n2502), .B(n2503), .Z(n2484) );
  ANDN U3050 ( .B(n2504), .A(n2505), .Z(n2478) );
  XNOR U3051 ( .A(n2471), .B(n2506), .Z(n2477) );
  XNOR U3052 ( .A(n2470), .B(n2472), .Z(n2506) );
  NAND U3053 ( .A(n2507), .B(n2508), .Z(n2472) );
  OR U3054 ( .A(n2509), .B(n2510), .Z(n2508) );
  OR U3055 ( .A(n2511), .B(n2512), .Z(n2507) );
  NAND U3056 ( .A(n2513), .B(n2514), .Z(n2470) );
  OR U3057 ( .A(n2515), .B(n2516), .Z(n2514) );
  OR U3058 ( .A(n2517), .B(n2518), .Z(n2513) );
  ANDN U3059 ( .B(n2519), .A(n2520), .Z(n2471) );
  IV U3060 ( .A(n2521), .Z(n2519) );
  ANDN U3061 ( .B(n2522), .A(n2523), .Z(n2463) );
  XOR U3062 ( .A(n2449), .B(n2524), .Z(n2461) );
  XOR U3063 ( .A(n2450), .B(n2451), .Z(n2524) );
  XOR U3064 ( .A(n2456), .B(n2525), .Z(n2451) );
  XOR U3065 ( .A(n2455), .B(n2458), .Z(n2525) );
  IV U3066 ( .A(n2457), .Z(n2458) );
  NAND U3067 ( .A(n2526), .B(n2527), .Z(n2457) );
  OR U3068 ( .A(n2528), .B(n2529), .Z(n2527) );
  OR U3069 ( .A(n2530), .B(n2531), .Z(n2526) );
  NAND U3070 ( .A(n2532), .B(n2533), .Z(n2455) );
  OR U3071 ( .A(n2534), .B(n2535), .Z(n2533) );
  OR U3072 ( .A(n2536), .B(n2537), .Z(n2532) );
  NOR U3073 ( .A(n2538), .B(n2539), .Z(n2456) );
  ANDN U3074 ( .B(n2540), .A(n2541), .Z(n2450) );
  IV U3075 ( .A(n2542), .Z(n2540) );
  XNOR U3076 ( .A(n2443), .B(n2543), .Z(n2449) );
  XNOR U3077 ( .A(n2442), .B(n2444), .Z(n2543) );
  NAND U3078 ( .A(n2544), .B(n2545), .Z(n2444) );
  OR U3079 ( .A(n2546), .B(n2547), .Z(n2545) );
  OR U3080 ( .A(n2548), .B(n2549), .Z(n2544) );
  NAND U3081 ( .A(n2550), .B(n2551), .Z(n2442) );
  OR U3082 ( .A(n2552), .B(n2553), .Z(n2551) );
  OR U3083 ( .A(n2554), .B(n2555), .Z(n2550) );
  ANDN U3084 ( .B(n2556), .A(n2557), .Z(n2443) );
  IV U3085 ( .A(n2558), .Z(n2556) );
  XNOR U3086 ( .A(n2523), .B(n2522), .Z(N2645) );
  XOR U3087 ( .A(n2542), .B(n2541), .Z(n2522) );
  XNOR U3088 ( .A(n2557), .B(n2558), .Z(n2541) );
  XNOR U3089 ( .A(n2552), .B(n2553), .Z(n2558) );
  XNOR U3090 ( .A(n2554), .B(n2555), .Z(n2553) );
  XNOR U3091 ( .A(y[157]), .B(x[157]), .Z(n2555) );
  XNOR U3092 ( .A(y[158]), .B(x[158]), .Z(n2554) );
  XNOR U3093 ( .A(y[156]), .B(x[156]), .Z(n2552) );
  XNOR U3094 ( .A(n2546), .B(n2547), .Z(n2557) );
  XNOR U3095 ( .A(y[153]), .B(x[153]), .Z(n2547) );
  XNOR U3096 ( .A(n2548), .B(n2549), .Z(n2546) );
  XNOR U3097 ( .A(y[154]), .B(x[154]), .Z(n2549) );
  XNOR U3098 ( .A(y[155]), .B(x[155]), .Z(n2548) );
  XNOR U3099 ( .A(n2539), .B(n2538), .Z(n2542) );
  XNOR U3100 ( .A(n2534), .B(n2535), .Z(n2538) );
  XNOR U3101 ( .A(y[150]), .B(x[150]), .Z(n2535) );
  XNOR U3102 ( .A(n2536), .B(n2537), .Z(n2534) );
  XNOR U3103 ( .A(y[151]), .B(x[151]), .Z(n2537) );
  XNOR U3104 ( .A(y[152]), .B(x[152]), .Z(n2536) );
  XNOR U3105 ( .A(n2528), .B(n2529), .Z(n2539) );
  XNOR U3106 ( .A(y[147]), .B(x[147]), .Z(n2529) );
  XNOR U3107 ( .A(n2530), .B(n2531), .Z(n2528) );
  XNOR U3108 ( .A(y[148]), .B(x[148]), .Z(n2531) );
  XNOR U3109 ( .A(y[149]), .B(x[149]), .Z(n2530) );
  XOR U3110 ( .A(n2504), .B(n2505), .Z(n2523) );
  XNOR U3111 ( .A(n2520), .B(n2521), .Z(n2505) );
  XNOR U3112 ( .A(n2515), .B(n2516), .Z(n2521) );
  XNOR U3113 ( .A(n2517), .B(n2518), .Z(n2516) );
  XNOR U3114 ( .A(y[145]), .B(x[145]), .Z(n2518) );
  XNOR U3115 ( .A(y[146]), .B(x[146]), .Z(n2517) );
  XNOR U3116 ( .A(y[144]), .B(x[144]), .Z(n2515) );
  XNOR U3117 ( .A(n2509), .B(n2510), .Z(n2520) );
  XNOR U3118 ( .A(y[141]), .B(x[141]), .Z(n2510) );
  XNOR U3119 ( .A(n2511), .B(n2512), .Z(n2509) );
  XNOR U3120 ( .A(y[142]), .B(x[142]), .Z(n2512) );
  XNOR U3121 ( .A(y[143]), .B(x[143]), .Z(n2511) );
  XOR U3122 ( .A(n2503), .B(n2502), .Z(n2504) );
  XNOR U3123 ( .A(n2498), .B(n2499), .Z(n2502) );
  XNOR U3124 ( .A(y[138]), .B(x[138]), .Z(n2499) );
  XNOR U3125 ( .A(n2500), .B(n2501), .Z(n2498) );
  XNOR U3126 ( .A(y[139]), .B(x[139]), .Z(n2501) );
  XNOR U3127 ( .A(y[140]), .B(x[140]), .Z(n2500) );
  XNOR U3128 ( .A(n2492), .B(n2493), .Z(n2503) );
  XNOR U3129 ( .A(y[135]), .B(x[135]), .Z(n2493) );
  XNOR U3130 ( .A(n2494), .B(n2495), .Z(n2492) );
  XNOR U3131 ( .A(y[136]), .B(x[136]), .Z(n2495) );
  XNOR U3132 ( .A(y[137]), .B(x[137]), .Z(n2494) );
  NAND U3133 ( .A(n2559), .B(n2560), .Z(N2640) );
  NANDN U3134 ( .A(n2561), .B(n2562), .Z(n2560) );
  OR U3135 ( .A(n2563), .B(n2564), .Z(n2562) );
  NAND U3136 ( .A(n2563), .B(n2564), .Z(n2559) );
  XOR U3137 ( .A(n2563), .B(n2565), .Z(N2639) );
  XNOR U3138 ( .A(n2561), .B(n2564), .Z(n2565) );
  AND U3139 ( .A(n2566), .B(n2567), .Z(n2564) );
  NANDN U3140 ( .A(n2568), .B(n2569), .Z(n2567) );
  NANDN U3141 ( .A(n2570), .B(n2571), .Z(n2569) );
  NANDN U3142 ( .A(n2571), .B(n2570), .Z(n2566) );
  NAND U3143 ( .A(n2572), .B(n2573), .Z(n2561) );
  NANDN U3144 ( .A(n2574), .B(n2575), .Z(n2573) );
  OR U3145 ( .A(n2576), .B(n2577), .Z(n2575) );
  NAND U3146 ( .A(n2577), .B(n2576), .Z(n2572) );
  AND U3147 ( .A(n2578), .B(n2579), .Z(n2563) );
  NANDN U3148 ( .A(n2580), .B(n2581), .Z(n2579) );
  NANDN U3149 ( .A(n2582), .B(n2583), .Z(n2581) );
  NANDN U3150 ( .A(n2583), .B(n2582), .Z(n2578) );
  XOR U3151 ( .A(n2577), .B(n2584), .Z(N2638) );
  XOR U3152 ( .A(n2574), .B(n2576), .Z(n2584) );
  XNOR U3153 ( .A(n2570), .B(n2585), .Z(n2576) );
  XNOR U3154 ( .A(n2568), .B(n2571), .Z(n2585) );
  NAND U3155 ( .A(n2586), .B(n2587), .Z(n2571) );
  NAND U3156 ( .A(n2588), .B(n2589), .Z(n2587) );
  OR U3157 ( .A(n2590), .B(n2591), .Z(n2588) );
  NANDN U3158 ( .A(n2592), .B(n2590), .Z(n2586) );
  IV U3159 ( .A(n2591), .Z(n2592) );
  NAND U3160 ( .A(n2593), .B(n2594), .Z(n2568) );
  NAND U3161 ( .A(n2595), .B(n2596), .Z(n2594) );
  NANDN U3162 ( .A(n2597), .B(n2598), .Z(n2595) );
  NANDN U3163 ( .A(n2598), .B(n2597), .Z(n2593) );
  AND U3164 ( .A(n2599), .B(n2600), .Z(n2570) );
  NAND U3165 ( .A(n2601), .B(n2602), .Z(n2600) );
  OR U3166 ( .A(n2603), .B(n2604), .Z(n2601) );
  NANDN U3167 ( .A(n2605), .B(n2603), .Z(n2599) );
  NAND U3168 ( .A(n2606), .B(n2607), .Z(n2574) );
  NANDN U3169 ( .A(n2608), .B(n2609), .Z(n2607) );
  OR U3170 ( .A(n2610), .B(n2611), .Z(n2609) );
  NANDN U3171 ( .A(n2612), .B(n2610), .Z(n2606) );
  IV U3172 ( .A(n2611), .Z(n2612) );
  XNOR U3173 ( .A(n2582), .B(n2613), .Z(n2577) );
  XNOR U3174 ( .A(n2580), .B(n2583), .Z(n2613) );
  NAND U3175 ( .A(n2614), .B(n2615), .Z(n2583) );
  NAND U3176 ( .A(n2616), .B(n2617), .Z(n2615) );
  OR U3177 ( .A(n2618), .B(n2619), .Z(n2616) );
  NANDN U3178 ( .A(n2620), .B(n2618), .Z(n2614) );
  IV U3179 ( .A(n2619), .Z(n2620) );
  NAND U3180 ( .A(n2621), .B(n2622), .Z(n2580) );
  NAND U3181 ( .A(n2623), .B(n2624), .Z(n2622) );
  NANDN U3182 ( .A(n2625), .B(n2626), .Z(n2623) );
  NANDN U3183 ( .A(n2626), .B(n2625), .Z(n2621) );
  AND U3184 ( .A(n2627), .B(n2628), .Z(n2582) );
  NAND U3185 ( .A(n2629), .B(n2630), .Z(n2628) );
  OR U3186 ( .A(n2631), .B(n2632), .Z(n2629) );
  NANDN U3187 ( .A(n2633), .B(n2631), .Z(n2627) );
  XNOR U3188 ( .A(n2608), .B(n2634), .Z(N2637) );
  XOR U3189 ( .A(n2610), .B(n2611), .Z(n2634) );
  XNOR U3190 ( .A(n2624), .B(n2635), .Z(n2611) );
  XOR U3191 ( .A(n2625), .B(n2626), .Z(n2635) );
  XOR U3192 ( .A(n2631), .B(n2636), .Z(n2626) );
  XOR U3193 ( .A(n2630), .B(n2633), .Z(n2636) );
  IV U3194 ( .A(n2632), .Z(n2633) );
  NAND U3195 ( .A(n2637), .B(n2638), .Z(n2632) );
  OR U3196 ( .A(n2639), .B(n2640), .Z(n2638) );
  OR U3197 ( .A(n2641), .B(n2642), .Z(n2637) );
  NAND U3198 ( .A(n2643), .B(n2644), .Z(n2630) );
  OR U3199 ( .A(n2645), .B(n2646), .Z(n2644) );
  OR U3200 ( .A(n2647), .B(n2648), .Z(n2643) );
  NOR U3201 ( .A(n2649), .B(n2650), .Z(n2631) );
  ANDN U3202 ( .B(n2651), .A(n2652), .Z(n2625) );
  XNOR U3203 ( .A(n2618), .B(n2653), .Z(n2624) );
  XNOR U3204 ( .A(n2617), .B(n2619), .Z(n2653) );
  NAND U3205 ( .A(n2654), .B(n2655), .Z(n2619) );
  OR U3206 ( .A(n2656), .B(n2657), .Z(n2655) );
  OR U3207 ( .A(n2658), .B(n2659), .Z(n2654) );
  NAND U3208 ( .A(n2660), .B(n2661), .Z(n2617) );
  OR U3209 ( .A(n2662), .B(n2663), .Z(n2661) );
  OR U3210 ( .A(n2664), .B(n2665), .Z(n2660) );
  ANDN U3211 ( .B(n2666), .A(n2667), .Z(n2618) );
  IV U3212 ( .A(n2668), .Z(n2666) );
  ANDN U3213 ( .B(n2669), .A(n2670), .Z(n2610) );
  XOR U3214 ( .A(n2596), .B(n2671), .Z(n2608) );
  XOR U3215 ( .A(n2597), .B(n2598), .Z(n2671) );
  XOR U3216 ( .A(n2603), .B(n2672), .Z(n2598) );
  XOR U3217 ( .A(n2602), .B(n2605), .Z(n2672) );
  IV U3218 ( .A(n2604), .Z(n2605) );
  NAND U3219 ( .A(n2673), .B(n2674), .Z(n2604) );
  OR U3220 ( .A(n2675), .B(n2676), .Z(n2674) );
  OR U3221 ( .A(n2677), .B(n2678), .Z(n2673) );
  NAND U3222 ( .A(n2679), .B(n2680), .Z(n2602) );
  OR U3223 ( .A(n2681), .B(n2682), .Z(n2680) );
  OR U3224 ( .A(n2683), .B(n2684), .Z(n2679) );
  NOR U3225 ( .A(n2685), .B(n2686), .Z(n2603) );
  ANDN U3226 ( .B(n2687), .A(n2688), .Z(n2597) );
  IV U3227 ( .A(n2689), .Z(n2687) );
  XNOR U3228 ( .A(n2590), .B(n2690), .Z(n2596) );
  XNOR U3229 ( .A(n2589), .B(n2591), .Z(n2690) );
  NAND U3230 ( .A(n2691), .B(n2692), .Z(n2591) );
  OR U3231 ( .A(n2693), .B(n2694), .Z(n2692) );
  OR U3232 ( .A(n2695), .B(n2696), .Z(n2691) );
  NAND U3233 ( .A(n2697), .B(n2698), .Z(n2589) );
  OR U3234 ( .A(n2699), .B(n2700), .Z(n2698) );
  OR U3235 ( .A(n2701), .B(n2702), .Z(n2697) );
  ANDN U3236 ( .B(n2703), .A(n2704), .Z(n2590) );
  IV U3237 ( .A(n2705), .Z(n2703) );
  XNOR U3238 ( .A(n2670), .B(n2669), .Z(N2636) );
  XOR U3239 ( .A(n2689), .B(n2688), .Z(n2669) );
  XNOR U3240 ( .A(n2704), .B(n2705), .Z(n2688) );
  XNOR U3241 ( .A(n2699), .B(n2700), .Z(n2705) );
  XNOR U3242 ( .A(n2701), .B(n2702), .Z(n2700) );
  XNOR U3243 ( .A(y[133]), .B(x[133]), .Z(n2702) );
  XNOR U3244 ( .A(y[134]), .B(x[134]), .Z(n2701) );
  XNOR U3245 ( .A(y[132]), .B(x[132]), .Z(n2699) );
  XNOR U3246 ( .A(n2693), .B(n2694), .Z(n2704) );
  XNOR U3247 ( .A(y[129]), .B(x[129]), .Z(n2694) );
  XNOR U3248 ( .A(n2695), .B(n2696), .Z(n2693) );
  XNOR U3249 ( .A(y[130]), .B(x[130]), .Z(n2696) );
  XNOR U3250 ( .A(y[131]), .B(x[131]), .Z(n2695) );
  XNOR U3251 ( .A(n2686), .B(n2685), .Z(n2689) );
  XNOR U3252 ( .A(n2681), .B(n2682), .Z(n2685) );
  XNOR U3253 ( .A(y[126]), .B(x[126]), .Z(n2682) );
  XNOR U3254 ( .A(n2683), .B(n2684), .Z(n2681) );
  XNOR U3255 ( .A(y[127]), .B(x[127]), .Z(n2684) );
  XNOR U3256 ( .A(y[128]), .B(x[128]), .Z(n2683) );
  XNOR U3257 ( .A(n2675), .B(n2676), .Z(n2686) );
  XNOR U3258 ( .A(y[123]), .B(x[123]), .Z(n2676) );
  XNOR U3259 ( .A(n2677), .B(n2678), .Z(n2675) );
  XNOR U3260 ( .A(y[124]), .B(x[124]), .Z(n2678) );
  XNOR U3261 ( .A(y[125]), .B(x[125]), .Z(n2677) );
  XOR U3262 ( .A(n2651), .B(n2652), .Z(n2670) );
  XNOR U3263 ( .A(n2667), .B(n2668), .Z(n2652) );
  XNOR U3264 ( .A(n2662), .B(n2663), .Z(n2668) );
  XNOR U3265 ( .A(n2664), .B(n2665), .Z(n2663) );
  XNOR U3266 ( .A(y[121]), .B(x[121]), .Z(n2665) );
  XNOR U3267 ( .A(y[122]), .B(x[122]), .Z(n2664) );
  XNOR U3268 ( .A(y[120]), .B(x[120]), .Z(n2662) );
  XNOR U3269 ( .A(n2656), .B(n2657), .Z(n2667) );
  XNOR U3270 ( .A(y[117]), .B(x[117]), .Z(n2657) );
  XNOR U3271 ( .A(n2658), .B(n2659), .Z(n2656) );
  XNOR U3272 ( .A(y[118]), .B(x[118]), .Z(n2659) );
  XNOR U3273 ( .A(y[119]), .B(x[119]), .Z(n2658) );
  XOR U3274 ( .A(n2650), .B(n2649), .Z(n2651) );
  XNOR U3275 ( .A(n2645), .B(n2646), .Z(n2649) );
  XNOR U3276 ( .A(y[114]), .B(x[114]), .Z(n2646) );
  XNOR U3277 ( .A(n2647), .B(n2648), .Z(n2645) );
  XNOR U3278 ( .A(y[115]), .B(x[115]), .Z(n2648) );
  XNOR U3279 ( .A(y[116]), .B(x[116]), .Z(n2647) );
  XNOR U3280 ( .A(n2639), .B(n2640), .Z(n2650) );
  XNOR U3281 ( .A(y[111]), .B(x[111]), .Z(n2640) );
  XNOR U3282 ( .A(n2641), .B(n2642), .Z(n2639) );
  XNOR U3283 ( .A(y[112]), .B(x[112]), .Z(n2642) );
  XNOR U3284 ( .A(y[113]), .B(x[113]), .Z(n2641) );
  NAND U3285 ( .A(n2706), .B(n2707), .Z(N2631) );
  NANDN U3286 ( .A(n2708), .B(n2709), .Z(n2707) );
  OR U3287 ( .A(n2710), .B(n2711), .Z(n2709) );
  NAND U3288 ( .A(n2710), .B(n2711), .Z(n2706) );
  XOR U3289 ( .A(n2710), .B(n2712), .Z(N2630) );
  XNOR U3290 ( .A(n2708), .B(n2711), .Z(n2712) );
  AND U3291 ( .A(n2713), .B(n2714), .Z(n2711) );
  NANDN U3292 ( .A(n2715), .B(n2716), .Z(n2714) );
  NANDN U3293 ( .A(n2717), .B(n2718), .Z(n2716) );
  NANDN U3294 ( .A(n2718), .B(n2717), .Z(n2713) );
  NAND U3295 ( .A(n2719), .B(n2720), .Z(n2708) );
  NANDN U3296 ( .A(n2721), .B(n2722), .Z(n2720) );
  OR U3297 ( .A(n2723), .B(n2724), .Z(n2722) );
  NAND U3298 ( .A(n2724), .B(n2723), .Z(n2719) );
  AND U3299 ( .A(n2725), .B(n2726), .Z(n2710) );
  NANDN U3300 ( .A(n2727), .B(n2728), .Z(n2726) );
  NANDN U3301 ( .A(n2729), .B(n2730), .Z(n2728) );
  NANDN U3302 ( .A(n2730), .B(n2729), .Z(n2725) );
  XOR U3303 ( .A(n2724), .B(n2731), .Z(N2629) );
  XOR U3304 ( .A(n2721), .B(n2723), .Z(n2731) );
  XNOR U3305 ( .A(n2717), .B(n2732), .Z(n2723) );
  XNOR U3306 ( .A(n2715), .B(n2718), .Z(n2732) );
  NAND U3307 ( .A(n2733), .B(n2734), .Z(n2718) );
  NAND U3308 ( .A(n2735), .B(n2736), .Z(n2734) );
  OR U3309 ( .A(n2737), .B(n2738), .Z(n2735) );
  NANDN U3310 ( .A(n2739), .B(n2737), .Z(n2733) );
  IV U3311 ( .A(n2738), .Z(n2739) );
  NAND U3312 ( .A(n2740), .B(n2741), .Z(n2715) );
  NAND U3313 ( .A(n2742), .B(n2743), .Z(n2741) );
  NANDN U3314 ( .A(n2744), .B(n2745), .Z(n2742) );
  NANDN U3315 ( .A(n2745), .B(n2744), .Z(n2740) );
  AND U3316 ( .A(n2746), .B(n2747), .Z(n2717) );
  NAND U3317 ( .A(n2748), .B(n2749), .Z(n2747) );
  OR U3318 ( .A(n2750), .B(n2751), .Z(n2748) );
  NANDN U3319 ( .A(n2752), .B(n2750), .Z(n2746) );
  NAND U3320 ( .A(n2753), .B(n2754), .Z(n2721) );
  NANDN U3321 ( .A(n2755), .B(n2756), .Z(n2754) );
  OR U3322 ( .A(n2757), .B(n2758), .Z(n2756) );
  NANDN U3323 ( .A(n2759), .B(n2757), .Z(n2753) );
  IV U3324 ( .A(n2758), .Z(n2759) );
  XNOR U3325 ( .A(n2729), .B(n2760), .Z(n2724) );
  XNOR U3326 ( .A(n2727), .B(n2730), .Z(n2760) );
  NAND U3327 ( .A(n2761), .B(n2762), .Z(n2730) );
  NAND U3328 ( .A(n2763), .B(n2764), .Z(n2762) );
  OR U3329 ( .A(n2765), .B(n2766), .Z(n2763) );
  NANDN U3330 ( .A(n2767), .B(n2765), .Z(n2761) );
  IV U3331 ( .A(n2766), .Z(n2767) );
  NAND U3332 ( .A(n2768), .B(n2769), .Z(n2727) );
  NAND U3333 ( .A(n2770), .B(n2771), .Z(n2769) );
  NANDN U3334 ( .A(n2772), .B(n2773), .Z(n2770) );
  NANDN U3335 ( .A(n2773), .B(n2772), .Z(n2768) );
  AND U3336 ( .A(n2774), .B(n2775), .Z(n2729) );
  NAND U3337 ( .A(n2776), .B(n2777), .Z(n2775) );
  OR U3338 ( .A(n2778), .B(n2779), .Z(n2776) );
  NANDN U3339 ( .A(n2780), .B(n2778), .Z(n2774) );
  XNOR U3340 ( .A(n2755), .B(n2781), .Z(N2628) );
  XOR U3341 ( .A(n2757), .B(n2758), .Z(n2781) );
  XNOR U3342 ( .A(n2771), .B(n2782), .Z(n2758) );
  XOR U3343 ( .A(n2772), .B(n2773), .Z(n2782) );
  XOR U3344 ( .A(n2778), .B(n2783), .Z(n2773) );
  XOR U3345 ( .A(n2777), .B(n2780), .Z(n2783) );
  IV U3346 ( .A(n2779), .Z(n2780) );
  NAND U3347 ( .A(n2784), .B(n2785), .Z(n2779) );
  OR U3348 ( .A(n2786), .B(n2787), .Z(n2785) );
  OR U3349 ( .A(n2788), .B(n2789), .Z(n2784) );
  NAND U3350 ( .A(n2790), .B(n2791), .Z(n2777) );
  OR U3351 ( .A(n2792), .B(n2793), .Z(n2791) );
  OR U3352 ( .A(n2794), .B(n2795), .Z(n2790) );
  NOR U3353 ( .A(n2796), .B(n2797), .Z(n2778) );
  ANDN U3354 ( .B(n2798), .A(n2799), .Z(n2772) );
  XNOR U3355 ( .A(n2765), .B(n2800), .Z(n2771) );
  XNOR U3356 ( .A(n2764), .B(n2766), .Z(n2800) );
  NAND U3357 ( .A(n2801), .B(n2802), .Z(n2766) );
  OR U3358 ( .A(n2803), .B(n2804), .Z(n2802) );
  OR U3359 ( .A(n2805), .B(n2806), .Z(n2801) );
  NAND U3360 ( .A(n2807), .B(n2808), .Z(n2764) );
  OR U3361 ( .A(n2809), .B(n2810), .Z(n2808) );
  OR U3362 ( .A(n2811), .B(n2812), .Z(n2807) );
  ANDN U3363 ( .B(n2813), .A(n2814), .Z(n2765) );
  IV U3364 ( .A(n2815), .Z(n2813) );
  ANDN U3365 ( .B(n2816), .A(n2817), .Z(n2757) );
  XOR U3366 ( .A(n2743), .B(n2818), .Z(n2755) );
  XOR U3367 ( .A(n2744), .B(n2745), .Z(n2818) );
  XOR U3368 ( .A(n2750), .B(n2819), .Z(n2745) );
  XOR U3369 ( .A(n2749), .B(n2752), .Z(n2819) );
  IV U3370 ( .A(n2751), .Z(n2752) );
  NAND U3371 ( .A(n2820), .B(n2821), .Z(n2751) );
  OR U3372 ( .A(n2822), .B(n2823), .Z(n2821) );
  OR U3373 ( .A(n2824), .B(n2825), .Z(n2820) );
  NAND U3374 ( .A(n2826), .B(n2827), .Z(n2749) );
  OR U3375 ( .A(n2828), .B(n2829), .Z(n2827) );
  OR U3376 ( .A(n2830), .B(n2831), .Z(n2826) );
  NOR U3377 ( .A(n2832), .B(n2833), .Z(n2750) );
  ANDN U3378 ( .B(n2834), .A(n2835), .Z(n2744) );
  IV U3379 ( .A(n2836), .Z(n2834) );
  XNOR U3380 ( .A(n2737), .B(n2837), .Z(n2743) );
  XNOR U3381 ( .A(n2736), .B(n2738), .Z(n2837) );
  NAND U3382 ( .A(n2838), .B(n2839), .Z(n2738) );
  OR U3383 ( .A(n2840), .B(n2841), .Z(n2839) );
  OR U3384 ( .A(n2842), .B(n2843), .Z(n2838) );
  NAND U3385 ( .A(n2844), .B(n2845), .Z(n2736) );
  OR U3386 ( .A(n2846), .B(n2847), .Z(n2845) );
  OR U3387 ( .A(n2848), .B(n2849), .Z(n2844) );
  ANDN U3388 ( .B(n2850), .A(n2851), .Z(n2737) );
  IV U3389 ( .A(n2852), .Z(n2850) );
  XNOR U3390 ( .A(n2817), .B(n2816), .Z(N2627) );
  XOR U3391 ( .A(n2836), .B(n2835), .Z(n2816) );
  XNOR U3392 ( .A(n2851), .B(n2852), .Z(n2835) );
  XNOR U3393 ( .A(n2846), .B(n2847), .Z(n2852) );
  XNOR U3394 ( .A(n2848), .B(n2849), .Z(n2847) );
  XNOR U3395 ( .A(y[109]), .B(x[109]), .Z(n2849) );
  XNOR U3396 ( .A(y[110]), .B(x[110]), .Z(n2848) );
  XNOR U3397 ( .A(y[108]), .B(x[108]), .Z(n2846) );
  XNOR U3398 ( .A(n2840), .B(n2841), .Z(n2851) );
  XNOR U3399 ( .A(y[105]), .B(x[105]), .Z(n2841) );
  XNOR U3400 ( .A(n2842), .B(n2843), .Z(n2840) );
  XNOR U3401 ( .A(y[106]), .B(x[106]), .Z(n2843) );
  XNOR U3402 ( .A(y[107]), .B(x[107]), .Z(n2842) );
  XNOR U3403 ( .A(n2833), .B(n2832), .Z(n2836) );
  XNOR U3404 ( .A(n2828), .B(n2829), .Z(n2832) );
  XNOR U3405 ( .A(y[102]), .B(x[102]), .Z(n2829) );
  XNOR U3406 ( .A(n2830), .B(n2831), .Z(n2828) );
  XNOR U3407 ( .A(y[103]), .B(x[103]), .Z(n2831) );
  XNOR U3408 ( .A(y[104]), .B(x[104]), .Z(n2830) );
  XNOR U3409 ( .A(n2822), .B(n2823), .Z(n2833) );
  XNOR U3410 ( .A(y[99]), .B(x[99]), .Z(n2823) );
  XNOR U3411 ( .A(n2824), .B(n2825), .Z(n2822) );
  XNOR U3412 ( .A(y[100]), .B(x[100]), .Z(n2825) );
  XNOR U3413 ( .A(y[101]), .B(x[101]), .Z(n2824) );
  XOR U3414 ( .A(n2798), .B(n2799), .Z(n2817) );
  XNOR U3415 ( .A(n2814), .B(n2815), .Z(n2799) );
  XNOR U3416 ( .A(n2809), .B(n2810), .Z(n2815) );
  XNOR U3417 ( .A(n2811), .B(n2812), .Z(n2810) );
  XNOR U3418 ( .A(y[97]), .B(x[97]), .Z(n2812) );
  XNOR U3419 ( .A(y[98]), .B(x[98]), .Z(n2811) );
  XNOR U3420 ( .A(y[96]), .B(x[96]), .Z(n2809) );
  XNOR U3421 ( .A(n2803), .B(n2804), .Z(n2814) );
  XNOR U3422 ( .A(y[93]), .B(x[93]), .Z(n2804) );
  XNOR U3423 ( .A(n2805), .B(n2806), .Z(n2803) );
  XNOR U3424 ( .A(y[94]), .B(x[94]), .Z(n2806) );
  XNOR U3425 ( .A(y[95]), .B(x[95]), .Z(n2805) );
  XOR U3426 ( .A(n2797), .B(n2796), .Z(n2798) );
  XNOR U3427 ( .A(n2792), .B(n2793), .Z(n2796) );
  XNOR U3428 ( .A(y[90]), .B(x[90]), .Z(n2793) );
  XNOR U3429 ( .A(n2794), .B(n2795), .Z(n2792) );
  XNOR U3430 ( .A(y[91]), .B(x[91]), .Z(n2795) );
  XNOR U3431 ( .A(y[92]), .B(x[92]), .Z(n2794) );
  XNOR U3432 ( .A(n2786), .B(n2787), .Z(n2797) );
  XNOR U3433 ( .A(y[87]), .B(x[87]), .Z(n2787) );
  XNOR U3434 ( .A(n2788), .B(n2789), .Z(n2786) );
  XNOR U3435 ( .A(y[88]), .B(x[88]), .Z(n2789) );
  XNOR U3436 ( .A(y[89]), .B(x[89]), .Z(n2788) );
  NAND U3437 ( .A(n2853), .B(n2854), .Z(N2622) );
  NANDN U3438 ( .A(n2855), .B(n2856), .Z(n2854) );
  OR U3439 ( .A(n2857), .B(n2858), .Z(n2856) );
  NAND U3440 ( .A(n2857), .B(n2858), .Z(n2853) );
  XOR U3441 ( .A(n2857), .B(n2859), .Z(N2621) );
  XNOR U3442 ( .A(n2855), .B(n2858), .Z(n2859) );
  AND U3443 ( .A(n2860), .B(n2861), .Z(n2858) );
  NANDN U3444 ( .A(n2862), .B(n2863), .Z(n2861) );
  NANDN U3445 ( .A(n2864), .B(n2865), .Z(n2863) );
  NANDN U3446 ( .A(n2865), .B(n2864), .Z(n2860) );
  NAND U3447 ( .A(n2866), .B(n2867), .Z(n2855) );
  NANDN U3448 ( .A(n2868), .B(n2869), .Z(n2867) );
  OR U3449 ( .A(n2870), .B(n2871), .Z(n2869) );
  NAND U3450 ( .A(n2871), .B(n2870), .Z(n2866) );
  AND U3451 ( .A(n2872), .B(n2873), .Z(n2857) );
  NANDN U3452 ( .A(n2874), .B(n2875), .Z(n2873) );
  NANDN U3453 ( .A(n2876), .B(n2877), .Z(n2875) );
  NANDN U3454 ( .A(n2877), .B(n2876), .Z(n2872) );
  XOR U3455 ( .A(n2871), .B(n2878), .Z(N2620) );
  XOR U3456 ( .A(n2868), .B(n2870), .Z(n2878) );
  XNOR U3457 ( .A(n2864), .B(n2879), .Z(n2870) );
  XNOR U3458 ( .A(n2862), .B(n2865), .Z(n2879) );
  NAND U3459 ( .A(n2880), .B(n2881), .Z(n2865) );
  NAND U3460 ( .A(n2882), .B(n2883), .Z(n2881) );
  OR U3461 ( .A(n2884), .B(n2885), .Z(n2882) );
  NANDN U3462 ( .A(n2886), .B(n2884), .Z(n2880) );
  IV U3463 ( .A(n2885), .Z(n2886) );
  NAND U3464 ( .A(n2887), .B(n2888), .Z(n2862) );
  NAND U3465 ( .A(n2889), .B(n2890), .Z(n2888) );
  NANDN U3466 ( .A(n2891), .B(n2892), .Z(n2889) );
  NANDN U3467 ( .A(n2892), .B(n2891), .Z(n2887) );
  AND U3468 ( .A(n2893), .B(n2894), .Z(n2864) );
  NAND U3469 ( .A(n2895), .B(n2896), .Z(n2894) );
  OR U3470 ( .A(n2897), .B(n2898), .Z(n2895) );
  NANDN U3471 ( .A(n2899), .B(n2897), .Z(n2893) );
  NAND U3472 ( .A(n2900), .B(n2901), .Z(n2868) );
  NANDN U3473 ( .A(n2902), .B(n2903), .Z(n2901) );
  OR U3474 ( .A(n2904), .B(n2905), .Z(n2903) );
  NANDN U3475 ( .A(n2906), .B(n2904), .Z(n2900) );
  IV U3476 ( .A(n2905), .Z(n2906) );
  XNOR U3477 ( .A(n2876), .B(n2907), .Z(n2871) );
  XNOR U3478 ( .A(n2874), .B(n2877), .Z(n2907) );
  NAND U3479 ( .A(n2908), .B(n2909), .Z(n2877) );
  NAND U3480 ( .A(n2910), .B(n2911), .Z(n2909) );
  OR U3481 ( .A(n2912), .B(n2913), .Z(n2910) );
  NANDN U3482 ( .A(n2914), .B(n2912), .Z(n2908) );
  IV U3483 ( .A(n2913), .Z(n2914) );
  NAND U3484 ( .A(n2915), .B(n2916), .Z(n2874) );
  NAND U3485 ( .A(n2917), .B(n2918), .Z(n2916) );
  NANDN U3486 ( .A(n2919), .B(n2920), .Z(n2917) );
  NANDN U3487 ( .A(n2920), .B(n2919), .Z(n2915) );
  AND U3488 ( .A(n2921), .B(n2922), .Z(n2876) );
  NAND U3489 ( .A(n2923), .B(n2924), .Z(n2922) );
  OR U3490 ( .A(n2925), .B(n2926), .Z(n2923) );
  NANDN U3491 ( .A(n2927), .B(n2925), .Z(n2921) );
  XNOR U3492 ( .A(n2902), .B(n2928), .Z(N2619) );
  XOR U3493 ( .A(n2904), .B(n2905), .Z(n2928) );
  XNOR U3494 ( .A(n2918), .B(n2929), .Z(n2905) );
  XOR U3495 ( .A(n2919), .B(n2920), .Z(n2929) );
  XOR U3496 ( .A(n2925), .B(n2930), .Z(n2920) );
  XOR U3497 ( .A(n2924), .B(n2927), .Z(n2930) );
  IV U3498 ( .A(n2926), .Z(n2927) );
  NAND U3499 ( .A(n2931), .B(n2932), .Z(n2926) );
  OR U3500 ( .A(n2933), .B(n2934), .Z(n2932) );
  OR U3501 ( .A(n2935), .B(n2936), .Z(n2931) );
  NAND U3502 ( .A(n2937), .B(n2938), .Z(n2924) );
  OR U3503 ( .A(n2939), .B(n2940), .Z(n2938) );
  OR U3504 ( .A(n2941), .B(n2942), .Z(n2937) );
  NOR U3505 ( .A(n2943), .B(n2944), .Z(n2925) );
  ANDN U3506 ( .B(n2945), .A(n2946), .Z(n2919) );
  XNOR U3507 ( .A(n2912), .B(n2947), .Z(n2918) );
  XNOR U3508 ( .A(n2911), .B(n2913), .Z(n2947) );
  NAND U3509 ( .A(n2948), .B(n2949), .Z(n2913) );
  OR U3510 ( .A(n2950), .B(n2951), .Z(n2949) );
  OR U3511 ( .A(n2952), .B(n2953), .Z(n2948) );
  NAND U3512 ( .A(n2954), .B(n2955), .Z(n2911) );
  OR U3513 ( .A(n2956), .B(n2957), .Z(n2955) );
  OR U3514 ( .A(n2958), .B(n2959), .Z(n2954) );
  ANDN U3515 ( .B(n2960), .A(n2961), .Z(n2912) );
  IV U3516 ( .A(n2962), .Z(n2960) );
  ANDN U3517 ( .B(n2963), .A(n2964), .Z(n2904) );
  XOR U3518 ( .A(n2890), .B(n2965), .Z(n2902) );
  XOR U3519 ( .A(n2891), .B(n2892), .Z(n2965) );
  XOR U3520 ( .A(n2897), .B(n2966), .Z(n2892) );
  XOR U3521 ( .A(n2896), .B(n2899), .Z(n2966) );
  IV U3522 ( .A(n2898), .Z(n2899) );
  NAND U3523 ( .A(n2967), .B(n2968), .Z(n2898) );
  OR U3524 ( .A(n2969), .B(n2970), .Z(n2968) );
  OR U3525 ( .A(n2971), .B(n2972), .Z(n2967) );
  NAND U3526 ( .A(n2973), .B(n2974), .Z(n2896) );
  OR U3527 ( .A(n2975), .B(n2976), .Z(n2974) );
  OR U3528 ( .A(n2977), .B(n2978), .Z(n2973) );
  NOR U3529 ( .A(n2979), .B(n2980), .Z(n2897) );
  ANDN U3530 ( .B(n2981), .A(n2982), .Z(n2891) );
  IV U3531 ( .A(n2983), .Z(n2981) );
  XNOR U3532 ( .A(n2884), .B(n2984), .Z(n2890) );
  XNOR U3533 ( .A(n2883), .B(n2885), .Z(n2984) );
  NAND U3534 ( .A(n2985), .B(n2986), .Z(n2885) );
  OR U3535 ( .A(n2987), .B(n2988), .Z(n2986) );
  OR U3536 ( .A(n2989), .B(n2990), .Z(n2985) );
  NAND U3537 ( .A(n2991), .B(n2992), .Z(n2883) );
  OR U3538 ( .A(n2993), .B(n2994), .Z(n2992) );
  OR U3539 ( .A(n2995), .B(n2996), .Z(n2991) );
  ANDN U3540 ( .B(n2997), .A(n2998), .Z(n2884) );
  IV U3541 ( .A(n2999), .Z(n2997) );
  XNOR U3542 ( .A(n2964), .B(n2963), .Z(N2618) );
  XOR U3543 ( .A(n2983), .B(n2982), .Z(n2963) );
  XNOR U3544 ( .A(n2998), .B(n2999), .Z(n2982) );
  XNOR U3545 ( .A(n2993), .B(n2994), .Z(n2999) );
  XNOR U3546 ( .A(n2995), .B(n2996), .Z(n2994) );
  XNOR U3547 ( .A(y[85]), .B(x[85]), .Z(n2996) );
  XNOR U3548 ( .A(y[86]), .B(x[86]), .Z(n2995) );
  XNOR U3549 ( .A(y[84]), .B(x[84]), .Z(n2993) );
  XNOR U3550 ( .A(n2987), .B(n2988), .Z(n2998) );
  XNOR U3551 ( .A(y[81]), .B(x[81]), .Z(n2988) );
  XNOR U3552 ( .A(n2989), .B(n2990), .Z(n2987) );
  XNOR U3553 ( .A(y[82]), .B(x[82]), .Z(n2990) );
  XNOR U3554 ( .A(y[83]), .B(x[83]), .Z(n2989) );
  XNOR U3555 ( .A(n2980), .B(n2979), .Z(n2983) );
  XNOR U3556 ( .A(n2975), .B(n2976), .Z(n2979) );
  XNOR U3557 ( .A(y[78]), .B(x[78]), .Z(n2976) );
  XNOR U3558 ( .A(n2977), .B(n2978), .Z(n2975) );
  XNOR U3559 ( .A(y[79]), .B(x[79]), .Z(n2978) );
  XNOR U3560 ( .A(y[80]), .B(x[80]), .Z(n2977) );
  XNOR U3561 ( .A(n2969), .B(n2970), .Z(n2980) );
  XNOR U3562 ( .A(y[75]), .B(x[75]), .Z(n2970) );
  XNOR U3563 ( .A(n2971), .B(n2972), .Z(n2969) );
  XNOR U3564 ( .A(y[76]), .B(x[76]), .Z(n2972) );
  XNOR U3565 ( .A(y[77]), .B(x[77]), .Z(n2971) );
  XOR U3566 ( .A(n2945), .B(n2946), .Z(n2964) );
  XNOR U3567 ( .A(n2961), .B(n2962), .Z(n2946) );
  XNOR U3568 ( .A(n2956), .B(n2957), .Z(n2962) );
  XNOR U3569 ( .A(n2958), .B(n2959), .Z(n2957) );
  XNOR U3570 ( .A(y[73]), .B(x[73]), .Z(n2959) );
  XNOR U3571 ( .A(y[74]), .B(x[74]), .Z(n2958) );
  XNOR U3572 ( .A(y[72]), .B(x[72]), .Z(n2956) );
  XNOR U3573 ( .A(n2950), .B(n2951), .Z(n2961) );
  XNOR U3574 ( .A(y[69]), .B(x[69]), .Z(n2951) );
  XNOR U3575 ( .A(n2952), .B(n2953), .Z(n2950) );
  XNOR U3576 ( .A(y[70]), .B(x[70]), .Z(n2953) );
  XNOR U3577 ( .A(y[71]), .B(x[71]), .Z(n2952) );
  XOR U3578 ( .A(n2944), .B(n2943), .Z(n2945) );
  XNOR U3579 ( .A(n2939), .B(n2940), .Z(n2943) );
  XNOR U3580 ( .A(y[66]), .B(x[66]), .Z(n2940) );
  XNOR U3581 ( .A(n2941), .B(n2942), .Z(n2939) );
  XNOR U3582 ( .A(y[67]), .B(x[67]), .Z(n2942) );
  XNOR U3583 ( .A(y[68]), .B(x[68]), .Z(n2941) );
  XNOR U3584 ( .A(n2933), .B(n2934), .Z(n2944) );
  XNOR U3585 ( .A(y[63]), .B(x[63]), .Z(n2934) );
  XNOR U3586 ( .A(n2935), .B(n2936), .Z(n2933) );
  XNOR U3587 ( .A(y[64]), .B(x[64]), .Z(n2936) );
  XNOR U3588 ( .A(y[65]), .B(x[65]), .Z(n2935) );
  NAND U3589 ( .A(n3000), .B(n3001), .Z(N2613) );
  NANDN U3590 ( .A(n3002), .B(n3003), .Z(n3001) );
  OR U3591 ( .A(n3004), .B(n3005), .Z(n3003) );
  NAND U3592 ( .A(n3004), .B(n3005), .Z(n3000) );
  XOR U3593 ( .A(n3004), .B(n3006), .Z(N2612) );
  XNOR U3594 ( .A(n3002), .B(n3005), .Z(n3006) );
  AND U3595 ( .A(n3007), .B(n3008), .Z(n3005) );
  NANDN U3596 ( .A(n3009), .B(n3010), .Z(n3008) );
  NANDN U3597 ( .A(n3011), .B(n3012), .Z(n3010) );
  NANDN U3598 ( .A(n3012), .B(n3011), .Z(n3007) );
  NAND U3599 ( .A(n3013), .B(n3014), .Z(n3002) );
  NANDN U3600 ( .A(n3015), .B(n3016), .Z(n3014) );
  OR U3601 ( .A(n3017), .B(n3018), .Z(n3016) );
  NAND U3602 ( .A(n3018), .B(n3017), .Z(n3013) );
  AND U3603 ( .A(n3019), .B(n3020), .Z(n3004) );
  NANDN U3604 ( .A(n3021), .B(n3022), .Z(n3020) );
  NANDN U3605 ( .A(n3023), .B(n3024), .Z(n3022) );
  NANDN U3606 ( .A(n3024), .B(n3023), .Z(n3019) );
  XOR U3607 ( .A(n3018), .B(n3025), .Z(N2611) );
  XOR U3608 ( .A(n3015), .B(n3017), .Z(n3025) );
  XNOR U3609 ( .A(n3011), .B(n3026), .Z(n3017) );
  XNOR U3610 ( .A(n3009), .B(n3012), .Z(n3026) );
  NAND U3611 ( .A(n3027), .B(n3028), .Z(n3012) );
  NAND U3612 ( .A(n3029), .B(n3030), .Z(n3028) );
  OR U3613 ( .A(n3031), .B(n3032), .Z(n3029) );
  NANDN U3614 ( .A(n3033), .B(n3031), .Z(n3027) );
  IV U3615 ( .A(n3032), .Z(n3033) );
  NAND U3616 ( .A(n3034), .B(n3035), .Z(n3009) );
  NAND U3617 ( .A(n3036), .B(n3037), .Z(n3035) );
  NANDN U3618 ( .A(n3038), .B(n3039), .Z(n3036) );
  NANDN U3619 ( .A(n3039), .B(n3038), .Z(n3034) );
  AND U3620 ( .A(n3040), .B(n3041), .Z(n3011) );
  NAND U3621 ( .A(n3042), .B(n3043), .Z(n3041) );
  OR U3622 ( .A(n3044), .B(n3045), .Z(n3042) );
  NANDN U3623 ( .A(n3046), .B(n3044), .Z(n3040) );
  NAND U3624 ( .A(n3047), .B(n3048), .Z(n3015) );
  NANDN U3625 ( .A(n3049), .B(n3050), .Z(n3048) );
  OR U3626 ( .A(n3051), .B(n3052), .Z(n3050) );
  NANDN U3627 ( .A(n3053), .B(n3051), .Z(n3047) );
  IV U3628 ( .A(n3052), .Z(n3053) );
  XNOR U3629 ( .A(n3023), .B(n3054), .Z(n3018) );
  XNOR U3630 ( .A(n3021), .B(n3024), .Z(n3054) );
  NAND U3631 ( .A(n3055), .B(n3056), .Z(n3024) );
  NAND U3632 ( .A(n3057), .B(n3058), .Z(n3056) );
  OR U3633 ( .A(n3059), .B(n3060), .Z(n3057) );
  NANDN U3634 ( .A(n3061), .B(n3059), .Z(n3055) );
  IV U3635 ( .A(n3060), .Z(n3061) );
  NAND U3636 ( .A(n3062), .B(n3063), .Z(n3021) );
  NAND U3637 ( .A(n3064), .B(n3065), .Z(n3063) );
  NANDN U3638 ( .A(n3066), .B(n3067), .Z(n3064) );
  NANDN U3639 ( .A(n3067), .B(n3066), .Z(n3062) );
  AND U3640 ( .A(n3068), .B(n3069), .Z(n3023) );
  NAND U3641 ( .A(n3070), .B(n3071), .Z(n3069) );
  OR U3642 ( .A(n3072), .B(n3073), .Z(n3070) );
  NANDN U3643 ( .A(n3074), .B(n3072), .Z(n3068) );
  XNOR U3644 ( .A(n3049), .B(n3075), .Z(N2610) );
  XOR U3645 ( .A(n3051), .B(n3052), .Z(n3075) );
  XNOR U3646 ( .A(n3065), .B(n3076), .Z(n3052) );
  XOR U3647 ( .A(n3066), .B(n3067), .Z(n3076) );
  XOR U3648 ( .A(n3072), .B(n3077), .Z(n3067) );
  XOR U3649 ( .A(n3071), .B(n3074), .Z(n3077) );
  IV U3650 ( .A(n3073), .Z(n3074) );
  NAND U3651 ( .A(n3078), .B(n3079), .Z(n3073) );
  OR U3652 ( .A(n3080), .B(n3081), .Z(n3079) );
  OR U3653 ( .A(n3082), .B(n3083), .Z(n3078) );
  NAND U3654 ( .A(n3084), .B(n3085), .Z(n3071) );
  OR U3655 ( .A(n3086), .B(n3087), .Z(n3085) );
  OR U3656 ( .A(n3088), .B(n3089), .Z(n3084) );
  NOR U3657 ( .A(n3090), .B(n3091), .Z(n3072) );
  ANDN U3658 ( .B(n3092), .A(n3093), .Z(n3066) );
  XNOR U3659 ( .A(n3059), .B(n3094), .Z(n3065) );
  XNOR U3660 ( .A(n3058), .B(n3060), .Z(n3094) );
  NAND U3661 ( .A(n3095), .B(n3096), .Z(n3060) );
  OR U3662 ( .A(n3097), .B(n3098), .Z(n3096) );
  OR U3663 ( .A(n3099), .B(n3100), .Z(n3095) );
  NAND U3664 ( .A(n3101), .B(n3102), .Z(n3058) );
  OR U3665 ( .A(n3103), .B(n3104), .Z(n3102) );
  OR U3666 ( .A(n3105), .B(n3106), .Z(n3101) );
  ANDN U3667 ( .B(n3107), .A(n3108), .Z(n3059) );
  IV U3668 ( .A(n3109), .Z(n3107) );
  ANDN U3669 ( .B(n3110), .A(n3111), .Z(n3051) );
  XOR U3670 ( .A(n3037), .B(n3112), .Z(n3049) );
  XOR U3671 ( .A(n3038), .B(n3039), .Z(n3112) );
  XOR U3672 ( .A(n3044), .B(n3113), .Z(n3039) );
  XOR U3673 ( .A(n3043), .B(n3046), .Z(n3113) );
  IV U3674 ( .A(n3045), .Z(n3046) );
  NAND U3675 ( .A(n3114), .B(n3115), .Z(n3045) );
  OR U3676 ( .A(n3116), .B(n3117), .Z(n3115) );
  OR U3677 ( .A(n3118), .B(n3119), .Z(n3114) );
  NAND U3678 ( .A(n3120), .B(n3121), .Z(n3043) );
  OR U3679 ( .A(n3122), .B(n3123), .Z(n3121) );
  OR U3680 ( .A(n3124), .B(n3125), .Z(n3120) );
  NOR U3681 ( .A(n3126), .B(n3127), .Z(n3044) );
  ANDN U3682 ( .B(n3128), .A(n3129), .Z(n3038) );
  IV U3683 ( .A(n3130), .Z(n3128) );
  XNOR U3684 ( .A(n3031), .B(n3131), .Z(n3037) );
  XNOR U3685 ( .A(n3030), .B(n3032), .Z(n3131) );
  NAND U3686 ( .A(n3132), .B(n3133), .Z(n3032) );
  OR U3687 ( .A(n3134), .B(n3135), .Z(n3133) );
  OR U3688 ( .A(n3136), .B(n3137), .Z(n3132) );
  NAND U3689 ( .A(n3138), .B(n3139), .Z(n3030) );
  OR U3690 ( .A(n3140), .B(n3141), .Z(n3139) );
  OR U3691 ( .A(n3142), .B(n3143), .Z(n3138) );
  ANDN U3692 ( .B(n3144), .A(n3145), .Z(n3031) );
  IV U3693 ( .A(n3146), .Z(n3144) );
  XNOR U3694 ( .A(n3111), .B(n3110), .Z(N2609) );
  XOR U3695 ( .A(n3130), .B(n3129), .Z(n3110) );
  XNOR U3696 ( .A(n3145), .B(n3146), .Z(n3129) );
  XNOR U3697 ( .A(n3140), .B(n3141), .Z(n3146) );
  XNOR U3698 ( .A(n3142), .B(n3143), .Z(n3141) );
  XNOR U3699 ( .A(y[61]), .B(x[61]), .Z(n3143) );
  XNOR U3700 ( .A(y[62]), .B(x[62]), .Z(n3142) );
  XNOR U3701 ( .A(y[60]), .B(x[60]), .Z(n3140) );
  XNOR U3702 ( .A(n3134), .B(n3135), .Z(n3145) );
  XNOR U3703 ( .A(y[57]), .B(x[57]), .Z(n3135) );
  XNOR U3704 ( .A(n3136), .B(n3137), .Z(n3134) );
  XNOR U3705 ( .A(y[58]), .B(x[58]), .Z(n3137) );
  XNOR U3706 ( .A(y[59]), .B(x[59]), .Z(n3136) );
  XNOR U3707 ( .A(n3127), .B(n3126), .Z(n3130) );
  XNOR U3708 ( .A(n3122), .B(n3123), .Z(n3126) );
  XNOR U3709 ( .A(y[54]), .B(x[54]), .Z(n3123) );
  XNOR U3710 ( .A(n3124), .B(n3125), .Z(n3122) );
  XNOR U3711 ( .A(y[55]), .B(x[55]), .Z(n3125) );
  XNOR U3712 ( .A(y[56]), .B(x[56]), .Z(n3124) );
  XNOR U3713 ( .A(n3116), .B(n3117), .Z(n3127) );
  XNOR U3714 ( .A(y[51]), .B(x[51]), .Z(n3117) );
  XNOR U3715 ( .A(n3118), .B(n3119), .Z(n3116) );
  XNOR U3716 ( .A(y[52]), .B(x[52]), .Z(n3119) );
  XNOR U3717 ( .A(y[53]), .B(x[53]), .Z(n3118) );
  XOR U3718 ( .A(n3092), .B(n3093), .Z(n3111) );
  XNOR U3719 ( .A(n3108), .B(n3109), .Z(n3093) );
  XNOR U3720 ( .A(n3103), .B(n3104), .Z(n3109) );
  XNOR U3721 ( .A(n3105), .B(n3106), .Z(n3104) );
  XNOR U3722 ( .A(y[49]), .B(x[49]), .Z(n3106) );
  XNOR U3723 ( .A(y[50]), .B(x[50]), .Z(n3105) );
  XNOR U3724 ( .A(y[48]), .B(x[48]), .Z(n3103) );
  XNOR U3725 ( .A(n3097), .B(n3098), .Z(n3108) );
  XNOR U3726 ( .A(y[45]), .B(x[45]), .Z(n3098) );
  XNOR U3727 ( .A(n3099), .B(n3100), .Z(n3097) );
  XNOR U3728 ( .A(y[46]), .B(x[46]), .Z(n3100) );
  XNOR U3729 ( .A(y[47]), .B(x[47]), .Z(n3099) );
  XOR U3730 ( .A(n3091), .B(n3090), .Z(n3092) );
  XNOR U3731 ( .A(n3086), .B(n3087), .Z(n3090) );
  XNOR U3732 ( .A(y[42]), .B(x[42]), .Z(n3087) );
  XNOR U3733 ( .A(n3088), .B(n3089), .Z(n3086) );
  XNOR U3734 ( .A(y[43]), .B(x[43]), .Z(n3089) );
  XNOR U3735 ( .A(y[44]), .B(x[44]), .Z(n3088) );
  XNOR U3736 ( .A(n3080), .B(n3081), .Z(n3091) );
  XNOR U3737 ( .A(y[39]), .B(x[39]), .Z(n3081) );
  XNOR U3738 ( .A(n3082), .B(n3083), .Z(n3080) );
  XNOR U3739 ( .A(y[40]), .B(x[40]), .Z(n3083) );
  XNOR U3740 ( .A(y[41]), .B(x[41]), .Z(n3082) );
  NAND U3741 ( .A(n3147), .B(n3148), .Z(N2604) );
  NANDN U3742 ( .A(n3149), .B(n3150), .Z(n3148) );
  OR U3743 ( .A(n3151), .B(n3152), .Z(n3150) );
  NAND U3744 ( .A(n3151), .B(n3152), .Z(n3147) );
  XOR U3745 ( .A(n3151), .B(n3153), .Z(N2603) );
  XNOR U3746 ( .A(n3149), .B(n3152), .Z(n3153) );
  AND U3747 ( .A(n3154), .B(n3155), .Z(n3152) );
  NANDN U3748 ( .A(n3156), .B(n3157), .Z(n3155) );
  NANDN U3749 ( .A(n3158), .B(n3159), .Z(n3157) );
  NANDN U3750 ( .A(n3159), .B(n3158), .Z(n3154) );
  NAND U3751 ( .A(n3160), .B(n3161), .Z(n3149) );
  NANDN U3752 ( .A(n3162), .B(n3163), .Z(n3161) );
  OR U3753 ( .A(n3164), .B(n3165), .Z(n3163) );
  NAND U3754 ( .A(n3165), .B(n3164), .Z(n3160) );
  AND U3755 ( .A(n3166), .B(n3167), .Z(n3151) );
  NANDN U3756 ( .A(n3168), .B(n3169), .Z(n3167) );
  NANDN U3757 ( .A(n3170), .B(n3171), .Z(n3169) );
  NANDN U3758 ( .A(n3171), .B(n3170), .Z(n3166) );
  XOR U3759 ( .A(n3165), .B(n3172), .Z(N2602) );
  XOR U3760 ( .A(n3162), .B(n3164), .Z(n3172) );
  XNOR U3761 ( .A(n3158), .B(n3173), .Z(n3164) );
  XNOR U3762 ( .A(n3156), .B(n3159), .Z(n3173) );
  NAND U3763 ( .A(n3174), .B(n3175), .Z(n3159) );
  NAND U3764 ( .A(n3176), .B(n3177), .Z(n3175) );
  OR U3765 ( .A(n3178), .B(n3179), .Z(n3176) );
  NANDN U3766 ( .A(n3180), .B(n3178), .Z(n3174) );
  IV U3767 ( .A(n3179), .Z(n3180) );
  NAND U3768 ( .A(n3181), .B(n3182), .Z(n3156) );
  NAND U3769 ( .A(n3183), .B(n3184), .Z(n3182) );
  NANDN U3770 ( .A(n3185), .B(n3186), .Z(n3183) );
  NANDN U3771 ( .A(n3186), .B(n3185), .Z(n3181) );
  AND U3772 ( .A(n3187), .B(n3188), .Z(n3158) );
  NAND U3773 ( .A(n3189), .B(n3190), .Z(n3188) );
  OR U3774 ( .A(n3191), .B(n3192), .Z(n3189) );
  NANDN U3775 ( .A(n3193), .B(n3191), .Z(n3187) );
  NAND U3776 ( .A(n3194), .B(n3195), .Z(n3162) );
  NANDN U3777 ( .A(n3196), .B(n3197), .Z(n3195) );
  OR U3778 ( .A(n3198), .B(n3199), .Z(n3197) );
  NANDN U3779 ( .A(n3200), .B(n3198), .Z(n3194) );
  IV U3780 ( .A(n3199), .Z(n3200) );
  XNOR U3781 ( .A(n3170), .B(n3201), .Z(n3165) );
  XNOR U3782 ( .A(n3168), .B(n3171), .Z(n3201) );
  NAND U3783 ( .A(n3202), .B(n3203), .Z(n3171) );
  NAND U3784 ( .A(n3204), .B(n3205), .Z(n3203) );
  OR U3785 ( .A(n3206), .B(n3207), .Z(n3204) );
  NANDN U3786 ( .A(n3208), .B(n3206), .Z(n3202) );
  IV U3787 ( .A(n3207), .Z(n3208) );
  NAND U3788 ( .A(n3209), .B(n3210), .Z(n3168) );
  NAND U3789 ( .A(n3211), .B(n3212), .Z(n3210) );
  NANDN U3790 ( .A(n3213), .B(n3214), .Z(n3211) );
  NANDN U3791 ( .A(n3214), .B(n3213), .Z(n3209) );
  AND U3792 ( .A(n3215), .B(n3216), .Z(n3170) );
  NAND U3793 ( .A(n3217), .B(n3218), .Z(n3216) );
  OR U3794 ( .A(n3219), .B(n3220), .Z(n3217) );
  NANDN U3795 ( .A(n3221), .B(n3219), .Z(n3215) );
  XNOR U3796 ( .A(n3196), .B(n3222), .Z(N2601) );
  XOR U3797 ( .A(n3198), .B(n3199), .Z(n3222) );
  XNOR U3798 ( .A(n3212), .B(n3223), .Z(n3199) );
  XOR U3799 ( .A(n3213), .B(n3214), .Z(n3223) );
  XOR U3800 ( .A(n3219), .B(n3224), .Z(n3214) );
  XOR U3801 ( .A(n3218), .B(n3221), .Z(n3224) );
  IV U3802 ( .A(n3220), .Z(n3221) );
  NAND U3803 ( .A(n3225), .B(n3226), .Z(n3220) );
  OR U3804 ( .A(n3227), .B(n3228), .Z(n3226) );
  OR U3805 ( .A(n3229), .B(n3230), .Z(n3225) );
  NAND U3806 ( .A(n3231), .B(n3232), .Z(n3218) );
  OR U3807 ( .A(n3233), .B(n3234), .Z(n3232) );
  OR U3808 ( .A(n3235), .B(n3236), .Z(n3231) );
  NOR U3809 ( .A(n3237), .B(n3238), .Z(n3219) );
  ANDN U3810 ( .B(n3239), .A(n3240), .Z(n3213) );
  XNOR U3811 ( .A(n3206), .B(n3241), .Z(n3212) );
  XNOR U3812 ( .A(n3205), .B(n3207), .Z(n3241) );
  NAND U3813 ( .A(n3242), .B(n3243), .Z(n3207) );
  OR U3814 ( .A(n3244), .B(n3245), .Z(n3243) );
  OR U3815 ( .A(n3246), .B(n3247), .Z(n3242) );
  NAND U3816 ( .A(n3248), .B(n3249), .Z(n3205) );
  OR U3817 ( .A(n3250), .B(n3251), .Z(n3249) );
  OR U3818 ( .A(n3252), .B(n3253), .Z(n3248) );
  ANDN U3819 ( .B(n3254), .A(n3255), .Z(n3206) );
  IV U3820 ( .A(n3256), .Z(n3254) );
  ANDN U3821 ( .B(n3257), .A(n3258), .Z(n3198) );
  XOR U3822 ( .A(n3184), .B(n3259), .Z(n3196) );
  XOR U3823 ( .A(n3185), .B(n3186), .Z(n3259) );
  XOR U3824 ( .A(n3191), .B(n3260), .Z(n3186) );
  XOR U3825 ( .A(n3190), .B(n3193), .Z(n3260) );
  IV U3826 ( .A(n3192), .Z(n3193) );
  NAND U3827 ( .A(n3261), .B(n3262), .Z(n3192) );
  OR U3828 ( .A(n3263), .B(n3264), .Z(n3262) );
  OR U3829 ( .A(n3265), .B(n3266), .Z(n3261) );
  NAND U3830 ( .A(n3267), .B(n3268), .Z(n3190) );
  OR U3831 ( .A(n3269), .B(n3270), .Z(n3268) );
  OR U3832 ( .A(n3271), .B(n3272), .Z(n3267) );
  NOR U3833 ( .A(n3273), .B(n3274), .Z(n3191) );
  ANDN U3834 ( .B(n3275), .A(n3276), .Z(n3185) );
  IV U3835 ( .A(n3277), .Z(n3275) );
  XNOR U3836 ( .A(n3178), .B(n3278), .Z(n3184) );
  XNOR U3837 ( .A(n3177), .B(n3179), .Z(n3278) );
  NAND U3838 ( .A(n3279), .B(n3280), .Z(n3179) );
  OR U3839 ( .A(n3281), .B(n3282), .Z(n3280) );
  OR U3840 ( .A(n3283), .B(n3284), .Z(n3279) );
  NAND U3841 ( .A(n3285), .B(n3286), .Z(n3177) );
  OR U3842 ( .A(n3287), .B(n3288), .Z(n3286) );
  OR U3843 ( .A(n3289), .B(n3290), .Z(n3285) );
  ANDN U3844 ( .B(n3291), .A(n3292), .Z(n3178) );
  IV U3845 ( .A(n3293), .Z(n3291) );
  XNOR U3846 ( .A(n3258), .B(n3257), .Z(N2600) );
  XOR U3847 ( .A(n3277), .B(n3276), .Z(n3257) );
  XNOR U3848 ( .A(n3292), .B(n3293), .Z(n3276) );
  XNOR U3849 ( .A(n3287), .B(n3288), .Z(n3293) );
  XNOR U3850 ( .A(n3289), .B(n3290), .Z(n3288) );
  XNOR U3851 ( .A(y[37]), .B(x[37]), .Z(n3290) );
  XNOR U3852 ( .A(y[38]), .B(x[38]), .Z(n3289) );
  XNOR U3853 ( .A(y[36]), .B(x[36]), .Z(n3287) );
  XNOR U3854 ( .A(n3281), .B(n3282), .Z(n3292) );
  XNOR U3855 ( .A(y[33]), .B(x[33]), .Z(n3282) );
  XNOR U3856 ( .A(n3283), .B(n3284), .Z(n3281) );
  XNOR U3857 ( .A(y[34]), .B(x[34]), .Z(n3284) );
  XNOR U3858 ( .A(y[35]), .B(x[35]), .Z(n3283) );
  XNOR U3859 ( .A(n3274), .B(n3273), .Z(n3277) );
  XNOR U3860 ( .A(n3269), .B(n3270), .Z(n3273) );
  XNOR U3861 ( .A(y[30]), .B(x[30]), .Z(n3270) );
  XNOR U3862 ( .A(n3271), .B(n3272), .Z(n3269) );
  XNOR U3863 ( .A(y[31]), .B(x[31]), .Z(n3272) );
  XNOR U3864 ( .A(y[32]), .B(x[32]), .Z(n3271) );
  XNOR U3865 ( .A(n3263), .B(n3264), .Z(n3274) );
  XNOR U3866 ( .A(y[27]), .B(x[27]), .Z(n3264) );
  XNOR U3867 ( .A(n3265), .B(n3266), .Z(n3263) );
  XNOR U3868 ( .A(y[28]), .B(x[28]), .Z(n3266) );
  XNOR U3869 ( .A(y[29]), .B(x[29]), .Z(n3265) );
  XOR U3870 ( .A(n3239), .B(n3240), .Z(n3258) );
  XNOR U3871 ( .A(n3255), .B(n3256), .Z(n3240) );
  XNOR U3872 ( .A(n3250), .B(n3251), .Z(n3256) );
  XNOR U3873 ( .A(n3252), .B(n3253), .Z(n3251) );
  XNOR U3874 ( .A(y[25]), .B(x[25]), .Z(n3253) );
  XNOR U3875 ( .A(y[26]), .B(x[26]), .Z(n3252) );
  XNOR U3876 ( .A(y[24]), .B(x[24]), .Z(n3250) );
  XNOR U3877 ( .A(n3244), .B(n3245), .Z(n3255) );
  XNOR U3878 ( .A(y[21]), .B(x[21]), .Z(n3245) );
  XNOR U3879 ( .A(n3246), .B(n3247), .Z(n3244) );
  XNOR U3880 ( .A(y[22]), .B(x[22]), .Z(n3247) );
  XNOR U3881 ( .A(y[23]), .B(x[23]), .Z(n3246) );
  XOR U3882 ( .A(n3238), .B(n3237), .Z(n3239) );
  XNOR U3883 ( .A(n3233), .B(n3234), .Z(n3237) );
  XNOR U3884 ( .A(y[18]), .B(x[18]), .Z(n3234) );
  XNOR U3885 ( .A(n3235), .B(n3236), .Z(n3233) );
  XNOR U3886 ( .A(y[19]), .B(x[19]), .Z(n3236) );
  XNOR U3887 ( .A(y[20]), .B(x[20]), .Z(n3235) );
  XNOR U3888 ( .A(n3227), .B(n3228), .Z(n3238) );
  XNOR U3889 ( .A(y[15]), .B(x[15]), .Z(n3228) );
  XNOR U3890 ( .A(n3229), .B(n3230), .Z(n3227) );
  XNOR U3891 ( .A(y[16]), .B(x[16]), .Z(n3230) );
  XNOR U3892 ( .A(y[17]), .B(x[17]), .Z(n3229) );
  NAND U3893 ( .A(n3294), .B(n3295), .Z(N2595) );
  OR U3894 ( .A(n3296), .B(n3297), .Z(n3295) );
  OR U3895 ( .A(n3297), .B(n3298), .Z(n3294) );
  XNOR U3896 ( .A(n3298), .B(n3299), .Z(N2594) );
  XOR U3897 ( .A(n3296), .B(n3297), .Z(n3299) );
  NAND U3898 ( .A(n3300), .B(n3301), .Z(n3297) );
  NANDN U3899 ( .A(n3302), .B(n3303), .Z(n3301) );
  NANDN U3900 ( .A(n3304), .B(n3305), .Z(n3303) );
  NANDN U3901 ( .A(n3305), .B(n3304), .Z(n3300) );
  NAND U3902 ( .A(n3306), .B(n3307), .Z(n3296) );
  NANDN U3903 ( .A(n3308), .B(n3309), .Z(n3307) );
  OR U3904 ( .A(n3310), .B(n3311), .Z(n3309) );
  NANDN U3905 ( .A(n3312), .B(n3310), .Z(n3306) );
  IV U3906 ( .A(n3311), .Z(n3312) );
  NANDN U3907 ( .A(n3313), .B(n3314), .Z(n3298) );
  XOR U3908 ( .A(n3311), .B(n3315), .Z(N2593) );
  XOR U3909 ( .A(n3308), .B(n3310), .Z(n3315) );
  XNOR U3910 ( .A(n3304), .B(n3316), .Z(n3310) );
  XNOR U3911 ( .A(n3302), .B(n3305), .Z(n3316) );
  NAND U3912 ( .A(n3317), .B(n3318), .Z(n3305) );
  NAND U3913 ( .A(n3319), .B(n3320), .Z(n3318) );
  OR U3914 ( .A(n3321), .B(n3322), .Z(n3319) );
  NANDN U3915 ( .A(n3323), .B(n3321), .Z(n3317) );
  IV U3916 ( .A(n3322), .Z(n3323) );
  NAND U3917 ( .A(n3324), .B(n3325), .Z(n3302) );
  NAND U3918 ( .A(n3326), .B(n3327), .Z(n3325) );
  NANDN U3919 ( .A(n3328), .B(n3329), .Z(n3326) );
  NANDN U3920 ( .A(n3329), .B(n3328), .Z(n3324) );
  AND U3921 ( .A(n3330), .B(n3331), .Z(n3304) );
  NAND U3922 ( .A(n3332), .B(n3333), .Z(n3331) );
  NANDN U3923 ( .A(n3334), .B(n3335), .Z(n3330) );
  NAND U3924 ( .A(n3336), .B(n3337), .Z(n3308) );
  NANDN U3925 ( .A(n3338), .B(n3339), .Z(n3337) );
  OR U3926 ( .A(n3340), .B(n3341), .Z(n3339) );
  NAND U3927 ( .A(n3341), .B(n3340), .Z(n3336) );
  XOR U3928 ( .A(n3314), .B(n3313), .Z(n3311) );
  NANDN U3929 ( .A(n3342), .B(n3343), .Z(n3313) );
  NAND U3930 ( .A(n3344), .B(n3345), .Z(n3314) );
  NAND U3931 ( .A(n3346), .B(n3347), .Z(n3345) );
  NAND U3932 ( .A(n3348), .B(n3349), .Z(n3346) );
  OR U3933 ( .A(n3348), .B(n3349), .Z(n3344) );
  XNOR U3934 ( .A(n3338), .B(n3350), .Z(N2592) );
  XOR U3935 ( .A(n3340), .B(n3341), .Z(n3350) );
  XOR U3936 ( .A(n3347), .B(n3351), .Z(n3341) );
  XOR U3937 ( .A(n3349), .B(n3348), .Z(n3351) );
  NANDN U3938 ( .A(n3352), .B(n3353), .Z(n3348) );
  AND U3939 ( .A(n3354), .B(n3355), .Z(n3349) );
  OR U3940 ( .A(n3356), .B(n3357), .Z(n3355) );
  OR U3941 ( .A(n3358), .B(n3359), .Z(n3354) );
  XNOR U3942 ( .A(n3343), .B(n3342), .Z(n3347) );
  AND U3943 ( .A(n3360), .B(n3361), .Z(n3342) );
  OR U3944 ( .A(n3362), .B(n3363), .Z(n3361) );
  OR U3945 ( .A(n3364), .B(n3365), .Z(n3360) );
  NAND U3946 ( .A(n3366), .B(n3367), .Z(n3343) );
  OR U3947 ( .A(n3368), .B(n3369), .Z(n3366) );
  IV U3948 ( .A(n3370), .Z(n3369) );
  ANDN U3949 ( .B(n3371), .A(n3372), .Z(n3340) );
  XOR U3950 ( .A(n3327), .B(n3373), .Z(n3338) );
  XOR U3951 ( .A(n3328), .B(n3329), .Z(n3373) );
  XNOR U3952 ( .A(n3332), .B(n3333), .Z(n3329) );
  XNOR U3953 ( .A(n3335), .B(n3334), .Z(n3333) );
  AND U3954 ( .A(n3374), .B(n3375), .Z(n3334) );
  NANDN U3955 ( .A(n3376), .B(n3377), .Z(n3375) );
  OR U3956 ( .A(n3378), .B(n3379), .Z(n3374) );
  IV U3957 ( .A(n3380), .Z(n3379) );
  NAND U3958 ( .A(n3381), .B(n3382), .Z(n3335) );
  NANDN U3959 ( .A(n3383), .B(n3384), .Z(n3382) );
  OR U3960 ( .A(n3385), .B(n3386), .Z(n3381) );
  IV U3961 ( .A(n3387), .Z(n3386) );
  ANDN U3962 ( .B(n3388), .A(n3389), .Z(n3332) );
  NOR U3963 ( .A(n3390), .B(n3391), .Z(n3328) );
  XNOR U3964 ( .A(n3321), .B(n3392), .Z(n3327) );
  XNOR U3965 ( .A(n3320), .B(n3322), .Z(n3392) );
  NAND U3966 ( .A(n3393), .B(n3394), .Z(n3322) );
  OR U3967 ( .A(n3395), .B(n3396), .Z(n3394) );
  OR U3968 ( .A(n3397), .B(n3398), .Z(n3393) );
  NAND U3969 ( .A(n3399), .B(n3400), .Z(n3320) );
  OR U3970 ( .A(n3401), .B(n3402), .Z(n3400) );
  OR U3971 ( .A(n3403), .B(n3404), .Z(n3399) );
  ANDN U3972 ( .B(n3405), .A(n3406), .Z(n3321) );
  IV U3973 ( .A(n3407), .Z(n3405) );
  XNOR U3974 ( .A(n3372), .B(n3371), .Z(N2591) );
  XOR U3975 ( .A(n3391), .B(n3390), .Z(n3371) );
  XNOR U3976 ( .A(n3406), .B(n3407), .Z(n3390) );
  XNOR U3977 ( .A(n3401), .B(n3402), .Z(n3407) );
  XNOR U3978 ( .A(n3403), .B(n3404), .Z(n3402) );
  XNOR U3979 ( .A(y[13]), .B(x[13]), .Z(n3404) );
  XNOR U3980 ( .A(y[14]), .B(x[14]), .Z(n3403) );
  XNOR U3981 ( .A(y[12]), .B(x[12]), .Z(n3401) );
  XNOR U3982 ( .A(n3395), .B(n3396), .Z(n3406) );
  XNOR U3983 ( .A(y[9]), .B(x[9]), .Z(n3396) );
  XNOR U3984 ( .A(n3397), .B(n3398), .Z(n3395) );
  XNOR U3985 ( .A(y[10]), .B(x[10]), .Z(n3398) );
  XNOR U3986 ( .A(y[11]), .B(x[11]), .Z(n3397) );
  XOR U3987 ( .A(n3388), .B(n3389), .Z(n3391) );
  XOR U3988 ( .A(n3376), .B(n3377), .Z(n3389) );
  XNOR U3989 ( .A(n3378), .B(n3380), .Z(n3377) );
  XOR U3990 ( .A(y[4]), .B(x[4]), .Z(n3380) );
  XNOR U3991 ( .A(y[5]), .B(x[5]), .Z(n3378) );
  XNOR U3992 ( .A(y[3]), .B(x[3]), .Z(n3376) );
  XNOR U3993 ( .A(n3383), .B(n3384), .Z(n3388) );
  XNOR U3994 ( .A(n3385), .B(n3387), .Z(n3384) );
  XOR U3995 ( .A(y[7]), .B(x[7]), .Z(n3387) );
  XNOR U3996 ( .A(y[8]), .B(x[8]), .Z(n3385) );
  XNOR U3997 ( .A(y[6]), .B(x[6]), .Z(n3383) );
  XOR U3998 ( .A(n3352), .B(n3353), .Z(n3372) );
  XNOR U3999 ( .A(n3368), .B(n3370), .Z(n3353) );
  XOR U4000 ( .A(y[498]), .B(x[498]), .Z(n3370) );
  NAND U4001 ( .A(n3408), .B(n3367), .Z(n3368) );
  OR U4002 ( .A(n3409), .B(n3410), .Z(n3367) );
  NAND U4003 ( .A(n3410), .B(n3409), .Z(n3408) );
  XNOR U4004 ( .A(y[499]), .B(x[499]), .Z(n3409) );
  XOR U4005 ( .A(n3411), .B(n3362), .Z(n3410) );
  XNOR U4006 ( .A(y[0]), .B(x[0]), .Z(n3362) );
  IV U4007 ( .A(n3363), .Z(n3411) );
  XNOR U4008 ( .A(n3365), .B(n3364), .Z(n3363) );
  XNOR U4009 ( .A(y[1]), .B(x[1]), .Z(n3364) );
  XNOR U4010 ( .A(y[2]), .B(x[2]), .Z(n3365) );
  XNOR U4011 ( .A(n3356), .B(n3357), .Z(n3352) );
  XNOR U4012 ( .A(y[495]), .B(x[495]), .Z(n3357) );
  XNOR U4013 ( .A(n3358), .B(n3359), .Z(n3356) );
  XNOR U4014 ( .A(y[496]), .B(x[496]), .Z(n3359) );
  XNOR U4015 ( .A(y[497]), .B(x[497]), .Z(n3358) );
endmodule

