
module mult_N256_CC64 ( clk, rst, a, b, c );
  input [255:0] a;
  input [3:0] b;
  output [511:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906;
  wire   [511:0] sreg;

  DFF \sreg_reg[507]  ( .D(c[511]), .CLK(clk), .RST(rst), .Q(sreg[507]) );
  DFF \sreg_reg[506]  ( .D(c[510]), .CLK(clk), .RST(rst), .Q(sreg[506]) );
  DFF \sreg_reg[505]  ( .D(c[509]), .CLK(clk), .RST(rst), .Q(sreg[505]) );
  DFF \sreg_reg[504]  ( .D(c[508]), .CLK(clk), .RST(rst), .Q(sreg[504]) );
  DFF \sreg_reg[503]  ( .D(c[507]), .CLK(clk), .RST(rst), .Q(sreg[503]) );
  DFF \sreg_reg[502]  ( .D(c[506]), .CLK(clk), .RST(rst), .Q(sreg[502]) );
  DFF \sreg_reg[501]  ( .D(c[505]), .CLK(clk), .RST(rst), .Q(sreg[501]) );
  DFF \sreg_reg[500]  ( .D(c[504]), .CLK(clk), .RST(rst), .Q(sreg[500]) );
  DFF \sreg_reg[499]  ( .D(c[503]), .CLK(clk), .RST(rst), .Q(sreg[499]) );
  DFF \sreg_reg[498]  ( .D(c[502]), .CLK(clk), .RST(rst), .Q(sreg[498]) );
  DFF \sreg_reg[497]  ( .D(c[501]), .CLK(clk), .RST(rst), .Q(sreg[497]) );
  DFF \sreg_reg[496]  ( .D(c[500]), .CLK(clk), .RST(rst), .Q(sreg[496]) );
  DFF \sreg_reg[495]  ( .D(c[499]), .CLK(clk), .RST(rst), .Q(sreg[495]) );
  DFF \sreg_reg[494]  ( .D(c[498]), .CLK(clk), .RST(rst), .Q(sreg[494]) );
  DFF \sreg_reg[493]  ( .D(c[497]), .CLK(clk), .RST(rst), .Q(sreg[493]) );
  DFF \sreg_reg[492]  ( .D(c[496]), .CLK(clk), .RST(rst), .Q(sreg[492]) );
  DFF \sreg_reg[491]  ( .D(c[495]), .CLK(clk), .RST(rst), .Q(sreg[491]) );
  DFF \sreg_reg[490]  ( .D(c[494]), .CLK(clk), .RST(rst), .Q(sreg[490]) );
  DFF \sreg_reg[489]  ( .D(c[493]), .CLK(clk), .RST(rst), .Q(sreg[489]) );
  DFF \sreg_reg[488]  ( .D(c[492]), .CLK(clk), .RST(rst), .Q(sreg[488]) );
  DFF \sreg_reg[487]  ( .D(c[491]), .CLK(clk), .RST(rst), .Q(sreg[487]) );
  DFF \sreg_reg[486]  ( .D(c[490]), .CLK(clk), .RST(rst), .Q(sreg[486]) );
  DFF \sreg_reg[485]  ( .D(c[489]), .CLK(clk), .RST(rst), .Q(sreg[485]) );
  DFF \sreg_reg[484]  ( .D(c[488]), .CLK(clk), .RST(rst), .Q(sreg[484]) );
  DFF \sreg_reg[483]  ( .D(c[487]), .CLK(clk), .RST(rst), .Q(sreg[483]) );
  DFF \sreg_reg[482]  ( .D(c[486]), .CLK(clk), .RST(rst), .Q(sreg[482]) );
  DFF \sreg_reg[481]  ( .D(c[485]), .CLK(clk), .RST(rst), .Q(sreg[481]) );
  DFF \sreg_reg[480]  ( .D(c[484]), .CLK(clk), .RST(rst), .Q(sreg[480]) );
  DFF \sreg_reg[479]  ( .D(c[483]), .CLK(clk), .RST(rst), .Q(sreg[479]) );
  DFF \sreg_reg[478]  ( .D(c[482]), .CLK(clk), .RST(rst), .Q(sreg[478]) );
  DFF \sreg_reg[477]  ( .D(c[481]), .CLK(clk), .RST(rst), .Q(sreg[477]) );
  DFF \sreg_reg[476]  ( .D(c[480]), .CLK(clk), .RST(rst), .Q(sreg[476]) );
  DFF \sreg_reg[475]  ( .D(c[479]), .CLK(clk), .RST(rst), .Q(sreg[475]) );
  DFF \sreg_reg[474]  ( .D(c[478]), .CLK(clk), .RST(rst), .Q(sreg[474]) );
  DFF \sreg_reg[473]  ( .D(c[477]), .CLK(clk), .RST(rst), .Q(sreg[473]) );
  DFF \sreg_reg[472]  ( .D(c[476]), .CLK(clk), .RST(rst), .Q(sreg[472]) );
  DFF \sreg_reg[471]  ( .D(c[475]), .CLK(clk), .RST(rst), .Q(sreg[471]) );
  DFF \sreg_reg[470]  ( .D(c[474]), .CLK(clk), .RST(rst), .Q(sreg[470]) );
  DFF \sreg_reg[469]  ( .D(c[473]), .CLK(clk), .RST(rst), .Q(sreg[469]) );
  DFF \sreg_reg[468]  ( .D(c[472]), .CLK(clk), .RST(rst), .Q(sreg[468]) );
  DFF \sreg_reg[467]  ( .D(c[471]), .CLK(clk), .RST(rst), .Q(sreg[467]) );
  DFF \sreg_reg[466]  ( .D(c[470]), .CLK(clk), .RST(rst), .Q(sreg[466]) );
  DFF \sreg_reg[465]  ( .D(c[469]), .CLK(clk), .RST(rst), .Q(sreg[465]) );
  DFF \sreg_reg[464]  ( .D(c[468]), .CLK(clk), .RST(rst), .Q(sreg[464]) );
  DFF \sreg_reg[463]  ( .D(c[467]), .CLK(clk), .RST(rst), .Q(sreg[463]) );
  DFF \sreg_reg[462]  ( .D(c[466]), .CLK(clk), .RST(rst), .Q(sreg[462]) );
  DFF \sreg_reg[461]  ( .D(c[465]), .CLK(clk), .RST(rst), .Q(sreg[461]) );
  DFF \sreg_reg[460]  ( .D(c[464]), .CLK(clk), .RST(rst), .Q(sreg[460]) );
  DFF \sreg_reg[459]  ( .D(c[463]), .CLK(clk), .RST(rst), .Q(sreg[459]) );
  DFF \sreg_reg[458]  ( .D(c[462]), .CLK(clk), .RST(rst), .Q(sreg[458]) );
  DFF \sreg_reg[457]  ( .D(c[461]), .CLK(clk), .RST(rst), .Q(sreg[457]) );
  DFF \sreg_reg[456]  ( .D(c[460]), .CLK(clk), .RST(rst), .Q(sreg[456]) );
  DFF \sreg_reg[455]  ( .D(c[459]), .CLK(clk), .RST(rst), .Q(sreg[455]) );
  DFF \sreg_reg[454]  ( .D(c[458]), .CLK(clk), .RST(rst), .Q(sreg[454]) );
  DFF \sreg_reg[453]  ( .D(c[457]), .CLK(clk), .RST(rst), .Q(sreg[453]) );
  DFF \sreg_reg[452]  ( .D(c[456]), .CLK(clk), .RST(rst), .Q(sreg[452]) );
  DFF \sreg_reg[451]  ( .D(c[455]), .CLK(clk), .RST(rst), .Q(sreg[451]) );
  DFF \sreg_reg[450]  ( .D(c[454]), .CLK(clk), .RST(rst), .Q(sreg[450]) );
  DFF \sreg_reg[449]  ( .D(c[453]), .CLK(clk), .RST(rst), .Q(sreg[449]) );
  DFF \sreg_reg[448]  ( .D(c[452]), .CLK(clk), .RST(rst), .Q(sreg[448]) );
  DFF \sreg_reg[447]  ( .D(c[451]), .CLK(clk), .RST(rst), .Q(sreg[447]) );
  DFF \sreg_reg[446]  ( .D(c[450]), .CLK(clk), .RST(rst), .Q(sreg[446]) );
  DFF \sreg_reg[445]  ( .D(c[449]), .CLK(clk), .RST(rst), .Q(sreg[445]) );
  DFF \sreg_reg[444]  ( .D(c[448]), .CLK(clk), .RST(rst), .Q(sreg[444]) );
  DFF \sreg_reg[443]  ( .D(c[447]), .CLK(clk), .RST(rst), .Q(sreg[443]) );
  DFF \sreg_reg[442]  ( .D(c[446]), .CLK(clk), .RST(rst), .Q(sreg[442]) );
  DFF \sreg_reg[441]  ( .D(c[445]), .CLK(clk), .RST(rst), .Q(sreg[441]) );
  DFF \sreg_reg[440]  ( .D(c[444]), .CLK(clk), .RST(rst), .Q(sreg[440]) );
  DFF \sreg_reg[439]  ( .D(c[443]), .CLK(clk), .RST(rst), .Q(sreg[439]) );
  DFF \sreg_reg[438]  ( .D(c[442]), .CLK(clk), .RST(rst), .Q(sreg[438]) );
  DFF \sreg_reg[437]  ( .D(c[441]), .CLK(clk), .RST(rst), .Q(sreg[437]) );
  DFF \sreg_reg[436]  ( .D(c[440]), .CLK(clk), .RST(rst), .Q(sreg[436]) );
  DFF \sreg_reg[435]  ( .D(c[439]), .CLK(clk), .RST(rst), .Q(sreg[435]) );
  DFF \sreg_reg[434]  ( .D(c[438]), .CLK(clk), .RST(rst), .Q(sreg[434]) );
  DFF \sreg_reg[433]  ( .D(c[437]), .CLK(clk), .RST(rst), .Q(sreg[433]) );
  DFF \sreg_reg[432]  ( .D(c[436]), .CLK(clk), .RST(rst), .Q(sreg[432]) );
  DFF \sreg_reg[431]  ( .D(c[435]), .CLK(clk), .RST(rst), .Q(sreg[431]) );
  DFF \sreg_reg[430]  ( .D(c[434]), .CLK(clk), .RST(rst), .Q(sreg[430]) );
  DFF \sreg_reg[429]  ( .D(c[433]), .CLK(clk), .RST(rst), .Q(sreg[429]) );
  DFF \sreg_reg[428]  ( .D(c[432]), .CLK(clk), .RST(rst), .Q(sreg[428]) );
  DFF \sreg_reg[427]  ( .D(c[431]), .CLK(clk), .RST(rst), .Q(sreg[427]) );
  DFF \sreg_reg[426]  ( .D(c[430]), .CLK(clk), .RST(rst), .Q(sreg[426]) );
  DFF \sreg_reg[425]  ( .D(c[429]), .CLK(clk), .RST(rst), .Q(sreg[425]) );
  DFF \sreg_reg[424]  ( .D(c[428]), .CLK(clk), .RST(rst), .Q(sreg[424]) );
  DFF \sreg_reg[423]  ( .D(c[427]), .CLK(clk), .RST(rst), .Q(sreg[423]) );
  DFF \sreg_reg[422]  ( .D(c[426]), .CLK(clk), .RST(rst), .Q(sreg[422]) );
  DFF \sreg_reg[421]  ( .D(c[425]), .CLK(clk), .RST(rst), .Q(sreg[421]) );
  DFF \sreg_reg[420]  ( .D(c[424]), .CLK(clk), .RST(rst), .Q(sreg[420]) );
  DFF \sreg_reg[419]  ( .D(c[423]), .CLK(clk), .RST(rst), .Q(sreg[419]) );
  DFF \sreg_reg[418]  ( .D(c[422]), .CLK(clk), .RST(rst), .Q(sreg[418]) );
  DFF \sreg_reg[417]  ( .D(c[421]), .CLK(clk), .RST(rst), .Q(sreg[417]) );
  DFF \sreg_reg[416]  ( .D(c[420]), .CLK(clk), .RST(rst), .Q(sreg[416]) );
  DFF \sreg_reg[415]  ( .D(c[419]), .CLK(clk), .RST(rst), .Q(sreg[415]) );
  DFF \sreg_reg[414]  ( .D(c[418]), .CLK(clk), .RST(rst), .Q(sreg[414]) );
  DFF \sreg_reg[413]  ( .D(c[417]), .CLK(clk), .RST(rst), .Q(sreg[413]) );
  DFF \sreg_reg[412]  ( .D(c[416]), .CLK(clk), .RST(rst), .Q(sreg[412]) );
  DFF \sreg_reg[411]  ( .D(c[415]), .CLK(clk), .RST(rst), .Q(sreg[411]) );
  DFF \sreg_reg[410]  ( .D(c[414]), .CLK(clk), .RST(rst), .Q(sreg[410]) );
  DFF \sreg_reg[409]  ( .D(c[413]), .CLK(clk), .RST(rst), .Q(sreg[409]) );
  DFF \sreg_reg[408]  ( .D(c[412]), .CLK(clk), .RST(rst), .Q(sreg[408]) );
  DFF \sreg_reg[407]  ( .D(c[411]), .CLK(clk), .RST(rst), .Q(sreg[407]) );
  DFF \sreg_reg[406]  ( .D(c[410]), .CLK(clk), .RST(rst), .Q(sreg[406]) );
  DFF \sreg_reg[405]  ( .D(c[409]), .CLK(clk), .RST(rst), .Q(sreg[405]) );
  DFF \sreg_reg[404]  ( .D(c[408]), .CLK(clk), .RST(rst), .Q(sreg[404]) );
  DFF \sreg_reg[403]  ( .D(c[407]), .CLK(clk), .RST(rst), .Q(sreg[403]) );
  DFF \sreg_reg[402]  ( .D(c[406]), .CLK(clk), .RST(rst), .Q(sreg[402]) );
  DFF \sreg_reg[401]  ( .D(c[405]), .CLK(clk), .RST(rst), .Q(sreg[401]) );
  DFF \sreg_reg[400]  ( .D(c[404]), .CLK(clk), .RST(rst), .Q(sreg[400]) );
  DFF \sreg_reg[399]  ( .D(c[403]), .CLK(clk), .RST(rst), .Q(sreg[399]) );
  DFF \sreg_reg[398]  ( .D(c[402]), .CLK(clk), .RST(rst), .Q(sreg[398]) );
  DFF \sreg_reg[397]  ( .D(c[401]), .CLK(clk), .RST(rst), .Q(sreg[397]) );
  DFF \sreg_reg[396]  ( .D(c[400]), .CLK(clk), .RST(rst), .Q(sreg[396]) );
  DFF \sreg_reg[395]  ( .D(c[399]), .CLK(clk), .RST(rst), .Q(sreg[395]) );
  DFF \sreg_reg[394]  ( .D(c[398]), .CLK(clk), .RST(rst), .Q(sreg[394]) );
  DFF \sreg_reg[393]  ( .D(c[397]), .CLK(clk), .RST(rst), .Q(sreg[393]) );
  DFF \sreg_reg[392]  ( .D(c[396]), .CLK(clk), .RST(rst), .Q(sreg[392]) );
  DFF \sreg_reg[391]  ( .D(c[395]), .CLK(clk), .RST(rst), .Q(sreg[391]) );
  DFF \sreg_reg[390]  ( .D(c[394]), .CLK(clk), .RST(rst), .Q(sreg[390]) );
  DFF \sreg_reg[389]  ( .D(c[393]), .CLK(clk), .RST(rst), .Q(sreg[389]) );
  DFF \sreg_reg[388]  ( .D(c[392]), .CLK(clk), .RST(rst), .Q(sreg[388]) );
  DFF \sreg_reg[387]  ( .D(c[391]), .CLK(clk), .RST(rst), .Q(sreg[387]) );
  DFF \sreg_reg[386]  ( .D(c[390]), .CLK(clk), .RST(rst), .Q(sreg[386]) );
  DFF \sreg_reg[385]  ( .D(c[389]), .CLK(clk), .RST(rst), .Q(sreg[385]) );
  DFF \sreg_reg[384]  ( .D(c[388]), .CLK(clk), .RST(rst), .Q(sreg[384]) );
  DFF \sreg_reg[383]  ( .D(c[387]), .CLK(clk), .RST(rst), .Q(sreg[383]) );
  DFF \sreg_reg[382]  ( .D(c[386]), .CLK(clk), .RST(rst), .Q(sreg[382]) );
  DFF \sreg_reg[381]  ( .D(c[385]), .CLK(clk), .RST(rst), .Q(sreg[381]) );
  DFF \sreg_reg[380]  ( .D(c[384]), .CLK(clk), .RST(rst), .Q(sreg[380]) );
  DFF \sreg_reg[379]  ( .D(c[383]), .CLK(clk), .RST(rst), .Q(sreg[379]) );
  DFF \sreg_reg[378]  ( .D(c[382]), .CLK(clk), .RST(rst), .Q(sreg[378]) );
  DFF \sreg_reg[377]  ( .D(c[381]), .CLK(clk), .RST(rst), .Q(sreg[377]) );
  DFF \sreg_reg[376]  ( .D(c[380]), .CLK(clk), .RST(rst), .Q(sreg[376]) );
  DFF \sreg_reg[375]  ( .D(c[379]), .CLK(clk), .RST(rst), .Q(sreg[375]) );
  DFF \sreg_reg[374]  ( .D(c[378]), .CLK(clk), .RST(rst), .Q(sreg[374]) );
  DFF \sreg_reg[373]  ( .D(c[377]), .CLK(clk), .RST(rst), .Q(sreg[373]) );
  DFF \sreg_reg[372]  ( .D(c[376]), .CLK(clk), .RST(rst), .Q(sreg[372]) );
  DFF \sreg_reg[371]  ( .D(c[375]), .CLK(clk), .RST(rst), .Q(sreg[371]) );
  DFF \sreg_reg[370]  ( .D(c[374]), .CLK(clk), .RST(rst), .Q(sreg[370]) );
  DFF \sreg_reg[369]  ( .D(c[373]), .CLK(clk), .RST(rst), .Q(sreg[369]) );
  DFF \sreg_reg[368]  ( .D(c[372]), .CLK(clk), .RST(rst), .Q(sreg[368]) );
  DFF \sreg_reg[367]  ( .D(c[371]), .CLK(clk), .RST(rst), .Q(sreg[367]) );
  DFF \sreg_reg[366]  ( .D(c[370]), .CLK(clk), .RST(rst), .Q(sreg[366]) );
  DFF \sreg_reg[365]  ( .D(c[369]), .CLK(clk), .RST(rst), .Q(sreg[365]) );
  DFF \sreg_reg[364]  ( .D(c[368]), .CLK(clk), .RST(rst), .Q(sreg[364]) );
  DFF \sreg_reg[363]  ( .D(c[367]), .CLK(clk), .RST(rst), .Q(sreg[363]) );
  DFF \sreg_reg[362]  ( .D(c[366]), .CLK(clk), .RST(rst), .Q(sreg[362]) );
  DFF \sreg_reg[361]  ( .D(c[365]), .CLK(clk), .RST(rst), .Q(sreg[361]) );
  DFF \sreg_reg[360]  ( .D(c[364]), .CLK(clk), .RST(rst), .Q(sreg[360]) );
  DFF \sreg_reg[359]  ( .D(c[363]), .CLK(clk), .RST(rst), .Q(sreg[359]) );
  DFF \sreg_reg[358]  ( .D(c[362]), .CLK(clk), .RST(rst), .Q(sreg[358]) );
  DFF \sreg_reg[357]  ( .D(c[361]), .CLK(clk), .RST(rst), .Q(sreg[357]) );
  DFF \sreg_reg[356]  ( .D(c[360]), .CLK(clk), .RST(rst), .Q(sreg[356]) );
  DFF \sreg_reg[355]  ( .D(c[359]), .CLK(clk), .RST(rst), .Q(sreg[355]) );
  DFF \sreg_reg[354]  ( .D(c[358]), .CLK(clk), .RST(rst), .Q(sreg[354]) );
  DFF \sreg_reg[353]  ( .D(c[357]), .CLK(clk), .RST(rst), .Q(sreg[353]) );
  DFF \sreg_reg[352]  ( .D(c[356]), .CLK(clk), .RST(rst), .Q(sreg[352]) );
  DFF \sreg_reg[351]  ( .D(c[355]), .CLK(clk), .RST(rst), .Q(sreg[351]) );
  DFF \sreg_reg[350]  ( .D(c[354]), .CLK(clk), .RST(rst), .Q(sreg[350]) );
  DFF \sreg_reg[349]  ( .D(c[353]), .CLK(clk), .RST(rst), .Q(sreg[349]) );
  DFF \sreg_reg[348]  ( .D(c[352]), .CLK(clk), .RST(rst), .Q(sreg[348]) );
  DFF \sreg_reg[347]  ( .D(c[351]), .CLK(clk), .RST(rst), .Q(sreg[347]) );
  DFF \sreg_reg[346]  ( .D(c[350]), .CLK(clk), .RST(rst), .Q(sreg[346]) );
  DFF \sreg_reg[345]  ( .D(c[349]), .CLK(clk), .RST(rst), .Q(sreg[345]) );
  DFF \sreg_reg[344]  ( .D(c[348]), .CLK(clk), .RST(rst), .Q(sreg[344]) );
  DFF \sreg_reg[343]  ( .D(c[347]), .CLK(clk), .RST(rst), .Q(sreg[343]) );
  DFF \sreg_reg[342]  ( .D(c[346]), .CLK(clk), .RST(rst), .Q(sreg[342]) );
  DFF \sreg_reg[341]  ( .D(c[345]), .CLK(clk), .RST(rst), .Q(sreg[341]) );
  DFF \sreg_reg[340]  ( .D(c[344]), .CLK(clk), .RST(rst), .Q(sreg[340]) );
  DFF \sreg_reg[339]  ( .D(c[343]), .CLK(clk), .RST(rst), .Q(sreg[339]) );
  DFF \sreg_reg[338]  ( .D(c[342]), .CLK(clk), .RST(rst), .Q(sreg[338]) );
  DFF \sreg_reg[337]  ( .D(c[341]), .CLK(clk), .RST(rst), .Q(sreg[337]) );
  DFF \sreg_reg[336]  ( .D(c[340]), .CLK(clk), .RST(rst), .Q(sreg[336]) );
  DFF \sreg_reg[335]  ( .D(c[339]), .CLK(clk), .RST(rst), .Q(sreg[335]) );
  DFF \sreg_reg[334]  ( .D(c[338]), .CLK(clk), .RST(rst), .Q(sreg[334]) );
  DFF \sreg_reg[333]  ( .D(c[337]), .CLK(clk), .RST(rst), .Q(sreg[333]) );
  DFF \sreg_reg[332]  ( .D(c[336]), .CLK(clk), .RST(rst), .Q(sreg[332]) );
  DFF \sreg_reg[331]  ( .D(c[335]), .CLK(clk), .RST(rst), .Q(sreg[331]) );
  DFF \sreg_reg[330]  ( .D(c[334]), .CLK(clk), .RST(rst), .Q(sreg[330]) );
  DFF \sreg_reg[329]  ( .D(c[333]), .CLK(clk), .RST(rst), .Q(sreg[329]) );
  DFF \sreg_reg[328]  ( .D(c[332]), .CLK(clk), .RST(rst), .Q(sreg[328]) );
  DFF \sreg_reg[327]  ( .D(c[331]), .CLK(clk), .RST(rst), .Q(sreg[327]) );
  DFF \sreg_reg[326]  ( .D(c[330]), .CLK(clk), .RST(rst), .Q(sreg[326]) );
  DFF \sreg_reg[325]  ( .D(c[329]), .CLK(clk), .RST(rst), .Q(sreg[325]) );
  DFF \sreg_reg[324]  ( .D(c[328]), .CLK(clk), .RST(rst), .Q(sreg[324]) );
  DFF \sreg_reg[323]  ( .D(c[327]), .CLK(clk), .RST(rst), .Q(sreg[323]) );
  DFF \sreg_reg[322]  ( .D(c[326]), .CLK(clk), .RST(rst), .Q(sreg[322]) );
  DFF \sreg_reg[321]  ( .D(c[325]), .CLK(clk), .RST(rst), .Q(sreg[321]) );
  DFF \sreg_reg[320]  ( .D(c[324]), .CLK(clk), .RST(rst), .Q(sreg[320]) );
  DFF \sreg_reg[319]  ( .D(c[323]), .CLK(clk), .RST(rst), .Q(sreg[319]) );
  DFF \sreg_reg[318]  ( .D(c[322]), .CLK(clk), .RST(rst), .Q(sreg[318]) );
  DFF \sreg_reg[317]  ( .D(c[321]), .CLK(clk), .RST(rst), .Q(sreg[317]) );
  DFF \sreg_reg[316]  ( .D(c[320]), .CLK(clk), .RST(rst), .Q(sreg[316]) );
  DFF \sreg_reg[315]  ( .D(c[319]), .CLK(clk), .RST(rst), .Q(sreg[315]) );
  DFF \sreg_reg[314]  ( .D(c[318]), .CLK(clk), .RST(rst), .Q(sreg[314]) );
  DFF \sreg_reg[313]  ( .D(c[317]), .CLK(clk), .RST(rst), .Q(sreg[313]) );
  DFF \sreg_reg[312]  ( .D(c[316]), .CLK(clk), .RST(rst), .Q(sreg[312]) );
  DFF \sreg_reg[311]  ( .D(c[315]), .CLK(clk), .RST(rst), .Q(sreg[311]) );
  DFF \sreg_reg[310]  ( .D(c[314]), .CLK(clk), .RST(rst), .Q(sreg[310]) );
  DFF \sreg_reg[309]  ( .D(c[313]), .CLK(clk), .RST(rst), .Q(sreg[309]) );
  DFF \sreg_reg[308]  ( .D(c[312]), .CLK(clk), .RST(rst), .Q(sreg[308]) );
  DFF \sreg_reg[307]  ( .D(c[311]), .CLK(clk), .RST(rst), .Q(sreg[307]) );
  DFF \sreg_reg[306]  ( .D(c[310]), .CLK(clk), .RST(rst), .Q(sreg[306]) );
  DFF \sreg_reg[305]  ( .D(c[309]), .CLK(clk), .RST(rst), .Q(sreg[305]) );
  DFF \sreg_reg[304]  ( .D(c[308]), .CLK(clk), .RST(rst), .Q(sreg[304]) );
  DFF \sreg_reg[303]  ( .D(c[307]), .CLK(clk), .RST(rst), .Q(sreg[303]) );
  DFF \sreg_reg[302]  ( .D(c[306]), .CLK(clk), .RST(rst), .Q(sreg[302]) );
  DFF \sreg_reg[301]  ( .D(c[305]), .CLK(clk), .RST(rst), .Q(sreg[301]) );
  DFF \sreg_reg[300]  ( .D(c[304]), .CLK(clk), .RST(rst), .Q(sreg[300]) );
  DFF \sreg_reg[299]  ( .D(c[303]), .CLK(clk), .RST(rst), .Q(sreg[299]) );
  DFF \sreg_reg[298]  ( .D(c[302]), .CLK(clk), .RST(rst), .Q(sreg[298]) );
  DFF \sreg_reg[297]  ( .D(c[301]), .CLK(clk), .RST(rst), .Q(sreg[297]) );
  DFF \sreg_reg[296]  ( .D(c[300]), .CLK(clk), .RST(rst), .Q(sreg[296]) );
  DFF \sreg_reg[295]  ( .D(c[299]), .CLK(clk), .RST(rst), .Q(sreg[295]) );
  DFF \sreg_reg[294]  ( .D(c[298]), .CLK(clk), .RST(rst), .Q(sreg[294]) );
  DFF \sreg_reg[293]  ( .D(c[297]), .CLK(clk), .RST(rst), .Q(sreg[293]) );
  DFF \sreg_reg[292]  ( .D(c[296]), .CLK(clk), .RST(rst), .Q(sreg[292]) );
  DFF \sreg_reg[291]  ( .D(c[295]), .CLK(clk), .RST(rst), .Q(sreg[291]) );
  DFF \sreg_reg[290]  ( .D(c[294]), .CLK(clk), .RST(rst), .Q(sreg[290]) );
  DFF \sreg_reg[289]  ( .D(c[293]), .CLK(clk), .RST(rst), .Q(sreg[289]) );
  DFF \sreg_reg[288]  ( .D(c[292]), .CLK(clk), .RST(rst), .Q(sreg[288]) );
  DFF \sreg_reg[287]  ( .D(c[291]), .CLK(clk), .RST(rst), .Q(sreg[287]) );
  DFF \sreg_reg[286]  ( .D(c[290]), .CLK(clk), .RST(rst), .Q(sreg[286]) );
  DFF \sreg_reg[285]  ( .D(c[289]), .CLK(clk), .RST(rst), .Q(sreg[285]) );
  DFF \sreg_reg[284]  ( .D(c[288]), .CLK(clk), .RST(rst), .Q(sreg[284]) );
  DFF \sreg_reg[283]  ( .D(c[287]), .CLK(clk), .RST(rst), .Q(sreg[283]) );
  DFF \sreg_reg[282]  ( .D(c[286]), .CLK(clk), .RST(rst), .Q(sreg[282]) );
  DFF \sreg_reg[281]  ( .D(c[285]), .CLK(clk), .RST(rst), .Q(sreg[281]) );
  DFF \sreg_reg[280]  ( .D(c[284]), .CLK(clk), .RST(rst), .Q(sreg[280]) );
  DFF \sreg_reg[279]  ( .D(c[283]), .CLK(clk), .RST(rst), .Q(sreg[279]) );
  DFF \sreg_reg[278]  ( .D(c[282]), .CLK(clk), .RST(rst), .Q(sreg[278]) );
  DFF \sreg_reg[277]  ( .D(c[281]), .CLK(clk), .RST(rst), .Q(sreg[277]) );
  DFF \sreg_reg[276]  ( .D(c[280]), .CLK(clk), .RST(rst), .Q(sreg[276]) );
  DFF \sreg_reg[275]  ( .D(c[279]), .CLK(clk), .RST(rst), .Q(sreg[275]) );
  DFF \sreg_reg[274]  ( .D(c[278]), .CLK(clk), .RST(rst), .Q(sreg[274]) );
  DFF \sreg_reg[273]  ( .D(c[277]), .CLK(clk), .RST(rst), .Q(sreg[273]) );
  DFF \sreg_reg[272]  ( .D(c[276]), .CLK(clk), .RST(rst), .Q(sreg[272]) );
  DFF \sreg_reg[271]  ( .D(c[275]), .CLK(clk), .RST(rst), .Q(sreg[271]) );
  DFF \sreg_reg[270]  ( .D(c[274]), .CLK(clk), .RST(rst), .Q(sreg[270]) );
  DFF \sreg_reg[269]  ( .D(c[273]), .CLK(clk), .RST(rst), .Q(sreg[269]) );
  DFF \sreg_reg[268]  ( .D(c[272]), .CLK(clk), .RST(rst), .Q(sreg[268]) );
  DFF \sreg_reg[267]  ( .D(c[271]), .CLK(clk), .RST(rst), .Q(sreg[267]) );
  DFF \sreg_reg[266]  ( .D(c[270]), .CLK(clk), .RST(rst), .Q(sreg[266]) );
  DFF \sreg_reg[265]  ( .D(c[269]), .CLK(clk), .RST(rst), .Q(sreg[265]) );
  DFF \sreg_reg[264]  ( .D(c[268]), .CLK(clk), .RST(rst), .Q(sreg[264]) );
  DFF \sreg_reg[263]  ( .D(c[267]), .CLK(clk), .RST(rst), .Q(sreg[263]) );
  DFF \sreg_reg[262]  ( .D(c[266]), .CLK(clk), .RST(rst), .Q(sreg[262]) );
  DFF \sreg_reg[261]  ( .D(c[265]), .CLK(clk), .RST(rst), .Q(sreg[261]) );
  DFF \sreg_reg[260]  ( .D(c[264]), .CLK(clk), .RST(rst), .Q(sreg[260]) );
  DFF \sreg_reg[259]  ( .D(c[263]), .CLK(clk), .RST(rst), .Q(sreg[259]) );
  DFF \sreg_reg[258]  ( .D(c[262]), .CLK(clk), .RST(rst), .Q(sreg[258]) );
  DFF \sreg_reg[257]  ( .D(c[261]), .CLK(clk), .RST(rst), .Q(sreg[257]) );
  DFF \sreg_reg[256]  ( .D(c[260]), .CLK(clk), .RST(rst), .Q(sreg[256]) );
  DFF \sreg_reg[255]  ( .D(c[259]), .CLK(clk), .RST(rst), .Q(sreg[255]) );
  DFF \sreg_reg[254]  ( .D(c[258]), .CLK(clk), .RST(rst), .Q(sreg[254]) );
  DFF \sreg_reg[253]  ( .D(c[257]), .CLK(clk), .RST(rst), .Q(sreg[253]) );
  DFF \sreg_reg[252]  ( .D(c[256]), .CLK(clk), .RST(rst), .Q(sreg[252]) );
  DFF \sreg_reg[251]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[251]) );
  DFF \sreg_reg[250]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[250]) );
  DFF \sreg_reg[249]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[249]) );
  DFF \sreg_reg[248]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[248]) );
  DFF \sreg_reg[247]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[247]) );
  DFF \sreg_reg[246]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[246]) );
  DFF \sreg_reg[245]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[245]) );
  DFF \sreg_reg[244]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[244]) );
  DFF \sreg_reg[243]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[243]) );
  DFF \sreg_reg[242]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[242]) );
  DFF \sreg_reg[241]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[241]) );
  DFF \sreg_reg[240]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[240]) );
  DFF \sreg_reg[239]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[239]) );
  DFF \sreg_reg[238]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[238]) );
  DFF \sreg_reg[237]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[237]) );
  DFF \sreg_reg[236]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[236]) );
  DFF \sreg_reg[235]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[235]) );
  DFF \sreg_reg[234]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[234]) );
  DFF \sreg_reg[233]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[233]) );
  DFF \sreg_reg[232]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[232]) );
  DFF \sreg_reg[231]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[231]) );
  DFF \sreg_reg[230]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[230]) );
  DFF \sreg_reg[229]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[229]) );
  DFF \sreg_reg[228]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[228]) );
  DFF \sreg_reg[227]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[227]) );
  DFF \sreg_reg[226]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[226]) );
  DFF \sreg_reg[225]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[225]) );
  DFF \sreg_reg[224]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[224]) );
  DFF \sreg_reg[223]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[222]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[221]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[220]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[219]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[218]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[217]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[216]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[215]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[214]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[213]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[212]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[211]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[210]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[209]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[208]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[207]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[206]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[205]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[204]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[203]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[202]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[201]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[200]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[199]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[198]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[197]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[196]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[195]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[194]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[193]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[192]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[191]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[190]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[189]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[188]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[187]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[186]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[185]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[184]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[183]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[182]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[181]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[180]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[179]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[178]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[177]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[176]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[175]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[174]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[173]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[172]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[171]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[170]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[169]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[168]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[167]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[166]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[165]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[164]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[163]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[162]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[161]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[160]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[159]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[158]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[157]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[156]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[155]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[154]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[153]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[152]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[151]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[150]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[149]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[148]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[147]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[146]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[145]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[144]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[143]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[142]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[141]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[140]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[139]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[138]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[137]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[136]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[135]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[134]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[133]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[132]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[131]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[130]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[129]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[128]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[127]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[126]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[125]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XOR U7 ( .A(n5887), .B(n5886), .Z(n5880) );
  NAND U8 ( .A(n5864), .B(n5863), .Z(n1) );
  NANDN U9 ( .A(n5862), .B(sreg[507]), .Z(n2) );
  NAND U10 ( .A(n1), .B(n2), .Z(n5865) );
  OR U11 ( .A(n5859), .B(n5858), .Z(n3) );
  NANDN U12 ( .A(n5861), .B(n5860), .Z(n4) );
  AND U13 ( .A(n3), .B(n4), .Z(n5867) );
  NANDN U14 ( .A(n5873), .B(n5874), .Z(n5) );
  NANDN U15 ( .A(n5875), .B(n5876), .Z(n6) );
  AND U16 ( .A(n5), .B(n6), .Z(n5881) );
  NAND U17 ( .A(n78), .B(n77), .Z(n7) );
  XOR U18 ( .A(n78), .B(n77), .Z(n8) );
  NANDN U19 ( .A(sreg[255]), .B(n8), .Z(n9) );
  NAND U20 ( .A(n7), .B(n9), .Z(n80) );
  XOR U21 ( .A(n5904), .B(n5905), .Z(n5899) );
  NANDN U22 ( .A(b[0]), .B(a[255]), .Z(n10) );
  NAND U23 ( .A(b[1]), .B(n10), .Z(n5875) );
  NANDN U24 ( .A(n5854), .B(n5853), .Z(n11) );
  NANDN U25 ( .A(n5851), .B(n5852), .Z(n12) );
  NAND U26 ( .A(n11), .B(n12), .Z(n5869) );
  NAND U27 ( .A(n80), .B(n81), .Z(n13) );
  XOR U28 ( .A(n80), .B(n81), .Z(n14) );
  NANDN U29 ( .A(sreg[256]), .B(n14), .Z(n15) );
  NAND U30 ( .A(n13), .B(n15), .Z(n120) );
  XNOR U31 ( .A(n5898), .B(n5899), .Z(n16) );
  NAND U32 ( .A(n5901), .B(n16), .Z(n17) );
  NANDN U33 ( .A(n5898), .B(n5899), .Z(n18) );
  AND U34 ( .A(n17), .B(n18), .Z(n19) );
  XOR U35 ( .A(n5901), .B(n16), .Z(n20) );
  NAND U36 ( .A(n20), .B(n5900), .Z(n21) );
  NAND U37 ( .A(n19), .B(n21), .Z(n22) );
  NAND U38 ( .A(n5904), .B(n5905), .Z(n23) );
  NAND U39 ( .A(n5903), .B(n5902), .Z(n24) );
  AND U40 ( .A(n23), .B(n24), .Z(n25) );
  XNOR U41 ( .A(a[255]), .B(a[253]), .Z(n26) );
  XNOR U42 ( .A(n5906), .B(n26), .Z(n27) );
  AND U43 ( .A(n27), .B(b[3]), .Z(n28) );
  XNOR U44 ( .A(n22), .B(n25), .Z(n29) );
  XNOR U45 ( .A(n28), .B(n29), .Z(c[511]) );
  NAND U46 ( .A(n49), .B(n5891), .Z(n30) );
  IV U47 ( .A(n30), .Z(n31) );
  AND U48 ( .A(b[0]), .B(a[0]), .Z(n33) );
  XOR U49 ( .A(n33), .B(sreg[252]), .Z(c[252]) );
  AND U50 ( .A(b[0]), .B(a[1]), .Z(n40) );
  NAND U51 ( .A(a[0]), .B(b[1]), .Z(n32) );
  XOR U52 ( .A(n40), .B(n32), .Z(n34) );
  XNOR U53 ( .A(sreg[253]), .B(n34), .Z(n36) );
  AND U54 ( .A(n33), .B(sreg[252]), .Z(n35) );
  XOR U55 ( .A(n36), .B(n35), .Z(c[253]) );
  NANDN U56 ( .A(n34), .B(sreg[253]), .Z(n38) );
  NAND U57 ( .A(n36), .B(n35), .Z(n37) );
  AND U58 ( .A(n38), .B(n37), .Z(n57) );
  XNOR U59 ( .A(n57), .B(sreg[254]), .Z(n59) );
  NAND U60 ( .A(a[0]), .B(b[2]), .Z(n39) );
  XNOR U61 ( .A(b[1]), .B(n39), .Z(n42) );
  NANDN U62 ( .A(a[0]), .B(n40), .Z(n41) );
  NAND U63 ( .A(n42), .B(n41), .Z(n56) );
  NAND U64 ( .A(b[0]), .B(a[2]), .Z(n43) );
  XNOR U65 ( .A(b[1]), .B(n43), .Z(n45) );
  NANDN U66 ( .A(b[0]), .B(a[1]), .Z(n44) );
  NAND U67 ( .A(n45), .B(n44), .Z(n55) );
  XOR U68 ( .A(n56), .B(n55), .Z(n58) );
  XOR U69 ( .A(n59), .B(n58), .Z(c[254]) );
  NAND U70 ( .A(b[0]), .B(a[3]), .Z(n46) );
  XNOR U71 ( .A(b[1]), .B(n46), .Z(n48) );
  NANDN U72 ( .A(b[0]), .B(a[2]), .Z(n47) );
  NAND U73 ( .A(n48), .B(n47), .Z(n76) );
  XOR U74 ( .A(b[3]), .B(a[1]), .Z(n69) );
  XNOR U75 ( .A(b[1]), .B(b[2]), .Z(n5891) );
  IV U76 ( .A(n5891), .Z(n5811) );
  AND U77 ( .A(n69), .B(n5811), .Z(n52) );
  XOR U78 ( .A(b[2]), .B(b[3]), .Z(n49) );
  XOR U79 ( .A(a[0]), .B(b[3]), .Z(n50) );
  NAND U80 ( .A(n31), .B(n50), .Z(n51) );
  NANDN U81 ( .A(n52), .B(n51), .Z(n75) );
  XNOR U82 ( .A(n76), .B(n75), .Z(n63) );
  NAND U83 ( .A(b[1]), .B(b[2]), .Z(n5906) );
  NAND U84 ( .A(n5811), .B(a[0]), .Z(n53) );
  AND U85 ( .A(n5906), .B(n53), .Z(n54) );
  NAND U86 ( .A(b[3]), .B(n54), .Z(n64) );
  XNOR U87 ( .A(n63), .B(n64), .Z(n66) );
  NOR U88 ( .A(n56), .B(n55), .Z(n65) );
  XNOR U89 ( .A(n66), .B(n65), .Z(n77) );
  NANDN U90 ( .A(n57), .B(sreg[254]), .Z(n61) );
  NAND U91 ( .A(n59), .B(n58), .Z(n60) );
  AND U92 ( .A(n61), .B(n60), .Z(n78) );
  XNOR U93 ( .A(sreg[255]), .B(n78), .Z(n62) );
  XNOR U94 ( .A(n77), .B(n62), .Z(c[255]) );
  NANDN U95 ( .A(n64), .B(n63), .Z(n68) );
  NAND U96 ( .A(n66), .B(n65), .Z(n67) );
  AND U97 ( .A(n68), .B(n67), .Z(n84) );
  NAND U98 ( .A(n31), .B(n69), .Z(n71) );
  XOR U99 ( .A(b[3]), .B(a[2]), .Z(n88) );
  NAND U100 ( .A(n5811), .B(n88), .Z(n70) );
  AND U101 ( .A(n71), .B(n70), .Z(n97) );
  AND U102 ( .A(b[3]), .B(a[0]), .Z(n94) );
  NAND U103 ( .A(b[0]), .B(a[4]), .Z(n72) );
  XNOR U104 ( .A(b[1]), .B(n72), .Z(n74) );
  NANDN U105 ( .A(b[0]), .B(a[3]), .Z(n73) );
  NAND U106 ( .A(n74), .B(n73), .Z(n95) );
  XNOR U107 ( .A(n94), .B(n95), .Z(n96) );
  XNOR U108 ( .A(n97), .B(n96), .Z(n82) );
  NANDN U109 ( .A(n76), .B(n75), .Z(n83) );
  XOR U110 ( .A(n82), .B(n83), .Z(n85) );
  XNOR U111 ( .A(n84), .B(n85), .Z(n81) );
  XNOR U112 ( .A(n80), .B(sreg[256]), .Z(n79) );
  XNOR U113 ( .A(n81), .B(n79), .Z(c[256]) );
  NANDN U114 ( .A(n83), .B(n82), .Z(n87) );
  OR U115 ( .A(n85), .B(n84), .Z(n86) );
  AND U116 ( .A(n87), .B(n86), .Z(n103) );
  NAND U117 ( .A(n31), .B(n88), .Z(n90) );
  XOR U118 ( .A(b[3]), .B(a[3]), .Z(n106) );
  NAND U119 ( .A(n5811), .B(n106), .Z(n89) );
  AND U120 ( .A(n90), .B(n89), .Z(n114) );
  AND U121 ( .A(b[0]), .B(a[5]), .Z(n91) );
  XOR U122 ( .A(b[1]), .B(n91), .Z(n93) );
  NANDN U123 ( .A(b[0]), .B(a[4]), .Z(n92) );
  AND U124 ( .A(n93), .B(n92), .Z(n112) );
  NAND U125 ( .A(b[3]), .B(a[1]), .Z(n113) );
  XOR U126 ( .A(n112), .B(n113), .Z(n115) );
  XOR U127 ( .A(n114), .B(n115), .Z(n101) );
  NANDN U128 ( .A(n95), .B(n94), .Z(n99) );
  NANDN U129 ( .A(n97), .B(n96), .Z(n98) );
  AND U130 ( .A(n99), .B(n98), .Z(n100) );
  XNOR U131 ( .A(n101), .B(n100), .Z(n102) );
  XOR U132 ( .A(n103), .B(n102), .Z(n118) );
  XNOR U133 ( .A(n118), .B(sreg[257]), .Z(n119) );
  XNOR U134 ( .A(n120), .B(n119), .Z(c[257]) );
  NANDN U135 ( .A(n101), .B(n100), .Z(n105) );
  NAND U136 ( .A(n103), .B(n102), .Z(n104) );
  AND U137 ( .A(n105), .B(n104), .Z(n125) );
  NAND U138 ( .A(n31), .B(n106), .Z(n108) );
  XOR U139 ( .A(b[3]), .B(a[4]), .Z(n129) );
  NAND U140 ( .A(n5811), .B(n129), .Z(n107) );
  AND U141 ( .A(n108), .B(n107), .Z(n137) );
  NAND U142 ( .A(b[0]), .B(a[6]), .Z(n109) );
  XNOR U143 ( .A(b[1]), .B(n109), .Z(n111) );
  NANDN U144 ( .A(b[0]), .B(a[5]), .Z(n110) );
  NAND U145 ( .A(n111), .B(n110), .Z(n136) );
  AND U146 ( .A(b[3]), .B(a[2]), .Z(n135) );
  XOR U147 ( .A(n136), .B(n135), .Z(n138) );
  XOR U148 ( .A(n137), .B(n138), .Z(n124) );
  NANDN U149 ( .A(n113), .B(n112), .Z(n117) );
  OR U150 ( .A(n115), .B(n114), .Z(n116) );
  AND U151 ( .A(n117), .B(n116), .Z(n123) );
  XOR U152 ( .A(n124), .B(n123), .Z(n126) );
  XOR U153 ( .A(n125), .B(n126), .Z(n141) );
  XNOR U154 ( .A(n141), .B(sreg[258]), .Z(n143) );
  NANDN U155 ( .A(n118), .B(sreg[257]), .Z(n122) );
  NANDN U156 ( .A(n120), .B(n119), .Z(n121) );
  NAND U157 ( .A(n122), .B(n121), .Z(n142) );
  XOR U158 ( .A(n143), .B(n142), .Z(c[258]) );
  NANDN U159 ( .A(n124), .B(n123), .Z(n128) );
  OR U160 ( .A(n126), .B(n125), .Z(n127) );
  AND U161 ( .A(n128), .B(n127), .Z(n148) );
  NAND U162 ( .A(n31), .B(n129), .Z(n131) );
  XOR U163 ( .A(b[3]), .B(a[5]), .Z(n152) );
  NAND U164 ( .A(n5811), .B(n152), .Z(n130) );
  AND U165 ( .A(n131), .B(n130), .Z(n160) );
  AND U166 ( .A(b[3]), .B(a[3]), .Z(n158) );
  NAND U167 ( .A(b[0]), .B(a[7]), .Z(n132) );
  XNOR U168 ( .A(b[1]), .B(n132), .Z(n134) );
  NANDN U169 ( .A(b[0]), .B(a[6]), .Z(n133) );
  NAND U170 ( .A(n134), .B(n133), .Z(n159) );
  XOR U171 ( .A(n158), .B(n159), .Z(n161) );
  XOR U172 ( .A(n160), .B(n161), .Z(n147) );
  NANDN U173 ( .A(n136), .B(n135), .Z(n140) );
  OR U174 ( .A(n138), .B(n137), .Z(n139) );
  AND U175 ( .A(n140), .B(n139), .Z(n146) );
  XOR U176 ( .A(n147), .B(n146), .Z(n149) );
  XOR U177 ( .A(n148), .B(n149), .Z(n164) );
  XNOR U178 ( .A(n164), .B(sreg[259]), .Z(n166) );
  NANDN U179 ( .A(n141), .B(sreg[258]), .Z(n145) );
  NAND U180 ( .A(n143), .B(n142), .Z(n144) );
  NAND U181 ( .A(n145), .B(n144), .Z(n165) );
  XOR U182 ( .A(n166), .B(n165), .Z(c[259]) );
  NANDN U183 ( .A(n147), .B(n146), .Z(n151) );
  OR U184 ( .A(n149), .B(n148), .Z(n150) );
  AND U185 ( .A(n151), .B(n150), .Z(n171) );
  NAND U186 ( .A(n31), .B(n152), .Z(n154) );
  XOR U187 ( .A(b[3]), .B(a[6]), .Z(n175) );
  NAND U188 ( .A(n5811), .B(n175), .Z(n153) );
  AND U189 ( .A(n154), .B(n153), .Z(n183) );
  NAND U190 ( .A(b[0]), .B(a[8]), .Z(n155) );
  XNOR U191 ( .A(b[1]), .B(n155), .Z(n157) );
  NANDN U192 ( .A(b[0]), .B(a[7]), .Z(n156) );
  NAND U193 ( .A(n157), .B(n156), .Z(n182) );
  AND U194 ( .A(b[3]), .B(a[4]), .Z(n181) );
  XOR U195 ( .A(n182), .B(n181), .Z(n184) );
  XOR U196 ( .A(n183), .B(n184), .Z(n170) );
  NANDN U197 ( .A(n159), .B(n158), .Z(n163) );
  OR U198 ( .A(n161), .B(n160), .Z(n162) );
  AND U199 ( .A(n163), .B(n162), .Z(n169) );
  XOR U200 ( .A(n170), .B(n169), .Z(n172) );
  XOR U201 ( .A(n171), .B(n172), .Z(n187) );
  XNOR U202 ( .A(n187), .B(sreg[260]), .Z(n189) );
  NANDN U203 ( .A(n164), .B(sreg[259]), .Z(n168) );
  NAND U204 ( .A(n166), .B(n165), .Z(n167) );
  NAND U205 ( .A(n168), .B(n167), .Z(n188) );
  XOR U206 ( .A(n189), .B(n188), .Z(c[260]) );
  NANDN U207 ( .A(n170), .B(n169), .Z(n174) );
  OR U208 ( .A(n172), .B(n171), .Z(n173) );
  AND U209 ( .A(n174), .B(n173), .Z(n194) );
  NAND U210 ( .A(n31), .B(n175), .Z(n177) );
  XOR U211 ( .A(b[3]), .B(a[7]), .Z(n198) );
  NAND U212 ( .A(n5811), .B(n198), .Z(n176) );
  AND U213 ( .A(n177), .B(n176), .Z(n206) );
  NAND U214 ( .A(b[0]), .B(a[9]), .Z(n178) );
  XNOR U215 ( .A(b[1]), .B(n178), .Z(n180) );
  NANDN U216 ( .A(b[0]), .B(a[8]), .Z(n179) );
  NAND U217 ( .A(n180), .B(n179), .Z(n205) );
  AND U218 ( .A(b[3]), .B(a[5]), .Z(n204) );
  XOR U219 ( .A(n205), .B(n204), .Z(n207) );
  XOR U220 ( .A(n206), .B(n207), .Z(n193) );
  NANDN U221 ( .A(n182), .B(n181), .Z(n186) );
  OR U222 ( .A(n184), .B(n183), .Z(n185) );
  AND U223 ( .A(n186), .B(n185), .Z(n192) );
  XOR U224 ( .A(n193), .B(n192), .Z(n195) );
  XOR U225 ( .A(n194), .B(n195), .Z(n210) );
  XNOR U226 ( .A(n210), .B(sreg[261]), .Z(n212) );
  NANDN U227 ( .A(n187), .B(sreg[260]), .Z(n191) );
  NAND U228 ( .A(n189), .B(n188), .Z(n190) );
  NAND U229 ( .A(n191), .B(n190), .Z(n211) );
  XOR U230 ( .A(n212), .B(n211), .Z(c[261]) );
  NANDN U231 ( .A(n193), .B(n192), .Z(n197) );
  OR U232 ( .A(n195), .B(n194), .Z(n196) );
  AND U233 ( .A(n197), .B(n196), .Z(n217) );
  NAND U234 ( .A(n31), .B(n198), .Z(n200) );
  XOR U235 ( .A(b[3]), .B(a[8]), .Z(n221) );
  NAND U236 ( .A(n5811), .B(n221), .Z(n199) );
  AND U237 ( .A(n200), .B(n199), .Z(n229) );
  AND U238 ( .A(b[3]), .B(a[6]), .Z(n227) );
  NAND U239 ( .A(b[0]), .B(a[10]), .Z(n201) );
  XNOR U240 ( .A(b[1]), .B(n201), .Z(n203) );
  NANDN U241 ( .A(b[0]), .B(a[9]), .Z(n202) );
  NAND U242 ( .A(n203), .B(n202), .Z(n228) );
  XOR U243 ( .A(n227), .B(n228), .Z(n230) );
  XOR U244 ( .A(n229), .B(n230), .Z(n216) );
  NANDN U245 ( .A(n205), .B(n204), .Z(n209) );
  OR U246 ( .A(n207), .B(n206), .Z(n208) );
  AND U247 ( .A(n209), .B(n208), .Z(n215) );
  XOR U248 ( .A(n216), .B(n215), .Z(n218) );
  XOR U249 ( .A(n217), .B(n218), .Z(n233) );
  XNOR U250 ( .A(n233), .B(sreg[262]), .Z(n235) );
  NANDN U251 ( .A(n210), .B(sreg[261]), .Z(n214) );
  NAND U252 ( .A(n212), .B(n211), .Z(n213) );
  NAND U253 ( .A(n214), .B(n213), .Z(n234) );
  XOR U254 ( .A(n235), .B(n234), .Z(c[262]) );
  NANDN U255 ( .A(n216), .B(n215), .Z(n220) );
  OR U256 ( .A(n218), .B(n217), .Z(n219) );
  AND U257 ( .A(n220), .B(n219), .Z(n240) );
  NAND U258 ( .A(n31), .B(n221), .Z(n223) );
  XOR U259 ( .A(b[3]), .B(a[9]), .Z(n244) );
  NAND U260 ( .A(n5811), .B(n244), .Z(n222) );
  AND U261 ( .A(n223), .B(n222), .Z(n252) );
  NAND U262 ( .A(b[0]), .B(a[11]), .Z(n224) );
  XNOR U263 ( .A(b[1]), .B(n224), .Z(n226) );
  NANDN U264 ( .A(b[0]), .B(a[10]), .Z(n225) );
  NAND U265 ( .A(n226), .B(n225), .Z(n251) );
  AND U266 ( .A(b[3]), .B(a[7]), .Z(n250) );
  XOR U267 ( .A(n251), .B(n250), .Z(n253) );
  XOR U268 ( .A(n252), .B(n253), .Z(n239) );
  NANDN U269 ( .A(n228), .B(n227), .Z(n232) );
  OR U270 ( .A(n230), .B(n229), .Z(n231) );
  AND U271 ( .A(n232), .B(n231), .Z(n238) );
  XOR U272 ( .A(n239), .B(n238), .Z(n241) );
  XOR U273 ( .A(n240), .B(n241), .Z(n256) );
  XNOR U274 ( .A(n256), .B(sreg[263]), .Z(n258) );
  NANDN U275 ( .A(n233), .B(sreg[262]), .Z(n237) );
  NAND U276 ( .A(n235), .B(n234), .Z(n236) );
  NAND U277 ( .A(n237), .B(n236), .Z(n257) );
  XOR U278 ( .A(n258), .B(n257), .Z(c[263]) );
  NANDN U279 ( .A(n239), .B(n238), .Z(n243) );
  OR U280 ( .A(n241), .B(n240), .Z(n242) );
  AND U281 ( .A(n243), .B(n242), .Z(n263) );
  NAND U282 ( .A(n31), .B(n244), .Z(n246) );
  XOR U283 ( .A(b[3]), .B(a[10]), .Z(n267) );
  NAND U284 ( .A(n5811), .B(n267), .Z(n245) );
  AND U285 ( .A(n246), .B(n245), .Z(n275) );
  NAND U286 ( .A(b[0]), .B(a[12]), .Z(n247) );
  XNOR U287 ( .A(b[1]), .B(n247), .Z(n249) );
  NANDN U288 ( .A(b[0]), .B(a[11]), .Z(n248) );
  NAND U289 ( .A(n249), .B(n248), .Z(n274) );
  AND U290 ( .A(b[3]), .B(a[8]), .Z(n273) );
  XOR U291 ( .A(n274), .B(n273), .Z(n276) );
  XOR U292 ( .A(n275), .B(n276), .Z(n262) );
  NANDN U293 ( .A(n251), .B(n250), .Z(n255) );
  OR U294 ( .A(n253), .B(n252), .Z(n254) );
  AND U295 ( .A(n255), .B(n254), .Z(n261) );
  XOR U296 ( .A(n262), .B(n261), .Z(n264) );
  XOR U297 ( .A(n263), .B(n264), .Z(n279) );
  XNOR U298 ( .A(n279), .B(sreg[264]), .Z(n281) );
  NANDN U299 ( .A(n256), .B(sreg[263]), .Z(n260) );
  NAND U300 ( .A(n258), .B(n257), .Z(n259) );
  NAND U301 ( .A(n260), .B(n259), .Z(n280) );
  XOR U302 ( .A(n281), .B(n280), .Z(c[264]) );
  NANDN U303 ( .A(n262), .B(n261), .Z(n266) );
  OR U304 ( .A(n264), .B(n263), .Z(n265) );
  AND U305 ( .A(n266), .B(n265), .Z(n286) );
  NAND U306 ( .A(n31), .B(n267), .Z(n269) );
  XOR U307 ( .A(b[3]), .B(a[11]), .Z(n290) );
  NAND U308 ( .A(n5811), .B(n290), .Z(n268) );
  AND U309 ( .A(n269), .B(n268), .Z(n298) );
  NAND U310 ( .A(b[0]), .B(a[13]), .Z(n270) );
  XNOR U311 ( .A(b[1]), .B(n270), .Z(n272) );
  NANDN U312 ( .A(b[0]), .B(a[12]), .Z(n271) );
  NAND U313 ( .A(n272), .B(n271), .Z(n297) );
  AND U314 ( .A(b[3]), .B(a[9]), .Z(n296) );
  XOR U315 ( .A(n297), .B(n296), .Z(n299) );
  XOR U316 ( .A(n298), .B(n299), .Z(n285) );
  NANDN U317 ( .A(n274), .B(n273), .Z(n278) );
  OR U318 ( .A(n276), .B(n275), .Z(n277) );
  AND U319 ( .A(n278), .B(n277), .Z(n284) );
  XOR U320 ( .A(n285), .B(n284), .Z(n287) );
  XOR U321 ( .A(n286), .B(n287), .Z(n302) );
  XNOR U322 ( .A(n302), .B(sreg[265]), .Z(n304) );
  NANDN U323 ( .A(n279), .B(sreg[264]), .Z(n283) );
  NAND U324 ( .A(n281), .B(n280), .Z(n282) );
  NAND U325 ( .A(n283), .B(n282), .Z(n303) );
  XOR U326 ( .A(n304), .B(n303), .Z(c[265]) );
  NANDN U327 ( .A(n285), .B(n284), .Z(n289) );
  OR U328 ( .A(n287), .B(n286), .Z(n288) );
  AND U329 ( .A(n289), .B(n288), .Z(n309) );
  NAND U330 ( .A(n31), .B(n290), .Z(n292) );
  XOR U331 ( .A(b[3]), .B(a[12]), .Z(n313) );
  NAND U332 ( .A(n5811), .B(n313), .Z(n291) );
  AND U333 ( .A(n292), .B(n291), .Z(n321) );
  NAND U334 ( .A(b[0]), .B(a[14]), .Z(n293) );
  XNOR U335 ( .A(b[1]), .B(n293), .Z(n295) );
  NANDN U336 ( .A(b[0]), .B(a[13]), .Z(n294) );
  NAND U337 ( .A(n295), .B(n294), .Z(n320) );
  AND U338 ( .A(b[3]), .B(a[10]), .Z(n319) );
  XOR U339 ( .A(n320), .B(n319), .Z(n322) );
  XOR U340 ( .A(n321), .B(n322), .Z(n308) );
  NANDN U341 ( .A(n297), .B(n296), .Z(n301) );
  OR U342 ( .A(n299), .B(n298), .Z(n300) );
  AND U343 ( .A(n301), .B(n300), .Z(n307) );
  XOR U344 ( .A(n308), .B(n307), .Z(n310) );
  XOR U345 ( .A(n309), .B(n310), .Z(n325) );
  XNOR U346 ( .A(n325), .B(sreg[266]), .Z(n327) );
  NANDN U347 ( .A(n302), .B(sreg[265]), .Z(n306) );
  NAND U348 ( .A(n304), .B(n303), .Z(n305) );
  NAND U349 ( .A(n306), .B(n305), .Z(n326) );
  XOR U350 ( .A(n327), .B(n326), .Z(c[266]) );
  NANDN U351 ( .A(n308), .B(n307), .Z(n312) );
  OR U352 ( .A(n310), .B(n309), .Z(n311) );
  AND U353 ( .A(n312), .B(n311), .Z(n332) );
  NAND U354 ( .A(n31), .B(n313), .Z(n315) );
  XOR U355 ( .A(b[3]), .B(a[13]), .Z(n336) );
  NAND U356 ( .A(n5811), .B(n336), .Z(n314) );
  AND U357 ( .A(n315), .B(n314), .Z(n344) );
  NAND U358 ( .A(b[0]), .B(a[15]), .Z(n316) );
  XNOR U359 ( .A(b[1]), .B(n316), .Z(n318) );
  NANDN U360 ( .A(b[0]), .B(a[14]), .Z(n317) );
  NAND U361 ( .A(n318), .B(n317), .Z(n343) );
  AND U362 ( .A(b[3]), .B(a[11]), .Z(n342) );
  XOR U363 ( .A(n343), .B(n342), .Z(n345) );
  XOR U364 ( .A(n344), .B(n345), .Z(n331) );
  NANDN U365 ( .A(n320), .B(n319), .Z(n324) );
  OR U366 ( .A(n322), .B(n321), .Z(n323) );
  AND U367 ( .A(n324), .B(n323), .Z(n330) );
  XOR U368 ( .A(n331), .B(n330), .Z(n333) );
  XOR U369 ( .A(n332), .B(n333), .Z(n348) );
  XNOR U370 ( .A(n348), .B(sreg[267]), .Z(n350) );
  NANDN U371 ( .A(n325), .B(sreg[266]), .Z(n329) );
  NAND U372 ( .A(n327), .B(n326), .Z(n328) );
  NAND U373 ( .A(n329), .B(n328), .Z(n349) );
  XOR U374 ( .A(n350), .B(n349), .Z(c[267]) );
  NANDN U375 ( .A(n331), .B(n330), .Z(n335) );
  OR U376 ( .A(n333), .B(n332), .Z(n334) );
  AND U377 ( .A(n335), .B(n334), .Z(n355) );
  NAND U378 ( .A(n31), .B(n336), .Z(n338) );
  XOR U379 ( .A(b[3]), .B(a[14]), .Z(n359) );
  NAND U380 ( .A(n5811), .B(n359), .Z(n337) );
  AND U381 ( .A(n338), .B(n337), .Z(n367) );
  AND U382 ( .A(b[3]), .B(a[12]), .Z(n365) );
  NAND U383 ( .A(b[0]), .B(a[16]), .Z(n339) );
  XNOR U384 ( .A(b[1]), .B(n339), .Z(n341) );
  NANDN U385 ( .A(b[0]), .B(a[15]), .Z(n340) );
  NAND U386 ( .A(n341), .B(n340), .Z(n366) );
  XOR U387 ( .A(n365), .B(n366), .Z(n368) );
  XOR U388 ( .A(n367), .B(n368), .Z(n354) );
  NANDN U389 ( .A(n343), .B(n342), .Z(n347) );
  OR U390 ( .A(n345), .B(n344), .Z(n346) );
  AND U391 ( .A(n347), .B(n346), .Z(n353) );
  XOR U392 ( .A(n354), .B(n353), .Z(n356) );
  XOR U393 ( .A(n355), .B(n356), .Z(n371) );
  XNOR U394 ( .A(n371), .B(sreg[268]), .Z(n373) );
  NANDN U395 ( .A(n348), .B(sreg[267]), .Z(n352) );
  NAND U396 ( .A(n350), .B(n349), .Z(n351) );
  NAND U397 ( .A(n352), .B(n351), .Z(n372) );
  XOR U398 ( .A(n373), .B(n372), .Z(c[268]) );
  NANDN U399 ( .A(n354), .B(n353), .Z(n358) );
  OR U400 ( .A(n356), .B(n355), .Z(n357) );
  AND U401 ( .A(n358), .B(n357), .Z(n378) );
  NAND U402 ( .A(n31), .B(n359), .Z(n361) );
  XOR U403 ( .A(b[3]), .B(a[15]), .Z(n382) );
  NAND U404 ( .A(n5811), .B(n382), .Z(n360) );
  AND U405 ( .A(n361), .B(n360), .Z(n390) );
  NAND U406 ( .A(b[0]), .B(a[17]), .Z(n362) );
  XNOR U407 ( .A(b[1]), .B(n362), .Z(n364) );
  NANDN U408 ( .A(b[0]), .B(a[16]), .Z(n363) );
  NAND U409 ( .A(n364), .B(n363), .Z(n389) );
  AND U410 ( .A(b[3]), .B(a[13]), .Z(n388) );
  XOR U411 ( .A(n389), .B(n388), .Z(n391) );
  XOR U412 ( .A(n390), .B(n391), .Z(n377) );
  NANDN U413 ( .A(n366), .B(n365), .Z(n370) );
  OR U414 ( .A(n368), .B(n367), .Z(n369) );
  AND U415 ( .A(n370), .B(n369), .Z(n376) );
  XOR U416 ( .A(n377), .B(n376), .Z(n379) );
  XOR U417 ( .A(n378), .B(n379), .Z(n394) );
  XNOR U418 ( .A(n394), .B(sreg[269]), .Z(n396) );
  NANDN U419 ( .A(n371), .B(sreg[268]), .Z(n375) );
  NAND U420 ( .A(n373), .B(n372), .Z(n374) );
  NAND U421 ( .A(n375), .B(n374), .Z(n395) );
  XOR U422 ( .A(n396), .B(n395), .Z(c[269]) );
  NANDN U423 ( .A(n377), .B(n376), .Z(n381) );
  OR U424 ( .A(n379), .B(n378), .Z(n380) );
  AND U425 ( .A(n381), .B(n380), .Z(n401) );
  NAND U426 ( .A(n31), .B(n382), .Z(n384) );
  XOR U427 ( .A(b[3]), .B(a[16]), .Z(n405) );
  NAND U428 ( .A(n5811), .B(n405), .Z(n383) );
  AND U429 ( .A(n384), .B(n383), .Z(n413) );
  NAND U430 ( .A(b[0]), .B(a[18]), .Z(n385) );
  XNOR U431 ( .A(b[1]), .B(n385), .Z(n387) );
  NANDN U432 ( .A(b[0]), .B(a[17]), .Z(n386) );
  NAND U433 ( .A(n387), .B(n386), .Z(n412) );
  AND U434 ( .A(b[3]), .B(a[14]), .Z(n411) );
  XOR U435 ( .A(n412), .B(n411), .Z(n414) );
  XOR U436 ( .A(n413), .B(n414), .Z(n400) );
  NANDN U437 ( .A(n389), .B(n388), .Z(n393) );
  OR U438 ( .A(n391), .B(n390), .Z(n392) );
  AND U439 ( .A(n393), .B(n392), .Z(n399) );
  XOR U440 ( .A(n400), .B(n399), .Z(n402) );
  XOR U441 ( .A(n401), .B(n402), .Z(n417) );
  XNOR U442 ( .A(n417), .B(sreg[270]), .Z(n419) );
  NANDN U443 ( .A(n394), .B(sreg[269]), .Z(n398) );
  NAND U444 ( .A(n396), .B(n395), .Z(n397) );
  NAND U445 ( .A(n398), .B(n397), .Z(n418) );
  XOR U446 ( .A(n419), .B(n418), .Z(c[270]) );
  NANDN U447 ( .A(n400), .B(n399), .Z(n404) );
  OR U448 ( .A(n402), .B(n401), .Z(n403) );
  AND U449 ( .A(n404), .B(n403), .Z(n424) );
  NAND U450 ( .A(n31), .B(n405), .Z(n407) );
  XOR U451 ( .A(b[3]), .B(a[17]), .Z(n428) );
  NAND U452 ( .A(n5811), .B(n428), .Z(n406) );
  AND U453 ( .A(n407), .B(n406), .Z(n436) );
  NAND U454 ( .A(b[0]), .B(a[19]), .Z(n408) );
  XNOR U455 ( .A(b[1]), .B(n408), .Z(n410) );
  NANDN U456 ( .A(b[0]), .B(a[18]), .Z(n409) );
  NAND U457 ( .A(n410), .B(n409), .Z(n435) );
  AND U458 ( .A(b[3]), .B(a[15]), .Z(n434) );
  XOR U459 ( .A(n435), .B(n434), .Z(n437) );
  XOR U460 ( .A(n436), .B(n437), .Z(n423) );
  NANDN U461 ( .A(n412), .B(n411), .Z(n416) );
  OR U462 ( .A(n414), .B(n413), .Z(n415) );
  AND U463 ( .A(n416), .B(n415), .Z(n422) );
  XOR U464 ( .A(n423), .B(n422), .Z(n425) );
  XOR U465 ( .A(n424), .B(n425), .Z(n440) );
  XNOR U466 ( .A(n440), .B(sreg[271]), .Z(n442) );
  NANDN U467 ( .A(n417), .B(sreg[270]), .Z(n421) );
  NAND U468 ( .A(n419), .B(n418), .Z(n420) );
  NAND U469 ( .A(n421), .B(n420), .Z(n441) );
  XOR U470 ( .A(n442), .B(n441), .Z(c[271]) );
  NANDN U471 ( .A(n423), .B(n422), .Z(n427) );
  OR U472 ( .A(n425), .B(n424), .Z(n426) );
  AND U473 ( .A(n427), .B(n426), .Z(n447) );
  NAND U474 ( .A(n31), .B(n428), .Z(n430) );
  XOR U475 ( .A(b[3]), .B(a[18]), .Z(n451) );
  NAND U476 ( .A(n5811), .B(n451), .Z(n429) );
  AND U477 ( .A(n430), .B(n429), .Z(n459) );
  AND U478 ( .A(b[3]), .B(a[16]), .Z(n457) );
  NAND U479 ( .A(b[0]), .B(a[20]), .Z(n431) );
  XNOR U480 ( .A(b[1]), .B(n431), .Z(n433) );
  NANDN U481 ( .A(b[0]), .B(a[19]), .Z(n432) );
  NAND U482 ( .A(n433), .B(n432), .Z(n458) );
  XOR U483 ( .A(n457), .B(n458), .Z(n460) );
  XOR U484 ( .A(n459), .B(n460), .Z(n446) );
  NANDN U485 ( .A(n435), .B(n434), .Z(n439) );
  OR U486 ( .A(n437), .B(n436), .Z(n438) );
  AND U487 ( .A(n439), .B(n438), .Z(n445) );
  XOR U488 ( .A(n446), .B(n445), .Z(n448) );
  XOR U489 ( .A(n447), .B(n448), .Z(n463) );
  XNOR U490 ( .A(n463), .B(sreg[272]), .Z(n465) );
  NANDN U491 ( .A(n440), .B(sreg[271]), .Z(n444) );
  NAND U492 ( .A(n442), .B(n441), .Z(n443) );
  NAND U493 ( .A(n444), .B(n443), .Z(n464) );
  XOR U494 ( .A(n465), .B(n464), .Z(c[272]) );
  NANDN U495 ( .A(n446), .B(n445), .Z(n450) );
  OR U496 ( .A(n448), .B(n447), .Z(n449) );
  AND U497 ( .A(n450), .B(n449), .Z(n470) );
  NAND U498 ( .A(n31), .B(n451), .Z(n453) );
  XOR U499 ( .A(b[3]), .B(a[19]), .Z(n474) );
  NAND U500 ( .A(n5811), .B(n474), .Z(n452) );
  AND U501 ( .A(n453), .B(n452), .Z(n482) );
  NAND U502 ( .A(b[0]), .B(a[21]), .Z(n454) );
  XNOR U503 ( .A(b[1]), .B(n454), .Z(n456) );
  NANDN U504 ( .A(b[0]), .B(a[20]), .Z(n455) );
  NAND U505 ( .A(n456), .B(n455), .Z(n481) );
  AND U506 ( .A(b[3]), .B(a[17]), .Z(n480) );
  XOR U507 ( .A(n481), .B(n480), .Z(n483) );
  XOR U508 ( .A(n482), .B(n483), .Z(n469) );
  NANDN U509 ( .A(n458), .B(n457), .Z(n462) );
  OR U510 ( .A(n460), .B(n459), .Z(n461) );
  AND U511 ( .A(n462), .B(n461), .Z(n468) );
  XOR U512 ( .A(n469), .B(n468), .Z(n471) );
  XOR U513 ( .A(n470), .B(n471), .Z(n486) );
  XNOR U514 ( .A(n486), .B(sreg[273]), .Z(n488) );
  NANDN U515 ( .A(n463), .B(sreg[272]), .Z(n467) );
  NAND U516 ( .A(n465), .B(n464), .Z(n466) );
  NAND U517 ( .A(n467), .B(n466), .Z(n487) );
  XOR U518 ( .A(n488), .B(n487), .Z(c[273]) );
  NANDN U519 ( .A(n469), .B(n468), .Z(n473) );
  OR U520 ( .A(n471), .B(n470), .Z(n472) );
  AND U521 ( .A(n473), .B(n472), .Z(n493) );
  NAND U522 ( .A(n31), .B(n474), .Z(n476) );
  XOR U523 ( .A(b[3]), .B(a[20]), .Z(n497) );
  NAND U524 ( .A(n5811), .B(n497), .Z(n475) );
  AND U525 ( .A(n476), .B(n475), .Z(n505) );
  NAND U526 ( .A(b[0]), .B(a[22]), .Z(n477) );
  XNOR U527 ( .A(b[1]), .B(n477), .Z(n479) );
  NANDN U528 ( .A(b[0]), .B(a[21]), .Z(n478) );
  NAND U529 ( .A(n479), .B(n478), .Z(n504) );
  AND U530 ( .A(b[3]), .B(a[18]), .Z(n503) );
  XOR U531 ( .A(n504), .B(n503), .Z(n506) );
  XOR U532 ( .A(n505), .B(n506), .Z(n492) );
  NANDN U533 ( .A(n481), .B(n480), .Z(n485) );
  OR U534 ( .A(n483), .B(n482), .Z(n484) );
  AND U535 ( .A(n485), .B(n484), .Z(n491) );
  XOR U536 ( .A(n492), .B(n491), .Z(n494) );
  XOR U537 ( .A(n493), .B(n494), .Z(n509) );
  XNOR U538 ( .A(n509), .B(sreg[274]), .Z(n511) );
  NANDN U539 ( .A(n486), .B(sreg[273]), .Z(n490) );
  NAND U540 ( .A(n488), .B(n487), .Z(n489) );
  NAND U541 ( .A(n490), .B(n489), .Z(n510) );
  XOR U542 ( .A(n511), .B(n510), .Z(c[274]) );
  NANDN U543 ( .A(n492), .B(n491), .Z(n496) );
  OR U544 ( .A(n494), .B(n493), .Z(n495) );
  AND U545 ( .A(n496), .B(n495), .Z(n516) );
  NAND U546 ( .A(n31), .B(n497), .Z(n499) );
  XOR U547 ( .A(b[3]), .B(a[21]), .Z(n520) );
  NAND U548 ( .A(n5811), .B(n520), .Z(n498) );
  AND U549 ( .A(n499), .B(n498), .Z(n528) );
  NAND U550 ( .A(b[0]), .B(a[23]), .Z(n500) );
  XNOR U551 ( .A(b[1]), .B(n500), .Z(n502) );
  NANDN U552 ( .A(b[0]), .B(a[22]), .Z(n501) );
  NAND U553 ( .A(n502), .B(n501), .Z(n527) );
  AND U554 ( .A(b[3]), .B(a[19]), .Z(n526) );
  XOR U555 ( .A(n527), .B(n526), .Z(n529) );
  XOR U556 ( .A(n528), .B(n529), .Z(n515) );
  NANDN U557 ( .A(n504), .B(n503), .Z(n508) );
  OR U558 ( .A(n506), .B(n505), .Z(n507) );
  AND U559 ( .A(n508), .B(n507), .Z(n514) );
  XOR U560 ( .A(n515), .B(n514), .Z(n517) );
  XOR U561 ( .A(n516), .B(n517), .Z(n532) );
  XNOR U562 ( .A(n532), .B(sreg[275]), .Z(n534) );
  NANDN U563 ( .A(n509), .B(sreg[274]), .Z(n513) );
  NAND U564 ( .A(n511), .B(n510), .Z(n512) );
  NAND U565 ( .A(n513), .B(n512), .Z(n533) );
  XOR U566 ( .A(n534), .B(n533), .Z(c[275]) );
  NANDN U567 ( .A(n515), .B(n514), .Z(n519) );
  OR U568 ( .A(n517), .B(n516), .Z(n518) );
  AND U569 ( .A(n519), .B(n518), .Z(n539) );
  NAND U570 ( .A(n31), .B(n520), .Z(n522) );
  XOR U571 ( .A(b[3]), .B(a[22]), .Z(n543) );
  NAND U572 ( .A(n5811), .B(n543), .Z(n521) );
  AND U573 ( .A(n522), .B(n521), .Z(n551) );
  NAND U574 ( .A(b[0]), .B(a[24]), .Z(n523) );
  XNOR U575 ( .A(b[1]), .B(n523), .Z(n525) );
  NANDN U576 ( .A(b[0]), .B(a[23]), .Z(n524) );
  NAND U577 ( .A(n525), .B(n524), .Z(n550) );
  AND U578 ( .A(b[3]), .B(a[20]), .Z(n549) );
  XOR U579 ( .A(n550), .B(n549), .Z(n552) );
  XOR U580 ( .A(n551), .B(n552), .Z(n538) );
  NANDN U581 ( .A(n527), .B(n526), .Z(n531) );
  OR U582 ( .A(n529), .B(n528), .Z(n530) );
  AND U583 ( .A(n531), .B(n530), .Z(n537) );
  XOR U584 ( .A(n538), .B(n537), .Z(n540) );
  XOR U585 ( .A(n539), .B(n540), .Z(n555) );
  XNOR U586 ( .A(n555), .B(sreg[276]), .Z(n557) );
  NANDN U587 ( .A(n532), .B(sreg[275]), .Z(n536) );
  NAND U588 ( .A(n534), .B(n533), .Z(n535) );
  NAND U589 ( .A(n536), .B(n535), .Z(n556) );
  XOR U590 ( .A(n557), .B(n556), .Z(c[276]) );
  NANDN U591 ( .A(n538), .B(n537), .Z(n542) );
  OR U592 ( .A(n540), .B(n539), .Z(n541) );
  AND U593 ( .A(n542), .B(n541), .Z(n562) );
  NAND U594 ( .A(n31), .B(n543), .Z(n545) );
  XOR U595 ( .A(b[3]), .B(a[23]), .Z(n566) );
  NAND U596 ( .A(n5811), .B(n566), .Z(n544) );
  AND U597 ( .A(n545), .B(n544), .Z(n574) );
  NAND U598 ( .A(b[0]), .B(a[25]), .Z(n546) );
  XNOR U599 ( .A(b[1]), .B(n546), .Z(n548) );
  NANDN U600 ( .A(b[0]), .B(a[24]), .Z(n547) );
  NAND U601 ( .A(n548), .B(n547), .Z(n573) );
  AND U602 ( .A(b[3]), .B(a[21]), .Z(n572) );
  XOR U603 ( .A(n573), .B(n572), .Z(n575) );
  XOR U604 ( .A(n574), .B(n575), .Z(n561) );
  NANDN U605 ( .A(n550), .B(n549), .Z(n554) );
  OR U606 ( .A(n552), .B(n551), .Z(n553) );
  AND U607 ( .A(n554), .B(n553), .Z(n560) );
  XOR U608 ( .A(n561), .B(n560), .Z(n563) );
  XOR U609 ( .A(n562), .B(n563), .Z(n578) );
  XNOR U610 ( .A(n578), .B(sreg[277]), .Z(n580) );
  NANDN U611 ( .A(n555), .B(sreg[276]), .Z(n559) );
  NAND U612 ( .A(n557), .B(n556), .Z(n558) );
  NAND U613 ( .A(n559), .B(n558), .Z(n579) );
  XOR U614 ( .A(n580), .B(n579), .Z(c[277]) );
  NANDN U615 ( .A(n561), .B(n560), .Z(n565) );
  OR U616 ( .A(n563), .B(n562), .Z(n564) );
  AND U617 ( .A(n565), .B(n564), .Z(n585) );
  NAND U618 ( .A(n31), .B(n566), .Z(n568) );
  XOR U619 ( .A(b[3]), .B(a[24]), .Z(n589) );
  NAND U620 ( .A(n5811), .B(n589), .Z(n567) );
  AND U621 ( .A(n568), .B(n567), .Z(n597) );
  AND U622 ( .A(b[3]), .B(a[22]), .Z(n595) );
  NAND U623 ( .A(b[0]), .B(a[26]), .Z(n569) );
  XNOR U624 ( .A(b[1]), .B(n569), .Z(n571) );
  NANDN U625 ( .A(b[0]), .B(a[25]), .Z(n570) );
  NAND U626 ( .A(n571), .B(n570), .Z(n596) );
  XOR U627 ( .A(n595), .B(n596), .Z(n598) );
  XOR U628 ( .A(n597), .B(n598), .Z(n584) );
  NANDN U629 ( .A(n573), .B(n572), .Z(n577) );
  OR U630 ( .A(n575), .B(n574), .Z(n576) );
  AND U631 ( .A(n577), .B(n576), .Z(n583) );
  XOR U632 ( .A(n584), .B(n583), .Z(n586) );
  XOR U633 ( .A(n585), .B(n586), .Z(n601) );
  XNOR U634 ( .A(n601), .B(sreg[278]), .Z(n603) );
  NANDN U635 ( .A(n578), .B(sreg[277]), .Z(n582) );
  NAND U636 ( .A(n580), .B(n579), .Z(n581) );
  NAND U637 ( .A(n582), .B(n581), .Z(n602) );
  XOR U638 ( .A(n603), .B(n602), .Z(c[278]) );
  NANDN U639 ( .A(n584), .B(n583), .Z(n588) );
  OR U640 ( .A(n586), .B(n585), .Z(n587) );
  AND U641 ( .A(n588), .B(n587), .Z(n608) );
  NAND U642 ( .A(n31), .B(n589), .Z(n591) );
  XOR U643 ( .A(b[3]), .B(a[25]), .Z(n612) );
  NAND U644 ( .A(n5811), .B(n612), .Z(n590) );
  AND U645 ( .A(n591), .B(n590), .Z(n620) );
  NAND U646 ( .A(b[0]), .B(a[27]), .Z(n592) );
  XNOR U647 ( .A(b[1]), .B(n592), .Z(n594) );
  NANDN U648 ( .A(b[0]), .B(a[26]), .Z(n593) );
  NAND U649 ( .A(n594), .B(n593), .Z(n619) );
  AND U650 ( .A(b[3]), .B(a[23]), .Z(n618) );
  XOR U651 ( .A(n619), .B(n618), .Z(n621) );
  XOR U652 ( .A(n620), .B(n621), .Z(n607) );
  NANDN U653 ( .A(n596), .B(n595), .Z(n600) );
  OR U654 ( .A(n598), .B(n597), .Z(n599) );
  AND U655 ( .A(n600), .B(n599), .Z(n606) );
  XOR U656 ( .A(n607), .B(n606), .Z(n609) );
  XOR U657 ( .A(n608), .B(n609), .Z(n624) );
  XNOR U658 ( .A(n624), .B(sreg[279]), .Z(n626) );
  NANDN U659 ( .A(n601), .B(sreg[278]), .Z(n605) );
  NAND U660 ( .A(n603), .B(n602), .Z(n604) );
  NAND U661 ( .A(n605), .B(n604), .Z(n625) );
  XOR U662 ( .A(n626), .B(n625), .Z(c[279]) );
  NANDN U663 ( .A(n607), .B(n606), .Z(n611) );
  OR U664 ( .A(n609), .B(n608), .Z(n610) );
  AND U665 ( .A(n611), .B(n610), .Z(n631) );
  NAND U666 ( .A(n31), .B(n612), .Z(n614) );
  XOR U667 ( .A(b[3]), .B(a[26]), .Z(n635) );
  NAND U668 ( .A(n5811), .B(n635), .Z(n613) );
  AND U669 ( .A(n614), .B(n613), .Z(n643) );
  AND U670 ( .A(b[3]), .B(a[24]), .Z(n641) );
  NAND U671 ( .A(b[0]), .B(a[28]), .Z(n615) );
  XNOR U672 ( .A(b[1]), .B(n615), .Z(n617) );
  NANDN U673 ( .A(b[0]), .B(a[27]), .Z(n616) );
  NAND U674 ( .A(n617), .B(n616), .Z(n642) );
  XOR U675 ( .A(n641), .B(n642), .Z(n644) );
  XOR U676 ( .A(n643), .B(n644), .Z(n630) );
  NANDN U677 ( .A(n619), .B(n618), .Z(n623) );
  OR U678 ( .A(n621), .B(n620), .Z(n622) );
  AND U679 ( .A(n623), .B(n622), .Z(n629) );
  XOR U680 ( .A(n630), .B(n629), .Z(n632) );
  XOR U681 ( .A(n631), .B(n632), .Z(n647) );
  XNOR U682 ( .A(n647), .B(sreg[280]), .Z(n649) );
  NANDN U683 ( .A(n624), .B(sreg[279]), .Z(n628) );
  NAND U684 ( .A(n626), .B(n625), .Z(n627) );
  NAND U685 ( .A(n628), .B(n627), .Z(n648) );
  XOR U686 ( .A(n649), .B(n648), .Z(c[280]) );
  NANDN U687 ( .A(n630), .B(n629), .Z(n634) );
  OR U688 ( .A(n632), .B(n631), .Z(n633) );
  AND U689 ( .A(n634), .B(n633), .Z(n654) );
  NAND U690 ( .A(n31), .B(n635), .Z(n637) );
  XOR U691 ( .A(b[3]), .B(a[27]), .Z(n658) );
  NAND U692 ( .A(n5811), .B(n658), .Z(n636) );
  AND U693 ( .A(n637), .B(n636), .Z(n666) );
  AND U694 ( .A(b[3]), .B(a[25]), .Z(n664) );
  NAND U695 ( .A(b[0]), .B(a[29]), .Z(n638) );
  XNOR U696 ( .A(b[1]), .B(n638), .Z(n640) );
  NANDN U697 ( .A(b[0]), .B(a[28]), .Z(n639) );
  NAND U698 ( .A(n640), .B(n639), .Z(n665) );
  XOR U699 ( .A(n664), .B(n665), .Z(n667) );
  XOR U700 ( .A(n666), .B(n667), .Z(n653) );
  NANDN U701 ( .A(n642), .B(n641), .Z(n646) );
  OR U702 ( .A(n644), .B(n643), .Z(n645) );
  AND U703 ( .A(n646), .B(n645), .Z(n652) );
  XOR U704 ( .A(n653), .B(n652), .Z(n655) );
  XOR U705 ( .A(n654), .B(n655), .Z(n670) );
  XNOR U706 ( .A(n670), .B(sreg[281]), .Z(n672) );
  NANDN U707 ( .A(n647), .B(sreg[280]), .Z(n651) );
  NAND U708 ( .A(n649), .B(n648), .Z(n650) );
  NAND U709 ( .A(n651), .B(n650), .Z(n671) );
  XOR U710 ( .A(n672), .B(n671), .Z(c[281]) );
  NANDN U711 ( .A(n653), .B(n652), .Z(n657) );
  OR U712 ( .A(n655), .B(n654), .Z(n656) );
  AND U713 ( .A(n657), .B(n656), .Z(n677) );
  NAND U714 ( .A(n31), .B(n658), .Z(n660) );
  XOR U715 ( .A(b[3]), .B(a[28]), .Z(n681) );
  NAND U716 ( .A(n5811), .B(n681), .Z(n659) );
  AND U717 ( .A(n660), .B(n659), .Z(n689) );
  NAND U718 ( .A(b[0]), .B(a[30]), .Z(n661) );
  XNOR U719 ( .A(b[1]), .B(n661), .Z(n663) );
  NANDN U720 ( .A(b[0]), .B(a[29]), .Z(n662) );
  NAND U721 ( .A(n663), .B(n662), .Z(n688) );
  AND U722 ( .A(b[3]), .B(a[26]), .Z(n687) );
  XOR U723 ( .A(n688), .B(n687), .Z(n690) );
  XOR U724 ( .A(n689), .B(n690), .Z(n676) );
  NANDN U725 ( .A(n665), .B(n664), .Z(n669) );
  OR U726 ( .A(n667), .B(n666), .Z(n668) );
  AND U727 ( .A(n669), .B(n668), .Z(n675) );
  XOR U728 ( .A(n676), .B(n675), .Z(n678) );
  XOR U729 ( .A(n677), .B(n678), .Z(n693) );
  XNOR U730 ( .A(n693), .B(sreg[282]), .Z(n695) );
  NANDN U731 ( .A(n670), .B(sreg[281]), .Z(n674) );
  NAND U732 ( .A(n672), .B(n671), .Z(n673) );
  NAND U733 ( .A(n674), .B(n673), .Z(n694) );
  XOR U734 ( .A(n695), .B(n694), .Z(c[282]) );
  NANDN U735 ( .A(n676), .B(n675), .Z(n680) );
  OR U736 ( .A(n678), .B(n677), .Z(n679) );
  AND U737 ( .A(n680), .B(n679), .Z(n700) );
  NAND U738 ( .A(n31), .B(n681), .Z(n683) );
  XOR U739 ( .A(b[3]), .B(a[29]), .Z(n704) );
  NAND U740 ( .A(n5811), .B(n704), .Z(n682) );
  AND U741 ( .A(n683), .B(n682), .Z(n712) );
  NAND U742 ( .A(b[0]), .B(a[31]), .Z(n684) );
  XNOR U743 ( .A(b[1]), .B(n684), .Z(n686) );
  NANDN U744 ( .A(b[0]), .B(a[30]), .Z(n685) );
  NAND U745 ( .A(n686), .B(n685), .Z(n711) );
  AND U746 ( .A(b[3]), .B(a[27]), .Z(n710) );
  XOR U747 ( .A(n711), .B(n710), .Z(n713) );
  XOR U748 ( .A(n712), .B(n713), .Z(n699) );
  NANDN U749 ( .A(n688), .B(n687), .Z(n692) );
  OR U750 ( .A(n690), .B(n689), .Z(n691) );
  AND U751 ( .A(n692), .B(n691), .Z(n698) );
  XOR U752 ( .A(n699), .B(n698), .Z(n701) );
  XOR U753 ( .A(n700), .B(n701), .Z(n716) );
  XNOR U754 ( .A(n716), .B(sreg[283]), .Z(n718) );
  NANDN U755 ( .A(n693), .B(sreg[282]), .Z(n697) );
  NAND U756 ( .A(n695), .B(n694), .Z(n696) );
  NAND U757 ( .A(n697), .B(n696), .Z(n717) );
  XOR U758 ( .A(n718), .B(n717), .Z(c[283]) );
  NANDN U759 ( .A(n699), .B(n698), .Z(n703) );
  OR U760 ( .A(n701), .B(n700), .Z(n702) );
  AND U761 ( .A(n703), .B(n702), .Z(n723) );
  NAND U762 ( .A(n31), .B(n704), .Z(n706) );
  XOR U763 ( .A(b[3]), .B(a[30]), .Z(n727) );
  NAND U764 ( .A(n5811), .B(n727), .Z(n705) );
  AND U765 ( .A(n706), .B(n705), .Z(n735) );
  NAND U766 ( .A(b[0]), .B(a[32]), .Z(n707) );
  XNOR U767 ( .A(b[1]), .B(n707), .Z(n709) );
  NANDN U768 ( .A(b[0]), .B(a[31]), .Z(n708) );
  NAND U769 ( .A(n709), .B(n708), .Z(n734) );
  AND U770 ( .A(b[3]), .B(a[28]), .Z(n733) );
  XOR U771 ( .A(n734), .B(n733), .Z(n736) );
  XOR U772 ( .A(n735), .B(n736), .Z(n722) );
  NANDN U773 ( .A(n711), .B(n710), .Z(n715) );
  OR U774 ( .A(n713), .B(n712), .Z(n714) );
  AND U775 ( .A(n715), .B(n714), .Z(n721) );
  XOR U776 ( .A(n722), .B(n721), .Z(n724) );
  XOR U777 ( .A(n723), .B(n724), .Z(n739) );
  XNOR U778 ( .A(n739), .B(sreg[284]), .Z(n741) );
  NANDN U779 ( .A(n716), .B(sreg[283]), .Z(n720) );
  NAND U780 ( .A(n718), .B(n717), .Z(n719) );
  NAND U781 ( .A(n720), .B(n719), .Z(n740) );
  XOR U782 ( .A(n741), .B(n740), .Z(c[284]) );
  NANDN U783 ( .A(n722), .B(n721), .Z(n726) );
  OR U784 ( .A(n724), .B(n723), .Z(n725) );
  AND U785 ( .A(n726), .B(n725), .Z(n746) );
  NAND U786 ( .A(n31), .B(n727), .Z(n729) );
  XOR U787 ( .A(b[3]), .B(a[31]), .Z(n750) );
  NAND U788 ( .A(n5811), .B(n750), .Z(n728) );
  AND U789 ( .A(n729), .B(n728), .Z(n758) );
  AND U790 ( .A(b[3]), .B(a[29]), .Z(n756) );
  NAND U791 ( .A(b[0]), .B(a[33]), .Z(n730) );
  XNOR U792 ( .A(b[1]), .B(n730), .Z(n732) );
  NANDN U793 ( .A(b[0]), .B(a[32]), .Z(n731) );
  NAND U794 ( .A(n732), .B(n731), .Z(n757) );
  XOR U795 ( .A(n756), .B(n757), .Z(n759) );
  XOR U796 ( .A(n758), .B(n759), .Z(n745) );
  NANDN U797 ( .A(n734), .B(n733), .Z(n738) );
  OR U798 ( .A(n736), .B(n735), .Z(n737) );
  AND U799 ( .A(n738), .B(n737), .Z(n744) );
  XOR U800 ( .A(n745), .B(n744), .Z(n747) );
  XOR U801 ( .A(n746), .B(n747), .Z(n762) );
  XNOR U802 ( .A(n762), .B(sreg[285]), .Z(n764) );
  NANDN U803 ( .A(n739), .B(sreg[284]), .Z(n743) );
  NAND U804 ( .A(n741), .B(n740), .Z(n742) );
  NAND U805 ( .A(n743), .B(n742), .Z(n763) );
  XOR U806 ( .A(n764), .B(n763), .Z(c[285]) );
  NANDN U807 ( .A(n745), .B(n744), .Z(n749) );
  OR U808 ( .A(n747), .B(n746), .Z(n748) );
  AND U809 ( .A(n749), .B(n748), .Z(n769) );
  NAND U810 ( .A(n31), .B(n750), .Z(n752) );
  XOR U811 ( .A(b[3]), .B(a[32]), .Z(n773) );
  NAND U812 ( .A(n5811), .B(n773), .Z(n751) );
  AND U813 ( .A(n752), .B(n751), .Z(n781) );
  NAND U814 ( .A(b[0]), .B(a[34]), .Z(n753) );
  XNOR U815 ( .A(b[1]), .B(n753), .Z(n755) );
  NANDN U816 ( .A(b[0]), .B(a[33]), .Z(n754) );
  NAND U817 ( .A(n755), .B(n754), .Z(n780) );
  AND U818 ( .A(b[3]), .B(a[30]), .Z(n779) );
  XOR U819 ( .A(n780), .B(n779), .Z(n782) );
  XOR U820 ( .A(n781), .B(n782), .Z(n768) );
  NANDN U821 ( .A(n757), .B(n756), .Z(n761) );
  OR U822 ( .A(n759), .B(n758), .Z(n760) );
  AND U823 ( .A(n761), .B(n760), .Z(n767) );
  XOR U824 ( .A(n768), .B(n767), .Z(n770) );
  XOR U825 ( .A(n769), .B(n770), .Z(n785) );
  XNOR U826 ( .A(n785), .B(sreg[286]), .Z(n787) );
  NANDN U827 ( .A(n762), .B(sreg[285]), .Z(n766) );
  NAND U828 ( .A(n764), .B(n763), .Z(n765) );
  NAND U829 ( .A(n766), .B(n765), .Z(n786) );
  XOR U830 ( .A(n787), .B(n786), .Z(c[286]) );
  NANDN U831 ( .A(n768), .B(n767), .Z(n772) );
  OR U832 ( .A(n770), .B(n769), .Z(n771) );
  AND U833 ( .A(n772), .B(n771), .Z(n792) );
  NAND U834 ( .A(n31), .B(n773), .Z(n775) );
  XOR U835 ( .A(b[3]), .B(a[33]), .Z(n796) );
  NAND U836 ( .A(n5811), .B(n796), .Z(n774) );
  AND U837 ( .A(n775), .B(n774), .Z(n804) );
  NAND U838 ( .A(b[0]), .B(a[35]), .Z(n776) );
  XNOR U839 ( .A(b[1]), .B(n776), .Z(n778) );
  NANDN U840 ( .A(b[0]), .B(a[34]), .Z(n777) );
  NAND U841 ( .A(n778), .B(n777), .Z(n803) );
  AND U842 ( .A(b[3]), .B(a[31]), .Z(n802) );
  XOR U843 ( .A(n803), .B(n802), .Z(n805) );
  XOR U844 ( .A(n804), .B(n805), .Z(n791) );
  NANDN U845 ( .A(n780), .B(n779), .Z(n784) );
  OR U846 ( .A(n782), .B(n781), .Z(n783) );
  AND U847 ( .A(n784), .B(n783), .Z(n790) );
  XOR U848 ( .A(n791), .B(n790), .Z(n793) );
  XOR U849 ( .A(n792), .B(n793), .Z(n808) );
  XNOR U850 ( .A(n808), .B(sreg[287]), .Z(n810) );
  NANDN U851 ( .A(n785), .B(sreg[286]), .Z(n789) );
  NAND U852 ( .A(n787), .B(n786), .Z(n788) );
  NAND U853 ( .A(n789), .B(n788), .Z(n809) );
  XOR U854 ( .A(n810), .B(n809), .Z(c[287]) );
  NANDN U855 ( .A(n791), .B(n790), .Z(n795) );
  OR U856 ( .A(n793), .B(n792), .Z(n794) );
  AND U857 ( .A(n795), .B(n794), .Z(n815) );
  NAND U858 ( .A(n31), .B(n796), .Z(n798) );
  XOR U859 ( .A(b[3]), .B(a[34]), .Z(n819) );
  NAND U860 ( .A(n5811), .B(n819), .Z(n797) );
  AND U861 ( .A(n798), .B(n797), .Z(n827) );
  AND U862 ( .A(b[3]), .B(a[32]), .Z(n825) );
  NAND U863 ( .A(b[0]), .B(a[36]), .Z(n799) );
  XNOR U864 ( .A(b[1]), .B(n799), .Z(n801) );
  NANDN U865 ( .A(b[0]), .B(a[35]), .Z(n800) );
  NAND U866 ( .A(n801), .B(n800), .Z(n826) );
  XOR U867 ( .A(n825), .B(n826), .Z(n828) );
  XOR U868 ( .A(n827), .B(n828), .Z(n814) );
  NANDN U869 ( .A(n803), .B(n802), .Z(n807) );
  OR U870 ( .A(n805), .B(n804), .Z(n806) );
  AND U871 ( .A(n807), .B(n806), .Z(n813) );
  XOR U872 ( .A(n814), .B(n813), .Z(n816) );
  XOR U873 ( .A(n815), .B(n816), .Z(n831) );
  XNOR U874 ( .A(n831), .B(sreg[288]), .Z(n833) );
  NANDN U875 ( .A(n808), .B(sreg[287]), .Z(n812) );
  NAND U876 ( .A(n810), .B(n809), .Z(n811) );
  NAND U877 ( .A(n812), .B(n811), .Z(n832) );
  XOR U878 ( .A(n833), .B(n832), .Z(c[288]) );
  NANDN U879 ( .A(n814), .B(n813), .Z(n818) );
  OR U880 ( .A(n816), .B(n815), .Z(n817) );
  AND U881 ( .A(n818), .B(n817), .Z(n838) );
  NAND U882 ( .A(n31), .B(n819), .Z(n821) );
  XOR U883 ( .A(b[3]), .B(a[35]), .Z(n842) );
  NAND U884 ( .A(n5811), .B(n842), .Z(n820) );
  AND U885 ( .A(n821), .B(n820), .Z(n850) );
  NAND U886 ( .A(b[0]), .B(a[37]), .Z(n822) );
  XNOR U887 ( .A(b[1]), .B(n822), .Z(n824) );
  NANDN U888 ( .A(b[0]), .B(a[36]), .Z(n823) );
  NAND U889 ( .A(n824), .B(n823), .Z(n849) );
  AND U890 ( .A(b[3]), .B(a[33]), .Z(n848) );
  XOR U891 ( .A(n849), .B(n848), .Z(n851) );
  XOR U892 ( .A(n850), .B(n851), .Z(n837) );
  NANDN U893 ( .A(n826), .B(n825), .Z(n830) );
  OR U894 ( .A(n828), .B(n827), .Z(n829) );
  AND U895 ( .A(n830), .B(n829), .Z(n836) );
  XOR U896 ( .A(n837), .B(n836), .Z(n839) );
  XOR U897 ( .A(n838), .B(n839), .Z(n854) );
  XNOR U898 ( .A(n854), .B(sreg[289]), .Z(n856) );
  NANDN U899 ( .A(n831), .B(sreg[288]), .Z(n835) );
  NAND U900 ( .A(n833), .B(n832), .Z(n834) );
  NAND U901 ( .A(n835), .B(n834), .Z(n855) );
  XOR U902 ( .A(n856), .B(n855), .Z(c[289]) );
  NANDN U903 ( .A(n837), .B(n836), .Z(n841) );
  OR U904 ( .A(n839), .B(n838), .Z(n840) );
  AND U905 ( .A(n841), .B(n840), .Z(n861) );
  NAND U906 ( .A(n31), .B(n842), .Z(n844) );
  XOR U907 ( .A(b[3]), .B(a[36]), .Z(n865) );
  NAND U908 ( .A(n5811), .B(n865), .Z(n843) );
  AND U909 ( .A(n844), .B(n843), .Z(n873) );
  NAND U910 ( .A(b[0]), .B(a[38]), .Z(n845) );
  XNOR U911 ( .A(b[1]), .B(n845), .Z(n847) );
  NANDN U912 ( .A(b[0]), .B(a[37]), .Z(n846) );
  NAND U913 ( .A(n847), .B(n846), .Z(n872) );
  AND U914 ( .A(b[3]), .B(a[34]), .Z(n871) );
  XOR U915 ( .A(n872), .B(n871), .Z(n874) );
  XOR U916 ( .A(n873), .B(n874), .Z(n860) );
  NANDN U917 ( .A(n849), .B(n848), .Z(n853) );
  OR U918 ( .A(n851), .B(n850), .Z(n852) );
  AND U919 ( .A(n853), .B(n852), .Z(n859) );
  XOR U920 ( .A(n860), .B(n859), .Z(n862) );
  XOR U921 ( .A(n861), .B(n862), .Z(n877) );
  XNOR U922 ( .A(n877), .B(sreg[290]), .Z(n879) );
  NANDN U923 ( .A(n854), .B(sreg[289]), .Z(n858) );
  NAND U924 ( .A(n856), .B(n855), .Z(n857) );
  NAND U925 ( .A(n858), .B(n857), .Z(n878) );
  XOR U926 ( .A(n879), .B(n878), .Z(c[290]) );
  NANDN U927 ( .A(n860), .B(n859), .Z(n864) );
  OR U928 ( .A(n862), .B(n861), .Z(n863) );
  AND U929 ( .A(n864), .B(n863), .Z(n884) );
  NAND U930 ( .A(n31), .B(n865), .Z(n867) );
  XOR U931 ( .A(b[3]), .B(a[37]), .Z(n888) );
  NAND U932 ( .A(n5811), .B(n888), .Z(n866) );
  AND U933 ( .A(n867), .B(n866), .Z(n896) );
  AND U934 ( .A(b[3]), .B(a[35]), .Z(n894) );
  NAND U935 ( .A(b[0]), .B(a[39]), .Z(n868) );
  XNOR U936 ( .A(b[1]), .B(n868), .Z(n870) );
  NANDN U937 ( .A(b[0]), .B(a[38]), .Z(n869) );
  NAND U938 ( .A(n870), .B(n869), .Z(n895) );
  XOR U939 ( .A(n894), .B(n895), .Z(n897) );
  XOR U940 ( .A(n896), .B(n897), .Z(n883) );
  NANDN U941 ( .A(n872), .B(n871), .Z(n876) );
  OR U942 ( .A(n874), .B(n873), .Z(n875) );
  AND U943 ( .A(n876), .B(n875), .Z(n882) );
  XOR U944 ( .A(n883), .B(n882), .Z(n885) );
  XOR U945 ( .A(n884), .B(n885), .Z(n900) );
  XNOR U946 ( .A(n900), .B(sreg[291]), .Z(n902) );
  NANDN U947 ( .A(n877), .B(sreg[290]), .Z(n881) );
  NAND U948 ( .A(n879), .B(n878), .Z(n880) );
  NAND U949 ( .A(n881), .B(n880), .Z(n901) );
  XOR U950 ( .A(n902), .B(n901), .Z(c[291]) );
  NANDN U951 ( .A(n883), .B(n882), .Z(n887) );
  OR U952 ( .A(n885), .B(n884), .Z(n886) );
  AND U953 ( .A(n887), .B(n886), .Z(n907) );
  NAND U954 ( .A(n31), .B(n888), .Z(n890) );
  XOR U955 ( .A(b[3]), .B(a[38]), .Z(n911) );
  NAND U956 ( .A(n5811), .B(n911), .Z(n889) );
  AND U957 ( .A(n890), .B(n889), .Z(n919) );
  NAND U958 ( .A(b[0]), .B(a[40]), .Z(n891) );
  XNOR U959 ( .A(b[1]), .B(n891), .Z(n893) );
  NANDN U960 ( .A(b[0]), .B(a[39]), .Z(n892) );
  NAND U961 ( .A(n893), .B(n892), .Z(n918) );
  AND U962 ( .A(b[3]), .B(a[36]), .Z(n917) );
  XOR U963 ( .A(n918), .B(n917), .Z(n920) );
  XOR U964 ( .A(n919), .B(n920), .Z(n906) );
  NANDN U965 ( .A(n895), .B(n894), .Z(n899) );
  OR U966 ( .A(n897), .B(n896), .Z(n898) );
  AND U967 ( .A(n899), .B(n898), .Z(n905) );
  XOR U968 ( .A(n906), .B(n905), .Z(n908) );
  XOR U969 ( .A(n907), .B(n908), .Z(n923) );
  XNOR U970 ( .A(n923), .B(sreg[292]), .Z(n925) );
  NANDN U971 ( .A(n900), .B(sreg[291]), .Z(n904) );
  NAND U972 ( .A(n902), .B(n901), .Z(n903) );
  NAND U973 ( .A(n904), .B(n903), .Z(n924) );
  XOR U974 ( .A(n925), .B(n924), .Z(c[292]) );
  NANDN U975 ( .A(n906), .B(n905), .Z(n910) );
  OR U976 ( .A(n908), .B(n907), .Z(n909) );
  AND U977 ( .A(n910), .B(n909), .Z(n930) );
  NAND U978 ( .A(n31), .B(n911), .Z(n913) );
  XOR U979 ( .A(b[3]), .B(a[39]), .Z(n934) );
  NAND U980 ( .A(n5811), .B(n934), .Z(n912) );
  AND U981 ( .A(n913), .B(n912), .Z(n942) );
  NAND U982 ( .A(b[0]), .B(a[41]), .Z(n914) );
  XNOR U983 ( .A(b[1]), .B(n914), .Z(n916) );
  NANDN U984 ( .A(b[0]), .B(a[40]), .Z(n915) );
  NAND U985 ( .A(n916), .B(n915), .Z(n941) );
  AND U986 ( .A(b[3]), .B(a[37]), .Z(n940) );
  XOR U987 ( .A(n941), .B(n940), .Z(n943) );
  XOR U988 ( .A(n942), .B(n943), .Z(n929) );
  NANDN U989 ( .A(n918), .B(n917), .Z(n922) );
  OR U990 ( .A(n920), .B(n919), .Z(n921) );
  AND U991 ( .A(n922), .B(n921), .Z(n928) );
  XOR U992 ( .A(n929), .B(n928), .Z(n931) );
  XOR U993 ( .A(n930), .B(n931), .Z(n946) );
  XNOR U994 ( .A(n946), .B(sreg[293]), .Z(n948) );
  NANDN U995 ( .A(n923), .B(sreg[292]), .Z(n927) );
  NAND U996 ( .A(n925), .B(n924), .Z(n926) );
  NAND U997 ( .A(n927), .B(n926), .Z(n947) );
  XOR U998 ( .A(n948), .B(n947), .Z(c[293]) );
  NANDN U999 ( .A(n929), .B(n928), .Z(n933) );
  OR U1000 ( .A(n931), .B(n930), .Z(n932) );
  AND U1001 ( .A(n933), .B(n932), .Z(n953) );
  NAND U1002 ( .A(n31), .B(n934), .Z(n936) );
  XOR U1003 ( .A(b[3]), .B(a[40]), .Z(n957) );
  NAND U1004 ( .A(n5811), .B(n957), .Z(n935) );
  AND U1005 ( .A(n936), .B(n935), .Z(n965) );
  NAND U1006 ( .A(b[0]), .B(a[42]), .Z(n937) );
  XNOR U1007 ( .A(b[1]), .B(n937), .Z(n939) );
  NANDN U1008 ( .A(b[0]), .B(a[41]), .Z(n938) );
  NAND U1009 ( .A(n939), .B(n938), .Z(n964) );
  AND U1010 ( .A(b[3]), .B(a[38]), .Z(n963) );
  XOR U1011 ( .A(n964), .B(n963), .Z(n966) );
  XOR U1012 ( .A(n965), .B(n966), .Z(n952) );
  NANDN U1013 ( .A(n941), .B(n940), .Z(n945) );
  OR U1014 ( .A(n943), .B(n942), .Z(n944) );
  AND U1015 ( .A(n945), .B(n944), .Z(n951) );
  XOR U1016 ( .A(n952), .B(n951), .Z(n954) );
  XOR U1017 ( .A(n953), .B(n954), .Z(n969) );
  XNOR U1018 ( .A(n969), .B(sreg[294]), .Z(n971) );
  NANDN U1019 ( .A(n946), .B(sreg[293]), .Z(n950) );
  NAND U1020 ( .A(n948), .B(n947), .Z(n949) );
  NAND U1021 ( .A(n950), .B(n949), .Z(n970) );
  XOR U1022 ( .A(n971), .B(n970), .Z(c[294]) );
  NANDN U1023 ( .A(n952), .B(n951), .Z(n956) );
  OR U1024 ( .A(n954), .B(n953), .Z(n955) );
  AND U1025 ( .A(n956), .B(n955), .Z(n976) );
  NAND U1026 ( .A(n31), .B(n957), .Z(n959) );
  XOR U1027 ( .A(b[3]), .B(a[41]), .Z(n980) );
  NAND U1028 ( .A(n5811), .B(n980), .Z(n958) );
  AND U1029 ( .A(n959), .B(n958), .Z(n988) );
  AND U1030 ( .A(b[3]), .B(a[39]), .Z(n986) );
  NAND U1031 ( .A(b[0]), .B(a[43]), .Z(n960) );
  XNOR U1032 ( .A(b[1]), .B(n960), .Z(n962) );
  NANDN U1033 ( .A(b[0]), .B(a[42]), .Z(n961) );
  NAND U1034 ( .A(n962), .B(n961), .Z(n987) );
  XOR U1035 ( .A(n986), .B(n987), .Z(n989) );
  XOR U1036 ( .A(n988), .B(n989), .Z(n975) );
  NANDN U1037 ( .A(n964), .B(n963), .Z(n968) );
  OR U1038 ( .A(n966), .B(n965), .Z(n967) );
  AND U1039 ( .A(n968), .B(n967), .Z(n974) );
  XOR U1040 ( .A(n975), .B(n974), .Z(n977) );
  XOR U1041 ( .A(n976), .B(n977), .Z(n992) );
  XNOR U1042 ( .A(n992), .B(sreg[295]), .Z(n994) );
  NANDN U1043 ( .A(n969), .B(sreg[294]), .Z(n973) );
  NAND U1044 ( .A(n971), .B(n970), .Z(n972) );
  NAND U1045 ( .A(n973), .B(n972), .Z(n993) );
  XOR U1046 ( .A(n994), .B(n993), .Z(c[295]) );
  NANDN U1047 ( .A(n975), .B(n974), .Z(n979) );
  OR U1048 ( .A(n977), .B(n976), .Z(n978) );
  AND U1049 ( .A(n979), .B(n978), .Z(n999) );
  NAND U1050 ( .A(n31), .B(n980), .Z(n982) );
  XOR U1051 ( .A(b[3]), .B(a[42]), .Z(n1003) );
  NAND U1052 ( .A(n5811), .B(n1003), .Z(n981) );
  AND U1053 ( .A(n982), .B(n981), .Z(n1011) );
  NAND U1054 ( .A(b[0]), .B(a[44]), .Z(n983) );
  XNOR U1055 ( .A(b[1]), .B(n983), .Z(n985) );
  NANDN U1056 ( .A(b[0]), .B(a[43]), .Z(n984) );
  NAND U1057 ( .A(n985), .B(n984), .Z(n1010) );
  AND U1058 ( .A(b[3]), .B(a[40]), .Z(n1009) );
  XOR U1059 ( .A(n1010), .B(n1009), .Z(n1012) );
  XOR U1060 ( .A(n1011), .B(n1012), .Z(n998) );
  NANDN U1061 ( .A(n987), .B(n986), .Z(n991) );
  OR U1062 ( .A(n989), .B(n988), .Z(n990) );
  AND U1063 ( .A(n991), .B(n990), .Z(n997) );
  XOR U1064 ( .A(n998), .B(n997), .Z(n1000) );
  XOR U1065 ( .A(n999), .B(n1000), .Z(n1015) );
  XNOR U1066 ( .A(n1015), .B(sreg[296]), .Z(n1017) );
  NANDN U1067 ( .A(n992), .B(sreg[295]), .Z(n996) );
  NAND U1068 ( .A(n994), .B(n993), .Z(n995) );
  NAND U1069 ( .A(n996), .B(n995), .Z(n1016) );
  XOR U1070 ( .A(n1017), .B(n1016), .Z(c[296]) );
  NANDN U1071 ( .A(n998), .B(n997), .Z(n1002) );
  OR U1072 ( .A(n1000), .B(n999), .Z(n1001) );
  AND U1073 ( .A(n1002), .B(n1001), .Z(n1022) );
  NAND U1074 ( .A(n31), .B(n1003), .Z(n1005) );
  XOR U1075 ( .A(b[3]), .B(a[43]), .Z(n1026) );
  NAND U1076 ( .A(n5811), .B(n1026), .Z(n1004) );
  AND U1077 ( .A(n1005), .B(n1004), .Z(n1034) );
  NAND U1078 ( .A(b[0]), .B(a[45]), .Z(n1006) );
  XNOR U1079 ( .A(b[1]), .B(n1006), .Z(n1008) );
  NANDN U1080 ( .A(b[0]), .B(a[44]), .Z(n1007) );
  NAND U1081 ( .A(n1008), .B(n1007), .Z(n1033) );
  AND U1082 ( .A(b[3]), .B(a[41]), .Z(n1032) );
  XOR U1083 ( .A(n1033), .B(n1032), .Z(n1035) );
  XOR U1084 ( .A(n1034), .B(n1035), .Z(n1021) );
  NANDN U1085 ( .A(n1010), .B(n1009), .Z(n1014) );
  OR U1086 ( .A(n1012), .B(n1011), .Z(n1013) );
  AND U1087 ( .A(n1014), .B(n1013), .Z(n1020) );
  XOR U1088 ( .A(n1021), .B(n1020), .Z(n1023) );
  XOR U1089 ( .A(n1022), .B(n1023), .Z(n1038) );
  XNOR U1090 ( .A(n1038), .B(sreg[297]), .Z(n1040) );
  NANDN U1091 ( .A(n1015), .B(sreg[296]), .Z(n1019) );
  NAND U1092 ( .A(n1017), .B(n1016), .Z(n1018) );
  NAND U1093 ( .A(n1019), .B(n1018), .Z(n1039) );
  XOR U1094 ( .A(n1040), .B(n1039), .Z(c[297]) );
  NANDN U1095 ( .A(n1021), .B(n1020), .Z(n1025) );
  OR U1096 ( .A(n1023), .B(n1022), .Z(n1024) );
  AND U1097 ( .A(n1025), .B(n1024), .Z(n1045) );
  NAND U1098 ( .A(n31), .B(n1026), .Z(n1028) );
  XOR U1099 ( .A(b[3]), .B(a[44]), .Z(n1049) );
  NAND U1100 ( .A(n5811), .B(n1049), .Z(n1027) );
  AND U1101 ( .A(n1028), .B(n1027), .Z(n1057) );
  NAND U1102 ( .A(b[0]), .B(a[46]), .Z(n1029) );
  XNOR U1103 ( .A(b[1]), .B(n1029), .Z(n1031) );
  NANDN U1104 ( .A(b[0]), .B(a[45]), .Z(n1030) );
  NAND U1105 ( .A(n1031), .B(n1030), .Z(n1056) );
  AND U1106 ( .A(b[3]), .B(a[42]), .Z(n1055) );
  XOR U1107 ( .A(n1056), .B(n1055), .Z(n1058) );
  XOR U1108 ( .A(n1057), .B(n1058), .Z(n1044) );
  NANDN U1109 ( .A(n1033), .B(n1032), .Z(n1037) );
  OR U1110 ( .A(n1035), .B(n1034), .Z(n1036) );
  AND U1111 ( .A(n1037), .B(n1036), .Z(n1043) );
  XOR U1112 ( .A(n1044), .B(n1043), .Z(n1046) );
  XOR U1113 ( .A(n1045), .B(n1046), .Z(n1061) );
  XNOR U1114 ( .A(n1061), .B(sreg[298]), .Z(n1063) );
  NANDN U1115 ( .A(n1038), .B(sreg[297]), .Z(n1042) );
  NAND U1116 ( .A(n1040), .B(n1039), .Z(n1041) );
  NAND U1117 ( .A(n1042), .B(n1041), .Z(n1062) );
  XOR U1118 ( .A(n1063), .B(n1062), .Z(c[298]) );
  NANDN U1119 ( .A(n1044), .B(n1043), .Z(n1048) );
  OR U1120 ( .A(n1046), .B(n1045), .Z(n1047) );
  AND U1121 ( .A(n1048), .B(n1047), .Z(n1068) );
  NAND U1122 ( .A(n31), .B(n1049), .Z(n1051) );
  XOR U1123 ( .A(b[3]), .B(a[45]), .Z(n1072) );
  NAND U1124 ( .A(n5811), .B(n1072), .Z(n1050) );
  AND U1125 ( .A(n1051), .B(n1050), .Z(n1080) );
  NAND U1126 ( .A(b[0]), .B(a[47]), .Z(n1052) );
  XNOR U1127 ( .A(b[1]), .B(n1052), .Z(n1054) );
  NANDN U1128 ( .A(b[0]), .B(a[46]), .Z(n1053) );
  NAND U1129 ( .A(n1054), .B(n1053), .Z(n1079) );
  AND U1130 ( .A(b[3]), .B(a[43]), .Z(n1078) );
  XOR U1131 ( .A(n1079), .B(n1078), .Z(n1081) );
  XOR U1132 ( .A(n1080), .B(n1081), .Z(n1067) );
  NANDN U1133 ( .A(n1056), .B(n1055), .Z(n1060) );
  OR U1134 ( .A(n1058), .B(n1057), .Z(n1059) );
  AND U1135 ( .A(n1060), .B(n1059), .Z(n1066) );
  XOR U1136 ( .A(n1067), .B(n1066), .Z(n1069) );
  XOR U1137 ( .A(n1068), .B(n1069), .Z(n1084) );
  XNOR U1138 ( .A(n1084), .B(sreg[299]), .Z(n1086) );
  NANDN U1139 ( .A(n1061), .B(sreg[298]), .Z(n1065) );
  NAND U1140 ( .A(n1063), .B(n1062), .Z(n1064) );
  NAND U1141 ( .A(n1065), .B(n1064), .Z(n1085) );
  XOR U1142 ( .A(n1086), .B(n1085), .Z(c[299]) );
  NANDN U1143 ( .A(n1067), .B(n1066), .Z(n1071) );
  OR U1144 ( .A(n1069), .B(n1068), .Z(n1070) );
  AND U1145 ( .A(n1071), .B(n1070), .Z(n1091) );
  NAND U1146 ( .A(n31), .B(n1072), .Z(n1074) );
  XOR U1147 ( .A(b[3]), .B(a[46]), .Z(n1095) );
  NAND U1148 ( .A(n5811), .B(n1095), .Z(n1073) );
  AND U1149 ( .A(n1074), .B(n1073), .Z(n1103) );
  AND U1150 ( .A(b[3]), .B(a[44]), .Z(n1101) );
  NAND U1151 ( .A(b[0]), .B(a[48]), .Z(n1075) );
  XNOR U1152 ( .A(b[1]), .B(n1075), .Z(n1077) );
  NANDN U1153 ( .A(b[0]), .B(a[47]), .Z(n1076) );
  NAND U1154 ( .A(n1077), .B(n1076), .Z(n1102) );
  XOR U1155 ( .A(n1101), .B(n1102), .Z(n1104) );
  XOR U1156 ( .A(n1103), .B(n1104), .Z(n1090) );
  NANDN U1157 ( .A(n1079), .B(n1078), .Z(n1083) );
  OR U1158 ( .A(n1081), .B(n1080), .Z(n1082) );
  AND U1159 ( .A(n1083), .B(n1082), .Z(n1089) );
  XOR U1160 ( .A(n1090), .B(n1089), .Z(n1092) );
  XOR U1161 ( .A(n1091), .B(n1092), .Z(n1107) );
  XNOR U1162 ( .A(n1107), .B(sreg[300]), .Z(n1109) );
  NANDN U1163 ( .A(n1084), .B(sreg[299]), .Z(n1088) );
  NAND U1164 ( .A(n1086), .B(n1085), .Z(n1087) );
  NAND U1165 ( .A(n1088), .B(n1087), .Z(n1108) );
  XOR U1166 ( .A(n1109), .B(n1108), .Z(c[300]) );
  NANDN U1167 ( .A(n1090), .B(n1089), .Z(n1094) );
  OR U1168 ( .A(n1092), .B(n1091), .Z(n1093) );
  AND U1169 ( .A(n1094), .B(n1093), .Z(n1114) );
  NAND U1170 ( .A(n31), .B(n1095), .Z(n1097) );
  XOR U1171 ( .A(b[3]), .B(a[47]), .Z(n1118) );
  NAND U1172 ( .A(n5811), .B(n1118), .Z(n1096) );
  AND U1173 ( .A(n1097), .B(n1096), .Z(n1126) );
  NAND U1174 ( .A(b[0]), .B(a[49]), .Z(n1098) );
  XNOR U1175 ( .A(b[1]), .B(n1098), .Z(n1100) );
  NANDN U1176 ( .A(b[0]), .B(a[48]), .Z(n1099) );
  NAND U1177 ( .A(n1100), .B(n1099), .Z(n1125) );
  AND U1178 ( .A(b[3]), .B(a[45]), .Z(n1124) );
  XOR U1179 ( .A(n1125), .B(n1124), .Z(n1127) );
  XOR U1180 ( .A(n1126), .B(n1127), .Z(n1113) );
  NANDN U1181 ( .A(n1102), .B(n1101), .Z(n1106) );
  OR U1182 ( .A(n1104), .B(n1103), .Z(n1105) );
  AND U1183 ( .A(n1106), .B(n1105), .Z(n1112) );
  XOR U1184 ( .A(n1113), .B(n1112), .Z(n1115) );
  XOR U1185 ( .A(n1114), .B(n1115), .Z(n1130) );
  XNOR U1186 ( .A(n1130), .B(sreg[301]), .Z(n1132) );
  NANDN U1187 ( .A(n1107), .B(sreg[300]), .Z(n1111) );
  NAND U1188 ( .A(n1109), .B(n1108), .Z(n1110) );
  NAND U1189 ( .A(n1111), .B(n1110), .Z(n1131) );
  XOR U1190 ( .A(n1132), .B(n1131), .Z(c[301]) );
  NANDN U1191 ( .A(n1113), .B(n1112), .Z(n1117) );
  OR U1192 ( .A(n1115), .B(n1114), .Z(n1116) );
  AND U1193 ( .A(n1117), .B(n1116), .Z(n1137) );
  NAND U1194 ( .A(n31), .B(n1118), .Z(n1120) );
  XOR U1195 ( .A(b[3]), .B(a[48]), .Z(n1141) );
  NAND U1196 ( .A(n5811), .B(n1141), .Z(n1119) );
  AND U1197 ( .A(n1120), .B(n1119), .Z(n1149) );
  NAND U1198 ( .A(b[0]), .B(a[50]), .Z(n1121) );
  XNOR U1199 ( .A(b[1]), .B(n1121), .Z(n1123) );
  NANDN U1200 ( .A(b[0]), .B(a[49]), .Z(n1122) );
  NAND U1201 ( .A(n1123), .B(n1122), .Z(n1148) );
  AND U1202 ( .A(b[3]), .B(a[46]), .Z(n1147) );
  XOR U1203 ( .A(n1148), .B(n1147), .Z(n1150) );
  XOR U1204 ( .A(n1149), .B(n1150), .Z(n1136) );
  NANDN U1205 ( .A(n1125), .B(n1124), .Z(n1129) );
  OR U1206 ( .A(n1127), .B(n1126), .Z(n1128) );
  AND U1207 ( .A(n1129), .B(n1128), .Z(n1135) );
  XOR U1208 ( .A(n1136), .B(n1135), .Z(n1138) );
  XOR U1209 ( .A(n1137), .B(n1138), .Z(n1153) );
  XNOR U1210 ( .A(n1153), .B(sreg[302]), .Z(n1155) );
  NANDN U1211 ( .A(n1130), .B(sreg[301]), .Z(n1134) );
  NAND U1212 ( .A(n1132), .B(n1131), .Z(n1133) );
  NAND U1213 ( .A(n1134), .B(n1133), .Z(n1154) );
  XOR U1214 ( .A(n1155), .B(n1154), .Z(c[302]) );
  NANDN U1215 ( .A(n1136), .B(n1135), .Z(n1140) );
  OR U1216 ( .A(n1138), .B(n1137), .Z(n1139) );
  AND U1217 ( .A(n1140), .B(n1139), .Z(n1160) );
  NAND U1218 ( .A(n31), .B(n1141), .Z(n1143) );
  XOR U1219 ( .A(b[3]), .B(a[49]), .Z(n1164) );
  NAND U1220 ( .A(n5811), .B(n1164), .Z(n1142) );
  AND U1221 ( .A(n1143), .B(n1142), .Z(n1172) );
  NAND U1222 ( .A(b[0]), .B(a[51]), .Z(n1144) );
  XNOR U1223 ( .A(b[1]), .B(n1144), .Z(n1146) );
  NANDN U1224 ( .A(b[0]), .B(a[50]), .Z(n1145) );
  NAND U1225 ( .A(n1146), .B(n1145), .Z(n1171) );
  AND U1226 ( .A(b[3]), .B(a[47]), .Z(n1170) );
  XOR U1227 ( .A(n1171), .B(n1170), .Z(n1173) );
  XOR U1228 ( .A(n1172), .B(n1173), .Z(n1159) );
  NANDN U1229 ( .A(n1148), .B(n1147), .Z(n1152) );
  OR U1230 ( .A(n1150), .B(n1149), .Z(n1151) );
  AND U1231 ( .A(n1152), .B(n1151), .Z(n1158) );
  XOR U1232 ( .A(n1159), .B(n1158), .Z(n1161) );
  XOR U1233 ( .A(n1160), .B(n1161), .Z(n1176) );
  XNOR U1234 ( .A(n1176), .B(sreg[303]), .Z(n1178) );
  NANDN U1235 ( .A(n1153), .B(sreg[302]), .Z(n1157) );
  NAND U1236 ( .A(n1155), .B(n1154), .Z(n1156) );
  NAND U1237 ( .A(n1157), .B(n1156), .Z(n1177) );
  XOR U1238 ( .A(n1178), .B(n1177), .Z(c[303]) );
  NANDN U1239 ( .A(n1159), .B(n1158), .Z(n1163) );
  OR U1240 ( .A(n1161), .B(n1160), .Z(n1162) );
  AND U1241 ( .A(n1163), .B(n1162), .Z(n1183) );
  NAND U1242 ( .A(n31), .B(n1164), .Z(n1166) );
  XOR U1243 ( .A(b[3]), .B(a[50]), .Z(n1187) );
  NAND U1244 ( .A(n5811), .B(n1187), .Z(n1165) );
  AND U1245 ( .A(n1166), .B(n1165), .Z(n1195) );
  AND U1246 ( .A(b[3]), .B(a[48]), .Z(n1193) );
  NAND U1247 ( .A(b[0]), .B(a[52]), .Z(n1167) );
  XNOR U1248 ( .A(b[1]), .B(n1167), .Z(n1169) );
  NANDN U1249 ( .A(b[0]), .B(a[51]), .Z(n1168) );
  NAND U1250 ( .A(n1169), .B(n1168), .Z(n1194) );
  XOR U1251 ( .A(n1193), .B(n1194), .Z(n1196) );
  XOR U1252 ( .A(n1195), .B(n1196), .Z(n1182) );
  NANDN U1253 ( .A(n1171), .B(n1170), .Z(n1175) );
  OR U1254 ( .A(n1173), .B(n1172), .Z(n1174) );
  AND U1255 ( .A(n1175), .B(n1174), .Z(n1181) );
  XOR U1256 ( .A(n1182), .B(n1181), .Z(n1184) );
  XOR U1257 ( .A(n1183), .B(n1184), .Z(n1199) );
  XNOR U1258 ( .A(n1199), .B(sreg[304]), .Z(n1201) );
  NANDN U1259 ( .A(n1176), .B(sreg[303]), .Z(n1180) );
  NAND U1260 ( .A(n1178), .B(n1177), .Z(n1179) );
  NAND U1261 ( .A(n1180), .B(n1179), .Z(n1200) );
  XOR U1262 ( .A(n1201), .B(n1200), .Z(c[304]) );
  NANDN U1263 ( .A(n1182), .B(n1181), .Z(n1186) );
  OR U1264 ( .A(n1184), .B(n1183), .Z(n1185) );
  AND U1265 ( .A(n1186), .B(n1185), .Z(n1206) );
  NAND U1266 ( .A(n31), .B(n1187), .Z(n1189) );
  XOR U1267 ( .A(b[3]), .B(a[51]), .Z(n1210) );
  NAND U1268 ( .A(n5811), .B(n1210), .Z(n1188) );
  AND U1269 ( .A(n1189), .B(n1188), .Z(n1218) );
  NAND U1270 ( .A(b[0]), .B(a[53]), .Z(n1190) );
  XNOR U1271 ( .A(b[1]), .B(n1190), .Z(n1192) );
  NANDN U1272 ( .A(b[0]), .B(a[52]), .Z(n1191) );
  NAND U1273 ( .A(n1192), .B(n1191), .Z(n1217) );
  AND U1274 ( .A(b[3]), .B(a[49]), .Z(n1216) );
  XOR U1275 ( .A(n1217), .B(n1216), .Z(n1219) );
  XOR U1276 ( .A(n1218), .B(n1219), .Z(n1205) );
  NANDN U1277 ( .A(n1194), .B(n1193), .Z(n1198) );
  OR U1278 ( .A(n1196), .B(n1195), .Z(n1197) );
  AND U1279 ( .A(n1198), .B(n1197), .Z(n1204) );
  XOR U1280 ( .A(n1205), .B(n1204), .Z(n1207) );
  XOR U1281 ( .A(n1206), .B(n1207), .Z(n1222) );
  XNOR U1282 ( .A(n1222), .B(sreg[305]), .Z(n1224) );
  NANDN U1283 ( .A(n1199), .B(sreg[304]), .Z(n1203) );
  NAND U1284 ( .A(n1201), .B(n1200), .Z(n1202) );
  NAND U1285 ( .A(n1203), .B(n1202), .Z(n1223) );
  XOR U1286 ( .A(n1224), .B(n1223), .Z(c[305]) );
  NANDN U1287 ( .A(n1205), .B(n1204), .Z(n1209) );
  OR U1288 ( .A(n1207), .B(n1206), .Z(n1208) );
  AND U1289 ( .A(n1209), .B(n1208), .Z(n1229) );
  NAND U1290 ( .A(n31), .B(n1210), .Z(n1212) );
  XOR U1291 ( .A(b[3]), .B(a[52]), .Z(n1233) );
  NAND U1292 ( .A(n5811), .B(n1233), .Z(n1211) );
  AND U1293 ( .A(n1212), .B(n1211), .Z(n1241) );
  NAND U1294 ( .A(b[0]), .B(a[54]), .Z(n1213) );
  XNOR U1295 ( .A(b[1]), .B(n1213), .Z(n1215) );
  NANDN U1296 ( .A(b[0]), .B(a[53]), .Z(n1214) );
  NAND U1297 ( .A(n1215), .B(n1214), .Z(n1240) );
  AND U1298 ( .A(b[3]), .B(a[50]), .Z(n1239) );
  XOR U1299 ( .A(n1240), .B(n1239), .Z(n1242) );
  XOR U1300 ( .A(n1241), .B(n1242), .Z(n1228) );
  NANDN U1301 ( .A(n1217), .B(n1216), .Z(n1221) );
  OR U1302 ( .A(n1219), .B(n1218), .Z(n1220) );
  AND U1303 ( .A(n1221), .B(n1220), .Z(n1227) );
  XOR U1304 ( .A(n1228), .B(n1227), .Z(n1230) );
  XOR U1305 ( .A(n1229), .B(n1230), .Z(n1245) );
  XNOR U1306 ( .A(n1245), .B(sreg[306]), .Z(n1247) );
  NANDN U1307 ( .A(n1222), .B(sreg[305]), .Z(n1226) );
  NAND U1308 ( .A(n1224), .B(n1223), .Z(n1225) );
  NAND U1309 ( .A(n1226), .B(n1225), .Z(n1246) );
  XOR U1310 ( .A(n1247), .B(n1246), .Z(c[306]) );
  NANDN U1311 ( .A(n1228), .B(n1227), .Z(n1232) );
  OR U1312 ( .A(n1230), .B(n1229), .Z(n1231) );
  AND U1313 ( .A(n1232), .B(n1231), .Z(n1252) );
  NAND U1314 ( .A(n31), .B(n1233), .Z(n1235) );
  XOR U1315 ( .A(b[3]), .B(a[53]), .Z(n1256) );
  NAND U1316 ( .A(n5811), .B(n1256), .Z(n1234) );
  AND U1317 ( .A(n1235), .B(n1234), .Z(n1264) );
  NAND U1318 ( .A(b[0]), .B(a[55]), .Z(n1236) );
  XNOR U1319 ( .A(b[1]), .B(n1236), .Z(n1238) );
  NANDN U1320 ( .A(b[0]), .B(a[54]), .Z(n1237) );
  NAND U1321 ( .A(n1238), .B(n1237), .Z(n1263) );
  AND U1322 ( .A(b[3]), .B(a[51]), .Z(n1262) );
  XOR U1323 ( .A(n1263), .B(n1262), .Z(n1265) );
  XOR U1324 ( .A(n1264), .B(n1265), .Z(n1251) );
  NANDN U1325 ( .A(n1240), .B(n1239), .Z(n1244) );
  OR U1326 ( .A(n1242), .B(n1241), .Z(n1243) );
  AND U1327 ( .A(n1244), .B(n1243), .Z(n1250) );
  XOR U1328 ( .A(n1251), .B(n1250), .Z(n1253) );
  XOR U1329 ( .A(n1252), .B(n1253), .Z(n1268) );
  XNOR U1330 ( .A(n1268), .B(sreg[307]), .Z(n1270) );
  NANDN U1331 ( .A(n1245), .B(sreg[306]), .Z(n1249) );
  NAND U1332 ( .A(n1247), .B(n1246), .Z(n1248) );
  NAND U1333 ( .A(n1249), .B(n1248), .Z(n1269) );
  XOR U1334 ( .A(n1270), .B(n1269), .Z(c[307]) );
  NANDN U1335 ( .A(n1251), .B(n1250), .Z(n1255) );
  OR U1336 ( .A(n1253), .B(n1252), .Z(n1254) );
  AND U1337 ( .A(n1255), .B(n1254), .Z(n1275) );
  NAND U1338 ( .A(n31), .B(n1256), .Z(n1258) );
  XOR U1339 ( .A(b[3]), .B(a[54]), .Z(n1279) );
  NAND U1340 ( .A(n5811), .B(n1279), .Z(n1257) );
  AND U1341 ( .A(n1258), .B(n1257), .Z(n1287) );
  AND U1342 ( .A(b[3]), .B(a[52]), .Z(n1285) );
  NAND U1343 ( .A(b[0]), .B(a[56]), .Z(n1259) );
  XNOR U1344 ( .A(b[1]), .B(n1259), .Z(n1261) );
  NANDN U1345 ( .A(b[0]), .B(a[55]), .Z(n1260) );
  NAND U1346 ( .A(n1261), .B(n1260), .Z(n1286) );
  XOR U1347 ( .A(n1285), .B(n1286), .Z(n1288) );
  XOR U1348 ( .A(n1287), .B(n1288), .Z(n1274) );
  NANDN U1349 ( .A(n1263), .B(n1262), .Z(n1267) );
  OR U1350 ( .A(n1265), .B(n1264), .Z(n1266) );
  AND U1351 ( .A(n1267), .B(n1266), .Z(n1273) );
  XOR U1352 ( .A(n1274), .B(n1273), .Z(n1276) );
  XOR U1353 ( .A(n1275), .B(n1276), .Z(n1291) );
  XNOR U1354 ( .A(n1291), .B(sreg[308]), .Z(n1293) );
  NANDN U1355 ( .A(n1268), .B(sreg[307]), .Z(n1272) );
  NAND U1356 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U1357 ( .A(n1272), .B(n1271), .Z(n1292) );
  XOR U1358 ( .A(n1293), .B(n1292), .Z(c[308]) );
  NANDN U1359 ( .A(n1274), .B(n1273), .Z(n1278) );
  OR U1360 ( .A(n1276), .B(n1275), .Z(n1277) );
  AND U1361 ( .A(n1278), .B(n1277), .Z(n1298) );
  NAND U1362 ( .A(n31), .B(n1279), .Z(n1281) );
  XOR U1363 ( .A(b[3]), .B(a[55]), .Z(n1302) );
  NAND U1364 ( .A(n5811), .B(n1302), .Z(n1280) );
  AND U1365 ( .A(n1281), .B(n1280), .Z(n1310) );
  NAND U1366 ( .A(b[0]), .B(a[57]), .Z(n1282) );
  XNOR U1367 ( .A(b[1]), .B(n1282), .Z(n1284) );
  NANDN U1368 ( .A(b[0]), .B(a[56]), .Z(n1283) );
  NAND U1369 ( .A(n1284), .B(n1283), .Z(n1309) );
  AND U1370 ( .A(b[3]), .B(a[53]), .Z(n1308) );
  XOR U1371 ( .A(n1309), .B(n1308), .Z(n1311) );
  XOR U1372 ( .A(n1310), .B(n1311), .Z(n1297) );
  NANDN U1373 ( .A(n1286), .B(n1285), .Z(n1290) );
  OR U1374 ( .A(n1288), .B(n1287), .Z(n1289) );
  AND U1375 ( .A(n1290), .B(n1289), .Z(n1296) );
  XOR U1376 ( .A(n1297), .B(n1296), .Z(n1299) );
  XOR U1377 ( .A(n1298), .B(n1299), .Z(n1314) );
  XNOR U1378 ( .A(n1314), .B(sreg[309]), .Z(n1316) );
  NANDN U1379 ( .A(n1291), .B(sreg[308]), .Z(n1295) );
  NAND U1380 ( .A(n1293), .B(n1292), .Z(n1294) );
  NAND U1381 ( .A(n1295), .B(n1294), .Z(n1315) );
  XOR U1382 ( .A(n1316), .B(n1315), .Z(c[309]) );
  NANDN U1383 ( .A(n1297), .B(n1296), .Z(n1301) );
  OR U1384 ( .A(n1299), .B(n1298), .Z(n1300) );
  AND U1385 ( .A(n1301), .B(n1300), .Z(n1321) );
  NAND U1386 ( .A(n31), .B(n1302), .Z(n1304) );
  XOR U1387 ( .A(b[3]), .B(a[56]), .Z(n1325) );
  NAND U1388 ( .A(n5811), .B(n1325), .Z(n1303) );
  AND U1389 ( .A(n1304), .B(n1303), .Z(n1333) );
  NAND U1390 ( .A(b[0]), .B(a[58]), .Z(n1305) );
  XNOR U1391 ( .A(b[1]), .B(n1305), .Z(n1307) );
  NANDN U1392 ( .A(b[0]), .B(a[57]), .Z(n1306) );
  NAND U1393 ( .A(n1307), .B(n1306), .Z(n1332) );
  AND U1394 ( .A(b[3]), .B(a[54]), .Z(n1331) );
  XOR U1395 ( .A(n1332), .B(n1331), .Z(n1334) );
  XOR U1396 ( .A(n1333), .B(n1334), .Z(n1320) );
  NANDN U1397 ( .A(n1309), .B(n1308), .Z(n1313) );
  OR U1398 ( .A(n1311), .B(n1310), .Z(n1312) );
  AND U1399 ( .A(n1313), .B(n1312), .Z(n1319) );
  XOR U1400 ( .A(n1320), .B(n1319), .Z(n1322) );
  XOR U1401 ( .A(n1321), .B(n1322), .Z(n1337) );
  XNOR U1402 ( .A(n1337), .B(sreg[310]), .Z(n1339) );
  NANDN U1403 ( .A(n1314), .B(sreg[309]), .Z(n1318) );
  NAND U1404 ( .A(n1316), .B(n1315), .Z(n1317) );
  NAND U1405 ( .A(n1318), .B(n1317), .Z(n1338) );
  XOR U1406 ( .A(n1339), .B(n1338), .Z(c[310]) );
  NANDN U1407 ( .A(n1320), .B(n1319), .Z(n1324) );
  OR U1408 ( .A(n1322), .B(n1321), .Z(n1323) );
  AND U1409 ( .A(n1324), .B(n1323), .Z(n1344) );
  NAND U1410 ( .A(n31), .B(n1325), .Z(n1327) );
  XOR U1411 ( .A(b[3]), .B(a[57]), .Z(n1348) );
  NAND U1412 ( .A(n5811), .B(n1348), .Z(n1326) );
  AND U1413 ( .A(n1327), .B(n1326), .Z(n1356) );
  NAND U1414 ( .A(b[0]), .B(a[59]), .Z(n1328) );
  XNOR U1415 ( .A(b[1]), .B(n1328), .Z(n1330) );
  NANDN U1416 ( .A(b[0]), .B(a[58]), .Z(n1329) );
  NAND U1417 ( .A(n1330), .B(n1329), .Z(n1355) );
  AND U1418 ( .A(b[3]), .B(a[55]), .Z(n1354) );
  XOR U1419 ( .A(n1355), .B(n1354), .Z(n1357) );
  XOR U1420 ( .A(n1356), .B(n1357), .Z(n1343) );
  NANDN U1421 ( .A(n1332), .B(n1331), .Z(n1336) );
  OR U1422 ( .A(n1334), .B(n1333), .Z(n1335) );
  AND U1423 ( .A(n1336), .B(n1335), .Z(n1342) );
  XOR U1424 ( .A(n1343), .B(n1342), .Z(n1345) );
  XOR U1425 ( .A(n1344), .B(n1345), .Z(n1360) );
  XNOR U1426 ( .A(n1360), .B(sreg[311]), .Z(n1362) );
  NANDN U1427 ( .A(n1337), .B(sreg[310]), .Z(n1341) );
  NAND U1428 ( .A(n1339), .B(n1338), .Z(n1340) );
  NAND U1429 ( .A(n1341), .B(n1340), .Z(n1361) );
  XOR U1430 ( .A(n1362), .B(n1361), .Z(c[311]) );
  NANDN U1431 ( .A(n1343), .B(n1342), .Z(n1347) );
  OR U1432 ( .A(n1345), .B(n1344), .Z(n1346) );
  AND U1433 ( .A(n1347), .B(n1346), .Z(n1367) );
  NAND U1434 ( .A(n31), .B(n1348), .Z(n1350) );
  XOR U1435 ( .A(b[3]), .B(a[58]), .Z(n1371) );
  NAND U1436 ( .A(n5811), .B(n1371), .Z(n1349) );
  AND U1437 ( .A(n1350), .B(n1349), .Z(n1379) );
  NAND U1438 ( .A(b[0]), .B(a[60]), .Z(n1351) );
  XNOR U1439 ( .A(b[1]), .B(n1351), .Z(n1353) );
  NANDN U1440 ( .A(b[0]), .B(a[59]), .Z(n1352) );
  NAND U1441 ( .A(n1353), .B(n1352), .Z(n1378) );
  AND U1442 ( .A(b[3]), .B(a[56]), .Z(n1377) );
  XOR U1443 ( .A(n1378), .B(n1377), .Z(n1380) );
  XOR U1444 ( .A(n1379), .B(n1380), .Z(n1366) );
  NANDN U1445 ( .A(n1355), .B(n1354), .Z(n1359) );
  OR U1446 ( .A(n1357), .B(n1356), .Z(n1358) );
  AND U1447 ( .A(n1359), .B(n1358), .Z(n1365) );
  XOR U1448 ( .A(n1366), .B(n1365), .Z(n1368) );
  XOR U1449 ( .A(n1367), .B(n1368), .Z(n1383) );
  XNOR U1450 ( .A(n1383), .B(sreg[312]), .Z(n1385) );
  NANDN U1451 ( .A(n1360), .B(sreg[311]), .Z(n1364) );
  NAND U1452 ( .A(n1362), .B(n1361), .Z(n1363) );
  NAND U1453 ( .A(n1364), .B(n1363), .Z(n1384) );
  XOR U1454 ( .A(n1385), .B(n1384), .Z(c[312]) );
  NANDN U1455 ( .A(n1366), .B(n1365), .Z(n1370) );
  OR U1456 ( .A(n1368), .B(n1367), .Z(n1369) );
  AND U1457 ( .A(n1370), .B(n1369), .Z(n1390) );
  NAND U1458 ( .A(n31), .B(n1371), .Z(n1373) );
  XOR U1459 ( .A(b[3]), .B(a[59]), .Z(n1394) );
  NAND U1460 ( .A(n5811), .B(n1394), .Z(n1372) );
  AND U1461 ( .A(n1373), .B(n1372), .Z(n1402) );
  NAND U1462 ( .A(b[0]), .B(a[61]), .Z(n1374) );
  XNOR U1463 ( .A(b[1]), .B(n1374), .Z(n1376) );
  NANDN U1464 ( .A(b[0]), .B(a[60]), .Z(n1375) );
  NAND U1465 ( .A(n1376), .B(n1375), .Z(n1401) );
  AND U1466 ( .A(b[3]), .B(a[57]), .Z(n1400) );
  XOR U1467 ( .A(n1401), .B(n1400), .Z(n1403) );
  XOR U1468 ( .A(n1402), .B(n1403), .Z(n1389) );
  NANDN U1469 ( .A(n1378), .B(n1377), .Z(n1382) );
  OR U1470 ( .A(n1380), .B(n1379), .Z(n1381) );
  AND U1471 ( .A(n1382), .B(n1381), .Z(n1388) );
  XOR U1472 ( .A(n1389), .B(n1388), .Z(n1391) );
  XOR U1473 ( .A(n1390), .B(n1391), .Z(n1406) );
  XNOR U1474 ( .A(n1406), .B(sreg[313]), .Z(n1408) );
  NANDN U1475 ( .A(n1383), .B(sreg[312]), .Z(n1387) );
  NAND U1476 ( .A(n1385), .B(n1384), .Z(n1386) );
  NAND U1477 ( .A(n1387), .B(n1386), .Z(n1407) );
  XOR U1478 ( .A(n1408), .B(n1407), .Z(c[313]) );
  NANDN U1479 ( .A(n1389), .B(n1388), .Z(n1393) );
  OR U1480 ( .A(n1391), .B(n1390), .Z(n1392) );
  AND U1481 ( .A(n1393), .B(n1392), .Z(n1413) );
  NAND U1482 ( .A(n31), .B(n1394), .Z(n1396) );
  XOR U1483 ( .A(b[3]), .B(a[60]), .Z(n1417) );
  NAND U1484 ( .A(n5811), .B(n1417), .Z(n1395) );
  AND U1485 ( .A(n1396), .B(n1395), .Z(n1425) );
  AND U1486 ( .A(b[3]), .B(a[58]), .Z(n1423) );
  NAND U1487 ( .A(b[0]), .B(a[62]), .Z(n1397) );
  XNOR U1488 ( .A(b[1]), .B(n1397), .Z(n1399) );
  NANDN U1489 ( .A(b[0]), .B(a[61]), .Z(n1398) );
  NAND U1490 ( .A(n1399), .B(n1398), .Z(n1424) );
  XOR U1491 ( .A(n1423), .B(n1424), .Z(n1426) );
  XOR U1492 ( .A(n1425), .B(n1426), .Z(n1412) );
  NANDN U1493 ( .A(n1401), .B(n1400), .Z(n1405) );
  OR U1494 ( .A(n1403), .B(n1402), .Z(n1404) );
  AND U1495 ( .A(n1405), .B(n1404), .Z(n1411) );
  XOR U1496 ( .A(n1412), .B(n1411), .Z(n1414) );
  XOR U1497 ( .A(n1413), .B(n1414), .Z(n1429) );
  XNOR U1498 ( .A(n1429), .B(sreg[314]), .Z(n1431) );
  NANDN U1499 ( .A(n1406), .B(sreg[313]), .Z(n1410) );
  NAND U1500 ( .A(n1408), .B(n1407), .Z(n1409) );
  NAND U1501 ( .A(n1410), .B(n1409), .Z(n1430) );
  XOR U1502 ( .A(n1431), .B(n1430), .Z(c[314]) );
  NANDN U1503 ( .A(n1412), .B(n1411), .Z(n1416) );
  OR U1504 ( .A(n1414), .B(n1413), .Z(n1415) );
  AND U1505 ( .A(n1416), .B(n1415), .Z(n1436) );
  NAND U1506 ( .A(n31), .B(n1417), .Z(n1419) );
  XOR U1507 ( .A(b[3]), .B(a[61]), .Z(n1440) );
  NAND U1508 ( .A(n5811), .B(n1440), .Z(n1418) );
  AND U1509 ( .A(n1419), .B(n1418), .Z(n1448) );
  NAND U1510 ( .A(b[0]), .B(a[63]), .Z(n1420) );
  XNOR U1511 ( .A(b[1]), .B(n1420), .Z(n1422) );
  NANDN U1512 ( .A(b[0]), .B(a[62]), .Z(n1421) );
  NAND U1513 ( .A(n1422), .B(n1421), .Z(n1447) );
  AND U1514 ( .A(b[3]), .B(a[59]), .Z(n1446) );
  XOR U1515 ( .A(n1447), .B(n1446), .Z(n1449) );
  XOR U1516 ( .A(n1448), .B(n1449), .Z(n1435) );
  NANDN U1517 ( .A(n1424), .B(n1423), .Z(n1428) );
  OR U1518 ( .A(n1426), .B(n1425), .Z(n1427) );
  AND U1519 ( .A(n1428), .B(n1427), .Z(n1434) );
  XOR U1520 ( .A(n1435), .B(n1434), .Z(n1437) );
  XOR U1521 ( .A(n1436), .B(n1437), .Z(n1452) );
  XNOR U1522 ( .A(n1452), .B(sreg[315]), .Z(n1454) );
  NANDN U1523 ( .A(n1429), .B(sreg[314]), .Z(n1433) );
  NAND U1524 ( .A(n1431), .B(n1430), .Z(n1432) );
  NAND U1525 ( .A(n1433), .B(n1432), .Z(n1453) );
  XOR U1526 ( .A(n1454), .B(n1453), .Z(c[315]) );
  NANDN U1527 ( .A(n1435), .B(n1434), .Z(n1439) );
  OR U1528 ( .A(n1437), .B(n1436), .Z(n1438) );
  AND U1529 ( .A(n1439), .B(n1438), .Z(n1459) );
  NAND U1530 ( .A(n31), .B(n1440), .Z(n1442) );
  XOR U1531 ( .A(b[3]), .B(a[62]), .Z(n1463) );
  NAND U1532 ( .A(n5811), .B(n1463), .Z(n1441) );
  AND U1533 ( .A(n1442), .B(n1441), .Z(n1471) );
  AND U1534 ( .A(b[3]), .B(a[60]), .Z(n1469) );
  NAND U1535 ( .A(b[0]), .B(a[64]), .Z(n1443) );
  XNOR U1536 ( .A(b[1]), .B(n1443), .Z(n1445) );
  NANDN U1537 ( .A(b[0]), .B(a[63]), .Z(n1444) );
  NAND U1538 ( .A(n1445), .B(n1444), .Z(n1470) );
  XOR U1539 ( .A(n1469), .B(n1470), .Z(n1472) );
  XOR U1540 ( .A(n1471), .B(n1472), .Z(n1458) );
  NANDN U1541 ( .A(n1447), .B(n1446), .Z(n1451) );
  OR U1542 ( .A(n1449), .B(n1448), .Z(n1450) );
  AND U1543 ( .A(n1451), .B(n1450), .Z(n1457) );
  XOR U1544 ( .A(n1458), .B(n1457), .Z(n1460) );
  XOR U1545 ( .A(n1459), .B(n1460), .Z(n1475) );
  XNOR U1546 ( .A(n1475), .B(sreg[316]), .Z(n1477) );
  NANDN U1547 ( .A(n1452), .B(sreg[315]), .Z(n1456) );
  NAND U1548 ( .A(n1454), .B(n1453), .Z(n1455) );
  NAND U1549 ( .A(n1456), .B(n1455), .Z(n1476) );
  XOR U1550 ( .A(n1477), .B(n1476), .Z(c[316]) );
  NANDN U1551 ( .A(n1458), .B(n1457), .Z(n1462) );
  OR U1552 ( .A(n1460), .B(n1459), .Z(n1461) );
  AND U1553 ( .A(n1462), .B(n1461), .Z(n1482) );
  NAND U1554 ( .A(n31), .B(n1463), .Z(n1465) );
  XOR U1555 ( .A(b[3]), .B(a[63]), .Z(n1486) );
  NAND U1556 ( .A(n5811), .B(n1486), .Z(n1464) );
  AND U1557 ( .A(n1465), .B(n1464), .Z(n1494) );
  NAND U1558 ( .A(b[0]), .B(a[65]), .Z(n1466) );
  XNOR U1559 ( .A(b[1]), .B(n1466), .Z(n1468) );
  NANDN U1560 ( .A(b[0]), .B(a[64]), .Z(n1467) );
  NAND U1561 ( .A(n1468), .B(n1467), .Z(n1493) );
  AND U1562 ( .A(b[3]), .B(a[61]), .Z(n1492) );
  XOR U1563 ( .A(n1493), .B(n1492), .Z(n1495) );
  XOR U1564 ( .A(n1494), .B(n1495), .Z(n1481) );
  NANDN U1565 ( .A(n1470), .B(n1469), .Z(n1474) );
  OR U1566 ( .A(n1472), .B(n1471), .Z(n1473) );
  AND U1567 ( .A(n1474), .B(n1473), .Z(n1480) );
  XOR U1568 ( .A(n1481), .B(n1480), .Z(n1483) );
  XOR U1569 ( .A(n1482), .B(n1483), .Z(n1498) );
  XNOR U1570 ( .A(n1498), .B(sreg[317]), .Z(n1500) );
  NANDN U1571 ( .A(n1475), .B(sreg[316]), .Z(n1479) );
  NAND U1572 ( .A(n1477), .B(n1476), .Z(n1478) );
  NAND U1573 ( .A(n1479), .B(n1478), .Z(n1499) );
  XOR U1574 ( .A(n1500), .B(n1499), .Z(c[317]) );
  NANDN U1575 ( .A(n1481), .B(n1480), .Z(n1485) );
  OR U1576 ( .A(n1483), .B(n1482), .Z(n1484) );
  AND U1577 ( .A(n1485), .B(n1484), .Z(n1505) );
  NAND U1578 ( .A(n31), .B(n1486), .Z(n1488) );
  XOR U1579 ( .A(b[3]), .B(a[64]), .Z(n1509) );
  NAND U1580 ( .A(n5811), .B(n1509), .Z(n1487) );
  AND U1581 ( .A(n1488), .B(n1487), .Z(n1517) );
  NAND U1582 ( .A(b[0]), .B(a[66]), .Z(n1489) );
  XNOR U1583 ( .A(b[1]), .B(n1489), .Z(n1491) );
  NANDN U1584 ( .A(b[0]), .B(a[65]), .Z(n1490) );
  NAND U1585 ( .A(n1491), .B(n1490), .Z(n1516) );
  AND U1586 ( .A(b[3]), .B(a[62]), .Z(n1515) );
  XOR U1587 ( .A(n1516), .B(n1515), .Z(n1518) );
  XOR U1588 ( .A(n1517), .B(n1518), .Z(n1504) );
  NANDN U1589 ( .A(n1493), .B(n1492), .Z(n1497) );
  OR U1590 ( .A(n1495), .B(n1494), .Z(n1496) );
  AND U1591 ( .A(n1497), .B(n1496), .Z(n1503) );
  XOR U1592 ( .A(n1504), .B(n1503), .Z(n1506) );
  XOR U1593 ( .A(n1505), .B(n1506), .Z(n1521) );
  XNOR U1594 ( .A(n1521), .B(sreg[318]), .Z(n1523) );
  NANDN U1595 ( .A(n1498), .B(sreg[317]), .Z(n1502) );
  NAND U1596 ( .A(n1500), .B(n1499), .Z(n1501) );
  NAND U1597 ( .A(n1502), .B(n1501), .Z(n1522) );
  XOR U1598 ( .A(n1523), .B(n1522), .Z(c[318]) );
  NANDN U1599 ( .A(n1504), .B(n1503), .Z(n1508) );
  OR U1600 ( .A(n1506), .B(n1505), .Z(n1507) );
  AND U1601 ( .A(n1508), .B(n1507), .Z(n1528) );
  NAND U1602 ( .A(n31), .B(n1509), .Z(n1511) );
  XOR U1603 ( .A(b[3]), .B(a[65]), .Z(n1532) );
  NAND U1604 ( .A(n5811), .B(n1532), .Z(n1510) );
  AND U1605 ( .A(n1511), .B(n1510), .Z(n1540) );
  AND U1606 ( .A(b[3]), .B(a[63]), .Z(n1538) );
  NAND U1607 ( .A(b[0]), .B(a[67]), .Z(n1512) );
  XNOR U1608 ( .A(b[1]), .B(n1512), .Z(n1514) );
  NANDN U1609 ( .A(b[0]), .B(a[66]), .Z(n1513) );
  NAND U1610 ( .A(n1514), .B(n1513), .Z(n1539) );
  XOR U1611 ( .A(n1538), .B(n1539), .Z(n1541) );
  XOR U1612 ( .A(n1540), .B(n1541), .Z(n1527) );
  NANDN U1613 ( .A(n1516), .B(n1515), .Z(n1520) );
  OR U1614 ( .A(n1518), .B(n1517), .Z(n1519) );
  AND U1615 ( .A(n1520), .B(n1519), .Z(n1526) );
  XOR U1616 ( .A(n1527), .B(n1526), .Z(n1529) );
  XOR U1617 ( .A(n1528), .B(n1529), .Z(n1544) );
  XNOR U1618 ( .A(n1544), .B(sreg[319]), .Z(n1546) );
  NANDN U1619 ( .A(n1521), .B(sreg[318]), .Z(n1525) );
  NAND U1620 ( .A(n1523), .B(n1522), .Z(n1524) );
  NAND U1621 ( .A(n1525), .B(n1524), .Z(n1545) );
  XOR U1622 ( .A(n1546), .B(n1545), .Z(c[319]) );
  NANDN U1623 ( .A(n1527), .B(n1526), .Z(n1531) );
  OR U1624 ( .A(n1529), .B(n1528), .Z(n1530) );
  AND U1625 ( .A(n1531), .B(n1530), .Z(n1551) );
  NAND U1626 ( .A(n31), .B(n1532), .Z(n1534) );
  XOR U1627 ( .A(b[3]), .B(a[66]), .Z(n1555) );
  NAND U1628 ( .A(n5811), .B(n1555), .Z(n1533) );
  AND U1629 ( .A(n1534), .B(n1533), .Z(n1563) );
  NAND U1630 ( .A(b[0]), .B(a[68]), .Z(n1535) );
  XNOR U1631 ( .A(b[1]), .B(n1535), .Z(n1537) );
  NANDN U1632 ( .A(b[0]), .B(a[67]), .Z(n1536) );
  NAND U1633 ( .A(n1537), .B(n1536), .Z(n1562) );
  AND U1634 ( .A(b[3]), .B(a[64]), .Z(n1561) );
  XOR U1635 ( .A(n1562), .B(n1561), .Z(n1564) );
  XOR U1636 ( .A(n1563), .B(n1564), .Z(n1550) );
  NANDN U1637 ( .A(n1539), .B(n1538), .Z(n1543) );
  OR U1638 ( .A(n1541), .B(n1540), .Z(n1542) );
  AND U1639 ( .A(n1543), .B(n1542), .Z(n1549) );
  XOR U1640 ( .A(n1550), .B(n1549), .Z(n1552) );
  XOR U1641 ( .A(n1551), .B(n1552), .Z(n1567) );
  XNOR U1642 ( .A(n1567), .B(sreg[320]), .Z(n1569) );
  NANDN U1643 ( .A(n1544), .B(sreg[319]), .Z(n1548) );
  NAND U1644 ( .A(n1546), .B(n1545), .Z(n1547) );
  NAND U1645 ( .A(n1548), .B(n1547), .Z(n1568) );
  XOR U1646 ( .A(n1569), .B(n1568), .Z(c[320]) );
  NANDN U1647 ( .A(n1550), .B(n1549), .Z(n1554) );
  OR U1648 ( .A(n1552), .B(n1551), .Z(n1553) );
  AND U1649 ( .A(n1554), .B(n1553), .Z(n1574) );
  NAND U1650 ( .A(n31), .B(n1555), .Z(n1557) );
  XOR U1651 ( .A(b[3]), .B(a[67]), .Z(n1578) );
  NAND U1652 ( .A(n5811), .B(n1578), .Z(n1556) );
  AND U1653 ( .A(n1557), .B(n1556), .Z(n1586) );
  NAND U1654 ( .A(b[0]), .B(a[69]), .Z(n1558) );
  XNOR U1655 ( .A(b[1]), .B(n1558), .Z(n1560) );
  NANDN U1656 ( .A(b[0]), .B(a[68]), .Z(n1559) );
  NAND U1657 ( .A(n1560), .B(n1559), .Z(n1585) );
  AND U1658 ( .A(b[3]), .B(a[65]), .Z(n1584) );
  XOR U1659 ( .A(n1585), .B(n1584), .Z(n1587) );
  XOR U1660 ( .A(n1586), .B(n1587), .Z(n1573) );
  NANDN U1661 ( .A(n1562), .B(n1561), .Z(n1566) );
  OR U1662 ( .A(n1564), .B(n1563), .Z(n1565) );
  AND U1663 ( .A(n1566), .B(n1565), .Z(n1572) );
  XOR U1664 ( .A(n1573), .B(n1572), .Z(n1575) );
  XOR U1665 ( .A(n1574), .B(n1575), .Z(n1590) );
  XNOR U1666 ( .A(n1590), .B(sreg[321]), .Z(n1592) );
  NANDN U1667 ( .A(n1567), .B(sreg[320]), .Z(n1571) );
  NAND U1668 ( .A(n1569), .B(n1568), .Z(n1570) );
  NAND U1669 ( .A(n1571), .B(n1570), .Z(n1591) );
  XOR U1670 ( .A(n1592), .B(n1591), .Z(c[321]) );
  NANDN U1671 ( .A(n1573), .B(n1572), .Z(n1577) );
  OR U1672 ( .A(n1575), .B(n1574), .Z(n1576) );
  AND U1673 ( .A(n1577), .B(n1576), .Z(n1597) );
  NAND U1674 ( .A(n31), .B(n1578), .Z(n1580) );
  XOR U1675 ( .A(b[3]), .B(a[68]), .Z(n1601) );
  NAND U1676 ( .A(n5811), .B(n1601), .Z(n1579) );
  AND U1677 ( .A(n1580), .B(n1579), .Z(n1609) );
  NAND U1678 ( .A(b[0]), .B(a[70]), .Z(n1581) );
  XNOR U1679 ( .A(b[1]), .B(n1581), .Z(n1583) );
  NANDN U1680 ( .A(b[0]), .B(a[69]), .Z(n1582) );
  NAND U1681 ( .A(n1583), .B(n1582), .Z(n1608) );
  AND U1682 ( .A(b[3]), .B(a[66]), .Z(n1607) );
  XOR U1683 ( .A(n1608), .B(n1607), .Z(n1610) );
  XOR U1684 ( .A(n1609), .B(n1610), .Z(n1596) );
  NANDN U1685 ( .A(n1585), .B(n1584), .Z(n1589) );
  OR U1686 ( .A(n1587), .B(n1586), .Z(n1588) );
  AND U1687 ( .A(n1589), .B(n1588), .Z(n1595) );
  XOR U1688 ( .A(n1596), .B(n1595), .Z(n1598) );
  XOR U1689 ( .A(n1597), .B(n1598), .Z(n1613) );
  XNOR U1690 ( .A(n1613), .B(sreg[322]), .Z(n1615) );
  NANDN U1691 ( .A(n1590), .B(sreg[321]), .Z(n1594) );
  NAND U1692 ( .A(n1592), .B(n1591), .Z(n1593) );
  NAND U1693 ( .A(n1594), .B(n1593), .Z(n1614) );
  XOR U1694 ( .A(n1615), .B(n1614), .Z(c[322]) );
  NANDN U1695 ( .A(n1596), .B(n1595), .Z(n1600) );
  OR U1696 ( .A(n1598), .B(n1597), .Z(n1599) );
  AND U1697 ( .A(n1600), .B(n1599), .Z(n1620) );
  NAND U1698 ( .A(n31), .B(n1601), .Z(n1603) );
  XOR U1699 ( .A(b[3]), .B(a[69]), .Z(n1624) );
  NAND U1700 ( .A(n5811), .B(n1624), .Z(n1602) );
  AND U1701 ( .A(n1603), .B(n1602), .Z(n1632) );
  AND U1702 ( .A(b[3]), .B(a[67]), .Z(n1630) );
  NAND U1703 ( .A(b[0]), .B(a[71]), .Z(n1604) );
  XNOR U1704 ( .A(b[1]), .B(n1604), .Z(n1606) );
  NANDN U1705 ( .A(b[0]), .B(a[70]), .Z(n1605) );
  NAND U1706 ( .A(n1606), .B(n1605), .Z(n1631) );
  XOR U1707 ( .A(n1630), .B(n1631), .Z(n1633) );
  XOR U1708 ( .A(n1632), .B(n1633), .Z(n1619) );
  NANDN U1709 ( .A(n1608), .B(n1607), .Z(n1612) );
  OR U1710 ( .A(n1610), .B(n1609), .Z(n1611) );
  AND U1711 ( .A(n1612), .B(n1611), .Z(n1618) );
  XOR U1712 ( .A(n1619), .B(n1618), .Z(n1621) );
  XOR U1713 ( .A(n1620), .B(n1621), .Z(n1636) );
  XNOR U1714 ( .A(n1636), .B(sreg[323]), .Z(n1638) );
  NANDN U1715 ( .A(n1613), .B(sreg[322]), .Z(n1617) );
  NAND U1716 ( .A(n1615), .B(n1614), .Z(n1616) );
  NAND U1717 ( .A(n1617), .B(n1616), .Z(n1637) );
  XOR U1718 ( .A(n1638), .B(n1637), .Z(c[323]) );
  NANDN U1719 ( .A(n1619), .B(n1618), .Z(n1623) );
  OR U1720 ( .A(n1621), .B(n1620), .Z(n1622) );
  AND U1721 ( .A(n1623), .B(n1622), .Z(n1643) );
  NAND U1722 ( .A(n31), .B(n1624), .Z(n1626) );
  XOR U1723 ( .A(b[3]), .B(a[70]), .Z(n1647) );
  NAND U1724 ( .A(n5811), .B(n1647), .Z(n1625) );
  AND U1725 ( .A(n1626), .B(n1625), .Z(n1655) );
  NAND U1726 ( .A(b[0]), .B(a[72]), .Z(n1627) );
  XNOR U1727 ( .A(b[1]), .B(n1627), .Z(n1629) );
  NANDN U1728 ( .A(b[0]), .B(a[71]), .Z(n1628) );
  NAND U1729 ( .A(n1629), .B(n1628), .Z(n1654) );
  AND U1730 ( .A(b[3]), .B(a[68]), .Z(n1653) );
  XOR U1731 ( .A(n1654), .B(n1653), .Z(n1656) );
  XOR U1732 ( .A(n1655), .B(n1656), .Z(n1642) );
  NANDN U1733 ( .A(n1631), .B(n1630), .Z(n1635) );
  OR U1734 ( .A(n1633), .B(n1632), .Z(n1634) );
  AND U1735 ( .A(n1635), .B(n1634), .Z(n1641) );
  XOR U1736 ( .A(n1642), .B(n1641), .Z(n1644) );
  XOR U1737 ( .A(n1643), .B(n1644), .Z(n1659) );
  XNOR U1738 ( .A(n1659), .B(sreg[324]), .Z(n1661) );
  NANDN U1739 ( .A(n1636), .B(sreg[323]), .Z(n1640) );
  NAND U1740 ( .A(n1638), .B(n1637), .Z(n1639) );
  NAND U1741 ( .A(n1640), .B(n1639), .Z(n1660) );
  XOR U1742 ( .A(n1661), .B(n1660), .Z(c[324]) );
  NANDN U1743 ( .A(n1642), .B(n1641), .Z(n1646) );
  OR U1744 ( .A(n1644), .B(n1643), .Z(n1645) );
  AND U1745 ( .A(n1646), .B(n1645), .Z(n1666) );
  NAND U1746 ( .A(n31), .B(n1647), .Z(n1649) );
  XOR U1747 ( .A(b[3]), .B(a[71]), .Z(n1670) );
  NAND U1748 ( .A(n5811), .B(n1670), .Z(n1648) );
  AND U1749 ( .A(n1649), .B(n1648), .Z(n1678) );
  NAND U1750 ( .A(b[0]), .B(a[73]), .Z(n1650) );
  XNOR U1751 ( .A(b[1]), .B(n1650), .Z(n1652) );
  NANDN U1752 ( .A(b[0]), .B(a[72]), .Z(n1651) );
  NAND U1753 ( .A(n1652), .B(n1651), .Z(n1677) );
  AND U1754 ( .A(b[3]), .B(a[69]), .Z(n1676) );
  XOR U1755 ( .A(n1677), .B(n1676), .Z(n1679) );
  XOR U1756 ( .A(n1678), .B(n1679), .Z(n1665) );
  NANDN U1757 ( .A(n1654), .B(n1653), .Z(n1658) );
  OR U1758 ( .A(n1656), .B(n1655), .Z(n1657) );
  AND U1759 ( .A(n1658), .B(n1657), .Z(n1664) );
  XOR U1760 ( .A(n1665), .B(n1664), .Z(n1667) );
  XOR U1761 ( .A(n1666), .B(n1667), .Z(n1682) );
  XNOR U1762 ( .A(n1682), .B(sreg[325]), .Z(n1684) );
  NANDN U1763 ( .A(n1659), .B(sreg[324]), .Z(n1663) );
  NAND U1764 ( .A(n1661), .B(n1660), .Z(n1662) );
  NAND U1765 ( .A(n1663), .B(n1662), .Z(n1683) );
  XOR U1766 ( .A(n1684), .B(n1683), .Z(c[325]) );
  NANDN U1767 ( .A(n1665), .B(n1664), .Z(n1669) );
  OR U1768 ( .A(n1667), .B(n1666), .Z(n1668) );
  AND U1769 ( .A(n1669), .B(n1668), .Z(n1689) );
  NAND U1770 ( .A(n31), .B(n1670), .Z(n1672) );
  XOR U1771 ( .A(b[3]), .B(a[72]), .Z(n1693) );
  NAND U1772 ( .A(n5811), .B(n1693), .Z(n1671) );
  AND U1773 ( .A(n1672), .B(n1671), .Z(n1701) );
  NAND U1774 ( .A(b[0]), .B(a[74]), .Z(n1673) );
  XNOR U1775 ( .A(b[1]), .B(n1673), .Z(n1675) );
  NANDN U1776 ( .A(b[0]), .B(a[73]), .Z(n1674) );
  NAND U1777 ( .A(n1675), .B(n1674), .Z(n1700) );
  AND U1778 ( .A(b[3]), .B(a[70]), .Z(n1699) );
  XOR U1779 ( .A(n1700), .B(n1699), .Z(n1702) );
  XOR U1780 ( .A(n1701), .B(n1702), .Z(n1688) );
  NANDN U1781 ( .A(n1677), .B(n1676), .Z(n1681) );
  OR U1782 ( .A(n1679), .B(n1678), .Z(n1680) );
  AND U1783 ( .A(n1681), .B(n1680), .Z(n1687) );
  XOR U1784 ( .A(n1688), .B(n1687), .Z(n1690) );
  XOR U1785 ( .A(n1689), .B(n1690), .Z(n1705) );
  XNOR U1786 ( .A(n1705), .B(sreg[326]), .Z(n1707) );
  NANDN U1787 ( .A(n1682), .B(sreg[325]), .Z(n1686) );
  NAND U1788 ( .A(n1684), .B(n1683), .Z(n1685) );
  NAND U1789 ( .A(n1686), .B(n1685), .Z(n1706) );
  XOR U1790 ( .A(n1707), .B(n1706), .Z(c[326]) );
  NANDN U1791 ( .A(n1688), .B(n1687), .Z(n1692) );
  OR U1792 ( .A(n1690), .B(n1689), .Z(n1691) );
  AND U1793 ( .A(n1692), .B(n1691), .Z(n1712) );
  NAND U1794 ( .A(n31), .B(n1693), .Z(n1695) );
  XOR U1795 ( .A(b[3]), .B(a[73]), .Z(n1716) );
  NAND U1796 ( .A(n5811), .B(n1716), .Z(n1694) );
  AND U1797 ( .A(n1695), .B(n1694), .Z(n1724) );
  NAND U1798 ( .A(b[0]), .B(a[75]), .Z(n1696) );
  XNOR U1799 ( .A(b[1]), .B(n1696), .Z(n1698) );
  NANDN U1800 ( .A(b[0]), .B(a[74]), .Z(n1697) );
  NAND U1801 ( .A(n1698), .B(n1697), .Z(n1723) );
  AND U1802 ( .A(b[3]), .B(a[71]), .Z(n1722) );
  XOR U1803 ( .A(n1723), .B(n1722), .Z(n1725) );
  XOR U1804 ( .A(n1724), .B(n1725), .Z(n1711) );
  NANDN U1805 ( .A(n1700), .B(n1699), .Z(n1704) );
  OR U1806 ( .A(n1702), .B(n1701), .Z(n1703) );
  AND U1807 ( .A(n1704), .B(n1703), .Z(n1710) );
  XOR U1808 ( .A(n1711), .B(n1710), .Z(n1713) );
  XOR U1809 ( .A(n1712), .B(n1713), .Z(n1728) );
  XNOR U1810 ( .A(n1728), .B(sreg[327]), .Z(n1730) );
  NANDN U1811 ( .A(n1705), .B(sreg[326]), .Z(n1709) );
  NAND U1812 ( .A(n1707), .B(n1706), .Z(n1708) );
  NAND U1813 ( .A(n1709), .B(n1708), .Z(n1729) );
  XOR U1814 ( .A(n1730), .B(n1729), .Z(c[327]) );
  NANDN U1815 ( .A(n1711), .B(n1710), .Z(n1715) );
  OR U1816 ( .A(n1713), .B(n1712), .Z(n1714) );
  AND U1817 ( .A(n1715), .B(n1714), .Z(n1735) );
  NAND U1818 ( .A(n31), .B(n1716), .Z(n1718) );
  XOR U1819 ( .A(b[3]), .B(a[74]), .Z(n1739) );
  NAND U1820 ( .A(n5811), .B(n1739), .Z(n1717) );
  AND U1821 ( .A(n1718), .B(n1717), .Z(n1747) );
  NAND U1822 ( .A(b[0]), .B(a[76]), .Z(n1719) );
  XNOR U1823 ( .A(b[1]), .B(n1719), .Z(n1721) );
  NANDN U1824 ( .A(b[0]), .B(a[75]), .Z(n1720) );
  NAND U1825 ( .A(n1721), .B(n1720), .Z(n1746) );
  AND U1826 ( .A(b[3]), .B(a[72]), .Z(n1745) );
  XOR U1827 ( .A(n1746), .B(n1745), .Z(n1748) );
  XOR U1828 ( .A(n1747), .B(n1748), .Z(n1734) );
  NANDN U1829 ( .A(n1723), .B(n1722), .Z(n1727) );
  OR U1830 ( .A(n1725), .B(n1724), .Z(n1726) );
  AND U1831 ( .A(n1727), .B(n1726), .Z(n1733) );
  XOR U1832 ( .A(n1734), .B(n1733), .Z(n1736) );
  XOR U1833 ( .A(n1735), .B(n1736), .Z(n1751) );
  XNOR U1834 ( .A(n1751), .B(sreg[328]), .Z(n1753) );
  NANDN U1835 ( .A(n1728), .B(sreg[327]), .Z(n1732) );
  NAND U1836 ( .A(n1730), .B(n1729), .Z(n1731) );
  NAND U1837 ( .A(n1732), .B(n1731), .Z(n1752) );
  XOR U1838 ( .A(n1753), .B(n1752), .Z(c[328]) );
  NANDN U1839 ( .A(n1734), .B(n1733), .Z(n1738) );
  OR U1840 ( .A(n1736), .B(n1735), .Z(n1737) );
  AND U1841 ( .A(n1738), .B(n1737), .Z(n1758) );
  NAND U1842 ( .A(n31), .B(n1739), .Z(n1741) );
  XOR U1843 ( .A(b[3]), .B(a[75]), .Z(n1762) );
  NAND U1844 ( .A(n5811), .B(n1762), .Z(n1740) );
  AND U1845 ( .A(n1741), .B(n1740), .Z(n1770) );
  NAND U1846 ( .A(b[0]), .B(a[77]), .Z(n1742) );
  XNOR U1847 ( .A(b[1]), .B(n1742), .Z(n1744) );
  NANDN U1848 ( .A(b[0]), .B(a[76]), .Z(n1743) );
  NAND U1849 ( .A(n1744), .B(n1743), .Z(n1769) );
  AND U1850 ( .A(b[3]), .B(a[73]), .Z(n1768) );
  XOR U1851 ( .A(n1769), .B(n1768), .Z(n1771) );
  XOR U1852 ( .A(n1770), .B(n1771), .Z(n1757) );
  NANDN U1853 ( .A(n1746), .B(n1745), .Z(n1750) );
  OR U1854 ( .A(n1748), .B(n1747), .Z(n1749) );
  AND U1855 ( .A(n1750), .B(n1749), .Z(n1756) );
  XOR U1856 ( .A(n1757), .B(n1756), .Z(n1759) );
  XOR U1857 ( .A(n1758), .B(n1759), .Z(n1774) );
  XNOR U1858 ( .A(n1774), .B(sreg[329]), .Z(n1776) );
  NANDN U1859 ( .A(n1751), .B(sreg[328]), .Z(n1755) );
  NAND U1860 ( .A(n1753), .B(n1752), .Z(n1754) );
  NAND U1861 ( .A(n1755), .B(n1754), .Z(n1775) );
  XOR U1862 ( .A(n1776), .B(n1775), .Z(c[329]) );
  NANDN U1863 ( .A(n1757), .B(n1756), .Z(n1761) );
  OR U1864 ( .A(n1759), .B(n1758), .Z(n1760) );
  AND U1865 ( .A(n1761), .B(n1760), .Z(n1781) );
  NAND U1866 ( .A(n31), .B(n1762), .Z(n1764) );
  XOR U1867 ( .A(b[3]), .B(a[76]), .Z(n1785) );
  NAND U1868 ( .A(n5811), .B(n1785), .Z(n1763) );
  AND U1869 ( .A(n1764), .B(n1763), .Z(n1793) );
  AND U1870 ( .A(b[3]), .B(a[74]), .Z(n1791) );
  NAND U1871 ( .A(b[0]), .B(a[78]), .Z(n1765) );
  XNOR U1872 ( .A(b[1]), .B(n1765), .Z(n1767) );
  NANDN U1873 ( .A(b[0]), .B(a[77]), .Z(n1766) );
  NAND U1874 ( .A(n1767), .B(n1766), .Z(n1792) );
  XOR U1875 ( .A(n1791), .B(n1792), .Z(n1794) );
  XOR U1876 ( .A(n1793), .B(n1794), .Z(n1780) );
  NANDN U1877 ( .A(n1769), .B(n1768), .Z(n1773) );
  OR U1878 ( .A(n1771), .B(n1770), .Z(n1772) );
  AND U1879 ( .A(n1773), .B(n1772), .Z(n1779) );
  XOR U1880 ( .A(n1780), .B(n1779), .Z(n1782) );
  XOR U1881 ( .A(n1781), .B(n1782), .Z(n1797) );
  XNOR U1882 ( .A(n1797), .B(sreg[330]), .Z(n1799) );
  NANDN U1883 ( .A(n1774), .B(sreg[329]), .Z(n1778) );
  NAND U1884 ( .A(n1776), .B(n1775), .Z(n1777) );
  NAND U1885 ( .A(n1778), .B(n1777), .Z(n1798) );
  XOR U1886 ( .A(n1799), .B(n1798), .Z(c[330]) );
  NANDN U1887 ( .A(n1780), .B(n1779), .Z(n1784) );
  OR U1888 ( .A(n1782), .B(n1781), .Z(n1783) );
  AND U1889 ( .A(n1784), .B(n1783), .Z(n1804) );
  NAND U1890 ( .A(n31), .B(n1785), .Z(n1787) );
  XOR U1891 ( .A(b[3]), .B(a[77]), .Z(n1808) );
  NAND U1892 ( .A(n5811), .B(n1808), .Z(n1786) );
  AND U1893 ( .A(n1787), .B(n1786), .Z(n1816) );
  NAND U1894 ( .A(b[0]), .B(a[79]), .Z(n1788) );
  XNOR U1895 ( .A(b[1]), .B(n1788), .Z(n1790) );
  NANDN U1896 ( .A(b[0]), .B(a[78]), .Z(n1789) );
  NAND U1897 ( .A(n1790), .B(n1789), .Z(n1815) );
  AND U1898 ( .A(b[3]), .B(a[75]), .Z(n1814) );
  XOR U1899 ( .A(n1815), .B(n1814), .Z(n1817) );
  XOR U1900 ( .A(n1816), .B(n1817), .Z(n1803) );
  NANDN U1901 ( .A(n1792), .B(n1791), .Z(n1796) );
  OR U1902 ( .A(n1794), .B(n1793), .Z(n1795) );
  AND U1903 ( .A(n1796), .B(n1795), .Z(n1802) );
  XOR U1904 ( .A(n1803), .B(n1802), .Z(n1805) );
  XOR U1905 ( .A(n1804), .B(n1805), .Z(n1820) );
  XNOR U1906 ( .A(n1820), .B(sreg[331]), .Z(n1822) );
  NANDN U1907 ( .A(n1797), .B(sreg[330]), .Z(n1801) );
  NAND U1908 ( .A(n1799), .B(n1798), .Z(n1800) );
  NAND U1909 ( .A(n1801), .B(n1800), .Z(n1821) );
  XOR U1910 ( .A(n1822), .B(n1821), .Z(c[331]) );
  NANDN U1911 ( .A(n1803), .B(n1802), .Z(n1807) );
  OR U1912 ( .A(n1805), .B(n1804), .Z(n1806) );
  AND U1913 ( .A(n1807), .B(n1806), .Z(n1827) );
  NAND U1914 ( .A(n31), .B(n1808), .Z(n1810) );
  XOR U1915 ( .A(b[3]), .B(a[78]), .Z(n1831) );
  NAND U1916 ( .A(n5811), .B(n1831), .Z(n1809) );
  AND U1917 ( .A(n1810), .B(n1809), .Z(n1839) );
  AND U1918 ( .A(b[3]), .B(a[76]), .Z(n1837) );
  NAND U1919 ( .A(b[0]), .B(a[80]), .Z(n1811) );
  XNOR U1920 ( .A(b[1]), .B(n1811), .Z(n1813) );
  NANDN U1921 ( .A(b[0]), .B(a[79]), .Z(n1812) );
  NAND U1922 ( .A(n1813), .B(n1812), .Z(n1838) );
  XOR U1923 ( .A(n1837), .B(n1838), .Z(n1840) );
  XOR U1924 ( .A(n1839), .B(n1840), .Z(n1826) );
  NANDN U1925 ( .A(n1815), .B(n1814), .Z(n1819) );
  OR U1926 ( .A(n1817), .B(n1816), .Z(n1818) );
  AND U1927 ( .A(n1819), .B(n1818), .Z(n1825) );
  XOR U1928 ( .A(n1826), .B(n1825), .Z(n1828) );
  XOR U1929 ( .A(n1827), .B(n1828), .Z(n1843) );
  XNOR U1930 ( .A(n1843), .B(sreg[332]), .Z(n1845) );
  NANDN U1931 ( .A(n1820), .B(sreg[331]), .Z(n1824) );
  NAND U1932 ( .A(n1822), .B(n1821), .Z(n1823) );
  NAND U1933 ( .A(n1824), .B(n1823), .Z(n1844) );
  XOR U1934 ( .A(n1845), .B(n1844), .Z(c[332]) );
  NANDN U1935 ( .A(n1826), .B(n1825), .Z(n1830) );
  OR U1936 ( .A(n1828), .B(n1827), .Z(n1829) );
  AND U1937 ( .A(n1830), .B(n1829), .Z(n1850) );
  NAND U1938 ( .A(n31), .B(n1831), .Z(n1833) );
  XOR U1939 ( .A(b[3]), .B(a[79]), .Z(n1854) );
  NAND U1940 ( .A(n5811), .B(n1854), .Z(n1832) );
  AND U1941 ( .A(n1833), .B(n1832), .Z(n1862) );
  NAND U1942 ( .A(b[0]), .B(a[81]), .Z(n1834) );
  XNOR U1943 ( .A(b[1]), .B(n1834), .Z(n1836) );
  NANDN U1944 ( .A(b[0]), .B(a[80]), .Z(n1835) );
  NAND U1945 ( .A(n1836), .B(n1835), .Z(n1861) );
  AND U1946 ( .A(b[3]), .B(a[77]), .Z(n1860) );
  XOR U1947 ( .A(n1861), .B(n1860), .Z(n1863) );
  XOR U1948 ( .A(n1862), .B(n1863), .Z(n1849) );
  NANDN U1949 ( .A(n1838), .B(n1837), .Z(n1842) );
  OR U1950 ( .A(n1840), .B(n1839), .Z(n1841) );
  AND U1951 ( .A(n1842), .B(n1841), .Z(n1848) );
  XOR U1952 ( .A(n1849), .B(n1848), .Z(n1851) );
  XOR U1953 ( .A(n1850), .B(n1851), .Z(n1866) );
  XNOR U1954 ( .A(n1866), .B(sreg[333]), .Z(n1868) );
  NANDN U1955 ( .A(n1843), .B(sreg[332]), .Z(n1847) );
  NAND U1956 ( .A(n1845), .B(n1844), .Z(n1846) );
  NAND U1957 ( .A(n1847), .B(n1846), .Z(n1867) );
  XOR U1958 ( .A(n1868), .B(n1867), .Z(c[333]) );
  NANDN U1959 ( .A(n1849), .B(n1848), .Z(n1853) );
  OR U1960 ( .A(n1851), .B(n1850), .Z(n1852) );
  AND U1961 ( .A(n1853), .B(n1852), .Z(n1873) );
  NAND U1962 ( .A(n31), .B(n1854), .Z(n1856) );
  XOR U1963 ( .A(b[3]), .B(a[80]), .Z(n1877) );
  NAND U1964 ( .A(n5811), .B(n1877), .Z(n1855) );
  AND U1965 ( .A(n1856), .B(n1855), .Z(n1885) );
  AND U1966 ( .A(b[3]), .B(a[78]), .Z(n1883) );
  NAND U1967 ( .A(b[0]), .B(a[82]), .Z(n1857) );
  XNOR U1968 ( .A(b[1]), .B(n1857), .Z(n1859) );
  NANDN U1969 ( .A(b[0]), .B(a[81]), .Z(n1858) );
  NAND U1970 ( .A(n1859), .B(n1858), .Z(n1884) );
  XOR U1971 ( .A(n1883), .B(n1884), .Z(n1886) );
  XOR U1972 ( .A(n1885), .B(n1886), .Z(n1872) );
  NANDN U1973 ( .A(n1861), .B(n1860), .Z(n1865) );
  OR U1974 ( .A(n1863), .B(n1862), .Z(n1864) );
  AND U1975 ( .A(n1865), .B(n1864), .Z(n1871) );
  XOR U1976 ( .A(n1872), .B(n1871), .Z(n1874) );
  XOR U1977 ( .A(n1873), .B(n1874), .Z(n1889) );
  XNOR U1978 ( .A(n1889), .B(sreg[334]), .Z(n1891) );
  NANDN U1979 ( .A(n1866), .B(sreg[333]), .Z(n1870) );
  NAND U1980 ( .A(n1868), .B(n1867), .Z(n1869) );
  NAND U1981 ( .A(n1870), .B(n1869), .Z(n1890) );
  XOR U1982 ( .A(n1891), .B(n1890), .Z(c[334]) );
  NANDN U1983 ( .A(n1872), .B(n1871), .Z(n1876) );
  OR U1984 ( .A(n1874), .B(n1873), .Z(n1875) );
  AND U1985 ( .A(n1876), .B(n1875), .Z(n1896) );
  NAND U1986 ( .A(n31), .B(n1877), .Z(n1879) );
  XOR U1987 ( .A(b[3]), .B(a[81]), .Z(n1900) );
  NAND U1988 ( .A(n5811), .B(n1900), .Z(n1878) );
  AND U1989 ( .A(n1879), .B(n1878), .Z(n1908) );
  NAND U1990 ( .A(b[0]), .B(a[83]), .Z(n1880) );
  XNOR U1991 ( .A(b[1]), .B(n1880), .Z(n1882) );
  NANDN U1992 ( .A(b[0]), .B(a[82]), .Z(n1881) );
  NAND U1993 ( .A(n1882), .B(n1881), .Z(n1907) );
  AND U1994 ( .A(b[3]), .B(a[79]), .Z(n1906) );
  XOR U1995 ( .A(n1907), .B(n1906), .Z(n1909) );
  XOR U1996 ( .A(n1908), .B(n1909), .Z(n1895) );
  NANDN U1997 ( .A(n1884), .B(n1883), .Z(n1888) );
  OR U1998 ( .A(n1886), .B(n1885), .Z(n1887) );
  AND U1999 ( .A(n1888), .B(n1887), .Z(n1894) );
  XOR U2000 ( .A(n1895), .B(n1894), .Z(n1897) );
  XOR U2001 ( .A(n1896), .B(n1897), .Z(n1912) );
  XNOR U2002 ( .A(n1912), .B(sreg[335]), .Z(n1914) );
  NANDN U2003 ( .A(n1889), .B(sreg[334]), .Z(n1893) );
  NAND U2004 ( .A(n1891), .B(n1890), .Z(n1892) );
  NAND U2005 ( .A(n1893), .B(n1892), .Z(n1913) );
  XOR U2006 ( .A(n1914), .B(n1913), .Z(c[335]) );
  NANDN U2007 ( .A(n1895), .B(n1894), .Z(n1899) );
  OR U2008 ( .A(n1897), .B(n1896), .Z(n1898) );
  AND U2009 ( .A(n1899), .B(n1898), .Z(n1919) );
  NAND U2010 ( .A(n31), .B(n1900), .Z(n1902) );
  XOR U2011 ( .A(b[3]), .B(a[82]), .Z(n1923) );
  NAND U2012 ( .A(n5811), .B(n1923), .Z(n1901) );
  AND U2013 ( .A(n1902), .B(n1901), .Z(n1931) );
  NAND U2014 ( .A(b[0]), .B(a[84]), .Z(n1903) );
  XNOR U2015 ( .A(b[1]), .B(n1903), .Z(n1905) );
  NANDN U2016 ( .A(b[0]), .B(a[83]), .Z(n1904) );
  NAND U2017 ( .A(n1905), .B(n1904), .Z(n1930) );
  AND U2018 ( .A(b[3]), .B(a[80]), .Z(n1929) );
  XOR U2019 ( .A(n1930), .B(n1929), .Z(n1932) );
  XOR U2020 ( .A(n1931), .B(n1932), .Z(n1918) );
  NANDN U2021 ( .A(n1907), .B(n1906), .Z(n1911) );
  OR U2022 ( .A(n1909), .B(n1908), .Z(n1910) );
  AND U2023 ( .A(n1911), .B(n1910), .Z(n1917) );
  XOR U2024 ( .A(n1918), .B(n1917), .Z(n1920) );
  XOR U2025 ( .A(n1919), .B(n1920), .Z(n1935) );
  XNOR U2026 ( .A(n1935), .B(sreg[336]), .Z(n1937) );
  NANDN U2027 ( .A(n1912), .B(sreg[335]), .Z(n1916) );
  NAND U2028 ( .A(n1914), .B(n1913), .Z(n1915) );
  NAND U2029 ( .A(n1916), .B(n1915), .Z(n1936) );
  XOR U2030 ( .A(n1937), .B(n1936), .Z(c[336]) );
  NANDN U2031 ( .A(n1918), .B(n1917), .Z(n1922) );
  OR U2032 ( .A(n1920), .B(n1919), .Z(n1921) );
  AND U2033 ( .A(n1922), .B(n1921), .Z(n1942) );
  NAND U2034 ( .A(n31), .B(n1923), .Z(n1925) );
  XOR U2035 ( .A(b[3]), .B(a[83]), .Z(n1946) );
  NAND U2036 ( .A(n5811), .B(n1946), .Z(n1924) );
  AND U2037 ( .A(n1925), .B(n1924), .Z(n1954) );
  AND U2038 ( .A(b[3]), .B(a[81]), .Z(n1952) );
  NAND U2039 ( .A(b[0]), .B(a[85]), .Z(n1926) );
  XNOR U2040 ( .A(b[1]), .B(n1926), .Z(n1928) );
  NANDN U2041 ( .A(b[0]), .B(a[84]), .Z(n1927) );
  NAND U2042 ( .A(n1928), .B(n1927), .Z(n1953) );
  XOR U2043 ( .A(n1952), .B(n1953), .Z(n1955) );
  XOR U2044 ( .A(n1954), .B(n1955), .Z(n1941) );
  NANDN U2045 ( .A(n1930), .B(n1929), .Z(n1934) );
  OR U2046 ( .A(n1932), .B(n1931), .Z(n1933) );
  AND U2047 ( .A(n1934), .B(n1933), .Z(n1940) );
  XOR U2048 ( .A(n1941), .B(n1940), .Z(n1943) );
  XOR U2049 ( .A(n1942), .B(n1943), .Z(n1958) );
  XNOR U2050 ( .A(n1958), .B(sreg[337]), .Z(n1960) );
  NANDN U2051 ( .A(n1935), .B(sreg[336]), .Z(n1939) );
  NAND U2052 ( .A(n1937), .B(n1936), .Z(n1938) );
  NAND U2053 ( .A(n1939), .B(n1938), .Z(n1959) );
  XOR U2054 ( .A(n1960), .B(n1959), .Z(c[337]) );
  NANDN U2055 ( .A(n1941), .B(n1940), .Z(n1945) );
  OR U2056 ( .A(n1943), .B(n1942), .Z(n1944) );
  AND U2057 ( .A(n1945), .B(n1944), .Z(n1965) );
  NAND U2058 ( .A(n31), .B(n1946), .Z(n1948) );
  XOR U2059 ( .A(b[3]), .B(a[84]), .Z(n1969) );
  NAND U2060 ( .A(n5811), .B(n1969), .Z(n1947) );
  AND U2061 ( .A(n1948), .B(n1947), .Z(n1977) );
  NAND U2062 ( .A(b[0]), .B(a[86]), .Z(n1949) );
  XNOR U2063 ( .A(b[1]), .B(n1949), .Z(n1951) );
  NANDN U2064 ( .A(b[0]), .B(a[85]), .Z(n1950) );
  NAND U2065 ( .A(n1951), .B(n1950), .Z(n1976) );
  AND U2066 ( .A(b[3]), .B(a[82]), .Z(n1975) );
  XOR U2067 ( .A(n1976), .B(n1975), .Z(n1978) );
  XOR U2068 ( .A(n1977), .B(n1978), .Z(n1964) );
  NANDN U2069 ( .A(n1953), .B(n1952), .Z(n1957) );
  OR U2070 ( .A(n1955), .B(n1954), .Z(n1956) );
  AND U2071 ( .A(n1957), .B(n1956), .Z(n1963) );
  XOR U2072 ( .A(n1964), .B(n1963), .Z(n1966) );
  XOR U2073 ( .A(n1965), .B(n1966), .Z(n1981) );
  XNOR U2074 ( .A(n1981), .B(sreg[338]), .Z(n1983) );
  NANDN U2075 ( .A(n1958), .B(sreg[337]), .Z(n1962) );
  NAND U2076 ( .A(n1960), .B(n1959), .Z(n1961) );
  NAND U2077 ( .A(n1962), .B(n1961), .Z(n1982) );
  XOR U2078 ( .A(n1983), .B(n1982), .Z(c[338]) );
  NANDN U2079 ( .A(n1964), .B(n1963), .Z(n1968) );
  OR U2080 ( .A(n1966), .B(n1965), .Z(n1967) );
  AND U2081 ( .A(n1968), .B(n1967), .Z(n1988) );
  NAND U2082 ( .A(n31), .B(n1969), .Z(n1971) );
  XOR U2083 ( .A(b[3]), .B(a[85]), .Z(n1992) );
  NAND U2084 ( .A(n5811), .B(n1992), .Z(n1970) );
  AND U2085 ( .A(n1971), .B(n1970), .Z(n2000) );
  NAND U2086 ( .A(b[0]), .B(a[87]), .Z(n1972) );
  XNOR U2087 ( .A(b[1]), .B(n1972), .Z(n1974) );
  NANDN U2088 ( .A(b[0]), .B(a[86]), .Z(n1973) );
  NAND U2089 ( .A(n1974), .B(n1973), .Z(n1999) );
  AND U2090 ( .A(b[3]), .B(a[83]), .Z(n1998) );
  XOR U2091 ( .A(n1999), .B(n1998), .Z(n2001) );
  XOR U2092 ( .A(n2000), .B(n2001), .Z(n1987) );
  NANDN U2093 ( .A(n1976), .B(n1975), .Z(n1980) );
  OR U2094 ( .A(n1978), .B(n1977), .Z(n1979) );
  AND U2095 ( .A(n1980), .B(n1979), .Z(n1986) );
  XOR U2096 ( .A(n1987), .B(n1986), .Z(n1989) );
  XOR U2097 ( .A(n1988), .B(n1989), .Z(n2004) );
  XNOR U2098 ( .A(n2004), .B(sreg[339]), .Z(n2006) );
  NANDN U2099 ( .A(n1981), .B(sreg[338]), .Z(n1985) );
  NAND U2100 ( .A(n1983), .B(n1982), .Z(n1984) );
  NAND U2101 ( .A(n1985), .B(n1984), .Z(n2005) );
  XOR U2102 ( .A(n2006), .B(n2005), .Z(c[339]) );
  NANDN U2103 ( .A(n1987), .B(n1986), .Z(n1991) );
  OR U2104 ( .A(n1989), .B(n1988), .Z(n1990) );
  AND U2105 ( .A(n1991), .B(n1990), .Z(n2011) );
  NAND U2106 ( .A(n31), .B(n1992), .Z(n1994) );
  XOR U2107 ( .A(b[3]), .B(a[86]), .Z(n2015) );
  NAND U2108 ( .A(n5811), .B(n2015), .Z(n1993) );
  AND U2109 ( .A(n1994), .B(n1993), .Z(n2023) );
  AND U2110 ( .A(b[3]), .B(a[84]), .Z(n2021) );
  NAND U2111 ( .A(b[0]), .B(a[88]), .Z(n1995) );
  XNOR U2112 ( .A(b[1]), .B(n1995), .Z(n1997) );
  NANDN U2113 ( .A(b[0]), .B(a[87]), .Z(n1996) );
  NAND U2114 ( .A(n1997), .B(n1996), .Z(n2022) );
  XOR U2115 ( .A(n2021), .B(n2022), .Z(n2024) );
  XOR U2116 ( .A(n2023), .B(n2024), .Z(n2010) );
  NANDN U2117 ( .A(n1999), .B(n1998), .Z(n2003) );
  OR U2118 ( .A(n2001), .B(n2000), .Z(n2002) );
  AND U2119 ( .A(n2003), .B(n2002), .Z(n2009) );
  XOR U2120 ( .A(n2010), .B(n2009), .Z(n2012) );
  XOR U2121 ( .A(n2011), .B(n2012), .Z(n2027) );
  XNOR U2122 ( .A(n2027), .B(sreg[340]), .Z(n2029) );
  NANDN U2123 ( .A(n2004), .B(sreg[339]), .Z(n2008) );
  NAND U2124 ( .A(n2006), .B(n2005), .Z(n2007) );
  NAND U2125 ( .A(n2008), .B(n2007), .Z(n2028) );
  XOR U2126 ( .A(n2029), .B(n2028), .Z(c[340]) );
  NANDN U2127 ( .A(n2010), .B(n2009), .Z(n2014) );
  OR U2128 ( .A(n2012), .B(n2011), .Z(n2013) );
  AND U2129 ( .A(n2014), .B(n2013), .Z(n2034) );
  NAND U2130 ( .A(n31), .B(n2015), .Z(n2017) );
  XOR U2131 ( .A(b[3]), .B(a[87]), .Z(n2038) );
  NAND U2132 ( .A(n5811), .B(n2038), .Z(n2016) );
  AND U2133 ( .A(n2017), .B(n2016), .Z(n2046) );
  NAND U2134 ( .A(b[0]), .B(a[89]), .Z(n2018) );
  XNOR U2135 ( .A(b[1]), .B(n2018), .Z(n2020) );
  NANDN U2136 ( .A(b[0]), .B(a[88]), .Z(n2019) );
  NAND U2137 ( .A(n2020), .B(n2019), .Z(n2045) );
  AND U2138 ( .A(b[3]), .B(a[85]), .Z(n2044) );
  XOR U2139 ( .A(n2045), .B(n2044), .Z(n2047) );
  XOR U2140 ( .A(n2046), .B(n2047), .Z(n2033) );
  NANDN U2141 ( .A(n2022), .B(n2021), .Z(n2026) );
  OR U2142 ( .A(n2024), .B(n2023), .Z(n2025) );
  AND U2143 ( .A(n2026), .B(n2025), .Z(n2032) );
  XOR U2144 ( .A(n2033), .B(n2032), .Z(n2035) );
  XOR U2145 ( .A(n2034), .B(n2035), .Z(n2050) );
  XNOR U2146 ( .A(n2050), .B(sreg[341]), .Z(n2052) );
  NANDN U2147 ( .A(n2027), .B(sreg[340]), .Z(n2031) );
  NAND U2148 ( .A(n2029), .B(n2028), .Z(n2030) );
  NAND U2149 ( .A(n2031), .B(n2030), .Z(n2051) );
  XOR U2150 ( .A(n2052), .B(n2051), .Z(c[341]) );
  NANDN U2151 ( .A(n2033), .B(n2032), .Z(n2037) );
  OR U2152 ( .A(n2035), .B(n2034), .Z(n2036) );
  AND U2153 ( .A(n2037), .B(n2036), .Z(n2057) );
  NAND U2154 ( .A(n31), .B(n2038), .Z(n2040) );
  XOR U2155 ( .A(b[3]), .B(a[88]), .Z(n2061) );
  NAND U2156 ( .A(n5811), .B(n2061), .Z(n2039) );
  AND U2157 ( .A(n2040), .B(n2039), .Z(n2069) );
  AND U2158 ( .A(b[3]), .B(a[86]), .Z(n2067) );
  NAND U2159 ( .A(b[0]), .B(a[90]), .Z(n2041) );
  XNOR U2160 ( .A(b[1]), .B(n2041), .Z(n2043) );
  NANDN U2161 ( .A(b[0]), .B(a[89]), .Z(n2042) );
  NAND U2162 ( .A(n2043), .B(n2042), .Z(n2068) );
  XOR U2163 ( .A(n2067), .B(n2068), .Z(n2070) );
  XOR U2164 ( .A(n2069), .B(n2070), .Z(n2056) );
  NANDN U2165 ( .A(n2045), .B(n2044), .Z(n2049) );
  OR U2166 ( .A(n2047), .B(n2046), .Z(n2048) );
  AND U2167 ( .A(n2049), .B(n2048), .Z(n2055) );
  XOR U2168 ( .A(n2056), .B(n2055), .Z(n2058) );
  XOR U2169 ( .A(n2057), .B(n2058), .Z(n2073) );
  XNOR U2170 ( .A(n2073), .B(sreg[342]), .Z(n2075) );
  NANDN U2171 ( .A(n2050), .B(sreg[341]), .Z(n2054) );
  NAND U2172 ( .A(n2052), .B(n2051), .Z(n2053) );
  NAND U2173 ( .A(n2054), .B(n2053), .Z(n2074) );
  XOR U2174 ( .A(n2075), .B(n2074), .Z(c[342]) );
  NANDN U2175 ( .A(n2056), .B(n2055), .Z(n2060) );
  OR U2176 ( .A(n2058), .B(n2057), .Z(n2059) );
  AND U2177 ( .A(n2060), .B(n2059), .Z(n2080) );
  NAND U2178 ( .A(n31), .B(n2061), .Z(n2063) );
  XOR U2179 ( .A(b[3]), .B(a[89]), .Z(n2084) );
  NAND U2180 ( .A(n5811), .B(n2084), .Z(n2062) );
  AND U2181 ( .A(n2063), .B(n2062), .Z(n2092) );
  NAND U2182 ( .A(b[0]), .B(a[91]), .Z(n2064) );
  XNOR U2183 ( .A(b[1]), .B(n2064), .Z(n2066) );
  NANDN U2184 ( .A(b[0]), .B(a[90]), .Z(n2065) );
  NAND U2185 ( .A(n2066), .B(n2065), .Z(n2091) );
  AND U2186 ( .A(b[3]), .B(a[87]), .Z(n2090) );
  XOR U2187 ( .A(n2091), .B(n2090), .Z(n2093) );
  XOR U2188 ( .A(n2092), .B(n2093), .Z(n2079) );
  NANDN U2189 ( .A(n2068), .B(n2067), .Z(n2072) );
  OR U2190 ( .A(n2070), .B(n2069), .Z(n2071) );
  AND U2191 ( .A(n2072), .B(n2071), .Z(n2078) );
  XOR U2192 ( .A(n2079), .B(n2078), .Z(n2081) );
  XOR U2193 ( .A(n2080), .B(n2081), .Z(n2096) );
  XNOR U2194 ( .A(n2096), .B(sreg[343]), .Z(n2098) );
  NANDN U2195 ( .A(n2073), .B(sreg[342]), .Z(n2077) );
  NAND U2196 ( .A(n2075), .B(n2074), .Z(n2076) );
  NAND U2197 ( .A(n2077), .B(n2076), .Z(n2097) );
  XOR U2198 ( .A(n2098), .B(n2097), .Z(c[343]) );
  NANDN U2199 ( .A(n2079), .B(n2078), .Z(n2083) );
  OR U2200 ( .A(n2081), .B(n2080), .Z(n2082) );
  AND U2201 ( .A(n2083), .B(n2082), .Z(n2103) );
  NAND U2202 ( .A(n31), .B(n2084), .Z(n2086) );
  XOR U2203 ( .A(b[3]), .B(a[90]), .Z(n2107) );
  NAND U2204 ( .A(n5811), .B(n2107), .Z(n2085) );
  AND U2205 ( .A(n2086), .B(n2085), .Z(n2115) );
  NAND U2206 ( .A(b[0]), .B(a[92]), .Z(n2087) );
  XNOR U2207 ( .A(b[1]), .B(n2087), .Z(n2089) );
  NANDN U2208 ( .A(b[0]), .B(a[91]), .Z(n2088) );
  NAND U2209 ( .A(n2089), .B(n2088), .Z(n2114) );
  AND U2210 ( .A(b[3]), .B(a[88]), .Z(n2113) );
  XOR U2211 ( .A(n2114), .B(n2113), .Z(n2116) );
  XOR U2212 ( .A(n2115), .B(n2116), .Z(n2102) );
  NANDN U2213 ( .A(n2091), .B(n2090), .Z(n2095) );
  OR U2214 ( .A(n2093), .B(n2092), .Z(n2094) );
  AND U2215 ( .A(n2095), .B(n2094), .Z(n2101) );
  XOR U2216 ( .A(n2102), .B(n2101), .Z(n2104) );
  XOR U2217 ( .A(n2103), .B(n2104), .Z(n2119) );
  XNOR U2218 ( .A(n2119), .B(sreg[344]), .Z(n2121) );
  NANDN U2219 ( .A(n2096), .B(sreg[343]), .Z(n2100) );
  NAND U2220 ( .A(n2098), .B(n2097), .Z(n2099) );
  NAND U2221 ( .A(n2100), .B(n2099), .Z(n2120) );
  XOR U2222 ( .A(n2121), .B(n2120), .Z(c[344]) );
  NANDN U2223 ( .A(n2102), .B(n2101), .Z(n2106) );
  OR U2224 ( .A(n2104), .B(n2103), .Z(n2105) );
  AND U2225 ( .A(n2106), .B(n2105), .Z(n2126) );
  NAND U2226 ( .A(n31), .B(n2107), .Z(n2109) );
  XOR U2227 ( .A(b[3]), .B(a[91]), .Z(n2130) );
  NAND U2228 ( .A(n5811), .B(n2130), .Z(n2108) );
  AND U2229 ( .A(n2109), .B(n2108), .Z(n2138) );
  NAND U2230 ( .A(b[0]), .B(a[93]), .Z(n2110) );
  XNOR U2231 ( .A(b[1]), .B(n2110), .Z(n2112) );
  NANDN U2232 ( .A(b[0]), .B(a[92]), .Z(n2111) );
  NAND U2233 ( .A(n2112), .B(n2111), .Z(n2137) );
  AND U2234 ( .A(b[3]), .B(a[89]), .Z(n2136) );
  XOR U2235 ( .A(n2137), .B(n2136), .Z(n2139) );
  XOR U2236 ( .A(n2138), .B(n2139), .Z(n2125) );
  NANDN U2237 ( .A(n2114), .B(n2113), .Z(n2118) );
  OR U2238 ( .A(n2116), .B(n2115), .Z(n2117) );
  AND U2239 ( .A(n2118), .B(n2117), .Z(n2124) );
  XOR U2240 ( .A(n2125), .B(n2124), .Z(n2127) );
  XOR U2241 ( .A(n2126), .B(n2127), .Z(n2142) );
  XNOR U2242 ( .A(n2142), .B(sreg[345]), .Z(n2144) );
  NANDN U2243 ( .A(n2119), .B(sreg[344]), .Z(n2123) );
  NAND U2244 ( .A(n2121), .B(n2120), .Z(n2122) );
  NAND U2245 ( .A(n2123), .B(n2122), .Z(n2143) );
  XOR U2246 ( .A(n2144), .B(n2143), .Z(c[345]) );
  NANDN U2247 ( .A(n2125), .B(n2124), .Z(n2129) );
  OR U2248 ( .A(n2127), .B(n2126), .Z(n2128) );
  AND U2249 ( .A(n2129), .B(n2128), .Z(n2149) );
  NAND U2250 ( .A(n31), .B(n2130), .Z(n2132) );
  XOR U2251 ( .A(b[3]), .B(a[92]), .Z(n2153) );
  NAND U2252 ( .A(n5811), .B(n2153), .Z(n2131) );
  AND U2253 ( .A(n2132), .B(n2131), .Z(n2161) );
  NAND U2254 ( .A(b[0]), .B(a[94]), .Z(n2133) );
  XNOR U2255 ( .A(b[1]), .B(n2133), .Z(n2135) );
  NANDN U2256 ( .A(b[0]), .B(a[93]), .Z(n2134) );
  NAND U2257 ( .A(n2135), .B(n2134), .Z(n2160) );
  AND U2258 ( .A(b[3]), .B(a[90]), .Z(n2159) );
  XOR U2259 ( .A(n2160), .B(n2159), .Z(n2162) );
  XOR U2260 ( .A(n2161), .B(n2162), .Z(n2148) );
  NANDN U2261 ( .A(n2137), .B(n2136), .Z(n2141) );
  OR U2262 ( .A(n2139), .B(n2138), .Z(n2140) );
  AND U2263 ( .A(n2141), .B(n2140), .Z(n2147) );
  XOR U2264 ( .A(n2148), .B(n2147), .Z(n2150) );
  XOR U2265 ( .A(n2149), .B(n2150), .Z(n2165) );
  XNOR U2266 ( .A(n2165), .B(sreg[346]), .Z(n2167) );
  NANDN U2267 ( .A(n2142), .B(sreg[345]), .Z(n2146) );
  NAND U2268 ( .A(n2144), .B(n2143), .Z(n2145) );
  NAND U2269 ( .A(n2146), .B(n2145), .Z(n2166) );
  XOR U2270 ( .A(n2167), .B(n2166), .Z(c[346]) );
  NANDN U2271 ( .A(n2148), .B(n2147), .Z(n2152) );
  OR U2272 ( .A(n2150), .B(n2149), .Z(n2151) );
  AND U2273 ( .A(n2152), .B(n2151), .Z(n2172) );
  NAND U2274 ( .A(n31), .B(n2153), .Z(n2155) );
  XOR U2275 ( .A(b[3]), .B(a[93]), .Z(n2176) );
  NAND U2276 ( .A(n5811), .B(n2176), .Z(n2154) );
  AND U2277 ( .A(n2155), .B(n2154), .Z(n2184) );
  NAND U2278 ( .A(b[0]), .B(a[95]), .Z(n2156) );
  XNOR U2279 ( .A(b[1]), .B(n2156), .Z(n2158) );
  NANDN U2280 ( .A(b[0]), .B(a[94]), .Z(n2157) );
  NAND U2281 ( .A(n2158), .B(n2157), .Z(n2183) );
  AND U2282 ( .A(b[3]), .B(a[91]), .Z(n2182) );
  XOR U2283 ( .A(n2183), .B(n2182), .Z(n2185) );
  XOR U2284 ( .A(n2184), .B(n2185), .Z(n2171) );
  NANDN U2285 ( .A(n2160), .B(n2159), .Z(n2164) );
  OR U2286 ( .A(n2162), .B(n2161), .Z(n2163) );
  AND U2287 ( .A(n2164), .B(n2163), .Z(n2170) );
  XOR U2288 ( .A(n2171), .B(n2170), .Z(n2173) );
  XOR U2289 ( .A(n2172), .B(n2173), .Z(n2188) );
  XNOR U2290 ( .A(n2188), .B(sreg[347]), .Z(n2190) );
  NANDN U2291 ( .A(n2165), .B(sreg[346]), .Z(n2169) );
  NAND U2292 ( .A(n2167), .B(n2166), .Z(n2168) );
  NAND U2293 ( .A(n2169), .B(n2168), .Z(n2189) );
  XOR U2294 ( .A(n2190), .B(n2189), .Z(c[347]) );
  NANDN U2295 ( .A(n2171), .B(n2170), .Z(n2175) );
  OR U2296 ( .A(n2173), .B(n2172), .Z(n2174) );
  AND U2297 ( .A(n2175), .B(n2174), .Z(n2195) );
  NAND U2298 ( .A(n31), .B(n2176), .Z(n2178) );
  XOR U2299 ( .A(b[3]), .B(a[94]), .Z(n2199) );
  NAND U2300 ( .A(n5811), .B(n2199), .Z(n2177) );
  AND U2301 ( .A(n2178), .B(n2177), .Z(n2207) );
  NAND U2302 ( .A(b[0]), .B(a[96]), .Z(n2179) );
  XNOR U2303 ( .A(b[1]), .B(n2179), .Z(n2181) );
  NANDN U2304 ( .A(b[0]), .B(a[95]), .Z(n2180) );
  NAND U2305 ( .A(n2181), .B(n2180), .Z(n2206) );
  AND U2306 ( .A(b[3]), .B(a[92]), .Z(n2205) );
  XOR U2307 ( .A(n2206), .B(n2205), .Z(n2208) );
  XOR U2308 ( .A(n2207), .B(n2208), .Z(n2194) );
  NANDN U2309 ( .A(n2183), .B(n2182), .Z(n2187) );
  OR U2310 ( .A(n2185), .B(n2184), .Z(n2186) );
  AND U2311 ( .A(n2187), .B(n2186), .Z(n2193) );
  XOR U2312 ( .A(n2194), .B(n2193), .Z(n2196) );
  XOR U2313 ( .A(n2195), .B(n2196), .Z(n2211) );
  XNOR U2314 ( .A(n2211), .B(sreg[348]), .Z(n2213) );
  NANDN U2315 ( .A(n2188), .B(sreg[347]), .Z(n2192) );
  NAND U2316 ( .A(n2190), .B(n2189), .Z(n2191) );
  NAND U2317 ( .A(n2192), .B(n2191), .Z(n2212) );
  XOR U2318 ( .A(n2213), .B(n2212), .Z(c[348]) );
  NANDN U2319 ( .A(n2194), .B(n2193), .Z(n2198) );
  OR U2320 ( .A(n2196), .B(n2195), .Z(n2197) );
  AND U2321 ( .A(n2198), .B(n2197), .Z(n2218) );
  NAND U2322 ( .A(n31), .B(n2199), .Z(n2201) );
  XOR U2323 ( .A(b[3]), .B(a[95]), .Z(n2222) );
  NAND U2324 ( .A(n5811), .B(n2222), .Z(n2200) );
  AND U2325 ( .A(n2201), .B(n2200), .Z(n2230) );
  AND U2326 ( .A(b[3]), .B(a[93]), .Z(n2228) );
  NAND U2327 ( .A(b[0]), .B(a[97]), .Z(n2202) );
  XNOR U2328 ( .A(b[1]), .B(n2202), .Z(n2204) );
  NANDN U2329 ( .A(b[0]), .B(a[96]), .Z(n2203) );
  NAND U2330 ( .A(n2204), .B(n2203), .Z(n2229) );
  XOR U2331 ( .A(n2228), .B(n2229), .Z(n2231) );
  XOR U2332 ( .A(n2230), .B(n2231), .Z(n2217) );
  NANDN U2333 ( .A(n2206), .B(n2205), .Z(n2210) );
  OR U2334 ( .A(n2208), .B(n2207), .Z(n2209) );
  AND U2335 ( .A(n2210), .B(n2209), .Z(n2216) );
  XOR U2336 ( .A(n2217), .B(n2216), .Z(n2219) );
  XOR U2337 ( .A(n2218), .B(n2219), .Z(n2234) );
  XNOR U2338 ( .A(n2234), .B(sreg[349]), .Z(n2236) );
  NANDN U2339 ( .A(n2211), .B(sreg[348]), .Z(n2215) );
  NAND U2340 ( .A(n2213), .B(n2212), .Z(n2214) );
  NAND U2341 ( .A(n2215), .B(n2214), .Z(n2235) );
  XOR U2342 ( .A(n2236), .B(n2235), .Z(c[349]) );
  NANDN U2343 ( .A(n2217), .B(n2216), .Z(n2221) );
  OR U2344 ( .A(n2219), .B(n2218), .Z(n2220) );
  AND U2345 ( .A(n2221), .B(n2220), .Z(n2241) );
  NAND U2346 ( .A(n31), .B(n2222), .Z(n2224) );
  XOR U2347 ( .A(b[3]), .B(a[96]), .Z(n2245) );
  NAND U2348 ( .A(n5811), .B(n2245), .Z(n2223) );
  AND U2349 ( .A(n2224), .B(n2223), .Z(n2253) );
  NAND U2350 ( .A(b[0]), .B(a[98]), .Z(n2225) );
  XNOR U2351 ( .A(b[1]), .B(n2225), .Z(n2227) );
  NANDN U2352 ( .A(b[0]), .B(a[97]), .Z(n2226) );
  NAND U2353 ( .A(n2227), .B(n2226), .Z(n2252) );
  AND U2354 ( .A(b[3]), .B(a[94]), .Z(n2251) );
  XOR U2355 ( .A(n2252), .B(n2251), .Z(n2254) );
  XOR U2356 ( .A(n2253), .B(n2254), .Z(n2240) );
  NANDN U2357 ( .A(n2229), .B(n2228), .Z(n2233) );
  OR U2358 ( .A(n2231), .B(n2230), .Z(n2232) );
  AND U2359 ( .A(n2233), .B(n2232), .Z(n2239) );
  XOR U2360 ( .A(n2240), .B(n2239), .Z(n2242) );
  XOR U2361 ( .A(n2241), .B(n2242), .Z(n2257) );
  XNOR U2362 ( .A(n2257), .B(sreg[350]), .Z(n2259) );
  NANDN U2363 ( .A(n2234), .B(sreg[349]), .Z(n2238) );
  NAND U2364 ( .A(n2236), .B(n2235), .Z(n2237) );
  NAND U2365 ( .A(n2238), .B(n2237), .Z(n2258) );
  XOR U2366 ( .A(n2259), .B(n2258), .Z(c[350]) );
  NANDN U2367 ( .A(n2240), .B(n2239), .Z(n2244) );
  OR U2368 ( .A(n2242), .B(n2241), .Z(n2243) );
  AND U2369 ( .A(n2244), .B(n2243), .Z(n2264) );
  NAND U2370 ( .A(n31), .B(n2245), .Z(n2247) );
  XOR U2371 ( .A(b[3]), .B(a[97]), .Z(n2268) );
  NAND U2372 ( .A(n5811), .B(n2268), .Z(n2246) );
  AND U2373 ( .A(n2247), .B(n2246), .Z(n2276) );
  AND U2374 ( .A(b[3]), .B(a[95]), .Z(n2274) );
  NAND U2375 ( .A(b[0]), .B(a[99]), .Z(n2248) );
  XNOR U2376 ( .A(b[1]), .B(n2248), .Z(n2250) );
  NANDN U2377 ( .A(b[0]), .B(a[98]), .Z(n2249) );
  NAND U2378 ( .A(n2250), .B(n2249), .Z(n2275) );
  XOR U2379 ( .A(n2274), .B(n2275), .Z(n2277) );
  XOR U2380 ( .A(n2276), .B(n2277), .Z(n2263) );
  NANDN U2381 ( .A(n2252), .B(n2251), .Z(n2256) );
  OR U2382 ( .A(n2254), .B(n2253), .Z(n2255) );
  AND U2383 ( .A(n2256), .B(n2255), .Z(n2262) );
  XOR U2384 ( .A(n2263), .B(n2262), .Z(n2265) );
  XOR U2385 ( .A(n2264), .B(n2265), .Z(n2280) );
  XNOR U2386 ( .A(n2280), .B(sreg[351]), .Z(n2282) );
  NANDN U2387 ( .A(n2257), .B(sreg[350]), .Z(n2261) );
  NAND U2388 ( .A(n2259), .B(n2258), .Z(n2260) );
  NAND U2389 ( .A(n2261), .B(n2260), .Z(n2281) );
  XOR U2390 ( .A(n2282), .B(n2281), .Z(c[351]) );
  NANDN U2391 ( .A(n2263), .B(n2262), .Z(n2267) );
  OR U2392 ( .A(n2265), .B(n2264), .Z(n2266) );
  AND U2393 ( .A(n2267), .B(n2266), .Z(n2287) );
  NAND U2394 ( .A(n31), .B(n2268), .Z(n2270) );
  XOR U2395 ( .A(b[3]), .B(a[98]), .Z(n2291) );
  NAND U2396 ( .A(n5811), .B(n2291), .Z(n2269) );
  AND U2397 ( .A(n2270), .B(n2269), .Z(n2299) );
  AND U2398 ( .A(b[3]), .B(a[96]), .Z(n2297) );
  NAND U2399 ( .A(b[0]), .B(a[100]), .Z(n2271) );
  XNOR U2400 ( .A(b[1]), .B(n2271), .Z(n2273) );
  NANDN U2401 ( .A(b[0]), .B(a[99]), .Z(n2272) );
  NAND U2402 ( .A(n2273), .B(n2272), .Z(n2298) );
  XOR U2403 ( .A(n2297), .B(n2298), .Z(n2300) );
  XOR U2404 ( .A(n2299), .B(n2300), .Z(n2286) );
  NANDN U2405 ( .A(n2275), .B(n2274), .Z(n2279) );
  OR U2406 ( .A(n2277), .B(n2276), .Z(n2278) );
  AND U2407 ( .A(n2279), .B(n2278), .Z(n2285) );
  XOR U2408 ( .A(n2286), .B(n2285), .Z(n2288) );
  XOR U2409 ( .A(n2287), .B(n2288), .Z(n2303) );
  XNOR U2410 ( .A(n2303), .B(sreg[352]), .Z(n2305) );
  NANDN U2411 ( .A(n2280), .B(sreg[351]), .Z(n2284) );
  NAND U2412 ( .A(n2282), .B(n2281), .Z(n2283) );
  NAND U2413 ( .A(n2284), .B(n2283), .Z(n2304) );
  XOR U2414 ( .A(n2305), .B(n2304), .Z(c[352]) );
  NANDN U2415 ( .A(n2286), .B(n2285), .Z(n2290) );
  OR U2416 ( .A(n2288), .B(n2287), .Z(n2289) );
  AND U2417 ( .A(n2290), .B(n2289), .Z(n2310) );
  NAND U2418 ( .A(n31), .B(n2291), .Z(n2293) );
  XOR U2419 ( .A(b[3]), .B(a[99]), .Z(n2314) );
  NAND U2420 ( .A(n5811), .B(n2314), .Z(n2292) );
  AND U2421 ( .A(n2293), .B(n2292), .Z(n2322) );
  NAND U2422 ( .A(b[0]), .B(a[101]), .Z(n2294) );
  XNOR U2423 ( .A(b[1]), .B(n2294), .Z(n2296) );
  NANDN U2424 ( .A(b[0]), .B(a[100]), .Z(n2295) );
  NAND U2425 ( .A(n2296), .B(n2295), .Z(n2321) );
  AND U2426 ( .A(b[3]), .B(a[97]), .Z(n2320) );
  XOR U2427 ( .A(n2321), .B(n2320), .Z(n2323) );
  XOR U2428 ( .A(n2322), .B(n2323), .Z(n2309) );
  NANDN U2429 ( .A(n2298), .B(n2297), .Z(n2302) );
  OR U2430 ( .A(n2300), .B(n2299), .Z(n2301) );
  AND U2431 ( .A(n2302), .B(n2301), .Z(n2308) );
  XOR U2432 ( .A(n2309), .B(n2308), .Z(n2311) );
  XOR U2433 ( .A(n2310), .B(n2311), .Z(n2326) );
  XNOR U2434 ( .A(n2326), .B(sreg[353]), .Z(n2328) );
  NANDN U2435 ( .A(n2303), .B(sreg[352]), .Z(n2307) );
  NAND U2436 ( .A(n2305), .B(n2304), .Z(n2306) );
  NAND U2437 ( .A(n2307), .B(n2306), .Z(n2327) );
  XOR U2438 ( .A(n2328), .B(n2327), .Z(c[353]) );
  NANDN U2439 ( .A(n2309), .B(n2308), .Z(n2313) );
  OR U2440 ( .A(n2311), .B(n2310), .Z(n2312) );
  AND U2441 ( .A(n2313), .B(n2312), .Z(n2333) );
  NAND U2442 ( .A(n31), .B(n2314), .Z(n2316) );
  XOR U2443 ( .A(b[3]), .B(a[100]), .Z(n2337) );
  NAND U2444 ( .A(n5811), .B(n2337), .Z(n2315) );
  AND U2445 ( .A(n2316), .B(n2315), .Z(n2345) );
  NAND U2446 ( .A(b[0]), .B(a[102]), .Z(n2317) );
  XNOR U2447 ( .A(b[1]), .B(n2317), .Z(n2319) );
  NANDN U2448 ( .A(b[0]), .B(a[101]), .Z(n2318) );
  NAND U2449 ( .A(n2319), .B(n2318), .Z(n2344) );
  AND U2450 ( .A(b[3]), .B(a[98]), .Z(n2343) );
  XOR U2451 ( .A(n2344), .B(n2343), .Z(n2346) );
  XOR U2452 ( .A(n2345), .B(n2346), .Z(n2332) );
  NANDN U2453 ( .A(n2321), .B(n2320), .Z(n2325) );
  OR U2454 ( .A(n2323), .B(n2322), .Z(n2324) );
  AND U2455 ( .A(n2325), .B(n2324), .Z(n2331) );
  XOR U2456 ( .A(n2332), .B(n2331), .Z(n2334) );
  XOR U2457 ( .A(n2333), .B(n2334), .Z(n2349) );
  XNOR U2458 ( .A(n2349), .B(sreg[354]), .Z(n2351) );
  NANDN U2459 ( .A(n2326), .B(sreg[353]), .Z(n2330) );
  NAND U2460 ( .A(n2328), .B(n2327), .Z(n2329) );
  NAND U2461 ( .A(n2330), .B(n2329), .Z(n2350) );
  XOR U2462 ( .A(n2351), .B(n2350), .Z(c[354]) );
  NANDN U2463 ( .A(n2332), .B(n2331), .Z(n2336) );
  OR U2464 ( .A(n2334), .B(n2333), .Z(n2335) );
  AND U2465 ( .A(n2336), .B(n2335), .Z(n2356) );
  NAND U2466 ( .A(n31), .B(n2337), .Z(n2339) );
  XOR U2467 ( .A(b[3]), .B(a[101]), .Z(n2360) );
  NAND U2468 ( .A(n5811), .B(n2360), .Z(n2338) );
  AND U2469 ( .A(n2339), .B(n2338), .Z(n2368) );
  NAND U2470 ( .A(b[0]), .B(a[103]), .Z(n2340) );
  XNOR U2471 ( .A(b[1]), .B(n2340), .Z(n2342) );
  NANDN U2472 ( .A(b[0]), .B(a[102]), .Z(n2341) );
  NAND U2473 ( .A(n2342), .B(n2341), .Z(n2367) );
  AND U2474 ( .A(b[3]), .B(a[99]), .Z(n2366) );
  XOR U2475 ( .A(n2367), .B(n2366), .Z(n2369) );
  XOR U2476 ( .A(n2368), .B(n2369), .Z(n2355) );
  NANDN U2477 ( .A(n2344), .B(n2343), .Z(n2348) );
  OR U2478 ( .A(n2346), .B(n2345), .Z(n2347) );
  AND U2479 ( .A(n2348), .B(n2347), .Z(n2354) );
  XOR U2480 ( .A(n2355), .B(n2354), .Z(n2357) );
  XOR U2481 ( .A(n2356), .B(n2357), .Z(n2372) );
  XNOR U2482 ( .A(n2372), .B(sreg[355]), .Z(n2374) );
  NANDN U2483 ( .A(n2349), .B(sreg[354]), .Z(n2353) );
  NAND U2484 ( .A(n2351), .B(n2350), .Z(n2352) );
  NAND U2485 ( .A(n2353), .B(n2352), .Z(n2373) );
  XOR U2486 ( .A(n2374), .B(n2373), .Z(c[355]) );
  NANDN U2487 ( .A(n2355), .B(n2354), .Z(n2359) );
  OR U2488 ( .A(n2357), .B(n2356), .Z(n2358) );
  AND U2489 ( .A(n2359), .B(n2358), .Z(n2379) );
  NAND U2490 ( .A(n31), .B(n2360), .Z(n2362) );
  XOR U2491 ( .A(b[3]), .B(a[102]), .Z(n2383) );
  NAND U2492 ( .A(n5811), .B(n2383), .Z(n2361) );
  AND U2493 ( .A(n2362), .B(n2361), .Z(n2391) );
  NAND U2494 ( .A(b[0]), .B(a[104]), .Z(n2363) );
  XNOR U2495 ( .A(b[1]), .B(n2363), .Z(n2365) );
  NANDN U2496 ( .A(b[0]), .B(a[103]), .Z(n2364) );
  NAND U2497 ( .A(n2365), .B(n2364), .Z(n2390) );
  AND U2498 ( .A(b[3]), .B(a[100]), .Z(n2389) );
  XOR U2499 ( .A(n2390), .B(n2389), .Z(n2392) );
  XOR U2500 ( .A(n2391), .B(n2392), .Z(n2378) );
  NANDN U2501 ( .A(n2367), .B(n2366), .Z(n2371) );
  OR U2502 ( .A(n2369), .B(n2368), .Z(n2370) );
  AND U2503 ( .A(n2371), .B(n2370), .Z(n2377) );
  XOR U2504 ( .A(n2378), .B(n2377), .Z(n2380) );
  XOR U2505 ( .A(n2379), .B(n2380), .Z(n2395) );
  XNOR U2506 ( .A(n2395), .B(sreg[356]), .Z(n2397) );
  NANDN U2507 ( .A(n2372), .B(sreg[355]), .Z(n2376) );
  NAND U2508 ( .A(n2374), .B(n2373), .Z(n2375) );
  NAND U2509 ( .A(n2376), .B(n2375), .Z(n2396) );
  XOR U2510 ( .A(n2397), .B(n2396), .Z(c[356]) );
  NANDN U2511 ( .A(n2378), .B(n2377), .Z(n2382) );
  OR U2512 ( .A(n2380), .B(n2379), .Z(n2381) );
  AND U2513 ( .A(n2382), .B(n2381), .Z(n2402) );
  NAND U2514 ( .A(n31), .B(n2383), .Z(n2385) );
  XOR U2515 ( .A(b[3]), .B(a[103]), .Z(n2406) );
  NAND U2516 ( .A(n5811), .B(n2406), .Z(n2384) );
  AND U2517 ( .A(n2385), .B(n2384), .Z(n2414) );
  NAND U2518 ( .A(b[0]), .B(a[105]), .Z(n2386) );
  XNOR U2519 ( .A(b[1]), .B(n2386), .Z(n2388) );
  NANDN U2520 ( .A(b[0]), .B(a[104]), .Z(n2387) );
  NAND U2521 ( .A(n2388), .B(n2387), .Z(n2413) );
  AND U2522 ( .A(b[3]), .B(a[101]), .Z(n2412) );
  XOR U2523 ( .A(n2413), .B(n2412), .Z(n2415) );
  XOR U2524 ( .A(n2414), .B(n2415), .Z(n2401) );
  NANDN U2525 ( .A(n2390), .B(n2389), .Z(n2394) );
  OR U2526 ( .A(n2392), .B(n2391), .Z(n2393) );
  AND U2527 ( .A(n2394), .B(n2393), .Z(n2400) );
  XOR U2528 ( .A(n2401), .B(n2400), .Z(n2403) );
  XOR U2529 ( .A(n2402), .B(n2403), .Z(n2418) );
  XNOR U2530 ( .A(n2418), .B(sreg[357]), .Z(n2420) );
  NANDN U2531 ( .A(n2395), .B(sreg[356]), .Z(n2399) );
  NAND U2532 ( .A(n2397), .B(n2396), .Z(n2398) );
  NAND U2533 ( .A(n2399), .B(n2398), .Z(n2419) );
  XOR U2534 ( .A(n2420), .B(n2419), .Z(c[357]) );
  NANDN U2535 ( .A(n2401), .B(n2400), .Z(n2405) );
  OR U2536 ( .A(n2403), .B(n2402), .Z(n2404) );
  AND U2537 ( .A(n2405), .B(n2404), .Z(n2425) );
  NAND U2538 ( .A(n31), .B(n2406), .Z(n2408) );
  XOR U2539 ( .A(b[3]), .B(a[104]), .Z(n2429) );
  NAND U2540 ( .A(n5811), .B(n2429), .Z(n2407) );
  AND U2541 ( .A(n2408), .B(n2407), .Z(n2437) );
  NAND U2542 ( .A(b[0]), .B(a[106]), .Z(n2409) );
  XNOR U2543 ( .A(b[1]), .B(n2409), .Z(n2411) );
  NANDN U2544 ( .A(b[0]), .B(a[105]), .Z(n2410) );
  NAND U2545 ( .A(n2411), .B(n2410), .Z(n2436) );
  AND U2546 ( .A(b[3]), .B(a[102]), .Z(n2435) );
  XOR U2547 ( .A(n2436), .B(n2435), .Z(n2438) );
  XOR U2548 ( .A(n2437), .B(n2438), .Z(n2424) );
  NANDN U2549 ( .A(n2413), .B(n2412), .Z(n2417) );
  OR U2550 ( .A(n2415), .B(n2414), .Z(n2416) );
  AND U2551 ( .A(n2417), .B(n2416), .Z(n2423) );
  XOR U2552 ( .A(n2424), .B(n2423), .Z(n2426) );
  XOR U2553 ( .A(n2425), .B(n2426), .Z(n2441) );
  XNOR U2554 ( .A(n2441), .B(sreg[358]), .Z(n2443) );
  NANDN U2555 ( .A(n2418), .B(sreg[357]), .Z(n2422) );
  NAND U2556 ( .A(n2420), .B(n2419), .Z(n2421) );
  NAND U2557 ( .A(n2422), .B(n2421), .Z(n2442) );
  XOR U2558 ( .A(n2443), .B(n2442), .Z(c[358]) );
  NANDN U2559 ( .A(n2424), .B(n2423), .Z(n2428) );
  OR U2560 ( .A(n2426), .B(n2425), .Z(n2427) );
  AND U2561 ( .A(n2428), .B(n2427), .Z(n2448) );
  NAND U2562 ( .A(n31), .B(n2429), .Z(n2431) );
  XOR U2563 ( .A(b[3]), .B(a[105]), .Z(n2452) );
  NAND U2564 ( .A(n5811), .B(n2452), .Z(n2430) );
  AND U2565 ( .A(n2431), .B(n2430), .Z(n2460) );
  NAND U2566 ( .A(b[0]), .B(a[107]), .Z(n2432) );
  XNOR U2567 ( .A(b[1]), .B(n2432), .Z(n2434) );
  NANDN U2568 ( .A(b[0]), .B(a[106]), .Z(n2433) );
  NAND U2569 ( .A(n2434), .B(n2433), .Z(n2459) );
  AND U2570 ( .A(b[3]), .B(a[103]), .Z(n2458) );
  XOR U2571 ( .A(n2459), .B(n2458), .Z(n2461) );
  XOR U2572 ( .A(n2460), .B(n2461), .Z(n2447) );
  NANDN U2573 ( .A(n2436), .B(n2435), .Z(n2440) );
  OR U2574 ( .A(n2438), .B(n2437), .Z(n2439) );
  AND U2575 ( .A(n2440), .B(n2439), .Z(n2446) );
  XOR U2576 ( .A(n2447), .B(n2446), .Z(n2449) );
  XOR U2577 ( .A(n2448), .B(n2449), .Z(n2464) );
  XNOR U2578 ( .A(n2464), .B(sreg[359]), .Z(n2466) );
  NANDN U2579 ( .A(n2441), .B(sreg[358]), .Z(n2445) );
  NAND U2580 ( .A(n2443), .B(n2442), .Z(n2444) );
  NAND U2581 ( .A(n2445), .B(n2444), .Z(n2465) );
  XOR U2582 ( .A(n2466), .B(n2465), .Z(c[359]) );
  NANDN U2583 ( .A(n2447), .B(n2446), .Z(n2451) );
  OR U2584 ( .A(n2449), .B(n2448), .Z(n2450) );
  AND U2585 ( .A(n2451), .B(n2450), .Z(n2471) );
  NAND U2586 ( .A(n31), .B(n2452), .Z(n2454) );
  XOR U2587 ( .A(b[3]), .B(a[106]), .Z(n2475) );
  NAND U2588 ( .A(n5811), .B(n2475), .Z(n2453) );
  AND U2589 ( .A(n2454), .B(n2453), .Z(n2483) );
  AND U2590 ( .A(b[3]), .B(a[104]), .Z(n2481) );
  NAND U2591 ( .A(b[0]), .B(a[108]), .Z(n2455) );
  XNOR U2592 ( .A(b[1]), .B(n2455), .Z(n2457) );
  NANDN U2593 ( .A(b[0]), .B(a[107]), .Z(n2456) );
  NAND U2594 ( .A(n2457), .B(n2456), .Z(n2482) );
  XOR U2595 ( .A(n2481), .B(n2482), .Z(n2484) );
  XOR U2596 ( .A(n2483), .B(n2484), .Z(n2470) );
  NANDN U2597 ( .A(n2459), .B(n2458), .Z(n2463) );
  OR U2598 ( .A(n2461), .B(n2460), .Z(n2462) );
  AND U2599 ( .A(n2463), .B(n2462), .Z(n2469) );
  XOR U2600 ( .A(n2470), .B(n2469), .Z(n2472) );
  XOR U2601 ( .A(n2471), .B(n2472), .Z(n2487) );
  XNOR U2602 ( .A(n2487), .B(sreg[360]), .Z(n2489) );
  NANDN U2603 ( .A(n2464), .B(sreg[359]), .Z(n2468) );
  NAND U2604 ( .A(n2466), .B(n2465), .Z(n2467) );
  NAND U2605 ( .A(n2468), .B(n2467), .Z(n2488) );
  XOR U2606 ( .A(n2489), .B(n2488), .Z(c[360]) );
  NANDN U2607 ( .A(n2470), .B(n2469), .Z(n2474) );
  OR U2608 ( .A(n2472), .B(n2471), .Z(n2473) );
  AND U2609 ( .A(n2474), .B(n2473), .Z(n2494) );
  NAND U2610 ( .A(n31), .B(n2475), .Z(n2477) );
  XOR U2611 ( .A(b[3]), .B(a[107]), .Z(n2498) );
  NAND U2612 ( .A(n5811), .B(n2498), .Z(n2476) );
  AND U2613 ( .A(n2477), .B(n2476), .Z(n2506) );
  NAND U2614 ( .A(b[0]), .B(a[109]), .Z(n2478) );
  XNOR U2615 ( .A(b[1]), .B(n2478), .Z(n2480) );
  NANDN U2616 ( .A(b[0]), .B(a[108]), .Z(n2479) );
  NAND U2617 ( .A(n2480), .B(n2479), .Z(n2505) );
  AND U2618 ( .A(b[3]), .B(a[105]), .Z(n2504) );
  XOR U2619 ( .A(n2505), .B(n2504), .Z(n2507) );
  XOR U2620 ( .A(n2506), .B(n2507), .Z(n2493) );
  NANDN U2621 ( .A(n2482), .B(n2481), .Z(n2486) );
  OR U2622 ( .A(n2484), .B(n2483), .Z(n2485) );
  AND U2623 ( .A(n2486), .B(n2485), .Z(n2492) );
  XOR U2624 ( .A(n2493), .B(n2492), .Z(n2495) );
  XOR U2625 ( .A(n2494), .B(n2495), .Z(n2510) );
  XNOR U2626 ( .A(n2510), .B(sreg[361]), .Z(n2512) );
  NANDN U2627 ( .A(n2487), .B(sreg[360]), .Z(n2491) );
  NAND U2628 ( .A(n2489), .B(n2488), .Z(n2490) );
  NAND U2629 ( .A(n2491), .B(n2490), .Z(n2511) );
  XOR U2630 ( .A(n2512), .B(n2511), .Z(c[361]) );
  NANDN U2631 ( .A(n2493), .B(n2492), .Z(n2497) );
  OR U2632 ( .A(n2495), .B(n2494), .Z(n2496) );
  AND U2633 ( .A(n2497), .B(n2496), .Z(n2517) );
  NAND U2634 ( .A(n31), .B(n2498), .Z(n2500) );
  XOR U2635 ( .A(b[3]), .B(a[108]), .Z(n2521) );
  NAND U2636 ( .A(n5811), .B(n2521), .Z(n2499) );
  AND U2637 ( .A(n2500), .B(n2499), .Z(n2529) );
  NAND U2638 ( .A(b[0]), .B(a[110]), .Z(n2501) );
  XNOR U2639 ( .A(b[1]), .B(n2501), .Z(n2503) );
  NANDN U2640 ( .A(b[0]), .B(a[109]), .Z(n2502) );
  NAND U2641 ( .A(n2503), .B(n2502), .Z(n2528) );
  AND U2642 ( .A(b[3]), .B(a[106]), .Z(n2527) );
  XOR U2643 ( .A(n2528), .B(n2527), .Z(n2530) );
  XOR U2644 ( .A(n2529), .B(n2530), .Z(n2516) );
  NANDN U2645 ( .A(n2505), .B(n2504), .Z(n2509) );
  OR U2646 ( .A(n2507), .B(n2506), .Z(n2508) );
  AND U2647 ( .A(n2509), .B(n2508), .Z(n2515) );
  XOR U2648 ( .A(n2516), .B(n2515), .Z(n2518) );
  XOR U2649 ( .A(n2517), .B(n2518), .Z(n2533) );
  XNOR U2650 ( .A(n2533), .B(sreg[362]), .Z(n2535) );
  NANDN U2651 ( .A(n2510), .B(sreg[361]), .Z(n2514) );
  NAND U2652 ( .A(n2512), .B(n2511), .Z(n2513) );
  NAND U2653 ( .A(n2514), .B(n2513), .Z(n2534) );
  XOR U2654 ( .A(n2535), .B(n2534), .Z(c[362]) );
  NANDN U2655 ( .A(n2516), .B(n2515), .Z(n2520) );
  OR U2656 ( .A(n2518), .B(n2517), .Z(n2519) );
  AND U2657 ( .A(n2520), .B(n2519), .Z(n2540) );
  NAND U2658 ( .A(n31), .B(n2521), .Z(n2523) );
  XOR U2659 ( .A(b[3]), .B(a[109]), .Z(n2544) );
  NAND U2660 ( .A(n5811), .B(n2544), .Z(n2522) );
  AND U2661 ( .A(n2523), .B(n2522), .Z(n2552) );
  NAND U2662 ( .A(b[0]), .B(a[111]), .Z(n2524) );
  XNOR U2663 ( .A(b[1]), .B(n2524), .Z(n2526) );
  NANDN U2664 ( .A(b[0]), .B(a[110]), .Z(n2525) );
  NAND U2665 ( .A(n2526), .B(n2525), .Z(n2551) );
  AND U2666 ( .A(b[3]), .B(a[107]), .Z(n2550) );
  XOR U2667 ( .A(n2551), .B(n2550), .Z(n2553) );
  XOR U2668 ( .A(n2552), .B(n2553), .Z(n2539) );
  NANDN U2669 ( .A(n2528), .B(n2527), .Z(n2532) );
  OR U2670 ( .A(n2530), .B(n2529), .Z(n2531) );
  AND U2671 ( .A(n2532), .B(n2531), .Z(n2538) );
  XOR U2672 ( .A(n2539), .B(n2538), .Z(n2541) );
  XOR U2673 ( .A(n2540), .B(n2541), .Z(n2556) );
  XNOR U2674 ( .A(n2556), .B(sreg[363]), .Z(n2558) );
  NANDN U2675 ( .A(n2533), .B(sreg[362]), .Z(n2537) );
  NAND U2676 ( .A(n2535), .B(n2534), .Z(n2536) );
  NAND U2677 ( .A(n2537), .B(n2536), .Z(n2557) );
  XOR U2678 ( .A(n2558), .B(n2557), .Z(c[363]) );
  NANDN U2679 ( .A(n2539), .B(n2538), .Z(n2543) );
  OR U2680 ( .A(n2541), .B(n2540), .Z(n2542) );
  AND U2681 ( .A(n2543), .B(n2542), .Z(n2563) );
  NAND U2682 ( .A(n31), .B(n2544), .Z(n2546) );
  XOR U2683 ( .A(b[3]), .B(a[110]), .Z(n2567) );
  NAND U2684 ( .A(n5811), .B(n2567), .Z(n2545) );
  AND U2685 ( .A(n2546), .B(n2545), .Z(n2575) );
  NAND U2686 ( .A(b[0]), .B(a[112]), .Z(n2547) );
  XNOR U2687 ( .A(b[1]), .B(n2547), .Z(n2549) );
  NANDN U2688 ( .A(b[0]), .B(a[111]), .Z(n2548) );
  NAND U2689 ( .A(n2549), .B(n2548), .Z(n2574) );
  AND U2690 ( .A(b[3]), .B(a[108]), .Z(n2573) );
  XOR U2691 ( .A(n2574), .B(n2573), .Z(n2576) );
  XOR U2692 ( .A(n2575), .B(n2576), .Z(n2562) );
  NANDN U2693 ( .A(n2551), .B(n2550), .Z(n2555) );
  OR U2694 ( .A(n2553), .B(n2552), .Z(n2554) );
  AND U2695 ( .A(n2555), .B(n2554), .Z(n2561) );
  XOR U2696 ( .A(n2562), .B(n2561), .Z(n2564) );
  XOR U2697 ( .A(n2563), .B(n2564), .Z(n2579) );
  XNOR U2698 ( .A(n2579), .B(sreg[364]), .Z(n2581) );
  NANDN U2699 ( .A(n2556), .B(sreg[363]), .Z(n2560) );
  NAND U2700 ( .A(n2558), .B(n2557), .Z(n2559) );
  NAND U2701 ( .A(n2560), .B(n2559), .Z(n2580) );
  XOR U2702 ( .A(n2581), .B(n2580), .Z(c[364]) );
  NANDN U2703 ( .A(n2562), .B(n2561), .Z(n2566) );
  OR U2704 ( .A(n2564), .B(n2563), .Z(n2565) );
  AND U2705 ( .A(n2566), .B(n2565), .Z(n2586) );
  NAND U2706 ( .A(n31), .B(n2567), .Z(n2569) );
  XOR U2707 ( .A(b[3]), .B(a[111]), .Z(n2590) );
  NAND U2708 ( .A(n5811), .B(n2590), .Z(n2568) );
  AND U2709 ( .A(n2569), .B(n2568), .Z(n2598) );
  NAND U2710 ( .A(b[0]), .B(a[113]), .Z(n2570) );
  XNOR U2711 ( .A(b[1]), .B(n2570), .Z(n2572) );
  NANDN U2712 ( .A(b[0]), .B(a[112]), .Z(n2571) );
  NAND U2713 ( .A(n2572), .B(n2571), .Z(n2597) );
  AND U2714 ( .A(b[3]), .B(a[109]), .Z(n2596) );
  XOR U2715 ( .A(n2597), .B(n2596), .Z(n2599) );
  XOR U2716 ( .A(n2598), .B(n2599), .Z(n2585) );
  NANDN U2717 ( .A(n2574), .B(n2573), .Z(n2578) );
  OR U2718 ( .A(n2576), .B(n2575), .Z(n2577) );
  AND U2719 ( .A(n2578), .B(n2577), .Z(n2584) );
  XOR U2720 ( .A(n2585), .B(n2584), .Z(n2587) );
  XOR U2721 ( .A(n2586), .B(n2587), .Z(n2602) );
  XNOR U2722 ( .A(n2602), .B(sreg[365]), .Z(n2604) );
  NANDN U2723 ( .A(n2579), .B(sreg[364]), .Z(n2583) );
  NAND U2724 ( .A(n2581), .B(n2580), .Z(n2582) );
  NAND U2725 ( .A(n2583), .B(n2582), .Z(n2603) );
  XOR U2726 ( .A(n2604), .B(n2603), .Z(c[365]) );
  NANDN U2727 ( .A(n2585), .B(n2584), .Z(n2589) );
  OR U2728 ( .A(n2587), .B(n2586), .Z(n2588) );
  AND U2729 ( .A(n2589), .B(n2588), .Z(n2609) );
  NAND U2730 ( .A(n31), .B(n2590), .Z(n2592) );
  XOR U2731 ( .A(b[3]), .B(a[112]), .Z(n2613) );
  NAND U2732 ( .A(n5811), .B(n2613), .Z(n2591) );
  AND U2733 ( .A(n2592), .B(n2591), .Z(n2621) );
  NAND U2734 ( .A(b[0]), .B(a[114]), .Z(n2593) );
  XNOR U2735 ( .A(b[1]), .B(n2593), .Z(n2595) );
  NANDN U2736 ( .A(b[0]), .B(a[113]), .Z(n2594) );
  NAND U2737 ( .A(n2595), .B(n2594), .Z(n2620) );
  AND U2738 ( .A(b[3]), .B(a[110]), .Z(n2619) );
  XOR U2739 ( .A(n2620), .B(n2619), .Z(n2622) );
  XOR U2740 ( .A(n2621), .B(n2622), .Z(n2608) );
  NANDN U2741 ( .A(n2597), .B(n2596), .Z(n2601) );
  OR U2742 ( .A(n2599), .B(n2598), .Z(n2600) );
  AND U2743 ( .A(n2601), .B(n2600), .Z(n2607) );
  XOR U2744 ( .A(n2608), .B(n2607), .Z(n2610) );
  XOR U2745 ( .A(n2609), .B(n2610), .Z(n2625) );
  XNOR U2746 ( .A(n2625), .B(sreg[366]), .Z(n2627) );
  NANDN U2747 ( .A(n2602), .B(sreg[365]), .Z(n2606) );
  NAND U2748 ( .A(n2604), .B(n2603), .Z(n2605) );
  NAND U2749 ( .A(n2606), .B(n2605), .Z(n2626) );
  XOR U2750 ( .A(n2627), .B(n2626), .Z(c[366]) );
  NANDN U2751 ( .A(n2608), .B(n2607), .Z(n2612) );
  OR U2752 ( .A(n2610), .B(n2609), .Z(n2611) );
  AND U2753 ( .A(n2612), .B(n2611), .Z(n2632) );
  NAND U2754 ( .A(n31), .B(n2613), .Z(n2615) );
  XOR U2755 ( .A(b[3]), .B(a[113]), .Z(n2636) );
  NAND U2756 ( .A(n5811), .B(n2636), .Z(n2614) );
  AND U2757 ( .A(n2615), .B(n2614), .Z(n2644) );
  NAND U2758 ( .A(b[0]), .B(a[115]), .Z(n2616) );
  XNOR U2759 ( .A(b[1]), .B(n2616), .Z(n2618) );
  NANDN U2760 ( .A(b[0]), .B(a[114]), .Z(n2617) );
  NAND U2761 ( .A(n2618), .B(n2617), .Z(n2643) );
  AND U2762 ( .A(b[3]), .B(a[111]), .Z(n2642) );
  XOR U2763 ( .A(n2643), .B(n2642), .Z(n2645) );
  XOR U2764 ( .A(n2644), .B(n2645), .Z(n2631) );
  NANDN U2765 ( .A(n2620), .B(n2619), .Z(n2624) );
  OR U2766 ( .A(n2622), .B(n2621), .Z(n2623) );
  AND U2767 ( .A(n2624), .B(n2623), .Z(n2630) );
  XOR U2768 ( .A(n2631), .B(n2630), .Z(n2633) );
  XOR U2769 ( .A(n2632), .B(n2633), .Z(n2648) );
  XNOR U2770 ( .A(n2648), .B(sreg[367]), .Z(n2650) );
  NANDN U2771 ( .A(n2625), .B(sreg[366]), .Z(n2629) );
  NAND U2772 ( .A(n2627), .B(n2626), .Z(n2628) );
  NAND U2773 ( .A(n2629), .B(n2628), .Z(n2649) );
  XOR U2774 ( .A(n2650), .B(n2649), .Z(c[367]) );
  NANDN U2775 ( .A(n2631), .B(n2630), .Z(n2635) );
  OR U2776 ( .A(n2633), .B(n2632), .Z(n2634) );
  AND U2777 ( .A(n2635), .B(n2634), .Z(n2655) );
  NAND U2778 ( .A(n31), .B(n2636), .Z(n2638) );
  XOR U2779 ( .A(b[3]), .B(a[114]), .Z(n2659) );
  NAND U2780 ( .A(n5811), .B(n2659), .Z(n2637) );
  AND U2781 ( .A(n2638), .B(n2637), .Z(n2667) );
  NAND U2782 ( .A(b[0]), .B(a[116]), .Z(n2639) );
  XNOR U2783 ( .A(b[1]), .B(n2639), .Z(n2641) );
  NANDN U2784 ( .A(b[0]), .B(a[115]), .Z(n2640) );
  NAND U2785 ( .A(n2641), .B(n2640), .Z(n2666) );
  AND U2786 ( .A(b[3]), .B(a[112]), .Z(n2665) );
  XOR U2787 ( .A(n2666), .B(n2665), .Z(n2668) );
  XOR U2788 ( .A(n2667), .B(n2668), .Z(n2654) );
  NANDN U2789 ( .A(n2643), .B(n2642), .Z(n2647) );
  OR U2790 ( .A(n2645), .B(n2644), .Z(n2646) );
  AND U2791 ( .A(n2647), .B(n2646), .Z(n2653) );
  XOR U2792 ( .A(n2654), .B(n2653), .Z(n2656) );
  XOR U2793 ( .A(n2655), .B(n2656), .Z(n2671) );
  XNOR U2794 ( .A(n2671), .B(sreg[368]), .Z(n2673) );
  NANDN U2795 ( .A(n2648), .B(sreg[367]), .Z(n2652) );
  NAND U2796 ( .A(n2650), .B(n2649), .Z(n2651) );
  NAND U2797 ( .A(n2652), .B(n2651), .Z(n2672) );
  XOR U2798 ( .A(n2673), .B(n2672), .Z(c[368]) );
  NANDN U2799 ( .A(n2654), .B(n2653), .Z(n2658) );
  OR U2800 ( .A(n2656), .B(n2655), .Z(n2657) );
  AND U2801 ( .A(n2658), .B(n2657), .Z(n2678) );
  NAND U2802 ( .A(n31), .B(n2659), .Z(n2661) );
  XOR U2803 ( .A(b[3]), .B(a[115]), .Z(n2682) );
  NAND U2804 ( .A(n5811), .B(n2682), .Z(n2660) );
  AND U2805 ( .A(n2661), .B(n2660), .Z(n2690) );
  AND U2806 ( .A(b[3]), .B(a[113]), .Z(n2688) );
  NAND U2807 ( .A(b[0]), .B(a[117]), .Z(n2662) );
  XNOR U2808 ( .A(b[1]), .B(n2662), .Z(n2664) );
  NANDN U2809 ( .A(b[0]), .B(a[116]), .Z(n2663) );
  NAND U2810 ( .A(n2664), .B(n2663), .Z(n2689) );
  XOR U2811 ( .A(n2688), .B(n2689), .Z(n2691) );
  XOR U2812 ( .A(n2690), .B(n2691), .Z(n2677) );
  NANDN U2813 ( .A(n2666), .B(n2665), .Z(n2670) );
  OR U2814 ( .A(n2668), .B(n2667), .Z(n2669) );
  AND U2815 ( .A(n2670), .B(n2669), .Z(n2676) );
  XOR U2816 ( .A(n2677), .B(n2676), .Z(n2679) );
  XOR U2817 ( .A(n2678), .B(n2679), .Z(n2694) );
  XNOR U2818 ( .A(n2694), .B(sreg[369]), .Z(n2696) );
  NANDN U2819 ( .A(n2671), .B(sreg[368]), .Z(n2675) );
  NAND U2820 ( .A(n2673), .B(n2672), .Z(n2674) );
  NAND U2821 ( .A(n2675), .B(n2674), .Z(n2695) );
  XOR U2822 ( .A(n2696), .B(n2695), .Z(c[369]) );
  NANDN U2823 ( .A(n2677), .B(n2676), .Z(n2681) );
  OR U2824 ( .A(n2679), .B(n2678), .Z(n2680) );
  AND U2825 ( .A(n2681), .B(n2680), .Z(n2701) );
  NAND U2826 ( .A(n31), .B(n2682), .Z(n2684) );
  XOR U2827 ( .A(b[3]), .B(a[116]), .Z(n2705) );
  NAND U2828 ( .A(n5811), .B(n2705), .Z(n2683) );
  AND U2829 ( .A(n2684), .B(n2683), .Z(n2713) );
  NAND U2830 ( .A(b[0]), .B(a[118]), .Z(n2685) );
  XNOR U2831 ( .A(b[1]), .B(n2685), .Z(n2687) );
  NANDN U2832 ( .A(b[0]), .B(a[117]), .Z(n2686) );
  NAND U2833 ( .A(n2687), .B(n2686), .Z(n2712) );
  AND U2834 ( .A(b[3]), .B(a[114]), .Z(n2711) );
  XOR U2835 ( .A(n2712), .B(n2711), .Z(n2714) );
  XOR U2836 ( .A(n2713), .B(n2714), .Z(n2700) );
  NANDN U2837 ( .A(n2689), .B(n2688), .Z(n2693) );
  OR U2838 ( .A(n2691), .B(n2690), .Z(n2692) );
  AND U2839 ( .A(n2693), .B(n2692), .Z(n2699) );
  XOR U2840 ( .A(n2700), .B(n2699), .Z(n2702) );
  XOR U2841 ( .A(n2701), .B(n2702), .Z(n2717) );
  XNOR U2842 ( .A(n2717), .B(sreg[370]), .Z(n2719) );
  NANDN U2843 ( .A(n2694), .B(sreg[369]), .Z(n2698) );
  NAND U2844 ( .A(n2696), .B(n2695), .Z(n2697) );
  NAND U2845 ( .A(n2698), .B(n2697), .Z(n2718) );
  XOR U2846 ( .A(n2719), .B(n2718), .Z(c[370]) );
  NANDN U2847 ( .A(n2700), .B(n2699), .Z(n2704) );
  OR U2848 ( .A(n2702), .B(n2701), .Z(n2703) );
  AND U2849 ( .A(n2704), .B(n2703), .Z(n2724) );
  NAND U2850 ( .A(n31), .B(n2705), .Z(n2707) );
  XOR U2851 ( .A(b[3]), .B(a[117]), .Z(n2728) );
  NAND U2852 ( .A(n5811), .B(n2728), .Z(n2706) );
  AND U2853 ( .A(n2707), .B(n2706), .Z(n2736) );
  NAND U2854 ( .A(b[0]), .B(a[119]), .Z(n2708) );
  XNOR U2855 ( .A(b[1]), .B(n2708), .Z(n2710) );
  NANDN U2856 ( .A(b[0]), .B(a[118]), .Z(n2709) );
  NAND U2857 ( .A(n2710), .B(n2709), .Z(n2735) );
  AND U2858 ( .A(b[3]), .B(a[115]), .Z(n2734) );
  XOR U2859 ( .A(n2735), .B(n2734), .Z(n2737) );
  XOR U2860 ( .A(n2736), .B(n2737), .Z(n2723) );
  NANDN U2861 ( .A(n2712), .B(n2711), .Z(n2716) );
  OR U2862 ( .A(n2714), .B(n2713), .Z(n2715) );
  AND U2863 ( .A(n2716), .B(n2715), .Z(n2722) );
  XOR U2864 ( .A(n2723), .B(n2722), .Z(n2725) );
  XOR U2865 ( .A(n2724), .B(n2725), .Z(n2740) );
  XNOR U2866 ( .A(n2740), .B(sreg[371]), .Z(n2742) );
  NANDN U2867 ( .A(n2717), .B(sreg[370]), .Z(n2721) );
  NAND U2868 ( .A(n2719), .B(n2718), .Z(n2720) );
  NAND U2869 ( .A(n2721), .B(n2720), .Z(n2741) );
  XOR U2870 ( .A(n2742), .B(n2741), .Z(c[371]) );
  NANDN U2871 ( .A(n2723), .B(n2722), .Z(n2727) );
  OR U2872 ( .A(n2725), .B(n2724), .Z(n2726) );
  AND U2873 ( .A(n2727), .B(n2726), .Z(n2747) );
  NAND U2874 ( .A(n31), .B(n2728), .Z(n2730) );
  XOR U2875 ( .A(b[3]), .B(a[118]), .Z(n2751) );
  NAND U2876 ( .A(n5811), .B(n2751), .Z(n2729) );
  AND U2877 ( .A(n2730), .B(n2729), .Z(n2759) );
  AND U2878 ( .A(b[3]), .B(a[116]), .Z(n2757) );
  NAND U2879 ( .A(b[0]), .B(a[120]), .Z(n2731) );
  XNOR U2880 ( .A(b[1]), .B(n2731), .Z(n2733) );
  NANDN U2881 ( .A(b[0]), .B(a[119]), .Z(n2732) );
  NAND U2882 ( .A(n2733), .B(n2732), .Z(n2758) );
  XOR U2883 ( .A(n2757), .B(n2758), .Z(n2760) );
  XOR U2884 ( .A(n2759), .B(n2760), .Z(n2746) );
  NANDN U2885 ( .A(n2735), .B(n2734), .Z(n2739) );
  OR U2886 ( .A(n2737), .B(n2736), .Z(n2738) );
  AND U2887 ( .A(n2739), .B(n2738), .Z(n2745) );
  XOR U2888 ( .A(n2746), .B(n2745), .Z(n2748) );
  XOR U2889 ( .A(n2747), .B(n2748), .Z(n2763) );
  XNOR U2890 ( .A(n2763), .B(sreg[372]), .Z(n2765) );
  NANDN U2891 ( .A(n2740), .B(sreg[371]), .Z(n2744) );
  NAND U2892 ( .A(n2742), .B(n2741), .Z(n2743) );
  NAND U2893 ( .A(n2744), .B(n2743), .Z(n2764) );
  XOR U2894 ( .A(n2765), .B(n2764), .Z(c[372]) );
  NANDN U2895 ( .A(n2746), .B(n2745), .Z(n2750) );
  OR U2896 ( .A(n2748), .B(n2747), .Z(n2749) );
  AND U2897 ( .A(n2750), .B(n2749), .Z(n2770) );
  NAND U2898 ( .A(n31), .B(n2751), .Z(n2753) );
  XOR U2899 ( .A(b[3]), .B(a[119]), .Z(n2774) );
  NAND U2900 ( .A(n5811), .B(n2774), .Z(n2752) );
  AND U2901 ( .A(n2753), .B(n2752), .Z(n2782) );
  AND U2902 ( .A(b[0]), .B(a[121]), .Z(n2754) );
  XOR U2903 ( .A(b[1]), .B(n2754), .Z(n2756) );
  NANDN U2904 ( .A(b[0]), .B(a[120]), .Z(n2755) );
  AND U2905 ( .A(n2756), .B(n2755), .Z(n2780) );
  NAND U2906 ( .A(b[3]), .B(a[117]), .Z(n2781) );
  XOR U2907 ( .A(n2780), .B(n2781), .Z(n2783) );
  XOR U2908 ( .A(n2782), .B(n2783), .Z(n2769) );
  NANDN U2909 ( .A(n2758), .B(n2757), .Z(n2762) );
  OR U2910 ( .A(n2760), .B(n2759), .Z(n2761) );
  AND U2911 ( .A(n2762), .B(n2761), .Z(n2768) );
  XOR U2912 ( .A(n2769), .B(n2768), .Z(n2771) );
  XOR U2913 ( .A(n2770), .B(n2771), .Z(n2786) );
  XNOR U2914 ( .A(n2786), .B(sreg[373]), .Z(n2788) );
  NANDN U2915 ( .A(n2763), .B(sreg[372]), .Z(n2767) );
  NAND U2916 ( .A(n2765), .B(n2764), .Z(n2766) );
  NAND U2917 ( .A(n2767), .B(n2766), .Z(n2787) );
  XOR U2918 ( .A(n2788), .B(n2787), .Z(c[373]) );
  NANDN U2919 ( .A(n2769), .B(n2768), .Z(n2773) );
  OR U2920 ( .A(n2771), .B(n2770), .Z(n2772) );
  AND U2921 ( .A(n2773), .B(n2772), .Z(n2793) );
  NAND U2922 ( .A(n31), .B(n2774), .Z(n2776) );
  XOR U2923 ( .A(b[3]), .B(a[120]), .Z(n2797) );
  NAND U2924 ( .A(n5811), .B(n2797), .Z(n2775) );
  AND U2925 ( .A(n2776), .B(n2775), .Z(n2805) );
  NAND U2926 ( .A(b[0]), .B(a[122]), .Z(n2777) );
  XNOR U2927 ( .A(b[1]), .B(n2777), .Z(n2779) );
  NANDN U2928 ( .A(b[0]), .B(a[121]), .Z(n2778) );
  NAND U2929 ( .A(n2779), .B(n2778), .Z(n2804) );
  AND U2930 ( .A(b[3]), .B(a[118]), .Z(n2803) );
  XOR U2931 ( .A(n2804), .B(n2803), .Z(n2806) );
  XOR U2932 ( .A(n2805), .B(n2806), .Z(n2792) );
  NANDN U2933 ( .A(n2781), .B(n2780), .Z(n2785) );
  OR U2934 ( .A(n2783), .B(n2782), .Z(n2784) );
  AND U2935 ( .A(n2785), .B(n2784), .Z(n2791) );
  XOR U2936 ( .A(n2792), .B(n2791), .Z(n2794) );
  XOR U2937 ( .A(n2793), .B(n2794), .Z(n2809) );
  XNOR U2938 ( .A(n2809), .B(sreg[374]), .Z(n2811) );
  NANDN U2939 ( .A(n2786), .B(sreg[373]), .Z(n2790) );
  NAND U2940 ( .A(n2788), .B(n2787), .Z(n2789) );
  NAND U2941 ( .A(n2790), .B(n2789), .Z(n2810) );
  XOR U2942 ( .A(n2811), .B(n2810), .Z(c[374]) );
  NANDN U2943 ( .A(n2792), .B(n2791), .Z(n2796) );
  OR U2944 ( .A(n2794), .B(n2793), .Z(n2795) );
  AND U2945 ( .A(n2796), .B(n2795), .Z(n2816) );
  NAND U2946 ( .A(n31), .B(n2797), .Z(n2799) );
  XOR U2947 ( .A(b[3]), .B(a[121]), .Z(n2820) );
  NAND U2948 ( .A(n5811), .B(n2820), .Z(n2798) );
  AND U2949 ( .A(n2799), .B(n2798), .Z(n2828) );
  AND U2950 ( .A(b[3]), .B(a[119]), .Z(n2826) );
  NAND U2951 ( .A(b[0]), .B(a[123]), .Z(n2800) );
  XNOR U2952 ( .A(b[1]), .B(n2800), .Z(n2802) );
  NANDN U2953 ( .A(b[0]), .B(a[122]), .Z(n2801) );
  NAND U2954 ( .A(n2802), .B(n2801), .Z(n2827) );
  XOR U2955 ( .A(n2826), .B(n2827), .Z(n2829) );
  XOR U2956 ( .A(n2828), .B(n2829), .Z(n2815) );
  NANDN U2957 ( .A(n2804), .B(n2803), .Z(n2808) );
  OR U2958 ( .A(n2806), .B(n2805), .Z(n2807) );
  AND U2959 ( .A(n2808), .B(n2807), .Z(n2814) );
  XOR U2960 ( .A(n2815), .B(n2814), .Z(n2817) );
  XOR U2961 ( .A(n2816), .B(n2817), .Z(n2832) );
  XNOR U2962 ( .A(n2832), .B(sreg[375]), .Z(n2834) );
  NANDN U2963 ( .A(n2809), .B(sreg[374]), .Z(n2813) );
  NAND U2964 ( .A(n2811), .B(n2810), .Z(n2812) );
  NAND U2965 ( .A(n2813), .B(n2812), .Z(n2833) );
  XOR U2966 ( .A(n2834), .B(n2833), .Z(c[375]) );
  NANDN U2967 ( .A(n2815), .B(n2814), .Z(n2819) );
  OR U2968 ( .A(n2817), .B(n2816), .Z(n2818) );
  AND U2969 ( .A(n2819), .B(n2818), .Z(n2839) );
  NAND U2970 ( .A(n31), .B(n2820), .Z(n2822) );
  XOR U2971 ( .A(b[3]), .B(a[122]), .Z(n2843) );
  NAND U2972 ( .A(n5811), .B(n2843), .Z(n2821) );
  AND U2973 ( .A(n2822), .B(n2821), .Z(n2851) );
  NAND U2974 ( .A(b[0]), .B(a[124]), .Z(n2823) );
  XNOR U2975 ( .A(b[1]), .B(n2823), .Z(n2825) );
  NANDN U2976 ( .A(b[0]), .B(a[123]), .Z(n2824) );
  NAND U2977 ( .A(n2825), .B(n2824), .Z(n2850) );
  AND U2978 ( .A(b[3]), .B(a[120]), .Z(n2849) );
  XOR U2979 ( .A(n2850), .B(n2849), .Z(n2852) );
  XOR U2980 ( .A(n2851), .B(n2852), .Z(n2838) );
  NANDN U2981 ( .A(n2827), .B(n2826), .Z(n2831) );
  OR U2982 ( .A(n2829), .B(n2828), .Z(n2830) );
  AND U2983 ( .A(n2831), .B(n2830), .Z(n2837) );
  XOR U2984 ( .A(n2838), .B(n2837), .Z(n2840) );
  XOR U2985 ( .A(n2839), .B(n2840), .Z(n2855) );
  XNOR U2986 ( .A(n2855), .B(sreg[376]), .Z(n2857) );
  NANDN U2987 ( .A(n2832), .B(sreg[375]), .Z(n2836) );
  NAND U2988 ( .A(n2834), .B(n2833), .Z(n2835) );
  NAND U2989 ( .A(n2836), .B(n2835), .Z(n2856) );
  XOR U2990 ( .A(n2857), .B(n2856), .Z(c[376]) );
  NANDN U2991 ( .A(n2838), .B(n2837), .Z(n2842) );
  OR U2992 ( .A(n2840), .B(n2839), .Z(n2841) );
  AND U2993 ( .A(n2842), .B(n2841), .Z(n2862) );
  NAND U2994 ( .A(n31), .B(n2843), .Z(n2845) );
  XOR U2995 ( .A(b[3]), .B(a[123]), .Z(n2866) );
  NAND U2996 ( .A(n5811), .B(n2866), .Z(n2844) );
  AND U2997 ( .A(n2845), .B(n2844), .Z(n2874) );
  AND U2998 ( .A(b[3]), .B(a[121]), .Z(n2872) );
  NAND U2999 ( .A(b[0]), .B(a[125]), .Z(n2846) );
  XNOR U3000 ( .A(b[1]), .B(n2846), .Z(n2848) );
  NANDN U3001 ( .A(b[0]), .B(a[124]), .Z(n2847) );
  NAND U3002 ( .A(n2848), .B(n2847), .Z(n2873) );
  XOR U3003 ( .A(n2872), .B(n2873), .Z(n2875) );
  XOR U3004 ( .A(n2874), .B(n2875), .Z(n2861) );
  NANDN U3005 ( .A(n2850), .B(n2849), .Z(n2854) );
  OR U3006 ( .A(n2852), .B(n2851), .Z(n2853) );
  AND U3007 ( .A(n2854), .B(n2853), .Z(n2860) );
  XOR U3008 ( .A(n2861), .B(n2860), .Z(n2863) );
  XOR U3009 ( .A(n2862), .B(n2863), .Z(n2878) );
  XNOR U3010 ( .A(n2878), .B(sreg[377]), .Z(n2880) );
  NANDN U3011 ( .A(n2855), .B(sreg[376]), .Z(n2859) );
  NAND U3012 ( .A(n2857), .B(n2856), .Z(n2858) );
  NAND U3013 ( .A(n2859), .B(n2858), .Z(n2879) );
  XOR U3014 ( .A(n2880), .B(n2879), .Z(c[377]) );
  NANDN U3015 ( .A(n2861), .B(n2860), .Z(n2865) );
  OR U3016 ( .A(n2863), .B(n2862), .Z(n2864) );
  AND U3017 ( .A(n2865), .B(n2864), .Z(n2885) );
  NAND U3018 ( .A(n31), .B(n2866), .Z(n2868) );
  XOR U3019 ( .A(b[3]), .B(a[124]), .Z(n2889) );
  NAND U3020 ( .A(n5811), .B(n2889), .Z(n2867) );
  AND U3021 ( .A(n2868), .B(n2867), .Z(n2897) );
  NAND U3022 ( .A(b[0]), .B(a[126]), .Z(n2869) );
  XNOR U3023 ( .A(b[1]), .B(n2869), .Z(n2871) );
  NANDN U3024 ( .A(b[0]), .B(a[125]), .Z(n2870) );
  NAND U3025 ( .A(n2871), .B(n2870), .Z(n2896) );
  AND U3026 ( .A(b[3]), .B(a[122]), .Z(n2895) );
  XOR U3027 ( .A(n2896), .B(n2895), .Z(n2898) );
  XOR U3028 ( .A(n2897), .B(n2898), .Z(n2884) );
  NANDN U3029 ( .A(n2873), .B(n2872), .Z(n2877) );
  OR U3030 ( .A(n2875), .B(n2874), .Z(n2876) );
  AND U3031 ( .A(n2877), .B(n2876), .Z(n2883) );
  XOR U3032 ( .A(n2884), .B(n2883), .Z(n2886) );
  XOR U3033 ( .A(n2885), .B(n2886), .Z(n2901) );
  XNOR U3034 ( .A(n2901), .B(sreg[378]), .Z(n2903) );
  NANDN U3035 ( .A(n2878), .B(sreg[377]), .Z(n2882) );
  NAND U3036 ( .A(n2880), .B(n2879), .Z(n2881) );
  NAND U3037 ( .A(n2882), .B(n2881), .Z(n2902) );
  XOR U3038 ( .A(n2903), .B(n2902), .Z(c[378]) );
  NANDN U3039 ( .A(n2884), .B(n2883), .Z(n2888) );
  OR U3040 ( .A(n2886), .B(n2885), .Z(n2887) );
  AND U3041 ( .A(n2888), .B(n2887), .Z(n2908) );
  NAND U3042 ( .A(n31), .B(n2889), .Z(n2891) );
  XOR U3043 ( .A(b[3]), .B(a[125]), .Z(n2912) );
  NAND U3044 ( .A(n5811), .B(n2912), .Z(n2890) );
  AND U3045 ( .A(n2891), .B(n2890), .Z(n2920) );
  AND U3046 ( .A(b[3]), .B(a[123]), .Z(n2918) );
  NAND U3047 ( .A(b[0]), .B(a[127]), .Z(n2892) );
  XNOR U3048 ( .A(b[1]), .B(n2892), .Z(n2894) );
  NANDN U3049 ( .A(b[0]), .B(a[126]), .Z(n2893) );
  NAND U3050 ( .A(n2894), .B(n2893), .Z(n2919) );
  XOR U3051 ( .A(n2918), .B(n2919), .Z(n2921) );
  XOR U3052 ( .A(n2920), .B(n2921), .Z(n2907) );
  NANDN U3053 ( .A(n2896), .B(n2895), .Z(n2900) );
  OR U3054 ( .A(n2898), .B(n2897), .Z(n2899) );
  AND U3055 ( .A(n2900), .B(n2899), .Z(n2906) );
  XOR U3056 ( .A(n2907), .B(n2906), .Z(n2909) );
  XOR U3057 ( .A(n2908), .B(n2909), .Z(n2924) );
  XNOR U3058 ( .A(n2924), .B(sreg[379]), .Z(n2926) );
  NANDN U3059 ( .A(n2901), .B(sreg[378]), .Z(n2905) );
  NAND U3060 ( .A(n2903), .B(n2902), .Z(n2904) );
  NAND U3061 ( .A(n2905), .B(n2904), .Z(n2925) );
  XOR U3062 ( .A(n2926), .B(n2925), .Z(c[379]) );
  NANDN U3063 ( .A(n2907), .B(n2906), .Z(n2911) );
  OR U3064 ( .A(n2909), .B(n2908), .Z(n2910) );
  AND U3065 ( .A(n2911), .B(n2910), .Z(n2931) );
  NAND U3066 ( .A(n31), .B(n2912), .Z(n2914) );
  XOR U3067 ( .A(b[3]), .B(a[126]), .Z(n2935) );
  NAND U3068 ( .A(n5811), .B(n2935), .Z(n2913) );
  AND U3069 ( .A(n2914), .B(n2913), .Z(n2943) );
  AND U3070 ( .A(b[3]), .B(a[124]), .Z(n2941) );
  NAND U3071 ( .A(b[0]), .B(a[128]), .Z(n2915) );
  XNOR U3072 ( .A(b[1]), .B(n2915), .Z(n2917) );
  NANDN U3073 ( .A(b[0]), .B(a[127]), .Z(n2916) );
  NAND U3074 ( .A(n2917), .B(n2916), .Z(n2942) );
  XOR U3075 ( .A(n2941), .B(n2942), .Z(n2944) );
  XOR U3076 ( .A(n2943), .B(n2944), .Z(n2930) );
  NANDN U3077 ( .A(n2919), .B(n2918), .Z(n2923) );
  OR U3078 ( .A(n2921), .B(n2920), .Z(n2922) );
  AND U3079 ( .A(n2923), .B(n2922), .Z(n2929) );
  XOR U3080 ( .A(n2930), .B(n2929), .Z(n2932) );
  XOR U3081 ( .A(n2931), .B(n2932), .Z(n2947) );
  XNOR U3082 ( .A(n2947), .B(sreg[380]), .Z(n2949) );
  NANDN U3083 ( .A(n2924), .B(sreg[379]), .Z(n2928) );
  NAND U3084 ( .A(n2926), .B(n2925), .Z(n2927) );
  NAND U3085 ( .A(n2928), .B(n2927), .Z(n2948) );
  XOR U3086 ( .A(n2949), .B(n2948), .Z(c[380]) );
  NANDN U3087 ( .A(n2930), .B(n2929), .Z(n2934) );
  OR U3088 ( .A(n2932), .B(n2931), .Z(n2933) );
  AND U3089 ( .A(n2934), .B(n2933), .Z(n2954) );
  NAND U3090 ( .A(n31), .B(n2935), .Z(n2937) );
  XOR U3091 ( .A(b[3]), .B(a[127]), .Z(n2958) );
  NAND U3092 ( .A(n5811), .B(n2958), .Z(n2936) );
  AND U3093 ( .A(n2937), .B(n2936), .Z(n2966) );
  NAND U3094 ( .A(b[0]), .B(a[129]), .Z(n2938) );
  XNOR U3095 ( .A(b[1]), .B(n2938), .Z(n2940) );
  NANDN U3096 ( .A(b[0]), .B(a[128]), .Z(n2939) );
  NAND U3097 ( .A(n2940), .B(n2939), .Z(n2965) );
  AND U3098 ( .A(b[3]), .B(a[125]), .Z(n2964) );
  XOR U3099 ( .A(n2965), .B(n2964), .Z(n2967) );
  XOR U3100 ( .A(n2966), .B(n2967), .Z(n2953) );
  NANDN U3101 ( .A(n2942), .B(n2941), .Z(n2946) );
  OR U3102 ( .A(n2944), .B(n2943), .Z(n2945) );
  AND U3103 ( .A(n2946), .B(n2945), .Z(n2952) );
  XOR U3104 ( .A(n2953), .B(n2952), .Z(n2955) );
  XOR U3105 ( .A(n2954), .B(n2955), .Z(n2970) );
  XNOR U3106 ( .A(n2970), .B(sreg[381]), .Z(n2972) );
  NANDN U3107 ( .A(n2947), .B(sreg[380]), .Z(n2951) );
  NAND U3108 ( .A(n2949), .B(n2948), .Z(n2950) );
  NAND U3109 ( .A(n2951), .B(n2950), .Z(n2971) );
  XOR U3110 ( .A(n2972), .B(n2971), .Z(c[381]) );
  NANDN U3111 ( .A(n2953), .B(n2952), .Z(n2957) );
  OR U3112 ( .A(n2955), .B(n2954), .Z(n2956) );
  AND U3113 ( .A(n2957), .B(n2956), .Z(n2977) );
  NAND U3114 ( .A(n31), .B(n2958), .Z(n2960) );
  XOR U3115 ( .A(b[3]), .B(a[128]), .Z(n2981) );
  NAND U3116 ( .A(n5811), .B(n2981), .Z(n2959) );
  AND U3117 ( .A(n2960), .B(n2959), .Z(n2989) );
  NAND U3118 ( .A(b[0]), .B(a[130]), .Z(n2961) );
  XNOR U3119 ( .A(b[1]), .B(n2961), .Z(n2963) );
  NANDN U3120 ( .A(b[0]), .B(a[129]), .Z(n2962) );
  NAND U3121 ( .A(n2963), .B(n2962), .Z(n2988) );
  AND U3122 ( .A(b[3]), .B(a[126]), .Z(n2987) );
  XOR U3123 ( .A(n2988), .B(n2987), .Z(n2990) );
  XOR U3124 ( .A(n2989), .B(n2990), .Z(n2976) );
  NANDN U3125 ( .A(n2965), .B(n2964), .Z(n2969) );
  OR U3126 ( .A(n2967), .B(n2966), .Z(n2968) );
  AND U3127 ( .A(n2969), .B(n2968), .Z(n2975) );
  XOR U3128 ( .A(n2976), .B(n2975), .Z(n2978) );
  XOR U3129 ( .A(n2977), .B(n2978), .Z(n2993) );
  XNOR U3130 ( .A(n2993), .B(sreg[382]), .Z(n2995) );
  NANDN U3131 ( .A(n2970), .B(sreg[381]), .Z(n2974) );
  NAND U3132 ( .A(n2972), .B(n2971), .Z(n2973) );
  NAND U3133 ( .A(n2974), .B(n2973), .Z(n2994) );
  XOR U3134 ( .A(n2995), .B(n2994), .Z(c[382]) );
  NANDN U3135 ( .A(n2976), .B(n2975), .Z(n2980) );
  OR U3136 ( .A(n2978), .B(n2977), .Z(n2979) );
  AND U3137 ( .A(n2980), .B(n2979), .Z(n3000) );
  NAND U3138 ( .A(n31), .B(n2981), .Z(n2983) );
  XOR U3139 ( .A(b[3]), .B(a[129]), .Z(n3004) );
  NAND U3140 ( .A(n5811), .B(n3004), .Z(n2982) );
  AND U3141 ( .A(n2983), .B(n2982), .Z(n3012) );
  NAND U3142 ( .A(b[0]), .B(a[131]), .Z(n2984) );
  XNOR U3143 ( .A(b[1]), .B(n2984), .Z(n2986) );
  NANDN U3144 ( .A(b[0]), .B(a[130]), .Z(n2985) );
  NAND U3145 ( .A(n2986), .B(n2985), .Z(n3011) );
  AND U3146 ( .A(b[3]), .B(a[127]), .Z(n3010) );
  XOR U3147 ( .A(n3011), .B(n3010), .Z(n3013) );
  XOR U3148 ( .A(n3012), .B(n3013), .Z(n2999) );
  NANDN U3149 ( .A(n2988), .B(n2987), .Z(n2992) );
  OR U3150 ( .A(n2990), .B(n2989), .Z(n2991) );
  AND U3151 ( .A(n2992), .B(n2991), .Z(n2998) );
  XOR U3152 ( .A(n2999), .B(n2998), .Z(n3001) );
  XOR U3153 ( .A(n3000), .B(n3001), .Z(n3016) );
  XNOR U3154 ( .A(n3016), .B(sreg[383]), .Z(n3018) );
  NANDN U3155 ( .A(n2993), .B(sreg[382]), .Z(n2997) );
  NAND U3156 ( .A(n2995), .B(n2994), .Z(n2996) );
  NAND U3157 ( .A(n2997), .B(n2996), .Z(n3017) );
  XOR U3158 ( .A(n3018), .B(n3017), .Z(c[383]) );
  NANDN U3159 ( .A(n2999), .B(n2998), .Z(n3003) );
  OR U3160 ( .A(n3001), .B(n3000), .Z(n3002) );
  AND U3161 ( .A(n3003), .B(n3002), .Z(n3023) );
  NAND U3162 ( .A(n31), .B(n3004), .Z(n3006) );
  XOR U3163 ( .A(b[3]), .B(a[130]), .Z(n3027) );
  NAND U3164 ( .A(n5811), .B(n3027), .Z(n3005) );
  AND U3165 ( .A(n3006), .B(n3005), .Z(n3035) );
  AND U3166 ( .A(b[3]), .B(a[128]), .Z(n3033) );
  NAND U3167 ( .A(b[0]), .B(a[132]), .Z(n3007) );
  XNOR U3168 ( .A(b[1]), .B(n3007), .Z(n3009) );
  NANDN U3169 ( .A(b[0]), .B(a[131]), .Z(n3008) );
  NAND U3170 ( .A(n3009), .B(n3008), .Z(n3034) );
  XOR U3171 ( .A(n3033), .B(n3034), .Z(n3036) );
  XOR U3172 ( .A(n3035), .B(n3036), .Z(n3022) );
  NANDN U3173 ( .A(n3011), .B(n3010), .Z(n3015) );
  OR U3174 ( .A(n3013), .B(n3012), .Z(n3014) );
  AND U3175 ( .A(n3015), .B(n3014), .Z(n3021) );
  XOR U3176 ( .A(n3022), .B(n3021), .Z(n3024) );
  XOR U3177 ( .A(n3023), .B(n3024), .Z(n3039) );
  XNOR U3178 ( .A(n3039), .B(sreg[384]), .Z(n3041) );
  NANDN U3179 ( .A(n3016), .B(sreg[383]), .Z(n3020) );
  NAND U3180 ( .A(n3018), .B(n3017), .Z(n3019) );
  NAND U3181 ( .A(n3020), .B(n3019), .Z(n3040) );
  XOR U3182 ( .A(n3041), .B(n3040), .Z(c[384]) );
  NANDN U3183 ( .A(n3022), .B(n3021), .Z(n3026) );
  OR U3184 ( .A(n3024), .B(n3023), .Z(n3025) );
  AND U3185 ( .A(n3026), .B(n3025), .Z(n3046) );
  NAND U3186 ( .A(n31), .B(n3027), .Z(n3029) );
  XOR U3187 ( .A(b[3]), .B(a[131]), .Z(n3050) );
  NAND U3188 ( .A(n5811), .B(n3050), .Z(n3028) );
  AND U3189 ( .A(n3029), .B(n3028), .Z(n3058) );
  AND U3190 ( .A(b[3]), .B(a[129]), .Z(n3056) );
  NAND U3191 ( .A(b[0]), .B(a[133]), .Z(n3030) );
  XNOR U3192 ( .A(b[1]), .B(n3030), .Z(n3032) );
  NANDN U3193 ( .A(b[0]), .B(a[132]), .Z(n3031) );
  NAND U3194 ( .A(n3032), .B(n3031), .Z(n3057) );
  XOR U3195 ( .A(n3056), .B(n3057), .Z(n3059) );
  XOR U3196 ( .A(n3058), .B(n3059), .Z(n3045) );
  NANDN U3197 ( .A(n3034), .B(n3033), .Z(n3038) );
  OR U3198 ( .A(n3036), .B(n3035), .Z(n3037) );
  AND U3199 ( .A(n3038), .B(n3037), .Z(n3044) );
  XOR U3200 ( .A(n3045), .B(n3044), .Z(n3047) );
  XOR U3201 ( .A(n3046), .B(n3047), .Z(n3062) );
  XNOR U3202 ( .A(n3062), .B(sreg[385]), .Z(n3064) );
  NANDN U3203 ( .A(n3039), .B(sreg[384]), .Z(n3043) );
  NAND U3204 ( .A(n3041), .B(n3040), .Z(n3042) );
  NAND U3205 ( .A(n3043), .B(n3042), .Z(n3063) );
  XOR U3206 ( .A(n3064), .B(n3063), .Z(c[385]) );
  NANDN U3207 ( .A(n3045), .B(n3044), .Z(n3049) );
  OR U3208 ( .A(n3047), .B(n3046), .Z(n3048) );
  AND U3209 ( .A(n3049), .B(n3048), .Z(n3069) );
  NAND U3210 ( .A(n31), .B(n3050), .Z(n3052) );
  XOR U3211 ( .A(b[3]), .B(a[132]), .Z(n3073) );
  NAND U3212 ( .A(n5811), .B(n3073), .Z(n3051) );
  AND U3213 ( .A(n3052), .B(n3051), .Z(n3081) );
  NAND U3214 ( .A(b[0]), .B(a[134]), .Z(n3053) );
  XNOR U3215 ( .A(b[1]), .B(n3053), .Z(n3055) );
  NANDN U3216 ( .A(b[0]), .B(a[133]), .Z(n3054) );
  NAND U3217 ( .A(n3055), .B(n3054), .Z(n3080) );
  AND U3218 ( .A(b[3]), .B(a[130]), .Z(n3079) );
  XOR U3219 ( .A(n3080), .B(n3079), .Z(n3082) );
  XOR U3220 ( .A(n3081), .B(n3082), .Z(n3068) );
  NANDN U3221 ( .A(n3057), .B(n3056), .Z(n3061) );
  OR U3222 ( .A(n3059), .B(n3058), .Z(n3060) );
  AND U3223 ( .A(n3061), .B(n3060), .Z(n3067) );
  XOR U3224 ( .A(n3068), .B(n3067), .Z(n3070) );
  XOR U3225 ( .A(n3069), .B(n3070), .Z(n3085) );
  XNOR U3226 ( .A(n3085), .B(sreg[386]), .Z(n3087) );
  NANDN U3227 ( .A(n3062), .B(sreg[385]), .Z(n3066) );
  NAND U3228 ( .A(n3064), .B(n3063), .Z(n3065) );
  NAND U3229 ( .A(n3066), .B(n3065), .Z(n3086) );
  XOR U3230 ( .A(n3087), .B(n3086), .Z(c[386]) );
  NANDN U3231 ( .A(n3068), .B(n3067), .Z(n3072) );
  OR U3232 ( .A(n3070), .B(n3069), .Z(n3071) );
  AND U3233 ( .A(n3072), .B(n3071), .Z(n3092) );
  NAND U3234 ( .A(n31), .B(n3073), .Z(n3075) );
  XOR U3235 ( .A(b[3]), .B(a[133]), .Z(n3096) );
  NAND U3236 ( .A(n5811), .B(n3096), .Z(n3074) );
  AND U3237 ( .A(n3075), .B(n3074), .Z(n3104) );
  AND U3238 ( .A(b[3]), .B(a[131]), .Z(n3102) );
  NAND U3239 ( .A(b[0]), .B(a[135]), .Z(n3076) );
  XNOR U3240 ( .A(b[1]), .B(n3076), .Z(n3078) );
  NANDN U3241 ( .A(b[0]), .B(a[134]), .Z(n3077) );
  NAND U3242 ( .A(n3078), .B(n3077), .Z(n3103) );
  XOR U3243 ( .A(n3102), .B(n3103), .Z(n3105) );
  XOR U3244 ( .A(n3104), .B(n3105), .Z(n3091) );
  NANDN U3245 ( .A(n3080), .B(n3079), .Z(n3084) );
  OR U3246 ( .A(n3082), .B(n3081), .Z(n3083) );
  AND U3247 ( .A(n3084), .B(n3083), .Z(n3090) );
  XOR U3248 ( .A(n3091), .B(n3090), .Z(n3093) );
  XOR U3249 ( .A(n3092), .B(n3093), .Z(n3108) );
  XNOR U3250 ( .A(n3108), .B(sreg[387]), .Z(n3110) );
  NANDN U3251 ( .A(n3085), .B(sreg[386]), .Z(n3089) );
  NAND U3252 ( .A(n3087), .B(n3086), .Z(n3088) );
  NAND U3253 ( .A(n3089), .B(n3088), .Z(n3109) );
  XOR U3254 ( .A(n3110), .B(n3109), .Z(c[387]) );
  NANDN U3255 ( .A(n3091), .B(n3090), .Z(n3095) );
  OR U3256 ( .A(n3093), .B(n3092), .Z(n3094) );
  AND U3257 ( .A(n3095), .B(n3094), .Z(n3115) );
  NAND U3258 ( .A(n31), .B(n3096), .Z(n3098) );
  XOR U3259 ( .A(b[3]), .B(a[134]), .Z(n3119) );
  NAND U3260 ( .A(n5811), .B(n3119), .Z(n3097) );
  AND U3261 ( .A(n3098), .B(n3097), .Z(n3127) );
  NAND U3262 ( .A(b[0]), .B(a[136]), .Z(n3099) );
  XNOR U3263 ( .A(b[1]), .B(n3099), .Z(n3101) );
  NANDN U3264 ( .A(b[0]), .B(a[135]), .Z(n3100) );
  NAND U3265 ( .A(n3101), .B(n3100), .Z(n3126) );
  AND U3266 ( .A(b[3]), .B(a[132]), .Z(n3125) );
  XOR U3267 ( .A(n3126), .B(n3125), .Z(n3128) );
  XOR U3268 ( .A(n3127), .B(n3128), .Z(n3114) );
  NANDN U3269 ( .A(n3103), .B(n3102), .Z(n3107) );
  OR U3270 ( .A(n3105), .B(n3104), .Z(n3106) );
  AND U3271 ( .A(n3107), .B(n3106), .Z(n3113) );
  XOR U3272 ( .A(n3114), .B(n3113), .Z(n3116) );
  XOR U3273 ( .A(n3115), .B(n3116), .Z(n3131) );
  XNOR U3274 ( .A(n3131), .B(sreg[388]), .Z(n3133) );
  NANDN U3275 ( .A(n3108), .B(sreg[387]), .Z(n3112) );
  NAND U3276 ( .A(n3110), .B(n3109), .Z(n3111) );
  NAND U3277 ( .A(n3112), .B(n3111), .Z(n3132) );
  XOR U3278 ( .A(n3133), .B(n3132), .Z(c[388]) );
  NANDN U3279 ( .A(n3114), .B(n3113), .Z(n3118) );
  OR U3280 ( .A(n3116), .B(n3115), .Z(n3117) );
  AND U3281 ( .A(n3118), .B(n3117), .Z(n3138) );
  NAND U3282 ( .A(n31), .B(n3119), .Z(n3121) );
  XOR U3283 ( .A(b[3]), .B(a[135]), .Z(n3142) );
  NAND U3284 ( .A(n5811), .B(n3142), .Z(n3120) );
  AND U3285 ( .A(n3121), .B(n3120), .Z(n3150) );
  NAND U3286 ( .A(b[0]), .B(a[137]), .Z(n3122) );
  XNOR U3287 ( .A(b[1]), .B(n3122), .Z(n3124) );
  NANDN U3288 ( .A(b[0]), .B(a[136]), .Z(n3123) );
  NAND U3289 ( .A(n3124), .B(n3123), .Z(n3149) );
  AND U3290 ( .A(b[3]), .B(a[133]), .Z(n3148) );
  XOR U3291 ( .A(n3149), .B(n3148), .Z(n3151) );
  XOR U3292 ( .A(n3150), .B(n3151), .Z(n3137) );
  NANDN U3293 ( .A(n3126), .B(n3125), .Z(n3130) );
  OR U3294 ( .A(n3128), .B(n3127), .Z(n3129) );
  AND U3295 ( .A(n3130), .B(n3129), .Z(n3136) );
  XOR U3296 ( .A(n3137), .B(n3136), .Z(n3139) );
  XOR U3297 ( .A(n3138), .B(n3139), .Z(n3154) );
  XNOR U3298 ( .A(n3154), .B(sreg[389]), .Z(n3156) );
  NANDN U3299 ( .A(n3131), .B(sreg[388]), .Z(n3135) );
  NAND U3300 ( .A(n3133), .B(n3132), .Z(n3134) );
  NAND U3301 ( .A(n3135), .B(n3134), .Z(n3155) );
  XOR U3302 ( .A(n3156), .B(n3155), .Z(c[389]) );
  NANDN U3303 ( .A(n3137), .B(n3136), .Z(n3141) );
  OR U3304 ( .A(n3139), .B(n3138), .Z(n3140) );
  AND U3305 ( .A(n3141), .B(n3140), .Z(n3161) );
  NAND U3306 ( .A(n31), .B(n3142), .Z(n3144) );
  XOR U3307 ( .A(b[3]), .B(a[136]), .Z(n3165) );
  NAND U3308 ( .A(n5811), .B(n3165), .Z(n3143) );
  AND U3309 ( .A(n3144), .B(n3143), .Z(n3173) );
  AND U3310 ( .A(b[3]), .B(a[134]), .Z(n3171) );
  NAND U3311 ( .A(b[0]), .B(a[138]), .Z(n3145) );
  XNOR U3312 ( .A(b[1]), .B(n3145), .Z(n3147) );
  NANDN U3313 ( .A(b[0]), .B(a[137]), .Z(n3146) );
  NAND U3314 ( .A(n3147), .B(n3146), .Z(n3172) );
  XOR U3315 ( .A(n3171), .B(n3172), .Z(n3174) );
  XOR U3316 ( .A(n3173), .B(n3174), .Z(n3160) );
  NANDN U3317 ( .A(n3149), .B(n3148), .Z(n3153) );
  OR U3318 ( .A(n3151), .B(n3150), .Z(n3152) );
  AND U3319 ( .A(n3153), .B(n3152), .Z(n3159) );
  XOR U3320 ( .A(n3160), .B(n3159), .Z(n3162) );
  XOR U3321 ( .A(n3161), .B(n3162), .Z(n3177) );
  XNOR U3322 ( .A(n3177), .B(sreg[390]), .Z(n3179) );
  NANDN U3323 ( .A(n3154), .B(sreg[389]), .Z(n3158) );
  NAND U3324 ( .A(n3156), .B(n3155), .Z(n3157) );
  NAND U3325 ( .A(n3158), .B(n3157), .Z(n3178) );
  XOR U3326 ( .A(n3179), .B(n3178), .Z(c[390]) );
  NANDN U3327 ( .A(n3160), .B(n3159), .Z(n3164) );
  OR U3328 ( .A(n3162), .B(n3161), .Z(n3163) );
  AND U3329 ( .A(n3164), .B(n3163), .Z(n3184) );
  NAND U3330 ( .A(n31), .B(n3165), .Z(n3167) );
  XOR U3331 ( .A(b[3]), .B(a[137]), .Z(n3188) );
  NAND U3332 ( .A(n5811), .B(n3188), .Z(n3166) );
  AND U3333 ( .A(n3167), .B(n3166), .Z(n3196) );
  NAND U3334 ( .A(b[0]), .B(a[139]), .Z(n3168) );
  XNOR U3335 ( .A(b[1]), .B(n3168), .Z(n3170) );
  NANDN U3336 ( .A(b[0]), .B(a[138]), .Z(n3169) );
  NAND U3337 ( .A(n3170), .B(n3169), .Z(n3195) );
  AND U3338 ( .A(b[3]), .B(a[135]), .Z(n3194) );
  XOR U3339 ( .A(n3195), .B(n3194), .Z(n3197) );
  XOR U3340 ( .A(n3196), .B(n3197), .Z(n3183) );
  NANDN U3341 ( .A(n3172), .B(n3171), .Z(n3176) );
  OR U3342 ( .A(n3174), .B(n3173), .Z(n3175) );
  AND U3343 ( .A(n3176), .B(n3175), .Z(n3182) );
  XOR U3344 ( .A(n3183), .B(n3182), .Z(n3185) );
  XOR U3345 ( .A(n3184), .B(n3185), .Z(n3200) );
  XNOR U3346 ( .A(n3200), .B(sreg[391]), .Z(n3202) );
  NANDN U3347 ( .A(n3177), .B(sreg[390]), .Z(n3181) );
  NAND U3348 ( .A(n3179), .B(n3178), .Z(n3180) );
  NAND U3349 ( .A(n3181), .B(n3180), .Z(n3201) );
  XOR U3350 ( .A(n3202), .B(n3201), .Z(c[391]) );
  NANDN U3351 ( .A(n3183), .B(n3182), .Z(n3187) );
  OR U3352 ( .A(n3185), .B(n3184), .Z(n3186) );
  AND U3353 ( .A(n3187), .B(n3186), .Z(n3207) );
  NAND U3354 ( .A(n31), .B(n3188), .Z(n3190) );
  XOR U3355 ( .A(b[3]), .B(a[138]), .Z(n3211) );
  NAND U3356 ( .A(n5811), .B(n3211), .Z(n3189) );
  AND U3357 ( .A(n3190), .B(n3189), .Z(n3219) );
  AND U3358 ( .A(b[3]), .B(a[136]), .Z(n3217) );
  NAND U3359 ( .A(b[0]), .B(a[140]), .Z(n3191) );
  XNOR U3360 ( .A(b[1]), .B(n3191), .Z(n3193) );
  NANDN U3361 ( .A(b[0]), .B(a[139]), .Z(n3192) );
  NAND U3362 ( .A(n3193), .B(n3192), .Z(n3218) );
  XOR U3363 ( .A(n3217), .B(n3218), .Z(n3220) );
  XOR U3364 ( .A(n3219), .B(n3220), .Z(n3206) );
  NANDN U3365 ( .A(n3195), .B(n3194), .Z(n3199) );
  OR U3366 ( .A(n3197), .B(n3196), .Z(n3198) );
  AND U3367 ( .A(n3199), .B(n3198), .Z(n3205) );
  XOR U3368 ( .A(n3206), .B(n3205), .Z(n3208) );
  XOR U3369 ( .A(n3207), .B(n3208), .Z(n3223) );
  XNOR U3370 ( .A(n3223), .B(sreg[392]), .Z(n3225) );
  NANDN U3371 ( .A(n3200), .B(sreg[391]), .Z(n3204) );
  NAND U3372 ( .A(n3202), .B(n3201), .Z(n3203) );
  NAND U3373 ( .A(n3204), .B(n3203), .Z(n3224) );
  XOR U3374 ( .A(n3225), .B(n3224), .Z(c[392]) );
  NANDN U3375 ( .A(n3206), .B(n3205), .Z(n3210) );
  OR U3376 ( .A(n3208), .B(n3207), .Z(n3209) );
  AND U3377 ( .A(n3210), .B(n3209), .Z(n3230) );
  NAND U3378 ( .A(n31), .B(n3211), .Z(n3213) );
  XOR U3379 ( .A(b[3]), .B(a[139]), .Z(n3234) );
  NAND U3380 ( .A(n5811), .B(n3234), .Z(n3212) );
  AND U3381 ( .A(n3213), .B(n3212), .Z(n3242) );
  NAND U3382 ( .A(b[0]), .B(a[141]), .Z(n3214) );
  XNOR U3383 ( .A(b[1]), .B(n3214), .Z(n3216) );
  NANDN U3384 ( .A(b[0]), .B(a[140]), .Z(n3215) );
  NAND U3385 ( .A(n3216), .B(n3215), .Z(n3241) );
  AND U3386 ( .A(b[3]), .B(a[137]), .Z(n3240) );
  XOR U3387 ( .A(n3241), .B(n3240), .Z(n3243) );
  XOR U3388 ( .A(n3242), .B(n3243), .Z(n3229) );
  NANDN U3389 ( .A(n3218), .B(n3217), .Z(n3222) );
  OR U3390 ( .A(n3220), .B(n3219), .Z(n3221) );
  AND U3391 ( .A(n3222), .B(n3221), .Z(n3228) );
  XOR U3392 ( .A(n3229), .B(n3228), .Z(n3231) );
  XOR U3393 ( .A(n3230), .B(n3231), .Z(n3246) );
  XNOR U3394 ( .A(n3246), .B(sreg[393]), .Z(n3248) );
  NANDN U3395 ( .A(n3223), .B(sreg[392]), .Z(n3227) );
  NAND U3396 ( .A(n3225), .B(n3224), .Z(n3226) );
  NAND U3397 ( .A(n3227), .B(n3226), .Z(n3247) );
  XOR U3398 ( .A(n3248), .B(n3247), .Z(c[393]) );
  NANDN U3399 ( .A(n3229), .B(n3228), .Z(n3233) );
  OR U3400 ( .A(n3231), .B(n3230), .Z(n3232) );
  AND U3401 ( .A(n3233), .B(n3232), .Z(n3253) );
  NAND U3402 ( .A(n31), .B(n3234), .Z(n3236) );
  XOR U3403 ( .A(b[3]), .B(a[140]), .Z(n3257) );
  NAND U3404 ( .A(n5811), .B(n3257), .Z(n3235) );
  AND U3405 ( .A(n3236), .B(n3235), .Z(n3265) );
  NAND U3406 ( .A(b[0]), .B(a[142]), .Z(n3237) );
  XNOR U3407 ( .A(b[1]), .B(n3237), .Z(n3239) );
  NANDN U3408 ( .A(b[0]), .B(a[141]), .Z(n3238) );
  NAND U3409 ( .A(n3239), .B(n3238), .Z(n3264) );
  AND U3410 ( .A(b[3]), .B(a[138]), .Z(n3263) );
  XOR U3411 ( .A(n3264), .B(n3263), .Z(n3266) );
  XOR U3412 ( .A(n3265), .B(n3266), .Z(n3252) );
  NANDN U3413 ( .A(n3241), .B(n3240), .Z(n3245) );
  OR U3414 ( .A(n3243), .B(n3242), .Z(n3244) );
  AND U3415 ( .A(n3245), .B(n3244), .Z(n3251) );
  XOR U3416 ( .A(n3252), .B(n3251), .Z(n3254) );
  XOR U3417 ( .A(n3253), .B(n3254), .Z(n3269) );
  XNOR U3418 ( .A(n3269), .B(sreg[394]), .Z(n3271) );
  NANDN U3419 ( .A(n3246), .B(sreg[393]), .Z(n3250) );
  NAND U3420 ( .A(n3248), .B(n3247), .Z(n3249) );
  NAND U3421 ( .A(n3250), .B(n3249), .Z(n3270) );
  XOR U3422 ( .A(n3271), .B(n3270), .Z(c[394]) );
  NANDN U3423 ( .A(n3252), .B(n3251), .Z(n3256) );
  OR U3424 ( .A(n3254), .B(n3253), .Z(n3255) );
  AND U3425 ( .A(n3256), .B(n3255), .Z(n3276) );
  NAND U3426 ( .A(n31), .B(n3257), .Z(n3259) );
  XOR U3427 ( .A(b[3]), .B(a[141]), .Z(n3280) );
  NAND U3428 ( .A(n5811), .B(n3280), .Z(n3258) );
  AND U3429 ( .A(n3259), .B(n3258), .Z(n3288) );
  NAND U3430 ( .A(b[0]), .B(a[143]), .Z(n3260) );
  XNOR U3431 ( .A(b[1]), .B(n3260), .Z(n3262) );
  NANDN U3432 ( .A(b[0]), .B(a[142]), .Z(n3261) );
  NAND U3433 ( .A(n3262), .B(n3261), .Z(n3287) );
  AND U3434 ( .A(b[3]), .B(a[139]), .Z(n3286) );
  XOR U3435 ( .A(n3287), .B(n3286), .Z(n3289) );
  XOR U3436 ( .A(n3288), .B(n3289), .Z(n3275) );
  NANDN U3437 ( .A(n3264), .B(n3263), .Z(n3268) );
  OR U3438 ( .A(n3266), .B(n3265), .Z(n3267) );
  AND U3439 ( .A(n3268), .B(n3267), .Z(n3274) );
  XOR U3440 ( .A(n3275), .B(n3274), .Z(n3277) );
  XOR U3441 ( .A(n3276), .B(n3277), .Z(n3292) );
  XNOR U3442 ( .A(n3292), .B(sreg[395]), .Z(n3294) );
  NANDN U3443 ( .A(n3269), .B(sreg[394]), .Z(n3273) );
  NAND U3444 ( .A(n3271), .B(n3270), .Z(n3272) );
  NAND U3445 ( .A(n3273), .B(n3272), .Z(n3293) );
  XOR U3446 ( .A(n3294), .B(n3293), .Z(c[395]) );
  NANDN U3447 ( .A(n3275), .B(n3274), .Z(n3279) );
  OR U3448 ( .A(n3277), .B(n3276), .Z(n3278) );
  AND U3449 ( .A(n3279), .B(n3278), .Z(n3299) );
  NAND U3450 ( .A(n31), .B(n3280), .Z(n3282) );
  XOR U3451 ( .A(b[3]), .B(a[142]), .Z(n3303) );
  NAND U3452 ( .A(n5811), .B(n3303), .Z(n3281) );
  AND U3453 ( .A(n3282), .B(n3281), .Z(n3311) );
  NAND U3454 ( .A(b[0]), .B(a[144]), .Z(n3283) );
  XNOR U3455 ( .A(b[1]), .B(n3283), .Z(n3285) );
  NANDN U3456 ( .A(b[0]), .B(a[143]), .Z(n3284) );
  NAND U3457 ( .A(n3285), .B(n3284), .Z(n3310) );
  AND U3458 ( .A(b[3]), .B(a[140]), .Z(n3309) );
  XOR U3459 ( .A(n3310), .B(n3309), .Z(n3312) );
  XOR U3460 ( .A(n3311), .B(n3312), .Z(n3298) );
  NANDN U3461 ( .A(n3287), .B(n3286), .Z(n3291) );
  OR U3462 ( .A(n3289), .B(n3288), .Z(n3290) );
  AND U3463 ( .A(n3291), .B(n3290), .Z(n3297) );
  XOR U3464 ( .A(n3298), .B(n3297), .Z(n3300) );
  XOR U3465 ( .A(n3299), .B(n3300), .Z(n3315) );
  XNOR U3466 ( .A(n3315), .B(sreg[396]), .Z(n3317) );
  NANDN U3467 ( .A(n3292), .B(sreg[395]), .Z(n3296) );
  NAND U3468 ( .A(n3294), .B(n3293), .Z(n3295) );
  NAND U3469 ( .A(n3296), .B(n3295), .Z(n3316) );
  XOR U3470 ( .A(n3317), .B(n3316), .Z(c[396]) );
  NANDN U3471 ( .A(n3298), .B(n3297), .Z(n3302) );
  OR U3472 ( .A(n3300), .B(n3299), .Z(n3301) );
  AND U3473 ( .A(n3302), .B(n3301), .Z(n3322) );
  NAND U3474 ( .A(n31), .B(n3303), .Z(n3305) );
  XOR U3475 ( .A(b[3]), .B(a[143]), .Z(n3326) );
  NAND U3476 ( .A(n5811), .B(n3326), .Z(n3304) );
  AND U3477 ( .A(n3305), .B(n3304), .Z(n3334) );
  NAND U3478 ( .A(b[0]), .B(a[145]), .Z(n3306) );
  XNOR U3479 ( .A(b[1]), .B(n3306), .Z(n3308) );
  NANDN U3480 ( .A(b[0]), .B(a[144]), .Z(n3307) );
  NAND U3481 ( .A(n3308), .B(n3307), .Z(n3333) );
  AND U3482 ( .A(b[3]), .B(a[141]), .Z(n3332) );
  XOR U3483 ( .A(n3333), .B(n3332), .Z(n3335) );
  XOR U3484 ( .A(n3334), .B(n3335), .Z(n3321) );
  NANDN U3485 ( .A(n3310), .B(n3309), .Z(n3314) );
  OR U3486 ( .A(n3312), .B(n3311), .Z(n3313) );
  AND U3487 ( .A(n3314), .B(n3313), .Z(n3320) );
  XOR U3488 ( .A(n3321), .B(n3320), .Z(n3323) );
  XOR U3489 ( .A(n3322), .B(n3323), .Z(n3338) );
  XNOR U3490 ( .A(n3338), .B(sreg[397]), .Z(n3340) );
  NANDN U3491 ( .A(n3315), .B(sreg[396]), .Z(n3319) );
  NAND U3492 ( .A(n3317), .B(n3316), .Z(n3318) );
  NAND U3493 ( .A(n3319), .B(n3318), .Z(n3339) );
  XOR U3494 ( .A(n3340), .B(n3339), .Z(c[397]) );
  NANDN U3495 ( .A(n3321), .B(n3320), .Z(n3325) );
  OR U3496 ( .A(n3323), .B(n3322), .Z(n3324) );
  AND U3497 ( .A(n3325), .B(n3324), .Z(n3345) );
  NAND U3498 ( .A(n31), .B(n3326), .Z(n3328) );
  XOR U3499 ( .A(b[3]), .B(a[144]), .Z(n3349) );
  NAND U3500 ( .A(n5811), .B(n3349), .Z(n3327) );
  AND U3501 ( .A(n3328), .B(n3327), .Z(n3357) );
  NAND U3502 ( .A(b[0]), .B(a[146]), .Z(n3329) );
  XNOR U3503 ( .A(b[1]), .B(n3329), .Z(n3331) );
  NANDN U3504 ( .A(b[0]), .B(a[145]), .Z(n3330) );
  NAND U3505 ( .A(n3331), .B(n3330), .Z(n3356) );
  AND U3506 ( .A(b[3]), .B(a[142]), .Z(n3355) );
  XOR U3507 ( .A(n3356), .B(n3355), .Z(n3358) );
  XOR U3508 ( .A(n3357), .B(n3358), .Z(n3344) );
  NANDN U3509 ( .A(n3333), .B(n3332), .Z(n3337) );
  OR U3510 ( .A(n3335), .B(n3334), .Z(n3336) );
  AND U3511 ( .A(n3337), .B(n3336), .Z(n3343) );
  XOR U3512 ( .A(n3344), .B(n3343), .Z(n3346) );
  XOR U3513 ( .A(n3345), .B(n3346), .Z(n3361) );
  XNOR U3514 ( .A(n3361), .B(sreg[398]), .Z(n3363) );
  NANDN U3515 ( .A(n3338), .B(sreg[397]), .Z(n3342) );
  NAND U3516 ( .A(n3340), .B(n3339), .Z(n3341) );
  NAND U3517 ( .A(n3342), .B(n3341), .Z(n3362) );
  XOR U3518 ( .A(n3363), .B(n3362), .Z(c[398]) );
  NANDN U3519 ( .A(n3344), .B(n3343), .Z(n3348) );
  OR U3520 ( .A(n3346), .B(n3345), .Z(n3347) );
  AND U3521 ( .A(n3348), .B(n3347), .Z(n3368) );
  NAND U3522 ( .A(n31), .B(n3349), .Z(n3351) );
  XOR U3523 ( .A(b[3]), .B(a[145]), .Z(n3372) );
  NAND U3524 ( .A(n5811), .B(n3372), .Z(n3350) );
  AND U3525 ( .A(n3351), .B(n3350), .Z(n3380) );
  NAND U3526 ( .A(b[0]), .B(a[147]), .Z(n3352) );
  XNOR U3527 ( .A(b[1]), .B(n3352), .Z(n3354) );
  NANDN U3528 ( .A(b[0]), .B(a[146]), .Z(n3353) );
  NAND U3529 ( .A(n3354), .B(n3353), .Z(n3379) );
  AND U3530 ( .A(b[3]), .B(a[143]), .Z(n3378) );
  XOR U3531 ( .A(n3379), .B(n3378), .Z(n3381) );
  XOR U3532 ( .A(n3380), .B(n3381), .Z(n3367) );
  NANDN U3533 ( .A(n3356), .B(n3355), .Z(n3360) );
  OR U3534 ( .A(n3358), .B(n3357), .Z(n3359) );
  AND U3535 ( .A(n3360), .B(n3359), .Z(n3366) );
  XOR U3536 ( .A(n3367), .B(n3366), .Z(n3369) );
  XOR U3537 ( .A(n3368), .B(n3369), .Z(n3384) );
  XNOR U3538 ( .A(n3384), .B(sreg[399]), .Z(n3386) );
  NANDN U3539 ( .A(n3361), .B(sreg[398]), .Z(n3365) );
  NAND U3540 ( .A(n3363), .B(n3362), .Z(n3364) );
  NAND U3541 ( .A(n3365), .B(n3364), .Z(n3385) );
  XOR U3542 ( .A(n3386), .B(n3385), .Z(c[399]) );
  NANDN U3543 ( .A(n3367), .B(n3366), .Z(n3371) );
  OR U3544 ( .A(n3369), .B(n3368), .Z(n3370) );
  AND U3545 ( .A(n3371), .B(n3370), .Z(n3391) );
  NAND U3546 ( .A(n31), .B(n3372), .Z(n3374) );
  XOR U3547 ( .A(b[3]), .B(a[146]), .Z(n3395) );
  NAND U3548 ( .A(n5811), .B(n3395), .Z(n3373) );
  AND U3549 ( .A(n3374), .B(n3373), .Z(n3403) );
  NAND U3550 ( .A(b[0]), .B(a[148]), .Z(n3375) );
  XNOR U3551 ( .A(b[1]), .B(n3375), .Z(n3377) );
  NANDN U3552 ( .A(b[0]), .B(a[147]), .Z(n3376) );
  NAND U3553 ( .A(n3377), .B(n3376), .Z(n3402) );
  AND U3554 ( .A(b[3]), .B(a[144]), .Z(n3401) );
  XOR U3555 ( .A(n3402), .B(n3401), .Z(n3404) );
  XOR U3556 ( .A(n3403), .B(n3404), .Z(n3390) );
  NANDN U3557 ( .A(n3379), .B(n3378), .Z(n3383) );
  OR U3558 ( .A(n3381), .B(n3380), .Z(n3382) );
  AND U3559 ( .A(n3383), .B(n3382), .Z(n3389) );
  XOR U3560 ( .A(n3390), .B(n3389), .Z(n3392) );
  XOR U3561 ( .A(n3391), .B(n3392), .Z(n3407) );
  XNOR U3562 ( .A(n3407), .B(sreg[400]), .Z(n3409) );
  NANDN U3563 ( .A(n3384), .B(sreg[399]), .Z(n3388) );
  NAND U3564 ( .A(n3386), .B(n3385), .Z(n3387) );
  NAND U3565 ( .A(n3388), .B(n3387), .Z(n3408) );
  XOR U3566 ( .A(n3409), .B(n3408), .Z(c[400]) );
  NANDN U3567 ( .A(n3390), .B(n3389), .Z(n3394) );
  OR U3568 ( .A(n3392), .B(n3391), .Z(n3393) );
  AND U3569 ( .A(n3394), .B(n3393), .Z(n3414) );
  NAND U3570 ( .A(n31), .B(n3395), .Z(n3397) );
  XOR U3571 ( .A(b[3]), .B(a[147]), .Z(n3418) );
  NAND U3572 ( .A(n5811), .B(n3418), .Z(n3396) );
  AND U3573 ( .A(n3397), .B(n3396), .Z(n3426) );
  NAND U3574 ( .A(b[0]), .B(a[149]), .Z(n3398) );
  XNOR U3575 ( .A(b[1]), .B(n3398), .Z(n3400) );
  NANDN U3576 ( .A(b[0]), .B(a[148]), .Z(n3399) );
  NAND U3577 ( .A(n3400), .B(n3399), .Z(n3425) );
  AND U3578 ( .A(b[3]), .B(a[145]), .Z(n3424) );
  XOR U3579 ( .A(n3425), .B(n3424), .Z(n3427) );
  XOR U3580 ( .A(n3426), .B(n3427), .Z(n3413) );
  NANDN U3581 ( .A(n3402), .B(n3401), .Z(n3406) );
  OR U3582 ( .A(n3404), .B(n3403), .Z(n3405) );
  AND U3583 ( .A(n3406), .B(n3405), .Z(n3412) );
  XOR U3584 ( .A(n3413), .B(n3412), .Z(n3415) );
  XOR U3585 ( .A(n3414), .B(n3415), .Z(n3430) );
  XNOR U3586 ( .A(n3430), .B(sreg[401]), .Z(n3432) );
  NANDN U3587 ( .A(n3407), .B(sreg[400]), .Z(n3411) );
  NAND U3588 ( .A(n3409), .B(n3408), .Z(n3410) );
  NAND U3589 ( .A(n3411), .B(n3410), .Z(n3431) );
  XOR U3590 ( .A(n3432), .B(n3431), .Z(c[401]) );
  NANDN U3591 ( .A(n3413), .B(n3412), .Z(n3417) );
  OR U3592 ( .A(n3415), .B(n3414), .Z(n3416) );
  AND U3593 ( .A(n3417), .B(n3416), .Z(n3437) );
  NAND U3594 ( .A(n31), .B(n3418), .Z(n3420) );
  XOR U3595 ( .A(b[3]), .B(a[148]), .Z(n3441) );
  NAND U3596 ( .A(n5811), .B(n3441), .Z(n3419) );
  AND U3597 ( .A(n3420), .B(n3419), .Z(n3449) );
  NAND U3598 ( .A(b[0]), .B(a[150]), .Z(n3421) );
  XNOR U3599 ( .A(b[1]), .B(n3421), .Z(n3423) );
  NANDN U3600 ( .A(b[0]), .B(a[149]), .Z(n3422) );
  NAND U3601 ( .A(n3423), .B(n3422), .Z(n3448) );
  AND U3602 ( .A(b[3]), .B(a[146]), .Z(n3447) );
  XOR U3603 ( .A(n3448), .B(n3447), .Z(n3450) );
  XOR U3604 ( .A(n3449), .B(n3450), .Z(n3436) );
  NANDN U3605 ( .A(n3425), .B(n3424), .Z(n3429) );
  OR U3606 ( .A(n3427), .B(n3426), .Z(n3428) );
  AND U3607 ( .A(n3429), .B(n3428), .Z(n3435) );
  XOR U3608 ( .A(n3436), .B(n3435), .Z(n3438) );
  XOR U3609 ( .A(n3437), .B(n3438), .Z(n3453) );
  XNOR U3610 ( .A(n3453), .B(sreg[402]), .Z(n3455) );
  NANDN U3611 ( .A(n3430), .B(sreg[401]), .Z(n3434) );
  NAND U3612 ( .A(n3432), .B(n3431), .Z(n3433) );
  NAND U3613 ( .A(n3434), .B(n3433), .Z(n3454) );
  XOR U3614 ( .A(n3455), .B(n3454), .Z(c[402]) );
  NANDN U3615 ( .A(n3436), .B(n3435), .Z(n3440) );
  OR U3616 ( .A(n3438), .B(n3437), .Z(n3439) );
  AND U3617 ( .A(n3440), .B(n3439), .Z(n3460) );
  NAND U3618 ( .A(n31), .B(n3441), .Z(n3443) );
  XOR U3619 ( .A(b[3]), .B(a[149]), .Z(n3464) );
  NAND U3620 ( .A(n5811), .B(n3464), .Z(n3442) );
  AND U3621 ( .A(n3443), .B(n3442), .Z(n3472) );
  NAND U3622 ( .A(b[0]), .B(a[151]), .Z(n3444) );
  XNOR U3623 ( .A(b[1]), .B(n3444), .Z(n3446) );
  NANDN U3624 ( .A(b[0]), .B(a[150]), .Z(n3445) );
  NAND U3625 ( .A(n3446), .B(n3445), .Z(n3471) );
  AND U3626 ( .A(b[3]), .B(a[147]), .Z(n3470) );
  XOR U3627 ( .A(n3471), .B(n3470), .Z(n3473) );
  XOR U3628 ( .A(n3472), .B(n3473), .Z(n3459) );
  NANDN U3629 ( .A(n3448), .B(n3447), .Z(n3452) );
  OR U3630 ( .A(n3450), .B(n3449), .Z(n3451) );
  AND U3631 ( .A(n3452), .B(n3451), .Z(n3458) );
  XOR U3632 ( .A(n3459), .B(n3458), .Z(n3461) );
  XOR U3633 ( .A(n3460), .B(n3461), .Z(n3476) );
  XNOR U3634 ( .A(n3476), .B(sreg[403]), .Z(n3478) );
  NANDN U3635 ( .A(n3453), .B(sreg[402]), .Z(n3457) );
  NAND U3636 ( .A(n3455), .B(n3454), .Z(n3456) );
  NAND U3637 ( .A(n3457), .B(n3456), .Z(n3477) );
  XOR U3638 ( .A(n3478), .B(n3477), .Z(c[403]) );
  NANDN U3639 ( .A(n3459), .B(n3458), .Z(n3463) );
  OR U3640 ( .A(n3461), .B(n3460), .Z(n3462) );
  AND U3641 ( .A(n3463), .B(n3462), .Z(n3483) );
  NAND U3642 ( .A(n31), .B(n3464), .Z(n3466) );
  XOR U3643 ( .A(b[3]), .B(a[150]), .Z(n3487) );
  NAND U3644 ( .A(n5811), .B(n3487), .Z(n3465) );
  AND U3645 ( .A(n3466), .B(n3465), .Z(n3495) );
  NAND U3646 ( .A(b[0]), .B(a[152]), .Z(n3467) );
  XNOR U3647 ( .A(b[1]), .B(n3467), .Z(n3469) );
  NANDN U3648 ( .A(b[0]), .B(a[151]), .Z(n3468) );
  NAND U3649 ( .A(n3469), .B(n3468), .Z(n3494) );
  AND U3650 ( .A(b[3]), .B(a[148]), .Z(n3493) );
  XOR U3651 ( .A(n3494), .B(n3493), .Z(n3496) );
  XOR U3652 ( .A(n3495), .B(n3496), .Z(n3482) );
  NANDN U3653 ( .A(n3471), .B(n3470), .Z(n3475) );
  OR U3654 ( .A(n3473), .B(n3472), .Z(n3474) );
  AND U3655 ( .A(n3475), .B(n3474), .Z(n3481) );
  XOR U3656 ( .A(n3482), .B(n3481), .Z(n3484) );
  XOR U3657 ( .A(n3483), .B(n3484), .Z(n3499) );
  XNOR U3658 ( .A(n3499), .B(sreg[404]), .Z(n3501) );
  NANDN U3659 ( .A(n3476), .B(sreg[403]), .Z(n3480) );
  NAND U3660 ( .A(n3478), .B(n3477), .Z(n3479) );
  NAND U3661 ( .A(n3480), .B(n3479), .Z(n3500) );
  XOR U3662 ( .A(n3501), .B(n3500), .Z(c[404]) );
  NANDN U3663 ( .A(n3482), .B(n3481), .Z(n3486) );
  OR U3664 ( .A(n3484), .B(n3483), .Z(n3485) );
  AND U3665 ( .A(n3486), .B(n3485), .Z(n3506) );
  NAND U3666 ( .A(n31), .B(n3487), .Z(n3489) );
  XOR U3667 ( .A(b[3]), .B(a[151]), .Z(n3510) );
  NAND U3668 ( .A(n5811), .B(n3510), .Z(n3488) );
  AND U3669 ( .A(n3489), .B(n3488), .Z(n3518) );
  NAND U3670 ( .A(b[0]), .B(a[153]), .Z(n3490) );
  XNOR U3671 ( .A(b[1]), .B(n3490), .Z(n3492) );
  NANDN U3672 ( .A(b[0]), .B(a[152]), .Z(n3491) );
  NAND U3673 ( .A(n3492), .B(n3491), .Z(n3517) );
  AND U3674 ( .A(b[3]), .B(a[149]), .Z(n3516) );
  XOR U3675 ( .A(n3517), .B(n3516), .Z(n3519) );
  XOR U3676 ( .A(n3518), .B(n3519), .Z(n3505) );
  NANDN U3677 ( .A(n3494), .B(n3493), .Z(n3498) );
  OR U3678 ( .A(n3496), .B(n3495), .Z(n3497) );
  AND U3679 ( .A(n3498), .B(n3497), .Z(n3504) );
  XOR U3680 ( .A(n3505), .B(n3504), .Z(n3507) );
  XOR U3681 ( .A(n3506), .B(n3507), .Z(n3522) );
  XNOR U3682 ( .A(n3522), .B(sreg[405]), .Z(n3524) );
  NANDN U3683 ( .A(n3499), .B(sreg[404]), .Z(n3503) );
  NAND U3684 ( .A(n3501), .B(n3500), .Z(n3502) );
  NAND U3685 ( .A(n3503), .B(n3502), .Z(n3523) );
  XOR U3686 ( .A(n3524), .B(n3523), .Z(c[405]) );
  NANDN U3687 ( .A(n3505), .B(n3504), .Z(n3509) );
  OR U3688 ( .A(n3507), .B(n3506), .Z(n3508) );
  AND U3689 ( .A(n3509), .B(n3508), .Z(n3529) );
  NAND U3690 ( .A(n31), .B(n3510), .Z(n3512) );
  XOR U3691 ( .A(b[3]), .B(a[152]), .Z(n3533) );
  NAND U3692 ( .A(n5811), .B(n3533), .Z(n3511) );
  AND U3693 ( .A(n3512), .B(n3511), .Z(n3541) );
  NAND U3694 ( .A(b[0]), .B(a[154]), .Z(n3513) );
  XNOR U3695 ( .A(b[1]), .B(n3513), .Z(n3515) );
  NANDN U3696 ( .A(b[0]), .B(a[153]), .Z(n3514) );
  NAND U3697 ( .A(n3515), .B(n3514), .Z(n3540) );
  AND U3698 ( .A(b[3]), .B(a[150]), .Z(n3539) );
  XOR U3699 ( .A(n3540), .B(n3539), .Z(n3542) );
  XOR U3700 ( .A(n3541), .B(n3542), .Z(n3528) );
  NANDN U3701 ( .A(n3517), .B(n3516), .Z(n3521) );
  OR U3702 ( .A(n3519), .B(n3518), .Z(n3520) );
  AND U3703 ( .A(n3521), .B(n3520), .Z(n3527) );
  XOR U3704 ( .A(n3528), .B(n3527), .Z(n3530) );
  XOR U3705 ( .A(n3529), .B(n3530), .Z(n3545) );
  XNOR U3706 ( .A(n3545), .B(sreg[406]), .Z(n3547) );
  NANDN U3707 ( .A(n3522), .B(sreg[405]), .Z(n3526) );
  NAND U3708 ( .A(n3524), .B(n3523), .Z(n3525) );
  NAND U3709 ( .A(n3526), .B(n3525), .Z(n3546) );
  XOR U3710 ( .A(n3547), .B(n3546), .Z(c[406]) );
  NANDN U3711 ( .A(n3528), .B(n3527), .Z(n3532) );
  OR U3712 ( .A(n3530), .B(n3529), .Z(n3531) );
  AND U3713 ( .A(n3532), .B(n3531), .Z(n3552) );
  NAND U3714 ( .A(n31), .B(n3533), .Z(n3535) );
  XOR U3715 ( .A(b[3]), .B(a[153]), .Z(n3556) );
  NAND U3716 ( .A(n5811), .B(n3556), .Z(n3534) );
  AND U3717 ( .A(n3535), .B(n3534), .Z(n3564) );
  AND U3718 ( .A(b[3]), .B(a[151]), .Z(n3562) );
  NAND U3719 ( .A(b[0]), .B(a[155]), .Z(n3536) );
  XNOR U3720 ( .A(b[1]), .B(n3536), .Z(n3538) );
  NANDN U3721 ( .A(b[0]), .B(a[154]), .Z(n3537) );
  NAND U3722 ( .A(n3538), .B(n3537), .Z(n3563) );
  XOR U3723 ( .A(n3562), .B(n3563), .Z(n3565) );
  XOR U3724 ( .A(n3564), .B(n3565), .Z(n3551) );
  NANDN U3725 ( .A(n3540), .B(n3539), .Z(n3544) );
  OR U3726 ( .A(n3542), .B(n3541), .Z(n3543) );
  AND U3727 ( .A(n3544), .B(n3543), .Z(n3550) );
  XOR U3728 ( .A(n3551), .B(n3550), .Z(n3553) );
  XOR U3729 ( .A(n3552), .B(n3553), .Z(n3568) );
  XNOR U3730 ( .A(n3568), .B(sreg[407]), .Z(n3570) );
  NANDN U3731 ( .A(n3545), .B(sreg[406]), .Z(n3549) );
  NAND U3732 ( .A(n3547), .B(n3546), .Z(n3548) );
  NAND U3733 ( .A(n3549), .B(n3548), .Z(n3569) );
  XOR U3734 ( .A(n3570), .B(n3569), .Z(c[407]) );
  NANDN U3735 ( .A(n3551), .B(n3550), .Z(n3555) );
  OR U3736 ( .A(n3553), .B(n3552), .Z(n3554) );
  AND U3737 ( .A(n3555), .B(n3554), .Z(n3575) );
  NAND U3738 ( .A(n31), .B(n3556), .Z(n3558) );
  XOR U3739 ( .A(b[3]), .B(a[154]), .Z(n3579) );
  NAND U3740 ( .A(n5811), .B(n3579), .Z(n3557) );
  AND U3741 ( .A(n3558), .B(n3557), .Z(n3587) );
  NAND U3742 ( .A(b[0]), .B(a[156]), .Z(n3559) );
  XNOR U3743 ( .A(b[1]), .B(n3559), .Z(n3561) );
  NANDN U3744 ( .A(b[0]), .B(a[155]), .Z(n3560) );
  NAND U3745 ( .A(n3561), .B(n3560), .Z(n3586) );
  AND U3746 ( .A(b[3]), .B(a[152]), .Z(n3585) );
  XOR U3747 ( .A(n3586), .B(n3585), .Z(n3588) );
  XOR U3748 ( .A(n3587), .B(n3588), .Z(n3574) );
  NANDN U3749 ( .A(n3563), .B(n3562), .Z(n3567) );
  OR U3750 ( .A(n3565), .B(n3564), .Z(n3566) );
  AND U3751 ( .A(n3567), .B(n3566), .Z(n3573) );
  XOR U3752 ( .A(n3574), .B(n3573), .Z(n3576) );
  XOR U3753 ( .A(n3575), .B(n3576), .Z(n3591) );
  XNOR U3754 ( .A(n3591), .B(sreg[408]), .Z(n3593) );
  NANDN U3755 ( .A(n3568), .B(sreg[407]), .Z(n3572) );
  NAND U3756 ( .A(n3570), .B(n3569), .Z(n3571) );
  NAND U3757 ( .A(n3572), .B(n3571), .Z(n3592) );
  XOR U3758 ( .A(n3593), .B(n3592), .Z(c[408]) );
  NANDN U3759 ( .A(n3574), .B(n3573), .Z(n3578) );
  OR U3760 ( .A(n3576), .B(n3575), .Z(n3577) );
  AND U3761 ( .A(n3578), .B(n3577), .Z(n3598) );
  NAND U3762 ( .A(n31), .B(n3579), .Z(n3581) );
  XOR U3763 ( .A(b[3]), .B(a[155]), .Z(n3602) );
  NAND U3764 ( .A(n5811), .B(n3602), .Z(n3580) );
  AND U3765 ( .A(n3581), .B(n3580), .Z(n3610) );
  NAND U3766 ( .A(b[0]), .B(a[157]), .Z(n3582) );
  XNOR U3767 ( .A(b[1]), .B(n3582), .Z(n3584) );
  NANDN U3768 ( .A(b[0]), .B(a[156]), .Z(n3583) );
  NAND U3769 ( .A(n3584), .B(n3583), .Z(n3609) );
  AND U3770 ( .A(b[3]), .B(a[153]), .Z(n3608) );
  XOR U3771 ( .A(n3609), .B(n3608), .Z(n3611) );
  XOR U3772 ( .A(n3610), .B(n3611), .Z(n3597) );
  NANDN U3773 ( .A(n3586), .B(n3585), .Z(n3590) );
  OR U3774 ( .A(n3588), .B(n3587), .Z(n3589) );
  AND U3775 ( .A(n3590), .B(n3589), .Z(n3596) );
  XOR U3776 ( .A(n3597), .B(n3596), .Z(n3599) );
  XOR U3777 ( .A(n3598), .B(n3599), .Z(n3614) );
  XNOR U3778 ( .A(n3614), .B(sreg[409]), .Z(n3616) );
  NANDN U3779 ( .A(n3591), .B(sreg[408]), .Z(n3595) );
  NAND U3780 ( .A(n3593), .B(n3592), .Z(n3594) );
  NAND U3781 ( .A(n3595), .B(n3594), .Z(n3615) );
  XOR U3782 ( .A(n3616), .B(n3615), .Z(c[409]) );
  NANDN U3783 ( .A(n3597), .B(n3596), .Z(n3601) );
  OR U3784 ( .A(n3599), .B(n3598), .Z(n3600) );
  AND U3785 ( .A(n3601), .B(n3600), .Z(n3621) );
  NAND U3786 ( .A(n31), .B(n3602), .Z(n3604) );
  XOR U3787 ( .A(b[3]), .B(a[156]), .Z(n3625) );
  NAND U3788 ( .A(n5811), .B(n3625), .Z(n3603) );
  AND U3789 ( .A(n3604), .B(n3603), .Z(n3633) );
  NAND U3790 ( .A(b[0]), .B(a[158]), .Z(n3605) );
  XNOR U3791 ( .A(b[1]), .B(n3605), .Z(n3607) );
  NANDN U3792 ( .A(b[0]), .B(a[157]), .Z(n3606) );
  NAND U3793 ( .A(n3607), .B(n3606), .Z(n3632) );
  AND U3794 ( .A(b[3]), .B(a[154]), .Z(n3631) );
  XOR U3795 ( .A(n3632), .B(n3631), .Z(n3634) );
  XOR U3796 ( .A(n3633), .B(n3634), .Z(n3620) );
  NANDN U3797 ( .A(n3609), .B(n3608), .Z(n3613) );
  OR U3798 ( .A(n3611), .B(n3610), .Z(n3612) );
  AND U3799 ( .A(n3613), .B(n3612), .Z(n3619) );
  XOR U3800 ( .A(n3620), .B(n3619), .Z(n3622) );
  XOR U3801 ( .A(n3621), .B(n3622), .Z(n3637) );
  XNOR U3802 ( .A(n3637), .B(sreg[410]), .Z(n3639) );
  NANDN U3803 ( .A(n3614), .B(sreg[409]), .Z(n3618) );
  NAND U3804 ( .A(n3616), .B(n3615), .Z(n3617) );
  NAND U3805 ( .A(n3618), .B(n3617), .Z(n3638) );
  XOR U3806 ( .A(n3639), .B(n3638), .Z(c[410]) );
  NANDN U3807 ( .A(n3620), .B(n3619), .Z(n3624) );
  OR U3808 ( .A(n3622), .B(n3621), .Z(n3623) );
  AND U3809 ( .A(n3624), .B(n3623), .Z(n3644) );
  NAND U3810 ( .A(n31), .B(n3625), .Z(n3627) );
  XOR U3811 ( .A(b[3]), .B(a[157]), .Z(n3648) );
  NAND U3812 ( .A(n5811), .B(n3648), .Z(n3626) );
  AND U3813 ( .A(n3627), .B(n3626), .Z(n3656) );
  AND U3814 ( .A(b[3]), .B(a[155]), .Z(n3654) );
  NAND U3815 ( .A(b[0]), .B(a[159]), .Z(n3628) );
  XNOR U3816 ( .A(b[1]), .B(n3628), .Z(n3630) );
  NANDN U3817 ( .A(b[0]), .B(a[158]), .Z(n3629) );
  NAND U3818 ( .A(n3630), .B(n3629), .Z(n3655) );
  XOR U3819 ( .A(n3654), .B(n3655), .Z(n3657) );
  XOR U3820 ( .A(n3656), .B(n3657), .Z(n3643) );
  NANDN U3821 ( .A(n3632), .B(n3631), .Z(n3636) );
  OR U3822 ( .A(n3634), .B(n3633), .Z(n3635) );
  AND U3823 ( .A(n3636), .B(n3635), .Z(n3642) );
  XOR U3824 ( .A(n3643), .B(n3642), .Z(n3645) );
  XOR U3825 ( .A(n3644), .B(n3645), .Z(n3660) );
  XNOR U3826 ( .A(n3660), .B(sreg[411]), .Z(n3662) );
  NANDN U3827 ( .A(n3637), .B(sreg[410]), .Z(n3641) );
  NAND U3828 ( .A(n3639), .B(n3638), .Z(n3640) );
  NAND U3829 ( .A(n3641), .B(n3640), .Z(n3661) );
  XOR U3830 ( .A(n3662), .B(n3661), .Z(c[411]) );
  NANDN U3831 ( .A(n3643), .B(n3642), .Z(n3647) );
  OR U3832 ( .A(n3645), .B(n3644), .Z(n3646) );
  AND U3833 ( .A(n3647), .B(n3646), .Z(n3667) );
  NAND U3834 ( .A(n31), .B(n3648), .Z(n3650) );
  XOR U3835 ( .A(b[3]), .B(a[158]), .Z(n3671) );
  NAND U3836 ( .A(n5811), .B(n3671), .Z(n3649) );
  AND U3837 ( .A(n3650), .B(n3649), .Z(n3679) );
  NAND U3838 ( .A(b[0]), .B(a[160]), .Z(n3651) );
  XNOR U3839 ( .A(b[1]), .B(n3651), .Z(n3653) );
  NANDN U3840 ( .A(b[0]), .B(a[159]), .Z(n3652) );
  NAND U3841 ( .A(n3653), .B(n3652), .Z(n3678) );
  AND U3842 ( .A(b[3]), .B(a[156]), .Z(n3677) );
  XOR U3843 ( .A(n3678), .B(n3677), .Z(n3680) );
  XOR U3844 ( .A(n3679), .B(n3680), .Z(n3666) );
  NANDN U3845 ( .A(n3655), .B(n3654), .Z(n3659) );
  OR U3846 ( .A(n3657), .B(n3656), .Z(n3658) );
  AND U3847 ( .A(n3659), .B(n3658), .Z(n3665) );
  XOR U3848 ( .A(n3666), .B(n3665), .Z(n3668) );
  XOR U3849 ( .A(n3667), .B(n3668), .Z(n3683) );
  XNOR U3850 ( .A(n3683), .B(sreg[412]), .Z(n3685) );
  NANDN U3851 ( .A(n3660), .B(sreg[411]), .Z(n3664) );
  NAND U3852 ( .A(n3662), .B(n3661), .Z(n3663) );
  NAND U3853 ( .A(n3664), .B(n3663), .Z(n3684) );
  XOR U3854 ( .A(n3685), .B(n3684), .Z(c[412]) );
  NANDN U3855 ( .A(n3666), .B(n3665), .Z(n3670) );
  OR U3856 ( .A(n3668), .B(n3667), .Z(n3669) );
  AND U3857 ( .A(n3670), .B(n3669), .Z(n3690) );
  NAND U3858 ( .A(n31), .B(n3671), .Z(n3673) );
  XOR U3859 ( .A(b[3]), .B(a[159]), .Z(n3694) );
  NAND U3860 ( .A(n5811), .B(n3694), .Z(n3672) );
  AND U3861 ( .A(n3673), .B(n3672), .Z(n3702) );
  NAND U3862 ( .A(b[0]), .B(a[161]), .Z(n3674) );
  XNOR U3863 ( .A(b[1]), .B(n3674), .Z(n3676) );
  NANDN U3864 ( .A(b[0]), .B(a[160]), .Z(n3675) );
  NAND U3865 ( .A(n3676), .B(n3675), .Z(n3701) );
  AND U3866 ( .A(b[3]), .B(a[157]), .Z(n3700) );
  XOR U3867 ( .A(n3701), .B(n3700), .Z(n3703) );
  XOR U3868 ( .A(n3702), .B(n3703), .Z(n3689) );
  NANDN U3869 ( .A(n3678), .B(n3677), .Z(n3682) );
  OR U3870 ( .A(n3680), .B(n3679), .Z(n3681) );
  AND U3871 ( .A(n3682), .B(n3681), .Z(n3688) );
  XOR U3872 ( .A(n3689), .B(n3688), .Z(n3691) );
  XOR U3873 ( .A(n3690), .B(n3691), .Z(n3706) );
  XNOR U3874 ( .A(n3706), .B(sreg[413]), .Z(n3708) );
  NANDN U3875 ( .A(n3683), .B(sreg[412]), .Z(n3687) );
  NAND U3876 ( .A(n3685), .B(n3684), .Z(n3686) );
  NAND U3877 ( .A(n3687), .B(n3686), .Z(n3707) );
  XOR U3878 ( .A(n3708), .B(n3707), .Z(c[413]) );
  NANDN U3879 ( .A(n3689), .B(n3688), .Z(n3693) );
  OR U3880 ( .A(n3691), .B(n3690), .Z(n3692) );
  AND U3881 ( .A(n3693), .B(n3692), .Z(n3713) );
  NAND U3882 ( .A(n31), .B(n3694), .Z(n3696) );
  XOR U3883 ( .A(b[3]), .B(a[160]), .Z(n3717) );
  NAND U3884 ( .A(n5811), .B(n3717), .Z(n3695) );
  AND U3885 ( .A(n3696), .B(n3695), .Z(n3725) );
  NAND U3886 ( .A(b[0]), .B(a[162]), .Z(n3697) );
  XNOR U3887 ( .A(b[1]), .B(n3697), .Z(n3699) );
  NANDN U3888 ( .A(b[0]), .B(a[161]), .Z(n3698) );
  NAND U3889 ( .A(n3699), .B(n3698), .Z(n3724) );
  AND U3890 ( .A(b[3]), .B(a[158]), .Z(n3723) );
  XOR U3891 ( .A(n3724), .B(n3723), .Z(n3726) );
  XOR U3892 ( .A(n3725), .B(n3726), .Z(n3712) );
  NANDN U3893 ( .A(n3701), .B(n3700), .Z(n3705) );
  OR U3894 ( .A(n3703), .B(n3702), .Z(n3704) );
  AND U3895 ( .A(n3705), .B(n3704), .Z(n3711) );
  XOR U3896 ( .A(n3712), .B(n3711), .Z(n3714) );
  XOR U3897 ( .A(n3713), .B(n3714), .Z(n3729) );
  XNOR U3898 ( .A(n3729), .B(sreg[414]), .Z(n3731) );
  NANDN U3899 ( .A(n3706), .B(sreg[413]), .Z(n3710) );
  NAND U3900 ( .A(n3708), .B(n3707), .Z(n3709) );
  NAND U3901 ( .A(n3710), .B(n3709), .Z(n3730) );
  XOR U3902 ( .A(n3731), .B(n3730), .Z(c[414]) );
  NANDN U3903 ( .A(n3712), .B(n3711), .Z(n3716) );
  OR U3904 ( .A(n3714), .B(n3713), .Z(n3715) );
  AND U3905 ( .A(n3716), .B(n3715), .Z(n3736) );
  NAND U3906 ( .A(n31), .B(n3717), .Z(n3719) );
  XOR U3907 ( .A(b[3]), .B(a[161]), .Z(n3740) );
  NAND U3908 ( .A(n5811), .B(n3740), .Z(n3718) );
  AND U3909 ( .A(n3719), .B(n3718), .Z(n3748) );
  NAND U3910 ( .A(b[0]), .B(a[163]), .Z(n3720) );
  XNOR U3911 ( .A(b[1]), .B(n3720), .Z(n3722) );
  NANDN U3912 ( .A(b[0]), .B(a[162]), .Z(n3721) );
  NAND U3913 ( .A(n3722), .B(n3721), .Z(n3747) );
  AND U3914 ( .A(b[3]), .B(a[159]), .Z(n3746) );
  XOR U3915 ( .A(n3747), .B(n3746), .Z(n3749) );
  XOR U3916 ( .A(n3748), .B(n3749), .Z(n3735) );
  NANDN U3917 ( .A(n3724), .B(n3723), .Z(n3728) );
  OR U3918 ( .A(n3726), .B(n3725), .Z(n3727) );
  AND U3919 ( .A(n3728), .B(n3727), .Z(n3734) );
  XOR U3920 ( .A(n3735), .B(n3734), .Z(n3737) );
  XOR U3921 ( .A(n3736), .B(n3737), .Z(n3752) );
  XNOR U3922 ( .A(n3752), .B(sreg[415]), .Z(n3754) );
  NANDN U3923 ( .A(n3729), .B(sreg[414]), .Z(n3733) );
  NAND U3924 ( .A(n3731), .B(n3730), .Z(n3732) );
  NAND U3925 ( .A(n3733), .B(n3732), .Z(n3753) );
  XOR U3926 ( .A(n3754), .B(n3753), .Z(c[415]) );
  NANDN U3927 ( .A(n3735), .B(n3734), .Z(n3739) );
  OR U3928 ( .A(n3737), .B(n3736), .Z(n3738) );
  AND U3929 ( .A(n3739), .B(n3738), .Z(n3759) );
  NAND U3930 ( .A(n31), .B(n3740), .Z(n3742) );
  XOR U3931 ( .A(b[3]), .B(a[162]), .Z(n3763) );
  NAND U3932 ( .A(n5811), .B(n3763), .Z(n3741) );
  AND U3933 ( .A(n3742), .B(n3741), .Z(n3771) );
  NAND U3934 ( .A(b[0]), .B(a[164]), .Z(n3743) );
  XNOR U3935 ( .A(b[1]), .B(n3743), .Z(n3745) );
  NANDN U3936 ( .A(b[0]), .B(a[163]), .Z(n3744) );
  NAND U3937 ( .A(n3745), .B(n3744), .Z(n3770) );
  AND U3938 ( .A(b[3]), .B(a[160]), .Z(n3769) );
  XOR U3939 ( .A(n3770), .B(n3769), .Z(n3772) );
  XOR U3940 ( .A(n3771), .B(n3772), .Z(n3758) );
  NANDN U3941 ( .A(n3747), .B(n3746), .Z(n3751) );
  OR U3942 ( .A(n3749), .B(n3748), .Z(n3750) );
  AND U3943 ( .A(n3751), .B(n3750), .Z(n3757) );
  XOR U3944 ( .A(n3758), .B(n3757), .Z(n3760) );
  XOR U3945 ( .A(n3759), .B(n3760), .Z(n3775) );
  XNOR U3946 ( .A(n3775), .B(sreg[416]), .Z(n3777) );
  NANDN U3947 ( .A(n3752), .B(sreg[415]), .Z(n3756) );
  NAND U3948 ( .A(n3754), .B(n3753), .Z(n3755) );
  NAND U3949 ( .A(n3756), .B(n3755), .Z(n3776) );
  XOR U3950 ( .A(n3777), .B(n3776), .Z(c[416]) );
  NANDN U3951 ( .A(n3758), .B(n3757), .Z(n3762) );
  OR U3952 ( .A(n3760), .B(n3759), .Z(n3761) );
  AND U3953 ( .A(n3762), .B(n3761), .Z(n3782) );
  NAND U3954 ( .A(n31), .B(n3763), .Z(n3765) );
  XOR U3955 ( .A(b[3]), .B(a[163]), .Z(n3786) );
  NAND U3956 ( .A(n5811), .B(n3786), .Z(n3764) );
  AND U3957 ( .A(n3765), .B(n3764), .Z(n3794) );
  AND U3958 ( .A(b[3]), .B(a[161]), .Z(n3792) );
  NAND U3959 ( .A(b[0]), .B(a[165]), .Z(n3766) );
  XNOR U3960 ( .A(b[1]), .B(n3766), .Z(n3768) );
  NANDN U3961 ( .A(b[0]), .B(a[164]), .Z(n3767) );
  NAND U3962 ( .A(n3768), .B(n3767), .Z(n3793) );
  XOR U3963 ( .A(n3792), .B(n3793), .Z(n3795) );
  XOR U3964 ( .A(n3794), .B(n3795), .Z(n3781) );
  NANDN U3965 ( .A(n3770), .B(n3769), .Z(n3774) );
  OR U3966 ( .A(n3772), .B(n3771), .Z(n3773) );
  AND U3967 ( .A(n3774), .B(n3773), .Z(n3780) );
  XOR U3968 ( .A(n3781), .B(n3780), .Z(n3783) );
  XOR U3969 ( .A(n3782), .B(n3783), .Z(n3798) );
  XNOR U3970 ( .A(n3798), .B(sreg[417]), .Z(n3800) );
  NANDN U3971 ( .A(n3775), .B(sreg[416]), .Z(n3779) );
  NAND U3972 ( .A(n3777), .B(n3776), .Z(n3778) );
  NAND U3973 ( .A(n3779), .B(n3778), .Z(n3799) );
  XOR U3974 ( .A(n3800), .B(n3799), .Z(c[417]) );
  NANDN U3975 ( .A(n3781), .B(n3780), .Z(n3785) );
  OR U3976 ( .A(n3783), .B(n3782), .Z(n3784) );
  AND U3977 ( .A(n3785), .B(n3784), .Z(n3805) );
  NAND U3978 ( .A(n31), .B(n3786), .Z(n3788) );
  XOR U3979 ( .A(b[3]), .B(a[164]), .Z(n3809) );
  NAND U3980 ( .A(n5811), .B(n3809), .Z(n3787) );
  AND U3981 ( .A(n3788), .B(n3787), .Z(n3817) );
  NAND U3982 ( .A(b[0]), .B(a[166]), .Z(n3789) );
  XNOR U3983 ( .A(b[1]), .B(n3789), .Z(n3791) );
  NANDN U3984 ( .A(b[0]), .B(a[165]), .Z(n3790) );
  NAND U3985 ( .A(n3791), .B(n3790), .Z(n3816) );
  AND U3986 ( .A(b[3]), .B(a[162]), .Z(n3815) );
  XOR U3987 ( .A(n3816), .B(n3815), .Z(n3818) );
  XOR U3988 ( .A(n3817), .B(n3818), .Z(n3804) );
  NANDN U3989 ( .A(n3793), .B(n3792), .Z(n3797) );
  OR U3990 ( .A(n3795), .B(n3794), .Z(n3796) );
  AND U3991 ( .A(n3797), .B(n3796), .Z(n3803) );
  XOR U3992 ( .A(n3804), .B(n3803), .Z(n3806) );
  XOR U3993 ( .A(n3805), .B(n3806), .Z(n3821) );
  XNOR U3994 ( .A(n3821), .B(sreg[418]), .Z(n3823) );
  NANDN U3995 ( .A(n3798), .B(sreg[417]), .Z(n3802) );
  NAND U3996 ( .A(n3800), .B(n3799), .Z(n3801) );
  NAND U3997 ( .A(n3802), .B(n3801), .Z(n3822) );
  XOR U3998 ( .A(n3823), .B(n3822), .Z(c[418]) );
  NANDN U3999 ( .A(n3804), .B(n3803), .Z(n3808) );
  OR U4000 ( .A(n3806), .B(n3805), .Z(n3807) );
  AND U4001 ( .A(n3808), .B(n3807), .Z(n3828) );
  NAND U4002 ( .A(n31), .B(n3809), .Z(n3811) );
  XOR U4003 ( .A(b[3]), .B(a[165]), .Z(n3832) );
  NAND U4004 ( .A(n5811), .B(n3832), .Z(n3810) );
  AND U4005 ( .A(n3811), .B(n3810), .Z(n3840) );
  NAND U4006 ( .A(b[0]), .B(a[167]), .Z(n3812) );
  XNOR U4007 ( .A(b[1]), .B(n3812), .Z(n3814) );
  NANDN U4008 ( .A(b[0]), .B(a[166]), .Z(n3813) );
  NAND U4009 ( .A(n3814), .B(n3813), .Z(n3839) );
  AND U4010 ( .A(b[3]), .B(a[163]), .Z(n3838) );
  XOR U4011 ( .A(n3839), .B(n3838), .Z(n3841) );
  XOR U4012 ( .A(n3840), .B(n3841), .Z(n3827) );
  NANDN U4013 ( .A(n3816), .B(n3815), .Z(n3820) );
  OR U4014 ( .A(n3818), .B(n3817), .Z(n3819) );
  AND U4015 ( .A(n3820), .B(n3819), .Z(n3826) );
  XOR U4016 ( .A(n3827), .B(n3826), .Z(n3829) );
  XOR U4017 ( .A(n3828), .B(n3829), .Z(n3844) );
  XNOR U4018 ( .A(n3844), .B(sreg[419]), .Z(n3846) );
  NANDN U4019 ( .A(n3821), .B(sreg[418]), .Z(n3825) );
  NAND U4020 ( .A(n3823), .B(n3822), .Z(n3824) );
  NAND U4021 ( .A(n3825), .B(n3824), .Z(n3845) );
  XOR U4022 ( .A(n3846), .B(n3845), .Z(c[419]) );
  NANDN U4023 ( .A(n3827), .B(n3826), .Z(n3831) );
  OR U4024 ( .A(n3829), .B(n3828), .Z(n3830) );
  AND U4025 ( .A(n3831), .B(n3830), .Z(n3851) );
  NAND U4026 ( .A(n31), .B(n3832), .Z(n3834) );
  XOR U4027 ( .A(b[3]), .B(a[166]), .Z(n3855) );
  NAND U4028 ( .A(n5811), .B(n3855), .Z(n3833) );
  AND U4029 ( .A(n3834), .B(n3833), .Z(n3863) );
  NAND U4030 ( .A(b[0]), .B(a[168]), .Z(n3835) );
  XNOR U4031 ( .A(b[1]), .B(n3835), .Z(n3837) );
  NANDN U4032 ( .A(b[0]), .B(a[167]), .Z(n3836) );
  NAND U4033 ( .A(n3837), .B(n3836), .Z(n3862) );
  AND U4034 ( .A(b[3]), .B(a[164]), .Z(n3861) );
  XOR U4035 ( .A(n3862), .B(n3861), .Z(n3864) );
  XOR U4036 ( .A(n3863), .B(n3864), .Z(n3850) );
  NANDN U4037 ( .A(n3839), .B(n3838), .Z(n3843) );
  OR U4038 ( .A(n3841), .B(n3840), .Z(n3842) );
  AND U4039 ( .A(n3843), .B(n3842), .Z(n3849) );
  XOR U4040 ( .A(n3850), .B(n3849), .Z(n3852) );
  XOR U4041 ( .A(n3851), .B(n3852), .Z(n3867) );
  XNOR U4042 ( .A(n3867), .B(sreg[420]), .Z(n3869) );
  NANDN U4043 ( .A(n3844), .B(sreg[419]), .Z(n3848) );
  NAND U4044 ( .A(n3846), .B(n3845), .Z(n3847) );
  NAND U4045 ( .A(n3848), .B(n3847), .Z(n3868) );
  XOR U4046 ( .A(n3869), .B(n3868), .Z(c[420]) );
  NANDN U4047 ( .A(n3850), .B(n3849), .Z(n3854) );
  OR U4048 ( .A(n3852), .B(n3851), .Z(n3853) );
  AND U4049 ( .A(n3854), .B(n3853), .Z(n3874) );
  NAND U4050 ( .A(n31), .B(n3855), .Z(n3857) );
  XOR U4051 ( .A(b[3]), .B(a[167]), .Z(n3878) );
  NAND U4052 ( .A(n5811), .B(n3878), .Z(n3856) );
  AND U4053 ( .A(n3857), .B(n3856), .Z(n3886) );
  NAND U4054 ( .A(b[0]), .B(a[169]), .Z(n3858) );
  XNOR U4055 ( .A(b[1]), .B(n3858), .Z(n3860) );
  NANDN U4056 ( .A(b[0]), .B(a[168]), .Z(n3859) );
  NAND U4057 ( .A(n3860), .B(n3859), .Z(n3885) );
  AND U4058 ( .A(b[3]), .B(a[165]), .Z(n3884) );
  XOR U4059 ( .A(n3885), .B(n3884), .Z(n3887) );
  XOR U4060 ( .A(n3886), .B(n3887), .Z(n3873) );
  NANDN U4061 ( .A(n3862), .B(n3861), .Z(n3866) );
  OR U4062 ( .A(n3864), .B(n3863), .Z(n3865) );
  AND U4063 ( .A(n3866), .B(n3865), .Z(n3872) );
  XOR U4064 ( .A(n3873), .B(n3872), .Z(n3875) );
  XOR U4065 ( .A(n3874), .B(n3875), .Z(n3890) );
  XNOR U4066 ( .A(n3890), .B(sreg[421]), .Z(n3892) );
  NANDN U4067 ( .A(n3867), .B(sreg[420]), .Z(n3871) );
  NAND U4068 ( .A(n3869), .B(n3868), .Z(n3870) );
  NAND U4069 ( .A(n3871), .B(n3870), .Z(n3891) );
  XOR U4070 ( .A(n3892), .B(n3891), .Z(c[421]) );
  NANDN U4071 ( .A(n3873), .B(n3872), .Z(n3877) );
  OR U4072 ( .A(n3875), .B(n3874), .Z(n3876) );
  AND U4073 ( .A(n3877), .B(n3876), .Z(n3897) );
  NAND U4074 ( .A(n31), .B(n3878), .Z(n3880) );
  XOR U4075 ( .A(b[3]), .B(a[168]), .Z(n3901) );
  NAND U4076 ( .A(n5811), .B(n3901), .Z(n3879) );
  AND U4077 ( .A(n3880), .B(n3879), .Z(n3909) );
  NAND U4078 ( .A(b[0]), .B(a[170]), .Z(n3881) );
  XNOR U4079 ( .A(b[1]), .B(n3881), .Z(n3883) );
  NANDN U4080 ( .A(b[0]), .B(a[169]), .Z(n3882) );
  NAND U4081 ( .A(n3883), .B(n3882), .Z(n3908) );
  AND U4082 ( .A(b[3]), .B(a[166]), .Z(n3907) );
  XOR U4083 ( .A(n3908), .B(n3907), .Z(n3910) );
  XOR U4084 ( .A(n3909), .B(n3910), .Z(n3896) );
  NANDN U4085 ( .A(n3885), .B(n3884), .Z(n3889) );
  OR U4086 ( .A(n3887), .B(n3886), .Z(n3888) );
  AND U4087 ( .A(n3889), .B(n3888), .Z(n3895) );
  XOR U4088 ( .A(n3896), .B(n3895), .Z(n3898) );
  XOR U4089 ( .A(n3897), .B(n3898), .Z(n3913) );
  XNOR U4090 ( .A(n3913), .B(sreg[422]), .Z(n3915) );
  NANDN U4091 ( .A(n3890), .B(sreg[421]), .Z(n3894) );
  NAND U4092 ( .A(n3892), .B(n3891), .Z(n3893) );
  NAND U4093 ( .A(n3894), .B(n3893), .Z(n3914) );
  XOR U4094 ( .A(n3915), .B(n3914), .Z(c[422]) );
  NANDN U4095 ( .A(n3896), .B(n3895), .Z(n3900) );
  OR U4096 ( .A(n3898), .B(n3897), .Z(n3899) );
  AND U4097 ( .A(n3900), .B(n3899), .Z(n3920) );
  NAND U4098 ( .A(n31), .B(n3901), .Z(n3903) );
  XOR U4099 ( .A(b[3]), .B(a[169]), .Z(n3924) );
  NAND U4100 ( .A(n5811), .B(n3924), .Z(n3902) );
  AND U4101 ( .A(n3903), .B(n3902), .Z(n3932) );
  AND U4102 ( .A(b[3]), .B(a[167]), .Z(n3930) );
  NAND U4103 ( .A(b[0]), .B(a[171]), .Z(n3904) );
  XNOR U4104 ( .A(b[1]), .B(n3904), .Z(n3906) );
  NANDN U4105 ( .A(b[0]), .B(a[170]), .Z(n3905) );
  NAND U4106 ( .A(n3906), .B(n3905), .Z(n3931) );
  XOR U4107 ( .A(n3930), .B(n3931), .Z(n3933) );
  XOR U4108 ( .A(n3932), .B(n3933), .Z(n3919) );
  NANDN U4109 ( .A(n3908), .B(n3907), .Z(n3912) );
  OR U4110 ( .A(n3910), .B(n3909), .Z(n3911) );
  AND U4111 ( .A(n3912), .B(n3911), .Z(n3918) );
  XOR U4112 ( .A(n3919), .B(n3918), .Z(n3921) );
  XOR U4113 ( .A(n3920), .B(n3921), .Z(n3936) );
  XNOR U4114 ( .A(n3936), .B(sreg[423]), .Z(n3938) );
  NANDN U4115 ( .A(n3913), .B(sreg[422]), .Z(n3917) );
  NAND U4116 ( .A(n3915), .B(n3914), .Z(n3916) );
  NAND U4117 ( .A(n3917), .B(n3916), .Z(n3937) );
  XOR U4118 ( .A(n3938), .B(n3937), .Z(c[423]) );
  NANDN U4119 ( .A(n3919), .B(n3918), .Z(n3923) );
  OR U4120 ( .A(n3921), .B(n3920), .Z(n3922) );
  AND U4121 ( .A(n3923), .B(n3922), .Z(n3943) );
  NAND U4122 ( .A(n31), .B(n3924), .Z(n3926) );
  XOR U4123 ( .A(b[3]), .B(a[170]), .Z(n3947) );
  NAND U4124 ( .A(n5811), .B(n3947), .Z(n3925) );
  AND U4125 ( .A(n3926), .B(n3925), .Z(n3955) );
  NAND U4126 ( .A(b[0]), .B(a[172]), .Z(n3927) );
  XNOR U4127 ( .A(b[1]), .B(n3927), .Z(n3929) );
  NANDN U4128 ( .A(b[0]), .B(a[171]), .Z(n3928) );
  NAND U4129 ( .A(n3929), .B(n3928), .Z(n3954) );
  AND U4130 ( .A(b[3]), .B(a[168]), .Z(n3953) );
  XOR U4131 ( .A(n3954), .B(n3953), .Z(n3956) );
  XOR U4132 ( .A(n3955), .B(n3956), .Z(n3942) );
  NANDN U4133 ( .A(n3931), .B(n3930), .Z(n3935) );
  OR U4134 ( .A(n3933), .B(n3932), .Z(n3934) );
  AND U4135 ( .A(n3935), .B(n3934), .Z(n3941) );
  XOR U4136 ( .A(n3942), .B(n3941), .Z(n3944) );
  XOR U4137 ( .A(n3943), .B(n3944), .Z(n3959) );
  XNOR U4138 ( .A(n3959), .B(sreg[424]), .Z(n3961) );
  NANDN U4139 ( .A(n3936), .B(sreg[423]), .Z(n3940) );
  NAND U4140 ( .A(n3938), .B(n3937), .Z(n3939) );
  NAND U4141 ( .A(n3940), .B(n3939), .Z(n3960) );
  XOR U4142 ( .A(n3961), .B(n3960), .Z(c[424]) );
  NANDN U4143 ( .A(n3942), .B(n3941), .Z(n3946) );
  OR U4144 ( .A(n3944), .B(n3943), .Z(n3945) );
  AND U4145 ( .A(n3946), .B(n3945), .Z(n3966) );
  NAND U4146 ( .A(n31), .B(n3947), .Z(n3949) );
  XOR U4147 ( .A(b[3]), .B(a[171]), .Z(n3970) );
  NAND U4148 ( .A(n5811), .B(n3970), .Z(n3948) );
  AND U4149 ( .A(n3949), .B(n3948), .Z(n3978) );
  NAND U4150 ( .A(b[0]), .B(a[173]), .Z(n3950) );
  XNOR U4151 ( .A(b[1]), .B(n3950), .Z(n3952) );
  NANDN U4152 ( .A(b[0]), .B(a[172]), .Z(n3951) );
  NAND U4153 ( .A(n3952), .B(n3951), .Z(n3977) );
  AND U4154 ( .A(b[3]), .B(a[169]), .Z(n3976) );
  XOR U4155 ( .A(n3977), .B(n3976), .Z(n3979) );
  XOR U4156 ( .A(n3978), .B(n3979), .Z(n3965) );
  NANDN U4157 ( .A(n3954), .B(n3953), .Z(n3958) );
  OR U4158 ( .A(n3956), .B(n3955), .Z(n3957) );
  AND U4159 ( .A(n3958), .B(n3957), .Z(n3964) );
  XOR U4160 ( .A(n3965), .B(n3964), .Z(n3967) );
  XOR U4161 ( .A(n3966), .B(n3967), .Z(n3982) );
  XNOR U4162 ( .A(n3982), .B(sreg[425]), .Z(n3984) );
  NANDN U4163 ( .A(n3959), .B(sreg[424]), .Z(n3963) );
  NAND U4164 ( .A(n3961), .B(n3960), .Z(n3962) );
  NAND U4165 ( .A(n3963), .B(n3962), .Z(n3983) );
  XOR U4166 ( .A(n3984), .B(n3983), .Z(c[425]) );
  NANDN U4167 ( .A(n3965), .B(n3964), .Z(n3969) );
  OR U4168 ( .A(n3967), .B(n3966), .Z(n3968) );
  AND U4169 ( .A(n3969), .B(n3968), .Z(n3989) );
  NAND U4170 ( .A(n31), .B(n3970), .Z(n3972) );
  XOR U4171 ( .A(b[3]), .B(a[172]), .Z(n3993) );
  NAND U4172 ( .A(n5811), .B(n3993), .Z(n3971) );
  AND U4173 ( .A(n3972), .B(n3971), .Z(n4001) );
  AND U4174 ( .A(b[3]), .B(a[170]), .Z(n3999) );
  NAND U4175 ( .A(b[0]), .B(a[174]), .Z(n3973) );
  XNOR U4176 ( .A(b[1]), .B(n3973), .Z(n3975) );
  NANDN U4177 ( .A(b[0]), .B(a[173]), .Z(n3974) );
  NAND U4178 ( .A(n3975), .B(n3974), .Z(n4000) );
  XOR U4179 ( .A(n3999), .B(n4000), .Z(n4002) );
  XOR U4180 ( .A(n4001), .B(n4002), .Z(n3988) );
  NANDN U4181 ( .A(n3977), .B(n3976), .Z(n3981) );
  OR U4182 ( .A(n3979), .B(n3978), .Z(n3980) );
  AND U4183 ( .A(n3981), .B(n3980), .Z(n3987) );
  XOR U4184 ( .A(n3988), .B(n3987), .Z(n3990) );
  XOR U4185 ( .A(n3989), .B(n3990), .Z(n4005) );
  XNOR U4186 ( .A(n4005), .B(sreg[426]), .Z(n4007) );
  NANDN U4187 ( .A(n3982), .B(sreg[425]), .Z(n3986) );
  NAND U4188 ( .A(n3984), .B(n3983), .Z(n3985) );
  NAND U4189 ( .A(n3986), .B(n3985), .Z(n4006) );
  XOR U4190 ( .A(n4007), .B(n4006), .Z(c[426]) );
  NANDN U4191 ( .A(n3988), .B(n3987), .Z(n3992) );
  OR U4192 ( .A(n3990), .B(n3989), .Z(n3991) );
  AND U4193 ( .A(n3992), .B(n3991), .Z(n4012) );
  NAND U4194 ( .A(n31), .B(n3993), .Z(n3995) );
  XOR U4195 ( .A(b[3]), .B(a[173]), .Z(n4016) );
  NAND U4196 ( .A(n5811), .B(n4016), .Z(n3994) );
  AND U4197 ( .A(n3995), .B(n3994), .Z(n4024) );
  NAND U4198 ( .A(b[0]), .B(a[175]), .Z(n3996) );
  XNOR U4199 ( .A(b[1]), .B(n3996), .Z(n3998) );
  NANDN U4200 ( .A(b[0]), .B(a[174]), .Z(n3997) );
  NAND U4201 ( .A(n3998), .B(n3997), .Z(n4023) );
  AND U4202 ( .A(b[3]), .B(a[171]), .Z(n4022) );
  XOR U4203 ( .A(n4023), .B(n4022), .Z(n4025) );
  XOR U4204 ( .A(n4024), .B(n4025), .Z(n4011) );
  NANDN U4205 ( .A(n4000), .B(n3999), .Z(n4004) );
  OR U4206 ( .A(n4002), .B(n4001), .Z(n4003) );
  AND U4207 ( .A(n4004), .B(n4003), .Z(n4010) );
  XOR U4208 ( .A(n4011), .B(n4010), .Z(n4013) );
  XOR U4209 ( .A(n4012), .B(n4013), .Z(n4028) );
  XNOR U4210 ( .A(n4028), .B(sreg[427]), .Z(n4030) );
  NANDN U4211 ( .A(n4005), .B(sreg[426]), .Z(n4009) );
  NAND U4212 ( .A(n4007), .B(n4006), .Z(n4008) );
  NAND U4213 ( .A(n4009), .B(n4008), .Z(n4029) );
  XOR U4214 ( .A(n4030), .B(n4029), .Z(c[427]) );
  NANDN U4215 ( .A(n4011), .B(n4010), .Z(n4015) );
  OR U4216 ( .A(n4013), .B(n4012), .Z(n4014) );
  AND U4217 ( .A(n4015), .B(n4014), .Z(n4035) );
  NAND U4218 ( .A(n31), .B(n4016), .Z(n4018) );
  XOR U4219 ( .A(b[3]), .B(a[174]), .Z(n4039) );
  NAND U4220 ( .A(n5811), .B(n4039), .Z(n4017) );
  AND U4221 ( .A(n4018), .B(n4017), .Z(n4047) );
  NAND U4222 ( .A(b[0]), .B(a[176]), .Z(n4019) );
  XNOR U4223 ( .A(b[1]), .B(n4019), .Z(n4021) );
  NANDN U4224 ( .A(b[0]), .B(a[175]), .Z(n4020) );
  NAND U4225 ( .A(n4021), .B(n4020), .Z(n4046) );
  AND U4226 ( .A(b[3]), .B(a[172]), .Z(n4045) );
  XOR U4227 ( .A(n4046), .B(n4045), .Z(n4048) );
  XOR U4228 ( .A(n4047), .B(n4048), .Z(n4034) );
  NANDN U4229 ( .A(n4023), .B(n4022), .Z(n4027) );
  OR U4230 ( .A(n4025), .B(n4024), .Z(n4026) );
  AND U4231 ( .A(n4027), .B(n4026), .Z(n4033) );
  XOR U4232 ( .A(n4034), .B(n4033), .Z(n4036) );
  XOR U4233 ( .A(n4035), .B(n4036), .Z(n4051) );
  XNOR U4234 ( .A(n4051), .B(sreg[428]), .Z(n4053) );
  NANDN U4235 ( .A(n4028), .B(sreg[427]), .Z(n4032) );
  NAND U4236 ( .A(n4030), .B(n4029), .Z(n4031) );
  NAND U4237 ( .A(n4032), .B(n4031), .Z(n4052) );
  XOR U4238 ( .A(n4053), .B(n4052), .Z(c[428]) );
  NANDN U4239 ( .A(n4034), .B(n4033), .Z(n4038) );
  OR U4240 ( .A(n4036), .B(n4035), .Z(n4037) );
  AND U4241 ( .A(n4038), .B(n4037), .Z(n4058) );
  NAND U4242 ( .A(n31), .B(n4039), .Z(n4041) );
  XOR U4243 ( .A(b[3]), .B(a[175]), .Z(n4062) );
  NAND U4244 ( .A(n5811), .B(n4062), .Z(n4040) );
  AND U4245 ( .A(n4041), .B(n4040), .Z(n4070) );
  NAND U4246 ( .A(b[0]), .B(a[177]), .Z(n4042) );
  XNOR U4247 ( .A(b[1]), .B(n4042), .Z(n4044) );
  NANDN U4248 ( .A(b[0]), .B(a[176]), .Z(n4043) );
  NAND U4249 ( .A(n4044), .B(n4043), .Z(n4069) );
  AND U4250 ( .A(b[3]), .B(a[173]), .Z(n4068) );
  XOR U4251 ( .A(n4069), .B(n4068), .Z(n4071) );
  XOR U4252 ( .A(n4070), .B(n4071), .Z(n4057) );
  NANDN U4253 ( .A(n4046), .B(n4045), .Z(n4050) );
  OR U4254 ( .A(n4048), .B(n4047), .Z(n4049) );
  AND U4255 ( .A(n4050), .B(n4049), .Z(n4056) );
  XOR U4256 ( .A(n4057), .B(n4056), .Z(n4059) );
  XOR U4257 ( .A(n4058), .B(n4059), .Z(n4074) );
  XNOR U4258 ( .A(n4074), .B(sreg[429]), .Z(n4076) );
  NANDN U4259 ( .A(n4051), .B(sreg[428]), .Z(n4055) );
  NAND U4260 ( .A(n4053), .B(n4052), .Z(n4054) );
  NAND U4261 ( .A(n4055), .B(n4054), .Z(n4075) );
  XOR U4262 ( .A(n4076), .B(n4075), .Z(c[429]) );
  NANDN U4263 ( .A(n4057), .B(n4056), .Z(n4061) );
  OR U4264 ( .A(n4059), .B(n4058), .Z(n4060) );
  AND U4265 ( .A(n4061), .B(n4060), .Z(n4081) );
  NAND U4266 ( .A(n31), .B(n4062), .Z(n4064) );
  XOR U4267 ( .A(b[3]), .B(a[176]), .Z(n4085) );
  NAND U4268 ( .A(n5811), .B(n4085), .Z(n4063) );
  AND U4269 ( .A(n4064), .B(n4063), .Z(n4093) );
  NAND U4270 ( .A(b[0]), .B(a[178]), .Z(n4065) );
  XNOR U4271 ( .A(b[1]), .B(n4065), .Z(n4067) );
  NANDN U4272 ( .A(b[0]), .B(a[177]), .Z(n4066) );
  NAND U4273 ( .A(n4067), .B(n4066), .Z(n4092) );
  AND U4274 ( .A(b[3]), .B(a[174]), .Z(n4091) );
  XOR U4275 ( .A(n4092), .B(n4091), .Z(n4094) );
  XOR U4276 ( .A(n4093), .B(n4094), .Z(n4080) );
  NANDN U4277 ( .A(n4069), .B(n4068), .Z(n4073) );
  OR U4278 ( .A(n4071), .B(n4070), .Z(n4072) );
  AND U4279 ( .A(n4073), .B(n4072), .Z(n4079) );
  XOR U4280 ( .A(n4080), .B(n4079), .Z(n4082) );
  XOR U4281 ( .A(n4081), .B(n4082), .Z(n4097) );
  XNOR U4282 ( .A(n4097), .B(sreg[430]), .Z(n4099) );
  NANDN U4283 ( .A(n4074), .B(sreg[429]), .Z(n4078) );
  NAND U4284 ( .A(n4076), .B(n4075), .Z(n4077) );
  NAND U4285 ( .A(n4078), .B(n4077), .Z(n4098) );
  XOR U4286 ( .A(n4099), .B(n4098), .Z(c[430]) );
  NANDN U4287 ( .A(n4080), .B(n4079), .Z(n4084) );
  OR U4288 ( .A(n4082), .B(n4081), .Z(n4083) );
  AND U4289 ( .A(n4084), .B(n4083), .Z(n4104) );
  NAND U4290 ( .A(n31), .B(n4085), .Z(n4087) );
  XOR U4291 ( .A(b[3]), .B(a[177]), .Z(n4108) );
  NAND U4292 ( .A(n5811), .B(n4108), .Z(n4086) );
  AND U4293 ( .A(n4087), .B(n4086), .Z(n4116) );
  NAND U4294 ( .A(b[0]), .B(a[179]), .Z(n4088) );
  XNOR U4295 ( .A(b[1]), .B(n4088), .Z(n4090) );
  NANDN U4296 ( .A(b[0]), .B(a[178]), .Z(n4089) );
  NAND U4297 ( .A(n4090), .B(n4089), .Z(n4115) );
  AND U4298 ( .A(b[3]), .B(a[175]), .Z(n4114) );
  XOR U4299 ( .A(n4115), .B(n4114), .Z(n4117) );
  XOR U4300 ( .A(n4116), .B(n4117), .Z(n4103) );
  NANDN U4301 ( .A(n4092), .B(n4091), .Z(n4096) );
  OR U4302 ( .A(n4094), .B(n4093), .Z(n4095) );
  AND U4303 ( .A(n4096), .B(n4095), .Z(n4102) );
  XOR U4304 ( .A(n4103), .B(n4102), .Z(n4105) );
  XOR U4305 ( .A(n4104), .B(n4105), .Z(n4120) );
  XNOR U4306 ( .A(n4120), .B(sreg[431]), .Z(n4122) );
  NANDN U4307 ( .A(n4097), .B(sreg[430]), .Z(n4101) );
  NAND U4308 ( .A(n4099), .B(n4098), .Z(n4100) );
  NAND U4309 ( .A(n4101), .B(n4100), .Z(n4121) );
  XOR U4310 ( .A(n4122), .B(n4121), .Z(c[431]) );
  NANDN U4311 ( .A(n4103), .B(n4102), .Z(n4107) );
  OR U4312 ( .A(n4105), .B(n4104), .Z(n4106) );
  AND U4313 ( .A(n4107), .B(n4106), .Z(n4127) );
  NAND U4314 ( .A(n31), .B(n4108), .Z(n4110) );
  XOR U4315 ( .A(b[3]), .B(a[178]), .Z(n4131) );
  NAND U4316 ( .A(n5811), .B(n4131), .Z(n4109) );
  AND U4317 ( .A(n4110), .B(n4109), .Z(n4139) );
  AND U4318 ( .A(b[3]), .B(a[176]), .Z(n4137) );
  NAND U4319 ( .A(b[0]), .B(a[180]), .Z(n4111) );
  XNOR U4320 ( .A(b[1]), .B(n4111), .Z(n4113) );
  NANDN U4321 ( .A(b[0]), .B(a[179]), .Z(n4112) );
  NAND U4322 ( .A(n4113), .B(n4112), .Z(n4138) );
  XOR U4323 ( .A(n4137), .B(n4138), .Z(n4140) );
  XOR U4324 ( .A(n4139), .B(n4140), .Z(n4126) );
  NANDN U4325 ( .A(n4115), .B(n4114), .Z(n4119) );
  OR U4326 ( .A(n4117), .B(n4116), .Z(n4118) );
  AND U4327 ( .A(n4119), .B(n4118), .Z(n4125) );
  XOR U4328 ( .A(n4126), .B(n4125), .Z(n4128) );
  XOR U4329 ( .A(n4127), .B(n4128), .Z(n4143) );
  XNOR U4330 ( .A(n4143), .B(sreg[432]), .Z(n4145) );
  NANDN U4331 ( .A(n4120), .B(sreg[431]), .Z(n4124) );
  NAND U4332 ( .A(n4122), .B(n4121), .Z(n4123) );
  NAND U4333 ( .A(n4124), .B(n4123), .Z(n4144) );
  XOR U4334 ( .A(n4145), .B(n4144), .Z(c[432]) );
  NANDN U4335 ( .A(n4126), .B(n4125), .Z(n4130) );
  OR U4336 ( .A(n4128), .B(n4127), .Z(n4129) );
  AND U4337 ( .A(n4130), .B(n4129), .Z(n4150) );
  NAND U4338 ( .A(n31), .B(n4131), .Z(n4133) );
  XOR U4339 ( .A(b[3]), .B(a[179]), .Z(n4154) );
  NAND U4340 ( .A(n5811), .B(n4154), .Z(n4132) );
  AND U4341 ( .A(n4133), .B(n4132), .Z(n4162) );
  NAND U4342 ( .A(b[0]), .B(a[181]), .Z(n4134) );
  XNOR U4343 ( .A(b[1]), .B(n4134), .Z(n4136) );
  NANDN U4344 ( .A(b[0]), .B(a[180]), .Z(n4135) );
  NAND U4345 ( .A(n4136), .B(n4135), .Z(n4161) );
  AND U4346 ( .A(b[3]), .B(a[177]), .Z(n4160) );
  XOR U4347 ( .A(n4161), .B(n4160), .Z(n4163) );
  XOR U4348 ( .A(n4162), .B(n4163), .Z(n4149) );
  NANDN U4349 ( .A(n4138), .B(n4137), .Z(n4142) );
  OR U4350 ( .A(n4140), .B(n4139), .Z(n4141) );
  AND U4351 ( .A(n4142), .B(n4141), .Z(n4148) );
  XOR U4352 ( .A(n4149), .B(n4148), .Z(n4151) );
  XOR U4353 ( .A(n4150), .B(n4151), .Z(n4166) );
  XNOR U4354 ( .A(n4166), .B(sreg[433]), .Z(n4168) );
  NANDN U4355 ( .A(n4143), .B(sreg[432]), .Z(n4147) );
  NAND U4356 ( .A(n4145), .B(n4144), .Z(n4146) );
  NAND U4357 ( .A(n4147), .B(n4146), .Z(n4167) );
  XOR U4358 ( .A(n4168), .B(n4167), .Z(c[433]) );
  NANDN U4359 ( .A(n4149), .B(n4148), .Z(n4153) );
  OR U4360 ( .A(n4151), .B(n4150), .Z(n4152) );
  AND U4361 ( .A(n4153), .B(n4152), .Z(n4173) );
  NAND U4362 ( .A(n31), .B(n4154), .Z(n4156) );
  XOR U4363 ( .A(b[3]), .B(a[180]), .Z(n4177) );
  NAND U4364 ( .A(n5811), .B(n4177), .Z(n4155) );
  AND U4365 ( .A(n4156), .B(n4155), .Z(n4185) );
  AND U4366 ( .A(b[3]), .B(a[178]), .Z(n4183) );
  NAND U4367 ( .A(b[0]), .B(a[182]), .Z(n4157) );
  XNOR U4368 ( .A(b[1]), .B(n4157), .Z(n4159) );
  NANDN U4369 ( .A(b[0]), .B(a[181]), .Z(n4158) );
  NAND U4370 ( .A(n4159), .B(n4158), .Z(n4184) );
  XOR U4371 ( .A(n4183), .B(n4184), .Z(n4186) );
  XOR U4372 ( .A(n4185), .B(n4186), .Z(n4172) );
  NANDN U4373 ( .A(n4161), .B(n4160), .Z(n4165) );
  OR U4374 ( .A(n4163), .B(n4162), .Z(n4164) );
  AND U4375 ( .A(n4165), .B(n4164), .Z(n4171) );
  XOR U4376 ( .A(n4172), .B(n4171), .Z(n4174) );
  XOR U4377 ( .A(n4173), .B(n4174), .Z(n4189) );
  XNOR U4378 ( .A(n4189), .B(sreg[434]), .Z(n4191) );
  NANDN U4379 ( .A(n4166), .B(sreg[433]), .Z(n4170) );
  NAND U4380 ( .A(n4168), .B(n4167), .Z(n4169) );
  NAND U4381 ( .A(n4170), .B(n4169), .Z(n4190) );
  XOR U4382 ( .A(n4191), .B(n4190), .Z(c[434]) );
  NANDN U4383 ( .A(n4172), .B(n4171), .Z(n4176) );
  OR U4384 ( .A(n4174), .B(n4173), .Z(n4175) );
  AND U4385 ( .A(n4176), .B(n4175), .Z(n4196) );
  NAND U4386 ( .A(n31), .B(n4177), .Z(n4179) );
  XOR U4387 ( .A(b[3]), .B(a[181]), .Z(n4200) );
  NAND U4388 ( .A(n5811), .B(n4200), .Z(n4178) );
  AND U4389 ( .A(n4179), .B(n4178), .Z(n4208) );
  AND U4390 ( .A(b[0]), .B(a[183]), .Z(n4180) );
  XOR U4391 ( .A(b[1]), .B(n4180), .Z(n4182) );
  NANDN U4392 ( .A(b[0]), .B(a[182]), .Z(n4181) );
  AND U4393 ( .A(n4182), .B(n4181), .Z(n4206) );
  NAND U4394 ( .A(b[3]), .B(a[179]), .Z(n4207) );
  XOR U4395 ( .A(n4206), .B(n4207), .Z(n4209) );
  XOR U4396 ( .A(n4208), .B(n4209), .Z(n4195) );
  NANDN U4397 ( .A(n4184), .B(n4183), .Z(n4188) );
  OR U4398 ( .A(n4186), .B(n4185), .Z(n4187) );
  AND U4399 ( .A(n4188), .B(n4187), .Z(n4194) );
  XOR U4400 ( .A(n4195), .B(n4194), .Z(n4197) );
  XOR U4401 ( .A(n4196), .B(n4197), .Z(n4212) );
  XNOR U4402 ( .A(n4212), .B(sreg[435]), .Z(n4214) );
  NANDN U4403 ( .A(n4189), .B(sreg[434]), .Z(n4193) );
  NAND U4404 ( .A(n4191), .B(n4190), .Z(n4192) );
  NAND U4405 ( .A(n4193), .B(n4192), .Z(n4213) );
  XOR U4406 ( .A(n4214), .B(n4213), .Z(c[435]) );
  NANDN U4407 ( .A(n4195), .B(n4194), .Z(n4199) );
  OR U4408 ( .A(n4197), .B(n4196), .Z(n4198) );
  AND U4409 ( .A(n4199), .B(n4198), .Z(n4219) );
  NAND U4410 ( .A(n31), .B(n4200), .Z(n4202) );
  XOR U4411 ( .A(b[3]), .B(a[182]), .Z(n4223) );
  NAND U4412 ( .A(n5811), .B(n4223), .Z(n4201) );
  AND U4413 ( .A(n4202), .B(n4201), .Z(n4231) );
  NAND U4414 ( .A(b[0]), .B(a[184]), .Z(n4203) );
  XNOR U4415 ( .A(b[1]), .B(n4203), .Z(n4205) );
  NANDN U4416 ( .A(b[0]), .B(a[183]), .Z(n4204) );
  NAND U4417 ( .A(n4205), .B(n4204), .Z(n4230) );
  AND U4418 ( .A(b[3]), .B(a[180]), .Z(n4229) );
  XOR U4419 ( .A(n4230), .B(n4229), .Z(n4232) );
  XOR U4420 ( .A(n4231), .B(n4232), .Z(n4218) );
  NANDN U4421 ( .A(n4207), .B(n4206), .Z(n4211) );
  OR U4422 ( .A(n4209), .B(n4208), .Z(n4210) );
  AND U4423 ( .A(n4211), .B(n4210), .Z(n4217) );
  XOR U4424 ( .A(n4218), .B(n4217), .Z(n4220) );
  XOR U4425 ( .A(n4219), .B(n4220), .Z(n4235) );
  XNOR U4426 ( .A(n4235), .B(sreg[436]), .Z(n4237) );
  NANDN U4427 ( .A(n4212), .B(sreg[435]), .Z(n4216) );
  NAND U4428 ( .A(n4214), .B(n4213), .Z(n4215) );
  NAND U4429 ( .A(n4216), .B(n4215), .Z(n4236) );
  XOR U4430 ( .A(n4237), .B(n4236), .Z(c[436]) );
  NANDN U4431 ( .A(n4218), .B(n4217), .Z(n4222) );
  OR U4432 ( .A(n4220), .B(n4219), .Z(n4221) );
  AND U4433 ( .A(n4222), .B(n4221), .Z(n4242) );
  NAND U4434 ( .A(n31), .B(n4223), .Z(n4225) );
  XOR U4435 ( .A(b[3]), .B(a[183]), .Z(n4246) );
  NAND U4436 ( .A(n5811), .B(n4246), .Z(n4224) );
  AND U4437 ( .A(n4225), .B(n4224), .Z(n4254) );
  NAND U4438 ( .A(b[0]), .B(a[185]), .Z(n4226) );
  XNOR U4439 ( .A(b[1]), .B(n4226), .Z(n4228) );
  NANDN U4440 ( .A(b[0]), .B(a[184]), .Z(n4227) );
  NAND U4441 ( .A(n4228), .B(n4227), .Z(n4253) );
  AND U4442 ( .A(b[3]), .B(a[181]), .Z(n4252) );
  XOR U4443 ( .A(n4253), .B(n4252), .Z(n4255) );
  XOR U4444 ( .A(n4254), .B(n4255), .Z(n4241) );
  NANDN U4445 ( .A(n4230), .B(n4229), .Z(n4234) );
  OR U4446 ( .A(n4232), .B(n4231), .Z(n4233) );
  AND U4447 ( .A(n4234), .B(n4233), .Z(n4240) );
  XOR U4448 ( .A(n4241), .B(n4240), .Z(n4243) );
  XOR U4449 ( .A(n4242), .B(n4243), .Z(n4258) );
  XNOR U4450 ( .A(n4258), .B(sreg[437]), .Z(n4260) );
  NANDN U4451 ( .A(n4235), .B(sreg[436]), .Z(n4239) );
  NAND U4452 ( .A(n4237), .B(n4236), .Z(n4238) );
  NAND U4453 ( .A(n4239), .B(n4238), .Z(n4259) );
  XOR U4454 ( .A(n4260), .B(n4259), .Z(c[437]) );
  NANDN U4455 ( .A(n4241), .B(n4240), .Z(n4245) );
  OR U4456 ( .A(n4243), .B(n4242), .Z(n4244) );
  AND U4457 ( .A(n4245), .B(n4244), .Z(n4265) );
  NAND U4458 ( .A(n31), .B(n4246), .Z(n4248) );
  XOR U4459 ( .A(b[3]), .B(a[184]), .Z(n4269) );
  NAND U4460 ( .A(n5811), .B(n4269), .Z(n4247) );
  AND U4461 ( .A(n4248), .B(n4247), .Z(n4277) );
  NAND U4462 ( .A(b[0]), .B(a[186]), .Z(n4249) );
  XNOR U4463 ( .A(b[1]), .B(n4249), .Z(n4251) );
  NANDN U4464 ( .A(b[0]), .B(a[185]), .Z(n4250) );
  NAND U4465 ( .A(n4251), .B(n4250), .Z(n4276) );
  AND U4466 ( .A(b[3]), .B(a[182]), .Z(n4275) );
  XOR U4467 ( .A(n4276), .B(n4275), .Z(n4278) );
  XOR U4468 ( .A(n4277), .B(n4278), .Z(n4264) );
  NANDN U4469 ( .A(n4253), .B(n4252), .Z(n4257) );
  OR U4470 ( .A(n4255), .B(n4254), .Z(n4256) );
  AND U4471 ( .A(n4257), .B(n4256), .Z(n4263) );
  XOR U4472 ( .A(n4264), .B(n4263), .Z(n4266) );
  XOR U4473 ( .A(n4265), .B(n4266), .Z(n4281) );
  XNOR U4474 ( .A(n4281), .B(sreg[438]), .Z(n4283) );
  NANDN U4475 ( .A(n4258), .B(sreg[437]), .Z(n4262) );
  NAND U4476 ( .A(n4260), .B(n4259), .Z(n4261) );
  NAND U4477 ( .A(n4262), .B(n4261), .Z(n4282) );
  XOR U4478 ( .A(n4283), .B(n4282), .Z(c[438]) );
  NANDN U4479 ( .A(n4264), .B(n4263), .Z(n4268) );
  OR U4480 ( .A(n4266), .B(n4265), .Z(n4267) );
  AND U4481 ( .A(n4268), .B(n4267), .Z(n4288) );
  NAND U4482 ( .A(n31), .B(n4269), .Z(n4271) );
  XOR U4483 ( .A(b[3]), .B(a[185]), .Z(n4292) );
  NAND U4484 ( .A(n5811), .B(n4292), .Z(n4270) );
  AND U4485 ( .A(n4271), .B(n4270), .Z(n4300) );
  NAND U4486 ( .A(b[0]), .B(a[187]), .Z(n4272) );
  XNOR U4487 ( .A(b[1]), .B(n4272), .Z(n4274) );
  NANDN U4488 ( .A(b[0]), .B(a[186]), .Z(n4273) );
  NAND U4489 ( .A(n4274), .B(n4273), .Z(n4299) );
  AND U4490 ( .A(b[3]), .B(a[183]), .Z(n4298) );
  XOR U4491 ( .A(n4299), .B(n4298), .Z(n4301) );
  XOR U4492 ( .A(n4300), .B(n4301), .Z(n4287) );
  NANDN U4493 ( .A(n4276), .B(n4275), .Z(n4280) );
  OR U4494 ( .A(n4278), .B(n4277), .Z(n4279) );
  AND U4495 ( .A(n4280), .B(n4279), .Z(n4286) );
  XOR U4496 ( .A(n4287), .B(n4286), .Z(n4289) );
  XOR U4497 ( .A(n4288), .B(n4289), .Z(n4304) );
  XNOR U4498 ( .A(n4304), .B(sreg[439]), .Z(n4306) );
  NANDN U4499 ( .A(n4281), .B(sreg[438]), .Z(n4285) );
  NAND U4500 ( .A(n4283), .B(n4282), .Z(n4284) );
  NAND U4501 ( .A(n4285), .B(n4284), .Z(n4305) );
  XOR U4502 ( .A(n4306), .B(n4305), .Z(c[439]) );
  NANDN U4503 ( .A(n4287), .B(n4286), .Z(n4291) );
  OR U4504 ( .A(n4289), .B(n4288), .Z(n4290) );
  AND U4505 ( .A(n4291), .B(n4290), .Z(n4311) );
  NAND U4506 ( .A(n31), .B(n4292), .Z(n4294) );
  XOR U4507 ( .A(b[3]), .B(a[186]), .Z(n4315) );
  NAND U4508 ( .A(n5811), .B(n4315), .Z(n4293) );
  AND U4509 ( .A(n4294), .B(n4293), .Z(n4323) );
  NAND U4510 ( .A(b[0]), .B(a[188]), .Z(n4295) );
  XNOR U4511 ( .A(b[1]), .B(n4295), .Z(n4297) );
  NANDN U4512 ( .A(b[0]), .B(a[187]), .Z(n4296) );
  NAND U4513 ( .A(n4297), .B(n4296), .Z(n4322) );
  AND U4514 ( .A(b[3]), .B(a[184]), .Z(n4321) );
  XOR U4515 ( .A(n4322), .B(n4321), .Z(n4324) );
  XOR U4516 ( .A(n4323), .B(n4324), .Z(n4310) );
  NANDN U4517 ( .A(n4299), .B(n4298), .Z(n4303) );
  OR U4518 ( .A(n4301), .B(n4300), .Z(n4302) );
  AND U4519 ( .A(n4303), .B(n4302), .Z(n4309) );
  XOR U4520 ( .A(n4310), .B(n4309), .Z(n4312) );
  XOR U4521 ( .A(n4311), .B(n4312), .Z(n4327) );
  XNOR U4522 ( .A(n4327), .B(sreg[440]), .Z(n4329) );
  NANDN U4523 ( .A(n4304), .B(sreg[439]), .Z(n4308) );
  NAND U4524 ( .A(n4306), .B(n4305), .Z(n4307) );
  NAND U4525 ( .A(n4308), .B(n4307), .Z(n4328) );
  XOR U4526 ( .A(n4329), .B(n4328), .Z(c[440]) );
  NANDN U4527 ( .A(n4310), .B(n4309), .Z(n4314) );
  OR U4528 ( .A(n4312), .B(n4311), .Z(n4313) );
  AND U4529 ( .A(n4314), .B(n4313), .Z(n4334) );
  NAND U4530 ( .A(n31), .B(n4315), .Z(n4317) );
  XOR U4531 ( .A(b[3]), .B(a[187]), .Z(n4338) );
  NAND U4532 ( .A(n5811), .B(n4338), .Z(n4316) );
  AND U4533 ( .A(n4317), .B(n4316), .Z(n4346) );
  NAND U4534 ( .A(b[0]), .B(a[189]), .Z(n4318) );
  XNOR U4535 ( .A(b[1]), .B(n4318), .Z(n4320) );
  NANDN U4536 ( .A(b[0]), .B(a[188]), .Z(n4319) );
  NAND U4537 ( .A(n4320), .B(n4319), .Z(n4345) );
  AND U4538 ( .A(b[3]), .B(a[185]), .Z(n4344) );
  XOR U4539 ( .A(n4345), .B(n4344), .Z(n4347) );
  XOR U4540 ( .A(n4346), .B(n4347), .Z(n4333) );
  NANDN U4541 ( .A(n4322), .B(n4321), .Z(n4326) );
  OR U4542 ( .A(n4324), .B(n4323), .Z(n4325) );
  AND U4543 ( .A(n4326), .B(n4325), .Z(n4332) );
  XOR U4544 ( .A(n4333), .B(n4332), .Z(n4335) );
  XOR U4545 ( .A(n4334), .B(n4335), .Z(n4350) );
  XNOR U4546 ( .A(n4350), .B(sreg[441]), .Z(n4352) );
  NANDN U4547 ( .A(n4327), .B(sreg[440]), .Z(n4331) );
  NAND U4548 ( .A(n4329), .B(n4328), .Z(n4330) );
  NAND U4549 ( .A(n4331), .B(n4330), .Z(n4351) );
  XOR U4550 ( .A(n4352), .B(n4351), .Z(c[441]) );
  NANDN U4551 ( .A(n4333), .B(n4332), .Z(n4337) );
  OR U4552 ( .A(n4335), .B(n4334), .Z(n4336) );
  AND U4553 ( .A(n4337), .B(n4336), .Z(n4357) );
  NAND U4554 ( .A(n31), .B(n4338), .Z(n4340) );
  XOR U4555 ( .A(b[3]), .B(a[188]), .Z(n4361) );
  NAND U4556 ( .A(n5811), .B(n4361), .Z(n4339) );
  AND U4557 ( .A(n4340), .B(n4339), .Z(n4369) );
  NAND U4558 ( .A(b[0]), .B(a[190]), .Z(n4341) );
  XNOR U4559 ( .A(b[1]), .B(n4341), .Z(n4343) );
  NANDN U4560 ( .A(b[0]), .B(a[189]), .Z(n4342) );
  NAND U4561 ( .A(n4343), .B(n4342), .Z(n4368) );
  AND U4562 ( .A(b[3]), .B(a[186]), .Z(n4367) );
  XOR U4563 ( .A(n4368), .B(n4367), .Z(n4370) );
  XOR U4564 ( .A(n4369), .B(n4370), .Z(n4356) );
  NANDN U4565 ( .A(n4345), .B(n4344), .Z(n4349) );
  OR U4566 ( .A(n4347), .B(n4346), .Z(n4348) );
  AND U4567 ( .A(n4349), .B(n4348), .Z(n4355) );
  XOR U4568 ( .A(n4356), .B(n4355), .Z(n4358) );
  XOR U4569 ( .A(n4357), .B(n4358), .Z(n4373) );
  XNOR U4570 ( .A(n4373), .B(sreg[442]), .Z(n4375) );
  NANDN U4571 ( .A(n4350), .B(sreg[441]), .Z(n4354) );
  NAND U4572 ( .A(n4352), .B(n4351), .Z(n4353) );
  NAND U4573 ( .A(n4354), .B(n4353), .Z(n4374) );
  XOR U4574 ( .A(n4375), .B(n4374), .Z(c[442]) );
  NANDN U4575 ( .A(n4356), .B(n4355), .Z(n4360) );
  OR U4576 ( .A(n4358), .B(n4357), .Z(n4359) );
  AND U4577 ( .A(n4360), .B(n4359), .Z(n4380) );
  NAND U4578 ( .A(n31), .B(n4361), .Z(n4363) );
  XOR U4579 ( .A(b[3]), .B(a[189]), .Z(n4384) );
  NAND U4580 ( .A(n5811), .B(n4384), .Z(n4362) );
  AND U4581 ( .A(n4363), .B(n4362), .Z(n4392) );
  NAND U4582 ( .A(b[0]), .B(a[191]), .Z(n4364) );
  XNOR U4583 ( .A(b[1]), .B(n4364), .Z(n4366) );
  NANDN U4584 ( .A(b[0]), .B(a[190]), .Z(n4365) );
  NAND U4585 ( .A(n4366), .B(n4365), .Z(n4391) );
  AND U4586 ( .A(b[3]), .B(a[187]), .Z(n4390) );
  XOR U4587 ( .A(n4391), .B(n4390), .Z(n4393) );
  XOR U4588 ( .A(n4392), .B(n4393), .Z(n4379) );
  NANDN U4589 ( .A(n4368), .B(n4367), .Z(n4372) );
  OR U4590 ( .A(n4370), .B(n4369), .Z(n4371) );
  AND U4591 ( .A(n4372), .B(n4371), .Z(n4378) );
  XOR U4592 ( .A(n4379), .B(n4378), .Z(n4381) );
  XOR U4593 ( .A(n4380), .B(n4381), .Z(n4396) );
  XNOR U4594 ( .A(n4396), .B(sreg[443]), .Z(n4398) );
  NANDN U4595 ( .A(n4373), .B(sreg[442]), .Z(n4377) );
  NAND U4596 ( .A(n4375), .B(n4374), .Z(n4376) );
  NAND U4597 ( .A(n4377), .B(n4376), .Z(n4397) );
  XOR U4598 ( .A(n4398), .B(n4397), .Z(c[443]) );
  NANDN U4599 ( .A(n4379), .B(n4378), .Z(n4383) );
  OR U4600 ( .A(n4381), .B(n4380), .Z(n4382) );
  AND U4601 ( .A(n4383), .B(n4382), .Z(n4403) );
  NAND U4602 ( .A(n31), .B(n4384), .Z(n4386) );
  XOR U4603 ( .A(b[3]), .B(a[190]), .Z(n4407) );
  NAND U4604 ( .A(n5811), .B(n4407), .Z(n4385) );
  AND U4605 ( .A(n4386), .B(n4385), .Z(n4415) );
  NAND U4606 ( .A(b[0]), .B(a[192]), .Z(n4387) );
  XNOR U4607 ( .A(b[1]), .B(n4387), .Z(n4389) );
  NANDN U4608 ( .A(b[0]), .B(a[191]), .Z(n4388) );
  NAND U4609 ( .A(n4389), .B(n4388), .Z(n4414) );
  AND U4610 ( .A(b[3]), .B(a[188]), .Z(n4413) );
  XOR U4611 ( .A(n4414), .B(n4413), .Z(n4416) );
  XOR U4612 ( .A(n4415), .B(n4416), .Z(n4402) );
  NANDN U4613 ( .A(n4391), .B(n4390), .Z(n4395) );
  OR U4614 ( .A(n4393), .B(n4392), .Z(n4394) );
  AND U4615 ( .A(n4395), .B(n4394), .Z(n4401) );
  XOR U4616 ( .A(n4402), .B(n4401), .Z(n4404) );
  XOR U4617 ( .A(n4403), .B(n4404), .Z(n4419) );
  XNOR U4618 ( .A(n4419), .B(sreg[444]), .Z(n4421) );
  NANDN U4619 ( .A(n4396), .B(sreg[443]), .Z(n4400) );
  NAND U4620 ( .A(n4398), .B(n4397), .Z(n4399) );
  NAND U4621 ( .A(n4400), .B(n4399), .Z(n4420) );
  XOR U4622 ( .A(n4421), .B(n4420), .Z(c[444]) );
  NANDN U4623 ( .A(n4402), .B(n4401), .Z(n4406) );
  OR U4624 ( .A(n4404), .B(n4403), .Z(n4405) );
  AND U4625 ( .A(n4406), .B(n4405), .Z(n4426) );
  NAND U4626 ( .A(n31), .B(n4407), .Z(n4409) );
  XOR U4627 ( .A(b[3]), .B(a[191]), .Z(n4430) );
  NAND U4628 ( .A(n5811), .B(n4430), .Z(n4408) );
  AND U4629 ( .A(n4409), .B(n4408), .Z(n4438) );
  NAND U4630 ( .A(b[0]), .B(a[193]), .Z(n4410) );
  XNOR U4631 ( .A(b[1]), .B(n4410), .Z(n4412) );
  NANDN U4632 ( .A(b[0]), .B(a[192]), .Z(n4411) );
  NAND U4633 ( .A(n4412), .B(n4411), .Z(n4437) );
  AND U4634 ( .A(b[3]), .B(a[189]), .Z(n4436) );
  XOR U4635 ( .A(n4437), .B(n4436), .Z(n4439) );
  XOR U4636 ( .A(n4438), .B(n4439), .Z(n4425) );
  NANDN U4637 ( .A(n4414), .B(n4413), .Z(n4418) );
  OR U4638 ( .A(n4416), .B(n4415), .Z(n4417) );
  AND U4639 ( .A(n4418), .B(n4417), .Z(n4424) );
  XOR U4640 ( .A(n4425), .B(n4424), .Z(n4427) );
  XOR U4641 ( .A(n4426), .B(n4427), .Z(n4442) );
  XNOR U4642 ( .A(n4442), .B(sreg[445]), .Z(n4444) );
  NANDN U4643 ( .A(n4419), .B(sreg[444]), .Z(n4423) );
  NAND U4644 ( .A(n4421), .B(n4420), .Z(n4422) );
  NAND U4645 ( .A(n4423), .B(n4422), .Z(n4443) );
  XOR U4646 ( .A(n4444), .B(n4443), .Z(c[445]) );
  NANDN U4647 ( .A(n4425), .B(n4424), .Z(n4429) );
  OR U4648 ( .A(n4427), .B(n4426), .Z(n4428) );
  AND U4649 ( .A(n4429), .B(n4428), .Z(n4449) );
  NAND U4650 ( .A(n31), .B(n4430), .Z(n4432) );
  XOR U4651 ( .A(b[3]), .B(a[192]), .Z(n4453) );
  NAND U4652 ( .A(n5811), .B(n4453), .Z(n4431) );
  AND U4653 ( .A(n4432), .B(n4431), .Z(n4461) );
  NAND U4654 ( .A(b[0]), .B(a[194]), .Z(n4433) );
  XNOR U4655 ( .A(b[1]), .B(n4433), .Z(n4435) );
  NANDN U4656 ( .A(b[0]), .B(a[193]), .Z(n4434) );
  NAND U4657 ( .A(n4435), .B(n4434), .Z(n4460) );
  AND U4658 ( .A(b[3]), .B(a[190]), .Z(n4459) );
  XOR U4659 ( .A(n4460), .B(n4459), .Z(n4462) );
  XOR U4660 ( .A(n4461), .B(n4462), .Z(n4448) );
  NANDN U4661 ( .A(n4437), .B(n4436), .Z(n4441) );
  OR U4662 ( .A(n4439), .B(n4438), .Z(n4440) );
  AND U4663 ( .A(n4441), .B(n4440), .Z(n4447) );
  XOR U4664 ( .A(n4448), .B(n4447), .Z(n4450) );
  XOR U4665 ( .A(n4449), .B(n4450), .Z(n4465) );
  XNOR U4666 ( .A(n4465), .B(sreg[446]), .Z(n4467) );
  NANDN U4667 ( .A(n4442), .B(sreg[445]), .Z(n4446) );
  NAND U4668 ( .A(n4444), .B(n4443), .Z(n4445) );
  NAND U4669 ( .A(n4446), .B(n4445), .Z(n4466) );
  XOR U4670 ( .A(n4467), .B(n4466), .Z(c[446]) );
  NANDN U4671 ( .A(n4448), .B(n4447), .Z(n4452) );
  OR U4672 ( .A(n4450), .B(n4449), .Z(n4451) );
  AND U4673 ( .A(n4452), .B(n4451), .Z(n4472) );
  NAND U4674 ( .A(n31), .B(n4453), .Z(n4455) );
  XOR U4675 ( .A(b[3]), .B(a[193]), .Z(n4476) );
  NAND U4676 ( .A(n5811), .B(n4476), .Z(n4454) );
  AND U4677 ( .A(n4455), .B(n4454), .Z(n4484) );
  AND U4678 ( .A(b[3]), .B(a[191]), .Z(n4482) );
  NAND U4679 ( .A(b[0]), .B(a[195]), .Z(n4456) );
  XNOR U4680 ( .A(b[1]), .B(n4456), .Z(n4458) );
  NANDN U4681 ( .A(b[0]), .B(a[194]), .Z(n4457) );
  NAND U4682 ( .A(n4458), .B(n4457), .Z(n4483) );
  XOR U4683 ( .A(n4482), .B(n4483), .Z(n4485) );
  XOR U4684 ( .A(n4484), .B(n4485), .Z(n4471) );
  NANDN U4685 ( .A(n4460), .B(n4459), .Z(n4464) );
  OR U4686 ( .A(n4462), .B(n4461), .Z(n4463) );
  AND U4687 ( .A(n4464), .B(n4463), .Z(n4470) );
  XOR U4688 ( .A(n4471), .B(n4470), .Z(n4473) );
  XOR U4689 ( .A(n4472), .B(n4473), .Z(n4488) );
  XNOR U4690 ( .A(n4488), .B(sreg[447]), .Z(n4490) );
  NANDN U4691 ( .A(n4465), .B(sreg[446]), .Z(n4469) );
  NAND U4692 ( .A(n4467), .B(n4466), .Z(n4468) );
  NAND U4693 ( .A(n4469), .B(n4468), .Z(n4489) );
  XOR U4694 ( .A(n4490), .B(n4489), .Z(c[447]) );
  NANDN U4695 ( .A(n4471), .B(n4470), .Z(n4475) );
  OR U4696 ( .A(n4473), .B(n4472), .Z(n4474) );
  AND U4697 ( .A(n4475), .B(n4474), .Z(n4495) );
  NAND U4698 ( .A(n31), .B(n4476), .Z(n4478) );
  XOR U4699 ( .A(b[3]), .B(a[194]), .Z(n4499) );
  NAND U4700 ( .A(n5811), .B(n4499), .Z(n4477) );
  AND U4701 ( .A(n4478), .B(n4477), .Z(n4507) );
  NAND U4702 ( .A(b[0]), .B(a[196]), .Z(n4479) );
  XNOR U4703 ( .A(b[1]), .B(n4479), .Z(n4481) );
  NANDN U4704 ( .A(b[0]), .B(a[195]), .Z(n4480) );
  NAND U4705 ( .A(n4481), .B(n4480), .Z(n4506) );
  AND U4706 ( .A(b[3]), .B(a[192]), .Z(n4505) );
  XOR U4707 ( .A(n4506), .B(n4505), .Z(n4508) );
  XOR U4708 ( .A(n4507), .B(n4508), .Z(n4494) );
  NANDN U4709 ( .A(n4483), .B(n4482), .Z(n4487) );
  OR U4710 ( .A(n4485), .B(n4484), .Z(n4486) );
  AND U4711 ( .A(n4487), .B(n4486), .Z(n4493) );
  XOR U4712 ( .A(n4494), .B(n4493), .Z(n4496) );
  XOR U4713 ( .A(n4495), .B(n4496), .Z(n4511) );
  XNOR U4714 ( .A(n4511), .B(sreg[448]), .Z(n4513) );
  NANDN U4715 ( .A(n4488), .B(sreg[447]), .Z(n4492) );
  NAND U4716 ( .A(n4490), .B(n4489), .Z(n4491) );
  NAND U4717 ( .A(n4492), .B(n4491), .Z(n4512) );
  XOR U4718 ( .A(n4513), .B(n4512), .Z(c[448]) );
  NANDN U4719 ( .A(n4494), .B(n4493), .Z(n4498) );
  OR U4720 ( .A(n4496), .B(n4495), .Z(n4497) );
  AND U4721 ( .A(n4498), .B(n4497), .Z(n4518) );
  NAND U4722 ( .A(n31), .B(n4499), .Z(n4501) );
  XOR U4723 ( .A(b[3]), .B(a[195]), .Z(n4522) );
  NAND U4724 ( .A(n5811), .B(n4522), .Z(n4500) );
  AND U4725 ( .A(n4501), .B(n4500), .Z(n4530) );
  AND U4726 ( .A(b[3]), .B(a[193]), .Z(n4528) );
  NAND U4727 ( .A(b[0]), .B(a[197]), .Z(n4502) );
  XNOR U4728 ( .A(b[1]), .B(n4502), .Z(n4504) );
  NANDN U4729 ( .A(b[0]), .B(a[196]), .Z(n4503) );
  NAND U4730 ( .A(n4504), .B(n4503), .Z(n4529) );
  XOR U4731 ( .A(n4528), .B(n4529), .Z(n4531) );
  XOR U4732 ( .A(n4530), .B(n4531), .Z(n4517) );
  NANDN U4733 ( .A(n4506), .B(n4505), .Z(n4510) );
  OR U4734 ( .A(n4508), .B(n4507), .Z(n4509) );
  AND U4735 ( .A(n4510), .B(n4509), .Z(n4516) );
  XOR U4736 ( .A(n4517), .B(n4516), .Z(n4519) );
  XOR U4737 ( .A(n4518), .B(n4519), .Z(n4534) );
  XNOR U4738 ( .A(n4534), .B(sreg[449]), .Z(n4536) );
  NANDN U4739 ( .A(n4511), .B(sreg[448]), .Z(n4515) );
  NAND U4740 ( .A(n4513), .B(n4512), .Z(n4514) );
  NAND U4741 ( .A(n4515), .B(n4514), .Z(n4535) );
  XOR U4742 ( .A(n4536), .B(n4535), .Z(c[449]) );
  NANDN U4743 ( .A(n4517), .B(n4516), .Z(n4521) );
  OR U4744 ( .A(n4519), .B(n4518), .Z(n4520) );
  AND U4745 ( .A(n4521), .B(n4520), .Z(n4541) );
  NAND U4746 ( .A(n31), .B(n4522), .Z(n4524) );
  XOR U4747 ( .A(b[3]), .B(a[196]), .Z(n4545) );
  NAND U4748 ( .A(n5811), .B(n4545), .Z(n4523) );
  AND U4749 ( .A(n4524), .B(n4523), .Z(n4553) );
  NAND U4750 ( .A(b[0]), .B(a[198]), .Z(n4525) );
  XNOR U4751 ( .A(b[1]), .B(n4525), .Z(n4527) );
  NANDN U4752 ( .A(b[0]), .B(a[197]), .Z(n4526) );
  NAND U4753 ( .A(n4527), .B(n4526), .Z(n4552) );
  AND U4754 ( .A(b[3]), .B(a[194]), .Z(n4551) );
  XOR U4755 ( .A(n4552), .B(n4551), .Z(n4554) );
  XOR U4756 ( .A(n4553), .B(n4554), .Z(n4540) );
  NANDN U4757 ( .A(n4529), .B(n4528), .Z(n4533) );
  OR U4758 ( .A(n4531), .B(n4530), .Z(n4532) );
  AND U4759 ( .A(n4533), .B(n4532), .Z(n4539) );
  XOR U4760 ( .A(n4540), .B(n4539), .Z(n4542) );
  XOR U4761 ( .A(n4541), .B(n4542), .Z(n4557) );
  XNOR U4762 ( .A(n4557), .B(sreg[450]), .Z(n4559) );
  NANDN U4763 ( .A(n4534), .B(sreg[449]), .Z(n4538) );
  NAND U4764 ( .A(n4536), .B(n4535), .Z(n4537) );
  NAND U4765 ( .A(n4538), .B(n4537), .Z(n4558) );
  XOR U4766 ( .A(n4559), .B(n4558), .Z(c[450]) );
  NANDN U4767 ( .A(n4540), .B(n4539), .Z(n4544) );
  OR U4768 ( .A(n4542), .B(n4541), .Z(n4543) );
  AND U4769 ( .A(n4544), .B(n4543), .Z(n4564) );
  NAND U4770 ( .A(n31), .B(n4545), .Z(n4547) );
  XOR U4771 ( .A(b[3]), .B(a[197]), .Z(n4568) );
  NAND U4772 ( .A(n5811), .B(n4568), .Z(n4546) );
  AND U4773 ( .A(n4547), .B(n4546), .Z(n4576) );
  AND U4774 ( .A(b[3]), .B(a[195]), .Z(n4574) );
  NAND U4775 ( .A(b[0]), .B(a[199]), .Z(n4548) );
  XNOR U4776 ( .A(b[1]), .B(n4548), .Z(n4550) );
  NANDN U4777 ( .A(b[0]), .B(a[198]), .Z(n4549) );
  NAND U4778 ( .A(n4550), .B(n4549), .Z(n4575) );
  XOR U4779 ( .A(n4574), .B(n4575), .Z(n4577) );
  XOR U4780 ( .A(n4576), .B(n4577), .Z(n4563) );
  NANDN U4781 ( .A(n4552), .B(n4551), .Z(n4556) );
  OR U4782 ( .A(n4554), .B(n4553), .Z(n4555) );
  AND U4783 ( .A(n4556), .B(n4555), .Z(n4562) );
  XOR U4784 ( .A(n4563), .B(n4562), .Z(n4565) );
  XOR U4785 ( .A(n4564), .B(n4565), .Z(n4580) );
  XNOR U4786 ( .A(n4580), .B(sreg[451]), .Z(n4582) );
  NANDN U4787 ( .A(n4557), .B(sreg[450]), .Z(n4561) );
  NAND U4788 ( .A(n4559), .B(n4558), .Z(n4560) );
  NAND U4789 ( .A(n4561), .B(n4560), .Z(n4581) );
  XOR U4790 ( .A(n4582), .B(n4581), .Z(c[451]) );
  NANDN U4791 ( .A(n4563), .B(n4562), .Z(n4567) );
  OR U4792 ( .A(n4565), .B(n4564), .Z(n4566) );
  AND U4793 ( .A(n4567), .B(n4566), .Z(n4587) );
  NAND U4794 ( .A(n31), .B(n4568), .Z(n4570) );
  XOR U4795 ( .A(b[3]), .B(a[198]), .Z(n4591) );
  NAND U4796 ( .A(n5811), .B(n4591), .Z(n4569) );
  AND U4797 ( .A(n4570), .B(n4569), .Z(n4599) );
  NAND U4798 ( .A(b[0]), .B(a[200]), .Z(n4571) );
  XNOR U4799 ( .A(b[1]), .B(n4571), .Z(n4573) );
  NANDN U4800 ( .A(b[0]), .B(a[199]), .Z(n4572) );
  NAND U4801 ( .A(n4573), .B(n4572), .Z(n4598) );
  AND U4802 ( .A(b[3]), .B(a[196]), .Z(n4597) );
  XOR U4803 ( .A(n4598), .B(n4597), .Z(n4600) );
  XOR U4804 ( .A(n4599), .B(n4600), .Z(n4586) );
  NANDN U4805 ( .A(n4575), .B(n4574), .Z(n4579) );
  OR U4806 ( .A(n4577), .B(n4576), .Z(n4578) );
  AND U4807 ( .A(n4579), .B(n4578), .Z(n4585) );
  XOR U4808 ( .A(n4586), .B(n4585), .Z(n4588) );
  XOR U4809 ( .A(n4587), .B(n4588), .Z(n4603) );
  XNOR U4810 ( .A(n4603), .B(sreg[452]), .Z(n4605) );
  NANDN U4811 ( .A(n4580), .B(sreg[451]), .Z(n4584) );
  NAND U4812 ( .A(n4582), .B(n4581), .Z(n4583) );
  NAND U4813 ( .A(n4584), .B(n4583), .Z(n4604) );
  XOR U4814 ( .A(n4605), .B(n4604), .Z(c[452]) );
  NANDN U4815 ( .A(n4586), .B(n4585), .Z(n4590) );
  OR U4816 ( .A(n4588), .B(n4587), .Z(n4589) );
  AND U4817 ( .A(n4590), .B(n4589), .Z(n4610) );
  NAND U4818 ( .A(n31), .B(n4591), .Z(n4593) );
  XOR U4819 ( .A(b[3]), .B(a[199]), .Z(n4614) );
  NAND U4820 ( .A(n5811), .B(n4614), .Z(n4592) );
  AND U4821 ( .A(n4593), .B(n4592), .Z(n4622) );
  NAND U4822 ( .A(b[0]), .B(a[201]), .Z(n4594) );
  XNOR U4823 ( .A(b[1]), .B(n4594), .Z(n4596) );
  NANDN U4824 ( .A(b[0]), .B(a[200]), .Z(n4595) );
  NAND U4825 ( .A(n4596), .B(n4595), .Z(n4621) );
  AND U4826 ( .A(b[3]), .B(a[197]), .Z(n4620) );
  XOR U4827 ( .A(n4621), .B(n4620), .Z(n4623) );
  XOR U4828 ( .A(n4622), .B(n4623), .Z(n4609) );
  NANDN U4829 ( .A(n4598), .B(n4597), .Z(n4602) );
  OR U4830 ( .A(n4600), .B(n4599), .Z(n4601) );
  AND U4831 ( .A(n4602), .B(n4601), .Z(n4608) );
  XOR U4832 ( .A(n4609), .B(n4608), .Z(n4611) );
  XOR U4833 ( .A(n4610), .B(n4611), .Z(n4626) );
  XNOR U4834 ( .A(n4626), .B(sreg[453]), .Z(n4628) );
  NANDN U4835 ( .A(n4603), .B(sreg[452]), .Z(n4607) );
  NAND U4836 ( .A(n4605), .B(n4604), .Z(n4606) );
  NAND U4837 ( .A(n4607), .B(n4606), .Z(n4627) );
  XOR U4838 ( .A(n4628), .B(n4627), .Z(c[453]) );
  NANDN U4839 ( .A(n4609), .B(n4608), .Z(n4613) );
  OR U4840 ( .A(n4611), .B(n4610), .Z(n4612) );
  AND U4841 ( .A(n4613), .B(n4612), .Z(n4633) );
  NAND U4842 ( .A(n31), .B(n4614), .Z(n4616) );
  XOR U4843 ( .A(b[3]), .B(a[200]), .Z(n4637) );
  NAND U4844 ( .A(n5811), .B(n4637), .Z(n4615) );
  AND U4845 ( .A(n4616), .B(n4615), .Z(n4645) );
  NAND U4846 ( .A(b[0]), .B(a[202]), .Z(n4617) );
  XNOR U4847 ( .A(b[1]), .B(n4617), .Z(n4619) );
  NANDN U4848 ( .A(b[0]), .B(a[201]), .Z(n4618) );
  NAND U4849 ( .A(n4619), .B(n4618), .Z(n4644) );
  AND U4850 ( .A(b[3]), .B(a[198]), .Z(n4643) );
  XOR U4851 ( .A(n4644), .B(n4643), .Z(n4646) );
  XOR U4852 ( .A(n4645), .B(n4646), .Z(n4632) );
  NANDN U4853 ( .A(n4621), .B(n4620), .Z(n4625) );
  OR U4854 ( .A(n4623), .B(n4622), .Z(n4624) );
  AND U4855 ( .A(n4625), .B(n4624), .Z(n4631) );
  XOR U4856 ( .A(n4632), .B(n4631), .Z(n4634) );
  XOR U4857 ( .A(n4633), .B(n4634), .Z(n4649) );
  XNOR U4858 ( .A(n4649), .B(sreg[454]), .Z(n4651) );
  NANDN U4859 ( .A(n4626), .B(sreg[453]), .Z(n4630) );
  NAND U4860 ( .A(n4628), .B(n4627), .Z(n4629) );
  NAND U4861 ( .A(n4630), .B(n4629), .Z(n4650) );
  XOR U4862 ( .A(n4651), .B(n4650), .Z(c[454]) );
  NANDN U4863 ( .A(n4632), .B(n4631), .Z(n4636) );
  OR U4864 ( .A(n4634), .B(n4633), .Z(n4635) );
  AND U4865 ( .A(n4636), .B(n4635), .Z(n4656) );
  NAND U4866 ( .A(n31), .B(n4637), .Z(n4639) );
  XOR U4867 ( .A(b[3]), .B(a[201]), .Z(n4660) );
  NAND U4868 ( .A(n5811), .B(n4660), .Z(n4638) );
  AND U4869 ( .A(n4639), .B(n4638), .Z(n4668) );
  NAND U4870 ( .A(b[0]), .B(a[203]), .Z(n4640) );
  XNOR U4871 ( .A(b[1]), .B(n4640), .Z(n4642) );
  NANDN U4872 ( .A(b[0]), .B(a[202]), .Z(n4641) );
  NAND U4873 ( .A(n4642), .B(n4641), .Z(n4667) );
  AND U4874 ( .A(b[3]), .B(a[199]), .Z(n4666) );
  XOR U4875 ( .A(n4667), .B(n4666), .Z(n4669) );
  XOR U4876 ( .A(n4668), .B(n4669), .Z(n4655) );
  NANDN U4877 ( .A(n4644), .B(n4643), .Z(n4648) );
  OR U4878 ( .A(n4646), .B(n4645), .Z(n4647) );
  AND U4879 ( .A(n4648), .B(n4647), .Z(n4654) );
  XOR U4880 ( .A(n4655), .B(n4654), .Z(n4657) );
  XOR U4881 ( .A(n4656), .B(n4657), .Z(n4672) );
  XNOR U4882 ( .A(n4672), .B(sreg[455]), .Z(n4674) );
  NANDN U4883 ( .A(n4649), .B(sreg[454]), .Z(n4653) );
  NAND U4884 ( .A(n4651), .B(n4650), .Z(n4652) );
  NAND U4885 ( .A(n4653), .B(n4652), .Z(n4673) );
  XOR U4886 ( .A(n4674), .B(n4673), .Z(c[455]) );
  NANDN U4887 ( .A(n4655), .B(n4654), .Z(n4659) );
  OR U4888 ( .A(n4657), .B(n4656), .Z(n4658) );
  AND U4889 ( .A(n4659), .B(n4658), .Z(n4679) );
  NAND U4890 ( .A(n31), .B(n4660), .Z(n4662) );
  XOR U4891 ( .A(b[3]), .B(a[202]), .Z(n4683) );
  NAND U4892 ( .A(n5811), .B(n4683), .Z(n4661) );
  AND U4893 ( .A(n4662), .B(n4661), .Z(n4691) );
  AND U4894 ( .A(b[3]), .B(a[200]), .Z(n4689) );
  NAND U4895 ( .A(b[0]), .B(a[204]), .Z(n4663) );
  XNOR U4896 ( .A(b[1]), .B(n4663), .Z(n4665) );
  NANDN U4897 ( .A(b[0]), .B(a[203]), .Z(n4664) );
  NAND U4898 ( .A(n4665), .B(n4664), .Z(n4690) );
  XOR U4899 ( .A(n4689), .B(n4690), .Z(n4692) );
  XOR U4900 ( .A(n4691), .B(n4692), .Z(n4678) );
  NANDN U4901 ( .A(n4667), .B(n4666), .Z(n4671) );
  OR U4902 ( .A(n4669), .B(n4668), .Z(n4670) );
  AND U4903 ( .A(n4671), .B(n4670), .Z(n4677) );
  XOR U4904 ( .A(n4678), .B(n4677), .Z(n4680) );
  XOR U4905 ( .A(n4679), .B(n4680), .Z(n4695) );
  XNOR U4906 ( .A(n4695), .B(sreg[456]), .Z(n4697) );
  NANDN U4907 ( .A(n4672), .B(sreg[455]), .Z(n4676) );
  NAND U4908 ( .A(n4674), .B(n4673), .Z(n4675) );
  NAND U4909 ( .A(n4676), .B(n4675), .Z(n4696) );
  XOR U4910 ( .A(n4697), .B(n4696), .Z(c[456]) );
  NANDN U4911 ( .A(n4678), .B(n4677), .Z(n4682) );
  OR U4912 ( .A(n4680), .B(n4679), .Z(n4681) );
  AND U4913 ( .A(n4682), .B(n4681), .Z(n4702) );
  NAND U4914 ( .A(n31), .B(n4683), .Z(n4685) );
  XOR U4915 ( .A(b[3]), .B(a[203]), .Z(n4706) );
  NAND U4916 ( .A(n5811), .B(n4706), .Z(n4684) );
  AND U4917 ( .A(n4685), .B(n4684), .Z(n4714) );
  NAND U4918 ( .A(b[0]), .B(a[205]), .Z(n4686) );
  XNOR U4919 ( .A(b[1]), .B(n4686), .Z(n4688) );
  NANDN U4920 ( .A(b[0]), .B(a[204]), .Z(n4687) );
  NAND U4921 ( .A(n4688), .B(n4687), .Z(n4713) );
  AND U4922 ( .A(b[3]), .B(a[201]), .Z(n4712) );
  XOR U4923 ( .A(n4713), .B(n4712), .Z(n4715) );
  XOR U4924 ( .A(n4714), .B(n4715), .Z(n4701) );
  NANDN U4925 ( .A(n4690), .B(n4689), .Z(n4694) );
  OR U4926 ( .A(n4692), .B(n4691), .Z(n4693) );
  AND U4927 ( .A(n4694), .B(n4693), .Z(n4700) );
  XOR U4928 ( .A(n4701), .B(n4700), .Z(n4703) );
  XOR U4929 ( .A(n4702), .B(n4703), .Z(n4718) );
  XNOR U4930 ( .A(n4718), .B(sreg[457]), .Z(n4720) );
  NANDN U4931 ( .A(n4695), .B(sreg[456]), .Z(n4699) );
  NAND U4932 ( .A(n4697), .B(n4696), .Z(n4698) );
  NAND U4933 ( .A(n4699), .B(n4698), .Z(n4719) );
  XOR U4934 ( .A(n4720), .B(n4719), .Z(c[457]) );
  NANDN U4935 ( .A(n4701), .B(n4700), .Z(n4705) );
  OR U4936 ( .A(n4703), .B(n4702), .Z(n4704) );
  AND U4937 ( .A(n4705), .B(n4704), .Z(n4725) );
  NAND U4938 ( .A(n31), .B(n4706), .Z(n4708) );
  XOR U4939 ( .A(b[3]), .B(a[204]), .Z(n4729) );
  NAND U4940 ( .A(n5811), .B(n4729), .Z(n4707) );
  AND U4941 ( .A(n4708), .B(n4707), .Z(n4737) );
  AND U4942 ( .A(b[3]), .B(a[202]), .Z(n4735) );
  NAND U4943 ( .A(b[0]), .B(a[206]), .Z(n4709) );
  XNOR U4944 ( .A(b[1]), .B(n4709), .Z(n4711) );
  NANDN U4945 ( .A(b[0]), .B(a[205]), .Z(n4710) );
  NAND U4946 ( .A(n4711), .B(n4710), .Z(n4736) );
  XOR U4947 ( .A(n4735), .B(n4736), .Z(n4738) );
  XOR U4948 ( .A(n4737), .B(n4738), .Z(n4724) );
  NANDN U4949 ( .A(n4713), .B(n4712), .Z(n4717) );
  OR U4950 ( .A(n4715), .B(n4714), .Z(n4716) );
  AND U4951 ( .A(n4717), .B(n4716), .Z(n4723) );
  XOR U4952 ( .A(n4724), .B(n4723), .Z(n4726) );
  XOR U4953 ( .A(n4725), .B(n4726), .Z(n4741) );
  XNOR U4954 ( .A(n4741), .B(sreg[458]), .Z(n4743) );
  NANDN U4955 ( .A(n4718), .B(sreg[457]), .Z(n4722) );
  NAND U4956 ( .A(n4720), .B(n4719), .Z(n4721) );
  NAND U4957 ( .A(n4722), .B(n4721), .Z(n4742) );
  XOR U4958 ( .A(n4743), .B(n4742), .Z(c[458]) );
  NANDN U4959 ( .A(n4724), .B(n4723), .Z(n4728) );
  OR U4960 ( .A(n4726), .B(n4725), .Z(n4727) );
  AND U4961 ( .A(n4728), .B(n4727), .Z(n4748) );
  NAND U4962 ( .A(n31), .B(n4729), .Z(n4731) );
  XOR U4963 ( .A(b[3]), .B(a[205]), .Z(n4752) );
  NAND U4964 ( .A(n5811), .B(n4752), .Z(n4730) );
  AND U4965 ( .A(n4731), .B(n4730), .Z(n4760) );
  NAND U4966 ( .A(b[0]), .B(a[207]), .Z(n4732) );
  XNOR U4967 ( .A(b[1]), .B(n4732), .Z(n4734) );
  NANDN U4968 ( .A(b[0]), .B(a[206]), .Z(n4733) );
  NAND U4969 ( .A(n4734), .B(n4733), .Z(n4759) );
  AND U4970 ( .A(b[3]), .B(a[203]), .Z(n4758) );
  XOR U4971 ( .A(n4759), .B(n4758), .Z(n4761) );
  XOR U4972 ( .A(n4760), .B(n4761), .Z(n4747) );
  NANDN U4973 ( .A(n4736), .B(n4735), .Z(n4740) );
  OR U4974 ( .A(n4738), .B(n4737), .Z(n4739) );
  AND U4975 ( .A(n4740), .B(n4739), .Z(n4746) );
  XOR U4976 ( .A(n4747), .B(n4746), .Z(n4749) );
  XOR U4977 ( .A(n4748), .B(n4749), .Z(n4764) );
  XNOR U4978 ( .A(n4764), .B(sreg[459]), .Z(n4766) );
  NANDN U4979 ( .A(n4741), .B(sreg[458]), .Z(n4745) );
  NAND U4980 ( .A(n4743), .B(n4742), .Z(n4744) );
  NAND U4981 ( .A(n4745), .B(n4744), .Z(n4765) );
  XOR U4982 ( .A(n4766), .B(n4765), .Z(c[459]) );
  NANDN U4983 ( .A(n4747), .B(n4746), .Z(n4751) );
  OR U4984 ( .A(n4749), .B(n4748), .Z(n4750) );
  AND U4985 ( .A(n4751), .B(n4750), .Z(n4771) );
  NAND U4986 ( .A(n31), .B(n4752), .Z(n4754) );
  XOR U4987 ( .A(b[3]), .B(a[206]), .Z(n4775) );
  NAND U4988 ( .A(n5811), .B(n4775), .Z(n4753) );
  AND U4989 ( .A(n4754), .B(n4753), .Z(n4783) );
  NAND U4990 ( .A(b[0]), .B(a[208]), .Z(n4755) );
  XNOR U4991 ( .A(b[1]), .B(n4755), .Z(n4757) );
  NANDN U4992 ( .A(b[0]), .B(a[207]), .Z(n4756) );
  NAND U4993 ( .A(n4757), .B(n4756), .Z(n4782) );
  AND U4994 ( .A(b[3]), .B(a[204]), .Z(n4781) );
  XOR U4995 ( .A(n4782), .B(n4781), .Z(n4784) );
  XOR U4996 ( .A(n4783), .B(n4784), .Z(n4770) );
  NANDN U4997 ( .A(n4759), .B(n4758), .Z(n4763) );
  OR U4998 ( .A(n4761), .B(n4760), .Z(n4762) );
  AND U4999 ( .A(n4763), .B(n4762), .Z(n4769) );
  XOR U5000 ( .A(n4770), .B(n4769), .Z(n4772) );
  XOR U5001 ( .A(n4771), .B(n4772), .Z(n4787) );
  XNOR U5002 ( .A(n4787), .B(sreg[460]), .Z(n4789) );
  NANDN U5003 ( .A(n4764), .B(sreg[459]), .Z(n4768) );
  NAND U5004 ( .A(n4766), .B(n4765), .Z(n4767) );
  NAND U5005 ( .A(n4768), .B(n4767), .Z(n4788) );
  XOR U5006 ( .A(n4789), .B(n4788), .Z(c[460]) );
  NANDN U5007 ( .A(n4770), .B(n4769), .Z(n4774) );
  OR U5008 ( .A(n4772), .B(n4771), .Z(n4773) );
  AND U5009 ( .A(n4774), .B(n4773), .Z(n4794) );
  NAND U5010 ( .A(n31), .B(n4775), .Z(n4777) );
  XOR U5011 ( .A(b[3]), .B(a[207]), .Z(n4798) );
  NAND U5012 ( .A(n5811), .B(n4798), .Z(n4776) );
  AND U5013 ( .A(n4777), .B(n4776), .Z(n4806) );
  NAND U5014 ( .A(b[0]), .B(a[209]), .Z(n4778) );
  XNOR U5015 ( .A(b[1]), .B(n4778), .Z(n4780) );
  NANDN U5016 ( .A(b[0]), .B(a[208]), .Z(n4779) );
  NAND U5017 ( .A(n4780), .B(n4779), .Z(n4805) );
  AND U5018 ( .A(b[3]), .B(a[205]), .Z(n4804) );
  XOR U5019 ( .A(n4805), .B(n4804), .Z(n4807) );
  XOR U5020 ( .A(n4806), .B(n4807), .Z(n4793) );
  NANDN U5021 ( .A(n4782), .B(n4781), .Z(n4786) );
  OR U5022 ( .A(n4784), .B(n4783), .Z(n4785) );
  AND U5023 ( .A(n4786), .B(n4785), .Z(n4792) );
  XOR U5024 ( .A(n4793), .B(n4792), .Z(n4795) );
  XOR U5025 ( .A(n4794), .B(n4795), .Z(n4810) );
  XNOR U5026 ( .A(n4810), .B(sreg[461]), .Z(n4812) );
  NANDN U5027 ( .A(n4787), .B(sreg[460]), .Z(n4791) );
  NAND U5028 ( .A(n4789), .B(n4788), .Z(n4790) );
  NAND U5029 ( .A(n4791), .B(n4790), .Z(n4811) );
  XOR U5030 ( .A(n4812), .B(n4811), .Z(c[461]) );
  NANDN U5031 ( .A(n4793), .B(n4792), .Z(n4797) );
  OR U5032 ( .A(n4795), .B(n4794), .Z(n4796) );
  AND U5033 ( .A(n4797), .B(n4796), .Z(n4817) );
  NAND U5034 ( .A(n31), .B(n4798), .Z(n4800) );
  XOR U5035 ( .A(b[3]), .B(a[208]), .Z(n4821) );
  NAND U5036 ( .A(n5811), .B(n4821), .Z(n4799) );
  AND U5037 ( .A(n4800), .B(n4799), .Z(n4829) );
  AND U5038 ( .A(b[3]), .B(a[206]), .Z(n4827) );
  NAND U5039 ( .A(b[0]), .B(a[210]), .Z(n4801) );
  XNOR U5040 ( .A(b[1]), .B(n4801), .Z(n4803) );
  NANDN U5041 ( .A(b[0]), .B(a[209]), .Z(n4802) );
  NAND U5042 ( .A(n4803), .B(n4802), .Z(n4828) );
  XOR U5043 ( .A(n4827), .B(n4828), .Z(n4830) );
  XOR U5044 ( .A(n4829), .B(n4830), .Z(n4816) );
  NANDN U5045 ( .A(n4805), .B(n4804), .Z(n4809) );
  OR U5046 ( .A(n4807), .B(n4806), .Z(n4808) );
  AND U5047 ( .A(n4809), .B(n4808), .Z(n4815) );
  XOR U5048 ( .A(n4816), .B(n4815), .Z(n4818) );
  XOR U5049 ( .A(n4817), .B(n4818), .Z(n4833) );
  XNOR U5050 ( .A(n4833), .B(sreg[462]), .Z(n4835) );
  NANDN U5051 ( .A(n4810), .B(sreg[461]), .Z(n4814) );
  NAND U5052 ( .A(n4812), .B(n4811), .Z(n4813) );
  NAND U5053 ( .A(n4814), .B(n4813), .Z(n4834) );
  XOR U5054 ( .A(n4835), .B(n4834), .Z(c[462]) );
  NANDN U5055 ( .A(n4816), .B(n4815), .Z(n4820) );
  OR U5056 ( .A(n4818), .B(n4817), .Z(n4819) );
  AND U5057 ( .A(n4820), .B(n4819), .Z(n4840) );
  NAND U5058 ( .A(n31), .B(n4821), .Z(n4823) );
  XOR U5059 ( .A(b[3]), .B(a[209]), .Z(n4844) );
  NAND U5060 ( .A(n5811), .B(n4844), .Z(n4822) );
  AND U5061 ( .A(n4823), .B(n4822), .Z(n4852) );
  NAND U5062 ( .A(b[0]), .B(a[211]), .Z(n4824) );
  XNOR U5063 ( .A(b[1]), .B(n4824), .Z(n4826) );
  NANDN U5064 ( .A(b[0]), .B(a[210]), .Z(n4825) );
  NAND U5065 ( .A(n4826), .B(n4825), .Z(n4851) );
  AND U5066 ( .A(b[3]), .B(a[207]), .Z(n4850) );
  XOR U5067 ( .A(n4851), .B(n4850), .Z(n4853) );
  XOR U5068 ( .A(n4852), .B(n4853), .Z(n4839) );
  NANDN U5069 ( .A(n4828), .B(n4827), .Z(n4832) );
  OR U5070 ( .A(n4830), .B(n4829), .Z(n4831) );
  AND U5071 ( .A(n4832), .B(n4831), .Z(n4838) );
  XOR U5072 ( .A(n4839), .B(n4838), .Z(n4841) );
  XOR U5073 ( .A(n4840), .B(n4841), .Z(n4856) );
  XNOR U5074 ( .A(n4856), .B(sreg[463]), .Z(n4858) );
  NANDN U5075 ( .A(n4833), .B(sreg[462]), .Z(n4837) );
  NAND U5076 ( .A(n4835), .B(n4834), .Z(n4836) );
  NAND U5077 ( .A(n4837), .B(n4836), .Z(n4857) );
  XOR U5078 ( .A(n4858), .B(n4857), .Z(c[463]) );
  NANDN U5079 ( .A(n4839), .B(n4838), .Z(n4843) );
  OR U5080 ( .A(n4841), .B(n4840), .Z(n4842) );
  AND U5081 ( .A(n4843), .B(n4842), .Z(n4863) );
  NAND U5082 ( .A(n31), .B(n4844), .Z(n4846) );
  XOR U5083 ( .A(b[3]), .B(a[210]), .Z(n4867) );
  NAND U5084 ( .A(n5811), .B(n4867), .Z(n4845) );
  AND U5085 ( .A(n4846), .B(n4845), .Z(n4875) );
  AND U5086 ( .A(b[3]), .B(a[208]), .Z(n4873) );
  NAND U5087 ( .A(b[0]), .B(a[212]), .Z(n4847) );
  XNOR U5088 ( .A(b[1]), .B(n4847), .Z(n4849) );
  NANDN U5089 ( .A(b[0]), .B(a[211]), .Z(n4848) );
  NAND U5090 ( .A(n4849), .B(n4848), .Z(n4874) );
  XOR U5091 ( .A(n4873), .B(n4874), .Z(n4876) );
  XOR U5092 ( .A(n4875), .B(n4876), .Z(n4862) );
  NANDN U5093 ( .A(n4851), .B(n4850), .Z(n4855) );
  OR U5094 ( .A(n4853), .B(n4852), .Z(n4854) );
  AND U5095 ( .A(n4855), .B(n4854), .Z(n4861) );
  XOR U5096 ( .A(n4862), .B(n4861), .Z(n4864) );
  XOR U5097 ( .A(n4863), .B(n4864), .Z(n4879) );
  XNOR U5098 ( .A(n4879), .B(sreg[464]), .Z(n4881) );
  NANDN U5099 ( .A(n4856), .B(sreg[463]), .Z(n4860) );
  NAND U5100 ( .A(n4858), .B(n4857), .Z(n4859) );
  NAND U5101 ( .A(n4860), .B(n4859), .Z(n4880) );
  XOR U5102 ( .A(n4881), .B(n4880), .Z(c[464]) );
  NANDN U5103 ( .A(n4862), .B(n4861), .Z(n4866) );
  OR U5104 ( .A(n4864), .B(n4863), .Z(n4865) );
  AND U5105 ( .A(n4866), .B(n4865), .Z(n4886) );
  NAND U5106 ( .A(n31), .B(n4867), .Z(n4869) );
  XOR U5107 ( .A(b[3]), .B(a[211]), .Z(n4890) );
  NAND U5108 ( .A(n5811), .B(n4890), .Z(n4868) );
  AND U5109 ( .A(n4869), .B(n4868), .Z(n4898) );
  NAND U5110 ( .A(b[0]), .B(a[213]), .Z(n4870) );
  XNOR U5111 ( .A(b[1]), .B(n4870), .Z(n4872) );
  NANDN U5112 ( .A(b[0]), .B(a[212]), .Z(n4871) );
  NAND U5113 ( .A(n4872), .B(n4871), .Z(n4897) );
  AND U5114 ( .A(b[3]), .B(a[209]), .Z(n4896) );
  XOR U5115 ( .A(n4897), .B(n4896), .Z(n4899) );
  XOR U5116 ( .A(n4898), .B(n4899), .Z(n4885) );
  NANDN U5117 ( .A(n4874), .B(n4873), .Z(n4878) );
  OR U5118 ( .A(n4876), .B(n4875), .Z(n4877) );
  AND U5119 ( .A(n4878), .B(n4877), .Z(n4884) );
  XOR U5120 ( .A(n4885), .B(n4884), .Z(n4887) );
  XOR U5121 ( .A(n4886), .B(n4887), .Z(n4902) );
  XNOR U5122 ( .A(n4902), .B(sreg[465]), .Z(n4904) );
  NANDN U5123 ( .A(n4879), .B(sreg[464]), .Z(n4883) );
  NAND U5124 ( .A(n4881), .B(n4880), .Z(n4882) );
  NAND U5125 ( .A(n4883), .B(n4882), .Z(n4903) );
  XOR U5126 ( .A(n4904), .B(n4903), .Z(c[465]) );
  NANDN U5127 ( .A(n4885), .B(n4884), .Z(n4889) );
  OR U5128 ( .A(n4887), .B(n4886), .Z(n4888) );
  AND U5129 ( .A(n4889), .B(n4888), .Z(n4909) );
  NAND U5130 ( .A(n31), .B(n4890), .Z(n4892) );
  XOR U5131 ( .A(b[3]), .B(a[212]), .Z(n4913) );
  NAND U5132 ( .A(n5811), .B(n4913), .Z(n4891) );
  AND U5133 ( .A(n4892), .B(n4891), .Z(n4921) );
  NAND U5134 ( .A(b[0]), .B(a[214]), .Z(n4893) );
  XNOR U5135 ( .A(b[1]), .B(n4893), .Z(n4895) );
  NANDN U5136 ( .A(b[0]), .B(a[213]), .Z(n4894) );
  NAND U5137 ( .A(n4895), .B(n4894), .Z(n4920) );
  AND U5138 ( .A(b[3]), .B(a[210]), .Z(n4919) );
  XOR U5139 ( .A(n4920), .B(n4919), .Z(n4922) );
  XOR U5140 ( .A(n4921), .B(n4922), .Z(n4908) );
  NANDN U5141 ( .A(n4897), .B(n4896), .Z(n4901) );
  OR U5142 ( .A(n4899), .B(n4898), .Z(n4900) );
  AND U5143 ( .A(n4901), .B(n4900), .Z(n4907) );
  XOR U5144 ( .A(n4908), .B(n4907), .Z(n4910) );
  XOR U5145 ( .A(n4909), .B(n4910), .Z(n4925) );
  XNOR U5146 ( .A(n4925), .B(sreg[466]), .Z(n4927) );
  NANDN U5147 ( .A(n4902), .B(sreg[465]), .Z(n4906) );
  NAND U5148 ( .A(n4904), .B(n4903), .Z(n4905) );
  NAND U5149 ( .A(n4906), .B(n4905), .Z(n4926) );
  XOR U5150 ( .A(n4927), .B(n4926), .Z(c[466]) );
  NANDN U5151 ( .A(n4908), .B(n4907), .Z(n4912) );
  OR U5152 ( .A(n4910), .B(n4909), .Z(n4911) );
  AND U5153 ( .A(n4912), .B(n4911), .Z(n4932) );
  NAND U5154 ( .A(n31), .B(n4913), .Z(n4915) );
  XOR U5155 ( .A(b[3]), .B(a[213]), .Z(n4936) );
  NAND U5156 ( .A(n5811), .B(n4936), .Z(n4914) );
  AND U5157 ( .A(n4915), .B(n4914), .Z(n4944) );
  AND U5158 ( .A(b[3]), .B(a[211]), .Z(n4942) );
  NAND U5159 ( .A(b[0]), .B(a[215]), .Z(n4916) );
  XNOR U5160 ( .A(b[1]), .B(n4916), .Z(n4918) );
  NANDN U5161 ( .A(b[0]), .B(a[214]), .Z(n4917) );
  NAND U5162 ( .A(n4918), .B(n4917), .Z(n4943) );
  XOR U5163 ( .A(n4942), .B(n4943), .Z(n4945) );
  XOR U5164 ( .A(n4944), .B(n4945), .Z(n4931) );
  NANDN U5165 ( .A(n4920), .B(n4919), .Z(n4924) );
  OR U5166 ( .A(n4922), .B(n4921), .Z(n4923) );
  AND U5167 ( .A(n4924), .B(n4923), .Z(n4930) );
  XOR U5168 ( .A(n4931), .B(n4930), .Z(n4933) );
  XOR U5169 ( .A(n4932), .B(n4933), .Z(n4948) );
  XNOR U5170 ( .A(n4948), .B(sreg[467]), .Z(n4950) );
  NANDN U5171 ( .A(n4925), .B(sreg[466]), .Z(n4929) );
  NAND U5172 ( .A(n4927), .B(n4926), .Z(n4928) );
  NAND U5173 ( .A(n4929), .B(n4928), .Z(n4949) );
  XOR U5174 ( .A(n4950), .B(n4949), .Z(c[467]) );
  NANDN U5175 ( .A(n4931), .B(n4930), .Z(n4935) );
  OR U5176 ( .A(n4933), .B(n4932), .Z(n4934) );
  AND U5177 ( .A(n4935), .B(n4934), .Z(n4955) );
  NAND U5178 ( .A(n31), .B(n4936), .Z(n4938) );
  XOR U5179 ( .A(b[3]), .B(a[214]), .Z(n4959) );
  NAND U5180 ( .A(n5811), .B(n4959), .Z(n4937) );
  AND U5181 ( .A(n4938), .B(n4937), .Z(n4967) );
  NAND U5182 ( .A(b[0]), .B(a[216]), .Z(n4939) );
  XNOR U5183 ( .A(b[1]), .B(n4939), .Z(n4941) );
  NANDN U5184 ( .A(b[0]), .B(a[215]), .Z(n4940) );
  NAND U5185 ( .A(n4941), .B(n4940), .Z(n4966) );
  AND U5186 ( .A(b[3]), .B(a[212]), .Z(n4965) );
  XOR U5187 ( .A(n4966), .B(n4965), .Z(n4968) );
  XOR U5188 ( .A(n4967), .B(n4968), .Z(n4954) );
  NANDN U5189 ( .A(n4943), .B(n4942), .Z(n4947) );
  OR U5190 ( .A(n4945), .B(n4944), .Z(n4946) );
  AND U5191 ( .A(n4947), .B(n4946), .Z(n4953) );
  XOR U5192 ( .A(n4954), .B(n4953), .Z(n4956) );
  XOR U5193 ( .A(n4955), .B(n4956), .Z(n4971) );
  XNOR U5194 ( .A(n4971), .B(sreg[468]), .Z(n4973) );
  NANDN U5195 ( .A(n4948), .B(sreg[467]), .Z(n4952) );
  NAND U5196 ( .A(n4950), .B(n4949), .Z(n4951) );
  NAND U5197 ( .A(n4952), .B(n4951), .Z(n4972) );
  XOR U5198 ( .A(n4973), .B(n4972), .Z(c[468]) );
  NANDN U5199 ( .A(n4954), .B(n4953), .Z(n4958) );
  OR U5200 ( .A(n4956), .B(n4955), .Z(n4957) );
  AND U5201 ( .A(n4958), .B(n4957), .Z(n4978) );
  NAND U5202 ( .A(n31), .B(n4959), .Z(n4961) );
  XOR U5203 ( .A(b[3]), .B(a[215]), .Z(n4982) );
  NAND U5204 ( .A(n5811), .B(n4982), .Z(n4960) );
  AND U5205 ( .A(n4961), .B(n4960), .Z(n4990) );
  AND U5206 ( .A(b[3]), .B(a[213]), .Z(n4988) );
  NAND U5207 ( .A(b[0]), .B(a[217]), .Z(n4962) );
  XNOR U5208 ( .A(b[1]), .B(n4962), .Z(n4964) );
  NANDN U5209 ( .A(b[0]), .B(a[216]), .Z(n4963) );
  NAND U5210 ( .A(n4964), .B(n4963), .Z(n4989) );
  XOR U5211 ( .A(n4988), .B(n4989), .Z(n4991) );
  XOR U5212 ( .A(n4990), .B(n4991), .Z(n4977) );
  NANDN U5213 ( .A(n4966), .B(n4965), .Z(n4970) );
  OR U5214 ( .A(n4968), .B(n4967), .Z(n4969) );
  AND U5215 ( .A(n4970), .B(n4969), .Z(n4976) );
  XOR U5216 ( .A(n4977), .B(n4976), .Z(n4979) );
  XOR U5217 ( .A(n4978), .B(n4979), .Z(n4994) );
  XNOR U5218 ( .A(n4994), .B(sreg[469]), .Z(n4996) );
  NANDN U5219 ( .A(n4971), .B(sreg[468]), .Z(n4975) );
  NAND U5220 ( .A(n4973), .B(n4972), .Z(n4974) );
  NAND U5221 ( .A(n4975), .B(n4974), .Z(n4995) );
  XOR U5222 ( .A(n4996), .B(n4995), .Z(c[469]) );
  NANDN U5223 ( .A(n4977), .B(n4976), .Z(n4981) );
  OR U5224 ( .A(n4979), .B(n4978), .Z(n4980) );
  AND U5225 ( .A(n4981), .B(n4980), .Z(n5001) );
  NAND U5226 ( .A(n31), .B(n4982), .Z(n4984) );
  XOR U5227 ( .A(b[3]), .B(a[216]), .Z(n5005) );
  NAND U5228 ( .A(n5811), .B(n5005), .Z(n4983) );
  AND U5229 ( .A(n4984), .B(n4983), .Z(n5013) );
  NAND U5230 ( .A(b[0]), .B(a[218]), .Z(n4985) );
  XNOR U5231 ( .A(b[1]), .B(n4985), .Z(n4987) );
  NANDN U5232 ( .A(b[0]), .B(a[217]), .Z(n4986) );
  NAND U5233 ( .A(n4987), .B(n4986), .Z(n5012) );
  AND U5234 ( .A(b[3]), .B(a[214]), .Z(n5011) );
  XOR U5235 ( .A(n5012), .B(n5011), .Z(n5014) );
  XOR U5236 ( .A(n5013), .B(n5014), .Z(n5000) );
  NANDN U5237 ( .A(n4989), .B(n4988), .Z(n4993) );
  OR U5238 ( .A(n4991), .B(n4990), .Z(n4992) );
  AND U5239 ( .A(n4993), .B(n4992), .Z(n4999) );
  XOR U5240 ( .A(n5000), .B(n4999), .Z(n5002) );
  XOR U5241 ( .A(n5001), .B(n5002), .Z(n5017) );
  XNOR U5242 ( .A(n5017), .B(sreg[470]), .Z(n5019) );
  NANDN U5243 ( .A(n4994), .B(sreg[469]), .Z(n4998) );
  NAND U5244 ( .A(n4996), .B(n4995), .Z(n4997) );
  NAND U5245 ( .A(n4998), .B(n4997), .Z(n5018) );
  XOR U5246 ( .A(n5019), .B(n5018), .Z(c[470]) );
  NANDN U5247 ( .A(n5000), .B(n4999), .Z(n5004) );
  OR U5248 ( .A(n5002), .B(n5001), .Z(n5003) );
  AND U5249 ( .A(n5004), .B(n5003), .Z(n5024) );
  NAND U5250 ( .A(n31), .B(n5005), .Z(n5007) );
  XOR U5251 ( .A(b[3]), .B(a[217]), .Z(n5028) );
  NAND U5252 ( .A(n5811), .B(n5028), .Z(n5006) );
  AND U5253 ( .A(n5007), .B(n5006), .Z(n5036) );
  NAND U5254 ( .A(b[0]), .B(a[219]), .Z(n5008) );
  XNOR U5255 ( .A(b[1]), .B(n5008), .Z(n5010) );
  NANDN U5256 ( .A(b[0]), .B(a[218]), .Z(n5009) );
  NAND U5257 ( .A(n5010), .B(n5009), .Z(n5035) );
  AND U5258 ( .A(b[3]), .B(a[215]), .Z(n5034) );
  XOR U5259 ( .A(n5035), .B(n5034), .Z(n5037) );
  XOR U5260 ( .A(n5036), .B(n5037), .Z(n5023) );
  NANDN U5261 ( .A(n5012), .B(n5011), .Z(n5016) );
  OR U5262 ( .A(n5014), .B(n5013), .Z(n5015) );
  AND U5263 ( .A(n5016), .B(n5015), .Z(n5022) );
  XOR U5264 ( .A(n5023), .B(n5022), .Z(n5025) );
  XOR U5265 ( .A(n5024), .B(n5025), .Z(n5040) );
  XNOR U5266 ( .A(n5040), .B(sreg[471]), .Z(n5042) );
  NANDN U5267 ( .A(n5017), .B(sreg[470]), .Z(n5021) );
  NAND U5268 ( .A(n5019), .B(n5018), .Z(n5020) );
  NAND U5269 ( .A(n5021), .B(n5020), .Z(n5041) );
  XOR U5270 ( .A(n5042), .B(n5041), .Z(c[471]) );
  NANDN U5271 ( .A(n5023), .B(n5022), .Z(n5027) );
  OR U5272 ( .A(n5025), .B(n5024), .Z(n5026) );
  AND U5273 ( .A(n5027), .B(n5026), .Z(n5047) );
  NAND U5274 ( .A(n31), .B(n5028), .Z(n5030) );
  XOR U5275 ( .A(b[3]), .B(a[218]), .Z(n5051) );
  NAND U5276 ( .A(n5811), .B(n5051), .Z(n5029) );
  AND U5277 ( .A(n5030), .B(n5029), .Z(n5059) );
  NAND U5278 ( .A(b[0]), .B(a[220]), .Z(n5031) );
  XNOR U5279 ( .A(b[1]), .B(n5031), .Z(n5033) );
  NANDN U5280 ( .A(b[0]), .B(a[219]), .Z(n5032) );
  NAND U5281 ( .A(n5033), .B(n5032), .Z(n5058) );
  AND U5282 ( .A(b[3]), .B(a[216]), .Z(n5057) );
  XOR U5283 ( .A(n5058), .B(n5057), .Z(n5060) );
  XOR U5284 ( .A(n5059), .B(n5060), .Z(n5046) );
  NANDN U5285 ( .A(n5035), .B(n5034), .Z(n5039) );
  OR U5286 ( .A(n5037), .B(n5036), .Z(n5038) );
  AND U5287 ( .A(n5039), .B(n5038), .Z(n5045) );
  XOR U5288 ( .A(n5046), .B(n5045), .Z(n5048) );
  XOR U5289 ( .A(n5047), .B(n5048), .Z(n5063) );
  XNOR U5290 ( .A(n5063), .B(sreg[472]), .Z(n5065) );
  NANDN U5291 ( .A(n5040), .B(sreg[471]), .Z(n5044) );
  NAND U5292 ( .A(n5042), .B(n5041), .Z(n5043) );
  NAND U5293 ( .A(n5044), .B(n5043), .Z(n5064) );
  XOR U5294 ( .A(n5065), .B(n5064), .Z(c[472]) );
  NANDN U5295 ( .A(n5046), .B(n5045), .Z(n5050) );
  OR U5296 ( .A(n5048), .B(n5047), .Z(n5049) );
  AND U5297 ( .A(n5050), .B(n5049), .Z(n5070) );
  NAND U5298 ( .A(n31), .B(n5051), .Z(n5053) );
  XOR U5299 ( .A(b[3]), .B(a[219]), .Z(n5074) );
  NAND U5300 ( .A(n5811), .B(n5074), .Z(n5052) );
  AND U5301 ( .A(n5053), .B(n5052), .Z(n5082) );
  NAND U5302 ( .A(b[0]), .B(a[221]), .Z(n5054) );
  XNOR U5303 ( .A(b[1]), .B(n5054), .Z(n5056) );
  NANDN U5304 ( .A(b[0]), .B(a[220]), .Z(n5055) );
  NAND U5305 ( .A(n5056), .B(n5055), .Z(n5081) );
  AND U5306 ( .A(b[3]), .B(a[217]), .Z(n5080) );
  XOR U5307 ( .A(n5081), .B(n5080), .Z(n5083) );
  XOR U5308 ( .A(n5082), .B(n5083), .Z(n5069) );
  NANDN U5309 ( .A(n5058), .B(n5057), .Z(n5062) );
  OR U5310 ( .A(n5060), .B(n5059), .Z(n5061) );
  AND U5311 ( .A(n5062), .B(n5061), .Z(n5068) );
  XOR U5312 ( .A(n5069), .B(n5068), .Z(n5071) );
  XOR U5313 ( .A(n5070), .B(n5071), .Z(n5086) );
  XNOR U5314 ( .A(n5086), .B(sreg[473]), .Z(n5088) );
  NANDN U5315 ( .A(n5063), .B(sreg[472]), .Z(n5067) );
  NAND U5316 ( .A(n5065), .B(n5064), .Z(n5066) );
  NAND U5317 ( .A(n5067), .B(n5066), .Z(n5087) );
  XOR U5318 ( .A(n5088), .B(n5087), .Z(c[473]) );
  NANDN U5319 ( .A(n5069), .B(n5068), .Z(n5073) );
  OR U5320 ( .A(n5071), .B(n5070), .Z(n5072) );
  AND U5321 ( .A(n5073), .B(n5072), .Z(n5093) );
  NAND U5322 ( .A(n31), .B(n5074), .Z(n5076) );
  XOR U5323 ( .A(b[3]), .B(a[220]), .Z(n5097) );
  NAND U5324 ( .A(n5811), .B(n5097), .Z(n5075) );
  AND U5325 ( .A(n5076), .B(n5075), .Z(n5105) );
  NAND U5326 ( .A(b[0]), .B(a[222]), .Z(n5077) );
  XNOR U5327 ( .A(b[1]), .B(n5077), .Z(n5079) );
  NANDN U5328 ( .A(b[0]), .B(a[221]), .Z(n5078) );
  NAND U5329 ( .A(n5079), .B(n5078), .Z(n5104) );
  AND U5330 ( .A(b[3]), .B(a[218]), .Z(n5103) );
  XOR U5331 ( .A(n5104), .B(n5103), .Z(n5106) );
  XOR U5332 ( .A(n5105), .B(n5106), .Z(n5092) );
  NANDN U5333 ( .A(n5081), .B(n5080), .Z(n5085) );
  OR U5334 ( .A(n5083), .B(n5082), .Z(n5084) );
  AND U5335 ( .A(n5085), .B(n5084), .Z(n5091) );
  XOR U5336 ( .A(n5092), .B(n5091), .Z(n5094) );
  XOR U5337 ( .A(n5093), .B(n5094), .Z(n5109) );
  XNOR U5338 ( .A(n5109), .B(sreg[474]), .Z(n5111) );
  NANDN U5339 ( .A(n5086), .B(sreg[473]), .Z(n5090) );
  NAND U5340 ( .A(n5088), .B(n5087), .Z(n5089) );
  NAND U5341 ( .A(n5090), .B(n5089), .Z(n5110) );
  XOR U5342 ( .A(n5111), .B(n5110), .Z(c[474]) );
  NANDN U5343 ( .A(n5092), .B(n5091), .Z(n5096) );
  OR U5344 ( .A(n5094), .B(n5093), .Z(n5095) );
  AND U5345 ( .A(n5096), .B(n5095), .Z(n5116) );
  NAND U5346 ( .A(n31), .B(n5097), .Z(n5099) );
  XOR U5347 ( .A(b[3]), .B(a[221]), .Z(n5120) );
  NAND U5348 ( .A(n5811), .B(n5120), .Z(n5098) );
  AND U5349 ( .A(n5099), .B(n5098), .Z(n5128) );
  AND U5350 ( .A(b[3]), .B(a[219]), .Z(n5126) );
  NAND U5351 ( .A(b[0]), .B(a[223]), .Z(n5100) );
  XNOR U5352 ( .A(b[1]), .B(n5100), .Z(n5102) );
  NANDN U5353 ( .A(b[0]), .B(a[222]), .Z(n5101) );
  NAND U5354 ( .A(n5102), .B(n5101), .Z(n5127) );
  XOR U5355 ( .A(n5126), .B(n5127), .Z(n5129) );
  XOR U5356 ( .A(n5128), .B(n5129), .Z(n5115) );
  NANDN U5357 ( .A(n5104), .B(n5103), .Z(n5108) );
  OR U5358 ( .A(n5106), .B(n5105), .Z(n5107) );
  AND U5359 ( .A(n5108), .B(n5107), .Z(n5114) );
  XOR U5360 ( .A(n5115), .B(n5114), .Z(n5117) );
  XOR U5361 ( .A(n5116), .B(n5117), .Z(n5132) );
  XNOR U5362 ( .A(n5132), .B(sreg[475]), .Z(n5134) );
  NANDN U5363 ( .A(n5109), .B(sreg[474]), .Z(n5113) );
  NAND U5364 ( .A(n5111), .B(n5110), .Z(n5112) );
  NAND U5365 ( .A(n5113), .B(n5112), .Z(n5133) );
  XOR U5366 ( .A(n5134), .B(n5133), .Z(c[475]) );
  NANDN U5367 ( .A(n5115), .B(n5114), .Z(n5119) );
  OR U5368 ( .A(n5117), .B(n5116), .Z(n5118) );
  AND U5369 ( .A(n5119), .B(n5118), .Z(n5139) );
  NAND U5370 ( .A(n31), .B(n5120), .Z(n5122) );
  XOR U5371 ( .A(b[3]), .B(a[222]), .Z(n5143) );
  NAND U5372 ( .A(n5811), .B(n5143), .Z(n5121) );
  AND U5373 ( .A(n5122), .B(n5121), .Z(n5151) );
  NAND U5374 ( .A(b[0]), .B(a[224]), .Z(n5123) );
  XNOR U5375 ( .A(b[1]), .B(n5123), .Z(n5125) );
  NANDN U5376 ( .A(b[0]), .B(a[223]), .Z(n5124) );
  NAND U5377 ( .A(n5125), .B(n5124), .Z(n5150) );
  AND U5378 ( .A(b[3]), .B(a[220]), .Z(n5149) );
  XOR U5379 ( .A(n5150), .B(n5149), .Z(n5152) );
  XOR U5380 ( .A(n5151), .B(n5152), .Z(n5138) );
  NANDN U5381 ( .A(n5127), .B(n5126), .Z(n5131) );
  OR U5382 ( .A(n5129), .B(n5128), .Z(n5130) );
  AND U5383 ( .A(n5131), .B(n5130), .Z(n5137) );
  XOR U5384 ( .A(n5138), .B(n5137), .Z(n5140) );
  XOR U5385 ( .A(n5139), .B(n5140), .Z(n5155) );
  XNOR U5386 ( .A(n5155), .B(sreg[476]), .Z(n5157) );
  NANDN U5387 ( .A(n5132), .B(sreg[475]), .Z(n5136) );
  NAND U5388 ( .A(n5134), .B(n5133), .Z(n5135) );
  NAND U5389 ( .A(n5136), .B(n5135), .Z(n5156) );
  XOR U5390 ( .A(n5157), .B(n5156), .Z(c[476]) );
  NANDN U5391 ( .A(n5138), .B(n5137), .Z(n5142) );
  OR U5392 ( .A(n5140), .B(n5139), .Z(n5141) );
  AND U5393 ( .A(n5142), .B(n5141), .Z(n5162) );
  NAND U5394 ( .A(n31), .B(n5143), .Z(n5145) );
  XOR U5395 ( .A(b[3]), .B(a[223]), .Z(n5166) );
  NAND U5396 ( .A(n5811), .B(n5166), .Z(n5144) );
  AND U5397 ( .A(n5145), .B(n5144), .Z(n5174) );
  NAND U5398 ( .A(b[0]), .B(a[225]), .Z(n5146) );
  XNOR U5399 ( .A(b[1]), .B(n5146), .Z(n5148) );
  NANDN U5400 ( .A(b[0]), .B(a[224]), .Z(n5147) );
  NAND U5401 ( .A(n5148), .B(n5147), .Z(n5173) );
  AND U5402 ( .A(b[3]), .B(a[221]), .Z(n5172) );
  XOR U5403 ( .A(n5173), .B(n5172), .Z(n5175) );
  XOR U5404 ( .A(n5174), .B(n5175), .Z(n5161) );
  NANDN U5405 ( .A(n5150), .B(n5149), .Z(n5154) );
  OR U5406 ( .A(n5152), .B(n5151), .Z(n5153) );
  AND U5407 ( .A(n5154), .B(n5153), .Z(n5160) );
  XOR U5408 ( .A(n5161), .B(n5160), .Z(n5163) );
  XOR U5409 ( .A(n5162), .B(n5163), .Z(n5178) );
  XNOR U5410 ( .A(n5178), .B(sreg[477]), .Z(n5180) );
  NANDN U5411 ( .A(n5155), .B(sreg[476]), .Z(n5159) );
  NAND U5412 ( .A(n5157), .B(n5156), .Z(n5158) );
  NAND U5413 ( .A(n5159), .B(n5158), .Z(n5179) );
  XOR U5414 ( .A(n5180), .B(n5179), .Z(c[477]) );
  NANDN U5415 ( .A(n5161), .B(n5160), .Z(n5165) );
  OR U5416 ( .A(n5163), .B(n5162), .Z(n5164) );
  AND U5417 ( .A(n5165), .B(n5164), .Z(n5185) );
  NAND U5418 ( .A(n31), .B(n5166), .Z(n5168) );
  XOR U5419 ( .A(b[3]), .B(a[224]), .Z(n5189) );
  NAND U5420 ( .A(n5811), .B(n5189), .Z(n5167) );
  AND U5421 ( .A(n5168), .B(n5167), .Z(n5197) );
  AND U5422 ( .A(b[3]), .B(a[222]), .Z(n5195) );
  NAND U5423 ( .A(b[0]), .B(a[226]), .Z(n5169) );
  XNOR U5424 ( .A(b[1]), .B(n5169), .Z(n5171) );
  NANDN U5425 ( .A(b[0]), .B(a[225]), .Z(n5170) );
  NAND U5426 ( .A(n5171), .B(n5170), .Z(n5196) );
  XOR U5427 ( .A(n5195), .B(n5196), .Z(n5198) );
  XOR U5428 ( .A(n5197), .B(n5198), .Z(n5184) );
  NANDN U5429 ( .A(n5173), .B(n5172), .Z(n5177) );
  OR U5430 ( .A(n5175), .B(n5174), .Z(n5176) );
  AND U5431 ( .A(n5177), .B(n5176), .Z(n5183) );
  XOR U5432 ( .A(n5184), .B(n5183), .Z(n5186) );
  XOR U5433 ( .A(n5185), .B(n5186), .Z(n5201) );
  XNOR U5434 ( .A(n5201), .B(sreg[478]), .Z(n5203) );
  NANDN U5435 ( .A(n5178), .B(sreg[477]), .Z(n5182) );
  NAND U5436 ( .A(n5180), .B(n5179), .Z(n5181) );
  NAND U5437 ( .A(n5182), .B(n5181), .Z(n5202) );
  XOR U5438 ( .A(n5203), .B(n5202), .Z(c[478]) );
  NANDN U5439 ( .A(n5184), .B(n5183), .Z(n5188) );
  OR U5440 ( .A(n5186), .B(n5185), .Z(n5187) );
  AND U5441 ( .A(n5188), .B(n5187), .Z(n5208) );
  NAND U5442 ( .A(n31), .B(n5189), .Z(n5191) );
  XOR U5443 ( .A(b[3]), .B(a[225]), .Z(n5212) );
  NAND U5444 ( .A(n5811), .B(n5212), .Z(n5190) );
  AND U5445 ( .A(n5191), .B(n5190), .Z(n5220) );
  NAND U5446 ( .A(b[0]), .B(a[227]), .Z(n5192) );
  XNOR U5447 ( .A(b[1]), .B(n5192), .Z(n5194) );
  NANDN U5448 ( .A(b[0]), .B(a[226]), .Z(n5193) );
  NAND U5449 ( .A(n5194), .B(n5193), .Z(n5219) );
  AND U5450 ( .A(b[3]), .B(a[223]), .Z(n5218) );
  XOR U5451 ( .A(n5219), .B(n5218), .Z(n5221) );
  XOR U5452 ( .A(n5220), .B(n5221), .Z(n5207) );
  NANDN U5453 ( .A(n5196), .B(n5195), .Z(n5200) );
  OR U5454 ( .A(n5198), .B(n5197), .Z(n5199) );
  AND U5455 ( .A(n5200), .B(n5199), .Z(n5206) );
  XOR U5456 ( .A(n5207), .B(n5206), .Z(n5209) );
  XOR U5457 ( .A(n5208), .B(n5209), .Z(n5224) );
  XNOR U5458 ( .A(n5224), .B(sreg[479]), .Z(n5226) );
  NANDN U5459 ( .A(n5201), .B(sreg[478]), .Z(n5205) );
  NAND U5460 ( .A(n5203), .B(n5202), .Z(n5204) );
  NAND U5461 ( .A(n5205), .B(n5204), .Z(n5225) );
  XOR U5462 ( .A(n5226), .B(n5225), .Z(c[479]) );
  NANDN U5463 ( .A(n5207), .B(n5206), .Z(n5211) );
  OR U5464 ( .A(n5209), .B(n5208), .Z(n5210) );
  AND U5465 ( .A(n5211), .B(n5210), .Z(n5231) );
  NAND U5466 ( .A(n31), .B(n5212), .Z(n5214) );
  XOR U5467 ( .A(b[3]), .B(a[226]), .Z(n5235) );
  NAND U5468 ( .A(n5811), .B(n5235), .Z(n5213) );
  AND U5469 ( .A(n5214), .B(n5213), .Z(n5243) );
  NAND U5470 ( .A(b[0]), .B(a[228]), .Z(n5215) );
  XNOR U5471 ( .A(b[1]), .B(n5215), .Z(n5217) );
  NANDN U5472 ( .A(b[0]), .B(a[227]), .Z(n5216) );
  NAND U5473 ( .A(n5217), .B(n5216), .Z(n5242) );
  AND U5474 ( .A(b[3]), .B(a[224]), .Z(n5241) );
  XOR U5475 ( .A(n5242), .B(n5241), .Z(n5244) );
  XOR U5476 ( .A(n5243), .B(n5244), .Z(n5230) );
  NANDN U5477 ( .A(n5219), .B(n5218), .Z(n5223) );
  OR U5478 ( .A(n5221), .B(n5220), .Z(n5222) );
  AND U5479 ( .A(n5223), .B(n5222), .Z(n5229) );
  XOR U5480 ( .A(n5230), .B(n5229), .Z(n5232) );
  XOR U5481 ( .A(n5231), .B(n5232), .Z(n5247) );
  XNOR U5482 ( .A(n5247), .B(sreg[480]), .Z(n5249) );
  NANDN U5483 ( .A(n5224), .B(sreg[479]), .Z(n5228) );
  NAND U5484 ( .A(n5226), .B(n5225), .Z(n5227) );
  NAND U5485 ( .A(n5228), .B(n5227), .Z(n5248) );
  XOR U5486 ( .A(n5249), .B(n5248), .Z(c[480]) );
  NANDN U5487 ( .A(n5230), .B(n5229), .Z(n5234) );
  OR U5488 ( .A(n5232), .B(n5231), .Z(n5233) );
  AND U5489 ( .A(n5234), .B(n5233), .Z(n5254) );
  NAND U5490 ( .A(n31), .B(n5235), .Z(n5237) );
  XOR U5491 ( .A(b[3]), .B(a[227]), .Z(n5258) );
  NAND U5492 ( .A(n5811), .B(n5258), .Z(n5236) );
  AND U5493 ( .A(n5237), .B(n5236), .Z(n5266) );
  NAND U5494 ( .A(b[0]), .B(a[229]), .Z(n5238) );
  XNOR U5495 ( .A(b[1]), .B(n5238), .Z(n5240) );
  NANDN U5496 ( .A(b[0]), .B(a[228]), .Z(n5239) );
  NAND U5497 ( .A(n5240), .B(n5239), .Z(n5265) );
  AND U5498 ( .A(b[3]), .B(a[225]), .Z(n5264) );
  XOR U5499 ( .A(n5265), .B(n5264), .Z(n5267) );
  XOR U5500 ( .A(n5266), .B(n5267), .Z(n5253) );
  NANDN U5501 ( .A(n5242), .B(n5241), .Z(n5246) );
  OR U5502 ( .A(n5244), .B(n5243), .Z(n5245) );
  AND U5503 ( .A(n5246), .B(n5245), .Z(n5252) );
  XOR U5504 ( .A(n5253), .B(n5252), .Z(n5255) );
  XOR U5505 ( .A(n5254), .B(n5255), .Z(n5270) );
  XNOR U5506 ( .A(n5270), .B(sreg[481]), .Z(n5272) );
  NANDN U5507 ( .A(n5247), .B(sreg[480]), .Z(n5251) );
  NAND U5508 ( .A(n5249), .B(n5248), .Z(n5250) );
  NAND U5509 ( .A(n5251), .B(n5250), .Z(n5271) );
  XOR U5510 ( .A(n5272), .B(n5271), .Z(c[481]) );
  NANDN U5511 ( .A(n5253), .B(n5252), .Z(n5257) );
  OR U5512 ( .A(n5255), .B(n5254), .Z(n5256) );
  AND U5513 ( .A(n5257), .B(n5256), .Z(n5277) );
  NAND U5514 ( .A(n31), .B(n5258), .Z(n5260) );
  XOR U5515 ( .A(b[3]), .B(a[228]), .Z(n5281) );
  NAND U5516 ( .A(n5811), .B(n5281), .Z(n5259) );
  AND U5517 ( .A(n5260), .B(n5259), .Z(n5289) );
  NAND U5518 ( .A(b[0]), .B(a[230]), .Z(n5261) );
  XNOR U5519 ( .A(b[1]), .B(n5261), .Z(n5263) );
  NANDN U5520 ( .A(b[0]), .B(a[229]), .Z(n5262) );
  NAND U5521 ( .A(n5263), .B(n5262), .Z(n5288) );
  AND U5522 ( .A(b[3]), .B(a[226]), .Z(n5287) );
  XOR U5523 ( .A(n5288), .B(n5287), .Z(n5290) );
  XOR U5524 ( .A(n5289), .B(n5290), .Z(n5276) );
  NANDN U5525 ( .A(n5265), .B(n5264), .Z(n5269) );
  OR U5526 ( .A(n5267), .B(n5266), .Z(n5268) );
  AND U5527 ( .A(n5269), .B(n5268), .Z(n5275) );
  XOR U5528 ( .A(n5276), .B(n5275), .Z(n5278) );
  XOR U5529 ( .A(n5277), .B(n5278), .Z(n5293) );
  XNOR U5530 ( .A(n5293), .B(sreg[482]), .Z(n5295) );
  NANDN U5531 ( .A(n5270), .B(sreg[481]), .Z(n5274) );
  NAND U5532 ( .A(n5272), .B(n5271), .Z(n5273) );
  NAND U5533 ( .A(n5274), .B(n5273), .Z(n5294) );
  XOR U5534 ( .A(n5295), .B(n5294), .Z(c[482]) );
  NANDN U5535 ( .A(n5276), .B(n5275), .Z(n5280) );
  OR U5536 ( .A(n5278), .B(n5277), .Z(n5279) );
  AND U5537 ( .A(n5280), .B(n5279), .Z(n5300) );
  NAND U5538 ( .A(n31), .B(n5281), .Z(n5283) );
  XOR U5539 ( .A(b[3]), .B(a[229]), .Z(n5304) );
  NAND U5540 ( .A(n5811), .B(n5304), .Z(n5282) );
  AND U5541 ( .A(n5283), .B(n5282), .Z(n5312) );
  AND U5542 ( .A(b[0]), .B(a[231]), .Z(n5284) );
  XOR U5543 ( .A(b[1]), .B(n5284), .Z(n5286) );
  NANDN U5544 ( .A(b[0]), .B(a[230]), .Z(n5285) );
  AND U5545 ( .A(n5286), .B(n5285), .Z(n5310) );
  NAND U5546 ( .A(b[3]), .B(a[227]), .Z(n5311) );
  XOR U5547 ( .A(n5310), .B(n5311), .Z(n5313) );
  XOR U5548 ( .A(n5312), .B(n5313), .Z(n5299) );
  NANDN U5549 ( .A(n5288), .B(n5287), .Z(n5292) );
  OR U5550 ( .A(n5290), .B(n5289), .Z(n5291) );
  AND U5551 ( .A(n5292), .B(n5291), .Z(n5298) );
  XOR U5552 ( .A(n5299), .B(n5298), .Z(n5301) );
  XOR U5553 ( .A(n5300), .B(n5301), .Z(n5316) );
  XNOR U5554 ( .A(n5316), .B(sreg[483]), .Z(n5318) );
  NANDN U5555 ( .A(n5293), .B(sreg[482]), .Z(n5297) );
  NAND U5556 ( .A(n5295), .B(n5294), .Z(n5296) );
  NAND U5557 ( .A(n5297), .B(n5296), .Z(n5317) );
  XOR U5558 ( .A(n5318), .B(n5317), .Z(c[483]) );
  NANDN U5559 ( .A(n5299), .B(n5298), .Z(n5303) );
  OR U5560 ( .A(n5301), .B(n5300), .Z(n5302) );
  AND U5561 ( .A(n5303), .B(n5302), .Z(n5323) );
  NAND U5562 ( .A(n31), .B(n5304), .Z(n5306) );
  XOR U5563 ( .A(b[3]), .B(a[230]), .Z(n5327) );
  NAND U5564 ( .A(n5811), .B(n5327), .Z(n5305) );
  AND U5565 ( .A(n5306), .B(n5305), .Z(n5335) );
  NAND U5566 ( .A(b[0]), .B(a[232]), .Z(n5307) );
  XNOR U5567 ( .A(b[1]), .B(n5307), .Z(n5309) );
  NANDN U5568 ( .A(b[0]), .B(a[231]), .Z(n5308) );
  NAND U5569 ( .A(n5309), .B(n5308), .Z(n5334) );
  AND U5570 ( .A(b[3]), .B(a[228]), .Z(n5333) );
  XOR U5571 ( .A(n5334), .B(n5333), .Z(n5336) );
  XOR U5572 ( .A(n5335), .B(n5336), .Z(n5322) );
  NANDN U5573 ( .A(n5311), .B(n5310), .Z(n5315) );
  OR U5574 ( .A(n5313), .B(n5312), .Z(n5314) );
  AND U5575 ( .A(n5315), .B(n5314), .Z(n5321) );
  XOR U5576 ( .A(n5322), .B(n5321), .Z(n5324) );
  XOR U5577 ( .A(n5323), .B(n5324), .Z(n5339) );
  XNOR U5578 ( .A(n5339), .B(sreg[484]), .Z(n5341) );
  NANDN U5579 ( .A(n5316), .B(sreg[483]), .Z(n5320) );
  NAND U5580 ( .A(n5318), .B(n5317), .Z(n5319) );
  NAND U5581 ( .A(n5320), .B(n5319), .Z(n5340) );
  XOR U5582 ( .A(n5341), .B(n5340), .Z(c[484]) );
  NANDN U5583 ( .A(n5322), .B(n5321), .Z(n5326) );
  OR U5584 ( .A(n5324), .B(n5323), .Z(n5325) );
  AND U5585 ( .A(n5326), .B(n5325), .Z(n5346) );
  NAND U5586 ( .A(n31), .B(n5327), .Z(n5329) );
  XOR U5587 ( .A(b[3]), .B(a[231]), .Z(n5350) );
  NAND U5588 ( .A(n5811), .B(n5350), .Z(n5328) );
  AND U5589 ( .A(n5329), .B(n5328), .Z(n5358) );
  NAND U5590 ( .A(b[0]), .B(a[233]), .Z(n5330) );
  XNOR U5591 ( .A(b[1]), .B(n5330), .Z(n5332) );
  NANDN U5592 ( .A(b[0]), .B(a[232]), .Z(n5331) );
  NAND U5593 ( .A(n5332), .B(n5331), .Z(n5357) );
  AND U5594 ( .A(b[3]), .B(a[229]), .Z(n5356) );
  XOR U5595 ( .A(n5357), .B(n5356), .Z(n5359) );
  XOR U5596 ( .A(n5358), .B(n5359), .Z(n5345) );
  NANDN U5597 ( .A(n5334), .B(n5333), .Z(n5338) );
  OR U5598 ( .A(n5336), .B(n5335), .Z(n5337) );
  AND U5599 ( .A(n5338), .B(n5337), .Z(n5344) );
  XOR U5600 ( .A(n5345), .B(n5344), .Z(n5347) );
  XOR U5601 ( .A(n5346), .B(n5347), .Z(n5362) );
  XNOR U5602 ( .A(n5362), .B(sreg[485]), .Z(n5364) );
  NANDN U5603 ( .A(n5339), .B(sreg[484]), .Z(n5343) );
  NAND U5604 ( .A(n5341), .B(n5340), .Z(n5342) );
  NAND U5605 ( .A(n5343), .B(n5342), .Z(n5363) );
  XOR U5606 ( .A(n5364), .B(n5363), .Z(c[485]) );
  NANDN U5607 ( .A(n5345), .B(n5344), .Z(n5349) );
  OR U5608 ( .A(n5347), .B(n5346), .Z(n5348) );
  AND U5609 ( .A(n5349), .B(n5348), .Z(n5369) );
  NAND U5610 ( .A(n31), .B(n5350), .Z(n5352) );
  XOR U5611 ( .A(b[3]), .B(a[232]), .Z(n5373) );
  NAND U5612 ( .A(n5811), .B(n5373), .Z(n5351) );
  AND U5613 ( .A(n5352), .B(n5351), .Z(n5381) );
  NAND U5614 ( .A(b[0]), .B(a[234]), .Z(n5353) );
  XNOR U5615 ( .A(b[1]), .B(n5353), .Z(n5355) );
  NANDN U5616 ( .A(b[0]), .B(a[233]), .Z(n5354) );
  NAND U5617 ( .A(n5355), .B(n5354), .Z(n5380) );
  AND U5618 ( .A(b[3]), .B(a[230]), .Z(n5379) );
  XOR U5619 ( .A(n5380), .B(n5379), .Z(n5382) );
  XOR U5620 ( .A(n5381), .B(n5382), .Z(n5368) );
  NANDN U5621 ( .A(n5357), .B(n5356), .Z(n5361) );
  OR U5622 ( .A(n5359), .B(n5358), .Z(n5360) );
  AND U5623 ( .A(n5361), .B(n5360), .Z(n5367) );
  XOR U5624 ( .A(n5368), .B(n5367), .Z(n5370) );
  XOR U5625 ( .A(n5369), .B(n5370), .Z(n5385) );
  XNOR U5626 ( .A(n5385), .B(sreg[486]), .Z(n5387) );
  NANDN U5627 ( .A(n5362), .B(sreg[485]), .Z(n5366) );
  NAND U5628 ( .A(n5364), .B(n5363), .Z(n5365) );
  NAND U5629 ( .A(n5366), .B(n5365), .Z(n5386) );
  XOR U5630 ( .A(n5387), .B(n5386), .Z(c[486]) );
  NANDN U5631 ( .A(n5368), .B(n5367), .Z(n5372) );
  OR U5632 ( .A(n5370), .B(n5369), .Z(n5371) );
  AND U5633 ( .A(n5372), .B(n5371), .Z(n5392) );
  NAND U5634 ( .A(n31), .B(n5373), .Z(n5375) );
  XOR U5635 ( .A(b[3]), .B(a[233]), .Z(n5396) );
  NAND U5636 ( .A(n5811), .B(n5396), .Z(n5374) );
  AND U5637 ( .A(n5375), .B(n5374), .Z(n5404) );
  AND U5638 ( .A(b[3]), .B(a[231]), .Z(n5402) );
  NAND U5639 ( .A(b[0]), .B(a[235]), .Z(n5376) );
  XNOR U5640 ( .A(b[1]), .B(n5376), .Z(n5378) );
  NANDN U5641 ( .A(b[0]), .B(a[234]), .Z(n5377) );
  NAND U5642 ( .A(n5378), .B(n5377), .Z(n5403) );
  XOR U5643 ( .A(n5402), .B(n5403), .Z(n5405) );
  XOR U5644 ( .A(n5404), .B(n5405), .Z(n5391) );
  NANDN U5645 ( .A(n5380), .B(n5379), .Z(n5384) );
  OR U5646 ( .A(n5382), .B(n5381), .Z(n5383) );
  AND U5647 ( .A(n5384), .B(n5383), .Z(n5390) );
  XOR U5648 ( .A(n5391), .B(n5390), .Z(n5393) );
  XOR U5649 ( .A(n5392), .B(n5393), .Z(n5408) );
  XNOR U5650 ( .A(n5408), .B(sreg[487]), .Z(n5410) );
  NANDN U5651 ( .A(n5385), .B(sreg[486]), .Z(n5389) );
  NAND U5652 ( .A(n5387), .B(n5386), .Z(n5388) );
  NAND U5653 ( .A(n5389), .B(n5388), .Z(n5409) );
  XOR U5654 ( .A(n5410), .B(n5409), .Z(c[487]) );
  NANDN U5655 ( .A(n5391), .B(n5390), .Z(n5395) );
  OR U5656 ( .A(n5393), .B(n5392), .Z(n5394) );
  AND U5657 ( .A(n5395), .B(n5394), .Z(n5415) );
  NAND U5658 ( .A(n31), .B(n5396), .Z(n5398) );
  XOR U5659 ( .A(b[3]), .B(a[234]), .Z(n5419) );
  NAND U5660 ( .A(n5811), .B(n5419), .Z(n5397) );
  AND U5661 ( .A(n5398), .B(n5397), .Z(n5427) );
  NAND U5662 ( .A(b[0]), .B(a[236]), .Z(n5399) );
  XNOR U5663 ( .A(b[1]), .B(n5399), .Z(n5401) );
  NANDN U5664 ( .A(b[0]), .B(a[235]), .Z(n5400) );
  NAND U5665 ( .A(n5401), .B(n5400), .Z(n5426) );
  AND U5666 ( .A(b[3]), .B(a[232]), .Z(n5425) );
  XOR U5667 ( .A(n5426), .B(n5425), .Z(n5428) );
  XOR U5668 ( .A(n5427), .B(n5428), .Z(n5414) );
  NANDN U5669 ( .A(n5403), .B(n5402), .Z(n5407) );
  OR U5670 ( .A(n5405), .B(n5404), .Z(n5406) );
  AND U5671 ( .A(n5407), .B(n5406), .Z(n5413) );
  XOR U5672 ( .A(n5414), .B(n5413), .Z(n5416) );
  XOR U5673 ( .A(n5415), .B(n5416), .Z(n5431) );
  XNOR U5674 ( .A(n5431), .B(sreg[488]), .Z(n5433) );
  NANDN U5675 ( .A(n5408), .B(sreg[487]), .Z(n5412) );
  NAND U5676 ( .A(n5410), .B(n5409), .Z(n5411) );
  NAND U5677 ( .A(n5412), .B(n5411), .Z(n5432) );
  XOR U5678 ( .A(n5433), .B(n5432), .Z(c[488]) );
  NANDN U5679 ( .A(n5414), .B(n5413), .Z(n5418) );
  OR U5680 ( .A(n5416), .B(n5415), .Z(n5417) );
  AND U5681 ( .A(n5418), .B(n5417), .Z(n5438) );
  NAND U5682 ( .A(n31), .B(n5419), .Z(n5421) );
  XOR U5683 ( .A(b[3]), .B(a[235]), .Z(n5442) );
  NAND U5684 ( .A(n5811), .B(n5442), .Z(n5420) );
  AND U5685 ( .A(n5421), .B(n5420), .Z(n5450) );
  NAND U5686 ( .A(b[0]), .B(a[237]), .Z(n5422) );
  XNOR U5687 ( .A(b[1]), .B(n5422), .Z(n5424) );
  NANDN U5688 ( .A(b[0]), .B(a[236]), .Z(n5423) );
  NAND U5689 ( .A(n5424), .B(n5423), .Z(n5449) );
  AND U5690 ( .A(b[3]), .B(a[233]), .Z(n5448) );
  XOR U5691 ( .A(n5449), .B(n5448), .Z(n5451) );
  XOR U5692 ( .A(n5450), .B(n5451), .Z(n5437) );
  NANDN U5693 ( .A(n5426), .B(n5425), .Z(n5430) );
  OR U5694 ( .A(n5428), .B(n5427), .Z(n5429) );
  AND U5695 ( .A(n5430), .B(n5429), .Z(n5436) );
  XOR U5696 ( .A(n5437), .B(n5436), .Z(n5439) );
  XOR U5697 ( .A(n5438), .B(n5439), .Z(n5454) );
  XNOR U5698 ( .A(n5454), .B(sreg[489]), .Z(n5456) );
  NANDN U5699 ( .A(n5431), .B(sreg[488]), .Z(n5435) );
  NAND U5700 ( .A(n5433), .B(n5432), .Z(n5434) );
  NAND U5701 ( .A(n5435), .B(n5434), .Z(n5455) );
  XOR U5702 ( .A(n5456), .B(n5455), .Z(c[489]) );
  NANDN U5703 ( .A(n5437), .B(n5436), .Z(n5441) );
  OR U5704 ( .A(n5439), .B(n5438), .Z(n5440) );
  AND U5705 ( .A(n5441), .B(n5440), .Z(n5461) );
  NAND U5706 ( .A(n31), .B(n5442), .Z(n5444) );
  XOR U5707 ( .A(b[3]), .B(a[236]), .Z(n5465) );
  NAND U5708 ( .A(n5811), .B(n5465), .Z(n5443) );
  AND U5709 ( .A(n5444), .B(n5443), .Z(n5473) );
  NAND U5710 ( .A(b[0]), .B(a[238]), .Z(n5445) );
  XNOR U5711 ( .A(b[1]), .B(n5445), .Z(n5447) );
  NANDN U5712 ( .A(b[0]), .B(a[237]), .Z(n5446) );
  NAND U5713 ( .A(n5447), .B(n5446), .Z(n5472) );
  AND U5714 ( .A(b[3]), .B(a[234]), .Z(n5471) );
  XOR U5715 ( .A(n5472), .B(n5471), .Z(n5474) );
  XOR U5716 ( .A(n5473), .B(n5474), .Z(n5460) );
  NANDN U5717 ( .A(n5449), .B(n5448), .Z(n5453) );
  OR U5718 ( .A(n5451), .B(n5450), .Z(n5452) );
  AND U5719 ( .A(n5453), .B(n5452), .Z(n5459) );
  XOR U5720 ( .A(n5460), .B(n5459), .Z(n5462) );
  XOR U5721 ( .A(n5461), .B(n5462), .Z(n5477) );
  XNOR U5722 ( .A(n5477), .B(sreg[490]), .Z(n5479) );
  NANDN U5723 ( .A(n5454), .B(sreg[489]), .Z(n5458) );
  NAND U5724 ( .A(n5456), .B(n5455), .Z(n5457) );
  NAND U5725 ( .A(n5458), .B(n5457), .Z(n5478) );
  XOR U5726 ( .A(n5479), .B(n5478), .Z(c[490]) );
  NANDN U5727 ( .A(n5460), .B(n5459), .Z(n5464) );
  OR U5728 ( .A(n5462), .B(n5461), .Z(n5463) );
  AND U5729 ( .A(n5464), .B(n5463), .Z(n5484) );
  NAND U5730 ( .A(n31), .B(n5465), .Z(n5467) );
  XOR U5731 ( .A(b[3]), .B(a[237]), .Z(n5488) );
  NAND U5732 ( .A(n5811), .B(n5488), .Z(n5466) );
  AND U5733 ( .A(n5467), .B(n5466), .Z(n5496) );
  AND U5734 ( .A(b[3]), .B(a[235]), .Z(n5494) );
  NAND U5735 ( .A(b[0]), .B(a[239]), .Z(n5468) );
  XNOR U5736 ( .A(b[1]), .B(n5468), .Z(n5470) );
  NANDN U5737 ( .A(b[0]), .B(a[238]), .Z(n5469) );
  NAND U5738 ( .A(n5470), .B(n5469), .Z(n5495) );
  XOR U5739 ( .A(n5494), .B(n5495), .Z(n5497) );
  XOR U5740 ( .A(n5496), .B(n5497), .Z(n5483) );
  NANDN U5741 ( .A(n5472), .B(n5471), .Z(n5476) );
  OR U5742 ( .A(n5474), .B(n5473), .Z(n5475) );
  AND U5743 ( .A(n5476), .B(n5475), .Z(n5482) );
  XOR U5744 ( .A(n5483), .B(n5482), .Z(n5485) );
  XOR U5745 ( .A(n5484), .B(n5485), .Z(n5500) );
  XNOR U5746 ( .A(n5500), .B(sreg[491]), .Z(n5502) );
  NANDN U5747 ( .A(n5477), .B(sreg[490]), .Z(n5481) );
  NAND U5748 ( .A(n5479), .B(n5478), .Z(n5480) );
  NAND U5749 ( .A(n5481), .B(n5480), .Z(n5501) );
  XOR U5750 ( .A(n5502), .B(n5501), .Z(c[491]) );
  NANDN U5751 ( .A(n5483), .B(n5482), .Z(n5487) );
  OR U5752 ( .A(n5485), .B(n5484), .Z(n5486) );
  AND U5753 ( .A(n5487), .B(n5486), .Z(n5507) );
  NAND U5754 ( .A(n31), .B(n5488), .Z(n5490) );
  XOR U5755 ( .A(b[3]), .B(a[238]), .Z(n5511) );
  NAND U5756 ( .A(n5811), .B(n5511), .Z(n5489) );
  AND U5757 ( .A(n5490), .B(n5489), .Z(n5519) );
  NAND U5758 ( .A(b[0]), .B(a[240]), .Z(n5491) );
  XNOR U5759 ( .A(b[1]), .B(n5491), .Z(n5493) );
  NANDN U5760 ( .A(b[0]), .B(a[239]), .Z(n5492) );
  NAND U5761 ( .A(n5493), .B(n5492), .Z(n5518) );
  AND U5762 ( .A(b[3]), .B(a[236]), .Z(n5517) );
  XOR U5763 ( .A(n5518), .B(n5517), .Z(n5520) );
  XOR U5764 ( .A(n5519), .B(n5520), .Z(n5506) );
  NANDN U5765 ( .A(n5495), .B(n5494), .Z(n5499) );
  OR U5766 ( .A(n5497), .B(n5496), .Z(n5498) );
  AND U5767 ( .A(n5499), .B(n5498), .Z(n5505) );
  XOR U5768 ( .A(n5506), .B(n5505), .Z(n5508) );
  XOR U5769 ( .A(n5507), .B(n5508), .Z(n5523) );
  XNOR U5770 ( .A(n5523), .B(sreg[492]), .Z(n5525) );
  NANDN U5771 ( .A(n5500), .B(sreg[491]), .Z(n5504) );
  NAND U5772 ( .A(n5502), .B(n5501), .Z(n5503) );
  NAND U5773 ( .A(n5504), .B(n5503), .Z(n5524) );
  XOR U5774 ( .A(n5525), .B(n5524), .Z(c[492]) );
  NANDN U5775 ( .A(n5506), .B(n5505), .Z(n5510) );
  OR U5776 ( .A(n5508), .B(n5507), .Z(n5509) );
  AND U5777 ( .A(n5510), .B(n5509), .Z(n5530) );
  NAND U5778 ( .A(n31), .B(n5511), .Z(n5513) );
  XOR U5779 ( .A(b[3]), .B(a[239]), .Z(n5534) );
  NAND U5780 ( .A(n5811), .B(n5534), .Z(n5512) );
  AND U5781 ( .A(n5513), .B(n5512), .Z(n5542) );
  NAND U5782 ( .A(b[0]), .B(a[241]), .Z(n5514) );
  XNOR U5783 ( .A(b[1]), .B(n5514), .Z(n5516) );
  NANDN U5784 ( .A(b[0]), .B(a[240]), .Z(n5515) );
  NAND U5785 ( .A(n5516), .B(n5515), .Z(n5541) );
  AND U5786 ( .A(b[3]), .B(a[237]), .Z(n5540) );
  XOR U5787 ( .A(n5541), .B(n5540), .Z(n5543) );
  XOR U5788 ( .A(n5542), .B(n5543), .Z(n5529) );
  NANDN U5789 ( .A(n5518), .B(n5517), .Z(n5522) );
  OR U5790 ( .A(n5520), .B(n5519), .Z(n5521) );
  AND U5791 ( .A(n5522), .B(n5521), .Z(n5528) );
  XOR U5792 ( .A(n5529), .B(n5528), .Z(n5531) );
  XOR U5793 ( .A(n5530), .B(n5531), .Z(n5546) );
  XNOR U5794 ( .A(n5546), .B(sreg[493]), .Z(n5548) );
  NANDN U5795 ( .A(n5523), .B(sreg[492]), .Z(n5527) );
  NAND U5796 ( .A(n5525), .B(n5524), .Z(n5526) );
  NAND U5797 ( .A(n5527), .B(n5526), .Z(n5547) );
  XOR U5798 ( .A(n5548), .B(n5547), .Z(c[493]) );
  NANDN U5799 ( .A(n5529), .B(n5528), .Z(n5533) );
  OR U5800 ( .A(n5531), .B(n5530), .Z(n5532) );
  AND U5801 ( .A(n5533), .B(n5532), .Z(n5553) );
  NAND U5802 ( .A(n31), .B(n5534), .Z(n5536) );
  XOR U5803 ( .A(b[3]), .B(a[240]), .Z(n5557) );
  NAND U5804 ( .A(n5811), .B(n5557), .Z(n5535) );
  AND U5805 ( .A(n5536), .B(n5535), .Z(n5565) );
  NAND U5806 ( .A(b[0]), .B(a[242]), .Z(n5537) );
  XNOR U5807 ( .A(b[1]), .B(n5537), .Z(n5539) );
  NANDN U5808 ( .A(b[0]), .B(a[241]), .Z(n5538) );
  NAND U5809 ( .A(n5539), .B(n5538), .Z(n5564) );
  AND U5810 ( .A(b[3]), .B(a[238]), .Z(n5563) );
  XOR U5811 ( .A(n5564), .B(n5563), .Z(n5566) );
  XOR U5812 ( .A(n5565), .B(n5566), .Z(n5552) );
  NANDN U5813 ( .A(n5541), .B(n5540), .Z(n5545) );
  OR U5814 ( .A(n5543), .B(n5542), .Z(n5544) );
  AND U5815 ( .A(n5545), .B(n5544), .Z(n5551) );
  XOR U5816 ( .A(n5552), .B(n5551), .Z(n5554) );
  XOR U5817 ( .A(n5553), .B(n5554), .Z(n5569) );
  XNOR U5818 ( .A(n5569), .B(sreg[494]), .Z(n5571) );
  NANDN U5819 ( .A(n5546), .B(sreg[493]), .Z(n5550) );
  NAND U5820 ( .A(n5548), .B(n5547), .Z(n5549) );
  NAND U5821 ( .A(n5550), .B(n5549), .Z(n5570) );
  XOR U5822 ( .A(n5571), .B(n5570), .Z(c[494]) );
  NANDN U5823 ( .A(n5552), .B(n5551), .Z(n5556) );
  OR U5824 ( .A(n5554), .B(n5553), .Z(n5555) );
  AND U5825 ( .A(n5556), .B(n5555), .Z(n5576) );
  NAND U5826 ( .A(n31), .B(n5557), .Z(n5559) );
  XOR U5827 ( .A(b[3]), .B(a[241]), .Z(n5580) );
  NAND U5828 ( .A(n5811), .B(n5580), .Z(n5558) );
  AND U5829 ( .A(n5559), .B(n5558), .Z(n5588) );
  NAND U5830 ( .A(b[0]), .B(a[243]), .Z(n5560) );
  XNOR U5831 ( .A(b[1]), .B(n5560), .Z(n5562) );
  NANDN U5832 ( .A(b[0]), .B(a[242]), .Z(n5561) );
  NAND U5833 ( .A(n5562), .B(n5561), .Z(n5587) );
  AND U5834 ( .A(b[3]), .B(a[239]), .Z(n5586) );
  XOR U5835 ( .A(n5587), .B(n5586), .Z(n5589) );
  XOR U5836 ( .A(n5588), .B(n5589), .Z(n5575) );
  NANDN U5837 ( .A(n5564), .B(n5563), .Z(n5568) );
  OR U5838 ( .A(n5566), .B(n5565), .Z(n5567) );
  AND U5839 ( .A(n5568), .B(n5567), .Z(n5574) );
  XOR U5840 ( .A(n5575), .B(n5574), .Z(n5577) );
  XOR U5841 ( .A(n5576), .B(n5577), .Z(n5592) );
  XNOR U5842 ( .A(n5592), .B(sreg[495]), .Z(n5594) );
  NANDN U5843 ( .A(n5569), .B(sreg[494]), .Z(n5573) );
  NAND U5844 ( .A(n5571), .B(n5570), .Z(n5572) );
  NAND U5845 ( .A(n5573), .B(n5572), .Z(n5593) );
  XOR U5846 ( .A(n5594), .B(n5593), .Z(c[495]) );
  NANDN U5847 ( .A(n5575), .B(n5574), .Z(n5579) );
  OR U5848 ( .A(n5577), .B(n5576), .Z(n5578) );
  AND U5849 ( .A(n5579), .B(n5578), .Z(n5599) );
  NAND U5850 ( .A(n31), .B(n5580), .Z(n5582) );
  XOR U5851 ( .A(b[3]), .B(a[242]), .Z(n5603) );
  NAND U5852 ( .A(n5811), .B(n5603), .Z(n5581) );
  AND U5853 ( .A(n5582), .B(n5581), .Z(n5611) );
  NAND U5854 ( .A(b[0]), .B(a[244]), .Z(n5583) );
  XNOR U5855 ( .A(b[1]), .B(n5583), .Z(n5585) );
  NANDN U5856 ( .A(b[0]), .B(a[243]), .Z(n5584) );
  NAND U5857 ( .A(n5585), .B(n5584), .Z(n5610) );
  AND U5858 ( .A(b[3]), .B(a[240]), .Z(n5609) );
  XOR U5859 ( .A(n5610), .B(n5609), .Z(n5612) );
  XOR U5860 ( .A(n5611), .B(n5612), .Z(n5598) );
  NANDN U5861 ( .A(n5587), .B(n5586), .Z(n5591) );
  OR U5862 ( .A(n5589), .B(n5588), .Z(n5590) );
  AND U5863 ( .A(n5591), .B(n5590), .Z(n5597) );
  XOR U5864 ( .A(n5598), .B(n5597), .Z(n5600) );
  XOR U5865 ( .A(n5599), .B(n5600), .Z(n5615) );
  XNOR U5866 ( .A(n5615), .B(sreg[496]), .Z(n5617) );
  NANDN U5867 ( .A(n5592), .B(sreg[495]), .Z(n5596) );
  NAND U5868 ( .A(n5594), .B(n5593), .Z(n5595) );
  NAND U5869 ( .A(n5596), .B(n5595), .Z(n5616) );
  XOR U5870 ( .A(n5617), .B(n5616), .Z(c[496]) );
  NANDN U5871 ( .A(n5598), .B(n5597), .Z(n5602) );
  OR U5872 ( .A(n5600), .B(n5599), .Z(n5601) );
  AND U5873 ( .A(n5602), .B(n5601), .Z(n5622) );
  NAND U5874 ( .A(n31), .B(n5603), .Z(n5605) );
  XOR U5875 ( .A(b[3]), .B(a[243]), .Z(n5626) );
  NAND U5876 ( .A(n5811), .B(n5626), .Z(n5604) );
  AND U5877 ( .A(n5605), .B(n5604), .Z(n5634) );
  AND U5878 ( .A(b[3]), .B(a[241]), .Z(n5632) );
  NAND U5879 ( .A(b[0]), .B(a[245]), .Z(n5606) );
  XNOR U5880 ( .A(b[1]), .B(n5606), .Z(n5608) );
  NANDN U5881 ( .A(b[0]), .B(a[244]), .Z(n5607) );
  NAND U5882 ( .A(n5608), .B(n5607), .Z(n5633) );
  XOR U5883 ( .A(n5632), .B(n5633), .Z(n5635) );
  XOR U5884 ( .A(n5634), .B(n5635), .Z(n5621) );
  NANDN U5885 ( .A(n5610), .B(n5609), .Z(n5614) );
  OR U5886 ( .A(n5612), .B(n5611), .Z(n5613) );
  AND U5887 ( .A(n5614), .B(n5613), .Z(n5620) );
  XOR U5888 ( .A(n5621), .B(n5620), .Z(n5623) );
  XOR U5889 ( .A(n5622), .B(n5623), .Z(n5638) );
  XNOR U5890 ( .A(n5638), .B(sreg[497]), .Z(n5640) );
  NANDN U5891 ( .A(n5615), .B(sreg[496]), .Z(n5619) );
  NAND U5892 ( .A(n5617), .B(n5616), .Z(n5618) );
  NAND U5893 ( .A(n5619), .B(n5618), .Z(n5639) );
  XOR U5894 ( .A(n5640), .B(n5639), .Z(c[497]) );
  NANDN U5895 ( .A(n5621), .B(n5620), .Z(n5625) );
  OR U5896 ( .A(n5623), .B(n5622), .Z(n5624) );
  AND U5897 ( .A(n5625), .B(n5624), .Z(n5645) );
  NAND U5898 ( .A(n31), .B(n5626), .Z(n5628) );
  XOR U5899 ( .A(b[3]), .B(a[244]), .Z(n5649) );
  NAND U5900 ( .A(n5811), .B(n5649), .Z(n5627) );
  AND U5901 ( .A(n5628), .B(n5627), .Z(n5657) );
  NAND U5902 ( .A(b[0]), .B(a[246]), .Z(n5629) );
  XNOR U5903 ( .A(b[1]), .B(n5629), .Z(n5631) );
  NANDN U5904 ( .A(b[0]), .B(a[245]), .Z(n5630) );
  NAND U5905 ( .A(n5631), .B(n5630), .Z(n5656) );
  AND U5906 ( .A(b[3]), .B(a[242]), .Z(n5655) );
  XOR U5907 ( .A(n5656), .B(n5655), .Z(n5658) );
  XOR U5908 ( .A(n5657), .B(n5658), .Z(n5644) );
  NANDN U5909 ( .A(n5633), .B(n5632), .Z(n5637) );
  OR U5910 ( .A(n5635), .B(n5634), .Z(n5636) );
  AND U5911 ( .A(n5637), .B(n5636), .Z(n5643) );
  XOR U5912 ( .A(n5644), .B(n5643), .Z(n5646) );
  XOR U5913 ( .A(n5645), .B(n5646), .Z(n5661) );
  XNOR U5914 ( .A(n5661), .B(sreg[498]), .Z(n5663) );
  NANDN U5915 ( .A(n5638), .B(sreg[497]), .Z(n5642) );
  NAND U5916 ( .A(n5640), .B(n5639), .Z(n5641) );
  NAND U5917 ( .A(n5642), .B(n5641), .Z(n5662) );
  XOR U5918 ( .A(n5663), .B(n5662), .Z(c[498]) );
  NANDN U5919 ( .A(n5644), .B(n5643), .Z(n5648) );
  OR U5920 ( .A(n5646), .B(n5645), .Z(n5647) );
  AND U5921 ( .A(n5648), .B(n5647), .Z(n5668) );
  NAND U5922 ( .A(n31), .B(n5649), .Z(n5651) );
  XOR U5923 ( .A(b[3]), .B(a[245]), .Z(n5672) );
  NAND U5924 ( .A(n5811), .B(n5672), .Z(n5650) );
  AND U5925 ( .A(n5651), .B(n5650), .Z(n5680) );
  AND U5926 ( .A(b[3]), .B(a[243]), .Z(n5678) );
  NAND U5927 ( .A(b[0]), .B(a[247]), .Z(n5652) );
  XNOR U5928 ( .A(b[1]), .B(n5652), .Z(n5654) );
  NANDN U5929 ( .A(b[0]), .B(a[246]), .Z(n5653) );
  NAND U5930 ( .A(n5654), .B(n5653), .Z(n5679) );
  XOR U5931 ( .A(n5678), .B(n5679), .Z(n5681) );
  XOR U5932 ( .A(n5680), .B(n5681), .Z(n5667) );
  NANDN U5933 ( .A(n5656), .B(n5655), .Z(n5660) );
  OR U5934 ( .A(n5658), .B(n5657), .Z(n5659) );
  AND U5935 ( .A(n5660), .B(n5659), .Z(n5666) );
  XOR U5936 ( .A(n5667), .B(n5666), .Z(n5669) );
  XOR U5937 ( .A(n5668), .B(n5669), .Z(n5684) );
  XNOR U5938 ( .A(n5684), .B(sreg[499]), .Z(n5686) );
  NANDN U5939 ( .A(n5661), .B(sreg[498]), .Z(n5665) );
  NAND U5940 ( .A(n5663), .B(n5662), .Z(n5664) );
  NAND U5941 ( .A(n5665), .B(n5664), .Z(n5685) );
  XOR U5942 ( .A(n5686), .B(n5685), .Z(c[499]) );
  NANDN U5943 ( .A(n5667), .B(n5666), .Z(n5671) );
  OR U5944 ( .A(n5669), .B(n5668), .Z(n5670) );
  AND U5945 ( .A(n5671), .B(n5670), .Z(n5691) );
  NAND U5946 ( .A(n31), .B(n5672), .Z(n5674) );
  XOR U5947 ( .A(b[3]), .B(a[246]), .Z(n5695) );
  NAND U5948 ( .A(n5811), .B(n5695), .Z(n5673) );
  AND U5949 ( .A(n5674), .B(n5673), .Z(n5703) );
  NAND U5950 ( .A(b[0]), .B(a[248]), .Z(n5675) );
  XNOR U5951 ( .A(b[1]), .B(n5675), .Z(n5677) );
  NANDN U5952 ( .A(b[0]), .B(a[247]), .Z(n5676) );
  NAND U5953 ( .A(n5677), .B(n5676), .Z(n5702) );
  AND U5954 ( .A(b[3]), .B(a[244]), .Z(n5701) );
  XOR U5955 ( .A(n5702), .B(n5701), .Z(n5704) );
  XOR U5956 ( .A(n5703), .B(n5704), .Z(n5690) );
  NANDN U5957 ( .A(n5679), .B(n5678), .Z(n5683) );
  OR U5958 ( .A(n5681), .B(n5680), .Z(n5682) );
  AND U5959 ( .A(n5683), .B(n5682), .Z(n5689) );
  XOR U5960 ( .A(n5690), .B(n5689), .Z(n5692) );
  XOR U5961 ( .A(n5691), .B(n5692), .Z(n5707) );
  XNOR U5962 ( .A(n5707), .B(sreg[500]), .Z(n5709) );
  NANDN U5963 ( .A(n5684), .B(sreg[499]), .Z(n5688) );
  NAND U5964 ( .A(n5686), .B(n5685), .Z(n5687) );
  NAND U5965 ( .A(n5688), .B(n5687), .Z(n5708) );
  XOR U5966 ( .A(n5709), .B(n5708), .Z(c[500]) );
  NANDN U5967 ( .A(n5690), .B(n5689), .Z(n5694) );
  OR U5968 ( .A(n5692), .B(n5691), .Z(n5693) );
  AND U5969 ( .A(n5694), .B(n5693), .Z(n5714) );
  NAND U5970 ( .A(n31), .B(n5695), .Z(n5697) );
  XOR U5971 ( .A(b[3]), .B(a[247]), .Z(n5718) );
  NAND U5972 ( .A(n5811), .B(n5718), .Z(n5696) );
  AND U5973 ( .A(n5697), .B(n5696), .Z(n5726) );
  NAND U5974 ( .A(b[0]), .B(a[249]), .Z(n5698) );
  XNOR U5975 ( .A(b[1]), .B(n5698), .Z(n5700) );
  NANDN U5976 ( .A(b[0]), .B(a[248]), .Z(n5699) );
  NAND U5977 ( .A(n5700), .B(n5699), .Z(n5725) );
  AND U5978 ( .A(b[3]), .B(a[245]), .Z(n5724) );
  XOR U5979 ( .A(n5725), .B(n5724), .Z(n5727) );
  XOR U5980 ( .A(n5726), .B(n5727), .Z(n5713) );
  NANDN U5981 ( .A(n5702), .B(n5701), .Z(n5706) );
  OR U5982 ( .A(n5704), .B(n5703), .Z(n5705) );
  AND U5983 ( .A(n5706), .B(n5705), .Z(n5712) );
  XOR U5984 ( .A(n5713), .B(n5712), .Z(n5715) );
  XOR U5985 ( .A(n5714), .B(n5715), .Z(n5730) );
  XNOR U5986 ( .A(n5730), .B(sreg[501]), .Z(n5732) );
  NANDN U5987 ( .A(n5707), .B(sreg[500]), .Z(n5711) );
  NAND U5988 ( .A(n5709), .B(n5708), .Z(n5710) );
  NAND U5989 ( .A(n5711), .B(n5710), .Z(n5731) );
  XOR U5990 ( .A(n5732), .B(n5731), .Z(c[501]) );
  NANDN U5991 ( .A(n5713), .B(n5712), .Z(n5717) );
  OR U5992 ( .A(n5715), .B(n5714), .Z(n5716) );
  AND U5993 ( .A(n5717), .B(n5716), .Z(n5737) );
  NAND U5994 ( .A(n31), .B(n5718), .Z(n5720) );
  XOR U5995 ( .A(b[3]), .B(a[248]), .Z(n5741) );
  NAND U5996 ( .A(n5811), .B(n5741), .Z(n5719) );
  AND U5997 ( .A(n5720), .B(n5719), .Z(n5749) );
  NAND U5998 ( .A(b[0]), .B(a[250]), .Z(n5721) );
  XNOR U5999 ( .A(b[1]), .B(n5721), .Z(n5723) );
  NANDN U6000 ( .A(b[0]), .B(a[249]), .Z(n5722) );
  NAND U6001 ( .A(n5723), .B(n5722), .Z(n5748) );
  AND U6002 ( .A(b[3]), .B(a[246]), .Z(n5747) );
  XOR U6003 ( .A(n5748), .B(n5747), .Z(n5750) );
  XOR U6004 ( .A(n5749), .B(n5750), .Z(n5736) );
  NANDN U6005 ( .A(n5725), .B(n5724), .Z(n5729) );
  OR U6006 ( .A(n5727), .B(n5726), .Z(n5728) );
  AND U6007 ( .A(n5729), .B(n5728), .Z(n5735) );
  XOR U6008 ( .A(n5736), .B(n5735), .Z(n5738) );
  XOR U6009 ( .A(n5737), .B(n5738), .Z(n5753) );
  XNOR U6010 ( .A(n5753), .B(sreg[502]), .Z(n5755) );
  NANDN U6011 ( .A(n5730), .B(sreg[501]), .Z(n5734) );
  NAND U6012 ( .A(n5732), .B(n5731), .Z(n5733) );
  NAND U6013 ( .A(n5734), .B(n5733), .Z(n5754) );
  XOR U6014 ( .A(n5755), .B(n5754), .Z(c[502]) );
  NANDN U6015 ( .A(n5736), .B(n5735), .Z(n5740) );
  OR U6016 ( .A(n5738), .B(n5737), .Z(n5739) );
  AND U6017 ( .A(n5740), .B(n5739), .Z(n5760) );
  NAND U6018 ( .A(n31), .B(n5741), .Z(n5743) );
  XOR U6019 ( .A(b[3]), .B(a[249]), .Z(n5764) );
  NAND U6020 ( .A(n5811), .B(n5764), .Z(n5742) );
  AND U6021 ( .A(n5743), .B(n5742), .Z(n5772) );
  NAND U6022 ( .A(b[0]), .B(a[251]), .Z(n5744) );
  XNOR U6023 ( .A(b[1]), .B(n5744), .Z(n5746) );
  NANDN U6024 ( .A(b[0]), .B(a[250]), .Z(n5745) );
  NAND U6025 ( .A(n5746), .B(n5745), .Z(n5771) );
  AND U6026 ( .A(b[3]), .B(a[247]), .Z(n5770) );
  XOR U6027 ( .A(n5771), .B(n5770), .Z(n5773) );
  XOR U6028 ( .A(n5772), .B(n5773), .Z(n5759) );
  NANDN U6029 ( .A(n5748), .B(n5747), .Z(n5752) );
  OR U6030 ( .A(n5750), .B(n5749), .Z(n5751) );
  AND U6031 ( .A(n5752), .B(n5751), .Z(n5758) );
  XOR U6032 ( .A(n5759), .B(n5758), .Z(n5761) );
  XOR U6033 ( .A(n5760), .B(n5761), .Z(n5776) );
  XNOR U6034 ( .A(n5776), .B(sreg[503]), .Z(n5778) );
  NANDN U6035 ( .A(n5753), .B(sreg[502]), .Z(n5757) );
  NAND U6036 ( .A(n5755), .B(n5754), .Z(n5756) );
  NAND U6037 ( .A(n5757), .B(n5756), .Z(n5777) );
  XOR U6038 ( .A(n5778), .B(n5777), .Z(c[503]) );
  NANDN U6039 ( .A(n5759), .B(n5758), .Z(n5763) );
  OR U6040 ( .A(n5761), .B(n5760), .Z(n5762) );
  AND U6041 ( .A(n5763), .B(n5762), .Z(n5783) );
  NAND U6042 ( .A(n31), .B(n5764), .Z(n5766) );
  XOR U6043 ( .A(b[3]), .B(a[250]), .Z(n5787) );
  NAND U6044 ( .A(n5811), .B(n5787), .Z(n5765) );
  AND U6045 ( .A(n5766), .B(n5765), .Z(n5795) );
  AND U6046 ( .A(b[3]), .B(a[248]), .Z(n5793) );
  NAND U6047 ( .A(b[0]), .B(a[252]), .Z(n5767) );
  XNOR U6048 ( .A(b[1]), .B(n5767), .Z(n5769) );
  NANDN U6049 ( .A(b[0]), .B(a[251]), .Z(n5768) );
  NAND U6050 ( .A(n5769), .B(n5768), .Z(n5794) );
  XOR U6051 ( .A(n5793), .B(n5794), .Z(n5796) );
  XOR U6052 ( .A(n5795), .B(n5796), .Z(n5782) );
  NANDN U6053 ( .A(n5771), .B(n5770), .Z(n5775) );
  OR U6054 ( .A(n5773), .B(n5772), .Z(n5774) );
  AND U6055 ( .A(n5775), .B(n5774), .Z(n5781) );
  XOR U6056 ( .A(n5782), .B(n5781), .Z(n5784) );
  XOR U6057 ( .A(n5783), .B(n5784), .Z(n5799) );
  XNOR U6058 ( .A(n5799), .B(sreg[504]), .Z(n5801) );
  NANDN U6059 ( .A(n5776), .B(sreg[503]), .Z(n5780) );
  NAND U6060 ( .A(n5778), .B(n5777), .Z(n5779) );
  NAND U6061 ( .A(n5780), .B(n5779), .Z(n5800) );
  XOR U6062 ( .A(n5801), .B(n5800), .Z(c[504]) );
  NANDN U6063 ( .A(n5782), .B(n5781), .Z(n5786) );
  OR U6064 ( .A(n5784), .B(n5783), .Z(n5785) );
  AND U6065 ( .A(n5786), .B(n5785), .Z(n5806) );
  NAND U6066 ( .A(n31), .B(n5787), .Z(n5789) );
  XOR U6067 ( .A(b[3]), .B(a[251]), .Z(n5810) );
  NAND U6068 ( .A(n5811), .B(n5810), .Z(n5788) );
  AND U6069 ( .A(n5789), .B(n5788), .Z(n5819) );
  NAND U6070 ( .A(b[0]), .B(a[253]), .Z(n5790) );
  XNOR U6071 ( .A(b[1]), .B(n5790), .Z(n5792) );
  NANDN U6072 ( .A(b[0]), .B(a[252]), .Z(n5791) );
  NAND U6073 ( .A(n5792), .B(n5791), .Z(n5818) );
  AND U6074 ( .A(b[3]), .B(a[249]), .Z(n5817) );
  XOR U6075 ( .A(n5818), .B(n5817), .Z(n5820) );
  XOR U6076 ( .A(n5819), .B(n5820), .Z(n5805) );
  NANDN U6077 ( .A(n5794), .B(n5793), .Z(n5798) );
  OR U6078 ( .A(n5796), .B(n5795), .Z(n5797) );
  AND U6079 ( .A(n5798), .B(n5797), .Z(n5804) );
  XOR U6080 ( .A(n5805), .B(n5804), .Z(n5807) );
  XOR U6081 ( .A(n5806), .B(n5807), .Z(n5823) );
  XNOR U6082 ( .A(n5823), .B(sreg[505]), .Z(n5825) );
  NANDN U6083 ( .A(n5799), .B(sreg[504]), .Z(n5803) );
  NAND U6084 ( .A(n5801), .B(n5800), .Z(n5802) );
  NAND U6085 ( .A(n5803), .B(n5802), .Z(n5824) );
  XOR U6086 ( .A(n5825), .B(n5824), .Z(c[505]) );
  NANDN U6087 ( .A(n5805), .B(n5804), .Z(n5809) );
  OR U6088 ( .A(n5807), .B(n5806), .Z(n5808) );
  AND U6089 ( .A(n5809), .B(n5808), .Z(n5830) );
  NAND U6090 ( .A(n31), .B(n5810), .Z(n5813) );
  XOR U6091 ( .A(b[3]), .B(a[252]), .Z(n5834) );
  NAND U6092 ( .A(n5811), .B(n5834), .Z(n5812) );
  AND U6093 ( .A(n5813), .B(n5812), .Z(n5842) );
  NAND U6094 ( .A(b[0]), .B(a[254]), .Z(n5814) );
  XNOR U6095 ( .A(b[1]), .B(n5814), .Z(n5816) );
  NANDN U6096 ( .A(b[0]), .B(a[253]), .Z(n5815) );
  NAND U6097 ( .A(n5816), .B(n5815), .Z(n5841) );
  AND U6098 ( .A(b[3]), .B(a[250]), .Z(n5840) );
  XOR U6099 ( .A(n5841), .B(n5840), .Z(n5843) );
  XOR U6100 ( .A(n5842), .B(n5843), .Z(n5829) );
  NANDN U6101 ( .A(n5818), .B(n5817), .Z(n5822) );
  OR U6102 ( .A(n5820), .B(n5819), .Z(n5821) );
  AND U6103 ( .A(n5822), .B(n5821), .Z(n5828) );
  XOR U6104 ( .A(n5829), .B(n5828), .Z(n5831) );
  XOR U6105 ( .A(n5830), .B(n5831), .Z(n5846) );
  XNOR U6106 ( .A(n5846), .B(sreg[506]), .Z(n5848) );
  NANDN U6107 ( .A(n5823), .B(sreg[505]), .Z(n5827) );
  NAND U6108 ( .A(n5825), .B(n5824), .Z(n5826) );
  NAND U6109 ( .A(n5827), .B(n5826), .Z(n5847) );
  XOR U6110 ( .A(n5848), .B(n5847), .Z(c[506]) );
  NANDN U6111 ( .A(n5829), .B(n5828), .Z(n5833) );
  OR U6112 ( .A(n5831), .B(n5830), .Z(n5832) );
  AND U6113 ( .A(n5833), .B(n5832), .Z(n5854) );
  NANDN U6114 ( .A(n30), .B(n5834), .Z(n5836) );
  XNOR U6115 ( .A(b[3]), .B(a[253]), .Z(n5855) );
  OR U6116 ( .A(n5855), .B(n5891), .Z(n5835) );
  NAND U6117 ( .A(n5836), .B(n5835), .Z(n5860) );
  NAND U6118 ( .A(b[0]), .B(a[255]), .Z(n5837) );
  XNOR U6119 ( .A(b[1]), .B(n5837), .Z(n5839) );
  NANDN U6120 ( .A(b[0]), .B(a[254]), .Z(n5838) );
  NAND U6121 ( .A(n5839), .B(n5838), .Z(n5859) );
  NAND U6122 ( .A(b[3]), .B(a[251]), .Z(n5858) );
  XNOR U6123 ( .A(n5859), .B(n5858), .Z(n5861) );
  XNOR U6124 ( .A(n5860), .B(n5861), .Z(n5851) );
  NANDN U6125 ( .A(n5841), .B(n5840), .Z(n5845) );
  OR U6126 ( .A(n5843), .B(n5842), .Z(n5844) );
  AND U6127 ( .A(n5845), .B(n5844), .Z(n5852) );
  XNOR U6128 ( .A(n5851), .B(n5852), .Z(n5853) );
  XNOR U6129 ( .A(n5854), .B(n5853), .Z(n5862) );
  XNOR U6130 ( .A(n5862), .B(sreg[507]), .Z(n5864) );
  NANDN U6131 ( .A(n5846), .B(sreg[506]), .Z(n5850) );
  NAND U6132 ( .A(n5848), .B(n5847), .Z(n5849) );
  NAND U6133 ( .A(n5850), .B(n5849), .Z(n5863) );
  XOR U6134 ( .A(n5864), .B(n5863), .Z(c[507]) );
  OR U6135 ( .A(n5855), .B(n30), .Z(n5857) );
  XNOR U6136 ( .A(b[3]), .B(a[254]), .Z(n5877) );
  OR U6137 ( .A(n5877), .B(n5891), .Z(n5856) );
  AND U6138 ( .A(n5857), .B(n5856), .Z(n5873) );
  AND U6139 ( .A(b[3]), .B(a[252]), .Z(n5874) );
  XNOR U6140 ( .A(n5873), .B(n5874), .Z(n5876) );
  XNOR U6141 ( .A(n5875), .B(n5876), .Z(n5868) );
  XOR U6142 ( .A(n5868), .B(n5867), .Z(n5870) );
  XOR U6143 ( .A(n5869), .B(n5870), .Z(n5866) );
  XOR U6144 ( .A(n5866), .B(n5865), .Z(c[508]) );
  AND U6145 ( .A(n5866), .B(n5865), .Z(n5895) );
  NANDN U6146 ( .A(n5868), .B(n5867), .Z(n5872) );
  NANDN U6147 ( .A(n5870), .B(n5869), .Z(n5871) );
  NAND U6148 ( .A(n5872), .B(n5871), .Z(n5882) );
  OR U6149 ( .A(n5877), .B(n30), .Z(n5879) );
  XNOR U6150 ( .A(a[255]), .B(b[3]), .Z(n5890) );
  OR U6151 ( .A(n5890), .B(n5891), .Z(n5878) );
  AND U6152 ( .A(n5879), .B(n5878), .Z(n5886) );
  NAND U6153 ( .A(b[3]), .B(a[253]), .Z(n5902) );
  XNOR U6154 ( .A(b[1]), .B(n5902), .Z(n5887) );
  XNOR U6155 ( .A(n5881), .B(n5880), .Z(n5883) );
  XOR U6156 ( .A(n5882), .B(n5883), .Z(n5894) );
  XOR U6157 ( .A(n5895), .B(n5894), .Z(c[509]) );
  NAND U6158 ( .A(n5881), .B(n5880), .Z(n5885) );
  NANDN U6159 ( .A(n5883), .B(n5882), .Z(n5884) );
  AND U6160 ( .A(n5885), .B(n5884), .Z(n5901) );
  NANDN U6161 ( .A(n5902), .B(b[1]), .Z(n5889) );
  NAND U6162 ( .A(n5887), .B(n5886), .Z(n5888) );
  AND U6163 ( .A(n5889), .B(n5888), .Z(n5900) );
  XOR U6164 ( .A(n5901), .B(n5900), .Z(n5897) );
  OR U6165 ( .A(n5890), .B(n30), .Z(n5893) );
  NANDN U6166 ( .A(n5891), .B(b[3]), .Z(n5892) );
  NAND U6167 ( .A(n5893), .B(n5892), .Z(n5905) );
  AND U6168 ( .A(b[3]), .B(a[254]), .Z(n5903) );
  XOR U6169 ( .A(n5902), .B(n5903), .Z(n5904) );
  NAND U6170 ( .A(n5895), .B(n5894), .Z(n5898) );
  XOR U6171 ( .A(n5899), .B(n5898), .Z(n5896) );
  XNOR U6172 ( .A(n5897), .B(n5896), .Z(c[510]) );
endmodule

