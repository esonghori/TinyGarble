
module mult_N128_CC128 ( clk, rst, a, b, c );
  input [127:0] a;
  input [0:0] b;
  output [255:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762;
  wire   [255:0] sreg;

  DFF \sreg_reg[254]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(sreg[254]) );
  DFF \sreg_reg[253]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(sreg[253]) );
  DFF \sreg_reg[252]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(sreg[252]) );
  DFF \sreg_reg[251]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(sreg[251]) );
  DFF \sreg_reg[250]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(sreg[250]) );
  DFF \sreg_reg[249]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(sreg[249]) );
  DFF \sreg_reg[248]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(sreg[248]) );
  DFF \sreg_reg[247]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(sreg[247]) );
  DFF \sreg_reg[246]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(sreg[246]) );
  DFF \sreg_reg[245]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(sreg[245]) );
  DFF \sreg_reg[244]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(sreg[244]) );
  DFF \sreg_reg[243]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(sreg[243]) );
  DFF \sreg_reg[242]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(sreg[242]) );
  DFF \sreg_reg[241]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(sreg[241]) );
  DFF \sreg_reg[240]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(sreg[240]) );
  DFF \sreg_reg[239]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(sreg[239]) );
  DFF \sreg_reg[238]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(sreg[238]) );
  DFF \sreg_reg[237]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(sreg[237]) );
  DFF \sreg_reg[236]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(sreg[236]) );
  DFF \sreg_reg[235]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(sreg[235]) );
  DFF \sreg_reg[234]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(sreg[234]) );
  DFF \sreg_reg[233]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(sreg[233]) );
  DFF \sreg_reg[232]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(sreg[232]) );
  DFF \sreg_reg[231]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(sreg[231]) );
  DFF \sreg_reg[230]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(sreg[230]) );
  DFF \sreg_reg[229]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(sreg[229]) );
  DFF \sreg_reg[228]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(sreg[228]) );
  DFF \sreg_reg[227]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(sreg[227]) );
  DFF \sreg_reg[226]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(sreg[226]) );
  DFF \sreg_reg[225]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(sreg[225]) );
  DFF \sreg_reg[224]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(sreg[224]) );
  DFF \sreg_reg[223]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(sreg[223]) );
  DFF \sreg_reg[222]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(sreg[222]) );
  DFF \sreg_reg[221]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(sreg[221]) );
  DFF \sreg_reg[220]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(sreg[220]) );
  DFF \sreg_reg[219]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(sreg[219]) );
  DFF \sreg_reg[218]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(sreg[218]) );
  DFF \sreg_reg[217]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(sreg[217]) );
  DFF \sreg_reg[216]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(sreg[216]) );
  DFF \sreg_reg[215]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(sreg[215]) );
  DFF \sreg_reg[214]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(sreg[214]) );
  DFF \sreg_reg[213]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(sreg[213]) );
  DFF \sreg_reg[212]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(sreg[212]) );
  DFF \sreg_reg[211]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(sreg[211]) );
  DFF \sreg_reg[210]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(sreg[210]) );
  DFF \sreg_reg[209]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(sreg[209]) );
  DFF \sreg_reg[208]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(sreg[208]) );
  DFF \sreg_reg[207]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(sreg[207]) );
  DFF \sreg_reg[206]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(sreg[206]) );
  DFF \sreg_reg[205]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(sreg[205]) );
  DFF \sreg_reg[204]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(sreg[204]) );
  DFF \sreg_reg[203]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(sreg[203]) );
  DFF \sreg_reg[202]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(sreg[202]) );
  DFF \sreg_reg[201]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(sreg[201]) );
  DFF \sreg_reg[200]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(sreg[200]) );
  DFF \sreg_reg[199]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(sreg[199]) );
  DFF \sreg_reg[198]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(sreg[198]) );
  DFF \sreg_reg[197]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(sreg[197]) );
  DFF \sreg_reg[196]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(sreg[196]) );
  DFF \sreg_reg[195]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(sreg[195]) );
  DFF \sreg_reg[194]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(sreg[194]) );
  DFF \sreg_reg[193]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(sreg[193]) );
  DFF \sreg_reg[192]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(sreg[192]) );
  DFF \sreg_reg[191]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(sreg[191]) );
  DFF \sreg_reg[190]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(sreg[190]) );
  DFF \sreg_reg[189]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(sreg[189]) );
  DFF \sreg_reg[188]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(sreg[188]) );
  DFF \sreg_reg[187]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(sreg[187]) );
  DFF \sreg_reg[186]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(sreg[186]) );
  DFF \sreg_reg[185]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(sreg[185]) );
  DFF \sreg_reg[184]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(sreg[184]) );
  DFF \sreg_reg[183]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(sreg[183]) );
  DFF \sreg_reg[182]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(sreg[182]) );
  DFF \sreg_reg[181]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(sreg[181]) );
  DFF \sreg_reg[180]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(sreg[180]) );
  DFF \sreg_reg[179]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(sreg[179]) );
  DFF \sreg_reg[178]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(sreg[178]) );
  DFF \sreg_reg[177]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(sreg[177]) );
  DFF \sreg_reg[176]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(sreg[176]) );
  DFF \sreg_reg[175]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(sreg[175]) );
  DFF \sreg_reg[174]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(sreg[174]) );
  DFF \sreg_reg[173]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(sreg[173]) );
  DFF \sreg_reg[172]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(sreg[172]) );
  DFF \sreg_reg[171]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(sreg[171]) );
  DFF \sreg_reg[170]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(sreg[170]) );
  DFF \sreg_reg[169]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(sreg[169]) );
  DFF \sreg_reg[168]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(sreg[168]) );
  DFF \sreg_reg[167]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(sreg[167]) );
  DFF \sreg_reg[166]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(sreg[166]) );
  DFF \sreg_reg[165]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(sreg[165]) );
  DFF \sreg_reg[164]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(sreg[164]) );
  DFF \sreg_reg[163]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(sreg[163]) );
  DFF \sreg_reg[162]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(sreg[162]) );
  DFF \sreg_reg[161]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(sreg[161]) );
  DFF \sreg_reg[160]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(sreg[160]) );
  DFF \sreg_reg[159]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(sreg[159]) );
  DFF \sreg_reg[158]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(sreg[158]) );
  DFF \sreg_reg[157]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(sreg[157]) );
  DFF \sreg_reg[156]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(sreg[156]) );
  DFF \sreg_reg[155]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(sreg[155]) );
  DFF \sreg_reg[154]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(sreg[154]) );
  DFF \sreg_reg[153]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(sreg[153]) );
  DFF \sreg_reg[152]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(sreg[152]) );
  DFF \sreg_reg[151]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(sreg[151]) );
  DFF \sreg_reg[150]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(sreg[150]) );
  DFF \sreg_reg[149]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(sreg[149]) );
  DFF \sreg_reg[148]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(sreg[148]) );
  DFF \sreg_reg[147]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(sreg[147]) );
  DFF \sreg_reg[146]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(sreg[146]) );
  DFF \sreg_reg[145]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(sreg[145]) );
  DFF \sreg_reg[144]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(sreg[144]) );
  DFF \sreg_reg[143]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(sreg[143]) );
  DFF \sreg_reg[142]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(sreg[142]) );
  DFF \sreg_reg[141]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(sreg[141]) );
  DFF \sreg_reg[140]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(sreg[140]) );
  DFF \sreg_reg[139]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(sreg[139]) );
  DFF \sreg_reg[138]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(sreg[138]) );
  DFF \sreg_reg[137]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(sreg[137]) );
  DFF \sreg_reg[136]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(sreg[136]) );
  DFF \sreg_reg[135]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(sreg[135]) );
  DFF \sreg_reg[134]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(sreg[134]) );
  DFF \sreg_reg[133]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(sreg[133]) );
  DFF \sreg_reg[132]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(sreg[132]) );
  DFF \sreg_reg[131]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(sreg[131]) );
  DFF \sreg_reg[130]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(sreg[130]) );
  DFF \sreg_reg[129]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(sreg[129]) );
  DFF \sreg_reg[128]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(sreg[128]) );
  DFF \sreg_reg[127]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(sreg[127]) );
  DFF \sreg_reg[126]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[125]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[1]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XOR U4 ( .A(n381), .B(sreg[128]), .Z(n1) );
  NANDN U5 ( .A(n382), .B(n1), .Z(n2) );
  NAND U6 ( .A(n381), .B(sreg[128]), .Z(n3) );
  AND U7 ( .A(n2), .B(n3), .Z(n385) );
  XOR U8 ( .A(sreg[131]), .B(n390), .Z(n4) );
  NANDN U9 ( .A(n391), .B(n4), .Z(n5) );
  NAND U10 ( .A(sreg[131]), .B(n390), .Z(n6) );
  AND U11 ( .A(n5), .B(n6), .Z(n394) );
  XOR U12 ( .A(sreg[134]), .B(n399), .Z(n7) );
  NANDN U13 ( .A(n400), .B(n7), .Z(n8) );
  NAND U14 ( .A(sreg[134]), .B(n399), .Z(n9) );
  AND U15 ( .A(n8), .B(n9), .Z(n403) );
  XOR U16 ( .A(sreg[137]), .B(n408), .Z(n10) );
  NANDN U17 ( .A(n409), .B(n10), .Z(n11) );
  NAND U18 ( .A(sreg[137]), .B(n408), .Z(n12) );
  AND U19 ( .A(n11), .B(n12), .Z(n412) );
  XOR U20 ( .A(sreg[140]), .B(n417), .Z(n13) );
  NANDN U21 ( .A(n418), .B(n13), .Z(n14) );
  NAND U22 ( .A(sreg[140]), .B(n417), .Z(n15) );
  AND U23 ( .A(n14), .B(n15), .Z(n421) );
  XOR U24 ( .A(sreg[143]), .B(n426), .Z(n16) );
  NANDN U25 ( .A(n427), .B(n16), .Z(n17) );
  NAND U26 ( .A(sreg[143]), .B(n426), .Z(n18) );
  AND U27 ( .A(n17), .B(n18), .Z(n430) );
  XOR U28 ( .A(sreg[146]), .B(n435), .Z(n19) );
  NANDN U29 ( .A(n436), .B(n19), .Z(n20) );
  NAND U30 ( .A(sreg[146]), .B(n435), .Z(n21) );
  AND U31 ( .A(n20), .B(n21), .Z(n439) );
  XOR U32 ( .A(sreg[149]), .B(n444), .Z(n22) );
  NANDN U33 ( .A(n445), .B(n22), .Z(n23) );
  NAND U34 ( .A(sreg[149]), .B(n444), .Z(n24) );
  AND U35 ( .A(n23), .B(n24), .Z(n448) );
  XOR U36 ( .A(sreg[152]), .B(n453), .Z(n25) );
  NANDN U37 ( .A(n454), .B(n25), .Z(n26) );
  NAND U38 ( .A(sreg[152]), .B(n453), .Z(n27) );
  AND U39 ( .A(n26), .B(n27), .Z(n457) );
  XOR U40 ( .A(sreg[155]), .B(n462), .Z(n28) );
  NANDN U41 ( .A(n463), .B(n28), .Z(n29) );
  NAND U42 ( .A(sreg[155]), .B(n462), .Z(n30) );
  AND U43 ( .A(n29), .B(n30), .Z(n466) );
  XOR U44 ( .A(sreg[158]), .B(n471), .Z(n31) );
  NANDN U45 ( .A(n472), .B(n31), .Z(n32) );
  NAND U46 ( .A(sreg[158]), .B(n471), .Z(n33) );
  AND U47 ( .A(n32), .B(n33), .Z(n475) );
  XOR U48 ( .A(sreg[161]), .B(n480), .Z(n34) );
  NANDN U49 ( .A(n481), .B(n34), .Z(n35) );
  NAND U50 ( .A(sreg[161]), .B(n480), .Z(n36) );
  AND U51 ( .A(n35), .B(n36), .Z(n484) );
  XOR U52 ( .A(sreg[164]), .B(n489), .Z(n37) );
  NANDN U53 ( .A(n490), .B(n37), .Z(n38) );
  NAND U54 ( .A(sreg[164]), .B(n489), .Z(n39) );
  AND U55 ( .A(n38), .B(n39), .Z(n493) );
  XOR U56 ( .A(sreg[167]), .B(n498), .Z(n40) );
  NANDN U57 ( .A(n499), .B(n40), .Z(n41) );
  NAND U58 ( .A(sreg[167]), .B(n498), .Z(n42) );
  AND U59 ( .A(n41), .B(n42), .Z(n502) );
  XOR U60 ( .A(sreg[170]), .B(n507), .Z(n43) );
  NANDN U61 ( .A(n508), .B(n43), .Z(n44) );
  NAND U62 ( .A(sreg[170]), .B(n507), .Z(n45) );
  AND U63 ( .A(n44), .B(n45), .Z(n511) );
  XOR U64 ( .A(sreg[173]), .B(n516), .Z(n46) );
  NANDN U65 ( .A(n517), .B(n46), .Z(n47) );
  NAND U66 ( .A(sreg[173]), .B(n516), .Z(n48) );
  AND U67 ( .A(n47), .B(n48), .Z(n520) );
  XOR U68 ( .A(sreg[176]), .B(n525), .Z(n49) );
  NANDN U69 ( .A(n526), .B(n49), .Z(n50) );
  NAND U70 ( .A(sreg[176]), .B(n525), .Z(n51) );
  AND U71 ( .A(n50), .B(n51), .Z(n529) );
  XOR U72 ( .A(sreg[179]), .B(n534), .Z(n52) );
  NANDN U73 ( .A(n535), .B(n52), .Z(n53) );
  NAND U74 ( .A(sreg[179]), .B(n534), .Z(n54) );
  AND U75 ( .A(n53), .B(n54), .Z(n538) );
  XOR U76 ( .A(sreg[182]), .B(n543), .Z(n55) );
  NANDN U77 ( .A(n544), .B(n55), .Z(n56) );
  NAND U78 ( .A(sreg[182]), .B(n543), .Z(n57) );
  AND U79 ( .A(n56), .B(n57), .Z(n547) );
  XOR U80 ( .A(sreg[185]), .B(n552), .Z(n58) );
  NANDN U81 ( .A(n553), .B(n58), .Z(n59) );
  NAND U82 ( .A(sreg[185]), .B(n552), .Z(n60) );
  AND U83 ( .A(n59), .B(n60), .Z(n556) );
  XOR U84 ( .A(sreg[188]), .B(n561), .Z(n61) );
  NANDN U85 ( .A(n562), .B(n61), .Z(n62) );
  NAND U86 ( .A(sreg[188]), .B(n561), .Z(n63) );
  AND U87 ( .A(n62), .B(n63), .Z(n565) );
  XOR U88 ( .A(sreg[191]), .B(n570), .Z(n64) );
  NANDN U89 ( .A(n571), .B(n64), .Z(n65) );
  NAND U90 ( .A(sreg[191]), .B(n570), .Z(n66) );
  AND U91 ( .A(n65), .B(n66), .Z(n574) );
  XOR U92 ( .A(sreg[194]), .B(n579), .Z(n67) );
  NANDN U93 ( .A(n580), .B(n67), .Z(n68) );
  NAND U94 ( .A(sreg[194]), .B(n579), .Z(n69) );
  AND U95 ( .A(n68), .B(n69), .Z(n583) );
  XOR U96 ( .A(sreg[197]), .B(n588), .Z(n70) );
  NANDN U97 ( .A(n589), .B(n70), .Z(n71) );
  NAND U98 ( .A(sreg[197]), .B(n588), .Z(n72) );
  AND U99 ( .A(n71), .B(n72), .Z(n592) );
  XOR U100 ( .A(sreg[200]), .B(n597), .Z(n73) );
  NANDN U101 ( .A(n598), .B(n73), .Z(n74) );
  NAND U102 ( .A(sreg[200]), .B(n597), .Z(n75) );
  AND U103 ( .A(n74), .B(n75), .Z(n601) );
  XOR U104 ( .A(sreg[203]), .B(n606), .Z(n76) );
  NANDN U105 ( .A(n607), .B(n76), .Z(n77) );
  NAND U106 ( .A(sreg[203]), .B(n606), .Z(n78) );
  AND U107 ( .A(n77), .B(n78), .Z(n610) );
  XOR U108 ( .A(sreg[206]), .B(n615), .Z(n79) );
  NANDN U109 ( .A(n616), .B(n79), .Z(n80) );
  NAND U110 ( .A(sreg[206]), .B(n615), .Z(n81) );
  AND U111 ( .A(n80), .B(n81), .Z(n619) );
  XOR U112 ( .A(sreg[209]), .B(n624), .Z(n82) );
  NANDN U113 ( .A(n625), .B(n82), .Z(n83) );
  NAND U114 ( .A(sreg[209]), .B(n624), .Z(n84) );
  AND U115 ( .A(n83), .B(n84), .Z(n628) );
  XOR U116 ( .A(sreg[212]), .B(n633), .Z(n85) );
  NANDN U117 ( .A(n634), .B(n85), .Z(n86) );
  NAND U118 ( .A(sreg[212]), .B(n633), .Z(n87) );
  AND U119 ( .A(n86), .B(n87), .Z(n637) );
  XOR U120 ( .A(sreg[215]), .B(n642), .Z(n88) );
  NANDN U121 ( .A(n643), .B(n88), .Z(n89) );
  NAND U122 ( .A(sreg[215]), .B(n642), .Z(n90) );
  AND U123 ( .A(n89), .B(n90), .Z(n646) );
  XOR U124 ( .A(sreg[218]), .B(n651), .Z(n91) );
  NANDN U125 ( .A(n652), .B(n91), .Z(n92) );
  NAND U126 ( .A(sreg[218]), .B(n651), .Z(n93) );
  AND U127 ( .A(n92), .B(n93), .Z(n655) );
  XOR U128 ( .A(sreg[221]), .B(n660), .Z(n94) );
  NANDN U129 ( .A(n661), .B(n94), .Z(n95) );
  NAND U130 ( .A(sreg[221]), .B(n660), .Z(n96) );
  AND U131 ( .A(n95), .B(n96), .Z(n664) );
  XOR U132 ( .A(sreg[224]), .B(n669), .Z(n97) );
  NANDN U133 ( .A(n670), .B(n97), .Z(n98) );
  NAND U134 ( .A(sreg[224]), .B(n669), .Z(n99) );
  AND U135 ( .A(n98), .B(n99), .Z(n673) );
  XOR U136 ( .A(sreg[227]), .B(n678), .Z(n100) );
  NANDN U137 ( .A(n679), .B(n100), .Z(n101) );
  NAND U138 ( .A(sreg[227]), .B(n678), .Z(n102) );
  AND U139 ( .A(n101), .B(n102), .Z(n682) );
  XOR U140 ( .A(sreg[230]), .B(n687), .Z(n103) );
  NANDN U141 ( .A(n688), .B(n103), .Z(n104) );
  NAND U142 ( .A(sreg[230]), .B(n687), .Z(n105) );
  AND U143 ( .A(n104), .B(n105), .Z(n691) );
  XOR U144 ( .A(sreg[233]), .B(n696), .Z(n106) );
  NANDN U145 ( .A(n697), .B(n106), .Z(n107) );
  NAND U146 ( .A(sreg[233]), .B(n696), .Z(n108) );
  AND U147 ( .A(n107), .B(n108), .Z(n700) );
  XOR U148 ( .A(sreg[236]), .B(n705), .Z(n109) );
  NANDN U149 ( .A(n706), .B(n109), .Z(n110) );
  NAND U150 ( .A(sreg[236]), .B(n705), .Z(n111) );
  AND U151 ( .A(n110), .B(n111), .Z(n709) );
  XOR U152 ( .A(sreg[239]), .B(n714), .Z(n112) );
  NANDN U153 ( .A(n715), .B(n112), .Z(n113) );
  NAND U154 ( .A(sreg[239]), .B(n714), .Z(n114) );
  AND U155 ( .A(n113), .B(n114), .Z(n718) );
  XOR U156 ( .A(sreg[242]), .B(n723), .Z(n115) );
  NANDN U157 ( .A(n724), .B(n115), .Z(n116) );
  NAND U158 ( .A(sreg[242]), .B(n723), .Z(n117) );
  AND U159 ( .A(n116), .B(n117), .Z(n727) );
  XOR U160 ( .A(sreg[245]), .B(n732), .Z(n118) );
  NANDN U161 ( .A(n733), .B(n118), .Z(n119) );
  NAND U162 ( .A(sreg[245]), .B(n732), .Z(n120) );
  AND U163 ( .A(n119), .B(n120), .Z(n736) );
  XOR U164 ( .A(sreg[248]), .B(n741), .Z(n121) );
  NANDN U165 ( .A(n742), .B(n121), .Z(n122) );
  NAND U166 ( .A(sreg[248]), .B(n741), .Z(n123) );
  AND U167 ( .A(n122), .B(n123), .Z(n745) );
  XOR U168 ( .A(sreg[251]), .B(n750), .Z(n124) );
  NANDN U169 ( .A(n751), .B(n124), .Z(n125) );
  NAND U170 ( .A(sreg[251]), .B(n750), .Z(n126) );
  AND U171 ( .A(n125), .B(n126), .Z(n754) );
  XOR U172 ( .A(sreg[129]), .B(n384), .Z(n127) );
  NANDN U173 ( .A(n385), .B(n127), .Z(n128) );
  NAND U174 ( .A(sreg[129]), .B(n384), .Z(n129) );
  AND U175 ( .A(n128), .B(n129), .Z(n388) );
  XOR U176 ( .A(sreg[132]), .B(n393), .Z(n130) );
  NANDN U177 ( .A(n394), .B(n130), .Z(n131) );
  NAND U178 ( .A(sreg[132]), .B(n393), .Z(n132) );
  AND U179 ( .A(n131), .B(n132), .Z(n397) );
  XOR U180 ( .A(sreg[135]), .B(n402), .Z(n133) );
  NANDN U181 ( .A(n403), .B(n133), .Z(n134) );
  NAND U182 ( .A(sreg[135]), .B(n402), .Z(n135) );
  AND U183 ( .A(n134), .B(n135), .Z(n406) );
  XOR U184 ( .A(sreg[138]), .B(n411), .Z(n136) );
  NANDN U185 ( .A(n412), .B(n136), .Z(n137) );
  NAND U186 ( .A(sreg[138]), .B(n411), .Z(n138) );
  AND U187 ( .A(n137), .B(n138), .Z(n415) );
  XOR U188 ( .A(sreg[141]), .B(n420), .Z(n139) );
  NANDN U189 ( .A(n421), .B(n139), .Z(n140) );
  NAND U190 ( .A(sreg[141]), .B(n420), .Z(n141) );
  AND U191 ( .A(n140), .B(n141), .Z(n424) );
  XOR U192 ( .A(sreg[144]), .B(n429), .Z(n142) );
  NANDN U193 ( .A(n430), .B(n142), .Z(n143) );
  NAND U194 ( .A(sreg[144]), .B(n429), .Z(n144) );
  AND U195 ( .A(n143), .B(n144), .Z(n433) );
  XOR U196 ( .A(sreg[147]), .B(n438), .Z(n145) );
  NANDN U197 ( .A(n439), .B(n145), .Z(n146) );
  NAND U198 ( .A(sreg[147]), .B(n438), .Z(n147) );
  AND U199 ( .A(n146), .B(n147), .Z(n442) );
  XOR U200 ( .A(sreg[150]), .B(n447), .Z(n148) );
  NANDN U201 ( .A(n448), .B(n148), .Z(n149) );
  NAND U202 ( .A(sreg[150]), .B(n447), .Z(n150) );
  AND U203 ( .A(n149), .B(n150), .Z(n451) );
  XOR U204 ( .A(sreg[153]), .B(n456), .Z(n151) );
  NANDN U205 ( .A(n457), .B(n151), .Z(n152) );
  NAND U206 ( .A(sreg[153]), .B(n456), .Z(n153) );
  AND U207 ( .A(n152), .B(n153), .Z(n460) );
  XOR U208 ( .A(sreg[156]), .B(n465), .Z(n154) );
  NANDN U209 ( .A(n466), .B(n154), .Z(n155) );
  NAND U210 ( .A(sreg[156]), .B(n465), .Z(n156) );
  AND U211 ( .A(n155), .B(n156), .Z(n469) );
  XOR U212 ( .A(sreg[159]), .B(n474), .Z(n157) );
  NANDN U213 ( .A(n475), .B(n157), .Z(n158) );
  NAND U214 ( .A(sreg[159]), .B(n474), .Z(n159) );
  AND U215 ( .A(n158), .B(n159), .Z(n478) );
  XOR U216 ( .A(sreg[162]), .B(n483), .Z(n160) );
  NANDN U217 ( .A(n484), .B(n160), .Z(n161) );
  NAND U218 ( .A(sreg[162]), .B(n483), .Z(n162) );
  AND U219 ( .A(n161), .B(n162), .Z(n487) );
  XOR U220 ( .A(sreg[165]), .B(n492), .Z(n163) );
  NANDN U221 ( .A(n493), .B(n163), .Z(n164) );
  NAND U222 ( .A(sreg[165]), .B(n492), .Z(n165) );
  AND U223 ( .A(n164), .B(n165), .Z(n496) );
  XOR U224 ( .A(sreg[168]), .B(n501), .Z(n166) );
  NANDN U225 ( .A(n502), .B(n166), .Z(n167) );
  NAND U226 ( .A(sreg[168]), .B(n501), .Z(n168) );
  AND U227 ( .A(n167), .B(n168), .Z(n505) );
  XOR U228 ( .A(sreg[171]), .B(n510), .Z(n169) );
  NANDN U229 ( .A(n511), .B(n169), .Z(n170) );
  NAND U230 ( .A(sreg[171]), .B(n510), .Z(n171) );
  AND U231 ( .A(n170), .B(n171), .Z(n514) );
  XOR U232 ( .A(sreg[174]), .B(n519), .Z(n172) );
  NANDN U233 ( .A(n520), .B(n172), .Z(n173) );
  NAND U234 ( .A(sreg[174]), .B(n519), .Z(n174) );
  AND U235 ( .A(n173), .B(n174), .Z(n523) );
  XOR U236 ( .A(sreg[177]), .B(n528), .Z(n175) );
  NANDN U237 ( .A(n529), .B(n175), .Z(n176) );
  NAND U238 ( .A(sreg[177]), .B(n528), .Z(n177) );
  AND U239 ( .A(n176), .B(n177), .Z(n532) );
  XOR U240 ( .A(sreg[180]), .B(n537), .Z(n178) );
  NANDN U241 ( .A(n538), .B(n178), .Z(n179) );
  NAND U242 ( .A(sreg[180]), .B(n537), .Z(n180) );
  AND U243 ( .A(n179), .B(n180), .Z(n541) );
  XOR U244 ( .A(sreg[183]), .B(n546), .Z(n181) );
  NANDN U245 ( .A(n547), .B(n181), .Z(n182) );
  NAND U246 ( .A(sreg[183]), .B(n546), .Z(n183) );
  AND U247 ( .A(n182), .B(n183), .Z(n550) );
  XOR U248 ( .A(sreg[186]), .B(n555), .Z(n184) );
  NANDN U249 ( .A(n556), .B(n184), .Z(n185) );
  NAND U250 ( .A(sreg[186]), .B(n555), .Z(n186) );
  AND U251 ( .A(n185), .B(n186), .Z(n559) );
  XOR U252 ( .A(sreg[189]), .B(n564), .Z(n187) );
  NANDN U253 ( .A(n565), .B(n187), .Z(n188) );
  NAND U254 ( .A(sreg[189]), .B(n564), .Z(n189) );
  AND U255 ( .A(n188), .B(n189), .Z(n568) );
  XOR U256 ( .A(sreg[192]), .B(n573), .Z(n190) );
  NANDN U257 ( .A(n574), .B(n190), .Z(n191) );
  NAND U258 ( .A(sreg[192]), .B(n573), .Z(n192) );
  AND U259 ( .A(n191), .B(n192), .Z(n577) );
  XOR U260 ( .A(sreg[195]), .B(n582), .Z(n193) );
  NANDN U261 ( .A(n583), .B(n193), .Z(n194) );
  NAND U262 ( .A(sreg[195]), .B(n582), .Z(n195) );
  AND U263 ( .A(n194), .B(n195), .Z(n586) );
  XOR U264 ( .A(sreg[198]), .B(n591), .Z(n196) );
  NANDN U265 ( .A(n592), .B(n196), .Z(n197) );
  NAND U266 ( .A(sreg[198]), .B(n591), .Z(n198) );
  AND U267 ( .A(n197), .B(n198), .Z(n595) );
  XOR U268 ( .A(sreg[201]), .B(n600), .Z(n199) );
  NANDN U269 ( .A(n601), .B(n199), .Z(n200) );
  NAND U270 ( .A(sreg[201]), .B(n600), .Z(n201) );
  AND U271 ( .A(n200), .B(n201), .Z(n604) );
  XOR U272 ( .A(sreg[204]), .B(n609), .Z(n202) );
  NANDN U273 ( .A(n610), .B(n202), .Z(n203) );
  NAND U274 ( .A(sreg[204]), .B(n609), .Z(n204) );
  AND U275 ( .A(n203), .B(n204), .Z(n613) );
  XOR U276 ( .A(sreg[207]), .B(n618), .Z(n205) );
  NANDN U277 ( .A(n619), .B(n205), .Z(n206) );
  NAND U278 ( .A(sreg[207]), .B(n618), .Z(n207) );
  AND U279 ( .A(n206), .B(n207), .Z(n622) );
  XOR U280 ( .A(sreg[210]), .B(n627), .Z(n208) );
  NANDN U281 ( .A(n628), .B(n208), .Z(n209) );
  NAND U282 ( .A(sreg[210]), .B(n627), .Z(n210) );
  AND U283 ( .A(n209), .B(n210), .Z(n631) );
  XOR U284 ( .A(sreg[213]), .B(n636), .Z(n211) );
  NANDN U285 ( .A(n637), .B(n211), .Z(n212) );
  NAND U286 ( .A(sreg[213]), .B(n636), .Z(n213) );
  AND U287 ( .A(n212), .B(n213), .Z(n640) );
  XOR U288 ( .A(sreg[216]), .B(n645), .Z(n214) );
  NANDN U289 ( .A(n646), .B(n214), .Z(n215) );
  NAND U290 ( .A(sreg[216]), .B(n645), .Z(n216) );
  AND U291 ( .A(n215), .B(n216), .Z(n649) );
  XOR U292 ( .A(sreg[219]), .B(n654), .Z(n217) );
  NANDN U293 ( .A(n655), .B(n217), .Z(n218) );
  NAND U294 ( .A(sreg[219]), .B(n654), .Z(n219) );
  AND U295 ( .A(n218), .B(n219), .Z(n658) );
  XOR U296 ( .A(sreg[222]), .B(n663), .Z(n220) );
  NANDN U297 ( .A(n664), .B(n220), .Z(n221) );
  NAND U298 ( .A(sreg[222]), .B(n663), .Z(n222) );
  AND U299 ( .A(n221), .B(n222), .Z(n667) );
  XOR U300 ( .A(sreg[225]), .B(n672), .Z(n223) );
  NANDN U301 ( .A(n673), .B(n223), .Z(n224) );
  NAND U302 ( .A(sreg[225]), .B(n672), .Z(n225) );
  AND U303 ( .A(n224), .B(n225), .Z(n676) );
  XOR U304 ( .A(sreg[228]), .B(n681), .Z(n226) );
  NANDN U305 ( .A(n682), .B(n226), .Z(n227) );
  NAND U306 ( .A(sreg[228]), .B(n681), .Z(n228) );
  AND U307 ( .A(n227), .B(n228), .Z(n685) );
  XOR U308 ( .A(sreg[231]), .B(n690), .Z(n229) );
  NANDN U309 ( .A(n691), .B(n229), .Z(n230) );
  NAND U310 ( .A(sreg[231]), .B(n690), .Z(n231) );
  AND U311 ( .A(n230), .B(n231), .Z(n694) );
  XOR U312 ( .A(sreg[234]), .B(n699), .Z(n232) );
  NANDN U313 ( .A(n700), .B(n232), .Z(n233) );
  NAND U314 ( .A(sreg[234]), .B(n699), .Z(n234) );
  AND U315 ( .A(n233), .B(n234), .Z(n703) );
  XOR U316 ( .A(sreg[237]), .B(n708), .Z(n235) );
  NANDN U317 ( .A(n709), .B(n235), .Z(n236) );
  NAND U318 ( .A(sreg[237]), .B(n708), .Z(n237) );
  AND U319 ( .A(n236), .B(n237), .Z(n712) );
  XOR U320 ( .A(sreg[240]), .B(n717), .Z(n238) );
  NANDN U321 ( .A(n718), .B(n238), .Z(n239) );
  NAND U322 ( .A(sreg[240]), .B(n717), .Z(n240) );
  AND U323 ( .A(n239), .B(n240), .Z(n721) );
  XOR U324 ( .A(sreg[243]), .B(n726), .Z(n241) );
  NANDN U325 ( .A(n727), .B(n241), .Z(n242) );
  NAND U326 ( .A(sreg[243]), .B(n726), .Z(n243) );
  AND U327 ( .A(n242), .B(n243), .Z(n730) );
  XOR U328 ( .A(sreg[246]), .B(n735), .Z(n244) );
  NANDN U329 ( .A(n736), .B(n244), .Z(n245) );
  NAND U330 ( .A(sreg[246]), .B(n735), .Z(n246) );
  AND U331 ( .A(n245), .B(n246), .Z(n739) );
  XOR U332 ( .A(sreg[249]), .B(n744), .Z(n247) );
  NANDN U333 ( .A(n745), .B(n247), .Z(n248) );
  NAND U334 ( .A(sreg[249]), .B(n744), .Z(n249) );
  AND U335 ( .A(n248), .B(n249), .Z(n748) );
  XOR U336 ( .A(sreg[252]), .B(n753), .Z(n250) );
  NANDN U337 ( .A(n754), .B(n250), .Z(n251) );
  NAND U338 ( .A(sreg[252]), .B(n753), .Z(n252) );
  AND U339 ( .A(n251), .B(n252), .Z(n757) );
  XOR U340 ( .A(sreg[130]), .B(n387), .Z(n253) );
  NANDN U341 ( .A(n388), .B(n253), .Z(n254) );
  NAND U342 ( .A(sreg[130]), .B(n387), .Z(n255) );
  AND U343 ( .A(n254), .B(n255), .Z(n391) );
  XOR U344 ( .A(sreg[133]), .B(n396), .Z(n256) );
  NANDN U345 ( .A(n397), .B(n256), .Z(n257) );
  NAND U346 ( .A(sreg[133]), .B(n396), .Z(n258) );
  AND U347 ( .A(n257), .B(n258), .Z(n400) );
  XOR U348 ( .A(sreg[136]), .B(n405), .Z(n259) );
  NANDN U349 ( .A(n406), .B(n259), .Z(n260) );
  NAND U350 ( .A(sreg[136]), .B(n405), .Z(n261) );
  AND U351 ( .A(n260), .B(n261), .Z(n409) );
  XOR U352 ( .A(sreg[139]), .B(n414), .Z(n262) );
  NANDN U353 ( .A(n415), .B(n262), .Z(n263) );
  NAND U354 ( .A(sreg[139]), .B(n414), .Z(n264) );
  AND U355 ( .A(n263), .B(n264), .Z(n418) );
  XOR U356 ( .A(sreg[142]), .B(n423), .Z(n265) );
  NANDN U357 ( .A(n424), .B(n265), .Z(n266) );
  NAND U358 ( .A(sreg[142]), .B(n423), .Z(n267) );
  AND U359 ( .A(n266), .B(n267), .Z(n427) );
  XOR U360 ( .A(sreg[145]), .B(n432), .Z(n268) );
  NANDN U361 ( .A(n433), .B(n268), .Z(n269) );
  NAND U362 ( .A(sreg[145]), .B(n432), .Z(n270) );
  AND U363 ( .A(n269), .B(n270), .Z(n436) );
  XOR U364 ( .A(sreg[148]), .B(n441), .Z(n271) );
  NANDN U365 ( .A(n442), .B(n271), .Z(n272) );
  NAND U366 ( .A(sreg[148]), .B(n441), .Z(n273) );
  AND U367 ( .A(n272), .B(n273), .Z(n445) );
  XOR U368 ( .A(sreg[151]), .B(n450), .Z(n274) );
  NANDN U369 ( .A(n451), .B(n274), .Z(n275) );
  NAND U370 ( .A(sreg[151]), .B(n450), .Z(n276) );
  AND U371 ( .A(n275), .B(n276), .Z(n454) );
  XOR U372 ( .A(sreg[154]), .B(n459), .Z(n277) );
  NANDN U373 ( .A(n460), .B(n277), .Z(n278) );
  NAND U374 ( .A(sreg[154]), .B(n459), .Z(n279) );
  AND U375 ( .A(n278), .B(n279), .Z(n463) );
  XOR U376 ( .A(sreg[157]), .B(n468), .Z(n280) );
  NANDN U377 ( .A(n469), .B(n280), .Z(n281) );
  NAND U378 ( .A(sreg[157]), .B(n468), .Z(n282) );
  AND U379 ( .A(n281), .B(n282), .Z(n472) );
  XOR U380 ( .A(sreg[160]), .B(n477), .Z(n283) );
  NANDN U381 ( .A(n478), .B(n283), .Z(n284) );
  NAND U382 ( .A(sreg[160]), .B(n477), .Z(n285) );
  AND U383 ( .A(n284), .B(n285), .Z(n481) );
  XOR U384 ( .A(sreg[163]), .B(n486), .Z(n286) );
  NANDN U385 ( .A(n487), .B(n286), .Z(n287) );
  NAND U386 ( .A(sreg[163]), .B(n486), .Z(n288) );
  AND U387 ( .A(n287), .B(n288), .Z(n490) );
  XOR U388 ( .A(sreg[166]), .B(n495), .Z(n289) );
  NANDN U389 ( .A(n496), .B(n289), .Z(n290) );
  NAND U390 ( .A(sreg[166]), .B(n495), .Z(n291) );
  AND U391 ( .A(n290), .B(n291), .Z(n499) );
  XOR U392 ( .A(sreg[169]), .B(n504), .Z(n292) );
  NANDN U393 ( .A(n505), .B(n292), .Z(n293) );
  NAND U394 ( .A(sreg[169]), .B(n504), .Z(n294) );
  AND U395 ( .A(n293), .B(n294), .Z(n508) );
  XOR U396 ( .A(sreg[172]), .B(n513), .Z(n295) );
  NANDN U397 ( .A(n514), .B(n295), .Z(n296) );
  NAND U398 ( .A(sreg[172]), .B(n513), .Z(n297) );
  AND U399 ( .A(n296), .B(n297), .Z(n517) );
  XOR U400 ( .A(sreg[175]), .B(n522), .Z(n298) );
  NANDN U401 ( .A(n523), .B(n298), .Z(n299) );
  NAND U402 ( .A(sreg[175]), .B(n522), .Z(n300) );
  AND U403 ( .A(n299), .B(n300), .Z(n526) );
  XOR U404 ( .A(sreg[178]), .B(n531), .Z(n301) );
  NANDN U405 ( .A(n532), .B(n301), .Z(n302) );
  NAND U406 ( .A(sreg[178]), .B(n531), .Z(n303) );
  AND U407 ( .A(n302), .B(n303), .Z(n535) );
  XOR U408 ( .A(sreg[181]), .B(n540), .Z(n304) );
  NANDN U409 ( .A(n541), .B(n304), .Z(n305) );
  NAND U410 ( .A(sreg[181]), .B(n540), .Z(n306) );
  AND U411 ( .A(n305), .B(n306), .Z(n544) );
  XOR U412 ( .A(sreg[184]), .B(n549), .Z(n307) );
  NANDN U413 ( .A(n550), .B(n307), .Z(n308) );
  NAND U414 ( .A(sreg[184]), .B(n549), .Z(n309) );
  AND U415 ( .A(n308), .B(n309), .Z(n553) );
  XOR U416 ( .A(sreg[187]), .B(n558), .Z(n310) );
  NANDN U417 ( .A(n559), .B(n310), .Z(n311) );
  NAND U418 ( .A(sreg[187]), .B(n558), .Z(n312) );
  AND U419 ( .A(n311), .B(n312), .Z(n562) );
  XOR U420 ( .A(sreg[190]), .B(n567), .Z(n313) );
  NANDN U421 ( .A(n568), .B(n313), .Z(n314) );
  NAND U422 ( .A(sreg[190]), .B(n567), .Z(n315) );
  AND U423 ( .A(n314), .B(n315), .Z(n571) );
  XOR U424 ( .A(sreg[193]), .B(n576), .Z(n316) );
  NANDN U425 ( .A(n577), .B(n316), .Z(n317) );
  NAND U426 ( .A(sreg[193]), .B(n576), .Z(n318) );
  AND U427 ( .A(n317), .B(n318), .Z(n580) );
  XOR U428 ( .A(sreg[196]), .B(n585), .Z(n319) );
  NANDN U429 ( .A(n586), .B(n319), .Z(n320) );
  NAND U430 ( .A(sreg[196]), .B(n585), .Z(n321) );
  AND U431 ( .A(n320), .B(n321), .Z(n589) );
  XOR U432 ( .A(sreg[199]), .B(n594), .Z(n322) );
  NANDN U433 ( .A(n595), .B(n322), .Z(n323) );
  NAND U434 ( .A(sreg[199]), .B(n594), .Z(n324) );
  AND U435 ( .A(n323), .B(n324), .Z(n598) );
  XOR U436 ( .A(sreg[202]), .B(n603), .Z(n325) );
  NANDN U437 ( .A(n604), .B(n325), .Z(n326) );
  NAND U438 ( .A(sreg[202]), .B(n603), .Z(n327) );
  AND U439 ( .A(n326), .B(n327), .Z(n607) );
  XOR U440 ( .A(sreg[205]), .B(n612), .Z(n328) );
  NANDN U441 ( .A(n613), .B(n328), .Z(n329) );
  NAND U442 ( .A(sreg[205]), .B(n612), .Z(n330) );
  AND U443 ( .A(n329), .B(n330), .Z(n616) );
  XOR U444 ( .A(sreg[208]), .B(n621), .Z(n331) );
  NANDN U445 ( .A(n622), .B(n331), .Z(n332) );
  NAND U446 ( .A(sreg[208]), .B(n621), .Z(n333) );
  AND U447 ( .A(n332), .B(n333), .Z(n625) );
  XOR U448 ( .A(sreg[211]), .B(n630), .Z(n334) );
  NANDN U449 ( .A(n631), .B(n334), .Z(n335) );
  NAND U450 ( .A(sreg[211]), .B(n630), .Z(n336) );
  AND U451 ( .A(n335), .B(n336), .Z(n634) );
  XOR U452 ( .A(sreg[214]), .B(n639), .Z(n337) );
  NANDN U453 ( .A(n640), .B(n337), .Z(n338) );
  NAND U454 ( .A(sreg[214]), .B(n639), .Z(n339) );
  AND U455 ( .A(n338), .B(n339), .Z(n643) );
  XOR U456 ( .A(sreg[217]), .B(n648), .Z(n340) );
  NANDN U457 ( .A(n649), .B(n340), .Z(n341) );
  NAND U458 ( .A(sreg[217]), .B(n648), .Z(n342) );
  AND U459 ( .A(n341), .B(n342), .Z(n652) );
  XOR U460 ( .A(sreg[220]), .B(n657), .Z(n343) );
  NANDN U461 ( .A(n658), .B(n343), .Z(n344) );
  NAND U462 ( .A(sreg[220]), .B(n657), .Z(n345) );
  AND U463 ( .A(n344), .B(n345), .Z(n661) );
  XOR U464 ( .A(sreg[223]), .B(n666), .Z(n346) );
  NANDN U465 ( .A(n667), .B(n346), .Z(n347) );
  NAND U466 ( .A(sreg[223]), .B(n666), .Z(n348) );
  AND U467 ( .A(n347), .B(n348), .Z(n670) );
  XOR U468 ( .A(sreg[226]), .B(n675), .Z(n349) );
  NANDN U469 ( .A(n676), .B(n349), .Z(n350) );
  NAND U470 ( .A(sreg[226]), .B(n675), .Z(n351) );
  AND U471 ( .A(n350), .B(n351), .Z(n679) );
  XOR U472 ( .A(sreg[229]), .B(n684), .Z(n352) );
  NANDN U473 ( .A(n685), .B(n352), .Z(n353) );
  NAND U474 ( .A(sreg[229]), .B(n684), .Z(n354) );
  AND U475 ( .A(n353), .B(n354), .Z(n688) );
  XOR U476 ( .A(sreg[232]), .B(n693), .Z(n355) );
  NANDN U477 ( .A(n694), .B(n355), .Z(n356) );
  NAND U478 ( .A(sreg[232]), .B(n693), .Z(n357) );
  AND U479 ( .A(n356), .B(n357), .Z(n697) );
  XOR U480 ( .A(sreg[235]), .B(n702), .Z(n358) );
  NANDN U481 ( .A(n703), .B(n358), .Z(n359) );
  NAND U482 ( .A(sreg[235]), .B(n702), .Z(n360) );
  AND U483 ( .A(n359), .B(n360), .Z(n706) );
  XOR U484 ( .A(sreg[238]), .B(n711), .Z(n361) );
  NANDN U485 ( .A(n712), .B(n361), .Z(n362) );
  NAND U486 ( .A(sreg[238]), .B(n711), .Z(n363) );
  AND U487 ( .A(n362), .B(n363), .Z(n715) );
  XOR U488 ( .A(sreg[241]), .B(n720), .Z(n364) );
  NANDN U489 ( .A(n721), .B(n364), .Z(n365) );
  NAND U490 ( .A(sreg[241]), .B(n720), .Z(n366) );
  AND U491 ( .A(n365), .B(n366), .Z(n724) );
  XOR U492 ( .A(sreg[244]), .B(n729), .Z(n367) );
  NANDN U493 ( .A(n730), .B(n367), .Z(n368) );
  NAND U494 ( .A(sreg[244]), .B(n729), .Z(n369) );
  AND U495 ( .A(n368), .B(n369), .Z(n733) );
  XOR U496 ( .A(sreg[247]), .B(n738), .Z(n370) );
  NANDN U497 ( .A(n739), .B(n370), .Z(n371) );
  NAND U498 ( .A(sreg[247]), .B(n738), .Z(n372) );
  AND U499 ( .A(n371), .B(n372), .Z(n742) );
  XOR U500 ( .A(sreg[250]), .B(n747), .Z(n373) );
  NANDN U501 ( .A(n748), .B(n373), .Z(n374) );
  NAND U502 ( .A(sreg[250]), .B(n747), .Z(n375) );
  AND U503 ( .A(n374), .B(n375), .Z(n751) );
  XOR U504 ( .A(sreg[253]), .B(n756), .Z(n376) );
  NANDN U505 ( .A(n757), .B(n376), .Z(n377) );
  NAND U506 ( .A(sreg[253]), .B(n756), .Z(n378) );
  AND U507 ( .A(n377), .B(n378), .Z(n760) );
  AND U508 ( .A(b[0]), .B(a[0]), .Z(n379) );
  XOR U509 ( .A(n379), .B(sreg[127]), .Z(c[127]) );
  NAND U510 ( .A(b[0]), .B(a[1]), .Z(n382) );
  AND U511 ( .A(n379), .B(sreg[127]), .Z(n381) );
  XOR U512 ( .A(sreg[128]), .B(n381), .Z(n380) );
  XNOR U513 ( .A(n382), .B(n380), .Z(c[128]) );
  AND U514 ( .A(b[0]), .B(a[2]), .Z(n384) );
  XNOR U515 ( .A(n385), .B(sreg[129]), .Z(n383) );
  XOR U516 ( .A(n384), .B(n383), .Z(c[129]) );
  AND U517 ( .A(b[0]), .B(a[3]), .Z(n387) );
  XNOR U518 ( .A(n388), .B(sreg[130]), .Z(n386) );
  XOR U519 ( .A(n387), .B(n386), .Z(c[130]) );
  AND U520 ( .A(b[0]), .B(a[4]), .Z(n390) );
  XNOR U521 ( .A(n391), .B(sreg[131]), .Z(n389) );
  XOR U522 ( .A(n390), .B(n389), .Z(c[131]) );
  AND U523 ( .A(b[0]), .B(a[5]), .Z(n393) );
  XNOR U524 ( .A(n394), .B(sreg[132]), .Z(n392) );
  XOR U525 ( .A(n393), .B(n392), .Z(c[132]) );
  AND U526 ( .A(b[0]), .B(a[6]), .Z(n396) );
  XNOR U527 ( .A(n397), .B(sreg[133]), .Z(n395) );
  XOR U528 ( .A(n396), .B(n395), .Z(c[133]) );
  AND U529 ( .A(b[0]), .B(a[7]), .Z(n399) );
  XNOR U530 ( .A(n400), .B(sreg[134]), .Z(n398) );
  XOR U531 ( .A(n399), .B(n398), .Z(c[134]) );
  AND U532 ( .A(b[0]), .B(a[8]), .Z(n402) );
  XNOR U533 ( .A(n403), .B(sreg[135]), .Z(n401) );
  XOR U534 ( .A(n402), .B(n401), .Z(c[135]) );
  AND U535 ( .A(b[0]), .B(a[9]), .Z(n405) );
  XNOR U536 ( .A(n406), .B(sreg[136]), .Z(n404) );
  XOR U537 ( .A(n405), .B(n404), .Z(c[136]) );
  AND U538 ( .A(b[0]), .B(a[10]), .Z(n408) );
  XNOR U539 ( .A(n409), .B(sreg[137]), .Z(n407) );
  XOR U540 ( .A(n408), .B(n407), .Z(c[137]) );
  AND U541 ( .A(b[0]), .B(a[11]), .Z(n411) );
  XNOR U542 ( .A(n412), .B(sreg[138]), .Z(n410) );
  XOR U543 ( .A(n411), .B(n410), .Z(c[138]) );
  AND U544 ( .A(b[0]), .B(a[12]), .Z(n414) );
  XNOR U545 ( .A(n415), .B(sreg[139]), .Z(n413) );
  XOR U546 ( .A(n414), .B(n413), .Z(c[139]) );
  AND U547 ( .A(b[0]), .B(a[13]), .Z(n417) );
  XNOR U548 ( .A(n418), .B(sreg[140]), .Z(n416) );
  XOR U549 ( .A(n417), .B(n416), .Z(c[140]) );
  AND U550 ( .A(b[0]), .B(a[14]), .Z(n420) );
  XNOR U551 ( .A(n421), .B(sreg[141]), .Z(n419) );
  XOR U552 ( .A(n420), .B(n419), .Z(c[141]) );
  AND U553 ( .A(b[0]), .B(a[15]), .Z(n423) );
  XNOR U554 ( .A(n424), .B(sreg[142]), .Z(n422) );
  XOR U555 ( .A(n423), .B(n422), .Z(c[142]) );
  AND U556 ( .A(b[0]), .B(a[16]), .Z(n426) );
  XNOR U557 ( .A(n427), .B(sreg[143]), .Z(n425) );
  XOR U558 ( .A(n426), .B(n425), .Z(c[143]) );
  AND U559 ( .A(b[0]), .B(a[17]), .Z(n429) );
  XNOR U560 ( .A(n430), .B(sreg[144]), .Z(n428) );
  XOR U561 ( .A(n429), .B(n428), .Z(c[144]) );
  AND U562 ( .A(b[0]), .B(a[18]), .Z(n432) );
  XNOR U563 ( .A(n433), .B(sreg[145]), .Z(n431) );
  XOR U564 ( .A(n432), .B(n431), .Z(c[145]) );
  AND U565 ( .A(b[0]), .B(a[19]), .Z(n435) );
  XNOR U566 ( .A(n436), .B(sreg[146]), .Z(n434) );
  XOR U567 ( .A(n435), .B(n434), .Z(c[146]) );
  AND U568 ( .A(b[0]), .B(a[20]), .Z(n438) );
  XNOR U569 ( .A(n439), .B(sreg[147]), .Z(n437) );
  XOR U570 ( .A(n438), .B(n437), .Z(c[147]) );
  AND U571 ( .A(b[0]), .B(a[21]), .Z(n441) );
  XNOR U572 ( .A(n442), .B(sreg[148]), .Z(n440) );
  XOR U573 ( .A(n441), .B(n440), .Z(c[148]) );
  AND U574 ( .A(b[0]), .B(a[22]), .Z(n444) );
  XNOR U575 ( .A(n445), .B(sreg[149]), .Z(n443) );
  XOR U576 ( .A(n444), .B(n443), .Z(c[149]) );
  AND U577 ( .A(b[0]), .B(a[23]), .Z(n447) );
  XNOR U578 ( .A(n448), .B(sreg[150]), .Z(n446) );
  XOR U579 ( .A(n447), .B(n446), .Z(c[150]) );
  AND U580 ( .A(b[0]), .B(a[24]), .Z(n450) );
  XNOR U581 ( .A(n451), .B(sreg[151]), .Z(n449) );
  XOR U582 ( .A(n450), .B(n449), .Z(c[151]) );
  AND U583 ( .A(b[0]), .B(a[25]), .Z(n453) );
  XNOR U584 ( .A(n454), .B(sreg[152]), .Z(n452) );
  XOR U585 ( .A(n453), .B(n452), .Z(c[152]) );
  AND U586 ( .A(b[0]), .B(a[26]), .Z(n456) );
  XNOR U587 ( .A(n457), .B(sreg[153]), .Z(n455) );
  XOR U588 ( .A(n456), .B(n455), .Z(c[153]) );
  AND U589 ( .A(b[0]), .B(a[27]), .Z(n459) );
  XNOR U590 ( .A(n460), .B(sreg[154]), .Z(n458) );
  XOR U591 ( .A(n459), .B(n458), .Z(c[154]) );
  AND U592 ( .A(b[0]), .B(a[28]), .Z(n462) );
  XNOR U593 ( .A(n463), .B(sreg[155]), .Z(n461) );
  XOR U594 ( .A(n462), .B(n461), .Z(c[155]) );
  AND U595 ( .A(b[0]), .B(a[29]), .Z(n465) );
  XNOR U596 ( .A(n466), .B(sreg[156]), .Z(n464) );
  XOR U597 ( .A(n465), .B(n464), .Z(c[156]) );
  AND U598 ( .A(b[0]), .B(a[30]), .Z(n468) );
  XNOR U599 ( .A(n469), .B(sreg[157]), .Z(n467) );
  XOR U600 ( .A(n468), .B(n467), .Z(c[157]) );
  AND U601 ( .A(b[0]), .B(a[31]), .Z(n471) );
  XNOR U602 ( .A(n472), .B(sreg[158]), .Z(n470) );
  XOR U603 ( .A(n471), .B(n470), .Z(c[158]) );
  AND U604 ( .A(b[0]), .B(a[32]), .Z(n474) );
  XNOR U605 ( .A(n475), .B(sreg[159]), .Z(n473) );
  XOR U606 ( .A(n474), .B(n473), .Z(c[159]) );
  AND U607 ( .A(b[0]), .B(a[33]), .Z(n477) );
  XNOR U608 ( .A(n478), .B(sreg[160]), .Z(n476) );
  XOR U609 ( .A(n477), .B(n476), .Z(c[160]) );
  AND U610 ( .A(b[0]), .B(a[34]), .Z(n480) );
  XNOR U611 ( .A(n481), .B(sreg[161]), .Z(n479) );
  XOR U612 ( .A(n480), .B(n479), .Z(c[161]) );
  AND U613 ( .A(b[0]), .B(a[35]), .Z(n483) );
  XNOR U614 ( .A(n484), .B(sreg[162]), .Z(n482) );
  XOR U615 ( .A(n483), .B(n482), .Z(c[162]) );
  AND U616 ( .A(b[0]), .B(a[36]), .Z(n486) );
  XNOR U617 ( .A(n487), .B(sreg[163]), .Z(n485) );
  XOR U618 ( .A(n486), .B(n485), .Z(c[163]) );
  AND U619 ( .A(b[0]), .B(a[37]), .Z(n489) );
  XNOR U620 ( .A(n490), .B(sreg[164]), .Z(n488) );
  XOR U621 ( .A(n489), .B(n488), .Z(c[164]) );
  AND U622 ( .A(b[0]), .B(a[38]), .Z(n492) );
  XNOR U623 ( .A(n493), .B(sreg[165]), .Z(n491) );
  XOR U624 ( .A(n492), .B(n491), .Z(c[165]) );
  AND U625 ( .A(b[0]), .B(a[39]), .Z(n495) );
  XNOR U626 ( .A(n496), .B(sreg[166]), .Z(n494) );
  XOR U627 ( .A(n495), .B(n494), .Z(c[166]) );
  AND U628 ( .A(b[0]), .B(a[40]), .Z(n498) );
  XNOR U629 ( .A(n499), .B(sreg[167]), .Z(n497) );
  XOR U630 ( .A(n498), .B(n497), .Z(c[167]) );
  AND U631 ( .A(b[0]), .B(a[41]), .Z(n501) );
  XNOR U632 ( .A(n502), .B(sreg[168]), .Z(n500) );
  XOR U633 ( .A(n501), .B(n500), .Z(c[168]) );
  AND U634 ( .A(b[0]), .B(a[42]), .Z(n504) );
  XNOR U635 ( .A(n505), .B(sreg[169]), .Z(n503) );
  XOR U636 ( .A(n504), .B(n503), .Z(c[169]) );
  AND U637 ( .A(b[0]), .B(a[43]), .Z(n507) );
  XNOR U638 ( .A(n508), .B(sreg[170]), .Z(n506) );
  XOR U639 ( .A(n507), .B(n506), .Z(c[170]) );
  AND U640 ( .A(b[0]), .B(a[44]), .Z(n510) );
  XNOR U641 ( .A(n511), .B(sreg[171]), .Z(n509) );
  XOR U642 ( .A(n510), .B(n509), .Z(c[171]) );
  AND U643 ( .A(b[0]), .B(a[45]), .Z(n513) );
  XNOR U644 ( .A(n514), .B(sreg[172]), .Z(n512) );
  XOR U645 ( .A(n513), .B(n512), .Z(c[172]) );
  AND U646 ( .A(b[0]), .B(a[46]), .Z(n516) );
  XNOR U647 ( .A(n517), .B(sreg[173]), .Z(n515) );
  XOR U648 ( .A(n516), .B(n515), .Z(c[173]) );
  AND U649 ( .A(b[0]), .B(a[47]), .Z(n519) );
  XNOR U650 ( .A(n520), .B(sreg[174]), .Z(n518) );
  XOR U651 ( .A(n519), .B(n518), .Z(c[174]) );
  AND U652 ( .A(b[0]), .B(a[48]), .Z(n522) );
  XNOR U653 ( .A(n523), .B(sreg[175]), .Z(n521) );
  XOR U654 ( .A(n522), .B(n521), .Z(c[175]) );
  AND U655 ( .A(b[0]), .B(a[49]), .Z(n525) );
  XNOR U656 ( .A(n526), .B(sreg[176]), .Z(n524) );
  XOR U657 ( .A(n525), .B(n524), .Z(c[176]) );
  AND U658 ( .A(b[0]), .B(a[50]), .Z(n528) );
  XNOR U659 ( .A(n529), .B(sreg[177]), .Z(n527) );
  XOR U660 ( .A(n528), .B(n527), .Z(c[177]) );
  AND U661 ( .A(b[0]), .B(a[51]), .Z(n531) );
  XNOR U662 ( .A(n532), .B(sreg[178]), .Z(n530) );
  XOR U663 ( .A(n531), .B(n530), .Z(c[178]) );
  AND U664 ( .A(b[0]), .B(a[52]), .Z(n534) );
  XNOR U665 ( .A(n535), .B(sreg[179]), .Z(n533) );
  XOR U666 ( .A(n534), .B(n533), .Z(c[179]) );
  AND U667 ( .A(b[0]), .B(a[53]), .Z(n537) );
  XNOR U668 ( .A(n538), .B(sreg[180]), .Z(n536) );
  XOR U669 ( .A(n537), .B(n536), .Z(c[180]) );
  AND U670 ( .A(b[0]), .B(a[54]), .Z(n540) );
  XNOR U671 ( .A(n541), .B(sreg[181]), .Z(n539) );
  XOR U672 ( .A(n540), .B(n539), .Z(c[181]) );
  AND U673 ( .A(b[0]), .B(a[55]), .Z(n543) );
  XNOR U674 ( .A(n544), .B(sreg[182]), .Z(n542) );
  XOR U675 ( .A(n543), .B(n542), .Z(c[182]) );
  AND U676 ( .A(b[0]), .B(a[56]), .Z(n546) );
  XNOR U677 ( .A(n547), .B(sreg[183]), .Z(n545) );
  XOR U678 ( .A(n546), .B(n545), .Z(c[183]) );
  AND U679 ( .A(b[0]), .B(a[57]), .Z(n549) );
  XNOR U680 ( .A(n550), .B(sreg[184]), .Z(n548) );
  XOR U681 ( .A(n549), .B(n548), .Z(c[184]) );
  AND U682 ( .A(b[0]), .B(a[58]), .Z(n552) );
  XNOR U683 ( .A(n553), .B(sreg[185]), .Z(n551) );
  XOR U684 ( .A(n552), .B(n551), .Z(c[185]) );
  AND U685 ( .A(b[0]), .B(a[59]), .Z(n555) );
  XNOR U686 ( .A(n556), .B(sreg[186]), .Z(n554) );
  XOR U687 ( .A(n555), .B(n554), .Z(c[186]) );
  AND U688 ( .A(b[0]), .B(a[60]), .Z(n558) );
  XNOR U689 ( .A(n559), .B(sreg[187]), .Z(n557) );
  XOR U690 ( .A(n558), .B(n557), .Z(c[187]) );
  AND U691 ( .A(b[0]), .B(a[61]), .Z(n561) );
  XNOR U692 ( .A(n562), .B(sreg[188]), .Z(n560) );
  XOR U693 ( .A(n561), .B(n560), .Z(c[188]) );
  AND U694 ( .A(b[0]), .B(a[62]), .Z(n564) );
  XNOR U695 ( .A(n565), .B(sreg[189]), .Z(n563) );
  XOR U696 ( .A(n564), .B(n563), .Z(c[189]) );
  AND U697 ( .A(b[0]), .B(a[63]), .Z(n567) );
  XNOR U698 ( .A(n568), .B(sreg[190]), .Z(n566) );
  XOR U699 ( .A(n567), .B(n566), .Z(c[190]) );
  AND U700 ( .A(b[0]), .B(a[64]), .Z(n570) );
  XNOR U701 ( .A(n571), .B(sreg[191]), .Z(n569) );
  XOR U702 ( .A(n570), .B(n569), .Z(c[191]) );
  AND U703 ( .A(b[0]), .B(a[65]), .Z(n573) );
  XNOR U704 ( .A(n574), .B(sreg[192]), .Z(n572) );
  XOR U705 ( .A(n573), .B(n572), .Z(c[192]) );
  AND U706 ( .A(b[0]), .B(a[66]), .Z(n576) );
  XNOR U707 ( .A(n577), .B(sreg[193]), .Z(n575) );
  XOR U708 ( .A(n576), .B(n575), .Z(c[193]) );
  AND U709 ( .A(b[0]), .B(a[67]), .Z(n579) );
  XNOR U710 ( .A(n580), .B(sreg[194]), .Z(n578) );
  XOR U711 ( .A(n579), .B(n578), .Z(c[194]) );
  AND U712 ( .A(b[0]), .B(a[68]), .Z(n582) );
  XNOR U713 ( .A(n583), .B(sreg[195]), .Z(n581) );
  XOR U714 ( .A(n582), .B(n581), .Z(c[195]) );
  AND U715 ( .A(b[0]), .B(a[69]), .Z(n585) );
  XNOR U716 ( .A(n586), .B(sreg[196]), .Z(n584) );
  XOR U717 ( .A(n585), .B(n584), .Z(c[196]) );
  AND U718 ( .A(b[0]), .B(a[70]), .Z(n588) );
  XNOR U719 ( .A(n589), .B(sreg[197]), .Z(n587) );
  XOR U720 ( .A(n588), .B(n587), .Z(c[197]) );
  AND U721 ( .A(b[0]), .B(a[71]), .Z(n591) );
  XNOR U722 ( .A(n592), .B(sreg[198]), .Z(n590) );
  XOR U723 ( .A(n591), .B(n590), .Z(c[198]) );
  AND U724 ( .A(b[0]), .B(a[72]), .Z(n594) );
  XNOR U725 ( .A(n595), .B(sreg[199]), .Z(n593) );
  XOR U726 ( .A(n594), .B(n593), .Z(c[199]) );
  AND U727 ( .A(b[0]), .B(a[73]), .Z(n597) );
  XNOR U728 ( .A(n598), .B(sreg[200]), .Z(n596) );
  XOR U729 ( .A(n597), .B(n596), .Z(c[200]) );
  AND U730 ( .A(b[0]), .B(a[74]), .Z(n600) );
  XNOR U731 ( .A(n601), .B(sreg[201]), .Z(n599) );
  XOR U732 ( .A(n600), .B(n599), .Z(c[201]) );
  AND U733 ( .A(b[0]), .B(a[75]), .Z(n603) );
  XNOR U734 ( .A(n604), .B(sreg[202]), .Z(n602) );
  XOR U735 ( .A(n603), .B(n602), .Z(c[202]) );
  AND U736 ( .A(b[0]), .B(a[76]), .Z(n606) );
  XNOR U737 ( .A(n607), .B(sreg[203]), .Z(n605) );
  XOR U738 ( .A(n606), .B(n605), .Z(c[203]) );
  AND U739 ( .A(b[0]), .B(a[77]), .Z(n609) );
  XNOR U740 ( .A(n610), .B(sreg[204]), .Z(n608) );
  XOR U741 ( .A(n609), .B(n608), .Z(c[204]) );
  AND U742 ( .A(b[0]), .B(a[78]), .Z(n612) );
  XNOR U743 ( .A(n613), .B(sreg[205]), .Z(n611) );
  XOR U744 ( .A(n612), .B(n611), .Z(c[205]) );
  AND U745 ( .A(b[0]), .B(a[79]), .Z(n615) );
  XNOR U746 ( .A(n616), .B(sreg[206]), .Z(n614) );
  XOR U747 ( .A(n615), .B(n614), .Z(c[206]) );
  AND U748 ( .A(b[0]), .B(a[80]), .Z(n618) );
  XNOR U749 ( .A(n619), .B(sreg[207]), .Z(n617) );
  XOR U750 ( .A(n618), .B(n617), .Z(c[207]) );
  AND U751 ( .A(b[0]), .B(a[81]), .Z(n621) );
  XNOR U752 ( .A(n622), .B(sreg[208]), .Z(n620) );
  XOR U753 ( .A(n621), .B(n620), .Z(c[208]) );
  AND U754 ( .A(b[0]), .B(a[82]), .Z(n624) );
  XNOR U755 ( .A(n625), .B(sreg[209]), .Z(n623) );
  XOR U756 ( .A(n624), .B(n623), .Z(c[209]) );
  AND U757 ( .A(b[0]), .B(a[83]), .Z(n627) );
  XNOR U758 ( .A(n628), .B(sreg[210]), .Z(n626) );
  XOR U759 ( .A(n627), .B(n626), .Z(c[210]) );
  AND U760 ( .A(b[0]), .B(a[84]), .Z(n630) );
  XNOR U761 ( .A(n631), .B(sreg[211]), .Z(n629) );
  XOR U762 ( .A(n630), .B(n629), .Z(c[211]) );
  AND U763 ( .A(b[0]), .B(a[85]), .Z(n633) );
  XNOR U764 ( .A(n634), .B(sreg[212]), .Z(n632) );
  XOR U765 ( .A(n633), .B(n632), .Z(c[212]) );
  AND U766 ( .A(b[0]), .B(a[86]), .Z(n636) );
  XNOR U767 ( .A(n637), .B(sreg[213]), .Z(n635) );
  XOR U768 ( .A(n636), .B(n635), .Z(c[213]) );
  AND U769 ( .A(b[0]), .B(a[87]), .Z(n639) );
  XNOR U770 ( .A(n640), .B(sreg[214]), .Z(n638) );
  XOR U771 ( .A(n639), .B(n638), .Z(c[214]) );
  AND U772 ( .A(b[0]), .B(a[88]), .Z(n642) );
  XNOR U773 ( .A(n643), .B(sreg[215]), .Z(n641) );
  XOR U774 ( .A(n642), .B(n641), .Z(c[215]) );
  AND U775 ( .A(b[0]), .B(a[89]), .Z(n645) );
  XNOR U776 ( .A(n646), .B(sreg[216]), .Z(n644) );
  XOR U777 ( .A(n645), .B(n644), .Z(c[216]) );
  AND U778 ( .A(b[0]), .B(a[90]), .Z(n648) );
  XNOR U779 ( .A(n649), .B(sreg[217]), .Z(n647) );
  XOR U780 ( .A(n648), .B(n647), .Z(c[217]) );
  AND U781 ( .A(b[0]), .B(a[91]), .Z(n651) );
  XNOR U782 ( .A(n652), .B(sreg[218]), .Z(n650) );
  XOR U783 ( .A(n651), .B(n650), .Z(c[218]) );
  AND U784 ( .A(b[0]), .B(a[92]), .Z(n654) );
  XNOR U785 ( .A(n655), .B(sreg[219]), .Z(n653) );
  XOR U786 ( .A(n654), .B(n653), .Z(c[219]) );
  AND U787 ( .A(b[0]), .B(a[93]), .Z(n657) );
  XNOR U788 ( .A(n658), .B(sreg[220]), .Z(n656) );
  XOR U789 ( .A(n657), .B(n656), .Z(c[220]) );
  AND U790 ( .A(b[0]), .B(a[94]), .Z(n660) );
  XNOR U791 ( .A(n661), .B(sreg[221]), .Z(n659) );
  XOR U792 ( .A(n660), .B(n659), .Z(c[221]) );
  AND U793 ( .A(b[0]), .B(a[95]), .Z(n663) );
  XNOR U794 ( .A(n664), .B(sreg[222]), .Z(n662) );
  XOR U795 ( .A(n663), .B(n662), .Z(c[222]) );
  AND U796 ( .A(b[0]), .B(a[96]), .Z(n666) );
  XNOR U797 ( .A(n667), .B(sreg[223]), .Z(n665) );
  XOR U798 ( .A(n666), .B(n665), .Z(c[223]) );
  AND U799 ( .A(b[0]), .B(a[97]), .Z(n669) );
  XNOR U800 ( .A(n670), .B(sreg[224]), .Z(n668) );
  XOR U801 ( .A(n669), .B(n668), .Z(c[224]) );
  AND U802 ( .A(b[0]), .B(a[98]), .Z(n672) );
  XNOR U803 ( .A(n673), .B(sreg[225]), .Z(n671) );
  XOR U804 ( .A(n672), .B(n671), .Z(c[225]) );
  AND U805 ( .A(b[0]), .B(a[99]), .Z(n675) );
  XNOR U806 ( .A(n676), .B(sreg[226]), .Z(n674) );
  XOR U807 ( .A(n675), .B(n674), .Z(c[226]) );
  AND U808 ( .A(b[0]), .B(a[100]), .Z(n678) );
  XNOR U809 ( .A(n679), .B(sreg[227]), .Z(n677) );
  XOR U810 ( .A(n678), .B(n677), .Z(c[227]) );
  AND U811 ( .A(b[0]), .B(a[101]), .Z(n681) );
  XNOR U812 ( .A(n682), .B(sreg[228]), .Z(n680) );
  XOR U813 ( .A(n681), .B(n680), .Z(c[228]) );
  AND U814 ( .A(b[0]), .B(a[102]), .Z(n684) );
  XNOR U815 ( .A(n685), .B(sreg[229]), .Z(n683) );
  XOR U816 ( .A(n684), .B(n683), .Z(c[229]) );
  AND U817 ( .A(b[0]), .B(a[103]), .Z(n687) );
  XNOR U818 ( .A(n688), .B(sreg[230]), .Z(n686) );
  XOR U819 ( .A(n687), .B(n686), .Z(c[230]) );
  AND U820 ( .A(b[0]), .B(a[104]), .Z(n690) );
  XNOR U821 ( .A(n691), .B(sreg[231]), .Z(n689) );
  XOR U822 ( .A(n690), .B(n689), .Z(c[231]) );
  AND U823 ( .A(b[0]), .B(a[105]), .Z(n693) );
  XNOR U824 ( .A(n694), .B(sreg[232]), .Z(n692) );
  XOR U825 ( .A(n693), .B(n692), .Z(c[232]) );
  AND U826 ( .A(b[0]), .B(a[106]), .Z(n696) );
  XNOR U827 ( .A(n697), .B(sreg[233]), .Z(n695) );
  XOR U828 ( .A(n696), .B(n695), .Z(c[233]) );
  AND U829 ( .A(b[0]), .B(a[107]), .Z(n699) );
  XNOR U830 ( .A(n700), .B(sreg[234]), .Z(n698) );
  XOR U831 ( .A(n699), .B(n698), .Z(c[234]) );
  AND U832 ( .A(b[0]), .B(a[108]), .Z(n702) );
  XNOR U833 ( .A(n703), .B(sreg[235]), .Z(n701) );
  XOR U834 ( .A(n702), .B(n701), .Z(c[235]) );
  AND U835 ( .A(b[0]), .B(a[109]), .Z(n705) );
  XNOR U836 ( .A(n706), .B(sreg[236]), .Z(n704) );
  XOR U837 ( .A(n705), .B(n704), .Z(c[236]) );
  AND U838 ( .A(b[0]), .B(a[110]), .Z(n708) );
  XNOR U839 ( .A(n709), .B(sreg[237]), .Z(n707) );
  XOR U840 ( .A(n708), .B(n707), .Z(c[237]) );
  AND U841 ( .A(b[0]), .B(a[111]), .Z(n711) );
  XNOR U842 ( .A(n712), .B(sreg[238]), .Z(n710) );
  XOR U843 ( .A(n711), .B(n710), .Z(c[238]) );
  AND U844 ( .A(b[0]), .B(a[112]), .Z(n714) );
  XNOR U845 ( .A(n715), .B(sreg[239]), .Z(n713) );
  XOR U846 ( .A(n714), .B(n713), .Z(c[239]) );
  AND U847 ( .A(b[0]), .B(a[113]), .Z(n717) );
  XNOR U848 ( .A(n718), .B(sreg[240]), .Z(n716) );
  XOR U849 ( .A(n717), .B(n716), .Z(c[240]) );
  AND U850 ( .A(b[0]), .B(a[114]), .Z(n720) );
  XNOR U851 ( .A(n721), .B(sreg[241]), .Z(n719) );
  XOR U852 ( .A(n720), .B(n719), .Z(c[241]) );
  AND U853 ( .A(b[0]), .B(a[115]), .Z(n723) );
  XNOR U854 ( .A(n724), .B(sreg[242]), .Z(n722) );
  XOR U855 ( .A(n723), .B(n722), .Z(c[242]) );
  AND U856 ( .A(b[0]), .B(a[116]), .Z(n726) );
  XNOR U857 ( .A(n727), .B(sreg[243]), .Z(n725) );
  XOR U858 ( .A(n726), .B(n725), .Z(c[243]) );
  AND U859 ( .A(b[0]), .B(a[117]), .Z(n729) );
  XNOR U860 ( .A(n730), .B(sreg[244]), .Z(n728) );
  XOR U861 ( .A(n729), .B(n728), .Z(c[244]) );
  AND U862 ( .A(b[0]), .B(a[118]), .Z(n732) );
  XNOR U863 ( .A(n733), .B(sreg[245]), .Z(n731) );
  XOR U864 ( .A(n732), .B(n731), .Z(c[245]) );
  AND U865 ( .A(b[0]), .B(a[119]), .Z(n735) );
  XNOR U866 ( .A(n736), .B(sreg[246]), .Z(n734) );
  XOR U867 ( .A(n735), .B(n734), .Z(c[246]) );
  AND U868 ( .A(b[0]), .B(a[120]), .Z(n738) );
  XNOR U869 ( .A(n739), .B(sreg[247]), .Z(n737) );
  XOR U870 ( .A(n738), .B(n737), .Z(c[247]) );
  AND U871 ( .A(b[0]), .B(a[121]), .Z(n741) );
  XNOR U872 ( .A(n742), .B(sreg[248]), .Z(n740) );
  XOR U873 ( .A(n741), .B(n740), .Z(c[248]) );
  AND U874 ( .A(b[0]), .B(a[122]), .Z(n744) );
  XNOR U875 ( .A(n745), .B(sreg[249]), .Z(n743) );
  XOR U876 ( .A(n744), .B(n743), .Z(c[249]) );
  AND U877 ( .A(b[0]), .B(a[123]), .Z(n747) );
  XNOR U878 ( .A(n748), .B(sreg[250]), .Z(n746) );
  XOR U879 ( .A(n747), .B(n746), .Z(c[250]) );
  AND U880 ( .A(b[0]), .B(a[124]), .Z(n750) );
  XNOR U881 ( .A(n751), .B(sreg[251]), .Z(n749) );
  XOR U882 ( .A(n750), .B(n749), .Z(c[251]) );
  AND U883 ( .A(b[0]), .B(a[125]), .Z(n753) );
  XNOR U884 ( .A(n754), .B(sreg[252]), .Z(n752) );
  XOR U885 ( .A(n753), .B(n752), .Z(c[252]) );
  AND U886 ( .A(b[0]), .B(a[126]), .Z(n756) );
  XNOR U887 ( .A(n757), .B(sreg[253]), .Z(n755) );
  XOR U888 ( .A(n756), .B(n755), .Z(c[253]) );
  NAND U889 ( .A(b[0]), .B(a[127]), .Z(n758) );
  XNOR U890 ( .A(sreg[254]), .B(n760), .Z(n759) );
  XNOR U891 ( .A(n758), .B(n759), .Z(c[254]) );
  NAND U892 ( .A(n759), .B(n758), .Z(n762) );
  NANDN U893 ( .A(sreg[254]), .B(n760), .Z(n761) );
  AND U894 ( .A(n762), .B(n761), .Z(c[255]) );
endmodule

