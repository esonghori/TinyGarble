
module mult_N1024_CC128 ( clk, rst, a, b, c );
  input [1023:0] a;
  input [7:0] b;
  output [2047:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593,
         n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
         n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
         n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
         n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
         n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
         n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
         n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665,
         n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
         n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
         n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
         n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
         n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713,
         n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737,
         n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
         n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
         n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
         n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
         n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857,
         n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
         n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
         n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
         n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
         n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
         n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929,
         n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
         n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
         n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
         n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
         n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
         n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
         n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
         n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
         n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
         n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
         n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
         n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
         n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097,
         n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
         n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
         n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
         n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
         n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
         n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
         n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
         n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169,
         n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
         n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
         n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
         n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201,
         n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
         n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217,
         n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
         n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
         n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
         n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
         n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
         n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
         n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273,
         n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
         n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
         n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
         n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
         n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313,
         n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
         n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
         n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337,
         n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345,
         n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
         n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361,
         n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
         n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377,
         n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385,
         n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393,
         n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
         n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409,
         n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417,
         n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
         n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433,
         n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
         n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449,
         n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
         n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
         n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
         n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
         n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489,
         n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
         n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505,
         n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
         n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521,
         n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529,
         n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537,
         n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
         n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553,
         n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
         n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
         n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577,
         n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
         n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593,
         n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601,
         n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609,
         n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
         n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625,
         n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633,
         n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641,
         n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649,
         n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
         n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
         n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673,
         n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681,
         n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
         n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697,
         n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705,
         n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
         n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721,
         n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
         n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737,
         n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745,
         n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753,
         n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
         n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769,
         n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777,
         n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785,
         n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793,
         n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
         n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809,
         n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817,
         n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825,
         n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
         n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841,
         n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849,
         n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857,
         n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865,
         n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
         n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881,
         n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889,
         n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897,
         n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
         n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913,
         n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921,
         n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
         n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937,
         n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
         n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953,
         n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961,
         n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
         n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
         n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985,
         n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993,
         n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
         n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009,
         n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017,
         n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025,
         n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033,
         n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
         n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049,
         n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057,
         n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065,
         n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
         n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081,
         n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089,
         n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097,
         n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105,
         n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113,
         n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121,
         n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129,
         n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137,
         n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
         n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153,
         n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
         n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169,
         n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177,
         n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185,
         n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
         n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201,
         n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209,
         n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217,
         n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225,
         n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233,
         n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241,
         n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249,
         n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257,
         n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265,
         n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273,
         n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281,
         n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289,
         n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297,
         n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305,
         n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313,
         n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321,
         n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
         n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
         n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345,
         n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353,
         n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361,
         n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369,
         n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377,
         n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385,
         n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393,
         n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
         n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409,
         n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417,
         n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425,
         n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433,
         n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441,
         n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449,
         n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457,
         n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465,
         n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
         n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481,
         n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489,
         n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497,
         n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
         n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513,
         n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521,
         n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529,
         n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537,
         n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545,
         n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553,
         n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561,
         n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569,
         n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577,
         n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585,
         n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593,
         n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601,
         n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609,
         n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617,
         n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625,
         n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633,
         n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641,
         n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
         n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657,
         n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665,
         n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
         n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681,
         n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
         n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697,
         n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705,
         n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713,
         n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
         n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729,
         n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
         n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745,
         n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
         n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761,
         n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
         n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777,
         n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785,
         n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
         n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801,
         n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
         n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
         n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825,
         n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
         n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841,
         n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849,
         n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857,
         n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865,
         n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873,
         n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
         n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889,
         n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897,
         n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905,
         n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913,
         n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921,
         n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929,
         n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
         n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945,
         n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
         n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961,
         n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969,
         n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977,
         n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985,
         n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993,
         n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001,
         n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009,
         n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017,
         n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025,
         n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
         n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041,
         n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
         n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
         n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065,
         n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073,
         n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081,
         n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089,
         n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097,
         n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105,
         n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113,
         n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121,
         n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129,
         n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137,
         n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145,
         n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153,
         n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161,
         n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169,
         n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177,
         n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185,
         n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193,
         n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201,
         n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209,
         n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217,
         n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225,
         n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233,
         n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241,
         n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249,
         n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257,
         n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265,
         n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273,
         n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281,
         n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289,
         n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
         n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305,
         n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313,
         n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321,
         n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329,
         n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337,
         n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345,
         n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353,
         n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361,
         n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369,
         n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377,
         n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385,
         n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
         n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401,
         n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409,
         n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417,
         n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425,
         n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433,
         n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441,
         n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449,
         n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457,
         n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
         n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473,
         n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481,
         n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
         n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497,
         n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505,
         n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513,
         n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521,
         n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529,
         n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537,
         n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545,
         n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553,
         n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561,
         n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569,
         n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577,
         n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
         n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593,
         n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
         n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609,
         n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617,
         n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625,
         n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633,
         n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641,
         n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649,
         n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657,
         n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665,
         n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
         n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681,
         n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689,
         n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697,
         n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705,
         n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713,
         n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721,
         n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
         n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737,
         n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
         n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753,
         n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761,
         n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769,
         n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777,
         n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785,
         n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793,
         n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801,
         n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809,
         n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
         n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825,
         n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833,
         n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841,
         n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849,
         n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857,
         n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865,
         n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873,
         n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881,
         n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
         n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897,
         n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905,
         n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913,
         n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921,
         n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929,
         n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937,
         n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945,
         n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
         n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
         n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969,
         n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977,
         n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985,
         n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993,
         n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001,
         n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009,
         n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
         n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
         n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
         n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041,
         n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049,
         n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057,
         n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065,
         n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073,
         n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081,
         n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
         n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097,
         n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105,
         n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113,
         n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121,
         n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129,
         n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137,
         n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145,
         n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153,
         n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
         n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
         n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177,
         n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185,
         n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193,
         n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201,
         n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209,
         n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217,
         n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225,
         n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
         n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241,
         n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249,
         n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257,
         n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265,
         n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273,
         n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281,
         n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289,
         n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297,
         n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
         n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313,
         n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
         n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329,
         n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337,
         n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345,
         n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353,
         n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361,
         n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369,
         n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
         n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385,
         n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393,
         n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401,
         n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409,
         n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417,
         n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425,
         n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433,
         n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441,
         n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
         n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457,
         n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465,
         n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473,
         n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481,
         n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489,
         n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497,
         n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505,
         n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513,
         n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
         n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529,
         n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537,
         n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545,
         n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553,
         n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561,
         n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569,
         n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577,
         n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585,
         n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593,
         n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601,
         n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609,
         n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617,
         n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625,
         n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633,
         n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641,
         n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649,
         n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657,
         n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665,
         n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673,
         n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681,
         n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689,
         n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697,
         n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705,
         n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713,
         n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721,
         n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729,
         n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737,
         n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745,
         n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753,
         n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761,
         n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769,
         n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777,
         n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785,
         n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793,
         n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801,
         n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809,
         n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817,
         n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825,
         n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833,
         n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841,
         n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849,
         n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857,
         n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865,
         n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873,
         n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881,
         n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889,
         n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897,
         n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905,
         n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913,
         n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921,
         n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929,
         n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937,
         n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945,
         n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953,
         n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961,
         n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969,
         n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977,
         n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985,
         n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993,
         n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001,
         n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009,
         n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017,
         n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025,
         n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033,
         n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041,
         n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049,
         n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057,
         n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065,
         n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073,
         n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081,
         n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089,
         n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097,
         n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105,
         n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113,
         n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121,
         n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129,
         n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137,
         n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145,
         n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153,
         n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161,
         n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169,
         n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177,
         n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185,
         n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193,
         n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201,
         n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209,
         n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217,
         n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225,
         n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233,
         n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241,
         n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249,
         n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257,
         n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265,
         n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273,
         n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281,
         n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289,
         n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297,
         n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305,
         n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313,
         n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321,
         n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329,
         n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337,
         n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345,
         n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353,
         n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361,
         n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369,
         n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377,
         n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385,
         n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393,
         n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401,
         n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409,
         n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417,
         n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425,
         n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433,
         n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441,
         n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449,
         n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457,
         n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465,
         n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473,
         n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481,
         n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489,
         n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497,
         n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505,
         n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513,
         n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521,
         n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529,
         n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537,
         n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545,
         n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553,
         n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561,
         n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569,
         n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577,
         n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585,
         n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593,
         n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601,
         n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609,
         n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617,
         n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625,
         n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633,
         n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641,
         n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649,
         n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657,
         n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665,
         n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673,
         n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681,
         n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689,
         n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697,
         n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705,
         n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713,
         n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721,
         n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729,
         n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737,
         n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745,
         n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753,
         n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761,
         n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769,
         n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777,
         n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785,
         n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793,
         n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801,
         n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809,
         n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817,
         n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825,
         n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833,
         n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841,
         n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849,
         n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857,
         n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865,
         n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873,
         n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881,
         n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889,
         n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897,
         n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905,
         n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913,
         n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921,
         n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929,
         n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937,
         n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945,
         n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953,
         n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961,
         n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969,
         n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977,
         n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985,
         n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993,
         n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001,
         n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009,
         n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017,
         n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025,
         n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033,
         n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041,
         n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049,
         n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057,
         n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065,
         n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073,
         n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081,
         n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089,
         n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097,
         n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105,
         n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113,
         n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121,
         n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129,
         n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137,
         n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145,
         n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153,
         n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161,
         n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169,
         n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177,
         n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185,
         n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193,
         n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201,
         n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209,
         n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217,
         n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225,
         n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233,
         n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241,
         n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249,
         n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257,
         n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265,
         n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273,
         n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281,
         n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289,
         n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297,
         n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305,
         n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313,
         n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321,
         n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329,
         n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337,
         n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345,
         n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353,
         n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361,
         n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369,
         n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377,
         n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385,
         n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393,
         n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401,
         n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409,
         n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417,
         n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425,
         n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433,
         n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441,
         n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449,
         n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457,
         n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465,
         n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473,
         n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481,
         n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489,
         n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497,
         n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505,
         n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513,
         n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521,
         n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529,
         n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537,
         n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545,
         n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553,
         n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561,
         n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569,
         n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577,
         n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585,
         n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593,
         n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601,
         n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609,
         n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617,
         n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625,
         n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633,
         n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641,
         n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649,
         n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657,
         n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665,
         n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673,
         n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681,
         n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689,
         n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697,
         n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705,
         n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713,
         n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721,
         n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729,
         n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737,
         n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745,
         n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753,
         n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761,
         n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769,
         n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777,
         n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785,
         n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793,
         n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801,
         n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809,
         n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817,
         n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825,
         n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833,
         n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841,
         n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849,
         n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857,
         n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865,
         n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873,
         n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881,
         n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889,
         n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897,
         n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905,
         n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913,
         n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921,
         n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929,
         n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937,
         n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945,
         n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953,
         n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961,
         n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969,
         n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977,
         n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985,
         n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993,
         n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001,
         n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009,
         n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017,
         n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025,
         n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033,
         n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041,
         n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049,
         n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057,
         n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065,
         n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073,
         n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081,
         n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089,
         n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097,
         n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105,
         n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113,
         n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121,
         n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129,
         n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137,
         n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145,
         n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153,
         n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161,
         n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169,
         n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177,
         n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185,
         n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193,
         n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201,
         n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209,
         n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217,
         n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225,
         n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233,
         n32234, n32235, n32236, n32237, n32238, n32239, n32240, n32241,
         n32242, n32243, n32244, n32245, n32246, n32247, n32248, n32249,
         n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257,
         n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265,
         n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273,
         n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281,
         n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289,
         n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297,
         n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305,
         n32306, n32307, n32308, n32309, n32310, n32311, n32312, n32313,
         n32314, n32315, n32316, n32317, n32318, n32319, n32320, n32321,
         n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329,
         n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337,
         n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345,
         n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353,
         n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361,
         n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369,
         n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377,
         n32378, n32379, n32380, n32381, n32382, n32383, n32384, n32385,
         n32386, n32387, n32388, n32389, n32390, n32391, n32392, n32393,
         n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401,
         n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409,
         n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417,
         n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425,
         n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433,
         n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441,
         n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449,
         n32450, n32451, n32452, n32453, n32454, n32455, n32456, n32457,
         n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465,
         n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473,
         n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481,
         n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489,
         n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497,
         n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505,
         n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513,
         n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521,
         n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529,
         n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537,
         n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545,
         n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553,
         n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561,
         n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569,
         n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577,
         n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585,
         n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593,
         n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601,
         n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609,
         n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617,
         n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625,
         n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633,
         n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641,
         n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649,
         n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657,
         n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665,
         n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673,
         n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681,
         n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689,
         n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697,
         n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705,
         n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713,
         n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721,
         n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729,
         n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737,
         n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745,
         n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753,
         n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761,
         n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769,
         n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777,
         n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785,
         n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793,
         n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801,
         n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809,
         n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817,
         n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825,
         n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833,
         n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841,
         n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849,
         n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857,
         n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865,
         n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873,
         n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881,
         n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889,
         n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897,
         n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905,
         n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913,
         n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921,
         n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929,
         n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937,
         n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945,
         n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953,
         n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961,
         n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969,
         n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977,
         n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985,
         n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993,
         n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001,
         n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009,
         n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017,
         n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025,
         n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033,
         n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041,
         n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049,
         n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057,
         n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065,
         n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073,
         n33074, n33075, n33076, n33077, n33078, n33079, n33080, n33081,
         n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089,
         n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097,
         n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105,
         n33106, n33107, n33108, n33109, n33110, n33111, n33112, n33113,
         n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121,
         n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129,
         n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137,
         n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145,
         n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153,
         n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161,
         n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169,
         n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177,
         n33178, n33179, n33180, n33181, n33182, n33183, n33184, n33185,
         n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193,
         n33194, n33195, n33196, n33197, n33198, n33199, n33200, n33201,
         n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209,
         n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217,
         n33218, n33219, n33220, n33221, n33222, n33223, n33224, n33225,
         n33226, n33227, n33228, n33229, n33230, n33231, n33232, n33233,
         n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241,
         n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249,
         n33250, n33251, n33252, n33253, n33254, n33255, n33256, n33257,
         n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265,
         n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273,
         n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281,
         n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289,
         n33290, n33291, n33292, n33293, n33294, n33295, n33296, n33297,
         n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305,
         n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313,
         n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321,
         n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329,
         n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337,
         n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345,
         n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33353,
         n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361,
         n33362, n33363, n33364, n33365, n33366, n33367, n33368, n33369,
         n33370, n33371, n33372, n33373, n33374, n33375, n33376, n33377,
         n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385,
         n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393,
         n33394, n33395, n33396, n33397, n33398, n33399, n33400, n33401,
         n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409,
         n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417,
         n33418, n33419, n33420, n33421, n33422, n33423, n33424, n33425,
         n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433,
         n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441,
         n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449,
         n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457,
         n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465,
         n33466, n33467, n33468, n33469, n33470, n33471, n33472, n33473,
         n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481,
         n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489,
         n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497,
         n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505,
         n33506, n33507, n33508, n33509, n33510, n33511, n33512, n33513,
         n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521,
         n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529,
         n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537,
         n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545,
         n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553,
         n33554, n33555, n33556, n33557, n33558, n33559, n33560, n33561,
         n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569,
         n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577,
         n33578, n33579, n33580, n33581, n33582, n33583, n33584, n33585,
         n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593,
         n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601,
         n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609,
         n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617,
         n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625,
         n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633,
         n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641,
         n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649,
         n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657,
         n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665,
         n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673,
         n33674, n33675, n33676, n33677, n33678, n33679, n33680, n33681,
         n33682, n33683, n33684, n33685, n33686, n33687, n33688, n33689,
         n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697,
         n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705,
         n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713,
         n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721,
         n33722, n33723, n33724, n33725, n33726, n33727, n33728, n33729,
         n33730, n33731, n33732, n33733, n33734, n33735, n33736, n33737,
         n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745,
         n33746, n33747, n33748, n33749, n33750, n33751, n33752, n33753,
         n33754, n33755, n33756, n33757, n33758, n33759, n33760, n33761,
         n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769,
         n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777,
         n33778, n33779, n33780, n33781, n33782, n33783, n33784, n33785,
         n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793,
         n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801,
         n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809,
         n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817,
         n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825,
         n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833,
         n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841,
         n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849,
         n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857,
         n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865,
         n33866, n33867, n33868, n33869, n33870, n33871, n33872, n33873,
         n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881,
         n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889,
         n33890, n33891, n33892, n33893, n33894, n33895, n33896, n33897,
         n33898, n33899, n33900, n33901, n33902, n33903, n33904, n33905,
         n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913,
         n33914, n33915, n33916, n33917, n33918, n33919, n33920, n33921,
         n33922, n33923, n33924, n33925, n33926, n33927, n33928, n33929,
         n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937,
         n33938, n33939, n33940, n33941, n33942, n33943, n33944, n33945,
         n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953,
         n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961,
         n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969,
         n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977,
         n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985,
         n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993,
         n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001,
         n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009,
         n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017,
         n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025,
         n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033,
         n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041,
         n34042, n34043, n34044, n34045, n34046, n34047, n34048, n34049,
         n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057,
         n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065,
         n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073,
         n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081,
         n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089,
         n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097,
         n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105,
         n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113,
         n34114, n34115, n34116, n34117, n34118, n34119, n34120, n34121,
         n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129,
         n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137,
         n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145,
         n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153,
         n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161,
         n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169,
         n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177,
         n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185,
         n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193,
         n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201,
         n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209,
         n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217,
         n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225,
         n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233,
         n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241,
         n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249,
         n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257,
         n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265,
         n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273,
         n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281,
         n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289,
         n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297,
         n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305,
         n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313,
         n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321,
         n34322, n34323, n34324, n34325, n34326, n34327, n34328, n34329,
         n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337,
         n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345,
         n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353,
         n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361,
         n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369,
         n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377,
         n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385,
         n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393,
         n34394, n34395, n34396, n34397, n34398, n34399, n34400, n34401,
         n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409,
         n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417,
         n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425,
         n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433,
         n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441,
         n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449,
         n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457,
         n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465,
         n34466, n34467, n34468, n34469, n34470, n34471, n34472, n34473,
         n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481,
         n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489,
         n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497,
         n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505,
         n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513,
         n34514, n34515, n34516, n34517, n34518, n34519, n34520, n34521,
         n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529,
         n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537,
         n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545,
         n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553,
         n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561,
         n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569,
         n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577,
         n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585,
         n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593,
         n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601,
         n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609,
         n34610, n34611, n34612, n34613, n34614, n34615, n34616, n34617,
         n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625,
         n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633,
         n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641,
         n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649,
         n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657,
         n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665,
         n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673,
         n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681,
         n34682, n34683, n34684, n34685, n34686, n34687, n34688, n34689,
         n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697,
         n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705,
         n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713,
         n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721,
         n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729,
         n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737,
         n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745,
         n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753,
         n34754, n34755, n34756, n34757, n34758, n34759, n34760, n34761,
         n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769,
         n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777,
         n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785,
         n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793,
         n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801,
         n34802, n34803, n34804, n34805, n34806, n34807, n34808, n34809,
         n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817,
         n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825,
         n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833,
         n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841,
         n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849,
         n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857,
         n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865,
         n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873,
         n34874, n34875, n34876, n34877, n34878, n34879, n34880, n34881,
         n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889,
         n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897,
         n34898, n34899, n34900, n34901, n34902, n34903, n34904, n34905,
         n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913,
         n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921,
         n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929,
         n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937,
         n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945,
         n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953,
         n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961,
         n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969,
         n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977,
         n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985,
         n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993,
         n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001,
         n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009,
         n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017,
         n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025,
         n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033,
         n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041,
         n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049,
         n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057,
         n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065,
         n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073,
         n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081,
         n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089,
         n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097,
         n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105,
         n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113,
         n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121,
         n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129,
         n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137,
         n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145,
         n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153,
         n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161,
         n35162, n35163, n35164, n35165, n35166, n35167, n35168, n35169,
         n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177,
         n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185,
         n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193,
         n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201,
         n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209,
         n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217,
         n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225,
         n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233,
         n35234, n35235, n35236, n35237, n35238, n35239, n35240, n35241,
         n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249,
         n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257,
         n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265,
         n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273,
         n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281,
         n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289,
         n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297,
         n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305,
         n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313,
         n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321,
         n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329,
         n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337,
         n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345,
         n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353,
         n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361,
         n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369,
         n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377,
         n35378, n35379, n35380, n35381, n35382, n35383, n35384, n35385,
         n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393,
         n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401,
         n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35409,
         n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417,
         n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425,
         n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433,
         n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441,
         n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449,
         n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457,
         n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465,
         n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473,
         n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481,
         n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489,
         n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497,
         n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505,
         n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513,
         n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521,
         n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529,
         n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537,
         n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545,
         n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553,
         n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561,
         n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569,
         n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577,
         n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585,
         n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593,
         n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601,
         n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609,
         n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617,
         n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625,
         n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633,
         n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641,
         n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649,
         n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657,
         n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665,
         n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673,
         n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681,
         n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689,
         n35690, n35691, n35692, n35693, n35694, n35695, n35696, n35697,
         n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705,
         n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713,
         n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721,
         n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729,
         n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737,
         n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745,
         n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753,
         n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761,
         n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769,
         n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777,
         n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785,
         n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793,
         n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801,
         n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809,
         n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817,
         n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825,
         n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833,
         n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841,
         n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849,
         n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857,
         n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865,
         n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873,
         n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881,
         n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889,
         n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897,
         n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905,
         n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913,
         n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921,
         n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929,
         n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937,
         n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945,
         n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953,
         n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961,
         n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969,
         n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977,
         n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985,
         n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993,
         n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001,
         n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009,
         n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017,
         n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025,
         n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033,
         n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041,
         n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049,
         n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057,
         n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065,
         n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073,
         n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081,
         n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089,
         n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097,
         n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105,
         n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113,
         n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121,
         n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129,
         n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137,
         n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145,
         n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153,
         n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161,
         n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169,
         n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177,
         n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185,
         n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193,
         n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201,
         n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209,
         n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217,
         n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225,
         n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233,
         n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241,
         n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249,
         n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257,
         n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265,
         n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273,
         n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281,
         n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289,
         n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297,
         n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305,
         n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313,
         n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321,
         n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329,
         n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337,
         n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345,
         n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353,
         n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361,
         n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369,
         n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377,
         n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385,
         n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393,
         n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401,
         n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409,
         n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417,
         n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425,
         n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433,
         n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441,
         n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449,
         n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457,
         n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465,
         n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473,
         n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481,
         n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489,
         n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497,
         n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505,
         n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513,
         n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521,
         n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529,
         n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537,
         n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545,
         n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553,
         n36554, n36555, n36556, n36557, n36558, n36559, n36560, n36561,
         n36562, n36563, n36564, n36565, n36566, n36567, n36568, n36569,
         n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577,
         n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585,
         n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593,
         n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601,
         n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609,
         n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617,
         n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625,
         n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633,
         n36634, n36635, n36636, n36637, n36638, n36639, n36640, n36641,
         n36642, n36643, n36644, n36645, n36646, n36647, n36648, n36649,
         n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657,
         n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665,
         n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673,
         n36674, n36675, n36676, n36677, n36678, n36679, n36680, n36681,
         n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689,
         n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697,
         n36698, n36699, n36700, n36701, n36702, n36703, n36704, n36705,
         n36706, n36707, n36708, n36709, n36710, n36711, n36712, n36713,
         n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721,
         n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729,
         n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737,
         n36738, n36739, n36740, n36741, n36742, n36743, n36744, n36745,
         n36746, n36747, n36748, n36749, n36750, n36751, n36752, n36753,
         n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761,
         n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769,
         n36770, n36771, n36772, n36773, n36774, n36775, n36776, n36777,
         n36778, n36779, n36780, n36781, n36782, n36783, n36784, n36785,
         n36786, n36787, n36788, n36789, n36790, n36791, n36792, n36793,
         n36794, n36795, n36796, n36797, n36798, n36799, n36800, n36801,
         n36802, n36803, n36804, n36805, n36806, n36807, n36808, n36809,
         n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817,
         n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825,
         n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833,
         n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841,
         n36842, n36843, n36844, n36845, n36846, n36847, n36848, n36849,
         n36850, n36851, n36852, n36853, n36854, n36855, n36856, n36857,
         n36858, n36859, n36860, n36861, n36862, n36863, n36864, n36865,
         n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873,
         n36874, n36875, n36876, n36877, n36878, n36879, n36880, n36881,
         n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889,
         n36890, n36891, n36892, n36893, n36894, n36895, n36896, n36897,
         n36898, n36899, n36900, n36901, n36902, n36903, n36904, n36905,
         n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913,
         n36914, n36915, n36916, n36917, n36918, n36919, n36920, n36921,
         n36922, n36923, n36924, n36925, n36926, n36927, n36928, n36929,
         n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937,
         n36938, n36939, n36940, n36941, n36942, n36943, n36944, n36945,
         n36946, n36947, n36948, n36949, n36950, n36951, n36952, n36953,
         n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961,
         n36962, n36963, n36964, n36965, n36966, n36967, n36968, n36969,
         n36970, n36971, n36972, n36973, n36974, n36975, n36976, n36977,
         n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985,
         n36986, n36987, n36988, n36989, n36990, n36991, n36992, n36993,
         n36994, n36995, n36996, n36997, n36998, n36999, n37000, n37001,
         n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009,
         n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017,
         n37018, n37019, n37020, n37021, n37022, n37023, n37024, n37025,
         n37026, n37027, n37028, n37029, n37030, n37031, n37032, n37033,
         n37034, n37035, n37036, n37037, n37038, n37039, n37040, n37041,
         n37042, n37043, n37044, n37045, n37046, n37047, n37048, n37049,
         n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057,
         n37058, n37059, n37060, n37061, n37062, n37063, n37064, n37065,
         n37066, n37067, n37068, n37069, n37070, n37071, n37072, n37073,
         n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081,
         n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089,
         n37090, n37091, n37092, n37093, n37094, n37095, n37096, n37097,
         n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105,
         n37106, n37107, n37108, n37109, n37110, n37111, n37112, n37113,
         n37114, n37115, n37116, n37117, n37118, n37119, n37120, n37121,
         n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129,
         n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137,
         n37138, n37139, n37140, n37141, n37142, n37143, n37144, n37145,
         n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153,
         n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161,
         n37162, n37163, n37164, n37165, n37166, n37167, n37168, n37169,
         n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177,
         n37178, n37179, n37180, n37181, n37182, n37183, n37184, n37185,
         n37186, n37187, n37188, n37189, n37190, n37191, n37192, n37193,
         n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201,
         n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209,
         n37210, n37211, n37212, n37213, n37214, n37215, n37216, n37217,
         n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225,
         n37226, n37227, n37228, n37229, n37230, n37231, n37232, n37233,
         n37234, n37235, n37236, n37237, n37238, n37239, n37240, n37241,
         n37242, n37243, n37244, n37245, n37246, n37247, n37248, n37249,
         n37250, n37251, n37252, n37253, n37254, n37255, n37256, n37257,
         n37258, n37259, n37260, n37261, n37262, n37263, n37264, n37265,
         n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273,
         n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281,
         n37282, n37283, n37284, n37285, n37286, n37287, n37288, n37289,
         n37290, n37291, n37292, n37293, n37294, n37295, n37296, n37297,
         n37298, n37299, n37300, n37301, n37302, n37303, n37304, n37305,
         n37306, n37307, n37308, n37309, n37310, n37311, n37312, n37313,
         n37314, n37315, n37316, n37317, n37318, n37319, n37320, n37321,
         n37322, n37323, n37324, n37325, n37326, n37327, n37328, n37329,
         n37330, n37331, n37332, n37333, n37334, n37335, n37336, n37337,
         n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345,
         n37346, n37347, n37348, n37349, n37350, n37351, n37352, n37353,
         n37354, n37355, n37356, n37357, n37358, n37359, n37360, n37361,
         n37362, n37363, n37364, n37365, n37366, n37367, n37368, n37369,
         n37370, n37371, n37372, n37373, n37374, n37375, n37376, n37377,
         n37378, n37379, n37380, n37381, n37382, n37383, n37384, n37385,
         n37386, n37387, n37388, n37389, n37390, n37391, n37392, n37393,
         n37394, n37395, n37396, n37397, n37398, n37399, n37400, n37401,
         n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409,
         n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417,
         n37418, n37419, n37420, n37421, n37422, n37423, n37424, n37425,
         n37426, n37427, n37428, n37429, n37430, n37431, n37432, n37433,
         n37434, n37435, n37436, n37437, n37438, n37439, n37440, n37441,
         n37442, n37443, n37444, n37445, n37446, n37447, n37448, n37449,
         n37450, n37451, n37452, n37453, n37454, n37455, n37456, n37457,
         n37458, n37459, n37460, n37461, n37462, n37463, n37464, n37465,
         n37466, n37467, n37468, n37469, n37470, n37471, n37472, n37473,
         n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481,
         n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489,
         n37490, n37491, n37492, n37493, n37494, n37495, n37496, n37497,
         n37498, n37499, n37500, n37501, n37502, n37503, n37504, n37505,
         n37506, n37507, n37508, n37509, n37510, n37511, n37512, n37513,
         n37514, n37515, n37516, n37517, n37518, n37519, n37520, n37521,
         n37522, n37523, n37524, n37525, n37526, n37527, n37528, n37529,
         n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537,
         n37538, n37539, n37540, n37541, n37542, n37543, n37544, n37545,
         n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553,
         n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561,
         n37562, n37563, n37564, n37565, n37566, n37567, n37568, n37569,
         n37570, n37571, n37572, n37573, n37574, n37575, n37576, n37577,
         n37578, n37579, n37580, n37581, n37582, n37583, n37584, n37585,
         n37586, n37587, n37588, n37589, n37590, n37591, n37592, n37593,
         n37594, n37595, n37596, n37597, n37598, n37599, n37600, n37601,
         n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609,
         n37610, n37611, n37612, n37613, n37614, n37615, n37616, n37617,
         n37618, n37619, n37620, n37621, n37622, n37623, n37624, n37625,
         n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633,
         n37634, n37635, n37636, n37637, n37638, n37639, n37640, n37641,
         n37642, n37643, n37644, n37645, n37646, n37647, n37648, n37649,
         n37650, n37651, n37652, n37653, n37654, n37655, n37656, n37657,
         n37658, n37659, n37660, n37661, n37662, n37663, n37664, n37665,
         n37666, n37667, n37668, n37669, n37670, n37671, n37672, n37673,
         n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681,
         n37682, n37683, n37684, n37685, n37686, n37687, n37688, n37689,
         n37690, n37691, n37692, n37693, n37694, n37695, n37696, n37697,
         n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705,
         n37706, n37707, n37708, n37709, n37710, n37711, n37712, n37713,
         n37714, n37715, n37716, n37717, n37718, n37719, n37720, n37721,
         n37722, n37723, n37724, n37725, n37726, n37727, n37728, n37729,
         n37730, n37731, n37732, n37733, n37734, n37735, n37736, n37737,
         n37738, n37739, n37740, n37741, n37742, n37743, n37744, n37745,
         n37746, n37747, n37748, n37749, n37750, n37751, n37752, n37753,
         n37754, n37755, n37756, n37757, n37758, n37759, n37760, n37761,
         n37762, n37763, n37764, n37765, n37766, n37767, n37768, n37769,
         n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777,
         n37778, n37779, n37780, n37781, n37782, n37783, n37784, n37785,
         n37786, n37787, n37788, n37789, n37790, n37791, n37792, n37793,
         n37794, n37795, n37796, n37797, n37798, n37799, n37800, n37801,
         n37802, n37803, n37804, n37805, n37806, n37807, n37808, n37809,
         n37810, n37811, n37812, n37813, n37814, n37815, n37816, n37817,
         n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825,
         n37826, n37827, n37828, n37829, n37830, n37831, n37832, n37833,
         n37834, n37835, n37836, n37837, n37838, n37839, n37840, n37841,
         n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849,
         n37850, n37851, n37852, n37853, n37854, n37855, n37856, n37857,
         n37858, n37859, n37860, n37861, n37862, n37863, n37864, n37865,
         n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873,
         n37874, n37875, n37876, n37877, n37878, n37879, n37880, n37881,
         n37882, n37883, n37884, n37885, n37886, n37887, n37888, n37889,
         n37890, n37891, n37892, n37893, n37894, n37895, n37896, n37897,
         n37898, n37899, n37900, n37901, n37902, n37903, n37904, n37905,
         n37906, n37907, n37908, n37909, n37910, n37911, n37912, n37913,
         n37914, n37915, n37916, n37917, n37918, n37919, n37920, n37921,
         n37922, n37923, n37924, n37925, n37926, n37927, n37928, n37929,
         n37930, n37931, n37932, n37933, n37934, n37935, n37936, n37937,
         n37938, n37939, n37940, n37941, n37942, n37943, n37944, n37945,
         n37946, n37947, n37948, n37949, n37950, n37951, n37952, n37953,
         n37954, n37955, n37956, n37957, n37958, n37959, n37960, n37961,
         n37962, n37963, n37964, n37965, n37966, n37967, n37968, n37969,
         n37970, n37971, n37972, n37973, n37974, n37975, n37976, n37977,
         n37978, n37979, n37980, n37981, n37982, n37983, n37984, n37985,
         n37986, n37987, n37988, n37989, n37990, n37991, n37992, n37993,
         n37994, n37995, n37996, n37997, n37998, n37999, n38000, n38001,
         n38002, n38003, n38004, n38005, n38006, n38007, n38008, n38009,
         n38010, n38011, n38012, n38013, n38014, n38015, n38016, n38017,
         n38018, n38019, n38020, n38021, n38022, n38023, n38024, n38025,
         n38026, n38027, n38028, n38029, n38030, n38031, n38032, n38033,
         n38034, n38035, n38036, n38037, n38038, n38039, n38040, n38041,
         n38042, n38043, n38044, n38045, n38046, n38047, n38048, n38049,
         n38050, n38051, n38052, n38053, n38054, n38055, n38056, n38057,
         n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065,
         n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073,
         n38074, n38075, n38076, n38077, n38078, n38079, n38080, n38081,
         n38082, n38083, n38084, n38085, n38086, n38087, n38088, n38089,
         n38090, n38091, n38092, n38093, n38094, n38095, n38096, n38097,
         n38098, n38099, n38100, n38101, n38102, n38103, n38104, n38105,
         n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113,
         n38114, n38115, n38116, n38117, n38118, n38119, n38120, n38121,
         n38122, n38123, n38124, n38125, n38126, n38127, n38128, n38129,
         n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137,
         n38138, n38139, n38140, n38141, n38142, n38143, n38144, n38145,
         n38146, n38147, n38148, n38149, n38150, n38151, n38152, n38153,
         n38154, n38155, n38156, n38157, n38158, n38159, n38160, n38161,
         n38162, n38163, n38164, n38165, n38166, n38167, n38168, n38169,
         n38170, n38171, n38172, n38173, n38174, n38175, n38176, n38177,
         n38178, n38179, n38180, n38181, n38182, n38183, n38184, n38185,
         n38186, n38187, n38188, n38189, n38190, n38191, n38192, n38193,
         n38194, n38195, n38196, n38197, n38198, n38199, n38200, n38201,
         n38202, n38203, n38204, n38205, n38206, n38207, n38208, n38209,
         n38210, n38211, n38212, n38213, n38214, n38215, n38216, n38217,
         n38218, n38219, n38220, n38221, n38222, n38223, n38224, n38225,
         n38226, n38227, n38228, n38229, n38230, n38231, n38232, n38233,
         n38234, n38235, n38236, n38237, n38238, n38239, n38240, n38241,
         n38242, n38243, n38244, n38245, n38246, n38247, n38248, n38249,
         n38250, n38251, n38252, n38253, n38254, n38255, n38256, n38257,
         n38258, n38259, n38260, n38261, n38262, n38263, n38264, n38265,
         n38266, n38267, n38268, n38269, n38270, n38271, n38272, n38273,
         n38274, n38275, n38276, n38277, n38278, n38279, n38280, n38281,
         n38282, n38283, n38284, n38285, n38286, n38287, n38288, n38289,
         n38290, n38291, n38292, n38293, n38294, n38295, n38296, n38297,
         n38298, n38299, n38300, n38301, n38302, n38303, n38304, n38305,
         n38306, n38307, n38308, n38309, n38310, n38311, n38312, n38313,
         n38314, n38315, n38316, n38317, n38318, n38319, n38320, n38321,
         n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329,
         n38330, n38331, n38332, n38333, n38334, n38335, n38336, n38337,
         n38338, n38339, n38340, n38341, n38342, n38343, n38344, n38345,
         n38346, n38347, n38348, n38349, n38350, n38351, n38352, n38353,
         n38354, n38355, n38356, n38357, n38358, n38359, n38360, n38361,
         n38362, n38363, n38364, n38365, n38366, n38367, n38368, n38369,
         n38370, n38371, n38372, n38373, n38374, n38375, n38376, n38377,
         n38378, n38379, n38380, n38381, n38382, n38383, n38384, n38385,
         n38386, n38387, n38388, n38389, n38390, n38391, n38392, n38393,
         n38394, n38395, n38396, n38397, n38398, n38399, n38400, n38401,
         n38402, n38403, n38404, n38405, n38406, n38407, n38408, n38409,
         n38410, n38411, n38412, n38413, n38414, n38415, n38416, n38417,
         n38418, n38419, n38420, n38421, n38422, n38423, n38424, n38425,
         n38426, n38427, n38428, n38429, n38430, n38431, n38432, n38433,
         n38434, n38435, n38436, n38437, n38438, n38439, n38440, n38441,
         n38442, n38443, n38444, n38445, n38446, n38447, n38448, n38449,
         n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457,
         n38458, n38459, n38460, n38461, n38462, n38463, n38464, n38465,
         n38466, n38467, n38468, n38469, n38470, n38471, n38472, n38473,
         n38474, n38475, n38476, n38477, n38478, n38479, n38480, n38481,
         n38482, n38483, n38484, n38485, n38486, n38487, n38488, n38489,
         n38490, n38491, n38492, n38493, n38494, n38495, n38496, n38497,
         n38498, n38499, n38500, n38501, n38502, n38503, n38504, n38505,
         n38506, n38507, n38508, n38509, n38510, n38511, n38512, n38513,
         n38514, n38515, n38516, n38517, n38518, n38519, n38520, n38521,
         n38522, n38523, n38524, n38525, n38526, n38527, n38528, n38529,
         n38530, n38531, n38532, n38533, n38534, n38535, n38536, n38537,
         n38538, n38539, n38540, n38541, n38542, n38543, n38544, n38545,
         n38546, n38547, n38548, n38549, n38550, n38551, n38552, n38553,
         n38554, n38555, n38556, n38557, n38558, n38559, n38560, n38561,
         n38562, n38563, n38564, n38565, n38566, n38567, n38568, n38569,
         n38570, n38571, n38572, n38573, n38574, n38575, n38576, n38577,
         n38578, n38579, n38580, n38581, n38582, n38583, n38584, n38585,
         n38586, n38587, n38588, n38589, n38590, n38591, n38592, n38593,
         n38594, n38595, n38596, n38597, n38598, n38599, n38600, n38601,
         n38602, n38603, n38604, n38605, n38606, n38607, n38608, n38609,
         n38610, n38611, n38612, n38613, n38614, n38615, n38616, n38617,
         n38618, n38619, n38620, n38621, n38622, n38623, n38624, n38625,
         n38626, n38627, n38628, n38629, n38630, n38631, n38632, n38633,
         n38634, n38635, n38636, n38637, n38638, n38639, n38640, n38641,
         n38642, n38643, n38644, n38645, n38646, n38647, n38648, n38649,
         n38650, n38651, n38652, n38653, n38654, n38655, n38656, n38657,
         n38658, n38659, n38660, n38661, n38662, n38663, n38664, n38665,
         n38666, n38667, n38668, n38669, n38670, n38671, n38672, n38673,
         n38674, n38675, n38676, n38677, n38678, n38679, n38680, n38681,
         n38682, n38683, n38684, n38685, n38686, n38687, n38688, n38689,
         n38690, n38691, n38692, n38693, n38694, n38695, n38696, n38697,
         n38698, n38699, n38700, n38701, n38702, n38703, n38704, n38705,
         n38706, n38707, n38708, n38709, n38710, n38711, n38712, n38713,
         n38714, n38715, n38716, n38717, n38718, n38719, n38720, n38721,
         n38722, n38723, n38724, n38725, n38726, n38727, n38728, n38729,
         n38730, n38731, n38732, n38733, n38734, n38735, n38736, n38737,
         n38738, n38739, n38740, n38741, n38742, n38743, n38744, n38745,
         n38746, n38747, n38748, n38749, n38750, n38751, n38752, n38753,
         n38754, n38755, n38756, n38757, n38758, n38759, n38760, n38761,
         n38762, n38763, n38764, n38765, n38766, n38767, n38768, n38769,
         n38770, n38771, n38772, n38773, n38774, n38775, n38776, n38777,
         n38778, n38779, n38780, n38781, n38782, n38783, n38784, n38785,
         n38786, n38787, n38788, n38789, n38790, n38791, n38792, n38793,
         n38794, n38795, n38796, n38797, n38798, n38799, n38800, n38801,
         n38802, n38803, n38804, n38805, n38806, n38807, n38808, n38809,
         n38810, n38811, n38812, n38813, n38814, n38815, n38816, n38817,
         n38818, n38819, n38820, n38821, n38822, n38823, n38824, n38825,
         n38826, n38827, n38828, n38829, n38830, n38831, n38832, n38833,
         n38834, n38835, n38836, n38837, n38838, n38839, n38840, n38841,
         n38842, n38843, n38844, n38845, n38846, n38847, n38848, n38849,
         n38850, n38851, n38852, n38853, n38854, n38855, n38856, n38857,
         n38858, n38859, n38860, n38861, n38862, n38863, n38864, n38865,
         n38866, n38867, n38868, n38869, n38870, n38871, n38872, n38873,
         n38874, n38875, n38876, n38877, n38878, n38879, n38880, n38881,
         n38882, n38883, n38884, n38885, n38886, n38887, n38888, n38889,
         n38890, n38891, n38892, n38893, n38894, n38895, n38896, n38897,
         n38898, n38899, n38900, n38901, n38902, n38903, n38904, n38905,
         n38906, n38907, n38908, n38909, n38910, n38911, n38912, n38913,
         n38914, n38915, n38916, n38917, n38918, n38919, n38920, n38921,
         n38922, n38923, n38924, n38925, n38926, n38927, n38928, n38929,
         n38930, n38931, n38932, n38933, n38934, n38935, n38936, n38937,
         n38938, n38939, n38940, n38941, n38942, n38943, n38944, n38945,
         n38946, n38947, n38948, n38949, n38950, n38951, n38952, n38953,
         n38954, n38955, n38956, n38957, n38958, n38959, n38960, n38961,
         n38962, n38963, n38964, n38965, n38966, n38967, n38968, n38969,
         n38970, n38971, n38972, n38973, n38974, n38975, n38976, n38977,
         n38978, n38979, n38980, n38981, n38982, n38983, n38984, n38985,
         n38986, n38987, n38988, n38989, n38990, n38991, n38992, n38993,
         n38994, n38995, n38996, n38997, n38998, n38999, n39000, n39001,
         n39002, n39003, n39004, n39005, n39006, n39007, n39008, n39009,
         n39010, n39011, n39012, n39013, n39014, n39015, n39016, n39017,
         n39018, n39019, n39020, n39021, n39022, n39023, n39024, n39025,
         n39026, n39027, n39028, n39029, n39030, n39031, n39032, n39033,
         n39034, n39035, n39036, n39037, n39038, n39039, n39040, n39041,
         n39042, n39043, n39044, n39045, n39046, n39047, n39048, n39049,
         n39050, n39051, n39052, n39053, n39054, n39055, n39056, n39057,
         n39058, n39059, n39060, n39061, n39062, n39063, n39064, n39065,
         n39066, n39067, n39068, n39069, n39070, n39071, n39072, n39073,
         n39074, n39075, n39076, n39077, n39078, n39079, n39080, n39081,
         n39082, n39083, n39084, n39085, n39086, n39087, n39088, n39089,
         n39090, n39091, n39092, n39093, n39094, n39095, n39096, n39097,
         n39098, n39099, n39100, n39101, n39102, n39103, n39104, n39105,
         n39106, n39107, n39108, n39109, n39110, n39111, n39112, n39113,
         n39114, n39115, n39116, n39117, n39118, n39119, n39120, n39121,
         n39122, n39123, n39124, n39125, n39126, n39127, n39128, n39129,
         n39130, n39131, n39132, n39133, n39134, n39135, n39136, n39137,
         n39138, n39139, n39140, n39141, n39142, n39143, n39144, n39145,
         n39146, n39147, n39148, n39149, n39150, n39151, n39152, n39153,
         n39154, n39155, n39156, n39157, n39158, n39159, n39160, n39161,
         n39162, n39163, n39164, n39165, n39166, n39167, n39168, n39169,
         n39170, n39171, n39172, n39173, n39174, n39175, n39176, n39177,
         n39178, n39179, n39180, n39181, n39182, n39183, n39184, n39185,
         n39186, n39187, n39188, n39189, n39190, n39191, n39192, n39193,
         n39194, n39195, n39196, n39197, n39198, n39199, n39200, n39201,
         n39202, n39203, n39204, n39205, n39206, n39207, n39208, n39209,
         n39210, n39211, n39212, n39213, n39214, n39215, n39216, n39217,
         n39218, n39219, n39220, n39221, n39222, n39223, n39224, n39225,
         n39226, n39227, n39228, n39229, n39230, n39231, n39232, n39233,
         n39234, n39235, n39236, n39237, n39238, n39239, n39240, n39241,
         n39242, n39243, n39244, n39245, n39246, n39247, n39248, n39249,
         n39250, n39251, n39252, n39253, n39254, n39255, n39256, n39257,
         n39258, n39259, n39260, n39261, n39262, n39263, n39264, n39265,
         n39266, n39267, n39268, n39269, n39270, n39271, n39272, n39273,
         n39274, n39275, n39276, n39277, n39278, n39279, n39280, n39281,
         n39282, n39283, n39284, n39285, n39286, n39287, n39288, n39289,
         n39290, n39291, n39292, n39293, n39294, n39295, n39296, n39297,
         n39298, n39299, n39300, n39301, n39302, n39303, n39304, n39305,
         n39306, n39307, n39308, n39309, n39310, n39311, n39312, n39313,
         n39314, n39315, n39316, n39317, n39318, n39319, n39320, n39321,
         n39322, n39323, n39324, n39325, n39326, n39327, n39328, n39329,
         n39330, n39331, n39332, n39333, n39334, n39335, n39336, n39337,
         n39338, n39339, n39340, n39341, n39342, n39343, n39344, n39345,
         n39346, n39347, n39348, n39349, n39350, n39351, n39352, n39353,
         n39354, n39355, n39356, n39357, n39358, n39359, n39360, n39361,
         n39362, n39363, n39364, n39365, n39366, n39367, n39368, n39369,
         n39370, n39371, n39372, n39373, n39374, n39375, n39376, n39377,
         n39378, n39379, n39380, n39381, n39382, n39383, n39384, n39385,
         n39386, n39387, n39388, n39389, n39390, n39391, n39392, n39393,
         n39394, n39395, n39396, n39397, n39398, n39399, n39400, n39401,
         n39402, n39403, n39404, n39405, n39406, n39407, n39408, n39409,
         n39410, n39411, n39412, n39413, n39414, n39415, n39416, n39417,
         n39418, n39419, n39420, n39421, n39422, n39423, n39424, n39425,
         n39426, n39427, n39428, n39429, n39430, n39431, n39432, n39433,
         n39434, n39435, n39436, n39437, n39438, n39439, n39440, n39441,
         n39442, n39443, n39444, n39445, n39446, n39447, n39448, n39449,
         n39450, n39451, n39452, n39453, n39454, n39455, n39456, n39457,
         n39458, n39459, n39460, n39461, n39462, n39463, n39464, n39465,
         n39466, n39467, n39468, n39469, n39470, n39471, n39472, n39473,
         n39474, n39475, n39476, n39477, n39478, n39479, n39480, n39481,
         n39482, n39483, n39484, n39485, n39486, n39487, n39488, n39489,
         n39490, n39491, n39492, n39493, n39494, n39495, n39496, n39497,
         n39498, n39499, n39500, n39501, n39502, n39503, n39504, n39505,
         n39506, n39507, n39508, n39509, n39510, n39511, n39512, n39513,
         n39514, n39515, n39516, n39517, n39518, n39519, n39520, n39521,
         n39522, n39523, n39524, n39525, n39526, n39527, n39528, n39529,
         n39530, n39531, n39532, n39533, n39534, n39535, n39536, n39537,
         n39538, n39539, n39540, n39541, n39542, n39543, n39544, n39545,
         n39546, n39547, n39548, n39549, n39550, n39551, n39552, n39553,
         n39554, n39555, n39556, n39557, n39558, n39559, n39560, n39561,
         n39562, n39563, n39564, n39565, n39566, n39567, n39568, n39569,
         n39570, n39571, n39572, n39573, n39574, n39575, n39576, n39577,
         n39578, n39579, n39580, n39581, n39582, n39583, n39584, n39585,
         n39586, n39587, n39588, n39589, n39590, n39591, n39592, n39593,
         n39594, n39595, n39596, n39597, n39598, n39599, n39600, n39601,
         n39602, n39603, n39604, n39605, n39606, n39607, n39608, n39609,
         n39610, n39611, n39612, n39613, n39614, n39615, n39616, n39617,
         n39618, n39619, n39620, n39621, n39622, n39623, n39624, n39625,
         n39626, n39627, n39628, n39629, n39630, n39631, n39632, n39633,
         n39634, n39635, n39636, n39637, n39638, n39639, n39640, n39641,
         n39642, n39643, n39644, n39645, n39646, n39647, n39648, n39649,
         n39650, n39651, n39652, n39653, n39654, n39655, n39656, n39657,
         n39658, n39659, n39660, n39661, n39662, n39663, n39664, n39665,
         n39666, n39667, n39668, n39669, n39670, n39671, n39672, n39673,
         n39674, n39675, n39676, n39677, n39678, n39679, n39680, n39681,
         n39682, n39683, n39684, n39685, n39686, n39687, n39688, n39689,
         n39690, n39691, n39692, n39693, n39694, n39695, n39696, n39697,
         n39698, n39699, n39700, n39701, n39702, n39703, n39704, n39705,
         n39706, n39707, n39708, n39709, n39710, n39711, n39712, n39713,
         n39714, n39715, n39716, n39717, n39718, n39719, n39720, n39721,
         n39722, n39723, n39724, n39725, n39726, n39727, n39728, n39729,
         n39730, n39731, n39732, n39733, n39734, n39735, n39736, n39737,
         n39738, n39739, n39740, n39741, n39742, n39743, n39744, n39745,
         n39746, n39747, n39748, n39749, n39750, n39751, n39752, n39753,
         n39754, n39755, n39756, n39757, n39758, n39759, n39760, n39761,
         n39762, n39763, n39764, n39765, n39766, n39767, n39768, n39769,
         n39770, n39771, n39772, n39773, n39774, n39775, n39776, n39777,
         n39778, n39779, n39780, n39781, n39782, n39783, n39784, n39785,
         n39786, n39787, n39788, n39789, n39790, n39791, n39792, n39793,
         n39794, n39795, n39796, n39797, n39798, n39799, n39800, n39801,
         n39802, n39803, n39804, n39805, n39806, n39807, n39808, n39809,
         n39810, n39811, n39812, n39813, n39814, n39815, n39816, n39817,
         n39818, n39819, n39820, n39821, n39822, n39823, n39824, n39825,
         n39826, n39827, n39828, n39829, n39830, n39831, n39832, n39833,
         n39834, n39835, n39836, n39837, n39838, n39839, n39840, n39841,
         n39842, n39843, n39844, n39845, n39846, n39847, n39848, n39849,
         n39850, n39851, n39852, n39853, n39854, n39855, n39856, n39857,
         n39858, n39859, n39860, n39861, n39862, n39863, n39864, n39865,
         n39866, n39867, n39868, n39869, n39870, n39871, n39872, n39873,
         n39874, n39875, n39876, n39877, n39878, n39879, n39880, n39881,
         n39882, n39883, n39884, n39885, n39886, n39887, n39888, n39889,
         n39890, n39891, n39892, n39893, n39894, n39895, n39896, n39897,
         n39898, n39899, n39900, n39901, n39902, n39903, n39904, n39905,
         n39906, n39907, n39908, n39909, n39910, n39911, n39912, n39913,
         n39914, n39915, n39916, n39917, n39918, n39919, n39920, n39921,
         n39922, n39923, n39924, n39925, n39926, n39927, n39928, n39929,
         n39930, n39931, n39932, n39933, n39934, n39935, n39936, n39937,
         n39938, n39939, n39940, n39941, n39942, n39943, n39944, n39945,
         n39946, n39947, n39948, n39949, n39950, n39951, n39952, n39953,
         n39954, n39955, n39956, n39957, n39958, n39959, n39960, n39961,
         n39962, n39963, n39964, n39965, n39966, n39967, n39968, n39969,
         n39970, n39971, n39972, n39973, n39974, n39975, n39976, n39977,
         n39978, n39979, n39980, n39981, n39982, n39983, n39984, n39985,
         n39986, n39987, n39988, n39989, n39990, n39991, n39992, n39993,
         n39994, n39995, n39996, n39997, n39998, n39999, n40000, n40001,
         n40002, n40003, n40004, n40005, n40006, n40007, n40008, n40009,
         n40010, n40011, n40012, n40013, n40014, n40015, n40016, n40017,
         n40018, n40019, n40020, n40021, n40022, n40023, n40024, n40025,
         n40026, n40027, n40028, n40029, n40030, n40031, n40032, n40033,
         n40034, n40035, n40036, n40037, n40038, n40039, n40040, n40041,
         n40042, n40043, n40044, n40045, n40046, n40047, n40048, n40049,
         n40050, n40051, n40052, n40053, n40054, n40055, n40056, n40057,
         n40058, n40059, n40060, n40061, n40062, n40063, n40064, n40065,
         n40066, n40067, n40068, n40069, n40070, n40071, n40072, n40073,
         n40074, n40075, n40076, n40077, n40078, n40079, n40080, n40081,
         n40082, n40083, n40084, n40085, n40086, n40087, n40088, n40089,
         n40090, n40091, n40092, n40093, n40094, n40095, n40096, n40097,
         n40098, n40099, n40100, n40101, n40102, n40103, n40104, n40105,
         n40106, n40107, n40108, n40109, n40110, n40111, n40112, n40113,
         n40114, n40115, n40116, n40117, n40118, n40119, n40120, n40121,
         n40122, n40123, n40124, n40125, n40126, n40127, n40128, n40129,
         n40130, n40131, n40132, n40133, n40134, n40135, n40136, n40137,
         n40138, n40139, n40140, n40141, n40142, n40143, n40144, n40145,
         n40146, n40147, n40148, n40149, n40150, n40151, n40152, n40153,
         n40154, n40155, n40156, n40157, n40158, n40159, n40160, n40161,
         n40162, n40163, n40164, n40165, n40166, n40167, n40168, n40169,
         n40170, n40171, n40172, n40173, n40174, n40175, n40176, n40177,
         n40178, n40179, n40180, n40181, n40182, n40183, n40184, n40185,
         n40186, n40187, n40188, n40189, n40190, n40191, n40192, n40193,
         n40194, n40195, n40196, n40197, n40198, n40199, n40200, n40201,
         n40202, n40203, n40204, n40205, n40206, n40207, n40208, n40209,
         n40210, n40211, n40212, n40213, n40214, n40215, n40216, n40217,
         n40218, n40219, n40220, n40221, n40222, n40223, n40224, n40225,
         n40226, n40227, n40228, n40229, n40230, n40231, n40232, n40233,
         n40234, n40235, n40236, n40237, n40238, n40239, n40240, n40241,
         n40242, n40243, n40244, n40245, n40246, n40247, n40248, n40249,
         n40250, n40251, n40252, n40253, n40254, n40255, n40256, n40257,
         n40258, n40259, n40260, n40261, n40262, n40263, n40264, n40265,
         n40266, n40267, n40268, n40269, n40270, n40271, n40272, n40273,
         n40274, n40275, n40276, n40277, n40278, n40279, n40280, n40281,
         n40282, n40283, n40284, n40285, n40286, n40287, n40288, n40289,
         n40290, n40291, n40292, n40293, n40294, n40295, n40296, n40297,
         n40298, n40299, n40300, n40301, n40302, n40303, n40304, n40305,
         n40306, n40307, n40308, n40309, n40310, n40311, n40312, n40313,
         n40314, n40315, n40316, n40317, n40318, n40319, n40320, n40321,
         n40322, n40323, n40324, n40325, n40326, n40327, n40328, n40329,
         n40330, n40331, n40332, n40333, n40334, n40335, n40336, n40337,
         n40338, n40339, n40340, n40341, n40342, n40343, n40344, n40345,
         n40346, n40347, n40348, n40349, n40350, n40351, n40352, n40353,
         n40354, n40355, n40356, n40357, n40358, n40359, n40360, n40361,
         n40362, n40363, n40364, n40365, n40366, n40367, n40368, n40369,
         n40370, n40371, n40372, n40373, n40374, n40375, n40376, n40377,
         n40378, n40379, n40380, n40381, n40382, n40383, n40384, n40385,
         n40386, n40387, n40388, n40389, n40390, n40391, n40392, n40393,
         n40394, n40395, n40396, n40397, n40398, n40399, n40400, n40401,
         n40402, n40403, n40404, n40405, n40406, n40407, n40408, n40409,
         n40410, n40411, n40412, n40413, n40414, n40415, n40416, n40417,
         n40418, n40419, n40420, n40421, n40422, n40423, n40424, n40425,
         n40426, n40427, n40428, n40429, n40430, n40431, n40432, n40433,
         n40434, n40435, n40436, n40437, n40438, n40439, n40440, n40441,
         n40442, n40443, n40444, n40445, n40446, n40447, n40448, n40449,
         n40450, n40451, n40452, n40453, n40454, n40455, n40456, n40457,
         n40458, n40459, n40460, n40461, n40462, n40463, n40464, n40465,
         n40466, n40467, n40468, n40469, n40470, n40471, n40472, n40473,
         n40474, n40475, n40476, n40477, n40478, n40479, n40480, n40481,
         n40482, n40483, n40484, n40485, n40486, n40487, n40488, n40489,
         n40490, n40491, n40492, n40493, n40494, n40495, n40496, n40497,
         n40498, n40499, n40500, n40501, n40502, n40503, n40504, n40505,
         n40506, n40507, n40508, n40509, n40510, n40511, n40512, n40513,
         n40514, n40515, n40516, n40517, n40518, n40519, n40520, n40521,
         n40522, n40523, n40524, n40525, n40526, n40527, n40528, n40529,
         n40530, n40531, n40532, n40533, n40534, n40535, n40536, n40537,
         n40538, n40539, n40540, n40541, n40542, n40543, n40544, n40545,
         n40546, n40547, n40548, n40549, n40550, n40551, n40552, n40553,
         n40554, n40555, n40556, n40557, n40558, n40559, n40560, n40561,
         n40562, n40563, n40564, n40565, n40566, n40567, n40568, n40569,
         n40570, n40571, n40572, n40573, n40574, n40575, n40576, n40577,
         n40578, n40579, n40580, n40581, n40582, n40583, n40584, n40585,
         n40586, n40587, n40588, n40589, n40590, n40591, n40592, n40593,
         n40594, n40595, n40596, n40597, n40598, n40599, n40600, n40601,
         n40602, n40603, n40604, n40605, n40606, n40607, n40608, n40609,
         n40610, n40611, n40612, n40613, n40614, n40615, n40616, n40617,
         n40618, n40619, n40620, n40621, n40622, n40623, n40624, n40625,
         n40626, n40627, n40628, n40629, n40630, n40631, n40632, n40633,
         n40634, n40635, n40636, n40637, n40638, n40639, n40640, n40641,
         n40642, n40643, n40644, n40645, n40646, n40647, n40648, n40649,
         n40650, n40651, n40652, n40653, n40654, n40655, n40656, n40657,
         n40658, n40659, n40660, n40661, n40662, n40663, n40664, n40665,
         n40666, n40667, n40668, n40669, n40670, n40671, n40672, n40673,
         n40674, n40675, n40676, n40677, n40678, n40679, n40680, n40681,
         n40682, n40683, n40684, n40685, n40686, n40687, n40688, n40689,
         n40690, n40691, n40692, n40693, n40694, n40695, n40696, n40697,
         n40698, n40699, n40700, n40701, n40702, n40703, n40704, n40705,
         n40706, n40707, n40708, n40709, n40710, n40711, n40712, n40713,
         n40714, n40715, n40716, n40717, n40718, n40719, n40720, n40721,
         n40722, n40723, n40724, n40725, n40726, n40727, n40728, n40729,
         n40730, n40731, n40732, n40733, n40734, n40735, n40736, n40737,
         n40738, n40739, n40740, n40741, n40742, n40743, n40744, n40745,
         n40746, n40747, n40748, n40749, n40750, n40751, n40752, n40753,
         n40754, n40755, n40756, n40757, n40758, n40759, n40760, n40761,
         n40762, n40763, n40764, n40765, n40766, n40767, n40768, n40769,
         n40770, n40771, n40772, n40773, n40774, n40775, n40776, n40777,
         n40778, n40779, n40780, n40781, n40782, n40783, n40784, n40785,
         n40786, n40787, n40788, n40789, n40790, n40791, n40792, n40793,
         n40794, n40795, n40796, n40797, n40798, n40799, n40800, n40801,
         n40802, n40803, n40804, n40805, n40806, n40807, n40808, n40809,
         n40810, n40811, n40812, n40813, n40814, n40815, n40816, n40817,
         n40818, n40819, n40820, n40821, n40822, n40823, n40824, n40825,
         n40826, n40827, n40828, n40829, n40830, n40831, n40832, n40833,
         n40834, n40835, n40836, n40837, n40838, n40839, n40840, n40841,
         n40842, n40843, n40844, n40845, n40846, n40847, n40848, n40849,
         n40850, n40851, n40852, n40853, n40854, n40855, n40856, n40857,
         n40858, n40859, n40860, n40861, n40862, n40863, n40864, n40865,
         n40866, n40867, n40868, n40869, n40870, n40871, n40872, n40873,
         n40874, n40875, n40876, n40877, n40878, n40879, n40880, n40881,
         n40882, n40883, n40884, n40885, n40886, n40887, n40888, n40889,
         n40890, n40891, n40892, n40893, n40894, n40895, n40896, n40897,
         n40898, n40899, n40900, n40901, n40902, n40903, n40904, n40905,
         n40906, n40907, n40908, n40909, n40910, n40911, n40912, n40913,
         n40914, n40915, n40916, n40917, n40918, n40919, n40920, n40921,
         n40922, n40923, n40924, n40925, n40926, n40927, n40928, n40929,
         n40930, n40931, n40932, n40933, n40934, n40935, n40936, n40937,
         n40938, n40939, n40940, n40941, n40942, n40943, n40944, n40945,
         n40946, n40947, n40948, n40949, n40950, n40951, n40952, n40953,
         n40954, n40955, n40956, n40957, n40958, n40959, n40960, n40961,
         n40962, n40963, n40964, n40965, n40966, n40967, n40968, n40969,
         n40970, n40971, n40972, n40973, n40974, n40975, n40976, n40977,
         n40978, n40979, n40980, n40981, n40982, n40983, n40984, n40985,
         n40986, n40987, n40988, n40989, n40990, n40991, n40992, n40993,
         n40994, n40995, n40996, n40997, n40998, n40999, n41000, n41001,
         n41002, n41003, n41004, n41005, n41006, n41007, n41008, n41009,
         n41010, n41011, n41012, n41013, n41014, n41015, n41016, n41017,
         n41018, n41019, n41020, n41021, n41022, n41023, n41024, n41025,
         n41026, n41027, n41028, n41029, n41030, n41031, n41032, n41033,
         n41034, n41035, n41036, n41037, n41038, n41039, n41040, n41041,
         n41042, n41043, n41044, n41045, n41046, n41047, n41048, n41049,
         n41050, n41051, n41052, n41053, n41054, n41055, n41056, n41057,
         n41058, n41059, n41060, n41061, n41062, n41063, n41064, n41065,
         n41066, n41067, n41068, n41069, n41070, n41071, n41072, n41073,
         n41074, n41075, n41076, n41077, n41078, n41079, n41080, n41081,
         n41082, n41083, n41084, n41085, n41086, n41087, n41088, n41089,
         n41090, n41091, n41092, n41093, n41094, n41095, n41096, n41097,
         n41098, n41099, n41100, n41101, n41102, n41103, n41104, n41105,
         n41106, n41107, n41108, n41109, n41110, n41111, n41112, n41113,
         n41114, n41115, n41116, n41117, n41118, n41119, n41120, n41121,
         n41122, n41123, n41124, n41125, n41126, n41127, n41128, n41129,
         n41130, n41131, n41132, n41133, n41134, n41135, n41136, n41137,
         n41138, n41139, n41140, n41141, n41142, n41143, n41144, n41145,
         n41146, n41147, n41148, n41149, n41150, n41151, n41152, n41153,
         n41154, n41155, n41156, n41157, n41158, n41159, n41160, n41161,
         n41162, n41163, n41164, n41165, n41166, n41167, n41168, n41169,
         n41170, n41171, n41172, n41173, n41174, n41175, n41176, n41177,
         n41178, n41179, n41180, n41181, n41182, n41183, n41184, n41185,
         n41186, n41187, n41188, n41189, n41190, n41191, n41192, n41193,
         n41194, n41195, n41196, n41197, n41198, n41199, n41200, n41201,
         n41202, n41203, n41204, n41205, n41206, n41207, n41208, n41209,
         n41210, n41211, n41212, n41213, n41214, n41215, n41216, n41217,
         n41218, n41219, n41220, n41221, n41222, n41223, n41224, n41225,
         n41226, n41227, n41228, n41229, n41230, n41231, n41232, n41233,
         n41234, n41235, n41236, n41237, n41238, n41239, n41240, n41241,
         n41242, n41243, n41244, n41245, n41246, n41247, n41248, n41249,
         n41250, n41251, n41252, n41253, n41254, n41255, n41256, n41257,
         n41258, n41259, n41260, n41261, n41262, n41263, n41264, n41265,
         n41266, n41267, n41268, n41269, n41270, n41271, n41272, n41273,
         n41274, n41275, n41276, n41277, n41278, n41279, n41280, n41281,
         n41282, n41283, n41284, n41285, n41286, n41287, n41288, n41289,
         n41290, n41291, n41292, n41293, n41294, n41295, n41296, n41297,
         n41298, n41299, n41300, n41301, n41302, n41303, n41304, n41305,
         n41306, n41307, n41308, n41309, n41310, n41311, n41312, n41313,
         n41314, n41315, n41316, n41317, n41318, n41319, n41320, n41321,
         n41322, n41323, n41324, n41325, n41326, n41327, n41328, n41329,
         n41330, n41331, n41332, n41333, n41334, n41335, n41336, n41337,
         n41338, n41339, n41340, n41341, n41342, n41343, n41344, n41345,
         n41346, n41347, n41348, n41349, n41350, n41351, n41352, n41353,
         n41354, n41355, n41356, n41357, n41358, n41359, n41360, n41361,
         n41362, n41363, n41364, n41365, n41366, n41367, n41368, n41369,
         n41370, n41371, n41372, n41373, n41374, n41375, n41376, n41377,
         n41378, n41379, n41380, n41381, n41382, n41383, n41384, n41385,
         n41386, n41387, n41388, n41389, n41390, n41391, n41392, n41393,
         n41394, n41395, n41396, n41397, n41398, n41399, n41400, n41401,
         n41402, n41403, n41404, n41405, n41406, n41407, n41408, n41409,
         n41410, n41411, n41412, n41413, n41414, n41415, n41416, n41417,
         n41418, n41419, n41420, n41421, n41422, n41423, n41424, n41425,
         n41426, n41427, n41428, n41429, n41430, n41431, n41432, n41433,
         n41434, n41435, n41436, n41437, n41438, n41439, n41440, n41441,
         n41442, n41443, n41444, n41445, n41446, n41447, n41448, n41449,
         n41450, n41451, n41452, n41453, n41454, n41455, n41456, n41457,
         n41458, n41459, n41460, n41461, n41462, n41463, n41464, n41465,
         n41466, n41467, n41468, n41469, n41470, n41471, n41472, n41473,
         n41474, n41475, n41476, n41477, n41478, n41479, n41480, n41481,
         n41482, n41483, n41484, n41485, n41486, n41487, n41488, n41489,
         n41490, n41491, n41492, n41493, n41494, n41495, n41496, n41497,
         n41498, n41499, n41500, n41501, n41502, n41503, n41504, n41505,
         n41506, n41507, n41508, n41509, n41510, n41511, n41512, n41513,
         n41514, n41515, n41516, n41517, n41518, n41519, n41520, n41521,
         n41522, n41523, n41524, n41525, n41526, n41527, n41528, n41529,
         n41530, n41531, n41532, n41533, n41534, n41535, n41536, n41537,
         n41538, n41539, n41540, n41541, n41542, n41543, n41544, n41545,
         n41546, n41547, n41548, n41549, n41550, n41551, n41552, n41553,
         n41554, n41555, n41556, n41557, n41558, n41559, n41560, n41561,
         n41562, n41563, n41564, n41565, n41566, n41567, n41568, n41569,
         n41570, n41571, n41572, n41573, n41574, n41575, n41576, n41577,
         n41578, n41579, n41580, n41581, n41582, n41583, n41584, n41585,
         n41586, n41587, n41588, n41589, n41590, n41591, n41592, n41593,
         n41594, n41595, n41596, n41597, n41598, n41599, n41600, n41601,
         n41602, n41603, n41604, n41605, n41606, n41607, n41608, n41609,
         n41610, n41611, n41612, n41613, n41614, n41615, n41616, n41617,
         n41618, n41619, n41620, n41621, n41622, n41623, n41624, n41625,
         n41626, n41627, n41628, n41629, n41630, n41631, n41632, n41633,
         n41634, n41635, n41636, n41637, n41638, n41639, n41640, n41641,
         n41642, n41643, n41644, n41645, n41646, n41647, n41648, n41649,
         n41650, n41651, n41652, n41653, n41654, n41655, n41656, n41657,
         n41658, n41659, n41660, n41661, n41662, n41663, n41664, n41665,
         n41666, n41667, n41668, n41669, n41670, n41671, n41672, n41673,
         n41674, n41675, n41676, n41677, n41678, n41679, n41680, n41681,
         n41682, n41683, n41684, n41685, n41686, n41687, n41688, n41689,
         n41690, n41691, n41692, n41693, n41694, n41695, n41696, n41697,
         n41698, n41699, n41700, n41701, n41702, n41703, n41704, n41705,
         n41706, n41707, n41708, n41709, n41710, n41711, n41712, n41713,
         n41714, n41715, n41716, n41717, n41718, n41719, n41720, n41721,
         n41722, n41723, n41724, n41725, n41726, n41727, n41728, n41729,
         n41730, n41731, n41732, n41733, n41734, n41735, n41736, n41737,
         n41738, n41739, n41740, n41741, n41742, n41743, n41744, n41745,
         n41746, n41747, n41748, n41749, n41750, n41751, n41752, n41753,
         n41754, n41755, n41756, n41757, n41758, n41759, n41760, n41761,
         n41762, n41763, n41764, n41765, n41766, n41767, n41768, n41769,
         n41770, n41771, n41772, n41773, n41774, n41775, n41776, n41777,
         n41778, n41779, n41780, n41781, n41782, n41783, n41784, n41785,
         n41786, n41787, n41788, n41789, n41790, n41791, n41792, n41793,
         n41794, n41795, n41796, n41797, n41798, n41799, n41800, n41801,
         n41802, n41803, n41804, n41805, n41806, n41807, n41808, n41809,
         n41810, n41811, n41812, n41813, n41814, n41815, n41816, n41817,
         n41818, n41819, n41820, n41821, n41822, n41823, n41824, n41825,
         n41826, n41827, n41828, n41829, n41830, n41831, n41832, n41833,
         n41834, n41835, n41836, n41837, n41838, n41839, n41840, n41841,
         n41842, n41843, n41844, n41845, n41846, n41847, n41848, n41849,
         n41850, n41851, n41852, n41853, n41854, n41855, n41856, n41857,
         n41858, n41859, n41860, n41861, n41862, n41863, n41864, n41865,
         n41866, n41867, n41868, n41869, n41870, n41871, n41872, n41873,
         n41874, n41875, n41876, n41877, n41878, n41879, n41880, n41881,
         n41882, n41883, n41884, n41885, n41886, n41887, n41888, n41889,
         n41890, n41891, n41892, n41893, n41894, n41895, n41896, n41897,
         n41898, n41899, n41900, n41901, n41902, n41903, n41904, n41905,
         n41906, n41907, n41908, n41909, n41910, n41911, n41912, n41913,
         n41914, n41915, n41916, n41917, n41918, n41919, n41920, n41921,
         n41922, n41923, n41924, n41925, n41926, n41927, n41928, n41929,
         n41930, n41931, n41932, n41933, n41934, n41935, n41936, n41937,
         n41938, n41939, n41940, n41941, n41942, n41943, n41944, n41945,
         n41946, n41947, n41948, n41949, n41950, n41951, n41952, n41953,
         n41954, n41955, n41956, n41957, n41958, n41959, n41960, n41961,
         n41962, n41963, n41964, n41965, n41966, n41967, n41968, n41969,
         n41970, n41971, n41972, n41973, n41974, n41975, n41976, n41977,
         n41978, n41979, n41980, n41981, n41982, n41983, n41984, n41985,
         n41986, n41987, n41988, n41989, n41990, n41991, n41992, n41993,
         n41994, n41995, n41996, n41997, n41998, n41999, n42000, n42001,
         n42002, n42003, n42004, n42005, n42006, n42007, n42008, n42009,
         n42010, n42011, n42012, n42013, n42014, n42015, n42016, n42017,
         n42018, n42019, n42020, n42021, n42022, n42023, n42024, n42025,
         n42026, n42027, n42028, n42029, n42030, n42031, n42032, n42033,
         n42034, n42035, n42036, n42037, n42038, n42039, n42040, n42041,
         n42042, n42043, n42044, n42045, n42046, n42047, n42048, n42049,
         n42050, n42051, n42052, n42053, n42054, n42055, n42056, n42057,
         n42058, n42059, n42060, n42061, n42062, n42063, n42064, n42065,
         n42066, n42067, n42068, n42069, n42070, n42071, n42072, n42073,
         n42074, n42075, n42076, n42077, n42078, n42079, n42080, n42081,
         n42082, n42083, n42084, n42085, n42086, n42087, n42088, n42089,
         n42090, n42091, n42092, n42093, n42094, n42095, n42096, n42097,
         n42098, n42099, n42100, n42101, n42102, n42103, n42104, n42105,
         n42106, n42107, n42108, n42109, n42110, n42111, n42112, n42113,
         n42114, n42115, n42116, n42117, n42118, n42119, n42120, n42121,
         n42122, n42123, n42124, n42125, n42126, n42127, n42128, n42129,
         n42130, n42131, n42132, n42133, n42134, n42135, n42136, n42137,
         n42138, n42139, n42140, n42141, n42142, n42143, n42144, n42145,
         n42146, n42147, n42148, n42149, n42150, n42151, n42152, n42153,
         n42154, n42155, n42156, n42157, n42158, n42159, n42160, n42161,
         n42162, n42163, n42164, n42165, n42166, n42167, n42168, n42169,
         n42170, n42171, n42172, n42173, n42174, n42175, n42176, n42177,
         n42178, n42179, n42180, n42181, n42182, n42183, n42184, n42185,
         n42186, n42187, n42188, n42189, n42190, n42191, n42192, n42193,
         n42194, n42195, n42196, n42197, n42198, n42199, n42200, n42201,
         n42202, n42203, n42204, n42205, n42206, n42207, n42208, n42209,
         n42210, n42211, n42212, n42213, n42214, n42215, n42216, n42217,
         n42218, n42219, n42220, n42221, n42222, n42223, n42224, n42225,
         n42226, n42227, n42228, n42229, n42230, n42231, n42232, n42233,
         n42234, n42235, n42236, n42237, n42238, n42239, n42240, n42241,
         n42242, n42243, n42244, n42245, n42246, n42247, n42248, n42249,
         n42250, n42251, n42252, n42253, n42254, n42255, n42256, n42257,
         n42258, n42259, n42260, n42261, n42262, n42263, n42264, n42265,
         n42266, n42267, n42268, n42269, n42270, n42271, n42272, n42273,
         n42274, n42275, n42276, n42277, n42278, n42279, n42280, n42281,
         n42282, n42283, n42284, n42285, n42286, n42287, n42288;
  wire   [2047:0] sreg;

  DFF \sreg_reg[2039]  ( .D(c[2047]), .CLK(clk), .RST(rst), .Q(sreg[2039]) );
  DFF \sreg_reg[2038]  ( .D(c[2046]), .CLK(clk), .RST(rst), .Q(sreg[2038]) );
  DFF \sreg_reg[2037]  ( .D(c[2045]), .CLK(clk), .RST(rst), .Q(sreg[2037]) );
  DFF \sreg_reg[2036]  ( .D(c[2044]), .CLK(clk), .RST(rst), .Q(sreg[2036]) );
  DFF \sreg_reg[2035]  ( .D(c[2043]), .CLK(clk), .RST(rst), .Q(sreg[2035]) );
  DFF \sreg_reg[2034]  ( .D(c[2042]), .CLK(clk), .RST(rst), .Q(sreg[2034]) );
  DFF \sreg_reg[2033]  ( .D(c[2041]), .CLK(clk), .RST(rst), .Q(sreg[2033]) );
  DFF \sreg_reg[2032]  ( .D(c[2040]), .CLK(clk), .RST(rst), .Q(sreg[2032]) );
  DFF \sreg_reg[2031]  ( .D(c[2039]), .CLK(clk), .RST(rst), .Q(sreg[2031]) );
  DFF \sreg_reg[2030]  ( .D(c[2038]), .CLK(clk), .RST(rst), .Q(sreg[2030]) );
  DFF \sreg_reg[2029]  ( .D(c[2037]), .CLK(clk), .RST(rst), .Q(sreg[2029]) );
  DFF \sreg_reg[2028]  ( .D(c[2036]), .CLK(clk), .RST(rst), .Q(sreg[2028]) );
  DFF \sreg_reg[2027]  ( .D(c[2035]), .CLK(clk), .RST(rst), .Q(sreg[2027]) );
  DFF \sreg_reg[2026]  ( .D(c[2034]), .CLK(clk), .RST(rst), .Q(sreg[2026]) );
  DFF \sreg_reg[2025]  ( .D(c[2033]), .CLK(clk), .RST(rst), .Q(sreg[2025]) );
  DFF \sreg_reg[2024]  ( .D(c[2032]), .CLK(clk), .RST(rst), .Q(sreg[2024]) );
  DFF \sreg_reg[2023]  ( .D(c[2031]), .CLK(clk), .RST(rst), .Q(sreg[2023]) );
  DFF \sreg_reg[2022]  ( .D(c[2030]), .CLK(clk), .RST(rst), .Q(sreg[2022]) );
  DFF \sreg_reg[2021]  ( .D(c[2029]), .CLK(clk), .RST(rst), .Q(sreg[2021]) );
  DFF \sreg_reg[2020]  ( .D(c[2028]), .CLK(clk), .RST(rst), .Q(sreg[2020]) );
  DFF \sreg_reg[2019]  ( .D(c[2027]), .CLK(clk), .RST(rst), .Q(sreg[2019]) );
  DFF \sreg_reg[2018]  ( .D(c[2026]), .CLK(clk), .RST(rst), .Q(sreg[2018]) );
  DFF \sreg_reg[2017]  ( .D(c[2025]), .CLK(clk), .RST(rst), .Q(sreg[2017]) );
  DFF \sreg_reg[2016]  ( .D(c[2024]), .CLK(clk), .RST(rst), .Q(sreg[2016]) );
  DFF \sreg_reg[2015]  ( .D(c[2023]), .CLK(clk), .RST(rst), .Q(sreg[2015]) );
  DFF \sreg_reg[2014]  ( .D(c[2022]), .CLK(clk), .RST(rst), .Q(sreg[2014]) );
  DFF \sreg_reg[2013]  ( .D(c[2021]), .CLK(clk), .RST(rst), .Q(sreg[2013]) );
  DFF \sreg_reg[2012]  ( .D(c[2020]), .CLK(clk), .RST(rst), .Q(sreg[2012]) );
  DFF \sreg_reg[2011]  ( .D(c[2019]), .CLK(clk), .RST(rst), .Q(sreg[2011]) );
  DFF \sreg_reg[2010]  ( .D(c[2018]), .CLK(clk), .RST(rst), .Q(sreg[2010]) );
  DFF \sreg_reg[2009]  ( .D(c[2017]), .CLK(clk), .RST(rst), .Q(sreg[2009]) );
  DFF \sreg_reg[2008]  ( .D(c[2016]), .CLK(clk), .RST(rst), .Q(sreg[2008]) );
  DFF \sreg_reg[2007]  ( .D(c[2015]), .CLK(clk), .RST(rst), .Q(sreg[2007]) );
  DFF \sreg_reg[2006]  ( .D(c[2014]), .CLK(clk), .RST(rst), .Q(sreg[2006]) );
  DFF \sreg_reg[2005]  ( .D(c[2013]), .CLK(clk), .RST(rst), .Q(sreg[2005]) );
  DFF \sreg_reg[2004]  ( .D(c[2012]), .CLK(clk), .RST(rst), .Q(sreg[2004]) );
  DFF \sreg_reg[2003]  ( .D(c[2011]), .CLK(clk), .RST(rst), .Q(sreg[2003]) );
  DFF \sreg_reg[2002]  ( .D(c[2010]), .CLK(clk), .RST(rst), .Q(sreg[2002]) );
  DFF \sreg_reg[2001]  ( .D(c[2009]), .CLK(clk), .RST(rst), .Q(sreg[2001]) );
  DFF \sreg_reg[2000]  ( .D(c[2008]), .CLK(clk), .RST(rst), .Q(sreg[2000]) );
  DFF \sreg_reg[1999]  ( .D(c[2007]), .CLK(clk), .RST(rst), .Q(sreg[1999]) );
  DFF \sreg_reg[1998]  ( .D(c[2006]), .CLK(clk), .RST(rst), .Q(sreg[1998]) );
  DFF \sreg_reg[1997]  ( .D(c[2005]), .CLK(clk), .RST(rst), .Q(sreg[1997]) );
  DFF \sreg_reg[1996]  ( .D(c[2004]), .CLK(clk), .RST(rst), .Q(sreg[1996]) );
  DFF \sreg_reg[1995]  ( .D(c[2003]), .CLK(clk), .RST(rst), .Q(sreg[1995]) );
  DFF \sreg_reg[1994]  ( .D(c[2002]), .CLK(clk), .RST(rst), .Q(sreg[1994]) );
  DFF \sreg_reg[1993]  ( .D(c[2001]), .CLK(clk), .RST(rst), .Q(sreg[1993]) );
  DFF \sreg_reg[1992]  ( .D(c[2000]), .CLK(clk), .RST(rst), .Q(sreg[1992]) );
  DFF \sreg_reg[1991]  ( .D(c[1999]), .CLK(clk), .RST(rst), .Q(sreg[1991]) );
  DFF \sreg_reg[1990]  ( .D(c[1998]), .CLK(clk), .RST(rst), .Q(sreg[1990]) );
  DFF \sreg_reg[1989]  ( .D(c[1997]), .CLK(clk), .RST(rst), .Q(sreg[1989]) );
  DFF \sreg_reg[1988]  ( .D(c[1996]), .CLK(clk), .RST(rst), .Q(sreg[1988]) );
  DFF \sreg_reg[1987]  ( .D(c[1995]), .CLK(clk), .RST(rst), .Q(sreg[1987]) );
  DFF \sreg_reg[1986]  ( .D(c[1994]), .CLK(clk), .RST(rst), .Q(sreg[1986]) );
  DFF \sreg_reg[1985]  ( .D(c[1993]), .CLK(clk), .RST(rst), .Q(sreg[1985]) );
  DFF \sreg_reg[1984]  ( .D(c[1992]), .CLK(clk), .RST(rst), .Q(sreg[1984]) );
  DFF \sreg_reg[1983]  ( .D(c[1991]), .CLK(clk), .RST(rst), .Q(sreg[1983]) );
  DFF \sreg_reg[1982]  ( .D(c[1990]), .CLK(clk), .RST(rst), .Q(sreg[1982]) );
  DFF \sreg_reg[1981]  ( .D(c[1989]), .CLK(clk), .RST(rst), .Q(sreg[1981]) );
  DFF \sreg_reg[1980]  ( .D(c[1988]), .CLK(clk), .RST(rst), .Q(sreg[1980]) );
  DFF \sreg_reg[1979]  ( .D(c[1987]), .CLK(clk), .RST(rst), .Q(sreg[1979]) );
  DFF \sreg_reg[1978]  ( .D(c[1986]), .CLK(clk), .RST(rst), .Q(sreg[1978]) );
  DFF \sreg_reg[1977]  ( .D(c[1985]), .CLK(clk), .RST(rst), .Q(sreg[1977]) );
  DFF \sreg_reg[1976]  ( .D(c[1984]), .CLK(clk), .RST(rst), .Q(sreg[1976]) );
  DFF \sreg_reg[1975]  ( .D(c[1983]), .CLK(clk), .RST(rst), .Q(sreg[1975]) );
  DFF \sreg_reg[1974]  ( .D(c[1982]), .CLK(clk), .RST(rst), .Q(sreg[1974]) );
  DFF \sreg_reg[1973]  ( .D(c[1981]), .CLK(clk), .RST(rst), .Q(sreg[1973]) );
  DFF \sreg_reg[1972]  ( .D(c[1980]), .CLK(clk), .RST(rst), .Q(sreg[1972]) );
  DFF \sreg_reg[1971]  ( .D(c[1979]), .CLK(clk), .RST(rst), .Q(sreg[1971]) );
  DFF \sreg_reg[1970]  ( .D(c[1978]), .CLK(clk), .RST(rst), .Q(sreg[1970]) );
  DFF \sreg_reg[1969]  ( .D(c[1977]), .CLK(clk), .RST(rst), .Q(sreg[1969]) );
  DFF \sreg_reg[1968]  ( .D(c[1976]), .CLK(clk), .RST(rst), .Q(sreg[1968]) );
  DFF \sreg_reg[1967]  ( .D(c[1975]), .CLK(clk), .RST(rst), .Q(sreg[1967]) );
  DFF \sreg_reg[1966]  ( .D(c[1974]), .CLK(clk), .RST(rst), .Q(sreg[1966]) );
  DFF \sreg_reg[1965]  ( .D(c[1973]), .CLK(clk), .RST(rst), .Q(sreg[1965]) );
  DFF \sreg_reg[1964]  ( .D(c[1972]), .CLK(clk), .RST(rst), .Q(sreg[1964]) );
  DFF \sreg_reg[1963]  ( .D(c[1971]), .CLK(clk), .RST(rst), .Q(sreg[1963]) );
  DFF \sreg_reg[1962]  ( .D(c[1970]), .CLK(clk), .RST(rst), .Q(sreg[1962]) );
  DFF \sreg_reg[1961]  ( .D(c[1969]), .CLK(clk), .RST(rst), .Q(sreg[1961]) );
  DFF \sreg_reg[1960]  ( .D(c[1968]), .CLK(clk), .RST(rst), .Q(sreg[1960]) );
  DFF \sreg_reg[1959]  ( .D(c[1967]), .CLK(clk), .RST(rst), .Q(sreg[1959]) );
  DFF \sreg_reg[1958]  ( .D(c[1966]), .CLK(clk), .RST(rst), .Q(sreg[1958]) );
  DFF \sreg_reg[1957]  ( .D(c[1965]), .CLK(clk), .RST(rst), .Q(sreg[1957]) );
  DFF \sreg_reg[1956]  ( .D(c[1964]), .CLK(clk), .RST(rst), .Q(sreg[1956]) );
  DFF \sreg_reg[1955]  ( .D(c[1963]), .CLK(clk), .RST(rst), .Q(sreg[1955]) );
  DFF \sreg_reg[1954]  ( .D(c[1962]), .CLK(clk), .RST(rst), .Q(sreg[1954]) );
  DFF \sreg_reg[1953]  ( .D(c[1961]), .CLK(clk), .RST(rst), .Q(sreg[1953]) );
  DFF \sreg_reg[1952]  ( .D(c[1960]), .CLK(clk), .RST(rst), .Q(sreg[1952]) );
  DFF \sreg_reg[1951]  ( .D(c[1959]), .CLK(clk), .RST(rst), .Q(sreg[1951]) );
  DFF \sreg_reg[1950]  ( .D(c[1958]), .CLK(clk), .RST(rst), .Q(sreg[1950]) );
  DFF \sreg_reg[1949]  ( .D(c[1957]), .CLK(clk), .RST(rst), .Q(sreg[1949]) );
  DFF \sreg_reg[1948]  ( .D(c[1956]), .CLK(clk), .RST(rst), .Q(sreg[1948]) );
  DFF \sreg_reg[1947]  ( .D(c[1955]), .CLK(clk), .RST(rst), .Q(sreg[1947]) );
  DFF \sreg_reg[1946]  ( .D(c[1954]), .CLK(clk), .RST(rst), .Q(sreg[1946]) );
  DFF \sreg_reg[1945]  ( .D(c[1953]), .CLK(clk), .RST(rst), .Q(sreg[1945]) );
  DFF \sreg_reg[1944]  ( .D(c[1952]), .CLK(clk), .RST(rst), .Q(sreg[1944]) );
  DFF \sreg_reg[1943]  ( .D(c[1951]), .CLK(clk), .RST(rst), .Q(sreg[1943]) );
  DFF \sreg_reg[1942]  ( .D(c[1950]), .CLK(clk), .RST(rst), .Q(sreg[1942]) );
  DFF \sreg_reg[1941]  ( .D(c[1949]), .CLK(clk), .RST(rst), .Q(sreg[1941]) );
  DFF \sreg_reg[1940]  ( .D(c[1948]), .CLK(clk), .RST(rst), .Q(sreg[1940]) );
  DFF \sreg_reg[1939]  ( .D(c[1947]), .CLK(clk), .RST(rst), .Q(sreg[1939]) );
  DFF \sreg_reg[1938]  ( .D(c[1946]), .CLK(clk), .RST(rst), .Q(sreg[1938]) );
  DFF \sreg_reg[1937]  ( .D(c[1945]), .CLK(clk), .RST(rst), .Q(sreg[1937]) );
  DFF \sreg_reg[1936]  ( .D(c[1944]), .CLK(clk), .RST(rst), .Q(sreg[1936]) );
  DFF \sreg_reg[1935]  ( .D(c[1943]), .CLK(clk), .RST(rst), .Q(sreg[1935]) );
  DFF \sreg_reg[1934]  ( .D(c[1942]), .CLK(clk), .RST(rst), .Q(sreg[1934]) );
  DFF \sreg_reg[1933]  ( .D(c[1941]), .CLK(clk), .RST(rst), .Q(sreg[1933]) );
  DFF \sreg_reg[1932]  ( .D(c[1940]), .CLK(clk), .RST(rst), .Q(sreg[1932]) );
  DFF \sreg_reg[1931]  ( .D(c[1939]), .CLK(clk), .RST(rst), .Q(sreg[1931]) );
  DFF \sreg_reg[1930]  ( .D(c[1938]), .CLK(clk), .RST(rst), .Q(sreg[1930]) );
  DFF \sreg_reg[1929]  ( .D(c[1937]), .CLK(clk), .RST(rst), .Q(sreg[1929]) );
  DFF \sreg_reg[1928]  ( .D(c[1936]), .CLK(clk), .RST(rst), .Q(sreg[1928]) );
  DFF \sreg_reg[1927]  ( .D(c[1935]), .CLK(clk), .RST(rst), .Q(sreg[1927]) );
  DFF \sreg_reg[1926]  ( .D(c[1934]), .CLK(clk), .RST(rst), .Q(sreg[1926]) );
  DFF \sreg_reg[1925]  ( .D(c[1933]), .CLK(clk), .RST(rst), .Q(sreg[1925]) );
  DFF \sreg_reg[1924]  ( .D(c[1932]), .CLK(clk), .RST(rst), .Q(sreg[1924]) );
  DFF \sreg_reg[1923]  ( .D(c[1931]), .CLK(clk), .RST(rst), .Q(sreg[1923]) );
  DFF \sreg_reg[1922]  ( .D(c[1930]), .CLK(clk), .RST(rst), .Q(sreg[1922]) );
  DFF \sreg_reg[1921]  ( .D(c[1929]), .CLK(clk), .RST(rst), .Q(sreg[1921]) );
  DFF \sreg_reg[1920]  ( .D(c[1928]), .CLK(clk), .RST(rst), .Q(sreg[1920]) );
  DFF \sreg_reg[1919]  ( .D(c[1927]), .CLK(clk), .RST(rst), .Q(sreg[1919]) );
  DFF \sreg_reg[1918]  ( .D(c[1926]), .CLK(clk), .RST(rst), .Q(sreg[1918]) );
  DFF \sreg_reg[1917]  ( .D(c[1925]), .CLK(clk), .RST(rst), .Q(sreg[1917]) );
  DFF \sreg_reg[1916]  ( .D(c[1924]), .CLK(clk), .RST(rst), .Q(sreg[1916]) );
  DFF \sreg_reg[1915]  ( .D(c[1923]), .CLK(clk), .RST(rst), .Q(sreg[1915]) );
  DFF \sreg_reg[1914]  ( .D(c[1922]), .CLK(clk), .RST(rst), .Q(sreg[1914]) );
  DFF \sreg_reg[1913]  ( .D(c[1921]), .CLK(clk), .RST(rst), .Q(sreg[1913]) );
  DFF \sreg_reg[1912]  ( .D(c[1920]), .CLK(clk), .RST(rst), .Q(sreg[1912]) );
  DFF \sreg_reg[1911]  ( .D(c[1919]), .CLK(clk), .RST(rst), .Q(sreg[1911]) );
  DFF \sreg_reg[1910]  ( .D(c[1918]), .CLK(clk), .RST(rst), .Q(sreg[1910]) );
  DFF \sreg_reg[1909]  ( .D(c[1917]), .CLK(clk), .RST(rst), .Q(sreg[1909]) );
  DFF \sreg_reg[1908]  ( .D(c[1916]), .CLK(clk), .RST(rst), .Q(sreg[1908]) );
  DFF \sreg_reg[1907]  ( .D(c[1915]), .CLK(clk), .RST(rst), .Q(sreg[1907]) );
  DFF \sreg_reg[1906]  ( .D(c[1914]), .CLK(clk), .RST(rst), .Q(sreg[1906]) );
  DFF \sreg_reg[1905]  ( .D(c[1913]), .CLK(clk), .RST(rst), .Q(sreg[1905]) );
  DFF \sreg_reg[1904]  ( .D(c[1912]), .CLK(clk), .RST(rst), .Q(sreg[1904]) );
  DFF \sreg_reg[1903]  ( .D(c[1911]), .CLK(clk), .RST(rst), .Q(sreg[1903]) );
  DFF \sreg_reg[1902]  ( .D(c[1910]), .CLK(clk), .RST(rst), .Q(sreg[1902]) );
  DFF \sreg_reg[1901]  ( .D(c[1909]), .CLK(clk), .RST(rst), .Q(sreg[1901]) );
  DFF \sreg_reg[1900]  ( .D(c[1908]), .CLK(clk), .RST(rst), .Q(sreg[1900]) );
  DFF \sreg_reg[1899]  ( .D(c[1907]), .CLK(clk), .RST(rst), .Q(sreg[1899]) );
  DFF \sreg_reg[1898]  ( .D(c[1906]), .CLK(clk), .RST(rst), .Q(sreg[1898]) );
  DFF \sreg_reg[1897]  ( .D(c[1905]), .CLK(clk), .RST(rst), .Q(sreg[1897]) );
  DFF \sreg_reg[1896]  ( .D(c[1904]), .CLK(clk), .RST(rst), .Q(sreg[1896]) );
  DFF \sreg_reg[1895]  ( .D(c[1903]), .CLK(clk), .RST(rst), .Q(sreg[1895]) );
  DFF \sreg_reg[1894]  ( .D(c[1902]), .CLK(clk), .RST(rst), .Q(sreg[1894]) );
  DFF \sreg_reg[1893]  ( .D(c[1901]), .CLK(clk), .RST(rst), .Q(sreg[1893]) );
  DFF \sreg_reg[1892]  ( .D(c[1900]), .CLK(clk), .RST(rst), .Q(sreg[1892]) );
  DFF \sreg_reg[1891]  ( .D(c[1899]), .CLK(clk), .RST(rst), .Q(sreg[1891]) );
  DFF \sreg_reg[1890]  ( .D(c[1898]), .CLK(clk), .RST(rst), .Q(sreg[1890]) );
  DFF \sreg_reg[1889]  ( .D(c[1897]), .CLK(clk), .RST(rst), .Q(sreg[1889]) );
  DFF \sreg_reg[1888]  ( .D(c[1896]), .CLK(clk), .RST(rst), .Q(sreg[1888]) );
  DFF \sreg_reg[1887]  ( .D(c[1895]), .CLK(clk), .RST(rst), .Q(sreg[1887]) );
  DFF \sreg_reg[1886]  ( .D(c[1894]), .CLK(clk), .RST(rst), .Q(sreg[1886]) );
  DFF \sreg_reg[1885]  ( .D(c[1893]), .CLK(clk), .RST(rst), .Q(sreg[1885]) );
  DFF \sreg_reg[1884]  ( .D(c[1892]), .CLK(clk), .RST(rst), .Q(sreg[1884]) );
  DFF \sreg_reg[1883]  ( .D(c[1891]), .CLK(clk), .RST(rst), .Q(sreg[1883]) );
  DFF \sreg_reg[1882]  ( .D(c[1890]), .CLK(clk), .RST(rst), .Q(sreg[1882]) );
  DFF \sreg_reg[1881]  ( .D(c[1889]), .CLK(clk), .RST(rst), .Q(sreg[1881]) );
  DFF \sreg_reg[1880]  ( .D(c[1888]), .CLK(clk), .RST(rst), .Q(sreg[1880]) );
  DFF \sreg_reg[1879]  ( .D(c[1887]), .CLK(clk), .RST(rst), .Q(sreg[1879]) );
  DFF \sreg_reg[1878]  ( .D(c[1886]), .CLK(clk), .RST(rst), .Q(sreg[1878]) );
  DFF \sreg_reg[1877]  ( .D(c[1885]), .CLK(clk), .RST(rst), .Q(sreg[1877]) );
  DFF \sreg_reg[1876]  ( .D(c[1884]), .CLK(clk), .RST(rst), .Q(sreg[1876]) );
  DFF \sreg_reg[1875]  ( .D(c[1883]), .CLK(clk), .RST(rst), .Q(sreg[1875]) );
  DFF \sreg_reg[1874]  ( .D(c[1882]), .CLK(clk), .RST(rst), .Q(sreg[1874]) );
  DFF \sreg_reg[1873]  ( .D(c[1881]), .CLK(clk), .RST(rst), .Q(sreg[1873]) );
  DFF \sreg_reg[1872]  ( .D(c[1880]), .CLK(clk), .RST(rst), .Q(sreg[1872]) );
  DFF \sreg_reg[1871]  ( .D(c[1879]), .CLK(clk), .RST(rst), .Q(sreg[1871]) );
  DFF \sreg_reg[1870]  ( .D(c[1878]), .CLK(clk), .RST(rst), .Q(sreg[1870]) );
  DFF \sreg_reg[1869]  ( .D(c[1877]), .CLK(clk), .RST(rst), .Q(sreg[1869]) );
  DFF \sreg_reg[1868]  ( .D(c[1876]), .CLK(clk), .RST(rst), .Q(sreg[1868]) );
  DFF \sreg_reg[1867]  ( .D(c[1875]), .CLK(clk), .RST(rst), .Q(sreg[1867]) );
  DFF \sreg_reg[1866]  ( .D(c[1874]), .CLK(clk), .RST(rst), .Q(sreg[1866]) );
  DFF \sreg_reg[1865]  ( .D(c[1873]), .CLK(clk), .RST(rst), .Q(sreg[1865]) );
  DFF \sreg_reg[1864]  ( .D(c[1872]), .CLK(clk), .RST(rst), .Q(sreg[1864]) );
  DFF \sreg_reg[1863]  ( .D(c[1871]), .CLK(clk), .RST(rst), .Q(sreg[1863]) );
  DFF \sreg_reg[1862]  ( .D(c[1870]), .CLK(clk), .RST(rst), .Q(sreg[1862]) );
  DFF \sreg_reg[1861]  ( .D(c[1869]), .CLK(clk), .RST(rst), .Q(sreg[1861]) );
  DFF \sreg_reg[1860]  ( .D(c[1868]), .CLK(clk), .RST(rst), .Q(sreg[1860]) );
  DFF \sreg_reg[1859]  ( .D(c[1867]), .CLK(clk), .RST(rst), .Q(sreg[1859]) );
  DFF \sreg_reg[1858]  ( .D(c[1866]), .CLK(clk), .RST(rst), .Q(sreg[1858]) );
  DFF \sreg_reg[1857]  ( .D(c[1865]), .CLK(clk), .RST(rst), .Q(sreg[1857]) );
  DFF \sreg_reg[1856]  ( .D(c[1864]), .CLK(clk), .RST(rst), .Q(sreg[1856]) );
  DFF \sreg_reg[1855]  ( .D(c[1863]), .CLK(clk), .RST(rst), .Q(sreg[1855]) );
  DFF \sreg_reg[1854]  ( .D(c[1862]), .CLK(clk), .RST(rst), .Q(sreg[1854]) );
  DFF \sreg_reg[1853]  ( .D(c[1861]), .CLK(clk), .RST(rst), .Q(sreg[1853]) );
  DFF \sreg_reg[1852]  ( .D(c[1860]), .CLK(clk), .RST(rst), .Q(sreg[1852]) );
  DFF \sreg_reg[1851]  ( .D(c[1859]), .CLK(clk), .RST(rst), .Q(sreg[1851]) );
  DFF \sreg_reg[1850]  ( .D(c[1858]), .CLK(clk), .RST(rst), .Q(sreg[1850]) );
  DFF \sreg_reg[1849]  ( .D(c[1857]), .CLK(clk), .RST(rst), .Q(sreg[1849]) );
  DFF \sreg_reg[1848]  ( .D(c[1856]), .CLK(clk), .RST(rst), .Q(sreg[1848]) );
  DFF \sreg_reg[1847]  ( .D(c[1855]), .CLK(clk), .RST(rst), .Q(sreg[1847]) );
  DFF \sreg_reg[1846]  ( .D(c[1854]), .CLK(clk), .RST(rst), .Q(sreg[1846]) );
  DFF \sreg_reg[1845]  ( .D(c[1853]), .CLK(clk), .RST(rst), .Q(sreg[1845]) );
  DFF \sreg_reg[1844]  ( .D(c[1852]), .CLK(clk), .RST(rst), .Q(sreg[1844]) );
  DFF \sreg_reg[1843]  ( .D(c[1851]), .CLK(clk), .RST(rst), .Q(sreg[1843]) );
  DFF \sreg_reg[1842]  ( .D(c[1850]), .CLK(clk), .RST(rst), .Q(sreg[1842]) );
  DFF \sreg_reg[1841]  ( .D(c[1849]), .CLK(clk), .RST(rst), .Q(sreg[1841]) );
  DFF \sreg_reg[1840]  ( .D(c[1848]), .CLK(clk), .RST(rst), .Q(sreg[1840]) );
  DFF \sreg_reg[1839]  ( .D(c[1847]), .CLK(clk), .RST(rst), .Q(sreg[1839]) );
  DFF \sreg_reg[1838]  ( .D(c[1846]), .CLK(clk), .RST(rst), .Q(sreg[1838]) );
  DFF \sreg_reg[1837]  ( .D(c[1845]), .CLK(clk), .RST(rst), .Q(sreg[1837]) );
  DFF \sreg_reg[1836]  ( .D(c[1844]), .CLK(clk), .RST(rst), .Q(sreg[1836]) );
  DFF \sreg_reg[1835]  ( .D(c[1843]), .CLK(clk), .RST(rst), .Q(sreg[1835]) );
  DFF \sreg_reg[1834]  ( .D(c[1842]), .CLK(clk), .RST(rst), .Q(sreg[1834]) );
  DFF \sreg_reg[1833]  ( .D(c[1841]), .CLK(clk), .RST(rst), .Q(sreg[1833]) );
  DFF \sreg_reg[1832]  ( .D(c[1840]), .CLK(clk), .RST(rst), .Q(sreg[1832]) );
  DFF \sreg_reg[1831]  ( .D(c[1839]), .CLK(clk), .RST(rst), .Q(sreg[1831]) );
  DFF \sreg_reg[1830]  ( .D(c[1838]), .CLK(clk), .RST(rst), .Q(sreg[1830]) );
  DFF \sreg_reg[1829]  ( .D(c[1837]), .CLK(clk), .RST(rst), .Q(sreg[1829]) );
  DFF \sreg_reg[1828]  ( .D(c[1836]), .CLK(clk), .RST(rst), .Q(sreg[1828]) );
  DFF \sreg_reg[1827]  ( .D(c[1835]), .CLK(clk), .RST(rst), .Q(sreg[1827]) );
  DFF \sreg_reg[1826]  ( .D(c[1834]), .CLK(clk), .RST(rst), .Q(sreg[1826]) );
  DFF \sreg_reg[1825]  ( .D(c[1833]), .CLK(clk), .RST(rst), .Q(sreg[1825]) );
  DFF \sreg_reg[1824]  ( .D(c[1832]), .CLK(clk), .RST(rst), .Q(sreg[1824]) );
  DFF \sreg_reg[1823]  ( .D(c[1831]), .CLK(clk), .RST(rst), .Q(sreg[1823]) );
  DFF \sreg_reg[1822]  ( .D(c[1830]), .CLK(clk), .RST(rst), .Q(sreg[1822]) );
  DFF \sreg_reg[1821]  ( .D(c[1829]), .CLK(clk), .RST(rst), .Q(sreg[1821]) );
  DFF \sreg_reg[1820]  ( .D(c[1828]), .CLK(clk), .RST(rst), .Q(sreg[1820]) );
  DFF \sreg_reg[1819]  ( .D(c[1827]), .CLK(clk), .RST(rst), .Q(sreg[1819]) );
  DFF \sreg_reg[1818]  ( .D(c[1826]), .CLK(clk), .RST(rst), .Q(sreg[1818]) );
  DFF \sreg_reg[1817]  ( .D(c[1825]), .CLK(clk), .RST(rst), .Q(sreg[1817]) );
  DFF \sreg_reg[1816]  ( .D(c[1824]), .CLK(clk), .RST(rst), .Q(sreg[1816]) );
  DFF \sreg_reg[1815]  ( .D(c[1823]), .CLK(clk), .RST(rst), .Q(sreg[1815]) );
  DFF \sreg_reg[1814]  ( .D(c[1822]), .CLK(clk), .RST(rst), .Q(sreg[1814]) );
  DFF \sreg_reg[1813]  ( .D(c[1821]), .CLK(clk), .RST(rst), .Q(sreg[1813]) );
  DFF \sreg_reg[1812]  ( .D(c[1820]), .CLK(clk), .RST(rst), .Q(sreg[1812]) );
  DFF \sreg_reg[1811]  ( .D(c[1819]), .CLK(clk), .RST(rst), .Q(sreg[1811]) );
  DFF \sreg_reg[1810]  ( .D(c[1818]), .CLK(clk), .RST(rst), .Q(sreg[1810]) );
  DFF \sreg_reg[1809]  ( .D(c[1817]), .CLK(clk), .RST(rst), .Q(sreg[1809]) );
  DFF \sreg_reg[1808]  ( .D(c[1816]), .CLK(clk), .RST(rst), .Q(sreg[1808]) );
  DFF \sreg_reg[1807]  ( .D(c[1815]), .CLK(clk), .RST(rst), .Q(sreg[1807]) );
  DFF \sreg_reg[1806]  ( .D(c[1814]), .CLK(clk), .RST(rst), .Q(sreg[1806]) );
  DFF \sreg_reg[1805]  ( .D(c[1813]), .CLK(clk), .RST(rst), .Q(sreg[1805]) );
  DFF \sreg_reg[1804]  ( .D(c[1812]), .CLK(clk), .RST(rst), .Q(sreg[1804]) );
  DFF \sreg_reg[1803]  ( .D(c[1811]), .CLK(clk), .RST(rst), .Q(sreg[1803]) );
  DFF \sreg_reg[1802]  ( .D(c[1810]), .CLK(clk), .RST(rst), .Q(sreg[1802]) );
  DFF \sreg_reg[1801]  ( .D(c[1809]), .CLK(clk), .RST(rst), .Q(sreg[1801]) );
  DFF \sreg_reg[1800]  ( .D(c[1808]), .CLK(clk), .RST(rst), .Q(sreg[1800]) );
  DFF \sreg_reg[1799]  ( .D(c[1807]), .CLK(clk), .RST(rst), .Q(sreg[1799]) );
  DFF \sreg_reg[1798]  ( .D(c[1806]), .CLK(clk), .RST(rst), .Q(sreg[1798]) );
  DFF \sreg_reg[1797]  ( .D(c[1805]), .CLK(clk), .RST(rst), .Q(sreg[1797]) );
  DFF \sreg_reg[1796]  ( .D(c[1804]), .CLK(clk), .RST(rst), .Q(sreg[1796]) );
  DFF \sreg_reg[1795]  ( .D(c[1803]), .CLK(clk), .RST(rst), .Q(sreg[1795]) );
  DFF \sreg_reg[1794]  ( .D(c[1802]), .CLK(clk), .RST(rst), .Q(sreg[1794]) );
  DFF \sreg_reg[1793]  ( .D(c[1801]), .CLK(clk), .RST(rst), .Q(sreg[1793]) );
  DFF \sreg_reg[1792]  ( .D(c[1800]), .CLK(clk), .RST(rst), .Q(sreg[1792]) );
  DFF \sreg_reg[1791]  ( .D(c[1799]), .CLK(clk), .RST(rst), .Q(sreg[1791]) );
  DFF \sreg_reg[1790]  ( .D(c[1798]), .CLK(clk), .RST(rst), .Q(sreg[1790]) );
  DFF \sreg_reg[1789]  ( .D(c[1797]), .CLK(clk), .RST(rst), .Q(sreg[1789]) );
  DFF \sreg_reg[1788]  ( .D(c[1796]), .CLK(clk), .RST(rst), .Q(sreg[1788]) );
  DFF \sreg_reg[1787]  ( .D(c[1795]), .CLK(clk), .RST(rst), .Q(sreg[1787]) );
  DFF \sreg_reg[1786]  ( .D(c[1794]), .CLK(clk), .RST(rst), .Q(sreg[1786]) );
  DFF \sreg_reg[1785]  ( .D(c[1793]), .CLK(clk), .RST(rst), .Q(sreg[1785]) );
  DFF \sreg_reg[1784]  ( .D(c[1792]), .CLK(clk), .RST(rst), .Q(sreg[1784]) );
  DFF \sreg_reg[1783]  ( .D(c[1791]), .CLK(clk), .RST(rst), .Q(sreg[1783]) );
  DFF \sreg_reg[1782]  ( .D(c[1790]), .CLK(clk), .RST(rst), .Q(sreg[1782]) );
  DFF \sreg_reg[1781]  ( .D(c[1789]), .CLK(clk), .RST(rst), .Q(sreg[1781]) );
  DFF \sreg_reg[1780]  ( .D(c[1788]), .CLK(clk), .RST(rst), .Q(sreg[1780]) );
  DFF \sreg_reg[1779]  ( .D(c[1787]), .CLK(clk), .RST(rst), .Q(sreg[1779]) );
  DFF \sreg_reg[1778]  ( .D(c[1786]), .CLK(clk), .RST(rst), .Q(sreg[1778]) );
  DFF \sreg_reg[1777]  ( .D(c[1785]), .CLK(clk), .RST(rst), .Q(sreg[1777]) );
  DFF \sreg_reg[1776]  ( .D(c[1784]), .CLK(clk), .RST(rst), .Q(sreg[1776]) );
  DFF \sreg_reg[1775]  ( .D(c[1783]), .CLK(clk), .RST(rst), .Q(sreg[1775]) );
  DFF \sreg_reg[1774]  ( .D(c[1782]), .CLK(clk), .RST(rst), .Q(sreg[1774]) );
  DFF \sreg_reg[1773]  ( .D(c[1781]), .CLK(clk), .RST(rst), .Q(sreg[1773]) );
  DFF \sreg_reg[1772]  ( .D(c[1780]), .CLK(clk), .RST(rst), .Q(sreg[1772]) );
  DFF \sreg_reg[1771]  ( .D(c[1779]), .CLK(clk), .RST(rst), .Q(sreg[1771]) );
  DFF \sreg_reg[1770]  ( .D(c[1778]), .CLK(clk), .RST(rst), .Q(sreg[1770]) );
  DFF \sreg_reg[1769]  ( .D(c[1777]), .CLK(clk), .RST(rst), .Q(sreg[1769]) );
  DFF \sreg_reg[1768]  ( .D(c[1776]), .CLK(clk), .RST(rst), .Q(sreg[1768]) );
  DFF \sreg_reg[1767]  ( .D(c[1775]), .CLK(clk), .RST(rst), .Q(sreg[1767]) );
  DFF \sreg_reg[1766]  ( .D(c[1774]), .CLK(clk), .RST(rst), .Q(sreg[1766]) );
  DFF \sreg_reg[1765]  ( .D(c[1773]), .CLK(clk), .RST(rst), .Q(sreg[1765]) );
  DFF \sreg_reg[1764]  ( .D(c[1772]), .CLK(clk), .RST(rst), .Q(sreg[1764]) );
  DFF \sreg_reg[1763]  ( .D(c[1771]), .CLK(clk), .RST(rst), .Q(sreg[1763]) );
  DFF \sreg_reg[1762]  ( .D(c[1770]), .CLK(clk), .RST(rst), .Q(sreg[1762]) );
  DFF \sreg_reg[1761]  ( .D(c[1769]), .CLK(clk), .RST(rst), .Q(sreg[1761]) );
  DFF \sreg_reg[1760]  ( .D(c[1768]), .CLK(clk), .RST(rst), .Q(sreg[1760]) );
  DFF \sreg_reg[1759]  ( .D(c[1767]), .CLK(clk), .RST(rst), .Q(sreg[1759]) );
  DFF \sreg_reg[1758]  ( .D(c[1766]), .CLK(clk), .RST(rst), .Q(sreg[1758]) );
  DFF \sreg_reg[1757]  ( .D(c[1765]), .CLK(clk), .RST(rst), .Q(sreg[1757]) );
  DFF \sreg_reg[1756]  ( .D(c[1764]), .CLK(clk), .RST(rst), .Q(sreg[1756]) );
  DFF \sreg_reg[1755]  ( .D(c[1763]), .CLK(clk), .RST(rst), .Q(sreg[1755]) );
  DFF \sreg_reg[1754]  ( .D(c[1762]), .CLK(clk), .RST(rst), .Q(sreg[1754]) );
  DFF \sreg_reg[1753]  ( .D(c[1761]), .CLK(clk), .RST(rst), .Q(sreg[1753]) );
  DFF \sreg_reg[1752]  ( .D(c[1760]), .CLK(clk), .RST(rst), .Q(sreg[1752]) );
  DFF \sreg_reg[1751]  ( .D(c[1759]), .CLK(clk), .RST(rst), .Q(sreg[1751]) );
  DFF \sreg_reg[1750]  ( .D(c[1758]), .CLK(clk), .RST(rst), .Q(sreg[1750]) );
  DFF \sreg_reg[1749]  ( .D(c[1757]), .CLK(clk), .RST(rst), .Q(sreg[1749]) );
  DFF \sreg_reg[1748]  ( .D(c[1756]), .CLK(clk), .RST(rst), .Q(sreg[1748]) );
  DFF \sreg_reg[1747]  ( .D(c[1755]), .CLK(clk), .RST(rst), .Q(sreg[1747]) );
  DFF \sreg_reg[1746]  ( .D(c[1754]), .CLK(clk), .RST(rst), .Q(sreg[1746]) );
  DFF \sreg_reg[1745]  ( .D(c[1753]), .CLK(clk), .RST(rst), .Q(sreg[1745]) );
  DFF \sreg_reg[1744]  ( .D(c[1752]), .CLK(clk), .RST(rst), .Q(sreg[1744]) );
  DFF \sreg_reg[1743]  ( .D(c[1751]), .CLK(clk), .RST(rst), .Q(sreg[1743]) );
  DFF \sreg_reg[1742]  ( .D(c[1750]), .CLK(clk), .RST(rst), .Q(sreg[1742]) );
  DFF \sreg_reg[1741]  ( .D(c[1749]), .CLK(clk), .RST(rst), .Q(sreg[1741]) );
  DFF \sreg_reg[1740]  ( .D(c[1748]), .CLK(clk), .RST(rst), .Q(sreg[1740]) );
  DFF \sreg_reg[1739]  ( .D(c[1747]), .CLK(clk), .RST(rst), .Q(sreg[1739]) );
  DFF \sreg_reg[1738]  ( .D(c[1746]), .CLK(clk), .RST(rst), .Q(sreg[1738]) );
  DFF \sreg_reg[1737]  ( .D(c[1745]), .CLK(clk), .RST(rst), .Q(sreg[1737]) );
  DFF \sreg_reg[1736]  ( .D(c[1744]), .CLK(clk), .RST(rst), .Q(sreg[1736]) );
  DFF \sreg_reg[1735]  ( .D(c[1743]), .CLK(clk), .RST(rst), .Q(sreg[1735]) );
  DFF \sreg_reg[1734]  ( .D(c[1742]), .CLK(clk), .RST(rst), .Q(sreg[1734]) );
  DFF \sreg_reg[1733]  ( .D(c[1741]), .CLK(clk), .RST(rst), .Q(sreg[1733]) );
  DFF \sreg_reg[1732]  ( .D(c[1740]), .CLK(clk), .RST(rst), .Q(sreg[1732]) );
  DFF \sreg_reg[1731]  ( .D(c[1739]), .CLK(clk), .RST(rst), .Q(sreg[1731]) );
  DFF \sreg_reg[1730]  ( .D(c[1738]), .CLK(clk), .RST(rst), .Q(sreg[1730]) );
  DFF \sreg_reg[1729]  ( .D(c[1737]), .CLK(clk), .RST(rst), .Q(sreg[1729]) );
  DFF \sreg_reg[1728]  ( .D(c[1736]), .CLK(clk), .RST(rst), .Q(sreg[1728]) );
  DFF \sreg_reg[1727]  ( .D(c[1735]), .CLK(clk), .RST(rst), .Q(sreg[1727]) );
  DFF \sreg_reg[1726]  ( .D(c[1734]), .CLK(clk), .RST(rst), .Q(sreg[1726]) );
  DFF \sreg_reg[1725]  ( .D(c[1733]), .CLK(clk), .RST(rst), .Q(sreg[1725]) );
  DFF \sreg_reg[1724]  ( .D(c[1732]), .CLK(clk), .RST(rst), .Q(sreg[1724]) );
  DFF \sreg_reg[1723]  ( .D(c[1731]), .CLK(clk), .RST(rst), .Q(sreg[1723]) );
  DFF \sreg_reg[1722]  ( .D(c[1730]), .CLK(clk), .RST(rst), .Q(sreg[1722]) );
  DFF \sreg_reg[1721]  ( .D(c[1729]), .CLK(clk), .RST(rst), .Q(sreg[1721]) );
  DFF \sreg_reg[1720]  ( .D(c[1728]), .CLK(clk), .RST(rst), .Q(sreg[1720]) );
  DFF \sreg_reg[1719]  ( .D(c[1727]), .CLK(clk), .RST(rst), .Q(sreg[1719]) );
  DFF \sreg_reg[1718]  ( .D(c[1726]), .CLK(clk), .RST(rst), .Q(sreg[1718]) );
  DFF \sreg_reg[1717]  ( .D(c[1725]), .CLK(clk), .RST(rst), .Q(sreg[1717]) );
  DFF \sreg_reg[1716]  ( .D(c[1724]), .CLK(clk), .RST(rst), .Q(sreg[1716]) );
  DFF \sreg_reg[1715]  ( .D(c[1723]), .CLK(clk), .RST(rst), .Q(sreg[1715]) );
  DFF \sreg_reg[1714]  ( .D(c[1722]), .CLK(clk), .RST(rst), .Q(sreg[1714]) );
  DFF \sreg_reg[1713]  ( .D(c[1721]), .CLK(clk), .RST(rst), .Q(sreg[1713]) );
  DFF \sreg_reg[1712]  ( .D(c[1720]), .CLK(clk), .RST(rst), .Q(sreg[1712]) );
  DFF \sreg_reg[1711]  ( .D(c[1719]), .CLK(clk), .RST(rst), .Q(sreg[1711]) );
  DFF \sreg_reg[1710]  ( .D(c[1718]), .CLK(clk), .RST(rst), .Q(sreg[1710]) );
  DFF \sreg_reg[1709]  ( .D(c[1717]), .CLK(clk), .RST(rst), .Q(sreg[1709]) );
  DFF \sreg_reg[1708]  ( .D(c[1716]), .CLK(clk), .RST(rst), .Q(sreg[1708]) );
  DFF \sreg_reg[1707]  ( .D(c[1715]), .CLK(clk), .RST(rst), .Q(sreg[1707]) );
  DFF \sreg_reg[1706]  ( .D(c[1714]), .CLK(clk), .RST(rst), .Q(sreg[1706]) );
  DFF \sreg_reg[1705]  ( .D(c[1713]), .CLK(clk), .RST(rst), .Q(sreg[1705]) );
  DFF \sreg_reg[1704]  ( .D(c[1712]), .CLK(clk), .RST(rst), .Q(sreg[1704]) );
  DFF \sreg_reg[1703]  ( .D(c[1711]), .CLK(clk), .RST(rst), .Q(sreg[1703]) );
  DFF \sreg_reg[1702]  ( .D(c[1710]), .CLK(clk), .RST(rst), .Q(sreg[1702]) );
  DFF \sreg_reg[1701]  ( .D(c[1709]), .CLK(clk), .RST(rst), .Q(sreg[1701]) );
  DFF \sreg_reg[1700]  ( .D(c[1708]), .CLK(clk), .RST(rst), .Q(sreg[1700]) );
  DFF \sreg_reg[1699]  ( .D(c[1707]), .CLK(clk), .RST(rst), .Q(sreg[1699]) );
  DFF \sreg_reg[1698]  ( .D(c[1706]), .CLK(clk), .RST(rst), .Q(sreg[1698]) );
  DFF \sreg_reg[1697]  ( .D(c[1705]), .CLK(clk), .RST(rst), .Q(sreg[1697]) );
  DFF \sreg_reg[1696]  ( .D(c[1704]), .CLK(clk), .RST(rst), .Q(sreg[1696]) );
  DFF \sreg_reg[1695]  ( .D(c[1703]), .CLK(clk), .RST(rst), .Q(sreg[1695]) );
  DFF \sreg_reg[1694]  ( .D(c[1702]), .CLK(clk), .RST(rst), .Q(sreg[1694]) );
  DFF \sreg_reg[1693]  ( .D(c[1701]), .CLK(clk), .RST(rst), .Q(sreg[1693]) );
  DFF \sreg_reg[1692]  ( .D(c[1700]), .CLK(clk), .RST(rst), .Q(sreg[1692]) );
  DFF \sreg_reg[1691]  ( .D(c[1699]), .CLK(clk), .RST(rst), .Q(sreg[1691]) );
  DFF \sreg_reg[1690]  ( .D(c[1698]), .CLK(clk), .RST(rst), .Q(sreg[1690]) );
  DFF \sreg_reg[1689]  ( .D(c[1697]), .CLK(clk), .RST(rst), .Q(sreg[1689]) );
  DFF \sreg_reg[1688]  ( .D(c[1696]), .CLK(clk), .RST(rst), .Q(sreg[1688]) );
  DFF \sreg_reg[1687]  ( .D(c[1695]), .CLK(clk), .RST(rst), .Q(sreg[1687]) );
  DFF \sreg_reg[1686]  ( .D(c[1694]), .CLK(clk), .RST(rst), .Q(sreg[1686]) );
  DFF \sreg_reg[1685]  ( .D(c[1693]), .CLK(clk), .RST(rst), .Q(sreg[1685]) );
  DFF \sreg_reg[1684]  ( .D(c[1692]), .CLK(clk), .RST(rst), .Q(sreg[1684]) );
  DFF \sreg_reg[1683]  ( .D(c[1691]), .CLK(clk), .RST(rst), .Q(sreg[1683]) );
  DFF \sreg_reg[1682]  ( .D(c[1690]), .CLK(clk), .RST(rst), .Q(sreg[1682]) );
  DFF \sreg_reg[1681]  ( .D(c[1689]), .CLK(clk), .RST(rst), .Q(sreg[1681]) );
  DFF \sreg_reg[1680]  ( .D(c[1688]), .CLK(clk), .RST(rst), .Q(sreg[1680]) );
  DFF \sreg_reg[1679]  ( .D(c[1687]), .CLK(clk), .RST(rst), .Q(sreg[1679]) );
  DFF \sreg_reg[1678]  ( .D(c[1686]), .CLK(clk), .RST(rst), .Q(sreg[1678]) );
  DFF \sreg_reg[1677]  ( .D(c[1685]), .CLK(clk), .RST(rst), .Q(sreg[1677]) );
  DFF \sreg_reg[1676]  ( .D(c[1684]), .CLK(clk), .RST(rst), .Q(sreg[1676]) );
  DFF \sreg_reg[1675]  ( .D(c[1683]), .CLK(clk), .RST(rst), .Q(sreg[1675]) );
  DFF \sreg_reg[1674]  ( .D(c[1682]), .CLK(clk), .RST(rst), .Q(sreg[1674]) );
  DFF \sreg_reg[1673]  ( .D(c[1681]), .CLK(clk), .RST(rst), .Q(sreg[1673]) );
  DFF \sreg_reg[1672]  ( .D(c[1680]), .CLK(clk), .RST(rst), .Q(sreg[1672]) );
  DFF \sreg_reg[1671]  ( .D(c[1679]), .CLK(clk), .RST(rst), .Q(sreg[1671]) );
  DFF \sreg_reg[1670]  ( .D(c[1678]), .CLK(clk), .RST(rst), .Q(sreg[1670]) );
  DFF \sreg_reg[1669]  ( .D(c[1677]), .CLK(clk), .RST(rst), .Q(sreg[1669]) );
  DFF \sreg_reg[1668]  ( .D(c[1676]), .CLK(clk), .RST(rst), .Q(sreg[1668]) );
  DFF \sreg_reg[1667]  ( .D(c[1675]), .CLK(clk), .RST(rst), .Q(sreg[1667]) );
  DFF \sreg_reg[1666]  ( .D(c[1674]), .CLK(clk), .RST(rst), .Q(sreg[1666]) );
  DFF \sreg_reg[1665]  ( .D(c[1673]), .CLK(clk), .RST(rst), .Q(sreg[1665]) );
  DFF \sreg_reg[1664]  ( .D(c[1672]), .CLK(clk), .RST(rst), .Q(sreg[1664]) );
  DFF \sreg_reg[1663]  ( .D(c[1671]), .CLK(clk), .RST(rst), .Q(sreg[1663]) );
  DFF \sreg_reg[1662]  ( .D(c[1670]), .CLK(clk), .RST(rst), .Q(sreg[1662]) );
  DFF \sreg_reg[1661]  ( .D(c[1669]), .CLK(clk), .RST(rst), .Q(sreg[1661]) );
  DFF \sreg_reg[1660]  ( .D(c[1668]), .CLK(clk), .RST(rst), .Q(sreg[1660]) );
  DFF \sreg_reg[1659]  ( .D(c[1667]), .CLK(clk), .RST(rst), .Q(sreg[1659]) );
  DFF \sreg_reg[1658]  ( .D(c[1666]), .CLK(clk), .RST(rst), .Q(sreg[1658]) );
  DFF \sreg_reg[1657]  ( .D(c[1665]), .CLK(clk), .RST(rst), .Q(sreg[1657]) );
  DFF \sreg_reg[1656]  ( .D(c[1664]), .CLK(clk), .RST(rst), .Q(sreg[1656]) );
  DFF \sreg_reg[1655]  ( .D(c[1663]), .CLK(clk), .RST(rst), .Q(sreg[1655]) );
  DFF \sreg_reg[1654]  ( .D(c[1662]), .CLK(clk), .RST(rst), .Q(sreg[1654]) );
  DFF \sreg_reg[1653]  ( .D(c[1661]), .CLK(clk), .RST(rst), .Q(sreg[1653]) );
  DFF \sreg_reg[1652]  ( .D(c[1660]), .CLK(clk), .RST(rst), .Q(sreg[1652]) );
  DFF \sreg_reg[1651]  ( .D(c[1659]), .CLK(clk), .RST(rst), .Q(sreg[1651]) );
  DFF \sreg_reg[1650]  ( .D(c[1658]), .CLK(clk), .RST(rst), .Q(sreg[1650]) );
  DFF \sreg_reg[1649]  ( .D(c[1657]), .CLK(clk), .RST(rst), .Q(sreg[1649]) );
  DFF \sreg_reg[1648]  ( .D(c[1656]), .CLK(clk), .RST(rst), .Q(sreg[1648]) );
  DFF \sreg_reg[1647]  ( .D(c[1655]), .CLK(clk), .RST(rst), .Q(sreg[1647]) );
  DFF \sreg_reg[1646]  ( .D(c[1654]), .CLK(clk), .RST(rst), .Q(sreg[1646]) );
  DFF \sreg_reg[1645]  ( .D(c[1653]), .CLK(clk), .RST(rst), .Q(sreg[1645]) );
  DFF \sreg_reg[1644]  ( .D(c[1652]), .CLK(clk), .RST(rst), .Q(sreg[1644]) );
  DFF \sreg_reg[1643]  ( .D(c[1651]), .CLK(clk), .RST(rst), .Q(sreg[1643]) );
  DFF \sreg_reg[1642]  ( .D(c[1650]), .CLK(clk), .RST(rst), .Q(sreg[1642]) );
  DFF \sreg_reg[1641]  ( .D(c[1649]), .CLK(clk), .RST(rst), .Q(sreg[1641]) );
  DFF \sreg_reg[1640]  ( .D(c[1648]), .CLK(clk), .RST(rst), .Q(sreg[1640]) );
  DFF \sreg_reg[1639]  ( .D(c[1647]), .CLK(clk), .RST(rst), .Q(sreg[1639]) );
  DFF \sreg_reg[1638]  ( .D(c[1646]), .CLK(clk), .RST(rst), .Q(sreg[1638]) );
  DFF \sreg_reg[1637]  ( .D(c[1645]), .CLK(clk), .RST(rst), .Q(sreg[1637]) );
  DFF \sreg_reg[1636]  ( .D(c[1644]), .CLK(clk), .RST(rst), .Q(sreg[1636]) );
  DFF \sreg_reg[1635]  ( .D(c[1643]), .CLK(clk), .RST(rst), .Q(sreg[1635]) );
  DFF \sreg_reg[1634]  ( .D(c[1642]), .CLK(clk), .RST(rst), .Q(sreg[1634]) );
  DFF \sreg_reg[1633]  ( .D(c[1641]), .CLK(clk), .RST(rst), .Q(sreg[1633]) );
  DFF \sreg_reg[1632]  ( .D(c[1640]), .CLK(clk), .RST(rst), .Q(sreg[1632]) );
  DFF \sreg_reg[1631]  ( .D(c[1639]), .CLK(clk), .RST(rst), .Q(sreg[1631]) );
  DFF \sreg_reg[1630]  ( .D(c[1638]), .CLK(clk), .RST(rst), .Q(sreg[1630]) );
  DFF \sreg_reg[1629]  ( .D(c[1637]), .CLK(clk), .RST(rst), .Q(sreg[1629]) );
  DFF \sreg_reg[1628]  ( .D(c[1636]), .CLK(clk), .RST(rst), .Q(sreg[1628]) );
  DFF \sreg_reg[1627]  ( .D(c[1635]), .CLK(clk), .RST(rst), .Q(sreg[1627]) );
  DFF \sreg_reg[1626]  ( .D(c[1634]), .CLK(clk), .RST(rst), .Q(sreg[1626]) );
  DFF \sreg_reg[1625]  ( .D(c[1633]), .CLK(clk), .RST(rst), .Q(sreg[1625]) );
  DFF \sreg_reg[1624]  ( .D(c[1632]), .CLK(clk), .RST(rst), .Q(sreg[1624]) );
  DFF \sreg_reg[1623]  ( .D(c[1631]), .CLK(clk), .RST(rst), .Q(sreg[1623]) );
  DFF \sreg_reg[1622]  ( .D(c[1630]), .CLK(clk), .RST(rst), .Q(sreg[1622]) );
  DFF \sreg_reg[1621]  ( .D(c[1629]), .CLK(clk), .RST(rst), .Q(sreg[1621]) );
  DFF \sreg_reg[1620]  ( .D(c[1628]), .CLK(clk), .RST(rst), .Q(sreg[1620]) );
  DFF \sreg_reg[1619]  ( .D(c[1627]), .CLK(clk), .RST(rst), .Q(sreg[1619]) );
  DFF \sreg_reg[1618]  ( .D(c[1626]), .CLK(clk), .RST(rst), .Q(sreg[1618]) );
  DFF \sreg_reg[1617]  ( .D(c[1625]), .CLK(clk), .RST(rst), .Q(sreg[1617]) );
  DFF \sreg_reg[1616]  ( .D(c[1624]), .CLK(clk), .RST(rst), .Q(sreg[1616]) );
  DFF \sreg_reg[1615]  ( .D(c[1623]), .CLK(clk), .RST(rst), .Q(sreg[1615]) );
  DFF \sreg_reg[1614]  ( .D(c[1622]), .CLK(clk), .RST(rst), .Q(sreg[1614]) );
  DFF \sreg_reg[1613]  ( .D(c[1621]), .CLK(clk), .RST(rst), .Q(sreg[1613]) );
  DFF \sreg_reg[1612]  ( .D(c[1620]), .CLK(clk), .RST(rst), .Q(sreg[1612]) );
  DFF \sreg_reg[1611]  ( .D(c[1619]), .CLK(clk), .RST(rst), .Q(sreg[1611]) );
  DFF \sreg_reg[1610]  ( .D(c[1618]), .CLK(clk), .RST(rst), .Q(sreg[1610]) );
  DFF \sreg_reg[1609]  ( .D(c[1617]), .CLK(clk), .RST(rst), .Q(sreg[1609]) );
  DFF \sreg_reg[1608]  ( .D(c[1616]), .CLK(clk), .RST(rst), .Q(sreg[1608]) );
  DFF \sreg_reg[1607]  ( .D(c[1615]), .CLK(clk), .RST(rst), .Q(sreg[1607]) );
  DFF \sreg_reg[1606]  ( .D(c[1614]), .CLK(clk), .RST(rst), .Q(sreg[1606]) );
  DFF \sreg_reg[1605]  ( .D(c[1613]), .CLK(clk), .RST(rst), .Q(sreg[1605]) );
  DFF \sreg_reg[1604]  ( .D(c[1612]), .CLK(clk), .RST(rst), .Q(sreg[1604]) );
  DFF \sreg_reg[1603]  ( .D(c[1611]), .CLK(clk), .RST(rst), .Q(sreg[1603]) );
  DFF \sreg_reg[1602]  ( .D(c[1610]), .CLK(clk), .RST(rst), .Q(sreg[1602]) );
  DFF \sreg_reg[1601]  ( .D(c[1609]), .CLK(clk), .RST(rst), .Q(sreg[1601]) );
  DFF \sreg_reg[1600]  ( .D(c[1608]), .CLK(clk), .RST(rst), .Q(sreg[1600]) );
  DFF \sreg_reg[1599]  ( .D(c[1607]), .CLK(clk), .RST(rst), .Q(sreg[1599]) );
  DFF \sreg_reg[1598]  ( .D(c[1606]), .CLK(clk), .RST(rst), .Q(sreg[1598]) );
  DFF \sreg_reg[1597]  ( .D(c[1605]), .CLK(clk), .RST(rst), .Q(sreg[1597]) );
  DFF \sreg_reg[1596]  ( .D(c[1604]), .CLK(clk), .RST(rst), .Q(sreg[1596]) );
  DFF \sreg_reg[1595]  ( .D(c[1603]), .CLK(clk), .RST(rst), .Q(sreg[1595]) );
  DFF \sreg_reg[1594]  ( .D(c[1602]), .CLK(clk), .RST(rst), .Q(sreg[1594]) );
  DFF \sreg_reg[1593]  ( .D(c[1601]), .CLK(clk), .RST(rst), .Q(sreg[1593]) );
  DFF \sreg_reg[1592]  ( .D(c[1600]), .CLK(clk), .RST(rst), .Q(sreg[1592]) );
  DFF \sreg_reg[1591]  ( .D(c[1599]), .CLK(clk), .RST(rst), .Q(sreg[1591]) );
  DFF \sreg_reg[1590]  ( .D(c[1598]), .CLK(clk), .RST(rst), .Q(sreg[1590]) );
  DFF \sreg_reg[1589]  ( .D(c[1597]), .CLK(clk), .RST(rst), .Q(sreg[1589]) );
  DFF \sreg_reg[1588]  ( .D(c[1596]), .CLK(clk), .RST(rst), .Q(sreg[1588]) );
  DFF \sreg_reg[1587]  ( .D(c[1595]), .CLK(clk), .RST(rst), .Q(sreg[1587]) );
  DFF \sreg_reg[1586]  ( .D(c[1594]), .CLK(clk), .RST(rst), .Q(sreg[1586]) );
  DFF \sreg_reg[1585]  ( .D(c[1593]), .CLK(clk), .RST(rst), .Q(sreg[1585]) );
  DFF \sreg_reg[1584]  ( .D(c[1592]), .CLK(clk), .RST(rst), .Q(sreg[1584]) );
  DFF \sreg_reg[1583]  ( .D(c[1591]), .CLK(clk), .RST(rst), .Q(sreg[1583]) );
  DFF \sreg_reg[1582]  ( .D(c[1590]), .CLK(clk), .RST(rst), .Q(sreg[1582]) );
  DFF \sreg_reg[1581]  ( .D(c[1589]), .CLK(clk), .RST(rst), .Q(sreg[1581]) );
  DFF \sreg_reg[1580]  ( .D(c[1588]), .CLK(clk), .RST(rst), .Q(sreg[1580]) );
  DFF \sreg_reg[1579]  ( .D(c[1587]), .CLK(clk), .RST(rst), .Q(sreg[1579]) );
  DFF \sreg_reg[1578]  ( .D(c[1586]), .CLK(clk), .RST(rst), .Q(sreg[1578]) );
  DFF \sreg_reg[1577]  ( .D(c[1585]), .CLK(clk), .RST(rst), .Q(sreg[1577]) );
  DFF \sreg_reg[1576]  ( .D(c[1584]), .CLK(clk), .RST(rst), .Q(sreg[1576]) );
  DFF \sreg_reg[1575]  ( .D(c[1583]), .CLK(clk), .RST(rst), .Q(sreg[1575]) );
  DFF \sreg_reg[1574]  ( .D(c[1582]), .CLK(clk), .RST(rst), .Q(sreg[1574]) );
  DFF \sreg_reg[1573]  ( .D(c[1581]), .CLK(clk), .RST(rst), .Q(sreg[1573]) );
  DFF \sreg_reg[1572]  ( .D(c[1580]), .CLK(clk), .RST(rst), .Q(sreg[1572]) );
  DFF \sreg_reg[1571]  ( .D(c[1579]), .CLK(clk), .RST(rst), .Q(sreg[1571]) );
  DFF \sreg_reg[1570]  ( .D(c[1578]), .CLK(clk), .RST(rst), .Q(sreg[1570]) );
  DFF \sreg_reg[1569]  ( .D(c[1577]), .CLK(clk), .RST(rst), .Q(sreg[1569]) );
  DFF \sreg_reg[1568]  ( .D(c[1576]), .CLK(clk), .RST(rst), .Q(sreg[1568]) );
  DFF \sreg_reg[1567]  ( .D(c[1575]), .CLK(clk), .RST(rst), .Q(sreg[1567]) );
  DFF \sreg_reg[1566]  ( .D(c[1574]), .CLK(clk), .RST(rst), .Q(sreg[1566]) );
  DFF \sreg_reg[1565]  ( .D(c[1573]), .CLK(clk), .RST(rst), .Q(sreg[1565]) );
  DFF \sreg_reg[1564]  ( .D(c[1572]), .CLK(clk), .RST(rst), .Q(sreg[1564]) );
  DFF \sreg_reg[1563]  ( .D(c[1571]), .CLK(clk), .RST(rst), .Q(sreg[1563]) );
  DFF \sreg_reg[1562]  ( .D(c[1570]), .CLK(clk), .RST(rst), .Q(sreg[1562]) );
  DFF \sreg_reg[1561]  ( .D(c[1569]), .CLK(clk), .RST(rst), .Q(sreg[1561]) );
  DFF \sreg_reg[1560]  ( .D(c[1568]), .CLK(clk), .RST(rst), .Q(sreg[1560]) );
  DFF \sreg_reg[1559]  ( .D(c[1567]), .CLK(clk), .RST(rst), .Q(sreg[1559]) );
  DFF \sreg_reg[1558]  ( .D(c[1566]), .CLK(clk), .RST(rst), .Q(sreg[1558]) );
  DFF \sreg_reg[1557]  ( .D(c[1565]), .CLK(clk), .RST(rst), .Q(sreg[1557]) );
  DFF \sreg_reg[1556]  ( .D(c[1564]), .CLK(clk), .RST(rst), .Q(sreg[1556]) );
  DFF \sreg_reg[1555]  ( .D(c[1563]), .CLK(clk), .RST(rst), .Q(sreg[1555]) );
  DFF \sreg_reg[1554]  ( .D(c[1562]), .CLK(clk), .RST(rst), .Q(sreg[1554]) );
  DFF \sreg_reg[1553]  ( .D(c[1561]), .CLK(clk), .RST(rst), .Q(sreg[1553]) );
  DFF \sreg_reg[1552]  ( .D(c[1560]), .CLK(clk), .RST(rst), .Q(sreg[1552]) );
  DFF \sreg_reg[1551]  ( .D(c[1559]), .CLK(clk), .RST(rst), .Q(sreg[1551]) );
  DFF \sreg_reg[1550]  ( .D(c[1558]), .CLK(clk), .RST(rst), .Q(sreg[1550]) );
  DFF \sreg_reg[1549]  ( .D(c[1557]), .CLK(clk), .RST(rst), .Q(sreg[1549]) );
  DFF \sreg_reg[1548]  ( .D(c[1556]), .CLK(clk), .RST(rst), .Q(sreg[1548]) );
  DFF \sreg_reg[1547]  ( .D(c[1555]), .CLK(clk), .RST(rst), .Q(sreg[1547]) );
  DFF \sreg_reg[1546]  ( .D(c[1554]), .CLK(clk), .RST(rst), .Q(sreg[1546]) );
  DFF \sreg_reg[1545]  ( .D(c[1553]), .CLK(clk), .RST(rst), .Q(sreg[1545]) );
  DFF \sreg_reg[1544]  ( .D(c[1552]), .CLK(clk), .RST(rst), .Q(sreg[1544]) );
  DFF \sreg_reg[1543]  ( .D(c[1551]), .CLK(clk), .RST(rst), .Q(sreg[1543]) );
  DFF \sreg_reg[1542]  ( .D(c[1550]), .CLK(clk), .RST(rst), .Q(sreg[1542]) );
  DFF \sreg_reg[1541]  ( .D(c[1549]), .CLK(clk), .RST(rst), .Q(sreg[1541]) );
  DFF \sreg_reg[1540]  ( .D(c[1548]), .CLK(clk), .RST(rst), .Q(sreg[1540]) );
  DFF \sreg_reg[1539]  ( .D(c[1547]), .CLK(clk), .RST(rst), .Q(sreg[1539]) );
  DFF \sreg_reg[1538]  ( .D(c[1546]), .CLK(clk), .RST(rst), .Q(sreg[1538]) );
  DFF \sreg_reg[1537]  ( .D(c[1545]), .CLK(clk), .RST(rst), .Q(sreg[1537]) );
  DFF \sreg_reg[1536]  ( .D(c[1544]), .CLK(clk), .RST(rst), .Q(sreg[1536]) );
  DFF \sreg_reg[1535]  ( .D(c[1543]), .CLK(clk), .RST(rst), .Q(sreg[1535]) );
  DFF \sreg_reg[1534]  ( .D(c[1542]), .CLK(clk), .RST(rst), .Q(sreg[1534]) );
  DFF \sreg_reg[1533]  ( .D(c[1541]), .CLK(clk), .RST(rst), .Q(sreg[1533]) );
  DFF \sreg_reg[1532]  ( .D(c[1540]), .CLK(clk), .RST(rst), .Q(sreg[1532]) );
  DFF \sreg_reg[1531]  ( .D(c[1539]), .CLK(clk), .RST(rst), .Q(sreg[1531]) );
  DFF \sreg_reg[1530]  ( .D(c[1538]), .CLK(clk), .RST(rst), .Q(sreg[1530]) );
  DFF \sreg_reg[1529]  ( .D(c[1537]), .CLK(clk), .RST(rst), .Q(sreg[1529]) );
  DFF \sreg_reg[1528]  ( .D(c[1536]), .CLK(clk), .RST(rst), .Q(sreg[1528]) );
  DFF \sreg_reg[1527]  ( .D(c[1535]), .CLK(clk), .RST(rst), .Q(sreg[1527]) );
  DFF \sreg_reg[1526]  ( .D(c[1534]), .CLK(clk), .RST(rst), .Q(sreg[1526]) );
  DFF \sreg_reg[1525]  ( .D(c[1533]), .CLK(clk), .RST(rst), .Q(sreg[1525]) );
  DFF \sreg_reg[1524]  ( .D(c[1532]), .CLK(clk), .RST(rst), .Q(sreg[1524]) );
  DFF \sreg_reg[1523]  ( .D(c[1531]), .CLK(clk), .RST(rst), .Q(sreg[1523]) );
  DFF \sreg_reg[1522]  ( .D(c[1530]), .CLK(clk), .RST(rst), .Q(sreg[1522]) );
  DFF \sreg_reg[1521]  ( .D(c[1529]), .CLK(clk), .RST(rst), .Q(sreg[1521]) );
  DFF \sreg_reg[1520]  ( .D(c[1528]), .CLK(clk), .RST(rst), .Q(sreg[1520]) );
  DFF \sreg_reg[1519]  ( .D(c[1527]), .CLK(clk), .RST(rst), .Q(sreg[1519]) );
  DFF \sreg_reg[1518]  ( .D(c[1526]), .CLK(clk), .RST(rst), .Q(sreg[1518]) );
  DFF \sreg_reg[1517]  ( .D(c[1525]), .CLK(clk), .RST(rst), .Q(sreg[1517]) );
  DFF \sreg_reg[1516]  ( .D(c[1524]), .CLK(clk), .RST(rst), .Q(sreg[1516]) );
  DFF \sreg_reg[1515]  ( .D(c[1523]), .CLK(clk), .RST(rst), .Q(sreg[1515]) );
  DFF \sreg_reg[1514]  ( .D(c[1522]), .CLK(clk), .RST(rst), .Q(sreg[1514]) );
  DFF \sreg_reg[1513]  ( .D(c[1521]), .CLK(clk), .RST(rst), .Q(sreg[1513]) );
  DFF \sreg_reg[1512]  ( .D(c[1520]), .CLK(clk), .RST(rst), .Q(sreg[1512]) );
  DFF \sreg_reg[1511]  ( .D(c[1519]), .CLK(clk), .RST(rst), .Q(sreg[1511]) );
  DFF \sreg_reg[1510]  ( .D(c[1518]), .CLK(clk), .RST(rst), .Q(sreg[1510]) );
  DFF \sreg_reg[1509]  ( .D(c[1517]), .CLK(clk), .RST(rst), .Q(sreg[1509]) );
  DFF \sreg_reg[1508]  ( .D(c[1516]), .CLK(clk), .RST(rst), .Q(sreg[1508]) );
  DFF \sreg_reg[1507]  ( .D(c[1515]), .CLK(clk), .RST(rst), .Q(sreg[1507]) );
  DFF \sreg_reg[1506]  ( .D(c[1514]), .CLK(clk), .RST(rst), .Q(sreg[1506]) );
  DFF \sreg_reg[1505]  ( .D(c[1513]), .CLK(clk), .RST(rst), .Q(sreg[1505]) );
  DFF \sreg_reg[1504]  ( .D(c[1512]), .CLK(clk), .RST(rst), .Q(sreg[1504]) );
  DFF \sreg_reg[1503]  ( .D(c[1511]), .CLK(clk), .RST(rst), .Q(sreg[1503]) );
  DFF \sreg_reg[1502]  ( .D(c[1510]), .CLK(clk), .RST(rst), .Q(sreg[1502]) );
  DFF \sreg_reg[1501]  ( .D(c[1509]), .CLK(clk), .RST(rst), .Q(sreg[1501]) );
  DFF \sreg_reg[1500]  ( .D(c[1508]), .CLK(clk), .RST(rst), .Q(sreg[1500]) );
  DFF \sreg_reg[1499]  ( .D(c[1507]), .CLK(clk), .RST(rst), .Q(sreg[1499]) );
  DFF \sreg_reg[1498]  ( .D(c[1506]), .CLK(clk), .RST(rst), .Q(sreg[1498]) );
  DFF \sreg_reg[1497]  ( .D(c[1505]), .CLK(clk), .RST(rst), .Q(sreg[1497]) );
  DFF \sreg_reg[1496]  ( .D(c[1504]), .CLK(clk), .RST(rst), .Q(sreg[1496]) );
  DFF \sreg_reg[1495]  ( .D(c[1503]), .CLK(clk), .RST(rst), .Q(sreg[1495]) );
  DFF \sreg_reg[1494]  ( .D(c[1502]), .CLK(clk), .RST(rst), .Q(sreg[1494]) );
  DFF \sreg_reg[1493]  ( .D(c[1501]), .CLK(clk), .RST(rst), .Q(sreg[1493]) );
  DFF \sreg_reg[1492]  ( .D(c[1500]), .CLK(clk), .RST(rst), .Q(sreg[1492]) );
  DFF \sreg_reg[1491]  ( .D(c[1499]), .CLK(clk), .RST(rst), .Q(sreg[1491]) );
  DFF \sreg_reg[1490]  ( .D(c[1498]), .CLK(clk), .RST(rst), .Q(sreg[1490]) );
  DFF \sreg_reg[1489]  ( .D(c[1497]), .CLK(clk), .RST(rst), .Q(sreg[1489]) );
  DFF \sreg_reg[1488]  ( .D(c[1496]), .CLK(clk), .RST(rst), .Q(sreg[1488]) );
  DFF \sreg_reg[1487]  ( .D(c[1495]), .CLK(clk), .RST(rst), .Q(sreg[1487]) );
  DFF \sreg_reg[1486]  ( .D(c[1494]), .CLK(clk), .RST(rst), .Q(sreg[1486]) );
  DFF \sreg_reg[1485]  ( .D(c[1493]), .CLK(clk), .RST(rst), .Q(sreg[1485]) );
  DFF \sreg_reg[1484]  ( .D(c[1492]), .CLK(clk), .RST(rst), .Q(sreg[1484]) );
  DFF \sreg_reg[1483]  ( .D(c[1491]), .CLK(clk), .RST(rst), .Q(sreg[1483]) );
  DFF \sreg_reg[1482]  ( .D(c[1490]), .CLK(clk), .RST(rst), .Q(sreg[1482]) );
  DFF \sreg_reg[1481]  ( .D(c[1489]), .CLK(clk), .RST(rst), .Q(sreg[1481]) );
  DFF \sreg_reg[1480]  ( .D(c[1488]), .CLK(clk), .RST(rst), .Q(sreg[1480]) );
  DFF \sreg_reg[1479]  ( .D(c[1487]), .CLK(clk), .RST(rst), .Q(sreg[1479]) );
  DFF \sreg_reg[1478]  ( .D(c[1486]), .CLK(clk), .RST(rst), .Q(sreg[1478]) );
  DFF \sreg_reg[1477]  ( .D(c[1485]), .CLK(clk), .RST(rst), .Q(sreg[1477]) );
  DFF \sreg_reg[1476]  ( .D(c[1484]), .CLK(clk), .RST(rst), .Q(sreg[1476]) );
  DFF \sreg_reg[1475]  ( .D(c[1483]), .CLK(clk), .RST(rst), .Q(sreg[1475]) );
  DFF \sreg_reg[1474]  ( .D(c[1482]), .CLK(clk), .RST(rst), .Q(sreg[1474]) );
  DFF \sreg_reg[1473]  ( .D(c[1481]), .CLK(clk), .RST(rst), .Q(sreg[1473]) );
  DFF \sreg_reg[1472]  ( .D(c[1480]), .CLK(clk), .RST(rst), .Q(sreg[1472]) );
  DFF \sreg_reg[1471]  ( .D(c[1479]), .CLK(clk), .RST(rst), .Q(sreg[1471]) );
  DFF \sreg_reg[1470]  ( .D(c[1478]), .CLK(clk), .RST(rst), .Q(sreg[1470]) );
  DFF \sreg_reg[1469]  ( .D(c[1477]), .CLK(clk), .RST(rst), .Q(sreg[1469]) );
  DFF \sreg_reg[1468]  ( .D(c[1476]), .CLK(clk), .RST(rst), .Q(sreg[1468]) );
  DFF \sreg_reg[1467]  ( .D(c[1475]), .CLK(clk), .RST(rst), .Q(sreg[1467]) );
  DFF \sreg_reg[1466]  ( .D(c[1474]), .CLK(clk), .RST(rst), .Q(sreg[1466]) );
  DFF \sreg_reg[1465]  ( .D(c[1473]), .CLK(clk), .RST(rst), .Q(sreg[1465]) );
  DFF \sreg_reg[1464]  ( .D(c[1472]), .CLK(clk), .RST(rst), .Q(sreg[1464]) );
  DFF \sreg_reg[1463]  ( .D(c[1471]), .CLK(clk), .RST(rst), .Q(sreg[1463]) );
  DFF \sreg_reg[1462]  ( .D(c[1470]), .CLK(clk), .RST(rst), .Q(sreg[1462]) );
  DFF \sreg_reg[1461]  ( .D(c[1469]), .CLK(clk), .RST(rst), .Q(sreg[1461]) );
  DFF \sreg_reg[1460]  ( .D(c[1468]), .CLK(clk), .RST(rst), .Q(sreg[1460]) );
  DFF \sreg_reg[1459]  ( .D(c[1467]), .CLK(clk), .RST(rst), .Q(sreg[1459]) );
  DFF \sreg_reg[1458]  ( .D(c[1466]), .CLK(clk), .RST(rst), .Q(sreg[1458]) );
  DFF \sreg_reg[1457]  ( .D(c[1465]), .CLK(clk), .RST(rst), .Q(sreg[1457]) );
  DFF \sreg_reg[1456]  ( .D(c[1464]), .CLK(clk), .RST(rst), .Q(sreg[1456]) );
  DFF \sreg_reg[1455]  ( .D(c[1463]), .CLK(clk), .RST(rst), .Q(sreg[1455]) );
  DFF \sreg_reg[1454]  ( .D(c[1462]), .CLK(clk), .RST(rst), .Q(sreg[1454]) );
  DFF \sreg_reg[1453]  ( .D(c[1461]), .CLK(clk), .RST(rst), .Q(sreg[1453]) );
  DFF \sreg_reg[1452]  ( .D(c[1460]), .CLK(clk), .RST(rst), .Q(sreg[1452]) );
  DFF \sreg_reg[1451]  ( .D(c[1459]), .CLK(clk), .RST(rst), .Q(sreg[1451]) );
  DFF \sreg_reg[1450]  ( .D(c[1458]), .CLK(clk), .RST(rst), .Q(sreg[1450]) );
  DFF \sreg_reg[1449]  ( .D(c[1457]), .CLK(clk), .RST(rst), .Q(sreg[1449]) );
  DFF \sreg_reg[1448]  ( .D(c[1456]), .CLK(clk), .RST(rst), .Q(sreg[1448]) );
  DFF \sreg_reg[1447]  ( .D(c[1455]), .CLK(clk), .RST(rst), .Q(sreg[1447]) );
  DFF \sreg_reg[1446]  ( .D(c[1454]), .CLK(clk), .RST(rst), .Q(sreg[1446]) );
  DFF \sreg_reg[1445]  ( .D(c[1453]), .CLK(clk), .RST(rst), .Q(sreg[1445]) );
  DFF \sreg_reg[1444]  ( .D(c[1452]), .CLK(clk), .RST(rst), .Q(sreg[1444]) );
  DFF \sreg_reg[1443]  ( .D(c[1451]), .CLK(clk), .RST(rst), .Q(sreg[1443]) );
  DFF \sreg_reg[1442]  ( .D(c[1450]), .CLK(clk), .RST(rst), .Q(sreg[1442]) );
  DFF \sreg_reg[1441]  ( .D(c[1449]), .CLK(clk), .RST(rst), .Q(sreg[1441]) );
  DFF \sreg_reg[1440]  ( .D(c[1448]), .CLK(clk), .RST(rst), .Q(sreg[1440]) );
  DFF \sreg_reg[1439]  ( .D(c[1447]), .CLK(clk), .RST(rst), .Q(sreg[1439]) );
  DFF \sreg_reg[1438]  ( .D(c[1446]), .CLK(clk), .RST(rst), .Q(sreg[1438]) );
  DFF \sreg_reg[1437]  ( .D(c[1445]), .CLK(clk), .RST(rst), .Q(sreg[1437]) );
  DFF \sreg_reg[1436]  ( .D(c[1444]), .CLK(clk), .RST(rst), .Q(sreg[1436]) );
  DFF \sreg_reg[1435]  ( .D(c[1443]), .CLK(clk), .RST(rst), .Q(sreg[1435]) );
  DFF \sreg_reg[1434]  ( .D(c[1442]), .CLK(clk), .RST(rst), .Q(sreg[1434]) );
  DFF \sreg_reg[1433]  ( .D(c[1441]), .CLK(clk), .RST(rst), .Q(sreg[1433]) );
  DFF \sreg_reg[1432]  ( .D(c[1440]), .CLK(clk), .RST(rst), .Q(sreg[1432]) );
  DFF \sreg_reg[1431]  ( .D(c[1439]), .CLK(clk), .RST(rst), .Q(sreg[1431]) );
  DFF \sreg_reg[1430]  ( .D(c[1438]), .CLK(clk), .RST(rst), .Q(sreg[1430]) );
  DFF \sreg_reg[1429]  ( .D(c[1437]), .CLK(clk), .RST(rst), .Q(sreg[1429]) );
  DFF \sreg_reg[1428]  ( .D(c[1436]), .CLK(clk), .RST(rst), .Q(sreg[1428]) );
  DFF \sreg_reg[1427]  ( .D(c[1435]), .CLK(clk), .RST(rst), .Q(sreg[1427]) );
  DFF \sreg_reg[1426]  ( .D(c[1434]), .CLK(clk), .RST(rst), .Q(sreg[1426]) );
  DFF \sreg_reg[1425]  ( .D(c[1433]), .CLK(clk), .RST(rst), .Q(sreg[1425]) );
  DFF \sreg_reg[1424]  ( .D(c[1432]), .CLK(clk), .RST(rst), .Q(sreg[1424]) );
  DFF \sreg_reg[1423]  ( .D(c[1431]), .CLK(clk), .RST(rst), .Q(sreg[1423]) );
  DFF \sreg_reg[1422]  ( .D(c[1430]), .CLK(clk), .RST(rst), .Q(sreg[1422]) );
  DFF \sreg_reg[1421]  ( .D(c[1429]), .CLK(clk), .RST(rst), .Q(sreg[1421]) );
  DFF \sreg_reg[1420]  ( .D(c[1428]), .CLK(clk), .RST(rst), .Q(sreg[1420]) );
  DFF \sreg_reg[1419]  ( .D(c[1427]), .CLK(clk), .RST(rst), .Q(sreg[1419]) );
  DFF \sreg_reg[1418]  ( .D(c[1426]), .CLK(clk), .RST(rst), .Q(sreg[1418]) );
  DFF \sreg_reg[1417]  ( .D(c[1425]), .CLK(clk), .RST(rst), .Q(sreg[1417]) );
  DFF \sreg_reg[1416]  ( .D(c[1424]), .CLK(clk), .RST(rst), .Q(sreg[1416]) );
  DFF \sreg_reg[1415]  ( .D(c[1423]), .CLK(clk), .RST(rst), .Q(sreg[1415]) );
  DFF \sreg_reg[1414]  ( .D(c[1422]), .CLK(clk), .RST(rst), .Q(sreg[1414]) );
  DFF \sreg_reg[1413]  ( .D(c[1421]), .CLK(clk), .RST(rst), .Q(sreg[1413]) );
  DFF \sreg_reg[1412]  ( .D(c[1420]), .CLK(clk), .RST(rst), .Q(sreg[1412]) );
  DFF \sreg_reg[1411]  ( .D(c[1419]), .CLK(clk), .RST(rst), .Q(sreg[1411]) );
  DFF \sreg_reg[1410]  ( .D(c[1418]), .CLK(clk), .RST(rst), .Q(sreg[1410]) );
  DFF \sreg_reg[1409]  ( .D(c[1417]), .CLK(clk), .RST(rst), .Q(sreg[1409]) );
  DFF \sreg_reg[1408]  ( .D(c[1416]), .CLK(clk), .RST(rst), .Q(sreg[1408]) );
  DFF \sreg_reg[1407]  ( .D(c[1415]), .CLK(clk), .RST(rst), .Q(sreg[1407]) );
  DFF \sreg_reg[1406]  ( .D(c[1414]), .CLK(clk), .RST(rst), .Q(sreg[1406]) );
  DFF \sreg_reg[1405]  ( .D(c[1413]), .CLK(clk), .RST(rst), .Q(sreg[1405]) );
  DFF \sreg_reg[1404]  ( .D(c[1412]), .CLK(clk), .RST(rst), .Q(sreg[1404]) );
  DFF \sreg_reg[1403]  ( .D(c[1411]), .CLK(clk), .RST(rst), .Q(sreg[1403]) );
  DFF \sreg_reg[1402]  ( .D(c[1410]), .CLK(clk), .RST(rst), .Q(sreg[1402]) );
  DFF \sreg_reg[1401]  ( .D(c[1409]), .CLK(clk), .RST(rst), .Q(sreg[1401]) );
  DFF \sreg_reg[1400]  ( .D(c[1408]), .CLK(clk), .RST(rst), .Q(sreg[1400]) );
  DFF \sreg_reg[1399]  ( .D(c[1407]), .CLK(clk), .RST(rst), .Q(sreg[1399]) );
  DFF \sreg_reg[1398]  ( .D(c[1406]), .CLK(clk), .RST(rst), .Q(sreg[1398]) );
  DFF \sreg_reg[1397]  ( .D(c[1405]), .CLK(clk), .RST(rst), .Q(sreg[1397]) );
  DFF \sreg_reg[1396]  ( .D(c[1404]), .CLK(clk), .RST(rst), .Q(sreg[1396]) );
  DFF \sreg_reg[1395]  ( .D(c[1403]), .CLK(clk), .RST(rst), .Q(sreg[1395]) );
  DFF \sreg_reg[1394]  ( .D(c[1402]), .CLK(clk), .RST(rst), .Q(sreg[1394]) );
  DFF \sreg_reg[1393]  ( .D(c[1401]), .CLK(clk), .RST(rst), .Q(sreg[1393]) );
  DFF \sreg_reg[1392]  ( .D(c[1400]), .CLK(clk), .RST(rst), .Q(sreg[1392]) );
  DFF \sreg_reg[1391]  ( .D(c[1399]), .CLK(clk), .RST(rst), .Q(sreg[1391]) );
  DFF \sreg_reg[1390]  ( .D(c[1398]), .CLK(clk), .RST(rst), .Q(sreg[1390]) );
  DFF \sreg_reg[1389]  ( .D(c[1397]), .CLK(clk), .RST(rst), .Q(sreg[1389]) );
  DFF \sreg_reg[1388]  ( .D(c[1396]), .CLK(clk), .RST(rst), .Q(sreg[1388]) );
  DFF \sreg_reg[1387]  ( .D(c[1395]), .CLK(clk), .RST(rst), .Q(sreg[1387]) );
  DFF \sreg_reg[1386]  ( .D(c[1394]), .CLK(clk), .RST(rst), .Q(sreg[1386]) );
  DFF \sreg_reg[1385]  ( .D(c[1393]), .CLK(clk), .RST(rst), .Q(sreg[1385]) );
  DFF \sreg_reg[1384]  ( .D(c[1392]), .CLK(clk), .RST(rst), .Q(sreg[1384]) );
  DFF \sreg_reg[1383]  ( .D(c[1391]), .CLK(clk), .RST(rst), .Q(sreg[1383]) );
  DFF \sreg_reg[1382]  ( .D(c[1390]), .CLK(clk), .RST(rst), .Q(sreg[1382]) );
  DFF \sreg_reg[1381]  ( .D(c[1389]), .CLK(clk), .RST(rst), .Q(sreg[1381]) );
  DFF \sreg_reg[1380]  ( .D(c[1388]), .CLK(clk), .RST(rst), .Q(sreg[1380]) );
  DFF \sreg_reg[1379]  ( .D(c[1387]), .CLK(clk), .RST(rst), .Q(sreg[1379]) );
  DFF \sreg_reg[1378]  ( .D(c[1386]), .CLK(clk), .RST(rst), .Q(sreg[1378]) );
  DFF \sreg_reg[1377]  ( .D(c[1385]), .CLK(clk), .RST(rst), .Q(sreg[1377]) );
  DFF \sreg_reg[1376]  ( .D(c[1384]), .CLK(clk), .RST(rst), .Q(sreg[1376]) );
  DFF \sreg_reg[1375]  ( .D(c[1383]), .CLK(clk), .RST(rst), .Q(sreg[1375]) );
  DFF \sreg_reg[1374]  ( .D(c[1382]), .CLK(clk), .RST(rst), .Q(sreg[1374]) );
  DFF \sreg_reg[1373]  ( .D(c[1381]), .CLK(clk), .RST(rst), .Q(sreg[1373]) );
  DFF \sreg_reg[1372]  ( .D(c[1380]), .CLK(clk), .RST(rst), .Q(sreg[1372]) );
  DFF \sreg_reg[1371]  ( .D(c[1379]), .CLK(clk), .RST(rst), .Q(sreg[1371]) );
  DFF \sreg_reg[1370]  ( .D(c[1378]), .CLK(clk), .RST(rst), .Q(sreg[1370]) );
  DFF \sreg_reg[1369]  ( .D(c[1377]), .CLK(clk), .RST(rst), .Q(sreg[1369]) );
  DFF \sreg_reg[1368]  ( .D(c[1376]), .CLK(clk), .RST(rst), .Q(sreg[1368]) );
  DFF \sreg_reg[1367]  ( .D(c[1375]), .CLK(clk), .RST(rst), .Q(sreg[1367]) );
  DFF \sreg_reg[1366]  ( .D(c[1374]), .CLK(clk), .RST(rst), .Q(sreg[1366]) );
  DFF \sreg_reg[1365]  ( .D(c[1373]), .CLK(clk), .RST(rst), .Q(sreg[1365]) );
  DFF \sreg_reg[1364]  ( .D(c[1372]), .CLK(clk), .RST(rst), .Q(sreg[1364]) );
  DFF \sreg_reg[1363]  ( .D(c[1371]), .CLK(clk), .RST(rst), .Q(sreg[1363]) );
  DFF \sreg_reg[1362]  ( .D(c[1370]), .CLK(clk), .RST(rst), .Q(sreg[1362]) );
  DFF \sreg_reg[1361]  ( .D(c[1369]), .CLK(clk), .RST(rst), .Q(sreg[1361]) );
  DFF \sreg_reg[1360]  ( .D(c[1368]), .CLK(clk), .RST(rst), .Q(sreg[1360]) );
  DFF \sreg_reg[1359]  ( .D(c[1367]), .CLK(clk), .RST(rst), .Q(sreg[1359]) );
  DFF \sreg_reg[1358]  ( .D(c[1366]), .CLK(clk), .RST(rst), .Q(sreg[1358]) );
  DFF \sreg_reg[1357]  ( .D(c[1365]), .CLK(clk), .RST(rst), .Q(sreg[1357]) );
  DFF \sreg_reg[1356]  ( .D(c[1364]), .CLK(clk), .RST(rst), .Q(sreg[1356]) );
  DFF \sreg_reg[1355]  ( .D(c[1363]), .CLK(clk), .RST(rst), .Q(sreg[1355]) );
  DFF \sreg_reg[1354]  ( .D(c[1362]), .CLK(clk), .RST(rst), .Q(sreg[1354]) );
  DFF \sreg_reg[1353]  ( .D(c[1361]), .CLK(clk), .RST(rst), .Q(sreg[1353]) );
  DFF \sreg_reg[1352]  ( .D(c[1360]), .CLK(clk), .RST(rst), .Q(sreg[1352]) );
  DFF \sreg_reg[1351]  ( .D(c[1359]), .CLK(clk), .RST(rst), .Q(sreg[1351]) );
  DFF \sreg_reg[1350]  ( .D(c[1358]), .CLK(clk), .RST(rst), .Q(sreg[1350]) );
  DFF \sreg_reg[1349]  ( .D(c[1357]), .CLK(clk), .RST(rst), .Q(sreg[1349]) );
  DFF \sreg_reg[1348]  ( .D(c[1356]), .CLK(clk), .RST(rst), .Q(sreg[1348]) );
  DFF \sreg_reg[1347]  ( .D(c[1355]), .CLK(clk), .RST(rst), .Q(sreg[1347]) );
  DFF \sreg_reg[1346]  ( .D(c[1354]), .CLK(clk), .RST(rst), .Q(sreg[1346]) );
  DFF \sreg_reg[1345]  ( .D(c[1353]), .CLK(clk), .RST(rst), .Q(sreg[1345]) );
  DFF \sreg_reg[1344]  ( .D(c[1352]), .CLK(clk), .RST(rst), .Q(sreg[1344]) );
  DFF \sreg_reg[1343]  ( .D(c[1351]), .CLK(clk), .RST(rst), .Q(sreg[1343]) );
  DFF \sreg_reg[1342]  ( .D(c[1350]), .CLK(clk), .RST(rst), .Q(sreg[1342]) );
  DFF \sreg_reg[1341]  ( .D(c[1349]), .CLK(clk), .RST(rst), .Q(sreg[1341]) );
  DFF \sreg_reg[1340]  ( .D(c[1348]), .CLK(clk), .RST(rst), .Q(sreg[1340]) );
  DFF \sreg_reg[1339]  ( .D(c[1347]), .CLK(clk), .RST(rst), .Q(sreg[1339]) );
  DFF \sreg_reg[1338]  ( .D(c[1346]), .CLK(clk), .RST(rst), .Q(sreg[1338]) );
  DFF \sreg_reg[1337]  ( .D(c[1345]), .CLK(clk), .RST(rst), .Q(sreg[1337]) );
  DFF \sreg_reg[1336]  ( .D(c[1344]), .CLK(clk), .RST(rst), .Q(sreg[1336]) );
  DFF \sreg_reg[1335]  ( .D(c[1343]), .CLK(clk), .RST(rst), .Q(sreg[1335]) );
  DFF \sreg_reg[1334]  ( .D(c[1342]), .CLK(clk), .RST(rst), .Q(sreg[1334]) );
  DFF \sreg_reg[1333]  ( .D(c[1341]), .CLK(clk), .RST(rst), .Q(sreg[1333]) );
  DFF \sreg_reg[1332]  ( .D(c[1340]), .CLK(clk), .RST(rst), .Q(sreg[1332]) );
  DFF \sreg_reg[1331]  ( .D(c[1339]), .CLK(clk), .RST(rst), .Q(sreg[1331]) );
  DFF \sreg_reg[1330]  ( .D(c[1338]), .CLK(clk), .RST(rst), .Q(sreg[1330]) );
  DFF \sreg_reg[1329]  ( .D(c[1337]), .CLK(clk), .RST(rst), .Q(sreg[1329]) );
  DFF \sreg_reg[1328]  ( .D(c[1336]), .CLK(clk), .RST(rst), .Q(sreg[1328]) );
  DFF \sreg_reg[1327]  ( .D(c[1335]), .CLK(clk), .RST(rst), .Q(sreg[1327]) );
  DFF \sreg_reg[1326]  ( .D(c[1334]), .CLK(clk), .RST(rst), .Q(sreg[1326]) );
  DFF \sreg_reg[1325]  ( .D(c[1333]), .CLK(clk), .RST(rst), .Q(sreg[1325]) );
  DFF \sreg_reg[1324]  ( .D(c[1332]), .CLK(clk), .RST(rst), .Q(sreg[1324]) );
  DFF \sreg_reg[1323]  ( .D(c[1331]), .CLK(clk), .RST(rst), .Q(sreg[1323]) );
  DFF \sreg_reg[1322]  ( .D(c[1330]), .CLK(clk), .RST(rst), .Q(sreg[1322]) );
  DFF \sreg_reg[1321]  ( .D(c[1329]), .CLK(clk), .RST(rst), .Q(sreg[1321]) );
  DFF \sreg_reg[1320]  ( .D(c[1328]), .CLK(clk), .RST(rst), .Q(sreg[1320]) );
  DFF \sreg_reg[1319]  ( .D(c[1327]), .CLK(clk), .RST(rst), .Q(sreg[1319]) );
  DFF \sreg_reg[1318]  ( .D(c[1326]), .CLK(clk), .RST(rst), .Q(sreg[1318]) );
  DFF \sreg_reg[1317]  ( .D(c[1325]), .CLK(clk), .RST(rst), .Q(sreg[1317]) );
  DFF \sreg_reg[1316]  ( .D(c[1324]), .CLK(clk), .RST(rst), .Q(sreg[1316]) );
  DFF \sreg_reg[1315]  ( .D(c[1323]), .CLK(clk), .RST(rst), .Q(sreg[1315]) );
  DFF \sreg_reg[1314]  ( .D(c[1322]), .CLK(clk), .RST(rst), .Q(sreg[1314]) );
  DFF \sreg_reg[1313]  ( .D(c[1321]), .CLK(clk), .RST(rst), .Q(sreg[1313]) );
  DFF \sreg_reg[1312]  ( .D(c[1320]), .CLK(clk), .RST(rst), .Q(sreg[1312]) );
  DFF \sreg_reg[1311]  ( .D(c[1319]), .CLK(clk), .RST(rst), .Q(sreg[1311]) );
  DFF \sreg_reg[1310]  ( .D(c[1318]), .CLK(clk), .RST(rst), .Q(sreg[1310]) );
  DFF \sreg_reg[1309]  ( .D(c[1317]), .CLK(clk), .RST(rst), .Q(sreg[1309]) );
  DFF \sreg_reg[1308]  ( .D(c[1316]), .CLK(clk), .RST(rst), .Q(sreg[1308]) );
  DFF \sreg_reg[1307]  ( .D(c[1315]), .CLK(clk), .RST(rst), .Q(sreg[1307]) );
  DFF \sreg_reg[1306]  ( .D(c[1314]), .CLK(clk), .RST(rst), .Q(sreg[1306]) );
  DFF \sreg_reg[1305]  ( .D(c[1313]), .CLK(clk), .RST(rst), .Q(sreg[1305]) );
  DFF \sreg_reg[1304]  ( .D(c[1312]), .CLK(clk), .RST(rst), .Q(sreg[1304]) );
  DFF \sreg_reg[1303]  ( .D(c[1311]), .CLK(clk), .RST(rst), .Q(sreg[1303]) );
  DFF \sreg_reg[1302]  ( .D(c[1310]), .CLK(clk), .RST(rst), .Q(sreg[1302]) );
  DFF \sreg_reg[1301]  ( .D(c[1309]), .CLK(clk), .RST(rst), .Q(sreg[1301]) );
  DFF \sreg_reg[1300]  ( .D(c[1308]), .CLK(clk), .RST(rst), .Q(sreg[1300]) );
  DFF \sreg_reg[1299]  ( .D(c[1307]), .CLK(clk), .RST(rst), .Q(sreg[1299]) );
  DFF \sreg_reg[1298]  ( .D(c[1306]), .CLK(clk), .RST(rst), .Q(sreg[1298]) );
  DFF \sreg_reg[1297]  ( .D(c[1305]), .CLK(clk), .RST(rst), .Q(sreg[1297]) );
  DFF \sreg_reg[1296]  ( .D(c[1304]), .CLK(clk), .RST(rst), .Q(sreg[1296]) );
  DFF \sreg_reg[1295]  ( .D(c[1303]), .CLK(clk), .RST(rst), .Q(sreg[1295]) );
  DFF \sreg_reg[1294]  ( .D(c[1302]), .CLK(clk), .RST(rst), .Q(sreg[1294]) );
  DFF \sreg_reg[1293]  ( .D(c[1301]), .CLK(clk), .RST(rst), .Q(sreg[1293]) );
  DFF \sreg_reg[1292]  ( .D(c[1300]), .CLK(clk), .RST(rst), .Q(sreg[1292]) );
  DFF \sreg_reg[1291]  ( .D(c[1299]), .CLK(clk), .RST(rst), .Q(sreg[1291]) );
  DFF \sreg_reg[1290]  ( .D(c[1298]), .CLK(clk), .RST(rst), .Q(sreg[1290]) );
  DFF \sreg_reg[1289]  ( .D(c[1297]), .CLK(clk), .RST(rst), .Q(sreg[1289]) );
  DFF \sreg_reg[1288]  ( .D(c[1296]), .CLK(clk), .RST(rst), .Q(sreg[1288]) );
  DFF \sreg_reg[1287]  ( .D(c[1295]), .CLK(clk), .RST(rst), .Q(sreg[1287]) );
  DFF \sreg_reg[1286]  ( .D(c[1294]), .CLK(clk), .RST(rst), .Q(sreg[1286]) );
  DFF \sreg_reg[1285]  ( .D(c[1293]), .CLK(clk), .RST(rst), .Q(sreg[1285]) );
  DFF \sreg_reg[1284]  ( .D(c[1292]), .CLK(clk), .RST(rst), .Q(sreg[1284]) );
  DFF \sreg_reg[1283]  ( .D(c[1291]), .CLK(clk), .RST(rst), .Q(sreg[1283]) );
  DFF \sreg_reg[1282]  ( .D(c[1290]), .CLK(clk), .RST(rst), .Q(sreg[1282]) );
  DFF \sreg_reg[1281]  ( .D(c[1289]), .CLK(clk), .RST(rst), .Q(sreg[1281]) );
  DFF \sreg_reg[1280]  ( .D(c[1288]), .CLK(clk), .RST(rst), .Q(sreg[1280]) );
  DFF \sreg_reg[1279]  ( .D(c[1287]), .CLK(clk), .RST(rst), .Q(sreg[1279]) );
  DFF \sreg_reg[1278]  ( .D(c[1286]), .CLK(clk), .RST(rst), .Q(sreg[1278]) );
  DFF \sreg_reg[1277]  ( .D(c[1285]), .CLK(clk), .RST(rst), .Q(sreg[1277]) );
  DFF \sreg_reg[1276]  ( .D(c[1284]), .CLK(clk), .RST(rst), .Q(sreg[1276]) );
  DFF \sreg_reg[1275]  ( .D(c[1283]), .CLK(clk), .RST(rst), .Q(sreg[1275]) );
  DFF \sreg_reg[1274]  ( .D(c[1282]), .CLK(clk), .RST(rst), .Q(sreg[1274]) );
  DFF \sreg_reg[1273]  ( .D(c[1281]), .CLK(clk), .RST(rst), .Q(sreg[1273]) );
  DFF \sreg_reg[1272]  ( .D(c[1280]), .CLK(clk), .RST(rst), .Q(sreg[1272]) );
  DFF \sreg_reg[1271]  ( .D(c[1279]), .CLK(clk), .RST(rst), .Q(sreg[1271]) );
  DFF \sreg_reg[1270]  ( .D(c[1278]), .CLK(clk), .RST(rst), .Q(sreg[1270]) );
  DFF \sreg_reg[1269]  ( .D(c[1277]), .CLK(clk), .RST(rst), .Q(sreg[1269]) );
  DFF \sreg_reg[1268]  ( .D(c[1276]), .CLK(clk), .RST(rst), .Q(sreg[1268]) );
  DFF \sreg_reg[1267]  ( .D(c[1275]), .CLK(clk), .RST(rst), .Q(sreg[1267]) );
  DFF \sreg_reg[1266]  ( .D(c[1274]), .CLK(clk), .RST(rst), .Q(sreg[1266]) );
  DFF \sreg_reg[1265]  ( .D(c[1273]), .CLK(clk), .RST(rst), .Q(sreg[1265]) );
  DFF \sreg_reg[1264]  ( .D(c[1272]), .CLK(clk), .RST(rst), .Q(sreg[1264]) );
  DFF \sreg_reg[1263]  ( .D(c[1271]), .CLK(clk), .RST(rst), .Q(sreg[1263]) );
  DFF \sreg_reg[1262]  ( .D(c[1270]), .CLK(clk), .RST(rst), .Q(sreg[1262]) );
  DFF \sreg_reg[1261]  ( .D(c[1269]), .CLK(clk), .RST(rst), .Q(sreg[1261]) );
  DFF \sreg_reg[1260]  ( .D(c[1268]), .CLK(clk), .RST(rst), .Q(sreg[1260]) );
  DFF \sreg_reg[1259]  ( .D(c[1267]), .CLK(clk), .RST(rst), .Q(sreg[1259]) );
  DFF \sreg_reg[1258]  ( .D(c[1266]), .CLK(clk), .RST(rst), .Q(sreg[1258]) );
  DFF \sreg_reg[1257]  ( .D(c[1265]), .CLK(clk), .RST(rst), .Q(sreg[1257]) );
  DFF \sreg_reg[1256]  ( .D(c[1264]), .CLK(clk), .RST(rst), .Q(sreg[1256]) );
  DFF \sreg_reg[1255]  ( .D(c[1263]), .CLK(clk), .RST(rst), .Q(sreg[1255]) );
  DFF \sreg_reg[1254]  ( .D(c[1262]), .CLK(clk), .RST(rst), .Q(sreg[1254]) );
  DFF \sreg_reg[1253]  ( .D(c[1261]), .CLK(clk), .RST(rst), .Q(sreg[1253]) );
  DFF \sreg_reg[1252]  ( .D(c[1260]), .CLK(clk), .RST(rst), .Q(sreg[1252]) );
  DFF \sreg_reg[1251]  ( .D(c[1259]), .CLK(clk), .RST(rst), .Q(sreg[1251]) );
  DFF \sreg_reg[1250]  ( .D(c[1258]), .CLK(clk), .RST(rst), .Q(sreg[1250]) );
  DFF \sreg_reg[1249]  ( .D(c[1257]), .CLK(clk), .RST(rst), .Q(sreg[1249]) );
  DFF \sreg_reg[1248]  ( .D(c[1256]), .CLK(clk), .RST(rst), .Q(sreg[1248]) );
  DFF \sreg_reg[1247]  ( .D(c[1255]), .CLK(clk), .RST(rst), .Q(sreg[1247]) );
  DFF \sreg_reg[1246]  ( .D(c[1254]), .CLK(clk), .RST(rst), .Q(sreg[1246]) );
  DFF \sreg_reg[1245]  ( .D(c[1253]), .CLK(clk), .RST(rst), .Q(sreg[1245]) );
  DFF \sreg_reg[1244]  ( .D(c[1252]), .CLK(clk), .RST(rst), .Q(sreg[1244]) );
  DFF \sreg_reg[1243]  ( .D(c[1251]), .CLK(clk), .RST(rst), .Q(sreg[1243]) );
  DFF \sreg_reg[1242]  ( .D(c[1250]), .CLK(clk), .RST(rst), .Q(sreg[1242]) );
  DFF \sreg_reg[1241]  ( .D(c[1249]), .CLK(clk), .RST(rst), .Q(sreg[1241]) );
  DFF \sreg_reg[1240]  ( .D(c[1248]), .CLK(clk), .RST(rst), .Q(sreg[1240]) );
  DFF \sreg_reg[1239]  ( .D(c[1247]), .CLK(clk), .RST(rst), .Q(sreg[1239]) );
  DFF \sreg_reg[1238]  ( .D(c[1246]), .CLK(clk), .RST(rst), .Q(sreg[1238]) );
  DFF \sreg_reg[1237]  ( .D(c[1245]), .CLK(clk), .RST(rst), .Q(sreg[1237]) );
  DFF \sreg_reg[1236]  ( .D(c[1244]), .CLK(clk), .RST(rst), .Q(sreg[1236]) );
  DFF \sreg_reg[1235]  ( .D(c[1243]), .CLK(clk), .RST(rst), .Q(sreg[1235]) );
  DFF \sreg_reg[1234]  ( .D(c[1242]), .CLK(clk), .RST(rst), .Q(sreg[1234]) );
  DFF \sreg_reg[1233]  ( .D(c[1241]), .CLK(clk), .RST(rst), .Q(sreg[1233]) );
  DFF \sreg_reg[1232]  ( .D(c[1240]), .CLK(clk), .RST(rst), .Q(sreg[1232]) );
  DFF \sreg_reg[1231]  ( .D(c[1239]), .CLK(clk), .RST(rst), .Q(sreg[1231]) );
  DFF \sreg_reg[1230]  ( .D(c[1238]), .CLK(clk), .RST(rst), .Q(sreg[1230]) );
  DFF \sreg_reg[1229]  ( .D(c[1237]), .CLK(clk), .RST(rst), .Q(sreg[1229]) );
  DFF \sreg_reg[1228]  ( .D(c[1236]), .CLK(clk), .RST(rst), .Q(sreg[1228]) );
  DFF \sreg_reg[1227]  ( .D(c[1235]), .CLK(clk), .RST(rst), .Q(sreg[1227]) );
  DFF \sreg_reg[1226]  ( .D(c[1234]), .CLK(clk), .RST(rst), .Q(sreg[1226]) );
  DFF \sreg_reg[1225]  ( .D(c[1233]), .CLK(clk), .RST(rst), .Q(sreg[1225]) );
  DFF \sreg_reg[1224]  ( .D(c[1232]), .CLK(clk), .RST(rst), .Q(sreg[1224]) );
  DFF \sreg_reg[1223]  ( .D(c[1231]), .CLK(clk), .RST(rst), .Q(sreg[1223]) );
  DFF \sreg_reg[1222]  ( .D(c[1230]), .CLK(clk), .RST(rst), .Q(sreg[1222]) );
  DFF \sreg_reg[1221]  ( .D(c[1229]), .CLK(clk), .RST(rst), .Q(sreg[1221]) );
  DFF \sreg_reg[1220]  ( .D(c[1228]), .CLK(clk), .RST(rst), .Q(sreg[1220]) );
  DFF \sreg_reg[1219]  ( .D(c[1227]), .CLK(clk), .RST(rst), .Q(sreg[1219]) );
  DFF \sreg_reg[1218]  ( .D(c[1226]), .CLK(clk), .RST(rst), .Q(sreg[1218]) );
  DFF \sreg_reg[1217]  ( .D(c[1225]), .CLK(clk), .RST(rst), .Q(sreg[1217]) );
  DFF \sreg_reg[1216]  ( .D(c[1224]), .CLK(clk), .RST(rst), .Q(sreg[1216]) );
  DFF \sreg_reg[1215]  ( .D(c[1223]), .CLK(clk), .RST(rst), .Q(sreg[1215]) );
  DFF \sreg_reg[1214]  ( .D(c[1222]), .CLK(clk), .RST(rst), .Q(sreg[1214]) );
  DFF \sreg_reg[1213]  ( .D(c[1221]), .CLK(clk), .RST(rst), .Q(sreg[1213]) );
  DFF \sreg_reg[1212]  ( .D(c[1220]), .CLK(clk), .RST(rst), .Q(sreg[1212]) );
  DFF \sreg_reg[1211]  ( .D(c[1219]), .CLK(clk), .RST(rst), .Q(sreg[1211]) );
  DFF \sreg_reg[1210]  ( .D(c[1218]), .CLK(clk), .RST(rst), .Q(sreg[1210]) );
  DFF \sreg_reg[1209]  ( .D(c[1217]), .CLK(clk), .RST(rst), .Q(sreg[1209]) );
  DFF \sreg_reg[1208]  ( .D(c[1216]), .CLK(clk), .RST(rst), .Q(sreg[1208]) );
  DFF \sreg_reg[1207]  ( .D(c[1215]), .CLK(clk), .RST(rst), .Q(sreg[1207]) );
  DFF \sreg_reg[1206]  ( .D(c[1214]), .CLK(clk), .RST(rst), .Q(sreg[1206]) );
  DFF \sreg_reg[1205]  ( .D(c[1213]), .CLK(clk), .RST(rst), .Q(sreg[1205]) );
  DFF \sreg_reg[1204]  ( .D(c[1212]), .CLK(clk), .RST(rst), .Q(sreg[1204]) );
  DFF \sreg_reg[1203]  ( .D(c[1211]), .CLK(clk), .RST(rst), .Q(sreg[1203]) );
  DFF \sreg_reg[1202]  ( .D(c[1210]), .CLK(clk), .RST(rst), .Q(sreg[1202]) );
  DFF \sreg_reg[1201]  ( .D(c[1209]), .CLK(clk), .RST(rst), .Q(sreg[1201]) );
  DFF \sreg_reg[1200]  ( .D(c[1208]), .CLK(clk), .RST(rst), .Q(sreg[1200]) );
  DFF \sreg_reg[1199]  ( .D(c[1207]), .CLK(clk), .RST(rst), .Q(sreg[1199]) );
  DFF \sreg_reg[1198]  ( .D(c[1206]), .CLK(clk), .RST(rst), .Q(sreg[1198]) );
  DFF \sreg_reg[1197]  ( .D(c[1205]), .CLK(clk), .RST(rst), .Q(sreg[1197]) );
  DFF \sreg_reg[1196]  ( .D(c[1204]), .CLK(clk), .RST(rst), .Q(sreg[1196]) );
  DFF \sreg_reg[1195]  ( .D(c[1203]), .CLK(clk), .RST(rst), .Q(sreg[1195]) );
  DFF \sreg_reg[1194]  ( .D(c[1202]), .CLK(clk), .RST(rst), .Q(sreg[1194]) );
  DFF \sreg_reg[1193]  ( .D(c[1201]), .CLK(clk), .RST(rst), .Q(sreg[1193]) );
  DFF \sreg_reg[1192]  ( .D(c[1200]), .CLK(clk), .RST(rst), .Q(sreg[1192]) );
  DFF \sreg_reg[1191]  ( .D(c[1199]), .CLK(clk), .RST(rst), .Q(sreg[1191]) );
  DFF \sreg_reg[1190]  ( .D(c[1198]), .CLK(clk), .RST(rst), .Q(sreg[1190]) );
  DFF \sreg_reg[1189]  ( .D(c[1197]), .CLK(clk), .RST(rst), .Q(sreg[1189]) );
  DFF \sreg_reg[1188]  ( .D(c[1196]), .CLK(clk), .RST(rst), .Q(sreg[1188]) );
  DFF \sreg_reg[1187]  ( .D(c[1195]), .CLK(clk), .RST(rst), .Q(sreg[1187]) );
  DFF \sreg_reg[1186]  ( .D(c[1194]), .CLK(clk), .RST(rst), .Q(sreg[1186]) );
  DFF \sreg_reg[1185]  ( .D(c[1193]), .CLK(clk), .RST(rst), .Q(sreg[1185]) );
  DFF \sreg_reg[1184]  ( .D(c[1192]), .CLK(clk), .RST(rst), .Q(sreg[1184]) );
  DFF \sreg_reg[1183]  ( .D(c[1191]), .CLK(clk), .RST(rst), .Q(sreg[1183]) );
  DFF \sreg_reg[1182]  ( .D(c[1190]), .CLK(clk), .RST(rst), .Q(sreg[1182]) );
  DFF \sreg_reg[1181]  ( .D(c[1189]), .CLK(clk), .RST(rst), .Q(sreg[1181]) );
  DFF \sreg_reg[1180]  ( .D(c[1188]), .CLK(clk), .RST(rst), .Q(sreg[1180]) );
  DFF \sreg_reg[1179]  ( .D(c[1187]), .CLK(clk), .RST(rst), .Q(sreg[1179]) );
  DFF \sreg_reg[1178]  ( .D(c[1186]), .CLK(clk), .RST(rst), .Q(sreg[1178]) );
  DFF \sreg_reg[1177]  ( .D(c[1185]), .CLK(clk), .RST(rst), .Q(sreg[1177]) );
  DFF \sreg_reg[1176]  ( .D(c[1184]), .CLK(clk), .RST(rst), .Q(sreg[1176]) );
  DFF \sreg_reg[1175]  ( .D(c[1183]), .CLK(clk), .RST(rst), .Q(sreg[1175]) );
  DFF \sreg_reg[1174]  ( .D(c[1182]), .CLK(clk), .RST(rst), .Q(sreg[1174]) );
  DFF \sreg_reg[1173]  ( .D(c[1181]), .CLK(clk), .RST(rst), .Q(sreg[1173]) );
  DFF \sreg_reg[1172]  ( .D(c[1180]), .CLK(clk), .RST(rst), .Q(sreg[1172]) );
  DFF \sreg_reg[1171]  ( .D(c[1179]), .CLK(clk), .RST(rst), .Q(sreg[1171]) );
  DFF \sreg_reg[1170]  ( .D(c[1178]), .CLK(clk), .RST(rst), .Q(sreg[1170]) );
  DFF \sreg_reg[1169]  ( .D(c[1177]), .CLK(clk), .RST(rst), .Q(sreg[1169]) );
  DFF \sreg_reg[1168]  ( .D(c[1176]), .CLK(clk), .RST(rst), .Q(sreg[1168]) );
  DFF \sreg_reg[1167]  ( .D(c[1175]), .CLK(clk), .RST(rst), .Q(sreg[1167]) );
  DFF \sreg_reg[1166]  ( .D(c[1174]), .CLK(clk), .RST(rst), .Q(sreg[1166]) );
  DFF \sreg_reg[1165]  ( .D(c[1173]), .CLK(clk), .RST(rst), .Q(sreg[1165]) );
  DFF \sreg_reg[1164]  ( .D(c[1172]), .CLK(clk), .RST(rst), .Q(sreg[1164]) );
  DFF \sreg_reg[1163]  ( .D(c[1171]), .CLK(clk), .RST(rst), .Q(sreg[1163]) );
  DFF \sreg_reg[1162]  ( .D(c[1170]), .CLK(clk), .RST(rst), .Q(sreg[1162]) );
  DFF \sreg_reg[1161]  ( .D(c[1169]), .CLK(clk), .RST(rst), .Q(sreg[1161]) );
  DFF \sreg_reg[1160]  ( .D(c[1168]), .CLK(clk), .RST(rst), .Q(sreg[1160]) );
  DFF \sreg_reg[1159]  ( .D(c[1167]), .CLK(clk), .RST(rst), .Q(sreg[1159]) );
  DFF \sreg_reg[1158]  ( .D(c[1166]), .CLK(clk), .RST(rst), .Q(sreg[1158]) );
  DFF \sreg_reg[1157]  ( .D(c[1165]), .CLK(clk), .RST(rst), .Q(sreg[1157]) );
  DFF \sreg_reg[1156]  ( .D(c[1164]), .CLK(clk), .RST(rst), .Q(sreg[1156]) );
  DFF \sreg_reg[1155]  ( .D(c[1163]), .CLK(clk), .RST(rst), .Q(sreg[1155]) );
  DFF \sreg_reg[1154]  ( .D(c[1162]), .CLK(clk), .RST(rst), .Q(sreg[1154]) );
  DFF \sreg_reg[1153]  ( .D(c[1161]), .CLK(clk), .RST(rst), .Q(sreg[1153]) );
  DFF \sreg_reg[1152]  ( .D(c[1160]), .CLK(clk), .RST(rst), .Q(sreg[1152]) );
  DFF \sreg_reg[1151]  ( .D(c[1159]), .CLK(clk), .RST(rst), .Q(sreg[1151]) );
  DFF \sreg_reg[1150]  ( .D(c[1158]), .CLK(clk), .RST(rst), .Q(sreg[1150]) );
  DFF \sreg_reg[1149]  ( .D(c[1157]), .CLK(clk), .RST(rst), .Q(sreg[1149]) );
  DFF \sreg_reg[1148]  ( .D(c[1156]), .CLK(clk), .RST(rst), .Q(sreg[1148]) );
  DFF \sreg_reg[1147]  ( .D(c[1155]), .CLK(clk), .RST(rst), .Q(sreg[1147]) );
  DFF \sreg_reg[1146]  ( .D(c[1154]), .CLK(clk), .RST(rst), .Q(sreg[1146]) );
  DFF \sreg_reg[1145]  ( .D(c[1153]), .CLK(clk), .RST(rst), .Q(sreg[1145]) );
  DFF \sreg_reg[1144]  ( .D(c[1152]), .CLK(clk), .RST(rst), .Q(sreg[1144]) );
  DFF \sreg_reg[1143]  ( .D(c[1151]), .CLK(clk), .RST(rst), .Q(sreg[1143]) );
  DFF \sreg_reg[1142]  ( .D(c[1150]), .CLK(clk), .RST(rst), .Q(sreg[1142]) );
  DFF \sreg_reg[1141]  ( .D(c[1149]), .CLK(clk), .RST(rst), .Q(sreg[1141]) );
  DFF \sreg_reg[1140]  ( .D(c[1148]), .CLK(clk), .RST(rst), .Q(sreg[1140]) );
  DFF \sreg_reg[1139]  ( .D(c[1147]), .CLK(clk), .RST(rst), .Q(sreg[1139]) );
  DFF \sreg_reg[1138]  ( .D(c[1146]), .CLK(clk), .RST(rst), .Q(sreg[1138]) );
  DFF \sreg_reg[1137]  ( .D(c[1145]), .CLK(clk), .RST(rst), .Q(sreg[1137]) );
  DFF \sreg_reg[1136]  ( .D(c[1144]), .CLK(clk), .RST(rst), .Q(sreg[1136]) );
  DFF \sreg_reg[1135]  ( .D(c[1143]), .CLK(clk), .RST(rst), .Q(sreg[1135]) );
  DFF \sreg_reg[1134]  ( .D(c[1142]), .CLK(clk), .RST(rst), .Q(sreg[1134]) );
  DFF \sreg_reg[1133]  ( .D(c[1141]), .CLK(clk), .RST(rst), .Q(sreg[1133]) );
  DFF \sreg_reg[1132]  ( .D(c[1140]), .CLK(clk), .RST(rst), .Q(sreg[1132]) );
  DFF \sreg_reg[1131]  ( .D(c[1139]), .CLK(clk), .RST(rst), .Q(sreg[1131]) );
  DFF \sreg_reg[1130]  ( .D(c[1138]), .CLK(clk), .RST(rst), .Q(sreg[1130]) );
  DFF \sreg_reg[1129]  ( .D(c[1137]), .CLK(clk), .RST(rst), .Q(sreg[1129]) );
  DFF \sreg_reg[1128]  ( .D(c[1136]), .CLK(clk), .RST(rst), .Q(sreg[1128]) );
  DFF \sreg_reg[1127]  ( .D(c[1135]), .CLK(clk), .RST(rst), .Q(sreg[1127]) );
  DFF \sreg_reg[1126]  ( .D(c[1134]), .CLK(clk), .RST(rst), .Q(sreg[1126]) );
  DFF \sreg_reg[1125]  ( .D(c[1133]), .CLK(clk), .RST(rst), .Q(sreg[1125]) );
  DFF \sreg_reg[1124]  ( .D(c[1132]), .CLK(clk), .RST(rst), .Q(sreg[1124]) );
  DFF \sreg_reg[1123]  ( .D(c[1131]), .CLK(clk), .RST(rst), .Q(sreg[1123]) );
  DFF \sreg_reg[1122]  ( .D(c[1130]), .CLK(clk), .RST(rst), .Q(sreg[1122]) );
  DFF \sreg_reg[1121]  ( .D(c[1129]), .CLK(clk), .RST(rst), .Q(sreg[1121]) );
  DFF \sreg_reg[1120]  ( .D(c[1128]), .CLK(clk), .RST(rst), .Q(sreg[1120]) );
  DFF \sreg_reg[1119]  ( .D(c[1127]), .CLK(clk), .RST(rst), .Q(sreg[1119]) );
  DFF \sreg_reg[1118]  ( .D(c[1126]), .CLK(clk), .RST(rst), .Q(sreg[1118]) );
  DFF \sreg_reg[1117]  ( .D(c[1125]), .CLK(clk), .RST(rst), .Q(sreg[1117]) );
  DFF \sreg_reg[1116]  ( .D(c[1124]), .CLK(clk), .RST(rst), .Q(sreg[1116]) );
  DFF \sreg_reg[1115]  ( .D(c[1123]), .CLK(clk), .RST(rst), .Q(sreg[1115]) );
  DFF \sreg_reg[1114]  ( .D(c[1122]), .CLK(clk), .RST(rst), .Q(sreg[1114]) );
  DFF \sreg_reg[1113]  ( .D(c[1121]), .CLK(clk), .RST(rst), .Q(sreg[1113]) );
  DFF \sreg_reg[1112]  ( .D(c[1120]), .CLK(clk), .RST(rst), .Q(sreg[1112]) );
  DFF \sreg_reg[1111]  ( .D(c[1119]), .CLK(clk), .RST(rst), .Q(sreg[1111]) );
  DFF \sreg_reg[1110]  ( .D(c[1118]), .CLK(clk), .RST(rst), .Q(sreg[1110]) );
  DFF \sreg_reg[1109]  ( .D(c[1117]), .CLK(clk), .RST(rst), .Q(sreg[1109]) );
  DFF \sreg_reg[1108]  ( .D(c[1116]), .CLK(clk), .RST(rst), .Q(sreg[1108]) );
  DFF \sreg_reg[1107]  ( .D(c[1115]), .CLK(clk), .RST(rst), .Q(sreg[1107]) );
  DFF \sreg_reg[1106]  ( .D(c[1114]), .CLK(clk), .RST(rst), .Q(sreg[1106]) );
  DFF \sreg_reg[1105]  ( .D(c[1113]), .CLK(clk), .RST(rst), .Q(sreg[1105]) );
  DFF \sreg_reg[1104]  ( .D(c[1112]), .CLK(clk), .RST(rst), .Q(sreg[1104]) );
  DFF \sreg_reg[1103]  ( .D(c[1111]), .CLK(clk), .RST(rst), .Q(sreg[1103]) );
  DFF \sreg_reg[1102]  ( .D(c[1110]), .CLK(clk), .RST(rst), .Q(sreg[1102]) );
  DFF \sreg_reg[1101]  ( .D(c[1109]), .CLK(clk), .RST(rst), .Q(sreg[1101]) );
  DFF \sreg_reg[1100]  ( .D(c[1108]), .CLK(clk), .RST(rst), .Q(sreg[1100]) );
  DFF \sreg_reg[1099]  ( .D(c[1107]), .CLK(clk), .RST(rst), .Q(sreg[1099]) );
  DFF \sreg_reg[1098]  ( .D(c[1106]), .CLK(clk), .RST(rst), .Q(sreg[1098]) );
  DFF \sreg_reg[1097]  ( .D(c[1105]), .CLK(clk), .RST(rst), .Q(sreg[1097]) );
  DFF \sreg_reg[1096]  ( .D(c[1104]), .CLK(clk), .RST(rst), .Q(sreg[1096]) );
  DFF \sreg_reg[1095]  ( .D(c[1103]), .CLK(clk), .RST(rst), .Q(sreg[1095]) );
  DFF \sreg_reg[1094]  ( .D(c[1102]), .CLK(clk), .RST(rst), .Q(sreg[1094]) );
  DFF \sreg_reg[1093]  ( .D(c[1101]), .CLK(clk), .RST(rst), .Q(sreg[1093]) );
  DFF \sreg_reg[1092]  ( .D(c[1100]), .CLK(clk), .RST(rst), .Q(sreg[1092]) );
  DFF \sreg_reg[1091]  ( .D(c[1099]), .CLK(clk), .RST(rst), .Q(sreg[1091]) );
  DFF \sreg_reg[1090]  ( .D(c[1098]), .CLK(clk), .RST(rst), .Q(sreg[1090]) );
  DFF \sreg_reg[1089]  ( .D(c[1097]), .CLK(clk), .RST(rst), .Q(sreg[1089]) );
  DFF \sreg_reg[1088]  ( .D(c[1096]), .CLK(clk), .RST(rst), .Q(sreg[1088]) );
  DFF \sreg_reg[1087]  ( .D(c[1095]), .CLK(clk), .RST(rst), .Q(sreg[1087]) );
  DFF \sreg_reg[1086]  ( .D(c[1094]), .CLK(clk), .RST(rst), .Q(sreg[1086]) );
  DFF \sreg_reg[1085]  ( .D(c[1093]), .CLK(clk), .RST(rst), .Q(sreg[1085]) );
  DFF \sreg_reg[1084]  ( .D(c[1092]), .CLK(clk), .RST(rst), .Q(sreg[1084]) );
  DFF \sreg_reg[1083]  ( .D(c[1091]), .CLK(clk), .RST(rst), .Q(sreg[1083]) );
  DFF \sreg_reg[1082]  ( .D(c[1090]), .CLK(clk), .RST(rst), .Q(sreg[1082]) );
  DFF \sreg_reg[1081]  ( .D(c[1089]), .CLK(clk), .RST(rst), .Q(sreg[1081]) );
  DFF \sreg_reg[1080]  ( .D(c[1088]), .CLK(clk), .RST(rst), .Q(sreg[1080]) );
  DFF \sreg_reg[1079]  ( .D(c[1087]), .CLK(clk), .RST(rst), .Q(sreg[1079]) );
  DFF \sreg_reg[1078]  ( .D(c[1086]), .CLK(clk), .RST(rst), .Q(sreg[1078]) );
  DFF \sreg_reg[1077]  ( .D(c[1085]), .CLK(clk), .RST(rst), .Q(sreg[1077]) );
  DFF \sreg_reg[1076]  ( .D(c[1084]), .CLK(clk), .RST(rst), .Q(sreg[1076]) );
  DFF \sreg_reg[1075]  ( .D(c[1083]), .CLK(clk), .RST(rst), .Q(sreg[1075]) );
  DFF \sreg_reg[1074]  ( .D(c[1082]), .CLK(clk), .RST(rst), .Q(sreg[1074]) );
  DFF \sreg_reg[1073]  ( .D(c[1081]), .CLK(clk), .RST(rst), .Q(sreg[1073]) );
  DFF \sreg_reg[1072]  ( .D(c[1080]), .CLK(clk), .RST(rst), .Q(sreg[1072]) );
  DFF \sreg_reg[1071]  ( .D(c[1079]), .CLK(clk), .RST(rst), .Q(sreg[1071]) );
  DFF \sreg_reg[1070]  ( .D(c[1078]), .CLK(clk), .RST(rst), .Q(sreg[1070]) );
  DFF \sreg_reg[1069]  ( .D(c[1077]), .CLK(clk), .RST(rst), .Q(sreg[1069]) );
  DFF \sreg_reg[1068]  ( .D(c[1076]), .CLK(clk), .RST(rst), .Q(sreg[1068]) );
  DFF \sreg_reg[1067]  ( .D(c[1075]), .CLK(clk), .RST(rst), .Q(sreg[1067]) );
  DFF \sreg_reg[1066]  ( .D(c[1074]), .CLK(clk), .RST(rst), .Q(sreg[1066]) );
  DFF \sreg_reg[1065]  ( .D(c[1073]), .CLK(clk), .RST(rst), .Q(sreg[1065]) );
  DFF \sreg_reg[1064]  ( .D(c[1072]), .CLK(clk), .RST(rst), .Q(sreg[1064]) );
  DFF \sreg_reg[1063]  ( .D(c[1071]), .CLK(clk), .RST(rst), .Q(sreg[1063]) );
  DFF \sreg_reg[1062]  ( .D(c[1070]), .CLK(clk), .RST(rst), .Q(sreg[1062]) );
  DFF \sreg_reg[1061]  ( .D(c[1069]), .CLK(clk), .RST(rst), .Q(sreg[1061]) );
  DFF \sreg_reg[1060]  ( .D(c[1068]), .CLK(clk), .RST(rst), .Q(sreg[1060]) );
  DFF \sreg_reg[1059]  ( .D(c[1067]), .CLK(clk), .RST(rst), .Q(sreg[1059]) );
  DFF \sreg_reg[1058]  ( .D(c[1066]), .CLK(clk), .RST(rst), .Q(sreg[1058]) );
  DFF \sreg_reg[1057]  ( .D(c[1065]), .CLK(clk), .RST(rst), .Q(sreg[1057]) );
  DFF \sreg_reg[1056]  ( .D(c[1064]), .CLK(clk), .RST(rst), .Q(sreg[1056]) );
  DFF \sreg_reg[1055]  ( .D(c[1063]), .CLK(clk), .RST(rst), .Q(sreg[1055]) );
  DFF \sreg_reg[1054]  ( .D(c[1062]), .CLK(clk), .RST(rst), .Q(sreg[1054]) );
  DFF \sreg_reg[1053]  ( .D(c[1061]), .CLK(clk), .RST(rst), .Q(sreg[1053]) );
  DFF \sreg_reg[1052]  ( .D(c[1060]), .CLK(clk), .RST(rst), .Q(sreg[1052]) );
  DFF \sreg_reg[1051]  ( .D(c[1059]), .CLK(clk), .RST(rst), .Q(sreg[1051]) );
  DFF \sreg_reg[1050]  ( .D(c[1058]), .CLK(clk), .RST(rst), .Q(sreg[1050]) );
  DFF \sreg_reg[1049]  ( .D(c[1057]), .CLK(clk), .RST(rst), .Q(sreg[1049]) );
  DFF \sreg_reg[1048]  ( .D(c[1056]), .CLK(clk), .RST(rst), .Q(sreg[1048]) );
  DFF \sreg_reg[1047]  ( .D(c[1055]), .CLK(clk), .RST(rst), .Q(sreg[1047]) );
  DFF \sreg_reg[1046]  ( .D(c[1054]), .CLK(clk), .RST(rst), .Q(sreg[1046]) );
  DFF \sreg_reg[1045]  ( .D(c[1053]), .CLK(clk), .RST(rst), .Q(sreg[1045]) );
  DFF \sreg_reg[1044]  ( .D(c[1052]), .CLK(clk), .RST(rst), .Q(sreg[1044]) );
  DFF \sreg_reg[1043]  ( .D(c[1051]), .CLK(clk), .RST(rst), .Q(sreg[1043]) );
  DFF \sreg_reg[1042]  ( .D(c[1050]), .CLK(clk), .RST(rst), .Q(sreg[1042]) );
  DFF \sreg_reg[1041]  ( .D(c[1049]), .CLK(clk), .RST(rst), .Q(sreg[1041]) );
  DFF \sreg_reg[1040]  ( .D(c[1048]), .CLK(clk), .RST(rst), .Q(sreg[1040]) );
  DFF \sreg_reg[1039]  ( .D(c[1047]), .CLK(clk), .RST(rst), .Q(sreg[1039]) );
  DFF \sreg_reg[1038]  ( .D(c[1046]), .CLK(clk), .RST(rst), .Q(sreg[1038]) );
  DFF \sreg_reg[1037]  ( .D(c[1045]), .CLK(clk), .RST(rst), .Q(sreg[1037]) );
  DFF \sreg_reg[1036]  ( .D(c[1044]), .CLK(clk), .RST(rst), .Q(sreg[1036]) );
  DFF \sreg_reg[1035]  ( .D(c[1043]), .CLK(clk), .RST(rst), .Q(sreg[1035]) );
  DFF \sreg_reg[1034]  ( .D(c[1042]), .CLK(clk), .RST(rst), .Q(sreg[1034]) );
  DFF \sreg_reg[1033]  ( .D(c[1041]), .CLK(clk), .RST(rst), .Q(sreg[1033]) );
  DFF \sreg_reg[1032]  ( .D(c[1040]), .CLK(clk), .RST(rst), .Q(sreg[1032]) );
  DFF \sreg_reg[1031]  ( .D(c[1039]), .CLK(clk), .RST(rst), .Q(sreg[1031]) );
  DFF \sreg_reg[1030]  ( .D(c[1038]), .CLK(clk), .RST(rst), .Q(sreg[1030]) );
  DFF \sreg_reg[1029]  ( .D(c[1037]), .CLK(clk), .RST(rst), .Q(sreg[1029]) );
  DFF \sreg_reg[1028]  ( .D(c[1036]), .CLK(clk), .RST(rst), .Q(sreg[1028]) );
  DFF \sreg_reg[1027]  ( .D(c[1035]), .CLK(clk), .RST(rst), .Q(sreg[1027]) );
  DFF \sreg_reg[1026]  ( .D(c[1034]), .CLK(clk), .RST(rst), .Q(sreg[1026]) );
  DFF \sreg_reg[1025]  ( .D(c[1033]), .CLK(clk), .RST(rst), .Q(sreg[1025]) );
  DFF \sreg_reg[1024]  ( .D(c[1032]), .CLK(clk), .RST(rst), .Q(sreg[1024]) );
  DFF \sreg_reg[1023]  ( .D(c[1031]), .CLK(clk), .RST(rst), .Q(sreg[1023]) );
  DFF \sreg_reg[1022]  ( .D(c[1030]), .CLK(clk), .RST(rst), .Q(sreg[1022]) );
  DFF \sreg_reg[1021]  ( .D(c[1029]), .CLK(clk), .RST(rst), .Q(sreg[1021]) );
  DFF \sreg_reg[1020]  ( .D(c[1028]), .CLK(clk), .RST(rst), .Q(sreg[1020]) );
  DFF \sreg_reg[1019]  ( .D(c[1027]), .CLK(clk), .RST(rst), .Q(sreg[1019]) );
  DFF \sreg_reg[1018]  ( .D(c[1026]), .CLK(clk), .RST(rst), .Q(sreg[1018]) );
  DFF \sreg_reg[1017]  ( .D(c[1025]), .CLK(clk), .RST(rst), .Q(sreg[1017]) );
  DFF \sreg_reg[1016]  ( .D(c[1024]), .CLK(clk), .RST(rst), .Q(sreg[1016]) );
  DFF \sreg_reg[1015]  ( .D(c[1023]), .CLK(clk), .RST(rst), .Q(c[1015]) );
  DFF \sreg_reg[1014]  ( .D(c[1022]), .CLK(clk), .RST(rst), .Q(c[1014]) );
  DFF \sreg_reg[1013]  ( .D(c[1021]), .CLK(clk), .RST(rst), .Q(c[1013]) );
  DFF \sreg_reg[1012]  ( .D(c[1020]), .CLK(clk), .RST(rst), .Q(c[1012]) );
  DFF \sreg_reg[1011]  ( .D(c[1019]), .CLK(clk), .RST(rst), .Q(c[1011]) );
  DFF \sreg_reg[1010]  ( .D(c[1018]), .CLK(clk), .RST(rst), .Q(c[1010]) );
  DFF \sreg_reg[1009]  ( .D(c[1017]), .CLK(clk), .RST(rst), .Q(c[1009]) );
  DFF \sreg_reg[1008]  ( .D(c[1016]), .CLK(clk), .RST(rst), .Q(c[1008]) );
  DFF \sreg_reg[1007]  ( .D(c[1015]), .CLK(clk), .RST(rst), .Q(c[1007]) );
  DFF \sreg_reg[1006]  ( .D(c[1014]), .CLK(clk), .RST(rst), .Q(c[1006]) );
  DFF \sreg_reg[1005]  ( .D(c[1013]), .CLK(clk), .RST(rst), .Q(c[1005]) );
  DFF \sreg_reg[1004]  ( .D(c[1012]), .CLK(clk), .RST(rst), .Q(c[1004]) );
  DFF \sreg_reg[1003]  ( .D(c[1011]), .CLK(clk), .RST(rst), .Q(c[1003]) );
  DFF \sreg_reg[1002]  ( .D(c[1010]), .CLK(clk), .RST(rst), .Q(c[1002]) );
  DFF \sreg_reg[1001]  ( .D(c[1009]), .CLK(clk), .RST(rst), .Q(c[1001]) );
  DFF \sreg_reg[1000]  ( .D(c[1008]), .CLK(clk), .RST(rst), .Q(c[1000]) );
  DFF \sreg_reg[999]  ( .D(c[1007]), .CLK(clk), .RST(rst), .Q(c[999]) );
  DFF \sreg_reg[998]  ( .D(c[1006]), .CLK(clk), .RST(rst), .Q(c[998]) );
  DFF \sreg_reg[997]  ( .D(c[1005]), .CLK(clk), .RST(rst), .Q(c[997]) );
  DFF \sreg_reg[996]  ( .D(c[1004]), .CLK(clk), .RST(rst), .Q(c[996]) );
  DFF \sreg_reg[995]  ( .D(c[1003]), .CLK(clk), .RST(rst), .Q(c[995]) );
  DFF \sreg_reg[994]  ( .D(c[1002]), .CLK(clk), .RST(rst), .Q(c[994]) );
  DFF \sreg_reg[993]  ( .D(c[1001]), .CLK(clk), .RST(rst), .Q(c[993]) );
  DFF \sreg_reg[992]  ( .D(c[1000]), .CLK(clk), .RST(rst), .Q(c[992]) );
  DFF \sreg_reg[991]  ( .D(c[999]), .CLK(clk), .RST(rst), .Q(c[991]) );
  DFF \sreg_reg[990]  ( .D(c[998]), .CLK(clk), .RST(rst), .Q(c[990]) );
  DFF \sreg_reg[989]  ( .D(c[997]), .CLK(clk), .RST(rst), .Q(c[989]) );
  DFF \sreg_reg[988]  ( .D(c[996]), .CLK(clk), .RST(rst), .Q(c[988]) );
  DFF \sreg_reg[987]  ( .D(c[995]), .CLK(clk), .RST(rst), .Q(c[987]) );
  DFF \sreg_reg[986]  ( .D(c[994]), .CLK(clk), .RST(rst), .Q(c[986]) );
  DFF \sreg_reg[985]  ( .D(c[993]), .CLK(clk), .RST(rst), .Q(c[985]) );
  DFF \sreg_reg[984]  ( .D(c[992]), .CLK(clk), .RST(rst), .Q(c[984]) );
  DFF \sreg_reg[983]  ( .D(c[991]), .CLK(clk), .RST(rst), .Q(c[983]) );
  DFF \sreg_reg[982]  ( .D(c[990]), .CLK(clk), .RST(rst), .Q(c[982]) );
  DFF \sreg_reg[981]  ( .D(c[989]), .CLK(clk), .RST(rst), .Q(c[981]) );
  DFF \sreg_reg[980]  ( .D(c[988]), .CLK(clk), .RST(rst), .Q(c[980]) );
  DFF \sreg_reg[979]  ( .D(c[987]), .CLK(clk), .RST(rst), .Q(c[979]) );
  DFF \sreg_reg[978]  ( .D(c[986]), .CLK(clk), .RST(rst), .Q(c[978]) );
  DFF \sreg_reg[977]  ( .D(c[985]), .CLK(clk), .RST(rst), .Q(c[977]) );
  DFF \sreg_reg[976]  ( .D(c[984]), .CLK(clk), .RST(rst), .Q(c[976]) );
  DFF \sreg_reg[975]  ( .D(c[983]), .CLK(clk), .RST(rst), .Q(c[975]) );
  DFF \sreg_reg[974]  ( .D(c[982]), .CLK(clk), .RST(rst), .Q(c[974]) );
  DFF \sreg_reg[973]  ( .D(c[981]), .CLK(clk), .RST(rst), .Q(c[973]) );
  DFF \sreg_reg[972]  ( .D(c[980]), .CLK(clk), .RST(rst), .Q(c[972]) );
  DFF \sreg_reg[971]  ( .D(c[979]), .CLK(clk), .RST(rst), .Q(c[971]) );
  DFF \sreg_reg[970]  ( .D(c[978]), .CLK(clk), .RST(rst), .Q(c[970]) );
  DFF \sreg_reg[969]  ( .D(c[977]), .CLK(clk), .RST(rst), .Q(c[969]) );
  DFF \sreg_reg[968]  ( .D(c[976]), .CLK(clk), .RST(rst), .Q(c[968]) );
  DFF \sreg_reg[967]  ( .D(c[975]), .CLK(clk), .RST(rst), .Q(c[967]) );
  DFF \sreg_reg[966]  ( .D(c[974]), .CLK(clk), .RST(rst), .Q(c[966]) );
  DFF \sreg_reg[965]  ( .D(c[973]), .CLK(clk), .RST(rst), .Q(c[965]) );
  DFF \sreg_reg[964]  ( .D(c[972]), .CLK(clk), .RST(rst), .Q(c[964]) );
  DFF \sreg_reg[963]  ( .D(c[971]), .CLK(clk), .RST(rst), .Q(c[963]) );
  DFF \sreg_reg[962]  ( .D(c[970]), .CLK(clk), .RST(rst), .Q(c[962]) );
  DFF \sreg_reg[961]  ( .D(c[969]), .CLK(clk), .RST(rst), .Q(c[961]) );
  DFF \sreg_reg[960]  ( .D(c[968]), .CLK(clk), .RST(rst), .Q(c[960]) );
  DFF \sreg_reg[959]  ( .D(c[967]), .CLK(clk), .RST(rst), .Q(c[959]) );
  DFF \sreg_reg[958]  ( .D(c[966]), .CLK(clk), .RST(rst), .Q(c[958]) );
  DFF \sreg_reg[957]  ( .D(c[965]), .CLK(clk), .RST(rst), .Q(c[957]) );
  DFF \sreg_reg[956]  ( .D(c[964]), .CLK(clk), .RST(rst), .Q(c[956]) );
  DFF \sreg_reg[955]  ( .D(c[963]), .CLK(clk), .RST(rst), .Q(c[955]) );
  DFF \sreg_reg[954]  ( .D(c[962]), .CLK(clk), .RST(rst), .Q(c[954]) );
  DFF \sreg_reg[953]  ( .D(c[961]), .CLK(clk), .RST(rst), .Q(c[953]) );
  DFF \sreg_reg[952]  ( .D(c[960]), .CLK(clk), .RST(rst), .Q(c[952]) );
  DFF \sreg_reg[951]  ( .D(c[959]), .CLK(clk), .RST(rst), .Q(c[951]) );
  DFF \sreg_reg[950]  ( .D(c[958]), .CLK(clk), .RST(rst), .Q(c[950]) );
  DFF \sreg_reg[949]  ( .D(c[957]), .CLK(clk), .RST(rst), .Q(c[949]) );
  DFF \sreg_reg[948]  ( .D(c[956]), .CLK(clk), .RST(rst), .Q(c[948]) );
  DFF \sreg_reg[947]  ( .D(c[955]), .CLK(clk), .RST(rst), .Q(c[947]) );
  DFF \sreg_reg[946]  ( .D(c[954]), .CLK(clk), .RST(rst), .Q(c[946]) );
  DFF \sreg_reg[945]  ( .D(c[953]), .CLK(clk), .RST(rst), .Q(c[945]) );
  DFF \sreg_reg[944]  ( .D(c[952]), .CLK(clk), .RST(rst), .Q(c[944]) );
  DFF \sreg_reg[943]  ( .D(c[951]), .CLK(clk), .RST(rst), .Q(c[943]) );
  DFF \sreg_reg[942]  ( .D(c[950]), .CLK(clk), .RST(rst), .Q(c[942]) );
  DFF \sreg_reg[941]  ( .D(c[949]), .CLK(clk), .RST(rst), .Q(c[941]) );
  DFF \sreg_reg[940]  ( .D(c[948]), .CLK(clk), .RST(rst), .Q(c[940]) );
  DFF \sreg_reg[939]  ( .D(c[947]), .CLK(clk), .RST(rst), .Q(c[939]) );
  DFF \sreg_reg[938]  ( .D(c[946]), .CLK(clk), .RST(rst), .Q(c[938]) );
  DFF \sreg_reg[937]  ( .D(c[945]), .CLK(clk), .RST(rst), .Q(c[937]) );
  DFF \sreg_reg[936]  ( .D(c[944]), .CLK(clk), .RST(rst), .Q(c[936]) );
  DFF \sreg_reg[935]  ( .D(c[943]), .CLK(clk), .RST(rst), .Q(c[935]) );
  DFF \sreg_reg[934]  ( .D(c[942]), .CLK(clk), .RST(rst), .Q(c[934]) );
  DFF \sreg_reg[933]  ( .D(c[941]), .CLK(clk), .RST(rst), .Q(c[933]) );
  DFF \sreg_reg[932]  ( .D(c[940]), .CLK(clk), .RST(rst), .Q(c[932]) );
  DFF \sreg_reg[931]  ( .D(c[939]), .CLK(clk), .RST(rst), .Q(c[931]) );
  DFF \sreg_reg[930]  ( .D(c[938]), .CLK(clk), .RST(rst), .Q(c[930]) );
  DFF \sreg_reg[929]  ( .D(c[937]), .CLK(clk), .RST(rst), .Q(c[929]) );
  DFF \sreg_reg[928]  ( .D(c[936]), .CLK(clk), .RST(rst), .Q(c[928]) );
  DFF \sreg_reg[927]  ( .D(c[935]), .CLK(clk), .RST(rst), .Q(c[927]) );
  DFF \sreg_reg[926]  ( .D(c[934]), .CLK(clk), .RST(rst), .Q(c[926]) );
  DFF \sreg_reg[925]  ( .D(c[933]), .CLK(clk), .RST(rst), .Q(c[925]) );
  DFF \sreg_reg[924]  ( .D(c[932]), .CLK(clk), .RST(rst), .Q(c[924]) );
  DFF \sreg_reg[923]  ( .D(c[931]), .CLK(clk), .RST(rst), .Q(c[923]) );
  DFF \sreg_reg[922]  ( .D(c[930]), .CLK(clk), .RST(rst), .Q(c[922]) );
  DFF \sreg_reg[921]  ( .D(c[929]), .CLK(clk), .RST(rst), .Q(c[921]) );
  DFF \sreg_reg[920]  ( .D(c[928]), .CLK(clk), .RST(rst), .Q(c[920]) );
  DFF \sreg_reg[919]  ( .D(c[927]), .CLK(clk), .RST(rst), .Q(c[919]) );
  DFF \sreg_reg[918]  ( .D(c[926]), .CLK(clk), .RST(rst), .Q(c[918]) );
  DFF \sreg_reg[917]  ( .D(c[925]), .CLK(clk), .RST(rst), .Q(c[917]) );
  DFF \sreg_reg[916]  ( .D(c[924]), .CLK(clk), .RST(rst), .Q(c[916]) );
  DFF \sreg_reg[915]  ( .D(c[923]), .CLK(clk), .RST(rst), .Q(c[915]) );
  DFF \sreg_reg[914]  ( .D(c[922]), .CLK(clk), .RST(rst), .Q(c[914]) );
  DFF \sreg_reg[913]  ( .D(c[921]), .CLK(clk), .RST(rst), .Q(c[913]) );
  DFF \sreg_reg[912]  ( .D(c[920]), .CLK(clk), .RST(rst), .Q(c[912]) );
  DFF \sreg_reg[911]  ( .D(c[919]), .CLK(clk), .RST(rst), .Q(c[911]) );
  DFF \sreg_reg[910]  ( .D(c[918]), .CLK(clk), .RST(rst), .Q(c[910]) );
  DFF \sreg_reg[909]  ( .D(c[917]), .CLK(clk), .RST(rst), .Q(c[909]) );
  DFF \sreg_reg[908]  ( .D(c[916]), .CLK(clk), .RST(rst), .Q(c[908]) );
  DFF \sreg_reg[907]  ( .D(c[915]), .CLK(clk), .RST(rst), .Q(c[907]) );
  DFF \sreg_reg[906]  ( .D(c[914]), .CLK(clk), .RST(rst), .Q(c[906]) );
  DFF \sreg_reg[905]  ( .D(c[913]), .CLK(clk), .RST(rst), .Q(c[905]) );
  DFF \sreg_reg[904]  ( .D(c[912]), .CLK(clk), .RST(rst), .Q(c[904]) );
  DFF \sreg_reg[903]  ( .D(c[911]), .CLK(clk), .RST(rst), .Q(c[903]) );
  DFF \sreg_reg[902]  ( .D(c[910]), .CLK(clk), .RST(rst), .Q(c[902]) );
  DFF \sreg_reg[901]  ( .D(c[909]), .CLK(clk), .RST(rst), .Q(c[901]) );
  DFF \sreg_reg[900]  ( .D(c[908]), .CLK(clk), .RST(rst), .Q(c[900]) );
  DFF \sreg_reg[899]  ( .D(c[907]), .CLK(clk), .RST(rst), .Q(c[899]) );
  DFF \sreg_reg[898]  ( .D(c[906]), .CLK(clk), .RST(rst), .Q(c[898]) );
  DFF \sreg_reg[897]  ( .D(c[905]), .CLK(clk), .RST(rst), .Q(c[897]) );
  DFF \sreg_reg[896]  ( .D(c[904]), .CLK(clk), .RST(rst), .Q(c[896]) );
  DFF \sreg_reg[895]  ( .D(c[903]), .CLK(clk), .RST(rst), .Q(c[895]) );
  DFF \sreg_reg[894]  ( .D(c[902]), .CLK(clk), .RST(rst), .Q(c[894]) );
  DFF \sreg_reg[893]  ( .D(c[901]), .CLK(clk), .RST(rst), .Q(c[893]) );
  DFF \sreg_reg[892]  ( .D(c[900]), .CLK(clk), .RST(rst), .Q(c[892]) );
  DFF \sreg_reg[891]  ( .D(c[899]), .CLK(clk), .RST(rst), .Q(c[891]) );
  DFF \sreg_reg[890]  ( .D(c[898]), .CLK(clk), .RST(rst), .Q(c[890]) );
  DFF \sreg_reg[889]  ( .D(c[897]), .CLK(clk), .RST(rst), .Q(c[889]) );
  DFF \sreg_reg[888]  ( .D(c[896]), .CLK(clk), .RST(rst), .Q(c[888]) );
  DFF \sreg_reg[887]  ( .D(c[895]), .CLK(clk), .RST(rst), .Q(c[887]) );
  DFF \sreg_reg[886]  ( .D(c[894]), .CLK(clk), .RST(rst), .Q(c[886]) );
  DFF \sreg_reg[885]  ( .D(c[893]), .CLK(clk), .RST(rst), .Q(c[885]) );
  DFF \sreg_reg[884]  ( .D(c[892]), .CLK(clk), .RST(rst), .Q(c[884]) );
  DFF \sreg_reg[883]  ( .D(c[891]), .CLK(clk), .RST(rst), .Q(c[883]) );
  DFF \sreg_reg[882]  ( .D(c[890]), .CLK(clk), .RST(rst), .Q(c[882]) );
  DFF \sreg_reg[881]  ( .D(c[889]), .CLK(clk), .RST(rst), .Q(c[881]) );
  DFF \sreg_reg[880]  ( .D(c[888]), .CLK(clk), .RST(rst), .Q(c[880]) );
  DFF \sreg_reg[879]  ( .D(c[887]), .CLK(clk), .RST(rst), .Q(c[879]) );
  DFF \sreg_reg[878]  ( .D(c[886]), .CLK(clk), .RST(rst), .Q(c[878]) );
  DFF \sreg_reg[877]  ( .D(c[885]), .CLK(clk), .RST(rst), .Q(c[877]) );
  DFF \sreg_reg[876]  ( .D(c[884]), .CLK(clk), .RST(rst), .Q(c[876]) );
  DFF \sreg_reg[875]  ( .D(c[883]), .CLK(clk), .RST(rst), .Q(c[875]) );
  DFF \sreg_reg[874]  ( .D(c[882]), .CLK(clk), .RST(rst), .Q(c[874]) );
  DFF \sreg_reg[873]  ( .D(c[881]), .CLK(clk), .RST(rst), .Q(c[873]) );
  DFF \sreg_reg[872]  ( .D(c[880]), .CLK(clk), .RST(rst), .Q(c[872]) );
  DFF \sreg_reg[871]  ( .D(c[879]), .CLK(clk), .RST(rst), .Q(c[871]) );
  DFF \sreg_reg[870]  ( .D(c[878]), .CLK(clk), .RST(rst), .Q(c[870]) );
  DFF \sreg_reg[869]  ( .D(c[877]), .CLK(clk), .RST(rst), .Q(c[869]) );
  DFF \sreg_reg[868]  ( .D(c[876]), .CLK(clk), .RST(rst), .Q(c[868]) );
  DFF \sreg_reg[867]  ( .D(c[875]), .CLK(clk), .RST(rst), .Q(c[867]) );
  DFF \sreg_reg[866]  ( .D(c[874]), .CLK(clk), .RST(rst), .Q(c[866]) );
  DFF \sreg_reg[865]  ( .D(c[873]), .CLK(clk), .RST(rst), .Q(c[865]) );
  DFF \sreg_reg[864]  ( .D(c[872]), .CLK(clk), .RST(rst), .Q(c[864]) );
  DFF \sreg_reg[863]  ( .D(c[871]), .CLK(clk), .RST(rst), .Q(c[863]) );
  DFF \sreg_reg[862]  ( .D(c[870]), .CLK(clk), .RST(rst), .Q(c[862]) );
  DFF \sreg_reg[861]  ( .D(c[869]), .CLK(clk), .RST(rst), .Q(c[861]) );
  DFF \sreg_reg[860]  ( .D(c[868]), .CLK(clk), .RST(rst), .Q(c[860]) );
  DFF \sreg_reg[859]  ( .D(c[867]), .CLK(clk), .RST(rst), .Q(c[859]) );
  DFF \sreg_reg[858]  ( .D(c[866]), .CLK(clk), .RST(rst), .Q(c[858]) );
  DFF \sreg_reg[857]  ( .D(c[865]), .CLK(clk), .RST(rst), .Q(c[857]) );
  DFF \sreg_reg[856]  ( .D(c[864]), .CLK(clk), .RST(rst), .Q(c[856]) );
  DFF \sreg_reg[855]  ( .D(c[863]), .CLK(clk), .RST(rst), .Q(c[855]) );
  DFF \sreg_reg[854]  ( .D(c[862]), .CLK(clk), .RST(rst), .Q(c[854]) );
  DFF \sreg_reg[853]  ( .D(c[861]), .CLK(clk), .RST(rst), .Q(c[853]) );
  DFF \sreg_reg[852]  ( .D(c[860]), .CLK(clk), .RST(rst), .Q(c[852]) );
  DFF \sreg_reg[851]  ( .D(c[859]), .CLK(clk), .RST(rst), .Q(c[851]) );
  DFF \sreg_reg[850]  ( .D(c[858]), .CLK(clk), .RST(rst), .Q(c[850]) );
  DFF \sreg_reg[849]  ( .D(c[857]), .CLK(clk), .RST(rst), .Q(c[849]) );
  DFF \sreg_reg[848]  ( .D(c[856]), .CLK(clk), .RST(rst), .Q(c[848]) );
  DFF \sreg_reg[847]  ( .D(c[855]), .CLK(clk), .RST(rst), .Q(c[847]) );
  DFF \sreg_reg[846]  ( .D(c[854]), .CLK(clk), .RST(rst), .Q(c[846]) );
  DFF \sreg_reg[845]  ( .D(c[853]), .CLK(clk), .RST(rst), .Q(c[845]) );
  DFF \sreg_reg[844]  ( .D(c[852]), .CLK(clk), .RST(rst), .Q(c[844]) );
  DFF \sreg_reg[843]  ( .D(c[851]), .CLK(clk), .RST(rst), .Q(c[843]) );
  DFF \sreg_reg[842]  ( .D(c[850]), .CLK(clk), .RST(rst), .Q(c[842]) );
  DFF \sreg_reg[841]  ( .D(c[849]), .CLK(clk), .RST(rst), .Q(c[841]) );
  DFF \sreg_reg[840]  ( .D(c[848]), .CLK(clk), .RST(rst), .Q(c[840]) );
  DFF \sreg_reg[839]  ( .D(c[847]), .CLK(clk), .RST(rst), .Q(c[839]) );
  DFF \sreg_reg[838]  ( .D(c[846]), .CLK(clk), .RST(rst), .Q(c[838]) );
  DFF \sreg_reg[837]  ( .D(c[845]), .CLK(clk), .RST(rst), .Q(c[837]) );
  DFF \sreg_reg[836]  ( .D(c[844]), .CLK(clk), .RST(rst), .Q(c[836]) );
  DFF \sreg_reg[835]  ( .D(c[843]), .CLK(clk), .RST(rst), .Q(c[835]) );
  DFF \sreg_reg[834]  ( .D(c[842]), .CLK(clk), .RST(rst), .Q(c[834]) );
  DFF \sreg_reg[833]  ( .D(c[841]), .CLK(clk), .RST(rst), .Q(c[833]) );
  DFF \sreg_reg[832]  ( .D(c[840]), .CLK(clk), .RST(rst), .Q(c[832]) );
  DFF \sreg_reg[831]  ( .D(c[839]), .CLK(clk), .RST(rst), .Q(c[831]) );
  DFF \sreg_reg[830]  ( .D(c[838]), .CLK(clk), .RST(rst), .Q(c[830]) );
  DFF \sreg_reg[829]  ( .D(c[837]), .CLK(clk), .RST(rst), .Q(c[829]) );
  DFF \sreg_reg[828]  ( .D(c[836]), .CLK(clk), .RST(rst), .Q(c[828]) );
  DFF \sreg_reg[827]  ( .D(c[835]), .CLK(clk), .RST(rst), .Q(c[827]) );
  DFF \sreg_reg[826]  ( .D(c[834]), .CLK(clk), .RST(rst), .Q(c[826]) );
  DFF \sreg_reg[825]  ( .D(c[833]), .CLK(clk), .RST(rst), .Q(c[825]) );
  DFF \sreg_reg[824]  ( .D(c[832]), .CLK(clk), .RST(rst), .Q(c[824]) );
  DFF \sreg_reg[823]  ( .D(c[831]), .CLK(clk), .RST(rst), .Q(c[823]) );
  DFF \sreg_reg[822]  ( .D(c[830]), .CLK(clk), .RST(rst), .Q(c[822]) );
  DFF \sreg_reg[821]  ( .D(c[829]), .CLK(clk), .RST(rst), .Q(c[821]) );
  DFF \sreg_reg[820]  ( .D(c[828]), .CLK(clk), .RST(rst), .Q(c[820]) );
  DFF \sreg_reg[819]  ( .D(c[827]), .CLK(clk), .RST(rst), .Q(c[819]) );
  DFF \sreg_reg[818]  ( .D(c[826]), .CLK(clk), .RST(rst), .Q(c[818]) );
  DFF \sreg_reg[817]  ( .D(c[825]), .CLK(clk), .RST(rst), .Q(c[817]) );
  DFF \sreg_reg[816]  ( .D(c[824]), .CLK(clk), .RST(rst), .Q(c[816]) );
  DFF \sreg_reg[815]  ( .D(c[823]), .CLK(clk), .RST(rst), .Q(c[815]) );
  DFF \sreg_reg[814]  ( .D(c[822]), .CLK(clk), .RST(rst), .Q(c[814]) );
  DFF \sreg_reg[813]  ( .D(c[821]), .CLK(clk), .RST(rst), .Q(c[813]) );
  DFF \sreg_reg[812]  ( .D(c[820]), .CLK(clk), .RST(rst), .Q(c[812]) );
  DFF \sreg_reg[811]  ( .D(c[819]), .CLK(clk), .RST(rst), .Q(c[811]) );
  DFF \sreg_reg[810]  ( .D(c[818]), .CLK(clk), .RST(rst), .Q(c[810]) );
  DFF \sreg_reg[809]  ( .D(c[817]), .CLK(clk), .RST(rst), .Q(c[809]) );
  DFF \sreg_reg[808]  ( .D(c[816]), .CLK(clk), .RST(rst), .Q(c[808]) );
  DFF \sreg_reg[807]  ( .D(c[815]), .CLK(clk), .RST(rst), .Q(c[807]) );
  DFF \sreg_reg[806]  ( .D(c[814]), .CLK(clk), .RST(rst), .Q(c[806]) );
  DFF \sreg_reg[805]  ( .D(c[813]), .CLK(clk), .RST(rst), .Q(c[805]) );
  DFF \sreg_reg[804]  ( .D(c[812]), .CLK(clk), .RST(rst), .Q(c[804]) );
  DFF \sreg_reg[803]  ( .D(c[811]), .CLK(clk), .RST(rst), .Q(c[803]) );
  DFF \sreg_reg[802]  ( .D(c[810]), .CLK(clk), .RST(rst), .Q(c[802]) );
  DFF \sreg_reg[801]  ( .D(c[809]), .CLK(clk), .RST(rst), .Q(c[801]) );
  DFF \sreg_reg[800]  ( .D(c[808]), .CLK(clk), .RST(rst), .Q(c[800]) );
  DFF \sreg_reg[799]  ( .D(c[807]), .CLK(clk), .RST(rst), .Q(c[799]) );
  DFF \sreg_reg[798]  ( .D(c[806]), .CLK(clk), .RST(rst), .Q(c[798]) );
  DFF \sreg_reg[797]  ( .D(c[805]), .CLK(clk), .RST(rst), .Q(c[797]) );
  DFF \sreg_reg[796]  ( .D(c[804]), .CLK(clk), .RST(rst), .Q(c[796]) );
  DFF \sreg_reg[795]  ( .D(c[803]), .CLK(clk), .RST(rst), .Q(c[795]) );
  DFF \sreg_reg[794]  ( .D(c[802]), .CLK(clk), .RST(rst), .Q(c[794]) );
  DFF \sreg_reg[793]  ( .D(c[801]), .CLK(clk), .RST(rst), .Q(c[793]) );
  DFF \sreg_reg[792]  ( .D(c[800]), .CLK(clk), .RST(rst), .Q(c[792]) );
  DFF \sreg_reg[791]  ( .D(c[799]), .CLK(clk), .RST(rst), .Q(c[791]) );
  DFF \sreg_reg[790]  ( .D(c[798]), .CLK(clk), .RST(rst), .Q(c[790]) );
  DFF \sreg_reg[789]  ( .D(c[797]), .CLK(clk), .RST(rst), .Q(c[789]) );
  DFF \sreg_reg[788]  ( .D(c[796]), .CLK(clk), .RST(rst), .Q(c[788]) );
  DFF \sreg_reg[787]  ( .D(c[795]), .CLK(clk), .RST(rst), .Q(c[787]) );
  DFF \sreg_reg[786]  ( .D(c[794]), .CLK(clk), .RST(rst), .Q(c[786]) );
  DFF \sreg_reg[785]  ( .D(c[793]), .CLK(clk), .RST(rst), .Q(c[785]) );
  DFF \sreg_reg[784]  ( .D(c[792]), .CLK(clk), .RST(rst), .Q(c[784]) );
  DFF \sreg_reg[783]  ( .D(c[791]), .CLK(clk), .RST(rst), .Q(c[783]) );
  DFF \sreg_reg[782]  ( .D(c[790]), .CLK(clk), .RST(rst), .Q(c[782]) );
  DFF \sreg_reg[781]  ( .D(c[789]), .CLK(clk), .RST(rst), .Q(c[781]) );
  DFF \sreg_reg[780]  ( .D(c[788]), .CLK(clk), .RST(rst), .Q(c[780]) );
  DFF \sreg_reg[779]  ( .D(c[787]), .CLK(clk), .RST(rst), .Q(c[779]) );
  DFF \sreg_reg[778]  ( .D(c[786]), .CLK(clk), .RST(rst), .Q(c[778]) );
  DFF \sreg_reg[777]  ( .D(c[785]), .CLK(clk), .RST(rst), .Q(c[777]) );
  DFF \sreg_reg[776]  ( .D(c[784]), .CLK(clk), .RST(rst), .Q(c[776]) );
  DFF \sreg_reg[775]  ( .D(c[783]), .CLK(clk), .RST(rst), .Q(c[775]) );
  DFF \sreg_reg[774]  ( .D(c[782]), .CLK(clk), .RST(rst), .Q(c[774]) );
  DFF \sreg_reg[773]  ( .D(c[781]), .CLK(clk), .RST(rst), .Q(c[773]) );
  DFF \sreg_reg[772]  ( .D(c[780]), .CLK(clk), .RST(rst), .Q(c[772]) );
  DFF \sreg_reg[771]  ( .D(c[779]), .CLK(clk), .RST(rst), .Q(c[771]) );
  DFF \sreg_reg[770]  ( .D(c[778]), .CLK(clk), .RST(rst), .Q(c[770]) );
  DFF \sreg_reg[769]  ( .D(c[777]), .CLK(clk), .RST(rst), .Q(c[769]) );
  DFF \sreg_reg[768]  ( .D(c[776]), .CLK(clk), .RST(rst), .Q(c[768]) );
  DFF \sreg_reg[767]  ( .D(c[775]), .CLK(clk), .RST(rst), .Q(c[767]) );
  DFF \sreg_reg[766]  ( .D(c[774]), .CLK(clk), .RST(rst), .Q(c[766]) );
  DFF \sreg_reg[765]  ( .D(c[773]), .CLK(clk), .RST(rst), .Q(c[765]) );
  DFF \sreg_reg[764]  ( .D(c[772]), .CLK(clk), .RST(rst), .Q(c[764]) );
  DFF \sreg_reg[763]  ( .D(c[771]), .CLK(clk), .RST(rst), .Q(c[763]) );
  DFF \sreg_reg[762]  ( .D(c[770]), .CLK(clk), .RST(rst), .Q(c[762]) );
  DFF \sreg_reg[761]  ( .D(c[769]), .CLK(clk), .RST(rst), .Q(c[761]) );
  DFF \sreg_reg[760]  ( .D(c[768]), .CLK(clk), .RST(rst), .Q(c[760]) );
  DFF \sreg_reg[759]  ( .D(c[767]), .CLK(clk), .RST(rst), .Q(c[759]) );
  DFF \sreg_reg[758]  ( .D(c[766]), .CLK(clk), .RST(rst), .Q(c[758]) );
  DFF \sreg_reg[757]  ( .D(c[765]), .CLK(clk), .RST(rst), .Q(c[757]) );
  DFF \sreg_reg[756]  ( .D(c[764]), .CLK(clk), .RST(rst), .Q(c[756]) );
  DFF \sreg_reg[755]  ( .D(c[763]), .CLK(clk), .RST(rst), .Q(c[755]) );
  DFF \sreg_reg[754]  ( .D(c[762]), .CLK(clk), .RST(rst), .Q(c[754]) );
  DFF \sreg_reg[753]  ( .D(c[761]), .CLK(clk), .RST(rst), .Q(c[753]) );
  DFF \sreg_reg[752]  ( .D(c[760]), .CLK(clk), .RST(rst), .Q(c[752]) );
  DFF \sreg_reg[751]  ( .D(c[759]), .CLK(clk), .RST(rst), .Q(c[751]) );
  DFF \sreg_reg[750]  ( .D(c[758]), .CLK(clk), .RST(rst), .Q(c[750]) );
  DFF \sreg_reg[749]  ( .D(c[757]), .CLK(clk), .RST(rst), .Q(c[749]) );
  DFF \sreg_reg[748]  ( .D(c[756]), .CLK(clk), .RST(rst), .Q(c[748]) );
  DFF \sreg_reg[747]  ( .D(c[755]), .CLK(clk), .RST(rst), .Q(c[747]) );
  DFF \sreg_reg[746]  ( .D(c[754]), .CLK(clk), .RST(rst), .Q(c[746]) );
  DFF \sreg_reg[745]  ( .D(c[753]), .CLK(clk), .RST(rst), .Q(c[745]) );
  DFF \sreg_reg[744]  ( .D(c[752]), .CLK(clk), .RST(rst), .Q(c[744]) );
  DFF \sreg_reg[743]  ( .D(c[751]), .CLK(clk), .RST(rst), .Q(c[743]) );
  DFF \sreg_reg[742]  ( .D(c[750]), .CLK(clk), .RST(rst), .Q(c[742]) );
  DFF \sreg_reg[741]  ( .D(c[749]), .CLK(clk), .RST(rst), .Q(c[741]) );
  DFF \sreg_reg[740]  ( .D(c[748]), .CLK(clk), .RST(rst), .Q(c[740]) );
  DFF \sreg_reg[739]  ( .D(c[747]), .CLK(clk), .RST(rst), .Q(c[739]) );
  DFF \sreg_reg[738]  ( .D(c[746]), .CLK(clk), .RST(rst), .Q(c[738]) );
  DFF \sreg_reg[737]  ( .D(c[745]), .CLK(clk), .RST(rst), .Q(c[737]) );
  DFF \sreg_reg[736]  ( .D(c[744]), .CLK(clk), .RST(rst), .Q(c[736]) );
  DFF \sreg_reg[735]  ( .D(c[743]), .CLK(clk), .RST(rst), .Q(c[735]) );
  DFF \sreg_reg[734]  ( .D(c[742]), .CLK(clk), .RST(rst), .Q(c[734]) );
  DFF \sreg_reg[733]  ( .D(c[741]), .CLK(clk), .RST(rst), .Q(c[733]) );
  DFF \sreg_reg[732]  ( .D(c[740]), .CLK(clk), .RST(rst), .Q(c[732]) );
  DFF \sreg_reg[731]  ( .D(c[739]), .CLK(clk), .RST(rst), .Q(c[731]) );
  DFF \sreg_reg[730]  ( .D(c[738]), .CLK(clk), .RST(rst), .Q(c[730]) );
  DFF \sreg_reg[729]  ( .D(c[737]), .CLK(clk), .RST(rst), .Q(c[729]) );
  DFF \sreg_reg[728]  ( .D(c[736]), .CLK(clk), .RST(rst), .Q(c[728]) );
  DFF \sreg_reg[727]  ( .D(c[735]), .CLK(clk), .RST(rst), .Q(c[727]) );
  DFF \sreg_reg[726]  ( .D(c[734]), .CLK(clk), .RST(rst), .Q(c[726]) );
  DFF \sreg_reg[725]  ( .D(c[733]), .CLK(clk), .RST(rst), .Q(c[725]) );
  DFF \sreg_reg[724]  ( .D(c[732]), .CLK(clk), .RST(rst), .Q(c[724]) );
  DFF \sreg_reg[723]  ( .D(c[731]), .CLK(clk), .RST(rst), .Q(c[723]) );
  DFF \sreg_reg[722]  ( .D(c[730]), .CLK(clk), .RST(rst), .Q(c[722]) );
  DFF \sreg_reg[721]  ( .D(c[729]), .CLK(clk), .RST(rst), .Q(c[721]) );
  DFF \sreg_reg[720]  ( .D(c[728]), .CLK(clk), .RST(rst), .Q(c[720]) );
  DFF \sreg_reg[719]  ( .D(c[727]), .CLK(clk), .RST(rst), .Q(c[719]) );
  DFF \sreg_reg[718]  ( .D(c[726]), .CLK(clk), .RST(rst), .Q(c[718]) );
  DFF \sreg_reg[717]  ( .D(c[725]), .CLK(clk), .RST(rst), .Q(c[717]) );
  DFF \sreg_reg[716]  ( .D(c[724]), .CLK(clk), .RST(rst), .Q(c[716]) );
  DFF \sreg_reg[715]  ( .D(c[723]), .CLK(clk), .RST(rst), .Q(c[715]) );
  DFF \sreg_reg[714]  ( .D(c[722]), .CLK(clk), .RST(rst), .Q(c[714]) );
  DFF \sreg_reg[713]  ( .D(c[721]), .CLK(clk), .RST(rst), .Q(c[713]) );
  DFF \sreg_reg[712]  ( .D(c[720]), .CLK(clk), .RST(rst), .Q(c[712]) );
  DFF \sreg_reg[711]  ( .D(c[719]), .CLK(clk), .RST(rst), .Q(c[711]) );
  DFF \sreg_reg[710]  ( .D(c[718]), .CLK(clk), .RST(rst), .Q(c[710]) );
  DFF \sreg_reg[709]  ( .D(c[717]), .CLK(clk), .RST(rst), .Q(c[709]) );
  DFF \sreg_reg[708]  ( .D(c[716]), .CLK(clk), .RST(rst), .Q(c[708]) );
  DFF \sreg_reg[707]  ( .D(c[715]), .CLK(clk), .RST(rst), .Q(c[707]) );
  DFF \sreg_reg[706]  ( .D(c[714]), .CLK(clk), .RST(rst), .Q(c[706]) );
  DFF \sreg_reg[705]  ( .D(c[713]), .CLK(clk), .RST(rst), .Q(c[705]) );
  DFF \sreg_reg[704]  ( .D(c[712]), .CLK(clk), .RST(rst), .Q(c[704]) );
  DFF \sreg_reg[703]  ( .D(c[711]), .CLK(clk), .RST(rst), .Q(c[703]) );
  DFF \sreg_reg[702]  ( .D(c[710]), .CLK(clk), .RST(rst), .Q(c[702]) );
  DFF \sreg_reg[701]  ( .D(c[709]), .CLK(clk), .RST(rst), .Q(c[701]) );
  DFF \sreg_reg[700]  ( .D(c[708]), .CLK(clk), .RST(rst), .Q(c[700]) );
  DFF \sreg_reg[699]  ( .D(c[707]), .CLK(clk), .RST(rst), .Q(c[699]) );
  DFF \sreg_reg[698]  ( .D(c[706]), .CLK(clk), .RST(rst), .Q(c[698]) );
  DFF \sreg_reg[697]  ( .D(c[705]), .CLK(clk), .RST(rst), .Q(c[697]) );
  DFF \sreg_reg[696]  ( .D(c[704]), .CLK(clk), .RST(rst), .Q(c[696]) );
  DFF \sreg_reg[695]  ( .D(c[703]), .CLK(clk), .RST(rst), .Q(c[695]) );
  DFF \sreg_reg[694]  ( .D(c[702]), .CLK(clk), .RST(rst), .Q(c[694]) );
  DFF \sreg_reg[693]  ( .D(c[701]), .CLK(clk), .RST(rst), .Q(c[693]) );
  DFF \sreg_reg[692]  ( .D(c[700]), .CLK(clk), .RST(rst), .Q(c[692]) );
  DFF \sreg_reg[691]  ( .D(c[699]), .CLK(clk), .RST(rst), .Q(c[691]) );
  DFF \sreg_reg[690]  ( .D(c[698]), .CLK(clk), .RST(rst), .Q(c[690]) );
  DFF \sreg_reg[689]  ( .D(c[697]), .CLK(clk), .RST(rst), .Q(c[689]) );
  DFF \sreg_reg[688]  ( .D(c[696]), .CLK(clk), .RST(rst), .Q(c[688]) );
  DFF \sreg_reg[687]  ( .D(c[695]), .CLK(clk), .RST(rst), .Q(c[687]) );
  DFF \sreg_reg[686]  ( .D(c[694]), .CLK(clk), .RST(rst), .Q(c[686]) );
  DFF \sreg_reg[685]  ( .D(c[693]), .CLK(clk), .RST(rst), .Q(c[685]) );
  DFF \sreg_reg[684]  ( .D(c[692]), .CLK(clk), .RST(rst), .Q(c[684]) );
  DFF \sreg_reg[683]  ( .D(c[691]), .CLK(clk), .RST(rst), .Q(c[683]) );
  DFF \sreg_reg[682]  ( .D(c[690]), .CLK(clk), .RST(rst), .Q(c[682]) );
  DFF \sreg_reg[681]  ( .D(c[689]), .CLK(clk), .RST(rst), .Q(c[681]) );
  DFF \sreg_reg[680]  ( .D(c[688]), .CLK(clk), .RST(rst), .Q(c[680]) );
  DFF \sreg_reg[679]  ( .D(c[687]), .CLK(clk), .RST(rst), .Q(c[679]) );
  DFF \sreg_reg[678]  ( .D(c[686]), .CLK(clk), .RST(rst), .Q(c[678]) );
  DFF \sreg_reg[677]  ( .D(c[685]), .CLK(clk), .RST(rst), .Q(c[677]) );
  DFF \sreg_reg[676]  ( .D(c[684]), .CLK(clk), .RST(rst), .Q(c[676]) );
  DFF \sreg_reg[675]  ( .D(c[683]), .CLK(clk), .RST(rst), .Q(c[675]) );
  DFF \sreg_reg[674]  ( .D(c[682]), .CLK(clk), .RST(rst), .Q(c[674]) );
  DFF \sreg_reg[673]  ( .D(c[681]), .CLK(clk), .RST(rst), .Q(c[673]) );
  DFF \sreg_reg[672]  ( .D(c[680]), .CLK(clk), .RST(rst), .Q(c[672]) );
  DFF \sreg_reg[671]  ( .D(c[679]), .CLK(clk), .RST(rst), .Q(c[671]) );
  DFF \sreg_reg[670]  ( .D(c[678]), .CLK(clk), .RST(rst), .Q(c[670]) );
  DFF \sreg_reg[669]  ( .D(c[677]), .CLK(clk), .RST(rst), .Q(c[669]) );
  DFF \sreg_reg[668]  ( .D(c[676]), .CLK(clk), .RST(rst), .Q(c[668]) );
  DFF \sreg_reg[667]  ( .D(c[675]), .CLK(clk), .RST(rst), .Q(c[667]) );
  DFF \sreg_reg[666]  ( .D(c[674]), .CLK(clk), .RST(rst), .Q(c[666]) );
  DFF \sreg_reg[665]  ( .D(c[673]), .CLK(clk), .RST(rst), .Q(c[665]) );
  DFF \sreg_reg[664]  ( .D(c[672]), .CLK(clk), .RST(rst), .Q(c[664]) );
  DFF \sreg_reg[663]  ( .D(c[671]), .CLK(clk), .RST(rst), .Q(c[663]) );
  DFF \sreg_reg[662]  ( .D(c[670]), .CLK(clk), .RST(rst), .Q(c[662]) );
  DFF \sreg_reg[661]  ( .D(c[669]), .CLK(clk), .RST(rst), .Q(c[661]) );
  DFF \sreg_reg[660]  ( .D(c[668]), .CLK(clk), .RST(rst), .Q(c[660]) );
  DFF \sreg_reg[659]  ( .D(c[667]), .CLK(clk), .RST(rst), .Q(c[659]) );
  DFF \sreg_reg[658]  ( .D(c[666]), .CLK(clk), .RST(rst), .Q(c[658]) );
  DFF \sreg_reg[657]  ( .D(c[665]), .CLK(clk), .RST(rst), .Q(c[657]) );
  DFF \sreg_reg[656]  ( .D(c[664]), .CLK(clk), .RST(rst), .Q(c[656]) );
  DFF \sreg_reg[655]  ( .D(c[663]), .CLK(clk), .RST(rst), .Q(c[655]) );
  DFF \sreg_reg[654]  ( .D(c[662]), .CLK(clk), .RST(rst), .Q(c[654]) );
  DFF \sreg_reg[653]  ( .D(c[661]), .CLK(clk), .RST(rst), .Q(c[653]) );
  DFF \sreg_reg[652]  ( .D(c[660]), .CLK(clk), .RST(rst), .Q(c[652]) );
  DFF \sreg_reg[651]  ( .D(c[659]), .CLK(clk), .RST(rst), .Q(c[651]) );
  DFF \sreg_reg[650]  ( .D(c[658]), .CLK(clk), .RST(rst), .Q(c[650]) );
  DFF \sreg_reg[649]  ( .D(c[657]), .CLK(clk), .RST(rst), .Q(c[649]) );
  DFF \sreg_reg[648]  ( .D(c[656]), .CLK(clk), .RST(rst), .Q(c[648]) );
  DFF \sreg_reg[647]  ( .D(c[655]), .CLK(clk), .RST(rst), .Q(c[647]) );
  DFF \sreg_reg[646]  ( .D(c[654]), .CLK(clk), .RST(rst), .Q(c[646]) );
  DFF \sreg_reg[645]  ( .D(c[653]), .CLK(clk), .RST(rst), .Q(c[645]) );
  DFF \sreg_reg[644]  ( .D(c[652]), .CLK(clk), .RST(rst), .Q(c[644]) );
  DFF \sreg_reg[643]  ( .D(c[651]), .CLK(clk), .RST(rst), .Q(c[643]) );
  DFF \sreg_reg[642]  ( .D(c[650]), .CLK(clk), .RST(rst), .Q(c[642]) );
  DFF \sreg_reg[641]  ( .D(c[649]), .CLK(clk), .RST(rst), .Q(c[641]) );
  DFF \sreg_reg[640]  ( .D(c[648]), .CLK(clk), .RST(rst), .Q(c[640]) );
  DFF \sreg_reg[639]  ( .D(c[647]), .CLK(clk), .RST(rst), .Q(c[639]) );
  DFF \sreg_reg[638]  ( .D(c[646]), .CLK(clk), .RST(rst), .Q(c[638]) );
  DFF \sreg_reg[637]  ( .D(c[645]), .CLK(clk), .RST(rst), .Q(c[637]) );
  DFF \sreg_reg[636]  ( .D(c[644]), .CLK(clk), .RST(rst), .Q(c[636]) );
  DFF \sreg_reg[635]  ( .D(c[643]), .CLK(clk), .RST(rst), .Q(c[635]) );
  DFF \sreg_reg[634]  ( .D(c[642]), .CLK(clk), .RST(rst), .Q(c[634]) );
  DFF \sreg_reg[633]  ( .D(c[641]), .CLK(clk), .RST(rst), .Q(c[633]) );
  DFF \sreg_reg[632]  ( .D(c[640]), .CLK(clk), .RST(rst), .Q(c[632]) );
  DFF \sreg_reg[631]  ( .D(c[639]), .CLK(clk), .RST(rst), .Q(c[631]) );
  DFF \sreg_reg[630]  ( .D(c[638]), .CLK(clk), .RST(rst), .Q(c[630]) );
  DFF \sreg_reg[629]  ( .D(c[637]), .CLK(clk), .RST(rst), .Q(c[629]) );
  DFF \sreg_reg[628]  ( .D(c[636]), .CLK(clk), .RST(rst), .Q(c[628]) );
  DFF \sreg_reg[627]  ( .D(c[635]), .CLK(clk), .RST(rst), .Q(c[627]) );
  DFF \sreg_reg[626]  ( .D(c[634]), .CLK(clk), .RST(rst), .Q(c[626]) );
  DFF \sreg_reg[625]  ( .D(c[633]), .CLK(clk), .RST(rst), .Q(c[625]) );
  DFF \sreg_reg[624]  ( .D(c[632]), .CLK(clk), .RST(rst), .Q(c[624]) );
  DFF \sreg_reg[623]  ( .D(c[631]), .CLK(clk), .RST(rst), .Q(c[623]) );
  DFF \sreg_reg[622]  ( .D(c[630]), .CLK(clk), .RST(rst), .Q(c[622]) );
  DFF \sreg_reg[621]  ( .D(c[629]), .CLK(clk), .RST(rst), .Q(c[621]) );
  DFF \sreg_reg[620]  ( .D(c[628]), .CLK(clk), .RST(rst), .Q(c[620]) );
  DFF \sreg_reg[619]  ( .D(c[627]), .CLK(clk), .RST(rst), .Q(c[619]) );
  DFF \sreg_reg[618]  ( .D(c[626]), .CLK(clk), .RST(rst), .Q(c[618]) );
  DFF \sreg_reg[617]  ( .D(c[625]), .CLK(clk), .RST(rst), .Q(c[617]) );
  DFF \sreg_reg[616]  ( .D(c[624]), .CLK(clk), .RST(rst), .Q(c[616]) );
  DFF \sreg_reg[615]  ( .D(c[623]), .CLK(clk), .RST(rst), .Q(c[615]) );
  DFF \sreg_reg[614]  ( .D(c[622]), .CLK(clk), .RST(rst), .Q(c[614]) );
  DFF \sreg_reg[613]  ( .D(c[621]), .CLK(clk), .RST(rst), .Q(c[613]) );
  DFF \sreg_reg[612]  ( .D(c[620]), .CLK(clk), .RST(rst), .Q(c[612]) );
  DFF \sreg_reg[611]  ( .D(c[619]), .CLK(clk), .RST(rst), .Q(c[611]) );
  DFF \sreg_reg[610]  ( .D(c[618]), .CLK(clk), .RST(rst), .Q(c[610]) );
  DFF \sreg_reg[609]  ( .D(c[617]), .CLK(clk), .RST(rst), .Q(c[609]) );
  DFF \sreg_reg[608]  ( .D(c[616]), .CLK(clk), .RST(rst), .Q(c[608]) );
  DFF \sreg_reg[607]  ( .D(c[615]), .CLK(clk), .RST(rst), .Q(c[607]) );
  DFF \sreg_reg[606]  ( .D(c[614]), .CLK(clk), .RST(rst), .Q(c[606]) );
  DFF \sreg_reg[605]  ( .D(c[613]), .CLK(clk), .RST(rst), .Q(c[605]) );
  DFF \sreg_reg[604]  ( .D(c[612]), .CLK(clk), .RST(rst), .Q(c[604]) );
  DFF \sreg_reg[603]  ( .D(c[611]), .CLK(clk), .RST(rst), .Q(c[603]) );
  DFF \sreg_reg[602]  ( .D(c[610]), .CLK(clk), .RST(rst), .Q(c[602]) );
  DFF \sreg_reg[601]  ( .D(c[609]), .CLK(clk), .RST(rst), .Q(c[601]) );
  DFF \sreg_reg[600]  ( .D(c[608]), .CLK(clk), .RST(rst), .Q(c[600]) );
  DFF \sreg_reg[599]  ( .D(c[607]), .CLK(clk), .RST(rst), .Q(c[599]) );
  DFF \sreg_reg[598]  ( .D(c[606]), .CLK(clk), .RST(rst), .Q(c[598]) );
  DFF \sreg_reg[597]  ( .D(c[605]), .CLK(clk), .RST(rst), .Q(c[597]) );
  DFF \sreg_reg[596]  ( .D(c[604]), .CLK(clk), .RST(rst), .Q(c[596]) );
  DFF \sreg_reg[595]  ( .D(c[603]), .CLK(clk), .RST(rst), .Q(c[595]) );
  DFF \sreg_reg[594]  ( .D(c[602]), .CLK(clk), .RST(rst), .Q(c[594]) );
  DFF \sreg_reg[593]  ( .D(c[601]), .CLK(clk), .RST(rst), .Q(c[593]) );
  DFF \sreg_reg[592]  ( .D(c[600]), .CLK(clk), .RST(rst), .Q(c[592]) );
  DFF \sreg_reg[591]  ( .D(c[599]), .CLK(clk), .RST(rst), .Q(c[591]) );
  DFF \sreg_reg[590]  ( .D(c[598]), .CLK(clk), .RST(rst), .Q(c[590]) );
  DFF \sreg_reg[589]  ( .D(c[597]), .CLK(clk), .RST(rst), .Q(c[589]) );
  DFF \sreg_reg[588]  ( .D(c[596]), .CLK(clk), .RST(rst), .Q(c[588]) );
  DFF \sreg_reg[587]  ( .D(c[595]), .CLK(clk), .RST(rst), .Q(c[587]) );
  DFF \sreg_reg[586]  ( .D(c[594]), .CLK(clk), .RST(rst), .Q(c[586]) );
  DFF \sreg_reg[585]  ( .D(c[593]), .CLK(clk), .RST(rst), .Q(c[585]) );
  DFF \sreg_reg[584]  ( .D(c[592]), .CLK(clk), .RST(rst), .Q(c[584]) );
  DFF \sreg_reg[583]  ( .D(c[591]), .CLK(clk), .RST(rst), .Q(c[583]) );
  DFF \sreg_reg[582]  ( .D(c[590]), .CLK(clk), .RST(rst), .Q(c[582]) );
  DFF \sreg_reg[581]  ( .D(c[589]), .CLK(clk), .RST(rst), .Q(c[581]) );
  DFF \sreg_reg[580]  ( .D(c[588]), .CLK(clk), .RST(rst), .Q(c[580]) );
  DFF \sreg_reg[579]  ( .D(c[587]), .CLK(clk), .RST(rst), .Q(c[579]) );
  DFF \sreg_reg[578]  ( .D(c[586]), .CLK(clk), .RST(rst), .Q(c[578]) );
  DFF \sreg_reg[577]  ( .D(c[585]), .CLK(clk), .RST(rst), .Q(c[577]) );
  DFF \sreg_reg[576]  ( .D(c[584]), .CLK(clk), .RST(rst), .Q(c[576]) );
  DFF \sreg_reg[575]  ( .D(c[583]), .CLK(clk), .RST(rst), .Q(c[575]) );
  DFF \sreg_reg[574]  ( .D(c[582]), .CLK(clk), .RST(rst), .Q(c[574]) );
  DFF \sreg_reg[573]  ( .D(c[581]), .CLK(clk), .RST(rst), .Q(c[573]) );
  DFF \sreg_reg[572]  ( .D(c[580]), .CLK(clk), .RST(rst), .Q(c[572]) );
  DFF \sreg_reg[571]  ( .D(c[579]), .CLK(clk), .RST(rst), .Q(c[571]) );
  DFF \sreg_reg[570]  ( .D(c[578]), .CLK(clk), .RST(rst), .Q(c[570]) );
  DFF \sreg_reg[569]  ( .D(c[577]), .CLK(clk), .RST(rst), .Q(c[569]) );
  DFF \sreg_reg[568]  ( .D(c[576]), .CLK(clk), .RST(rst), .Q(c[568]) );
  DFF \sreg_reg[567]  ( .D(c[575]), .CLK(clk), .RST(rst), .Q(c[567]) );
  DFF \sreg_reg[566]  ( .D(c[574]), .CLK(clk), .RST(rst), .Q(c[566]) );
  DFF \sreg_reg[565]  ( .D(c[573]), .CLK(clk), .RST(rst), .Q(c[565]) );
  DFF \sreg_reg[564]  ( .D(c[572]), .CLK(clk), .RST(rst), .Q(c[564]) );
  DFF \sreg_reg[563]  ( .D(c[571]), .CLK(clk), .RST(rst), .Q(c[563]) );
  DFF \sreg_reg[562]  ( .D(c[570]), .CLK(clk), .RST(rst), .Q(c[562]) );
  DFF \sreg_reg[561]  ( .D(c[569]), .CLK(clk), .RST(rst), .Q(c[561]) );
  DFF \sreg_reg[560]  ( .D(c[568]), .CLK(clk), .RST(rst), .Q(c[560]) );
  DFF \sreg_reg[559]  ( .D(c[567]), .CLK(clk), .RST(rst), .Q(c[559]) );
  DFF \sreg_reg[558]  ( .D(c[566]), .CLK(clk), .RST(rst), .Q(c[558]) );
  DFF \sreg_reg[557]  ( .D(c[565]), .CLK(clk), .RST(rst), .Q(c[557]) );
  DFF \sreg_reg[556]  ( .D(c[564]), .CLK(clk), .RST(rst), .Q(c[556]) );
  DFF \sreg_reg[555]  ( .D(c[563]), .CLK(clk), .RST(rst), .Q(c[555]) );
  DFF \sreg_reg[554]  ( .D(c[562]), .CLK(clk), .RST(rst), .Q(c[554]) );
  DFF \sreg_reg[553]  ( .D(c[561]), .CLK(clk), .RST(rst), .Q(c[553]) );
  DFF \sreg_reg[552]  ( .D(c[560]), .CLK(clk), .RST(rst), .Q(c[552]) );
  DFF \sreg_reg[551]  ( .D(c[559]), .CLK(clk), .RST(rst), .Q(c[551]) );
  DFF \sreg_reg[550]  ( .D(c[558]), .CLK(clk), .RST(rst), .Q(c[550]) );
  DFF \sreg_reg[549]  ( .D(c[557]), .CLK(clk), .RST(rst), .Q(c[549]) );
  DFF \sreg_reg[548]  ( .D(c[556]), .CLK(clk), .RST(rst), .Q(c[548]) );
  DFF \sreg_reg[547]  ( .D(c[555]), .CLK(clk), .RST(rst), .Q(c[547]) );
  DFF \sreg_reg[546]  ( .D(c[554]), .CLK(clk), .RST(rst), .Q(c[546]) );
  DFF \sreg_reg[545]  ( .D(c[553]), .CLK(clk), .RST(rst), .Q(c[545]) );
  DFF \sreg_reg[544]  ( .D(c[552]), .CLK(clk), .RST(rst), .Q(c[544]) );
  DFF \sreg_reg[543]  ( .D(c[551]), .CLK(clk), .RST(rst), .Q(c[543]) );
  DFF \sreg_reg[542]  ( .D(c[550]), .CLK(clk), .RST(rst), .Q(c[542]) );
  DFF \sreg_reg[541]  ( .D(c[549]), .CLK(clk), .RST(rst), .Q(c[541]) );
  DFF \sreg_reg[540]  ( .D(c[548]), .CLK(clk), .RST(rst), .Q(c[540]) );
  DFF \sreg_reg[539]  ( .D(c[547]), .CLK(clk), .RST(rst), .Q(c[539]) );
  DFF \sreg_reg[538]  ( .D(c[546]), .CLK(clk), .RST(rst), .Q(c[538]) );
  DFF \sreg_reg[537]  ( .D(c[545]), .CLK(clk), .RST(rst), .Q(c[537]) );
  DFF \sreg_reg[536]  ( .D(c[544]), .CLK(clk), .RST(rst), .Q(c[536]) );
  DFF \sreg_reg[535]  ( .D(c[543]), .CLK(clk), .RST(rst), .Q(c[535]) );
  DFF \sreg_reg[534]  ( .D(c[542]), .CLK(clk), .RST(rst), .Q(c[534]) );
  DFF \sreg_reg[533]  ( .D(c[541]), .CLK(clk), .RST(rst), .Q(c[533]) );
  DFF \sreg_reg[532]  ( .D(c[540]), .CLK(clk), .RST(rst), .Q(c[532]) );
  DFF \sreg_reg[531]  ( .D(c[539]), .CLK(clk), .RST(rst), .Q(c[531]) );
  DFF \sreg_reg[530]  ( .D(c[538]), .CLK(clk), .RST(rst), .Q(c[530]) );
  DFF \sreg_reg[529]  ( .D(c[537]), .CLK(clk), .RST(rst), .Q(c[529]) );
  DFF \sreg_reg[528]  ( .D(c[536]), .CLK(clk), .RST(rst), .Q(c[528]) );
  DFF \sreg_reg[527]  ( .D(c[535]), .CLK(clk), .RST(rst), .Q(c[527]) );
  DFF \sreg_reg[526]  ( .D(c[534]), .CLK(clk), .RST(rst), .Q(c[526]) );
  DFF \sreg_reg[525]  ( .D(c[533]), .CLK(clk), .RST(rst), .Q(c[525]) );
  DFF \sreg_reg[524]  ( .D(c[532]), .CLK(clk), .RST(rst), .Q(c[524]) );
  DFF \sreg_reg[523]  ( .D(c[531]), .CLK(clk), .RST(rst), .Q(c[523]) );
  DFF \sreg_reg[522]  ( .D(c[530]), .CLK(clk), .RST(rst), .Q(c[522]) );
  DFF \sreg_reg[521]  ( .D(c[529]), .CLK(clk), .RST(rst), .Q(c[521]) );
  DFF \sreg_reg[520]  ( .D(c[528]), .CLK(clk), .RST(rst), .Q(c[520]) );
  DFF \sreg_reg[519]  ( .D(c[527]), .CLK(clk), .RST(rst), .Q(c[519]) );
  DFF \sreg_reg[518]  ( .D(c[526]), .CLK(clk), .RST(rst), .Q(c[518]) );
  DFF \sreg_reg[517]  ( .D(c[525]), .CLK(clk), .RST(rst), .Q(c[517]) );
  DFF \sreg_reg[516]  ( .D(c[524]), .CLK(clk), .RST(rst), .Q(c[516]) );
  DFF \sreg_reg[515]  ( .D(c[523]), .CLK(clk), .RST(rst), .Q(c[515]) );
  DFF \sreg_reg[514]  ( .D(c[522]), .CLK(clk), .RST(rst), .Q(c[514]) );
  DFF \sreg_reg[513]  ( .D(c[521]), .CLK(clk), .RST(rst), .Q(c[513]) );
  DFF \sreg_reg[512]  ( .D(c[520]), .CLK(clk), .RST(rst), .Q(c[512]) );
  DFF \sreg_reg[511]  ( .D(c[519]), .CLK(clk), .RST(rst), .Q(c[511]) );
  DFF \sreg_reg[510]  ( .D(c[518]), .CLK(clk), .RST(rst), .Q(c[510]) );
  DFF \sreg_reg[509]  ( .D(c[517]), .CLK(clk), .RST(rst), .Q(c[509]) );
  DFF \sreg_reg[508]  ( .D(c[516]), .CLK(clk), .RST(rst), .Q(c[508]) );
  DFF \sreg_reg[507]  ( .D(c[515]), .CLK(clk), .RST(rst), .Q(c[507]) );
  DFF \sreg_reg[506]  ( .D(c[514]), .CLK(clk), .RST(rst), .Q(c[506]) );
  DFF \sreg_reg[505]  ( .D(c[513]), .CLK(clk), .RST(rst), .Q(c[505]) );
  DFF \sreg_reg[504]  ( .D(c[512]), .CLK(clk), .RST(rst), .Q(c[504]) );
  DFF \sreg_reg[503]  ( .D(c[511]), .CLK(clk), .RST(rst), .Q(c[503]) );
  DFF \sreg_reg[502]  ( .D(c[510]), .CLK(clk), .RST(rst), .Q(c[502]) );
  DFF \sreg_reg[501]  ( .D(c[509]), .CLK(clk), .RST(rst), .Q(c[501]) );
  DFF \sreg_reg[500]  ( .D(c[508]), .CLK(clk), .RST(rst), .Q(c[500]) );
  DFF \sreg_reg[499]  ( .D(c[507]), .CLK(clk), .RST(rst), .Q(c[499]) );
  DFF \sreg_reg[498]  ( .D(c[506]), .CLK(clk), .RST(rst), .Q(c[498]) );
  DFF \sreg_reg[497]  ( .D(c[505]), .CLK(clk), .RST(rst), .Q(c[497]) );
  DFF \sreg_reg[496]  ( .D(c[504]), .CLK(clk), .RST(rst), .Q(c[496]) );
  DFF \sreg_reg[495]  ( .D(c[503]), .CLK(clk), .RST(rst), .Q(c[495]) );
  DFF \sreg_reg[494]  ( .D(c[502]), .CLK(clk), .RST(rst), .Q(c[494]) );
  DFF \sreg_reg[493]  ( .D(c[501]), .CLK(clk), .RST(rst), .Q(c[493]) );
  DFF \sreg_reg[492]  ( .D(c[500]), .CLK(clk), .RST(rst), .Q(c[492]) );
  DFF \sreg_reg[491]  ( .D(c[499]), .CLK(clk), .RST(rst), .Q(c[491]) );
  DFF \sreg_reg[490]  ( .D(c[498]), .CLK(clk), .RST(rst), .Q(c[490]) );
  DFF \sreg_reg[489]  ( .D(c[497]), .CLK(clk), .RST(rst), .Q(c[489]) );
  DFF \sreg_reg[488]  ( .D(c[496]), .CLK(clk), .RST(rst), .Q(c[488]) );
  DFF \sreg_reg[487]  ( .D(c[495]), .CLK(clk), .RST(rst), .Q(c[487]) );
  DFF \sreg_reg[486]  ( .D(c[494]), .CLK(clk), .RST(rst), .Q(c[486]) );
  DFF \sreg_reg[485]  ( .D(c[493]), .CLK(clk), .RST(rst), .Q(c[485]) );
  DFF \sreg_reg[484]  ( .D(c[492]), .CLK(clk), .RST(rst), .Q(c[484]) );
  DFF \sreg_reg[483]  ( .D(c[491]), .CLK(clk), .RST(rst), .Q(c[483]) );
  DFF \sreg_reg[482]  ( .D(c[490]), .CLK(clk), .RST(rst), .Q(c[482]) );
  DFF \sreg_reg[481]  ( .D(c[489]), .CLK(clk), .RST(rst), .Q(c[481]) );
  DFF \sreg_reg[480]  ( .D(c[488]), .CLK(clk), .RST(rst), .Q(c[480]) );
  DFF \sreg_reg[479]  ( .D(c[487]), .CLK(clk), .RST(rst), .Q(c[479]) );
  DFF \sreg_reg[478]  ( .D(c[486]), .CLK(clk), .RST(rst), .Q(c[478]) );
  DFF \sreg_reg[477]  ( .D(c[485]), .CLK(clk), .RST(rst), .Q(c[477]) );
  DFF \sreg_reg[476]  ( .D(c[484]), .CLK(clk), .RST(rst), .Q(c[476]) );
  DFF \sreg_reg[475]  ( .D(c[483]), .CLK(clk), .RST(rst), .Q(c[475]) );
  DFF \sreg_reg[474]  ( .D(c[482]), .CLK(clk), .RST(rst), .Q(c[474]) );
  DFF \sreg_reg[473]  ( .D(c[481]), .CLK(clk), .RST(rst), .Q(c[473]) );
  DFF \sreg_reg[472]  ( .D(c[480]), .CLK(clk), .RST(rst), .Q(c[472]) );
  DFF \sreg_reg[471]  ( .D(c[479]), .CLK(clk), .RST(rst), .Q(c[471]) );
  DFF \sreg_reg[470]  ( .D(c[478]), .CLK(clk), .RST(rst), .Q(c[470]) );
  DFF \sreg_reg[469]  ( .D(c[477]), .CLK(clk), .RST(rst), .Q(c[469]) );
  DFF \sreg_reg[468]  ( .D(c[476]), .CLK(clk), .RST(rst), .Q(c[468]) );
  DFF \sreg_reg[467]  ( .D(c[475]), .CLK(clk), .RST(rst), .Q(c[467]) );
  DFF \sreg_reg[466]  ( .D(c[474]), .CLK(clk), .RST(rst), .Q(c[466]) );
  DFF \sreg_reg[465]  ( .D(c[473]), .CLK(clk), .RST(rst), .Q(c[465]) );
  DFF \sreg_reg[464]  ( .D(c[472]), .CLK(clk), .RST(rst), .Q(c[464]) );
  DFF \sreg_reg[463]  ( .D(c[471]), .CLK(clk), .RST(rst), .Q(c[463]) );
  DFF \sreg_reg[462]  ( .D(c[470]), .CLK(clk), .RST(rst), .Q(c[462]) );
  DFF \sreg_reg[461]  ( .D(c[469]), .CLK(clk), .RST(rst), .Q(c[461]) );
  DFF \sreg_reg[460]  ( .D(c[468]), .CLK(clk), .RST(rst), .Q(c[460]) );
  DFF \sreg_reg[459]  ( .D(c[467]), .CLK(clk), .RST(rst), .Q(c[459]) );
  DFF \sreg_reg[458]  ( .D(c[466]), .CLK(clk), .RST(rst), .Q(c[458]) );
  DFF \sreg_reg[457]  ( .D(c[465]), .CLK(clk), .RST(rst), .Q(c[457]) );
  DFF \sreg_reg[456]  ( .D(c[464]), .CLK(clk), .RST(rst), .Q(c[456]) );
  DFF \sreg_reg[455]  ( .D(c[463]), .CLK(clk), .RST(rst), .Q(c[455]) );
  DFF \sreg_reg[454]  ( .D(c[462]), .CLK(clk), .RST(rst), .Q(c[454]) );
  DFF \sreg_reg[453]  ( .D(c[461]), .CLK(clk), .RST(rst), .Q(c[453]) );
  DFF \sreg_reg[452]  ( .D(c[460]), .CLK(clk), .RST(rst), .Q(c[452]) );
  DFF \sreg_reg[451]  ( .D(c[459]), .CLK(clk), .RST(rst), .Q(c[451]) );
  DFF \sreg_reg[450]  ( .D(c[458]), .CLK(clk), .RST(rst), .Q(c[450]) );
  DFF \sreg_reg[449]  ( .D(c[457]), .CLK(clk), .RST(rst), .Q(c[449]) );
  DFF \sreg_reg[448]  ( .D(c[456]), .CLK(clk), .RST(rst), .Q(c[448]) );
  DFF \sreg_reg[447]  ( .D(c[455]), .CLK(clk), .RST(rst), .Q(c[447]) );
  DFF \sreg_reg[446]  ( .D(c[454]), .CLK(clk), .RST(rst), .Q(c[446]) );
  DFF \sreg_reg[445]  ( .D(c[453]), .CLK(clk), .RST(rst), .Q(c[445]) );
  DFF \sreg_reg[444]  ( .D(c[452]), .CLK(clk), .RST(rst), .Q(c[444]) );
  DFF \sreg_reg[443]  ( .D(c[451]), .CLK(clk), .RST(rst), .Q(c[443]) );
  DFF \sreg_reg[442]  ( .D(c[450]), .CLK(clk), .RST(rst), .Q(c[442]) );
  DFF \sreg_reg[441]  ( .D(c[449]), .CLK(clk), .RST(rst), .Q(c[441]) );
  DFF \sreg_reg[440]  ( .D(c[448]), .CLK(clk), .RST(rst), .Q(c[440]) );
  DFF \sreg_reg[439]  ( .D(c[447]), .CLK(clk), .RST(rst), .Q(c[439]) );
  DFF \sreg_reg[438]  ( .D(c[446]), .CLK(clk), .RST(rst), .Q(c[438]) );
  DFF \sreg_reg[437]  ( .D(c[445]), .CLK(clk), .RST(rst), .Q(c[437]) );
  DFF \sreg_reg[436]  ( .D(c[444]), .CLK(clk), .RST(rst), .Q(c[436]) );
  DFF \sreg_reg[435]  ( .D(c[443]), .CLK(clk), .RST(rst), .Q(c[435]) );
  DFF \sreg_reg[434]  ( .D(c[442]), .CLK(clk), .RST(rst), .Q(c[434]) );
  DFF \sreg_reg[433]  ( .D(c[441]), .CLK(clk), .RST(rst), .Q(c[433]) );
  DFF \sreg_reg[432]  ( .D(c[440]), .CLK(clk), .RST(rst), .Q(c[432]) );
  DFF \sreg_reg[431]  ( .D(c[439]), .CLK(clk), .RST(rst), .Q(c[431]) );
  DFF \sreg_reg[430]  ( .D(c[438]), .CLK(clk), .RST(rst), .Q(c[430]) );
  DFF \sreg_reg[429]  ( .D(c[437]), .CLK(clk), .RST(rst), .Q(c[429]) );
  DFF \sreg_reg[428]  ( .D(c[436]), .CLK(clk), .RST(rst), .Q(c[428]) );
  DFF \sreg_reg[427]  ( .D(c[435]), .CLK(clk), .RST(rst), .Q(c[427]) );
  DFF \sreg_reg[426]  ( .D(c[434]), .CLK(clk), .RST(rst), .Q(c[426]) );
  DFF \sreg_reg[425]  ( .D(c[433]), .CLK(clk), .RST(rst), .Q(c[425]) );
  DFF \sreg_reg[424]  ( .D(c[432]), .CLK(clk), .RST(rst), .Q(c[424]) );
  DFF \sreg_reg[423]  ( .D(c[431]), .CLK(clk), .RST(rst), .Q(c[423]) );
  DFF \sreg_reg[422]  ( .D(c[430]), .CLK(clk), .RST(rst), .Q(c[422]) );
  DFF \sreg_reg[421]  ( .D(c[429]), .CLK(clk), .RST(rst), .Q(c[421]) );
  DFF \sreg_reg[420]  ( .D(c[428]), .CLK(clk), .RST(rst), .Q(c[420]) );
  DFF \sreg_reg[419]  ( .D(c[427]), .CLK(clk), .RST(rst), .Q(c[419]) );
  DFF \sreg_reg[418]  ( .D(c[426]), .CLK(clk), .RST(rst), .Q(c[418]) );
  DFF \sreg_reg[417]  ( .D(c[425]), .CLK(clk), .RST(rst), .Q(c[417]) );
  DFF \sreg_reg[416]  ( .D(c[424]), .CLK(clk), .RST(rst), .Q(c[416]) );
  DFF \sreg_reg[415]  ( .D(c[423]), .CLK(clk), .RST(rst), .Q(c[415]) );
  DFF \sreg_reg[414]  ( .D(c[422]), .CLK(clk), .RST(rst), .Q(c[414]) );
  DFF \sreg_reg[413]  ( .D(c[421]), .CLK(clk), .RST(rst), .Q(c[413]) );
  DFF \sreg_reg[412]  ( .D(c[420]), .CLK(clk), .RST(rst), .Q(c[412]) );
  DFF \sreg_reg[411]  ( .D(c[419]), .CLK(clk), .RST(rst), .Q(c[411]) );
  DFF \sreg_reg[410]  ( .D(c[418]), .CLK(clk), .RST(rst), .Q(c[410]) );
  DFF \sreg_reg[409]  ( .D(c[417]), .CLK(clk), .RST(rst), .Q(c[409]) );
  DFF \sreg_reg[408]  ( .D(c[416]), .CLK(clk), .RST(rst), .Q(c[408]) );
  DFF \sreg_reg[407]  ( .D(c[415]), .CLK(clk), .RST(rst), .Q(c[407]) );
  DFF \sreg_reg[406]  ( .D(c[414]), .CLK(clk), .RST(rst), .Q(c[406]) );
  DFF \sreg_reg[405]  ( .D(c[413]), .CLK(clk), .RST(rst), .Q(c[405]) );
  DFF \sreg_reg[404]  ( .D(c[412]), .CLK(clk), .RST(rst), .Q(c[404]) );
  DFF \sreg_reg[403]  ( .D(c[411]), .CLK(clk), .RST(rst), .Q(c[403]) );
  DFF \sreg_reg[402]  ( .D(c[410]), .CLK(clk), .RST(rst), .Q(c[402]) );
  DFF \sreg_reg[401]  ( .D(c[409]), .CLK(clk), .RST(rst), .Q(c[401]) );
  DFF \sreg_reg[400]  ( .D(c[408]), .CLK(clk), .RST(rst), .Q(c[400]) );
  DFF \sreg_reg[399]  ( .D(c[407]), .CLK(clk), .RST(rst), .Q(c[399]) );
  DFF \sreg_reg[398]  ( .D(c[406]), .CLK(clk), .RST(rst), .Q(c[398]) );
  DFF \sreg_reg[397]  ( .D(c[405]), .CLK(clk), .RST(rst), .Q(c[397]) );
  DFF \sreg_reg[396]  ( .D(c[404]), .CLK(clk), .RST(rst), .Q(c[396]) );
  DFF \sreg_reg[395]  ( .D(c[403]), .CLK(clk), .RST(rst), .Q(c[395]) );
  DFF \sreg_reg[394]  ( .D(c[402]), .CLK(clk), .RST(rst), .Q(c[394]) );
  DFF \sreg_reg[393]  ( .D(c[401]), .CLK(clk), .RST(rst), .Q(c[393]) );
  DFF \sreg_reg[392]  ( .D(c[400]), .CLK(clk), .RST(rst), .Q(c[392]) );
  DFF \sreg_reg[391]  ( .D(c[399]), .CLK(clk), .RST(rst), .Q(c[391]) );
  DFF \sreg_reg[390]  ( .D(c[398]), .CLK(clk), .RST(rst), .Q(c[390]) );
  DFF \sreg_reg[389]  ( .D(c[397]), .CLK(clk), .RST(rst), .Q(c[389]) );
  DFF \sreg_reg[388]  ( .D(c[396]), .CLK(clk), .RST(rst), .Q(c[388]) );
  DFF \sreg_reg[387]  ( .D(c[395]), .CLK(clk), .RST(rst), .Q(c[387]) );
  DFF \sreg_reg[386]  ( .D(c[394]), .CLK(clk), .RST(rst), .Q(c[386]) );
  DFF \sreg_reg[385]  ( .D(c[393]), .CLK(clk), .RST(rst), .Q(c[385]) );
  DFF \sreg_reg[384]  ( .D(c[392]), .CLK(clk), .RST(rst), .Q(c[384]) );
  DFF \sreg_reg[383]  ( .D(c[391]), .CLK(clk), .RST(rst), .Q(c[383]) );
  DFF \sreg_reg[382]  ( .D(c[390]), .CLK(clk), .RST(rst), .Q(c[382]) );
  DFF \sreg_reg[381]  ( .D(c[389]), .CLK(clk), .RST(rst), .Q(c[381]) );
  DFF \sreg_reg[380]  ( .D(c[388]), .CLK(clk), .RST(rst), .Q(c[380]) );
  DFF \sreg_reg[379]  ( .D(c[387]), .CLK(clk), .RST(rst), .Q(c[379]) );
  DFF \sreg_reg[378]  ( .D(c[386]), .CLK(clk), .RST(rst), .Q(c[378]) );
  DFF \sreg_reg[377]  ( .D(c[385]), .CLK(clk), .RST(rst), .Q(c[377]) );
  DFF \sreg_reg[376]  ( .D(c[384]), .CLK(clk), .RST(rst), .Q(c[376]) );
  DFF \sreg_reg[375]  ( .D(c[383]), .CLK(clk), .RST(rst), .Q(c[375]) );
  DFF \sreg_reg[374]  ( .D(c[382]), .CLK(clk), .RST(rst), .Q(c[374]) );
  DFF \sreg_reg[373]  ( .D(c[381]), .CLK(clk), .RST(rst), .Q(c[373]) );
  DFF \sreg_reg[372]  ( .D(c[380]), .CLK(clk), .RST(rst), .Q(c[372]) );
  DFF \sreg_reg[371]  ( .D(c[379]), .CLK(clk), .RST(rst), .Q(c[371]) );
  DFF \sreg_reg[370]  ( .D(c[378]), .CLK(clk), .RST(rst), .Q(c[370]) );
  DFF \sreg_reg[369]  ( .D(c[377]), .CLK(clk), .RST(rst), .Q(c[369]) );
  DFF \sreg_reg[368]  ( .D(c[376]), .CLK(clk), .RST(rst), .Q(c[368]) );
  DFF \sreg_reg[367]  ( .D(c[375]), .CLK(clk), .RST(rst), .Q(c[367]) );
  DFF \sreg_reg[366]  ( .D(c[374]), .CLK(clk), .RST(rst), .Q(c[366]) );
  DFF \sreg_reg[365]  ( .D(c[373]), .CLK(clk), .RST(rst), .Q(c[365]) );
  DFF \sreg_reg[364]  ( .D(c[372]), .CLK(clk), .RST(rst), .Q(c[364]) );
  DFF \sreg_reg[363]  ( .D(c[371]), .CLK(clk), .RST(rst), .Q(c[363]) );
  DFF \sreg_reg[362]  ( .D(c[370]), .CLK(clk), .RST(rst), .Q(c[362]) );
  DFF \sreg_reg[361]  ( .D(c[369]), .CLK(clk), .RST(rst), .Q(c[361]) );
  DFF \sreg_reg[360]  ( .D(c[368]), .CLK(clk), .RST(rst), .Q(c[360]) );
  DFF \sreg_reg[359]  ( .D(c[367]), .CLK(clk), .RST(rst), .Q(c[359]) );
  DFF \sreg_reg[358]  ( .D(c[366]), .CLK(clk), .RST(rst), .Q(c[358]) );
  DFF \sreg_reg[357]  ( .D(c[365]), .CLK(clk), .RST(rst), .Q(c[357]) );
  DFF \sreg_reg[356]  ( .D(c[364]), .CLK(clk), .RST(rst), .Q(c[356]) );
  DFF \sreg_reg[355]  ( .D(c[363]), .CLK(clk), .RST(rst), .Q(c[355]) );
  DFF \sreg_reg[354]  ( .D(c[362]), .CLK(clk), .RST(rst), .Q(c[354]) );
  DFF \sreg_reg[353]  ( .D(c[361]), .CLK(clk), .RST(rst), .Q(c[353]) );
  DFF \sreg_reg[352]  ( .D(c[360]), .CLK(clk), .RST(rst), .Q(c[352]) );
  DFF \sreg_reg[351]  ( .D(c[359]), .CLK(clk), .RST(rst), .Q(c[351]) );
  DFF \sreg_reg[350]  ( .D(c[358]), .CLK(clk), .RST(rst), .Q(c[350]) );
  DFF \sreg_reg[349]  ( .D(c[357]), .CLK(clk), .RST(rst), .Q(c[349]) );
  DFF \sreg_reg[348]  ( .D(c[356]), .CLK(clk), .RST(rst), .Q(c[348]) );
  DFF \sreg_reg[347]  ( .D(c[355]), .CLK(clk), .RST(rst), .Q(c[347]) );
  DFF \sreg_reg[346]  ( .D(c[354]), .CLK(clk), .RST(rst), .Q(c[346]) );
  DFF \sreg_reg[345]  ( .D(c[353]), .CLK(clk), .RST(rst), .Q(c[345]) );
  DFF \sreg_reg[344]  ( .D(c[352]), .CLK(clk), .RST(rst), .Q(c[344]) );
  DFF \sreg_reg[343]  ( .D(c[351]), .CLK(clk), .RST(rst), .Q(c[343]) );
  DFF \sreg_reg[342]  ( .D(c[350]), .CLK(clk), .RST(rst), .Q(c[342]) );
  DFF \sreg_reg[341]  ( .D(c[349]), .CLK(clk), .RST(rst), .Q(c[341]) );
  DFF \sreg_reg[340]  ( .D(c[348]), .CLK(clk), .RST(rst), .Q(c[340]) );
  DFF \sreg_reg[339]  ( .D(c[347]), .CLK(clk), .RST(rst), .Q(c[339]) );
  DFF \sreg_reg[338]  ( .D(c[346]), .CLK(clk), .RST(rst), .Q(c[338]) );
  DFF \sreg_reg[337]  ( .D(c[345]), .CLK(clk), .RST(rst), .Q(c[337]) );
  DFF \sreg_reg[336]  ( .D(c[344]), .CLK(clk), .RST(rst), .Q(c[336]) );
  DFF \sreg_reg[335]  ( .D(c[343]), .CLK(clk), .RST(rst), .Q(c[335]) );
  DFF \sreg_reg[334]  ( .D(c[342]), .CLK(clk), .RST(rst), .Q(c[334]) );
  DFF \sreg_reg[333]  ( .D(c[341]), .CLK(clk), .RST(rst), .Q(c[333]) );
  DFF \sreg_reg[332]  ( .D(c[340]), .CLK(clk), .RST(rst), .Q(c[332]) );
  DFF \sreg_reg[331]  ( .D(c[339]), .CLK(clk), .RST(rst), .Q(c[331]) );
  DFF \sreg_reg[330]  ( .D(c[338]), .CLK(clk), .RST(rst), .Q(c[330]) );
  DFF \sreg_reg[329]  ( .D(c[337]), .CLK(clk), .RST(rst), .Q(c[329]) );
  DFF \sreg_reg[328]  ( .D(c[336]), .CLK(clk), .RST(rst), .Q(c[328]) );
  DFF \sreg_reg[327]  ( .D(c[335]), .CLK(clk), .RST(rst), .Q(c[327]) );
  DFF \sreg_reg[326]  ( .D(c[334]), .CLK(clk), .RST(rst), .Q(c[326]) );
  DFF \sreg_reg[325]  ( .D(c[333]), .CLK(clk), .RST(rst), .Q(c[325]) );
  DFF \sreg_reg[324]  ( .D(c[332]), .CLK(clk), .RST(rst), .Q(c[324]) );
  DFF \sreg_reg[323]  ( .D(c[331]), .CLK(clk), .RST(rst), .Q(c[323]) );
  DFF \sreg_reg[322]  ( .D(c[330]), .CLK(clk), .RST(rst), .Q(c[322]) );
  DFF \sreg_reg[321]  ( .D(c[329]), .CLK(clk), .RST(rst), .Q(c[321]) );
  DFF \sreg_reg[320]  ( .D(c[328]), .CLK(clk), .RST(rst), .Q(c[320]) );
  DFF \sreg_reg[319]  ( .D(c[327]), .CLK(clk), .RST(rst), .Q(c[319]) );
  DFF \sreg_reg[318]  ( .D(c[326]), .CLK(clk), .RST(rst), .Q(c[318]) );
  DFF \sreg_reg[317]  ( .D(c[325]), .CLK(clk), .RST(rst), .Q(c[317]) );
  DFF \sreg_reg[316]  ( .D(c[324]), .CLK(clk), .RST(rst), .Q(c[316]) );
  DFF \sreg_reg[315]  ( .D(c[323]), .CLK(clk), .RST(rst), .Q(c[315]) );
  DFF \sreg_reg[314]  ( .D(c[322]), .CLK(clk), .RST(rst), .Q(c[314]) );
  DFF \sreg_reg[313]  ( .D(c[321]), .CLK(clk), .RST(rst), .Q(c[313]) );
  DFF \sreg_reg[312]  ( .D(c[320]), .CLK(clk), .RST(rst), .Q(c[312]) );
  DFF \sreg_reg[311]  ( .D(c[319]), .CLK(clk), .RST(rst), .Q(c[311]) );
  DFF \sreg_reg[310]  ( .D(c[318]), .CLK(clk), .RST(rst), .Q(c[310]) );
  DFF \sreg_reg[309]  ( .D(c[317]), .CLK(clk), .RST(rst), .Q(c[309]) );
  DFF \sreg_reg[308]  ( .D(c[316]), .CLK(clk), .RST(rst), .Q(c[308]) );
  DFF \sreg_reg[307]  ( .D(c[315]), .CLK(clk), .RST(rst), .Q(c[307]) );
  DFF \sreg_reg[306]  ( .D(c[314]), .CLK(clk), .RST(rst), .Q(c[306]) );
  DFF \sreg_reg[305]  ( .D(c[313]), .CLK(clk), .RST(rst), .Q(c[305]) );
  DFF \sreg_reg[304]  ( .D(c[312]), .CLK(clk), .RST(rst), .Q(c[304]) );
  DFF \sreg_reg[303]  ( .D(c[311]), .CLK(clk), .RST(rst), .Q(c[303]) );
  DFF \sreg_reg[302]  ( .D(c[310]), .CLK(clk), .RST(rst), .Q(c[302]) );
  DFF \sreg_reg[301]  ( .D(c[309]), .CLK(clk), .RST(rst), .Q(c[301]) );
  DFF \sreg_reg[300]  ( .D(c[308]), .CLK(clk), .RST(rst), .Q(c[300]) );
  DFF \sreg_reg[299]  ( .D(c[307]), .CLK(clk), .RST(rst), .Q(c[299]) );
  DFF \sreg_reg[298]  ( .D(c[306]), .CLK(clk), .RST(rst), .Q(c[298]) );
  DFF \sreg_reg[297]  ( .D(c[305]), .CLK(clk), .RST(rst), .Q(c[297]) );
  DFF \sreg_reg[296]  ( .D(c[304]), .CLK(clk), .RST(rst), .Q(c[296]) );
  DFF \sreg_reg[295]  ( .D(c[303]), .CLK(clk), .RST(rst), .Q(c[295]) );
  DFF \sreg_reg[294]  ( .D(c[302]), .CLK(clk), .RST(rst), .Q(c[294]) );
  DFF \sreg_reg[293]  ( .D(c[301]), .CLK(clk), .RST(rst), .Q(c[293]) );
  DFF \sreg_reg[292]  ( .D(c[300]), .CLK(clk), .RST(rst), .Q(c[292]) );
  DFF \sreg_reg[291]  ( .D(c[299]), .CLK(clk), .RST(rst), .Q(c[291]) );
  DFF \sreg_reg[290]  ( .D(c[298]), .CLK(clk), .RST(rst), .Q(c[290]) );
  DFF \sreg_reg[289]  ( .D(c[297]), .CLK(clk), .RST(rst), .Q(c[289]) );
  DFF \sreg_reg[288]  ( .D(c[296]), .CLK(clk), .RST(rst), .Q(c[288]) );
  DFF \sreg_reg[287]  ( .D(c[295]), .CLK(clk), .RST(rst), .Q(c[287]) );
  DFF \sreg_reg[286]  ( .D(c[294]), .CLK(clk), .RST(rst), .Q(c[286]) );
  DFF \sreg_reg[285]  ( .D(c[293]), .CLK(clk), .RST(rst), .Q(c[285]) );
  DFF \sreg_reg[284]  ( .D(c[292]), .CLK(clk), .RST(rst), .Q(c[284]) );
  DFF \sreg_reg[283]  ( .D(c[291]), .CLK(clk), .RST(rst), .Q(c[283]) );
  DFF \sreg_reg[282]  ( .D(c[290]), .CLK(clk), .RST(rst), .Q(c[282]) );
  DFF \sreg_reg[281]  ( .D(c[289]), .CLK(clk), .RST(rst), .Q(c[281]) );
  DFF \sreg_reg[280]  ( .D(c[288]), .CLK(clk), .RST(rst), .Q(c[280]) );
  DFF \sreg_reg[279]  ( .D(c[287]), .CLK(clk), .RST(rst), .Q(c[279]) );
  DFF \sreg_reg[278]  ( .D(c[286]), .CLK(clk), .RST(rst), .Q(c[278]) );
  DFF \sreg_reg[277]  ( .D(c[285]), .CLK(clk), .RST(rst), .Q(c[277]) );
  DFF \sreg_reg[276]  ( .D(c[284]), .CLK(clk), .RST(rst), .Q(c[276]) );
  DFF \sreg_reg[275]  ( .D(c[283]), .CLK(clk), .RST(rst), .Q(c[275]) );
  DFF \sreg_reg[274]  ( .D(c[282]), .CLK(clk), .RST(rst), .Q(c[274]) );
  DFF \sreg_reg[273]  ( .D(c[281]), .CLK(clk), .RST(rst), .Q(c[273]) );
  DFF \sreg_reg[272]  ( .D(c[280]), .CLK(clk), .RST(rst), .Q(c[272]) );
  DFF \sreg_reg[271]  ( .D(c[279]), .CLK(clk), .RST(rst), .Q(c[271]) );
  DFF \sreg_reg[270]  ( .D(c[278]), .CLK(clk), .RST(rst), .Q(c[270]) );
  DFF \sreg_reg[269]  ( .D(c[277]), .CLK(clk), .RST(rst), .Q(c[269]) );
  DFF \sreg_reg[268]  ( .D(c[276]), .CLK(clk), .RST(rst), .Q(c[268]) );
  DFF \sreg_reg[267]  ( .D(c[275]), .CLK(clk), .RST(rst), .Q(c[267]) );
  DFF \sreg_reg[266]  ( .D(c[274]), .CLK(clk), .RST(rst), .Q(c[266]) );
  DFF \sreg_reg[265]  ( .D(c[273]), .CLK(clk), .RST(rst), .Q(c[265]) );
  DFF \sreg_reg[264]  ( .D(c[272]), .CLK(clk), .RST(rst), .Q(c[264]) );
  DFF \sreg_reg[263]  ( .D(c[271]), .CLK(clk), .RST(rst), .Q(c[263]) );
  DFF \sreg_reg[262]  ( .D(c[270]), .CLK(clk), .RST(rst), .Q(c[262]) );
  DFF \sreg_reg[261]  ( .D(c[269]), .CLK(clk), .RST(rst), .Q(c[261]) );
  DFF \sreg_reg[260]  ( .D(c[268]), .CLK(clk), .RST(rst), .Q(c[260]) );
  DFF \sreg_reg[259]  ( .D(c[267]), .CLK(clk), .RST(rst), .Q(c[259]) );
  DFF \sreg_reg[258]  ( .D(c[266]), .CLK(clk), .RST(rst), .Q(c[258]) );
  DFF \sreg_reg[257]  ( .D(c[265]), .CLK(clk), .RST(rst), .Q(c[257]) );
  DFF \sreg_reg[256]  ( .D(c[264]), .CLK(clk), .RST(rst), .Q(c[256]) );
  DFF \sreg_reg[255]  ( .D(c[263]), .CLK(clk), .RST(rst), .Q(c[255]) );
  DFF \sreg_reg[254]  ( .D(c[262]), .CLK(clk), .RST(rst), .Q(c[254]) );
  DFF \sreg_reg[253]  ( .D(c[261]), .CLK(clk), .RST(rst), .Q(c[253]) );
  DFF \sreg_reg[252]  ( .D(c[260]), .CLK(clk), .RST(rst), .Q(c[252]) );
  DFF \sreg_reg[251]  ( .D(c[259]), .CLK(clk), .RST(rst), .Q(c[251]) );
  DFF \sreg_reg[250]  ( .D(c[258]), .CLK(clk), .RST(rst), .Q(c[250]) );
  DFF \sreg_reg[249]  ( .D(c[257]), .CLK(clk), .RST(rst), .Q(c[249]) );
  DFF \sreg_reg[248]  ( .D(c[256]), .CLK(clk), .RST(rst), .Q(c[248]) );
  DFF \sreg_reg[247]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[247]) );
  DFF \sreg_reg[246]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[246]) );
  DFF \sreg_reg[245]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[245]) );
  DFF \sreg_reg[244]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[244]) );
  DFF \sreg_reg[243]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[243]) );
  DFF \sreg_reg[242]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[242]) );
  DFF \sreg_reg[241]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[241]) );
  DFF \sreg_reg[240]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[240]) );
  DFF \sreg_reg[239]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[239]) );
  DFF \sreg_reg[238]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[238]) );
  DFF \sreg_reg[237]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[237]) );
  DFF \sreg_reg[236]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[236]) );
  DFF \sreg_reg[235]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[235]) );
  DFF \sreg_reg[234]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[234]) );
  DFF \sreg_reg[233]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[233]) );
  DFF \sreg_reg[232]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[232]) );
  DFF \sreg_reg[231]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[231]) );
  DFF \sreg_reg[230]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[230]) );
  DFF \sreg_reg[229]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[229]) );
  DFF \sreg_reg[228]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[228]) );
  DFF \sreg_reg[227]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[227]) );
  DFF \sreg_reg[226]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[226]) );
  DFF \sreg_reg[225]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[225]) );
  DFF \sreg_reg[224]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[224]) );
  DFF \sreg_reg[223]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[222]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[221]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[220]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[219]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[218]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[217]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[216]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[215]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[214]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[213]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[212]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[211]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[210]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[209]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[208]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[207]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[206]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[205]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[204]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[203]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[202]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[201]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[200]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[199]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[198]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[197]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[196]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[195]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[194]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[193]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[192]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[191]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[190]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[189]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[188]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[187]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[186]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[185]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[184]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[183]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[182]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[181]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[180]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[179]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[178]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[177]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[176]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[175]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[174]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[173]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[172]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[171]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[170]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[169]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[168]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[167]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[166]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[165]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[164]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[163]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[162]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[161]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[160]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[159]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[158]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[157]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[156]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[155]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[154]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[153]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[152]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[151]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[150]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[149]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[148]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[147]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[146]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[145]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[144]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[143]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[142]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[141]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[140]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[139]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[138]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[137]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[136]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[135]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[134]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[133]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[132]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[131]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[130]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[129]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[128]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[127]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[126]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[125]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[0]) );
  OR U11 ( .A(b[0]), .B(n42233), .Z(n1) );
  NAND U12 ( .A(n1), .B(b[1]), .Z(n42112) );
  NANDN U13 ( .A(n288), .B(n287), .Z(n296) );
  OR U14 ( .A(n340), .B(n341), .Z(n2) );
  NANDN U15 ( .A(n343), .B(n342), .Z(n3) );
  NAND U16 ( .A(n2), .B(n3), .Z(n350) );
  NANDN U17 ( .A(n286), .B(n285), .Z(n4) );
  NANDN U18 ( .A(n283), .B(n284), .Z(n5) );
  NAND U19 ( .A(n4), .B(n5), .Z(n298) );
  NANDN U20 ( .A(n42148), .B(n42149), .Z(n6) );
  NANDN U21 ( .A(n42147), .B(n42146), .Z(n7) );
  AND U22 ( .A(n6), .B(n7), .Z(n42156) );
  XNOR U23 ( .A(n42029), .B(n42030), .Z(n42032) );
  XOR U24 ( .A(b[1]), .B(b[2]), .Z(n42095) );
  XNOR U25 ( .A(n42111), .B(n42112), .Z(n42113) );
  OR U26 ( .A(n42208), .B(n42160), .Z(n8) );
  NAND U27 ( .A(n42159), .B(n42158), .Z(n9) );
  NAND U28 ( .A(n8), .B(n9), .Z(n42212) );
  NANDN U29 ( .A(n324), .B(n325), .Z(n10) );
  NANDN U30 ( .A(n326), .B(n327), .Z(n11) );
  NAND U31 ( .A(n10), .B(n11), .Z(n351) );
  NAND U32 ( .A(n42157), .B(n42156), .Z(n12) );
  XOR U33 ( .A(n42156), .B(n42157), .Z(n13) );
  NAND U34 ( .A(n13), .B(n42155), .Z(n14) );
  NAND U35 ( .A(n12), .B(n14), .Z(n42187) );
  IV U36 ( .A(b[0]), .Z(n15) );
  IV U37 ( .A(b[0]), .Z(n16) );
  IV U38 ( .A(b[0]), .Z(n17) );
  IV U39 ( .A(b[0]), .Z(n18) );
  IV U40 ( .A(b[0]), .Z(n19) );
  IV U41 ( .A(b[0]), .Z(n20) );
  IV U42 ( .A(b[0]), .Z(n21) );
  IV U43 ( .A(b[0]), .Z(n22) );
  IV U44 ( .A(b[0]), .Z(n23) );
  IV U45 ( .A(b[0]), .Z(n24) );
  IV U46 ( .A(b[0]), .Z(n25) );
  IV U47 ( .A(b[0]), .Z(n26) );
  IV U48 ( .A(b[0]), .Z(n27) );
  IV U49 ( .A(b[0]), .Z(n28) );
  IV U50 ( .A(b[0]), .Z(n29) );
  IV U51 ( .A(b[0]), .Z(n30) );
  IV U52 ( .A(b[0]), .Z(n31) );
  IV U53 ( .A(b[0]), .Z(n32) );
  IV U54 ( .A(b[0]), .Z(n33) );
  IV U55 ( .A(b[0]), .Z(n34) );
  IV U56 ( .A(b[0]), .Z(n35) );
  IV U57 ( .A(b[0]), .Z(n36) );
  IV U58 ( .A(b[0]), .Z(n37) );
  IV U59 ( .A(b[0]), .Z(n38) );
  IV U60 ( .A(b[0]), .Z(n39) );
  IV U61 ( .A(b[0]), .Z(n40) );
  IV U62 ( .A(b[0]), .Z(n41) );
  IV U63 ( .A(b[0]), .Z(n42) );
  IV U64 ( .A(b[0]), .Z(n43) );
  IV U65 ( .A(b[0]), .Z(n44) );
  IV U66 ( .A(b[0]), .Z(n45) );
  IV U67 ( .A(b[0]), .Z(n46) );
  IV U68 ( .A(b[0]), .Z(n47) );
  IV U69 ( .A(b[0]), .Z(n48) );
  IV U70 ( .A(b[0]), .Z(n49) );
  IV U71 ( .A(b[0]), .Z(n50) );
  IV U72 ( .A(b[0]), .Z(n51) );
  IV U73 ( .A(b[0]), .Z(n52) );
  IV U74 ( .A(b[0]), .Z(n53) );
  IV U75 ( .A(b[0]), .Z(n54) );
  IV U76 ( .A(b[0]), .Z(n55) );
  IV U77 ( .A(b[0]), .Z(n56) );
  IV U78 ( .A(b[0]), .Z(n57) );
  IV U79 ( .A(b[0]), .Z(n58) );
  IV U80 ( .A(b[0]), .Z(n59) );
  IV U81 ( .A(b[0]), .Z(n60) );
  IV U82 ( .A(b[0]), .Z(n61) );
  IV U83 ( .A(b[0]), .Z(n62) );
  IV U84 ( .A(b[0]), .Z(n63) );
  IV U85 ( .A(b[0]), .Z(n64) );
  IV U86 ( .A(b[0]), .Z(n65) );
  IV U87 ( .A(b[0]), .Z(n66) );
  IV U88 ( .A(b[0]), .Z(n67) );
  IV U89 ( .A(b[0]), .Z(n68) );
  IV U90 ( .A(b[0]), .Z(n69) );
  IV U91 ( .A(b[0]), .Z(n70) );
  IV U92 ( .A(b[0]), .Z(n71) );
  IV U93 ( .A(b[0]), .Z(n72) );
  IV U94 ( .A(b[0]), .Z(n73) );
  IV U95 ( .A(b[0]), .Z(n74) );
  IV U96 ( .A(b[0]), .Z(n75) );
  IV U97 ( .A(b[0]), .Z(n76) );
  IV U98 ( .A(b[0]), .Z(n77) );
  IV U99 ( .A(b[0]), .Z(n78) );
  IV U100 ( .A(b[0]), .Z(n79) );
  IV U101 ( .A(b[0]), .Z(n80) );
  IV U102 ( .A(b[0]), .Z(n81) );
  IV U103 ( .A(b[0]), .Z(n82) );
  IV U104 ( .A(b[0]), .Z(n83) );
  IV U105 ( .A(b[0]), .Z(n84) );
  IV U106 ( .A(b[0]), .Z(n85) );
  IV U107 ( .A(b[0]), .Z(n86) );
  IV U108 ( .A(b[0]), .Z(n87) );
  IV U109 ( .A(b[0]), .Z(n88) );
  IV U110 ( .A(b[0]), .Z(n89) );
  IV U111 ( .A(b[0]), .Z(n90) );
  IV U112 ( .A(b[0]), .Z(n91) );
  IV U113 ( .A(b[0]), .Z(n92) );
  IV U114 ( .A(b[0]), .Z(n93) );
  IV U115 ( .A(b[0]), .Z(n94) );
  IV U116 ( .A(b[0]), .Z(n95) );
  IV U117 ( .A(b[0]), .Z(n96) );
  IV U118 ( .A(b[0]), .Z(n97) );
  IV U119 ( .A(b[0]), .Z(n98) );
  IV U120 ( .A(b[0]), .Z(n99) );
  IV U121 ( .A(b[0]), .Z(n100) );
  IV U122 ( .A(b[0]), .Z(n101) );
  IV U123 ( .A(b[0]), .Z(n102) );
  IV U124 ( .A(b[0]), .Z(n103) );
  IV U125 ( .A(b[0]), .Z(n104) );
  IV U126 ( .A(b[0]), .Z(n105) );
  IV U127 ( .A(b[0]), .Z(n106) );
  IV U128 ( .A(b[0]), .Z(n107) );
  IV U129 ( .A(b[0]), .Z(n108) );
  IV U130 ( .A(b[0]), .Z(n109) );
  IV U131 ( .A(b[0]), .Z(n110) );
  IV U132 ( .A(b[0]), .Z(n111) );
  IV U133 ( .A(b[0]), .Z(n112) );
  IV U134 ( .A(b[0]), .Z(n113) );
  IV U135 ( .A(b[0]), .Z(n114) );
  IV U136 ( .A(b[0]), .Z(n115) );
  IV U137 ( .A(b[0]), .Z(n116) );
  IV U138 ( .A(b[0]), .Z(n117) );
  IV U139 ( .A(b[0]), .Z(n118) );
  IV U140 ( .A(b[0]), .Z(n119) );
  IV U141 ( .A(b[0]), .Z(n120) );
  IV U142 ( .A(b[0]), .Z(n121) );
  IV U143 ( .A(b[0]), .Z(n122) );
  IV U144 ( .A(b[0]), .Z(n123) );
  IV U145 ( .A(b[0]), .Z(n124) );
  IV U146 ( .A(b[0]), .Z(n125) );
  IV U147 ( .A(b[0]), .Z(n126) );
  IV U148 ( .A(b[0]), .Z(n127) );
  IV U149 ( .A(b[0]), .Z(n128) );
  IV U150 ( .A(b[0]), .Z(n129) );
  IV U151 ( .A(b[0]), .Z(n130) );
  IV U152 ( .A(b[0]), .Z(n131) );
  IV U153 ( .A(b[0]), .Z(n132) );
  IV U154 ( .A(b[0]), .Z(n133) );
  IV U155 ( .A(b[0]), .Z(n134) );
  IV U156 ( .A(b[0]), .Z(n135) );
  IV U157 ( .A(b[0]), .Z(n136) );
  IV U158 ( .A(b[0]), .Z(n137) );
  IV U159 ( .A(b[0]), .Z(n138) );
  IV U160 ( .A(b[0]), .Z(n139) );
  IV U161 ( .A(b[0]), .Z(n140) );
  IV U162 ( .A(b[0]), .Z(n141) );
  IV U163 ( .A(b[0]), .Z(n142) );
  IV U164 ( .A(b[0]), .Z(n143) );
  IV U165 ( .A(b[0]), .Z(n144) );
  IV U166 ( .A(b[0]), .Z(n145) );
  IV U167 ( .A(b[0]), .Z(n146) );
  IV U168 ( .A(b[0]), .Z(n147) );
  IV U169 ( .A(b[0]), .Z(n148) );
  IV U170 ( .A(b[0]), .Z(n149) );
  IV U171 ( .A(b[0]), .Z(n150) );
  IV U172 ( .A(b[0]), .Z(n151) );
  IV U173 ( .A(b[0]), .Z(n152) );
  IV U174 ( .A(b[0]), .Z(n153) );
  IV U175 ( .A(b[0]), .Z(n154) );
  IV U176 ( .A(b[0]), .Z(n155) );
  IV U177 ( .A(b[0]), .Z(n156) );
  IV U178 ( .A(b[0]), .Z(n157) );
  IV U179 ( .A(b[0]), .Z(n158) );
  IV U180 ( .A(b[0]), .Z(n159) );
  IV U181 ( .A(b[0]), .Z(n160) );
  IV U182 ( .A(b[0]), .Z(n161) );
  IV U183 ( .A(b[7]), .Z(n162) );
  IV U184 ( .A(b[7]), .Z(n163) );
  IV U185 ( .A(b[7]), .Z(n164) );
  IV U186 ( .A(b[7]), .Z(n165) );
  IV U187 ( .A(b[7]), .Z(n166) );
  IV U188 ( .A(b[7]), .Z(n167) );
  IV U189 ( .A(b[7]), .Z(n168) );
  IV U190 ( .A(b[7]), .Z(n169) );
  IV U191 ( .A(b[7]), .Z(n170) );
  IV U192 ( .A(b[7]), .Z(n171) );
  IV U193 ( .A(b[7]), .Z(n172) );
  IV U194 ( .A(b[7]), .Z(n173) );
  IV U195 ( .A(b[7]), .Z(n174) );
  IV U196 ( .A(b[7]), .Z(n175) );
  IV U197 ( .A(b[7]), .Z(n176) );
  IV U198 ( .A(b[7]), .Z(n177) );
  IV U199 ( .A(b[7]), .Z(n178) );
  IV U200 ( .A(b[7]), .Z(n179) );
  IV U201 ( .A(b[7]), .Z(n180) );
  IV U202 ( .A(b[7]), .Z(n181) );
  IV U203 ( .A(b[7]), .Z(n182) );
  IV U204 ( .A(b[7]), .Z(n183) );
  IV U205 ( .A(b[7]), .Z(n184) );
  IV U206 ( .A(b[7]), .Z(n185) );
  IV U207 ( .A(b[7]), .Z(n186) );
  IV U208 ( .A(b[7]), .Z(n187) );
  IV U209 ( .A(b[7]), .Z(n188) );
  IV U210 ( .A(b[7]), .Z(n189) );
  IV U211 ( .A(b[7]), .Z(n190) );
  IV U212 ( .A(b[7]), .Z(n191) );
  IV U213 ( .A(b[7]), .Z(n192) );
  IV U214 ( .A(b[7]), .Z(n193) );
  IV U215 ( .A(b[7]), .Z(n194) );
  IV U216 ( .A(b[7]), .Z(n195) );
  IV U217 ( .A(b[7]), .Z(n196) );
  IV U218 ( .A(b[7]), .Z(n197) );
  IV U219 ( .A(b[7]), .Z(n198) );
  IV U220 ( .A(b[7]), .Z(n199) );
  IV U221 ( .A(b[7]), .Z(n200) );
  IV U222 ( .A(b[7]), .Z(n201) );
  IV U223 ( .A(b[7]), .Z(n202) );
  IV U224 ( .A(b[7]), .Z(n203) );
  IV U225 ( .A(b[7]), .Z(n204) );
  IV U226 ( .A(b[7]), .Z(n205) );
  IV U227 ( .A(b[7]), .Z(n206) );
  IV U228 ( .A(b[7]), .Z(n207) );
  IV U229 ( .A(b[7]), .Z(n208) );
  IV U230 ( .A(b[7]), .Z(n209) );
  IV U231 ( .A(b[7]), .Z(n210) );
  IV U232 ( .A(b[7]), .Z(n211) );
  IV U233 ( .A(b[7]), .Z(n212) );
  IV U234 ( .A(b[7]), .Z(n213) );
  IV U235 ( .A(b[7]), .Z(n214) );
  IV U236 ( .A(b[7]), .Z(n215) );
  IV U237 ( .A(b[7]), .Z(n216) );
  IV U238 ( .A(b[7]), .Z(n217) );
  IV U239 ( .A(b[7]), .Z(n218) );
  IV U240 ( .A(b[7]), .Z(n219) );
  IV U241 ( .A(b[7]), .Z(n220) );
  IV U242 ( .A(b[7]), .Z(n221) );
  IV U243 ( .A(b[7]), .Z(n222) );
  IV U244 ( .A(b[7]), .Z(n223) );
  IV U245 ( .A(b[7]), .Z(n224) );
  IV U246 ( .A(b[7]), .Z(n225) );
  IV U247 ( .A(b[7]), .Z(n226) );
  IV U248 ( .A(b[7]), .Z(n227) );
  IV U249 ( .A(b[7]), .Z(n228) );
  IV U250 ( .A(b[7]), .Z(n229) );
  IV U251 ( .A(b[7]), .Z(n230) );
  IV U252 ( .A(b[7]), .Z(n231) );
  IV U253 ( .A(b[7]), .Z(n232) );
  IV U254 ( .A(b[7]), .Z(n233) );
  IV U255 ( .A(b[7]), .Z(n234) );
  IV U256 ( .A(b[7]), .Z(n235) );
  IV U257 ( .A(b[7]), .Z(n236) );
  IV U258 ( .A(b[7]), .Z(n237) );
  IV U259 ( .A(b[7]), .Z(n238) );
  IV U260 ( .A(b[7]), .Z(n239) );
  IV U261 ( .A(b[7]), .Z(n240) );
  IV U262 ( .A(b[7]), .Z(n241) );
  IV U263 ( .A(b[7]), .Z(n242) );
  IV U264 ( .A(b[7]), .Z(n243) );
  IV U265 ( .A(b[7]), .Z(n244) );
  IV U266 ( .A(b[7]), .Z(n245) );
  IV U267 ( .A(b[7]), .Z(n246) );
  IV U268 ( .A(b[7]), .Z(n247) );
  NAND U269 ( .A(b[0]), .B(a[0]), .Z(n249) );
  XNOR U270 ( .A(n249), .B(sreg[1016]), .Z(c[1016]) );
  NAND U271 ( .A(b[0]), .B(a[1]), .Z(n254) );
  NAND U272 ( .A(b[1]), .B(a[0]), .Z(n248) );
  XOR U273 ( .A(n254), .B(n248), .Z(n257) );
  XNOR U274 ( .A(sreg[1017]), .B(n257), .Z(n259) );
  NANDN U275 ( .A(n249), .B(sreg[1016]), .Z(n258) );
  XOR U276 ( .A(n259), .B(n258), .Z(c[1017]) );
  NAND U277 ( .A(b[0]), .B(a[2]), .Z(n250) );
  XNOR U278 ( .A(b[1]), .B(n250), .Z(n252) );
  NAND U279 ( .A(a[1]), .B(n15), .Z(n251) );
  AND U280 ( .A(n252), .B(n251), .Z(n271) );
  NAND U281 ( .A(a[0]), .B(b[2]), .Z(n253) );
  XNOR U282 ( .A(b[1]), .B(n253), .Z(n256) );
  OR U283 ( .A(n254), .B(a[0]), .Z(n255) );
  AND U284 ( .A(n256), .B(n255), .Z(n272) );
  XNOR U285 ( .A(n271), .B(n272), .Z(n275) );
  NAND U286 ( .A(n257), .B(sreg[1017]), .Z(n261) );
  OR U287 ( .A(n259), .B(n258), .Z(n260) );
  NAND U288 ( .A(n261), .B(n260), .Z(n273) );
  XNOR U289 ( .A(n273), .B(sreg[1018]), .Z(n274) );
  XOR U290 ( .A(n275), .B(n274), .Z(c[1018]) );
  NAND U291 ( .A(b[0]), .B(a[3]), .Z(n262) );
  XNOR U292 ( .A(b[1]), .B(n262), .Z(n264) );
  NAND U293 ( .A(n15), .B(a[2]), .Z(n263) );
  AND U294 ( .A(n264), .B(n263), .Z(n287) );
  XOR U295 ( .A(a[0]), .B(b[3]), .Z(n266) );
  XOR U296 ( .A(b[2]), .B(b[3]), .Z(n265) );
  ANDN U297 ( .B(n265), .A(n42095), .Z(n42093) );
  NAND U298 ( .A(n266), .B(n42093), .Z(n268) );
  IV U299 ( .A(b[3]), .Z(n42134) );
  IV U300 ( .A(a[1]), .Z(n372) );
  XNOR U301 ( .A(n42134), .B(n372), .Z(n292) );
  ANDN U302 ( .B(n42095), .A(n292), .Z(n267) );
  ANDN U303 ( .B(n268), .A(n267), .Z(n288) );
  XOR U304 ( .A(n287), .B(n288), .Z(n283) );
  NAND U305 ( .A(a[0]), .B(n42095), .Z(n270) );
  NAND U306 ( .A(b[1]), .B(b[2]), .Z(n269) );
  NANDN U307 ( .A(n42134), .B(n269), .Z(n42206) );
  ANDN U308 ( .B(n270), .A(n42206), .Z(n284) );
  XNOR U309 ( .A(n283), .B(n284), .Z(n285) );
  NAND U310 ( .A(n272), .B(n271), .Z(n286) );
  XNOR U311 ( .A(n285), .B(n286), .Z(n278) );
  XNOR U312 ( .A(sreg[1019]), .B(n278), .Z(n280) );
  NAND U313 ( .A(n273), .B(sreg[1018]), .Z(n277) );
  OR U314 ( .A(n275), .B(n274), .Z(n276) );
  AND U315 ( .A(n277), .B(n276), .Z(n279) );
  XOR U316 ( .A(n280), .B(n279), .Z(c[1019]) );
  NAND U317 ( .A(sreg[1019]), .B(n278), .Z(n282) );
  OR U318 ( .A(n280), .B(n279), .Z(n281) );
  NAND U319 ( .A(n282), .B(n281), .Z(n319) );
  XNOR U320 ( .A(n319), .B(sreg[1020]), .Z(n321) );
  XOR U321 ( .A(n42134), .B(b[4]), .Z(n308) );
  ANDN U322 ( .B(a[0]), .A(n308), .Z(n315) );
  NAND U323 ( .A(b[0]), .B(a[4]), .Z(n289) );
  XNOR U324 ( .A(b[1]), .B(n289), .Z(n291) );
  NAND U325 ( .A(n15), .B(a[3]), .Z(n290) );
  AND U326 ( .A(n291), .B(n290), .Z(n302) );
  NANDN U327 ( .A(n292), .B(n42093), .Z(n294) );
  XOR U328 ( .A(n42134), .B(a[2]), .Z(n316) );
  NANDN U329 ( .A(n316), .B(n42095), .Z(n293) );
  AND U330 ( .A(n294), .B(n293), .Z(n301) );
  XNOR U331 ( .A(n302), .B(n301), .Z(n303) );
  XNOR U332 ( .A(n315), .B(n303), .Z(n295) );
  XNOR U333 ( .A(n296), .B(n295), .Z(n297) );
  XOR U334 ( .A(n298), .B(n297), .Z(n320) );
  XOR U335 ( .A(n321), .B(n320), .Z(c[1020]) );
  NAND U336 ( .A(n296), .B(n295), .Z(n300) );
  OR U337 ( .A(n298), .B(n297), .Z(n299) );
  NAND U338 ( .A(n300), .B(n299), .Z(n327) );
  NANDN U339 ( .A(n302), .B(n301), .Z(n305) );
  NANDN U340 ( .A(n315), .B(n303), .Z(n304) );
  NAND U341 ( .A(n305), .B(n304), .Z(n325) );
  XOR U342 ( .A(b[5]), .B(a[0]), .Z(n307) );
  XOR U343 ( .A(b[5]), .B(b[3]), .Z(n336) );
  AND U344 ( .A(n336), .B(n308), .Z(n306) );
  NAND U345 ( .A(n307), .B(n306), .Z(n310) );
  IV U346 ( .A(b[5]), .Z(n42197) );
  XNOR U347 ( .A(n42197), .B(n372), .Z(n337) );
  IV U348 ( .A(n308), .Z(n42173) );
  NANDN U349 ( .A(n337), .B(n42173), .Z(n309) );
  NAND U350 ( .A(n310), .B(n309), .Z(n329) );
  NAND U351 ( .A(b[0]), .B(a[5]), .Z(n311) );
  XNOR U352 ( .A(b[1]), .B(n311), .Z(n313) );
  NAND U353 ( .A(n15), .B(a[4]), .Z(n312) );
  NAND U354 ( .A(n313), .B(n312), .Z(n328) );
  XNOR U355 ( .A(n329), .B(n328), .Z(n343) );
  NAND U356 ( .A(b[3]), .B(b[4]), .Z(n314) );
  NANDN U357 ( .A(n42197), .B(n314), .Z(n42250) );
  NOR U358 ( .A(n315), .B(n42250), .Z(n340) );
  NANDN U359 ( .A(n316), .B(n42093), .Z(n318) );
  XOR U360 ( .A(a[3]), .B(b[3]), .Z(n330) );
  NAND U361 ( .A(n42095), .B(n330), .Z(n317) );
  NAND U362 ( .A(n318), .B(n317), .Z(n341) );
  XOR U363 ( .A(n340), .B(n341), .Z(n342) );
  XOR U364 ( .A(n343), .B(n342), .Z(n324) );
  XOR U365 ( .A(n325), .B(n324), .Z(n326) );
  XOR U366 ( .A(n327), .B(n326), .Z(n344) );
  XNOR U367 ( .A(n344), .B(sreg[1021]), .Z(n346) );
  NAND U368 ( .A(n319), .B(sreg[1020]), .Z(n323) );
  OR U369 ( .A(n321), .B(n320), .Z(n322) );
  AND U370 ( .A(n323), .B(n322), .Z(n345) );
  XOR U371 ( .A(n346), .B(n345), .Z(c[1021]) );
  ANDN U372 ( .B(n329), .A(n328), .Z(n358) );
  XOR U373 ( .A(n42134), .B(a[4]), .Z(n366) );
  NANDN U374 ( .A(n366), .B(n42095), .Z(n332) );
  NAND U375 ( .A(n330), .B(n42093), .Z(n331) );
  NAND U376 ( .A(n332), .B(n331), .Z(n363) );
  XNOR U377 ( .A(n42197), .B(b[6]), .Z(n42234) );
  AND U378 ( .A(n42234), .B(a[0]), .Z(n377) );
  NAND U379 ( .A(b[0]), .B(a[6]), .Z(n333) );
  XNOR U380 ( .A(b[1]), .B(n333), .Z(n335) );
  NAND U381 ( .A(n15), .B(a[5]), .Z(n334) );
  AND U382 ( .A(n335), .B(n334), .Z(n361) );
  XOR U383 ( .A(n377), .B(n361), .Z(n362) );
  XNOR U384 ( .A(n363), .B(n362), .Z(n355) );
  ANDN U385 ( .B(n336), .A(n42173), .Z(n42172) );
  NANDN U386 ( .A(n337), .B(n42172), .Z(n339) );
  XOR U387 ( .A(a[2]), .B(b[5]), .Z(n369) );
  NAND U388 ( .A(n42173), .B(n369), .Z(n338) );
  NAND U389 ( .A(n339), .B(n338), .Z(n356) );
  XNOR U390 ( .A(n355), .B(n356), .Z(n357) );
  XOR U391 ( .A(n358), .B(n357), .Z(n349) );
  XOR U392 ( .A(n349), .B(n350), .Z(n352) );
  XOR U393 ( .A(n351), .B(n352), .Z(n383) );
  NAND U394 ( .A(n344), .B(sreg[1021]), .Z(n348) );
  OR U395 ( .A(n346), .B(n345), .Z(n347) );
  NAND U396 ( .A(n348), .B(n347), .Z(n382) );
  XNOR U397 ( .A(n382), .B(sreg[1022]), .Z(n384) );
  XNOR U398 ( .A(n383), .B(n384), .Z(c[1022]) );
  NANDN U399 ( .A(n350), .B(n349), .Z(n354) );
  OR U400 ( .A(n352), .B(n351), .Z(n353) );
  NAND U401 ( .A(n354), .B(n353), .Z(n395) );
  NANDN U402 ( .A(n356), .B(n355), .Z(n360) );
  NANDN U403 ( .A(n358), .B(n357), .Z(n359) );
  NAND U404 ( .A(n360), .B(n359), .Z(n393) );
  NAND U405 ( .A(n377), .B(n361), .Z(n365) );
  NAND U406 ( .A(n363), .B(n362), .Z(n364) );
  NAND U407 ( .A(n365), .B(n364), .Z(n399) );
  NANDN U408 ( .A(n366), .B(n42093), .Z(n368) );
  XOR U409 ( .A(n42134), .B(a[5]), .Z(n412) );
  NANDN U410 ( .A(n412), .B(n42095), .Z(n367) );
  AND U411 ( .A(n368), .B(n367), .Z(n398) );
  XNOR U412 ( .A(n399), .B(n398), .Z(n400) );
  XOR U413 ( .A(n42197), .B(a[3]), .Z(n421) );
  NANDN U414 ( .A(n421), .B(n42173), .Z(n371) );
  NAND U415 ( .A(n42172), .B(n369), .Z(n370) );
  NAND U416 ( .A(n371), .B(n370), .Z(n411) );
  XNOR U417 ( .A(n162), .B(n372), .Z(n415) );
  NANDN U418 ( .A(n415), .B(n42234), .Z(n376) );
  XNOR U419 ( .A(a[0]), .B(n162), .Z(n374) );
  XNOR U420 ( .A(b[5]), .B(n162), .Z(n373) );
  ANDN U421 ( .B(n373), .A(n42234), .Z(n42231) );
  NAND U422 ( .A(n374), .B(n42231), .Z(n375) );
  NAND U423 ( .A(n376), .B(n375), .Z(n410) );
  XNOR U424 ( .A(n411), .B(n410), .Z(n407) );
  ANDN U425 ( .B(b[6]), .A(n42197), .Z(n42273) );
  ANDN U426 ( .B(b[7]), .A(n42273), .Z(n378) );
  ANDN U427 ( .B(n378), .A(n377), .Z(n404) );
  NAND U428 ( .A(b[0]), .B(a[7]), .Z(n379) );
  XNOR U429 ( .A(b[1]), .B(n379), .Z(n381) );
  NAND U430 ( .A(n16), .B(a[6]), .Z(n380) );
  AND U431 ( .A(n381), .B(n380), .Z(n405) );
  XOR U432 ( .A(n404), .B(n405), .Z(n406) );
  XOR U433 ( .A(n407), .B(n406), .Z(n401) );
  XOR U434 ( .A(n400), .B(n401), .Z(n392) );
  XNOR U435 ( .A(n393), .B(n392), .Z(n394) );
  XNOR U436 ( .A(n395), .B(n394), .Z(n387) );
  XNOR U437 ( .A(n387), .B(sreg[1023]), .Z(n389) );
  NAND U438 ( .A(n382), .B(sreg[1022]), .Z(n386) );
  NANDN U439 ( .A(n384), .B(n383), .Z(n385) );
  AND U440 ( .A(n386), .B(n385), .Z(n388) );
  XOR U441 ( .A(n389), .B(n388), .Z(c[1023]) );
  NAND U442 ( .A(n387), .B(sreg[1023]), .Z(n391) );
  OR U443 ( .A(n389), .B(n388), .Z(n390) );
  NAND U444 ( .A(n391), .B(n390), .Z(n460) );
  XNOR U445 ( .A(n460), .B(sreg[1024]), .Z(n462) );
  NAND U446 ( .A(n393), .B(n392), .Z(n397) );
  OR U447 ( .A(n395), .B(n394), .Z(n396) );
  NAND U448 ( .A(n397), .B(n396), .Z(n427) );
  NANDN U449 ( .A(n399), .B(n398), .Z(n403) );
  NAND U450 ( .A(n401), .B(n400), .Z(n402) );
  NAND U451 ( .A(n403), .B(n402), .Z(n425) );
  OR U452 ( .A(n405), .B(n404), .Z(n409) );
  NAND U453 ( .A(n407), .B(n406), .Z(n408) );
  NAND U454 ( .A(n409), .B(n408), .Z(n454) );
  NAND U455 ( .A(n411), .B(n410), .Z(n451) );
  NANDN U456 ( .A(n412), .B(n42093), .Z(n414) );
  XOR U457 ( .A(n42134), .B(a[6]), .Z(n436) );
  NANDN U458 ( .A(n436), .B(n42095), .Z(n413) );
  NAND U459 ( .A(n414), .B(n413), .Z(n449) );
  NANDN U460 ( .A(n415), .B(n42231), .Z(n417) );
  XOR U461 ( .A(n162), .B(a[2]), .Z(n439) );
  NANDN U462 ( .A(n439), .B(n42234), .Z(n416) );
  AND U463 ( .A(n417), .B(n416), .Z(n448) );
  XNOR U464 ( .A(n449), .B(n448), .Z(n450) );
  XNOR U465 ( .A(n451), .B(n450), .Z(n455) );
  XNOR U466 ( .A(n454), .B(n455), .Z(n456) );
  NAND U467 ( .A(b[0]), .B(a[8]), .Z(n418) );
  XNOR U468 ( .A(b[1]), .B(n418), .Z(n420) );
  NAND U469 ( .A(n16), .B(a[7]), .Z(n419) );
  AND U470 ( .A(n420), .B(n419), .Z(n445) );
  AND U471 ( .A(a[0]), .B(b[7]), .Z(n442) );
  NANDN U472 ( .A(n421), .B(n42172), .Z(n423) );
  XOR U473 ( .A(a[4]), .B(b[5]), .Z(n433) );
  NAND U474 ( .A(n42173), .B(n433), .Z(n422) );
  NAND U475 ( .A(n423), .B(n422), .Z(n443) );
  XOR U476 ( .A(n442), .B(n443), .Z(n444) );
  XOR U477 ( .A(n445), .B(n444), .Z(n457) );
  XNOR U478 ( .A(n456), .B(n457), .Z(n424) );
  XOR U479 ( .A(n425), .B(n424), .Z(n426) );
  XOR U480 ( .A(n427), .B(n426), .Z(n461) );
  XOR U481 ( .A(n462), .B(n461), .Z(c[1024]) );
  NAND U482 ( .A(n425), .B(n424), .Z(n429) );
  NAND U483 ( .A(n427), .B(n426), .Z(n428) );
  NAND U484 ( .A(n429), .B(n428), .Z(n468) );
  NAND U485 ( .A(b[0]), .B(a[9]), .Z(n430) );
  XNOR U486 ( .A(b[1]), .B(n430), .Z(n432) );
  NAND U487 ( .A(n16), .B(a[8]), .Z(n431) );
  AND U488 ( .A(n432), .B(n431), .Z(n485) );
  XOR U489 ( .A(a[5]), .B(n42197), .Z(n474) );
  NANDN U490 ( .A(n474), .B(n42173), .Z(n435) );
  NAND U491 ( .A(n42172), .B(n433), .Z(n434) );
  NAND U492 ( .A(n435), .B(n434), .Z(n483) );
  NAND U493 ( .A(b[7]), .B(a[1]), .Z(n484) );
  XNOR U494 ( .A(n483), .B(n484), .Z(n486) );
  XOR U495 ( .A(n485), .B(n486), .Z(n492) );
  NANDN U496 ( .A(n436), .B(n42093), .Z(n438) );
  XOR U497 ( .A(n42134), .B(a[7]), .Z(n477) );
  NANDN U498 ( .A(n477), .B(n42095), .Z(n437) );
  NAND U499 ( .A(n438), .B(n437), .Z(n490) );
  NANDN U500 ( .A(n439), .B(n42231), .Z(n441) );
  XOR U501 ( .A(n162), .B(a[3]), .Z(n480) );
  NANDN U502 ( .A(n480), .B(n42234), .Z(n440) );
  AND U503 ( .A(n441), .B(n440), .Z(n489) );
  XNOR U504 ( .A(n490), .B(n489), .Z(n491) );
  XNOR U505 ( .A(n492), .B(n491), .Z(n495) );
  OR U506 ( .A(n443), .B(n442), .Z(n447) );
  NANDN U507 ( .A(n445), .B(n444), .Z(n446) );
  NAND U508 ( .A(n447), .B(n446), .Z(n496) );
  XOR U509 ( .A(n495), .B(n496), .Z(n497) );
  NANDN U510 ( .A(n449), .B(n448), .Z(n453) );
  NAND U511 ( .A(n451), .B(n450), .Z(n452) );
  NAND U512 ( .A(n453), .B(n452), .Z(n498) );
  XOR U513 ( .A(n497), .B(n498), .Z(n465) );
  NANDN U514 ( .A(n455), .B(n454), .Z(n459) );
  NANDN U515 ( .A(n457), .B(n456), .Z(n458) );
  AND U516 ( .A(n459), .B(n458), .Z(n466) );
  XNOR U517 ( .A(n465), .B(n466), .Z(n467) );
  XNOR U518 ( .A(n468), .B(n467), .Z(n501) );
  XNOR U519 ( .A(n501), .B(sreg[1025]), .Z(n503) );
  NAND U520 ( .A(n460), .B(sreg[1024]), .Z(n464) );
  OR U521 ( .A(n462), .B(n461), .Z(n463) );
  AND U522 ( .A(n464), .B(n463), .Z(n502) );
  XOR U523 ( .A(n503), .B(n502), .Z(c[1025]) );
  NANDN U524 ( .A(n466), .B(n465), .Z(n470) );
  NAND U525 ( .A(n468), .B(n467), .Z(n469) );
  NAND U526 ( .A(n470), .B(n469), .Z(n509) );
  NAND U527 ( .A(b[0]), .B(a[10]), .Z(n471) );
  XNOR U528 ( .A(b[1]), .B(n471), .Z(n473) );
  NAND U529 ( .A(n16), .B(a[9]), .Z(n472) );
  AND U530 ( .A(n473), .B(n472), .Z(n526) );
  XOR U531 ( .A(a[6]), .B(n42197), .Z(n515) );
  NANDN U532 ( .A(n515), .B(n42173), .Z(n476) );
  NANDN U533 ( .A(n474), .B(n42172), .Z(n475) );
  NAND U534 ( .A(n476), .B(n475), .Z(n524) );
  NAND U535 ( .A(b[7]), .B(a[2]), .Z(n525) );
  XNOR U536 ( .A(n524), .B(n525), .Z(n527) );
  XOR U537 ( .A(n526), .B(n527), .Z(n533) );
  NANDN U538 ( .A(n477), .B(n42093), .Z(n479) );
  XOR U539 ( .A(n42134), .B(a[8]), .Z(n518) );
  NANDN U540 ( .A(n518), .B(n42095), .Z(n478) );
  NAND U541 ( .A(n479), .B(n478), .Z(n531) );
  NANDN U542 ( .A(n480), .B(n42231), .Z(n482) );
  XOR U543 ( .A(n162), .B(a[4]), .Z(n521) );
  NANDN U544 ( .A(n521), .B(n42234), .Z(n481) );
  AND U545 ( .A(n482), .B(n481), .Z(n530) );
  XNOR U546 ( .A(n531), .B(n530), .Z(n532) );
  XNOR U547 ( .A(n533), .B(n532), .Z(n537) );
  NANDN U548 ( .A(n484), .B(n483), .Z(n488) );
  NAND U549 ( .A(n486), .B(n485), .Z(n487) );
  AND U550 ( .A(n488), .B(n487), .Z(n536) );
  XOR U551 ( .A(n537), .B(n536), .Z(n538) );
  NANDN U552 ( .A(n490), .B(n489), .Z(n494) );
  NANDN U553 ( .A(n492), .B(n491), .Z(n493) );
  NAND U554 ( .A(n494), .B(n493), .Z(n539) );
  XOR U555 ( .A(n538), .B(n539), .Z(n506) );
  OR U556 ( .A(n496), .B(n495), .Z(n500) );
  NANDN U557 ( .A(n498), .B(n497), .Z(n499) );
  NAND U558 ( .A(n500), .B(n499), .Z(n507) );
  XNOR U559 ( .A(n506), .B(n507), .Z(n508) );
  XNOR U560 ( .A(n509), .B(n508), .Z(n542) );
  XNOR U561 ( .A(n542), .B(sreg[1026]), .Z(n544) );
  NAND U562 ( .A(n501), .B(sreg[1025]), .Z(n505) );
  OR U563 ( .A(n503), .B(n502), .Z(n504) );
  AND U564 ( .A(n505), .B(n504), .Z(n543) );
  XOR U565 ( .A(n544), .B(n543), .Z(c[1026]) );
  NANDN U566 ( .A(n507), .B(n506), .Z(n511) );
  NAND U567 ( .A(n509), .B(n508), .Z(n510) );
  NAND U568 ( .A(n511), .B(n510), .Z(n550) );
  NAND U569 ( .A(b[0]), .B(a[11]), .Z(n512) );
  XNOR U570 ( .A(b[1]), .B(n512), .Z(n514) );
  NAND U571 ( .A(n16), .B(a[10]), .Z(n513) );
  AND U572 ( .A(n514), .B(n513), .Z(n567) );
  XOR U573 ( .A(a[7]), .B(n42197), .Z(n556) );
  NANDN U574 ( .A(n556), .B(n42173), .Z(n517) );
  NANDN U575 ( .A(n515), .B(n42172), .Z(n516) );
  NAND U576 ( .A(n517), .B(n516), .Z(n565) );
  NAND U577 ( .A(b[7]), .B(a[3]), .Z(n566) );
  XNOR U578 ( .A(n565), .B(n566), .Z(n568) );
  XOR U579 ( .A(n567), .B(n568), .Z(n574) );
  NANDN U580 ( .A(n518), .B(n42093), .Z(n520) );
  XOR U581 ( .A(n42134), .B(a[9]), .Z(n559) );
  NANDN U582 ( .A(n559), .B(n42095), .Z(n519) );
  NAND U583 ( .A(n520), .B(n519), .Z(n572) );
  NANDN U584 ( .A(n521), .B(n42231), .Z(n523) );
  XOR U585 ( .A(n162), .B(a[5]), .Z(n562) );
  NANDN U586 ( .A(n562), .B(n42234), .Z(n522) );
  AND U587 ( .A(n523), .B(n522), .Z(n571) );
  XNOR U588 ( .A(n572), .B(n571), .Z(n573) );
  XNOR U589 ( .A(n574), .B(n573), .Z(n578) );
  NANDN U590 ( .A(n525), .B(n524), .Z(n529) );
  NAND U591 ( .A(n527), .B(n526), .Z(n528) );
  AND U592 ( .A(n529), .B(n528), .Z(n577) );
  XOR U593 ( .A(n578), .B(n577), .Z(n579) );
  NANDN U594 ( .A(n531), .B(n530), .Z(n535) );
  NANDN U595 ( .A(n533), .B(n532), .Z(n534) );
  NAND U596 ( .A(n535), .B(n534), .Z(n580) );
  XOR U597 ( .A(n579), .B(n580), .Z(n547) );
  OR U598 ( .A(n537), .B(n536), .Z(n541) );
  NANDN U599 ( .A(n539), .B(n538), .Z(n540) );
  NAND U600 ( .A(n541), .B(n540), .Z(n548) );
  XNOR U601 ( .A(n547), .B(n548), .Z(n549) );
  XNOR U602 ( .A(n550), .B(n549), .Z(n583) );
  XNOR U603 ( .A(n583), .B(sreg[1027]), .Z(n585) );
  NAND U604 ( .A(n542), .B(sreg[1026]), .Z(n546) );
  OR U605 ( .A(n544), .B(n543), .Z(n545) );
  AND U606 ( .A(n546), .B(n545), .Z(n584) );
  XOR U607 ( .A(n585), .B(n584), .Z(c[1027]) );
  NANDN U608 ( .A(n548), .B(n547), .Z(n552) );
  NAND U609 ( .A(n550), .B(n549), .Z(n551) );
  NAND U610 ( .A(n552), .B(n551), .Z(n591) );
  NAND U611 ( .A(b[0]), .B(a[12]), .Z(n553) );
  XNOR U612 ( .A(b[1]), .B(n553), .Z(n555) );
  NAND U613 ( .A(n16), .B(a[11]), .Z(n554) );
  AND U614 ( .A(n555), .B(n554), .Z(n608) );
  XOR U615 ( .A(a[8]), .B(n42197), .Z(n597) );
  NANDN U616 ( .A(n597), .B(n42173), .Z(n558) );
  NANDN U617 ( .A(n556), .B(n42172), .Z(n557) );
  NAND U618 ( .A(n558), .B(n557), .Z(n606) );
  NAND U619 ( .A(b[7]), .B(a[4]), .Z(n607) );
  XNOR U620 ( .A(n606), .B(n607), .Z(n609) );
  XOR U621 ( .A(n608), .B(n609), .Z(n615) );
  NANDN U622 ( .A(n559), .B(n42093), .Z(n561) );
  XOR U623 ( .A(n42134), .B(a[10]), .Z(n600) );
  NANDN U624 ( .A(n600), .B(n42095), .Z(n560) );
  NAND U625 ( .A(n561), .B(n560), .Z(n613) );
  NANDN U626 ( .A(n562), .B(n42231), .Z(n564) );
  XOR U627 ( .A(n162), .B(a[6]), .Z(n603) );
  NANDN U628 ( .A(n603), .B(n42234), .Z(n563) );
  AND U629 ( .A(n564), .B(n563), .Z(n612) );
  XNOR U630 ( .A(n613), .B(n612), .Z(n614) );
  XNOR U631 ( .A(n615), .B(n614), .Z(n619) );
  NANDN U632 ( .A(n566), .B(n565), .Z(n570) );
  NAND U633 ( .A(n568), .B(n567), .Z(n569) );
  AND U634 ( .A(n570), .B(n569), .Z(n618) );
  XOR U635 ( .A(n619), .B(n618), .Z(n620) );
  NANDN U636 ( .A(n572), .B(n571), .Z(n576) );
  NANDN U637 ( .A(n574), .B(n573), .Z(n575) );
  NAND U638 ( .A(n576), .B(n575), .Z(n621) );
  XOR U639 ( .A(n620), .B(n621), .Z(n588) );
  OR U640 ( .A(n578), .B(n577), .Z(n582) );
  NANDN U641 ( .A(n580), .B(n579), .Z(n581) );
  NAND U642 ( .A(n582), .B(n581), .Z(n589) );
  XNOR U643 ( .A(n588), .B(n589), .Z(n590) );
  XNOR U644 ( .A(n591), .B(n590), .Z(n624) );
  XNOR U645 ( .A(n624), .B(sreg[1028]), .Z(n626) );
  NAND U646 ( .A(n583), .B(sreg[1027]), .Z(n587) );
  OR U647 ( .A(n585), .B(n584), .Z(n586) );
  AND U648 ( .A(n587), .B(n586), .Z(n625) );
  XOR U649 ( .A(n626), .B(n625), .Z(c[1028]) );
  NANDN U650 ( .A(n589), .B(n588), .Z(n593) );
  NAND U651 ( .A(n591), .B(n590), .Z(n592) );
  NAND U652 ( .A(n593), .B(n592), .Z(n632) );
  NAND U653 ( .A(b[0]), .B(a[13]), .Z(n594) );
  XNOR U654 ( .A(b[1]), .B(n594), .Z(n596) );
  NAND U655 ( .A(n16), .B(a[12]), .Z(n595) );
  AND U656 ( .A(n596), .B(n595), .Z(n649) );
  XOR U657 ( .A(a[9]), .B(n42197), .Z(n638) );
  NANDN U658 ( .A(n638), .B(n42173), .Z(n599) );
  NANDN U659 ( .A(n597), .B(n42172), .Z(n598) );
  NAND U660 ( .A(n599), .B(n598), .Z(n647) );
  NAND U661 ( .A(b[7]), .B(a[5]), .Z(n648) );
  XNOR U662 ( .A(n647), .B(n648), .Z(n650) );
  XOR U663 ( .A(n649), .B(n650), .Z(n656) );
  NANDN U664 ( .A(n600), .B(n42093), .Z(n602) );
  XOR U665 ( .A(n42134), .B(a[11]), .Z(n641) );
  NANDN U666 ( .A(n641), .B(n42095), .Z(n601) );
  NAND U667 ( .A(n602), .B(n601), .Z(n654) );
  NANDN U668 ( .A(n603), .B(n42231), .Z(n605) );
  XOR U669 ( .A(n162), .B(a[7]), .Z(n644) );
  NANDN U670 ( .A(n644), .B(n42234), .Z(n604) );
  AND U671 ( .A(n605), .B(n604), .Z(n653) );
  XNOR U672 ( .A(n654), .B(n653), .Z(n655) );
  XNOR U673 ( .A(n656), .B(n655), .Z(n660) );
  NANDN U674 ( .A(n607), .B(n606), .Z(n611) );
  NAND U675 ( .A(n609), .B(n608), .Z(n610) );
  AND U676 ( .A(n611), .B(n610), .Z(n659) );
  XOR U677 ( .A(n660), .B(n659), .Z(n661) );
  NANDN U678 ( .A(n613), .B(n612), .Z(n617) );
  NANDN U679 ( .A(n615), .B(n614), .Z(n616) );
  NAND U680 ( .A(n617), .B(n616), .Z(n662) );
  XOR U681 ( .A(n661), .B(n662), .Z(n629) );
  OR U682 ( .A(n619), .B(n618), .Z(n623) );
  NANDN U683 ( .A(n621), .B(n620), .Z(n622) );
  NAND U684 ( .A(n623), .B(n622), .Z(n630) );
  XNOR U685 ( .A(n629), .B(n630), .Z(n631) );
  XNOR U686 ( .A(n632), .B(n631), .Z(n665) );
  XNOR U687 ( .A(n665), .B(sreg[1029]), .Z(n667) );
  NAND U688 ( .A(n624), .B(sreg[1028]), .Z(n628) );
  OR U689 ( .A(n626), .B(n625), .Z(n627) );
  AND U690 ( .A(n628), .B(n627), .Z(n666) );
  XOR U691 ( .A(n667), .B(n666), .Z(c[1029]) );
  NANDN U692 ( .A(n630), .B(n629), .Z(n634) );
  NAND U693 ( .A(n632), .B(n631), .Z(n633) );
  NAND U694 ( .A(n634), .B(n633), .Z(n673) );
  NAND U695 ( .A(b[0]), .B(a[14]), .Z(n635) );
  XNOR U696 ( .A(b[1]), .B(n635), .Z(n637) );
  NAND U697 ( .A(n17), .B(a[13]), .Z(n636) );
  AND U698 ( .A(n637), .B(n636), .Z(n690) );
  XOR U699 ( .A(a[10]), .B(n42197), .Z(n679) );
  NANDN U700 ( .A(n679), .B(n42173), .Z(n640) );
  NANDN U701 ( .A(n638), .B(n42172), .Z(n639) );
  NAND U702 ( .A(n640), .B(n639), .Z(n688) );
  NAND U703 ( .A(b[7]), .B(a[6]), .Z(n689) );
  XNOR U704 ( .A(n688), .B(n689), .Z(n691) );
  XOR U705 ( .A(n690), .B(n691), .Z(n697) );
  NANDN U706 ( .A(n641), .B(n42093), .Z(n643) );
  XOR U707 ( .A(n42134), .B(a[12]), .Z(n682) );
  NANDN U708 ( .A(n682), .B(n42095), .Z(n642) );
  NAND U709 ( .A(n643), .B(n642), .Z(n695) );
  NANDN U710 ( .A(n644), .B(n42231), .Z(n646) );
  XOR U711 ( .A(n162), .B(a[8]), .Z(n685) );
  NANDN U712 ( .A(n685), .B(n42234), .Z(n645) );
  AND U713 ( .A(n646), .B(n645), .Z(n694) );
  XNOR U714 ( .A(n695), .B(n694), .Z(n696) );
  XNOR U715 ( .A(n697), .B(n696), .Z(n701) );
  NANDN U716 ( .A(n648), .B(n647), .Z(n652) );
  NAND U717 ( .A(n650), .B(n649), .Z(n651) );
  AND U718 ( .A(n652), .B(n651), .Z(n700) );
  XOR U719 ( .A(n701), .B(n700), .Z(n702) );
  NANDN U720 ( .A(n654), .B(n653), .Z(n658) );
  NANDN U721 ( .A(n656), .B(n655), .Z(n657) );
  NAND U722 ( .A(n658), .B(n657), .Z(n703) );
  XOR U723 ( .A(n702), .B(n703), .Z(n670) );
  OR U724 ( .A(n660), .B(n659), .Z(n664) );
  NANDN U725 ( .A(n662), .B(n661), .Z(n663) );
  NAND U726 ( .A(n664), .B(n663), .Z(n671) );
  XNOR U727 ( .A(n670), .B(n671), .Z(n672) );
  XNOR U728 ( .A(n673), .B(n672), .Z(n706) );
  XNOR U729 ( .A(n706), .B(sreg[1030]), .Z(n708) );
  NAND U730 ( .A(n665), .B(sreg[1029]), .Z(n669) );
  OR U731 ( .A(n667), .B(n666), .Z(n668) );
  AND U732 ( .A(n669), .B(n668), .Z(n707) );
  XOR U733 ( .A(n708), .B(n707), .Z(c[1030]) );
  NANDN U734 ( .A(n671), .B(n670), .Z(n675) );
  NAND U735 ( .A(n673), .B(n672), .Z(n674) );
  NAND U736 ( .A(n675), .B(n674), .Z(n714) );
  NAND U737 ( .A(b[0]), .B(a[15]), .Z(n676) );
  XNOR U738 ( .A(b[1]), .B(n676), .Z(n678) );
  NAND U739 ( .A(n17), .B(a[14]), .Z(n677) );
  AND U740 ( .A(n678), .B(n677), .Z(n731) );
  XOR U741 ( .A(a[11]), .B(n42197), .Z(n720) );
  NANDN U742 ( .A(n720), .B(n42173), .Z(n681) );
  NANDN U743 ( .A(n679), .B(n42172), .Z(n680) );
  NAND U744 ( .A(n681), .B(n680), .Z(n729) );
  NAND U745 ( .A(b[7]), .B(a[7]), .Z(n730) );
  XNOR U746 ( .A(n729), .B(n730), .Z(n732) );
  XOR U747 ( .A(n731), .B(n732), .Z(n738) );
  NANDN U748 ( .A(n682), .B(n42093), .Z(n684) );
  XOR U749 ( .A(n42134), .B(a[13]), .Z(n723) );
  NANDN U750 ( .A(n723), .B(n42095), .Z(n683) );
  NAND U751 ( .A(n684), .B(n683), .Z(n736) );
  NANDN U752 ( .A(n685), .B(n42231), .Z(n687) );
  XOR U753 ( .A(n162), .B(a[9]), .Z(n726) );
  NANDN U754 ( .A(n726), .B(n42234), .Z(n686) );
  AND U755 ( .A(n687), .B(n686), .Z(n735) );
  XNOR U756 ( .A(n736), .B(n735), .Z(n737) );
  XNOR U757 ( .A(n738), .B(n737), .Z(n742) );
  NANDN U758 ( .A(n689), .B(n688), .Z(n693) );
  NAND U759 ( .A(n691), .B(n690), .Z(n692) );
  AND U760 ( .A(n693), .B(n692), .Z(n741) );
  XOR U761 ( .A(n742), .B(n741), .Z(n743) );
  NANDN U762 ( .A(n695), .B(n694), .Z(n699) );
  NANDN U763 ( .A(n697), .B(n696), .Z(n698) );
  NAND U764 ( .A(n699), .B(n698), .Z(n744) );
  XOR U765 ( .A(n743), .B(n744), .Z(n711) );
  OR U766 ( .A(n701), .B(n700), .Z(n705) );
  NANDN U767 ( .A(n703), .B(n702), .Z(n704) );
  NAND U768 ( .A(n705), .B(n704), .Z(n712) );
  XNOR U769 ( .A(n711), .B(n712), .Z(n713) );
  XNOR U770 ( .A(n714), .B(n713), .Z(n747) );
  XNOR U771 ( .A(n747), .B(sreg[1031]), .Z(n749) );
  NAND U772 ( .A(n706), .B(sreg[1030]), .Z(n710) );
  OR U773 ( .A(n708), .B(n707), .Z(n709) );
  AND U774 ( .A(n710), .B(n709), .Z(n748) );
  XOR U775 ( .A(n749), .B(n748), .Z(c[1031]) );
  NANDN U776 ( .A(n712), .B(n711), .Z(n716) );
  NAND U777 ( .A(n714), .B(n713), .Z(n715) );
  NAND U778 ( .A(n716), .B(n715), .Z(n755) );
  NAND U779 ( .A(b[0]), .B(a[16]), .Z(n717) );
  XNOR U780 ( .A(b[1]), .B(n717), .Z(n719) );
  NAND U781 ( .A(n17), .B(a[15]), .Z(n718) );
  AND U782 ( .A(n719), .B(n718), .Z(n772) );
  XOR U783 ( .A(a[12]), .B(n42197), .Z(n761) );
  NANDN U784 ( .A(n761), .B(n42173), .Z(n722) );
  NANDN U785 ( .A(n720), .B(n42172), .Z(n721) );
  NAND U786 ( .A(n722), .B(n721), .Z(n770) );
  NAND U787 ( .A(b[7]), .B(a[8]), .Z(n771) );
  XNOR U788 ( .A(n770), .B(n771), .Z(n773) );
  XOR U789 ( .A(n772), .B(n773), .Z(n779) );
  NANDN U790 ( .A(n723), .B(n42093), .Z(n725) );
  XOR U791 ( .A(n42134), .B(a[14]), .Z(n764) );
  NANDN U792 ( .A(n764), .B(n42095), .Z(n724) );
  NAND U793 ( .A(n725), .B(n724), .Z(n777) );
  NANDN U794 ( .A(n726), .B(n42231), .Z(n728) );
  XOR U795 ( .A(n162), .B(a[10]), .Z(n767) );
  NANDN U796 ( .A(n767), .B(n42234), .Z(n727) );
  AND U797 ( .A(n728), .B(n727), .Z(n776) );
  XNOR U798 ( .A(n777), .B(n776), .Z(n778) );
  XNOR U799 ( .A(n779), .B(n778), .Z(n783) );
  NANDN U800 ( .A(n730), .B(n729), .Z(n734) );
  NAND U801 ( .A(n732), .B(n731), .Z(n733) );
  AND U802 ( .A(n734), .B(n733), .Z(n782) );
  XOR U803 ( .A(n783), .B(n782), .Z(n784) );
  NANDN U804 ( .A(n736), .B(n735), .Z(n740) );
  NANDN U805 ( .A(n738), .B(n737), .Z(n739) );
  NAND U806 ( .A(n740), .B(n739), .Z(n785) );
  XOR U807 ( .A(n784), .B(n785), .Z(n752) );
  OR U808 ( .A(n742), .B(n741), .Z(n746) );
  NANDN U809 ( .A(n744), .B(n743), .Z(n745) );
  NAND U810 ( .A(n746), .B(n745), .Z(n753) );
  XNOR U811 ( .A(n752), .B(n753), .Z(n754) );
  XNOR U812 ( .A(n755), .B(n754), .Z(n788) );
  XNOR U813 ( .A(n788), .B(sreg[1032]), .Z(n790) );
  NAND U814 ( .A(n747), .B(sreg[1031]), .Z(n751) );
  OR U815 ( .A(n749), .B(n748), .Z(n750) );
  AND U816 ( .A(n751), .B(n750), .Z(n789) );
  XOR U817 ( .A(n790), .B(n789), .Z(c[1032]) );
  NANDN U818 ( .A(n753), .B(n752), .Z(n757) );
  NAND U819 ( .A(n755), .B(n754), .Z(n756) );
  NAND U820 ( .A(n757), .B(n756), .Z(n796) );
  NAND U821 ( .A(b[0]), .B(a[17]), .Z(n758) );
  XNOR U822 ( .A(b[1]), .B(n758), .Z(n760) );
  NAND U823 ( .A(n17), .B(a[16]), .Z(n759) );
  AND U824 ( .A(n760), .B(n759), .Z(n813) );
  XOR U825 ( .A(a[13]), .B(n42197), .Z(n802) );
  NANDN U826 ( .A(n802), .B(n42173), .Z(n763) );
  NANDN U827 ( .A(n761), .B(n42172), .Z(n762) );
  NAND U828 ( .A(n763), .B(n762), .Z(n811) );
  NAND U829 ( .A(b[7]), .B(a[9]), .Z(n812) );
  XNOR U830 ( .A(n811), .B(n812), .Z(n814) );
  XOR U831 ( .A(n813), .B(n814), .Z(n820) );
  NANDN U832 ( .A(n764), .B(n42093), .Z(n766) );
  XOR U833 ( .A(n42134), .B(a[15]), .Z(n805) );
  NANDN U834 ( .A(n805), .B(n42095), .Z(n765) );
  NAND U835 ( .A(n766), .B(n765), .Z(n818) );
  NANDN U836 ( .A(n767), .B(n42231), .Z(n769) );
  XOR U837 ( .A(n163), .B(a[11]), .Z(n808) );
  NANDN U838 ( .A(n808), .B(n42234), .Z(n768) );
  AND U839 ( .A(n769), .B(n768), .Z(n817) );
  XNOR U840 ( .A(n818), .B(n817), .Z(n819) );
  XNOR U841 ( .A(n820), .B(n819), .Z(n824) );
  NANDN U842 ( .A(n771), .B(n770), .Z(n775) );
  NAND U843 ( .A(n773), .B(n772), .Z(n774) );
  AND U844 ( .A(n775), .B(n774), .Z(n823) );
  XOR U845 ( .A(n824), .B(n823), .Z(n825) );
  NANDN U846 ( .A(n777), .B(n776), .Z(n781) );
  NANDN U847 ( .A(n779), .B(n778), .Z(n780) );
  NAND U848 ( .A(n781), .B(n780), .Z(n826) );
  XOR U849 ( .A(n825), .B(n826), .Z(n793) );
  OR U850 ( .A(n783), .B(n782), .Z(n787) );
  NANDN U851 ( .A(n785), .B(n784), .Z(n786) );
  NAND U852 ( .A(n787), .B(n786), .Z(n794) );
  XNOR U853 ( .A(n793), .B(n794), .Z(n795) );
  XNOR U854 ( .A(n796), .B(n795), .Z(n829) );
  XNOR U855 ( .A(n829), .B(sreg[1033]), .Z(n831) );
  NAND U856 ( .A(n788), .B(sreg[1032]), .Z(n792) );
  OR U857 ( .A(n790), .B(n789), .Z(n791) );
  AND U858 ( .A(n792), .B(n791), .Z(n830) );
  XOR U859 ( .A(n831), .B(n830), .Z(c[1033]) );
  NANDN U860 ( .A(n794), .B(n793), .Z(n798) );
  NAND U861 ( .A(n796), .B(n795), .Z(n797) );
  NAND U862 ( .A(n798), .B(n797), .Z(n837) );
  NAND U863 ( .A(b[0]), .B(a[18]), .Z(n799) );
  XNOR U864 ( .A(b[1]), .B(n799), .Z(n801) );
  NAND U865 ( .A(n17), .B(a[17]), .Z(n800) );
  AND U866 ( .A(n801), .B(n800), .Z(n854) );
  XOR U867 ( .A(a[14]), .B(n42197), .Z(n843) );
  NANDN U868 ( .A(n843), .B(n42173), .Z(n804) );
  NANDN U869 ( .A(n802), .B(n42172), .Z(n803) );
  NAND U870 ( .A(n804), .B(n803), .Z(n852) );
  NAND U871 ( .A(b[7]), .B(a[10]), .Z(n853) );
  XNOR U872 ( .A(n852), .B(n853), .Z(n855) );
  XOR U873 ( .A(n854), .B(n855), .Z(n861) );
  NANDN U874 ( .A(n805), .B(n42093), .Z(n807) );
  XOR U875 ( .A(n42134), .B(a[16]), .Z(n846) );
  NANDN U876 ( .A(n846), .B(n42095), .Z(n806) );
  NAND U877 ( .A(n807), .B(n806), .Z(n859) );
  NANDN U878 ( .A(n808), .B(n42231), .Z(n810) );
  XOR U879 ( .A(n163), .B(a[12]), .Z(n849) );
  NANDN U880 ( .A(n849), .B(n42234), .Z(n809) );
  AND U881 ( .A(n810), .B(n809), .Z(n858) );
  XNOR U882 ( .A(n859), .B(n858), .Z(n860) );
  XNOR U883 ( .A(n861), .B(n860), .Z(n865) );
  NANDN U884 ( .A(n812), .B(n811), .Z(n816) );
  NAND U885 ( .A(n814), .B(n813), .Z(n815) );
  AND U886 ( .A(n816), .B(n815), .Z(n864) );
  XOR U887 ( .A(n865), .B(n864), .Z(n866) );
  NANDN U888 ( .A(n818), .B(n817), .Z(n822) );
  NANDN U889 ( .A(n820), .B(n819), .Z(n821) );
  NAND U890 ( .A(n822), .B(n821), .Z(n867) );
  XOR U891 ( .A(n866), .B(n867), .Z(n834) );
  OR U892 ( .A(n824), .B(n823), .Z(n828) );
  NANDN U893 ( .A(n826), .B(n825), .Z(n827) );
  NAND U894 ( .A(n828), .B(n827), .Z(n835) );
  XNOR U895 ( .A(n834), .B(n835), .Z(n836) );
  XNOR U896 ( .A(n837), .B(n836), .Z(n870) );
  XNOR U897 ( .A(n870), .B(sreg[1034]), .Z(n872) );
  NAND U898 ( .A(n829), .B(sreg[1033]), .Z(n833) );
  OR U899 ( .A(n831), .B(n830), .Z(n832) );
  AND U900 ( .A(n833), .B(n832), .Z(n871) );
  XOR U901 ( .A(n872), .B(n871), .Z(c[1034]) );
  NANDN U902 ( .A(n835), .B(n834), .Z(n839) );
  NAND U903 ( .A(n837), .B(n836), .Z(n838) );
  NAND U904 ( .A(n839), .B(n838), .Z(n878) );
  NAND U905 ( .A(b[0]), .B(a[19]), .Z(n840) );
  XNOR U906 ( .A(b[1]), .B(n840), .Z(n842) );
  NAND U907 ( .A(n17), .B(a[18]), .Z(n841) );
  AND U908 ( .A(n842), .B(n841), .Z(n895) );
  XOR U909 ( .A(a[15]), .B(n42197), .Z(n884) );
  NANDN U910 ( .A(n884), .B(n42173), .Z(n845) );
  NANDN U911 ( .A(n843), .B(n42172), .Z(n844) );
  NAND U912 ( .A(n845), .B(n844), .Z(n893) );
  NAND U913 ( .A(b[7]), .B(a[11]), .Z(n894) );
  XNOR U914 ( .A(n893), .B(n894), .Z(n896) );
  XOR U915 ( .A(n895), .B(n896), .Z(n902) );
  NANDN U916 ( .A(n846), .B(n42093), .Z(n848) );
  XOR U917 ( .A(n42134), .B(a[17]), .Z(n887) );
  NANDN U918 ( .A(n887), .B(n42095), .Z(n847) );
  NAND U919 ( .A(n848), .B(n847), .Z(n900) );
  NANDN U920 ( .A(n849), .B(n42231), .Z(n851) );
  XOR U921 ( .A(n163), .B(a[13]), .Z(n890) );
  NANDN U922 ( .A(n890), .B(n42234), .Z(n850) );
  AND U923 ( .A(n851), .B(n850), .Z(n899) );
  XNOR U924 ( .A(n900), .B(n899), .Z(n901) );
  XNOR U925 ( .A(n902), .B(n901), .Z(n906) );
  NANDN U926 ( .A(n853), .B(n852), .Z(n857) );
  NAND U927 ( .A(n855), .B(n854), .Z(n856) );
  AND U928 ( .A(n857), .B(n856), .Z(n905) );
  XOR U929 ( .A(n906), .B(n905), .Z(n907) );
  NANDN U930 ( .A(n859), .B(n858), .Z(n863) );
  NANDN U931 ( .A(n861), .B(n860), .Z(n862) );
  NAND U932 ( .A(n863), .B(n862), .Z(n908) );
  XOR U933 ( .A(n907), .B(n908), .Z(n875) );
  OR U934 ( .A(n865), .B(n864), .Z(n869) );
  NANDN U935 ( .A(n867), .B(n866), .Z(n868) );
  NAND U936 ( .A(n869), .B(n868), .Z(n876) );
  XNOR U937 ( .A(n875), .B(n876), .Z(n877) );
  XNOR U938 ( .A(n878), .B(n877), .Z(n911) );
  XNOR U939 ( .A(n911), .B(sreg[1035]), .Z(n913) );
  NAND U940 ( .A(n870), .B(sreg[1034]), .Z(n874) );
  OR U941 ( .A(n872), .B(n871), .Z(n873) );
  AND U942 ( .A(n874), .B(n873), .Z(n912) );
  XOR U943 ( .A(n913), .B(n912), .Z(c[1035]) );
  NANDN U944 ( .A(n876), .B(n875), .Z(n880) );
  NAND U945 ( .A(n878), .B(n877), .Z(n879) );
  NAND U946 ( .A(n880), .B(n879), .Z(n919) );
  NAND U947 ( .A(b[0]), .B(a[20]), .Z(n881) );
  XNOR U948 ( .A(b[1]), .B(n881), .Z(n883) );
  NAND U949 ( .A(n17), .B(a[19]), .Z(n882) );
  AND U950 ( .A(n883), .B(n882), .Z(n936) );
  XOR U951 ( .A(a[16]), .B(n42197), .Z(n925) );
  NANDN U952 ( .A(n925), .B(n42173), .Z(n886) );
  NANDN U953 ( .A(n884), .B(n42172), .Z(n885) );
  NAND U954 ( .A(n886), .B(n885), .Z(n934) );
  NAND U955 ( .A(b[7]), .B(a[12]), .Z(n935) );
  XNOR U956 ( .A(n934), .B(n935), .Z(n937) );
  XOR U957 ( .A(n936), .B(n937), .Z(n943) );
  NANDN U958 ( .A(n887), .B(n42093), .Z(n889) );
  XOR U959 ( .A(n42134), .B(a[18]), .Z(n928) );
  NANDN U960 ( .A(n928), .B(n42095), .Z(n888) );
  NAND U961 ( .A(n889), .B(n888), .Z(n941) );
  NANDN U962 ( .A(n890), .B(n42231), .Z(n892) );
  XOR U963 ( .A(n163), .B(a[14]), .Z(n931) );
  NANDN U964 ( .A(n931), .B(n42234), .Z(n891) );
  AND U965 ( .A(n892), .B(n891), .Z(n940) );
  XNOR U966 ( .A(n941), .B(n940), .Z(n942) );
  XNOR U967 ( .A(n943), .B(n942), .Z(n947) );
  NANDN U968 ( .A(n894), .B(n893), .Z(n898) );
  NAND U969 ( .A(n896), .B(n895), .Z(n897) );
  AND U970 ( .A(n898), .B(n897), .Z(n946) );
  XOR U971 ( .A(n947), .B(n946), .Z(n948) );
  NANDN U972 ( .A(n900), .B(n899), .Z(n904) );
  NANDN U973 ( .A(n902), .B(n901), .Z(n903) );
  NAND U974 ( .A(n904), .B(n903), .Z(n949) );
  XOR U975 ( .A(n948), .B(n949), .Z(n916) );
  OR U976 ( .A(n906), .B(n905), .Z(n910) );
  NANDN U977 ( .A(n908), .B(n907), .Z(n909) );
  NAND U978 ( .A(n910), .B(n909), .Z(n917) );
  XNOR U979 ( .A(n916), .B(n917), .Z(n918) );
  XNOR U980 ( .A(n919), .B(n918), .Z(n952) );
  XNOR U981 ( .A(n952), .B(sreg[1036]), .Z(n954) );
  NAND U982 ( .A(n911), .B(sreg[1035]), .Z(n915) );
  OR U983 ( .A(n913), .B(n912), .Z(n914) );
  AND U984 ( .A(n915), .B(n914), .Z(n953) );
  XOR U985 ( .A(n954), .B(n953), .Z(c[1036]) );
  NANDN U986 ( .A(n917), .B(n916), .Z(n921) );
  NAND U987 ( .A(n919), .B(n918), .Z(n920) );
  NAND U988 ( .A(n921), .B(n920), .Z(n960) );
  NAND U989 ( .A(b[0]), .B(a[21]), .Z(n922) );
  XNOR U990 ( .A(b[1]), .B(n922), .Z(n924) );
  NAND U991 ( .A(n18), .B(a[20]), .Z(n923) );
  AND U992 ( .A(n924), .B(n923), .Z(n977) );
  XOR U993 ( .A(a[17]), .B(n42197), .Z(n966) );
  NANDN U994 ( .A(n966), .B(n42173), .Z(n927) );
  NANDN U995 ( .A(n925), .B(n42172), .Z(n926) );
  NAND U996 ( .A(n927), .B(n926), .Z(n975) );
  NAND U997 ( .A(b[7]), .B(a[13]), .Z(n976) );
  XNOR U998 ( .A(n975), .B(n976), .Z(n978) );
  XOR U999 ( .A(n977), .B(n978), .Z(n984) );
  NANDN U1000 ( .A(n928), .B(n42093), .Z(n930) );
  XOR U1001 ( .A(n42134), .B(a[19]), .Z(n969) );
  NANDN U1002 ( .A(n969), .B(n42095), .Z(n929) );
  NAND U1003 ( .A(n930), .B(n929), .Z(n982) );
  NANDN U1004 ( .A(n931), .B(n42231), .Z(n933) );
  XOR U1005 ( .A(n163), .B(a[15]), .Z(n972) );
  NANDN U1006 ( .A(n972), .B(n42234), .Z(n932) );
  AND U1007 ( .A(n933), .B(n932), .Z(n981) );
  XNOR U1008 ( .A(n982), .B(n981), .Z(n983) );
  XNOR U1009 ( .A(n984), .B(n983), .Z(n988) );
  NANDN U1010 ( .A(n935), .B(n934), .Z(n939) );
  NAND U1011 ( .A(n937), .B(n936), .Z(n938) );
  AND U1012 ( .A(n939), .B(n938), .Z(n987) );
  XOR U1013 ( .A(n988), .B(n987), .Z(n989) );
  NANDN U1014 ( .A(n941), .B(n940), .Z(n945) );
  NANDN U1015 ( .A(n943), .B(n942), .Z(n944) );
  NAND U1016 ( .A(n945), .B(n944), .Z(n990) );
  XOR U1017 ( .A(n989), .B(n990), .Z(n957) );
  OR U1018 ( .A(n947), .B(n946), .Z(n951) );
  NANDN U1019 ( .A(n949), .B(n948), .Z(n950) );
  NAND U1020 ( .A(n951), .B(n950), .Z(n958) );
  XNOR U1021 ( .A(n957), .B(n958), .Z(n959) );
  XNOR U1022 ( .A(n960), .B(n959), .Z(n993) );
  XNOR U1023 ( .A(n993), .B(sreg[1037]), .Z(n995) );
  NAND U1024 ( .A(n952), .B(sreg[1036]), .Z(n956) );
  OR U1025 ( .A(n954), .B(n953), .Z(n955) );
  AND U1026 ( .A(n956), .B(n955), .Z(n994) );
  XOR U1027 ( .A(n995), .B(n994), .Z(c[1037]) );
  NANDN U1028 ( .A(n958), .B(n957), .Z(n962) );
  NAND U1029 ( .A(n960), .B(n959), .Z(n961) );
  NAND U1030 ( .A(n962), .B(n961), .Z(n1001) );
  NAND U1031 ( .A(b[0]), .B(a[22]), .Z(n963) );
  XNOR U1032 ( .A(b[1]), .B(n963), .Z(n965) );
  NAND U1033 ( .A(n18), .B(a[21]), .Z(n964) );
  AND U1034 ( .A(n965), .B(n964), .Z(n1018) );
  XOR U1035 ( .A(a[18]), .B(n42197), .Z(n1007) );
  NANDN U1036 ( .A(n1007), .B(n42173), .Z(n968) );
  NANDN U1037 ( .A(n966), .B(n42172), .Z(n967) );
  NAND U1038 ( .A(n968), .B(n967), .Z(n1016) );
  NAND U1039 ( .A(b[7]), .B(a[14]), .Z(n1017) );
  XNOR U1040 ( .A(n1016), .B(n1017), .Z(n1019) );
  XOR U1041 ( .A(n1018), .B(n1019), .Z(n1025) );
  NANDN U1042 ( .A(n969), .B(n42093), .Z(n971) );
  XOR U1043 ( .A(n42134), .B(a[20]), .Z(n1010) );
  NANDN U1044 ( .A(n1010), .B(n42095), .Z(n970) );
  NAND U1045 ( .A(n971), .B(n970), .Z(n1023) );
  NANDN U1046 ( .A(n972), .B(n42231), .Z(n974) );
  XOR U1047 ( .A(n163), .B(a[16]), .Z(n1013) );
  NANDN U1048 ( .A(n1013), .B(n42234), .Z(n973) );
  AND U1049 ( .A(n974), .B(n973), .Z(n1022) );
  XNOR U1050 ( .A(n1023), .B(n1022), .Z(n1024) );
  XNOR U1051 ( .A(n1025), .B(n1024), .Z(n1029) );
  NANDN U1052 ( .A(n976), .B(n975), .Z(n980) );
  NAND U1053 ( .A(n978), .B(n977), .Z(n979) );
  AND U1054 ( .A(n980), .B(n979), .Z(n1028) );
  XOR U1055 ( .A(n1029), .B(n1028), .Z(n1030) );
  NANDN U1056 ( .A(n982), .B(n981), .Z(n986) );
  NANDN U1057 ( .A(n984), .B(n983), .Z(n985) );
  NAND U1058 ( .A(n986), .B(n985), .Z(n1031) );
  XOR U1059 ( .A(n1030), .B(n1031), .Z(n998) );
  OR U1060 ( .A(n988), .B(n987), .Z(n992) );
  NANDN U1061 ( .A(n990), .B(n989), .Z(n991) );
  NAND U1062 ( .A(n992), .B(n991), .Z(n999) );
  XNOR U1063 ( .A(n998), .B(n999), .Z(n1000) );
  XNOR U1064 ( .A(n1001), .B(n1000), .Z(n1034) );
  XNOR U1065 ( .A(n1034), .B(sreg[1038]), .Z(n1036) );
  NAND U1066 ( .A(n993), .B(sreg[1037]), .Z(n997) );
  OR U1067 ( .A(n995), .B(n994), .Z(n996) );
  AND U1068 ( .A(n997), .B(n996), .Z(n1035) );
  XOR U1069 ( .A(n1036), .B(n1035), .Z(c[1038]) );
  NANDN U1070 ( .A(n999), .B(n998), .Z(n1003) );
  NAND U1071 ( .A(n1001), .B(n1000), .Z(n1002) );
  NAND U1072 ( .A(n1003), .B(n1002), .Z(n1042) );
  NAND U1073 ( .A(b[0]), .B(a[23]), .Z(n1004) );
  XNOR U1074 ( .A(b[1]), .B(n1004), .Z(n1006) );
  NAND U1075 ( .A(n18), .B(a[22]), .Z(n1005) );
  AND U1076 ( .A(n1006), .B(n1005), .Z(n1059) );
  XOR U1077 ( .A(a[19]), .B(n42197), .Z(n1048) );
  NANDN U1078 ( .A(n1048), .B(n42173), .Z(n1009) );
  NANDN U1079 ( .A(n1007), .B(n42172), .Z(n1008) );
  NAND U1080 ( .A(n1009), .B(n1008), .Z(n1057) );
  NAND U1081 ( .A(b[7]), .B(a[15]), .Z(n1058) );
  XNOR U1082 ( .A(n1057), .B(n1058), .Z(n1060) );
  XOR U1083 ( .A(n1059), .B(n1060), .Z(n1066) );
  NANDN U1084 ( .A(n1010), .B(n42093), .Z(n1012) );
  XOR U1085 ( .A(n42134), .B(a[21]), .Z(n1051) );
  NANDN U1086 ( .A(n1051), .B(n42095), .Z(n1011) );
  NAND U1087 ( .A(n1012), .B(n1011), .Z(n1064) );
  NANDN U1088 ( .A(n1013), .B(n42231), .Z(n1015) );
  XOR U1089 ( .A(n163), .B(a[17]), .Z(n1054) );
  NANDN U1090 ( .A(n1054), .B(n42234), .Z(n1014) );
  AND U1091 ( .A(n1015), .B(n1014), .Z(n1063) );
  XNOR U1092 ( .A(n1064), .B(n1063), .Z(n1065) );
  XNOR U1093 ( .A(n1066), .B(n1065), .Z(n1070) );
  NANDN U1094 ( .A(n1017), .B(n1016), .Z(n1021) );
  NAND U1095 ( .A(n1019), .B(n1018), .Z(n1020) );
  AND U1096 ( .A(n1021), .B(n1020), .Z(n1069) );
  XOR U1097 ( .A(n1070), .B(n1069), .Z(n1071) );
  NANDN U1098 ( .A(n1023), .B(n1022), .Z(n1027) );
  NANDN U1099 ( .A(n1025), .B(n1024), .Z(n1026) );
  NAND U1100 ( .A(n1027), .B(n1026), .Z(n1072) );
  XOR U1101 ( .A(n1071), .B(n1072), .Z(n1039) );
  OR U1102 ( .A(n1029), .B(n1028), .Z(n1033) );
  NANDN U1103 ( .A(n1031), .B(n1030), .Z(n1032) );
  NAND U1104 ( .A(n1033), .B(n1032), .Z(n1040) );
  XNOR U1105 ( .A(n1039), .B(n1040), .Z(n1041) );
  XNOR U1106 ( .A(n1042), .B(n1041), .Z(n1075) );
  XNOR U1107 ( .A(n1075), .B(sreg[1039]), .Z(n1077) );
  NAND U1108 ( .A(n1034), .B(sreg[1038]), .Z(n1038) );
  OR U1109 ( .A(n1036), .B(n1035), .Z(n1037) );
  AND U1110 ( .A(n1038), .B(n1037), .Z(n1076) );
  XOR U1111 ( .A(n1077), .B(n1076), .Z(c[1039]) );
  NANDN U1112 ( .A(n1040), .B(n1039), .Z(n1044) );
  NAND U1113 ( .A(n1042), .B(n1041), .Z(n1043) );
  NAND U1114 ( .A(n1044), .B(n1043), .Z(n1083) );
  NAND U1115 ( .A(b[0]), .B(a[24]), .Z(n1045) );
  XNOR U1116 ( .A(b[1]), .B(n1045), .Z(n1047) );
  NAND U1117 ( .A(n18), .B(a[23]), .Z(n1046) );
  AND U1118 ( .A(n1047), .B(n1046), .Z(n1100) );
  XOR U1119 ( .A(a[20]), .B(n42197), .Z(n1089) );
  NANDN U1120 ( .A(n1089), .B(n42173), .Z(n1050) );
  NANDN U1121 ( .A(n1048), .B(n42172), .Z(n1049) );
  NAND U1122 ( .A(n1050), .B(n1049), .Z(n1098) );
  NAND U1123 ( .A(b[7]), .B(a[16]), .Z(n1099) );
  XNOR U1124 ( .A(n1098), .B(n1099), .Z(n1101) );
  XOR U1125 ( .A(n1100), .B(n1101), .Z(n1107) );
  NANDN U1126 ( .A(n1051), .B(n42093), .Z(n1053) );
  XOR U1127 ( .A(n42134), .B(a[22]), .Z(n1092) );
  NANDN U1128 ( .A(n1092), .B(n42095), .Z(n1052) );
  NAND U1129 ( .A(n1053), .B(n1052), .Z(n1105) );
  NANDN U1130 ( .A(n1054), .B(n42231), .Z(n1056) );
  XOR U1131 ( .A(n163), .B(a[18]), .Z(n1095) );
  NANDN U1132 ( .A(n1095), .B(n42234), .Z(n1055) );
  AND U1133 ( .A(n1056), .B(n1055), .Z(n1104) );
  XNOR U1134 ( .A(n1105), .B(n1104), .Z(n1106) );
  XNOR U1135 ( .A(n1107), .B(n1106), .Z(n1111) );
  NANDN U1136 ( .A(n1058), .B(n1057), .Z(n1062) );
  NAND U1137 ( .A(n1060), .B(n1059), .Z(n1061) );
  AND U1138 ( .A(n1062), .B(n1061), .Z(n1110) );
  XOR U1139 ( .A(n1111), .B(n1110), .Z(n1112) );
  NANDN U1140 ( .A(n1064), .B(n1063), .Z(n1068) );
  NANDN U1141 ( .A(n1066), .B(n1065), .Z(n1067) );
  NAND U1142 ( .A(n1068), .B(n1067), .Z(n1113) );
  XOR U1143 ( .A(n1112), .B(n1113), .Z(n1080) );
  OR U1144 ( .A(n1070), .B(n1069), .Z(n1074) );
  NANDN U1145 ( .A(n1072), .B(n1071), .Z(n1073) );
  NAND U1146 ( .A(n1074), .B(n1073), .Z(n1081) );
  XNOR U1147 ( .A(n1080), .B(n1081), .Z(n1082) );
  XNOR U1148 ( .A(n1083), .B(n1082), .Z(n1116) );
  XNOR U1149 ( .A(n1116), .B(sreg[1040]), .Z(n1118) );
  NAND U1150 ( .A(n1075), .B(sreg[1039]), .Z(n1079) );
  OR U1151 ( .A(n1077), .B(n1076), .Z(n1078) );
  AND U1152 ( .A(n1079), .B(n1078), .Z(n1117) );
  XOR U1153 ( .A(n1118), .B(n1117), .Z(c[1040]) );
  NANDN U1154 ( .A(n1081), .B(n1080), .Z(n1085) );
  NAND U1155 ( .A(n1083), .B(n1082), .Z(n1084) );
  NAND U1156 ( .A(n1085), .B(n1084), .Z(n1124) );
  NAND U1157 ( .A(b[0]), .B(a[25]), .Z(n1086) );
  XNOR U1158 ( .A(b[1]), .B(n1086), .Z(n1088) );
  NAND U1159 ( .A(n18), .B(a[24]), .Z(n1087) );
  AND U1160 ( .A(n1088), .B(n1087), .Z(n1141) );
  XOR U1161 ( .A(a[21]), .B(n42197), .Z(n1130) );
  NANDN U1162 ( .A(n1130), .B(n42173), .Z(n1091) );
  NANDN U1163 ( .A(n1089), .B(n42172), .Z(n1090) );
  NAND U1164 ( .A(n1091), .B(n1090), .Z(n1139) );
  NAND U1165 ( .A(b[7]), .B(a[17]), .Z(n1140) );
  XNOR U1166 ( .A(n1139), .B(n1140), .Z(n1142) );
  XOR U1167 ( .A(n1141), .B(n1142), .Z(n1148) );
  NANDN U1168 ( .A(n1092), .B(n42093), .Z(n1094) );
  XOR U1169 ( .A(n42134), .B(a[23]), .Z(n1133) );
  NANDN U1170 ( .A(n1133), .B(n42095), .Z(n1093) );
  NAND U1171 ( .A(n1094), .B(n1093), .Z(n1146) );
  NANDN U1172 ( .A(n1095), .B(n42231), .Z(n1097) );
  XOR U1173 ( .A(n163), .B(a[19]), .Z(n1136) );
  NANDN U1174 ( .A(n1136), .B(n42234), .Z(n1096) );
  AND U1175 ( .A(n1097), .B(n1096), .Z(n1145) );
  XNOR U1176 ( .A(n1146), .B(n1145), .Z(n1147) );
  XNOR U1177 ( .A(n1148), .B(n1147), .Z(n1152) );
  NANDN U1178 ( .A(n1099), .B(n1098), .Z(n1103) );
  NAND U1179 ( .A(n1101), .B(n1100), .Z(n1102) );
  AND U1180 ( .A(n1103), .B(n1102), .Z(n1151) );
  XOR U1181 ( .A(n1152), .B(n1151), .Z(n1153) );
  NANDN U1182 ( .A(n1105), .B(n1104), .Z(n1109) );
  NANDN U1183 ( .A(n1107), .B(n1106), .Z(n1108) );
  NAND U1184 ( .A(n1109), .B(n1108), .Z(n1154) );
  XOR U1185 ( .A(n1153), .B(n1154), .Z(n1121) );
  OR U1186 ( .A(n1111), .B(n1110), .Z(n1115) );
  NANDN U1187 ( .A(n1113), .B(n1112), .Z(n1114) );
  NAND U1188 ( .A(n1115), .B(n1114), .Z(n1122) );
  XNOR U1189 ( .A(n1121), .B(n1122), .Z(n1123) );
  XNOR U1190 ( .A(n1124), .B(n1123), .Z(n1157) );
  XNOR U1191 ( .A(n1157), .B(sreg[1041]), .Z(n1159) );
  NAND U1192 ( .A(n1116), .B(sreg[1040]), .Z(n1120) );
  OR U1193 ( .A(n1118), .B(n1117), .Z(n1119) );
  AND U1194 ( .A(n1120), .B(n1119), .Z(n1158) );
  XOR U1195 ( .A(n1159), .B(n1158), .Z(c[1041]) );
  NANDN U1196 ( .A(n1122), .B(n1121), .Z(n1126) );
  NAND U1197 ( .A(n1124), .B(n1123), .Z(n1125) );
  NAND U1198 ( .A(n1126), .B(n1125), .Z(n1165) );
  NAND U1199 ( .A(b[0]), .B(a[26]), .Z(n1127) );
  XNOR U1200 ( .A(b[1]), .B(n1127), .Z(n1129) );
  NAND U1201 ( .A(n18), .B(a[25]), .Z(n1128) );
  AND U1202 ( .A(n1129), .B(n1128), .Z(n1182) );
  XOR U1203 ( .A(a[22]), .B(n42197), .Z(n1171) );
  NANDN U1204 ( .A(n1171), .B(n42173), .Z(n1132) );
  NANDN U1205 ( .A(n1130), .B(n42172), .Z(n1131) );
  NAND U1206 ( .A(n1132), .B(n1131), .Z(n1180) );
  NAND U1207 ( .A(b[7]), .B(a[18]), .Z(n1181) );
  XNOR U1208 ( .A(n1180), .B(n1181), .Z(n1183) );
  XOR U1209 ( .A(n1182), .B(n1183), .Z(n1189) );
  NANDN U1210 ( .A(n1133), .B(n42093), .Z(n1135) );
  XOR U1211 ( .A(n42134), .B(a[24]), .Z(n1174) );
  NANDN U1212 ( .A(n1174), .B(n42095), .Z(n1134) );
  NAND U1213 ( .A(n1135), .B(n1134), .Z(n1187) );
  NANDN U1214 ( .A(n1136), .B(n42231), .Z(n1138) );
  XOR U1215 ( .A(n163), .B(a[20]), .Z(n1177) );
  NANDN U1216 ( .A(n1177), .B(n42234), .Z(n1137) );
  AND U1217 ( .A(n1138), .B(n1137), .Z(n1186) );
  XNOR U1218 ( .A(n1187), .B(n1186), .Z(n1188) );
  XNOR U1219 ( .A(n1189), .B(n1188), .Z(n1193) );
  NANDN U1220 ( .A(n1140), .B(n1139), .Z(n1144) );
  NAND U1221 ( .A(n1142), .B(n1141), .Z(n1143) );
  AND U1222 ( .A(n1144), .B(n1143), .Z(n1192) );
  XOR U1223 ( .A(n1193), .B(n1192), .Z(n1194) );
  NANDN U1224 ( .A(n1146), .B(n1145), .Z(n1150) );
  NANDN U1225 ( .A(n1148), .B(n1147), .Z(n1149) );
  NAND U1226 ( .A(n1150), .B(n1149), .Z(n1195) );
  XOR U1227 ( .A(n1194), .B(n1195), .Z(n1162) );
  OR U1228 ( .A(n1152), .B(n1151), .Z(n1156) );
  NANDN U1229 ( .A(n1154), .B(n1153), .Z(n1155) );
  NAND U1230 ( .A(n1156), .B(n1155), .Z(n1163) );
  XNOR U1231 ( .A(n1162), .B(n1163), .Z(n1164) );
  XNOR U1232 ( .A(n1165), .B(n1164), .Z(n1198) );
  XNOR U1233 ( .A(n1198), .B(sreg[1042]), .Z(n1200) );
  NAND U1234 ( .A(n1157), .B(sreg[1041]), .Z(n1161) );
  OR U1235 ( .A(n1159), .B(n1158), .Z(n1160) );
  AND U1236 ( .A(n1161), .B(n1160), .Z(n1199) );
  XOR U1237 ( .A(n1200), .B(n1199), .Z(c[1042]) );
  NANDN U1238 ( .A(n1163), .B(n1162), .Z(n1167) );
  NAND U1239 ( .A(n1165), .B(n1164), .Z(n1166) );
  NAND U1240 ( .A(n1167), .B(n1166), .Z(n1206) );
  NAND U1241 ( .A(b[0]), .B(a[27]), .Z(n1168) );
  XNOR U1242 ( .A(b[1]), .B(n1168), .Z(n1170) );
  NAND U1243 ( .A(n18), .B(a[26]), .Z(n1169) );
  AND U1244 ( .A(n1170), .B(n1169), .Z(n1223) );
  XOR U1245 ( .A(a[23]), .B(n42197), .Z(n1212) );
  NANDN U1246 ( .A(n1212), .B(n42173), .Z(n1173) );
  NANDN U1247 ( .A(n1171), .B(n42172), .Z(n1172) );
  NAND U1248 ( .A(n1173), .B(n1172), .Z(n1221) );
  NAND U1249 ( .A(b[7]), .B(a[19]), .Z(n1222) );
  XNOR U1250 ( .A(n1221), .B(n1222), .Z(n1224) );
  XOR U1251 ( .A(n1223), .B(n1224), .Z(n1230) );
  NANDN U1252 ( .A(n1174), .B(n42093), .Z(n1176) );
  XOR U1253 ( .A(n42134), .B(a[25]), .Z(n1215) );
  NANDN U1254 ( .A(n1215), .B(n42095), .Z(n1175) );
  NAND U1255 ( .A(n1176), .B(n1175), .Z(n1228) );
  NANDN U1256 ( .A(n1177), .B(n42231), .Z(n1179) );
  XOR U1257 ( .A(n163), .B(a[21]), .Z(n1218) );
  NANDN U1258 ( .A(n1218), .B(n42234), .Z(n1178) );
  AND U1259 ( .A(n1179), .B(n1178), .Z(n1227) );
  XNOR U1260 ( .A(n1228), .B(n1227), .Z(n1229) );
  XNOR U1261 ( .A(n1230), .B(n1229), .Z(n1234) );
  NANDN U1262 ( .A(n1181), .B(n1180), .Z(n1185) );
  NAND U1263 ( .A(n1183), .B(n1182), .Z(n1184) );
  AND U1264 ( .A(n1185), .B(n1184), .Z(n1233) );
  XOR U1265 ( .A(n1234), .B(n1233), .Z(n1235) );
  NANDN U1266 ( .A(n1187), .B(n1186), .Z(n1191) );
  NANDN U1267 ( .A(n1189), .B(n1188), .Z(n1190) );
  NAND U1268 ( .A(n1191), .B(n1190), .Z(n1236) );
  XOR U1269 ( .A(n1235), .B(n1236), .Z(n1203) );
  OR U1270 ( .A(n1193), .B(n1192), .Z(n1197) );
  NANDN U1271 ( .A(n1195), .B(n1194), .Z(n1196) );
  NAND U1272 ( .A(n1197), .B(n1196), .Z(n1204) );
  XNOR U1273 ( .A(n1203), .B(n1204), .Z(n1205) );
  XNOR U1274 ( .A(n1206), .B(n1205), .Z(n1239) );
  XNOR U1275 ( .A(n1239), .B(sreg[1043]), .Z(n1241) );
  NAND U1276 ( .A(n1198), .B(sreg[1042]), .Z(n1202) );
  OR U1277 ( .A(n1200), .B(n1199), .Z(n1201) );
  AND U1278 ( .A(n1202), .B(n1201), .Z(n1240) );
  XOR U1279 ( .A(n1241), .B(n1240), .Z(c[1043]) );
  NANDN U1280 ( .A(n1204), .B(n1203), .Z(n1208) );
  NAND U1281 ( .A(n1206), .B(n1205), .Z(n1207) );
  NAND U1282 ( .A(n1208), .B(n1207), .Z(n1247) );
  NAND U1283 ( .A(b[0]), .B(a[28]), .Z(n1209) );
  XNOR U1284 ( .A(b[1]), .B(n1209), .Z(n1211) );
  NAND U1285 ( .A(n19), .B(a[27]), .Z(n1210) );
  AND U1286 ( .A(n1211), .B(n1210), .Z(n1264) );
  XOR U1287 ( .A(a[24]), .B(n42197), .Z(n1253) );
  NANDN U1288 ( .A(n1253), .B(n42173), .Z(n1214) );
  NANDN U1289 ( .A(n1212), .B(n42172), .Z(n1213) );
  NAND U1290 ( .A(n1214), .B(n1213), .Z(n1262) );
  NAND U1291 ( .A(b[7]), .B(a[20]), .Z(n1263) );
  XNOR U1292 ( .A(n1262), .B(n1263), .Z(n1265) );
  XOR U1293 ( .A(n1264), .B(n1265), .Z(n1271) );
  NANDN U1294 ( .A(n1215), .B(n42093), .Z(n1217) );
  XOR U1295 ( .A(n42134), .B(a[26]), .Z(n1256) );
  NANDN U1296 ( .A(n1256), .B(n42095), .Z(n1216) );
  NAND U1297 ( .A(n1217), .B(n1216), .Z(n1269) );
  NANDN U1298 ( .A(n1218), .B(n42231), .Z(n1220) );
  XOR U1299 ( .A(n163), .B(a[22]), .Z(n1259) );
  NANDN U1300 ( .A(n1259), .B(n42234), .Z(n1219) );
  AND U1301 ( .A(n1220), .B(n1219), .Z(n1268) );
  XNOR U1302 ( .A(n1269), .B(n1268), .Z(n1270) );
  XNOR U1303 ( .A(n1271), .B(n1270), .Z(n1275) );
  NANDN U1304 ( .A(n1222), .B(n1221), .Z(n1226) );
  NAND U1305 ( .A(n1224), .B(n1223), .Z(n1225) );
  AND U1306 ( .A(n1226), .B(n1225), .Z(n1274) );
  XOR U1307 ( .A(n1275), .B(n1274), .Z(n1276) );
  NANDN U1308 ( .A(n1228), .B(n1227), .Z(n1232) );
  NANDN U1309 ( .A(n1230), .B(n1229), .Z(n1231) );
  NAND U1310 ( .A(n1232), .B(n1231), .Z(n1277) );
  XOR U1311 ( .A(n1276), .B(n1277), .Z(n1244) );
  OR U1312 ( .A(n1234), .B(n1233), .Z(n1238) );
  NANDN U1313 ( .A(n1236), .B(n1235), .Z(n1237) );
  NAND U1314 ( .A(n1238), .B(n1237), .Z(n1245) );
  XNOR U1315 ( .A(n1244), .B(n1245), .Z(n1246) );
  XNOR U1316 ( .A(n1247), .B(n1246), .Z(n1280) );
  XNOR U1317 ( .A(n1280), .B(sreg[1044]), .Z(n1282) );
  NAND U1318 ( .A(n1239), .B(sreg[1043]), .Z(n1243) );
  OR U1319 ( .A(n1241), .B(n1240), .Z(n1242) );
  AND U1320 ( .A(n1243), .B(n1242), .Z(n1281) );
  XOR U1321 ( .A(n1282), .B(n1281), .Z(c[1044]) );
  NANDN U1322 ( .A(n1245), .B(n1244), .Z(n1249) );
  NAND U1323 ( .A(n1247), .B(n1246), .Z(n1248) );
  NAND U1324 ( .A(n1249), .B(n1248), .Z(n1288) );
  NAND U1325 ( .A(b[0]), .B(a[29]), .Z(n1250) );
  XNOR U1326 ( .A(b[1]), .B(n1250), .Z(n1252) );
  NAND U1327 ( .A(n19), .B(a[28]), .Z(n1251) );
  AND U1328 ( .A(n1252), .B(n1251), .Z(n1305) );
  XOR U1329 ( .A(a[25]), .B(n42197), .Z(n1294) );
  NANDN U1330 ( .A(n1294), .B(n42173), .Z(n1255) );
  NANDN U1331 ( .A(n1253), .B(n42172), .Z(n1254) );
  NAND U1332 ( .A(n1255), .B(n1254), .Z(n1303) );
  NAND U1333 ( .A(b[7]), .B(a[21]), .Z(n1304) );
  XNOR U1334 ( .A(n1303), .B(n1304), .Z(n1306) );
  XOR U1335 ( .A(n1305), .B(n1306), .Z(n1312) );
  NANDN U1336 ( .A(n1256), .B(n42093), .Z(n1258) );
  XOR U1337 ( .A(n42134), .B(a[27]), .Z(n1297) );
  NANDN U1338 ( .A(n1297), .B(n42095), .Z(n1257) );
  NAND U1339 ( .A(n1258), .B(n1257), .Z(n1310) );
  NANDN U1340 ( .A(n1259), .B(n42231), .Z(n1261) );
  XOR U1341 ( .A(n164), .B(a[23]), .Z(n1300) );
  NANDN U1342 ( .A(n1300), .B(n42234), .Z(n1260) );
  AND U1343 ( .A(n1261), .B(n1260), .Z(n1309) );
  XNOR U1344 ( .A(n1310), .B(n1309), .Z(n1311) );
  XNOR U1345 ( .A(n1312), .B(n1311), .Z(n1316) );
  NANDN U1346 ( .A(n1263), .B(n1262), .Z(n1267) );
  NAND U1347 ( .A(n1265), .B(n1264), .Z(n1266) );
  AND U1348 ( .A(n1267), .B(n1266), .Z(n1315) );
  XOR U1349 ( .A(n1316), .B(n1315), .Z(n1317) );
  NANDN U1350 ( .A(n1269), .B(n1268), .Z(n1273) );
  NANDN U1351 ( .A(n1271), .B(n1270), .Z(n1272) );
  NAND U1352 ( .A(n1273), .B(n1272), .Z(n1318) );
  XOR U1353 ( .A(n1317), .B(n1318), .Z(n1285) );
  OR U1354 ( .A(n1275), .B(n1274), .Z(n1279) );
  NANDN U1355 ( .A(n1277), .B(n1276), .Z(n1278) );
  NAND U1356 ( .A(n1279), .B(n1278), .Z(n1286) );
  XNOR U1357 ( .A(n1285), .B(n1286), .Z(n1287) );
  XNOR U1358 ( .A(n1288), .B(n1287), .Z(n1321) );
  XNOR U1359 ( .A(n1321), .B(sreg[1045]), .Z(n1323) );
  NAND U1360 ( .A(n1280), .B(sreg[1044]), .Z(n1284) );
  OR U1361 ( .A(n1282), .B(n1281), .Z(n1283) );
  AND U1362 ( .A(n1284), .B(n1283), .Z(n1322) );
  XOR U1363 ( .A(n1323), .B(n1322), .Z(c[1045]) );
  NANDN U1364 ( .A(n1286), .B(n1285), .Z(n1290) );
  NAND U1365 ( .A(n1288), .B(n1287), .Z(n1289) );
  NAND U1366 ( .A(n1290), .B(n1289), .Z(n1329) );
  NAND U1367 ( .A(b[0]), .B(a[30]), .Z(n1291) );
  XNOR U1368 ( .A(b[1]), .B(n1291), .Z(n1293) );
  NAND U1369 ( .A(n19), .B(a[29]), .Z(n1292) );
  AND U1370 ( .A(n1293), .B(n1292), .Z(n1346) );
  XOR U1371 ( .A(a[26]), .B(n42197), .Z(n1335) );
  NANDN U1372 ( .A(n1335), .B(n42173), .Z(n1296) );
  NANDN U1373 ( .A(n1294), .B(n42172), .Z(n1295) );
  NAND U1374 ( .A(n1296), .B(n1295), .Z(n1344) );
  NAND U1375 ( .A(b[7]), .B(a[22]), .Z(n1345) );
  XNOR U1376 ( .A(n1344), .B(n1345), .Z(n1347) );
  XOR U1377 ( .A(n1346), .B(n1347), .Z(n1353) );
  NANDN U1378 ( .A(n1297), .B(n42093), .Z(n1299) );
  XOR U1379 ( .A(n42134), .B(a[28]), .Z(n1338) );
  NANDN U1380 ( .A(n1338), .B(n42095), .Z(n1298) );
  NAND U1381 ( .A(n1299), .B(n1298), .Z(n1351) );
  NANDN U1382 ( .A(n1300), .B(n42231), .Z(n1302) );
  XOR U1383 ( .A(n164), .B(a[24]), .Z(n1341) );
  NANDN U1384 ( .A(n1341), .B(n42234), .Z(n1301) );
  AND U1385 ( .A(n1302), .B(n1301), .Z(n1350) );
  XNOR U1386 ( .A(n1351), .B(n1350), .Z(n1352) );
  XNOR U1387 ( .A(n1353), .B(n1352), .Z(n1357) );
  NANDN U1388 ( .A(n1304), .B(n1303), .Z(n1308) );
  NAND U1389 ( .A(n1306), .B(n1305), .Z(n1307) );
  AND U1390 ( .A(n1308), .B(n1307), .Z(n1356) );
  XOR U1391 ( .A(n1357), .B(n1356), .Z(n1358) );
  NANDN U1392 ( .A(n1310), .B(n1309), .Z(n1314) );
  NANDN U1393 ( .A(n1312), .B(n1311), .Z(n1313) );
  NAND U1394 ( .A(n1314), .B(n1313), .Z(n1359) );
  XOR U1395 ( .A(n1358), .B(n1359), .Z(n1326) );
  OR U1396 ( .A(n1316), .B(n1315), .Z(n1320) );
  NANDN U1397 ( .A(n1318), .B(n1317), .Z(n1319) );
  NAND U1398 ( .A(n1320), .B(n1319), .Z(n1327) );
  XNOR U1399 ( .A(n1326), .B(n1327), .Z(n1328) );
  XNOR U1400 ( .A(n1329), .B(n1328), .Z(n1362) );
  XNOR U1401 ( .A(n1362), .B(sreg[1046]), .Z(n1364) );
  NAND U1402 ( .A(n1321), .B(sreg[1045]), .Z(n1325) );
  OR U1403 ( .A(n1323), .B(n1322), .Z(n1324) );
  AND U1404 ( .A(n1325), .B(n1324), .Z(n1363) );
  XOR U1405 ( .A(n1364), .B(n1363), .Z(c[1046]) );
  NANDN U1406 ( .A(n1327), .B(n1326), .Z(n1331) );
  NAND U1407 ( .A(n1329), .B(n1328), .Z(n1330) );
  NAND U1408 ( .A(n1331), .B(n1330), .Z(n1370) );
  NAND U1409 ( .A(b[0]), .B(a[31]), .Z(n1332) );
  XNOR U1410 ( .A(b[1]), .B(n1332), .Z(n1334) );
  NAND U1411 ( .A(n19), .B(a[30]), .Z(n1333) );
  AND U1412 ( .A(n1334), .B(n1333), .Z(n1387) );
  XOR U1413 ( .A(a[27]), .B(n42197), .Z(n1376) );
  NANDN U1414 ( .A(n1376), .B(n42173), .Z(n1337) );
  NANDN U1415 ( .A(n1335), .B(n42172), .Z(n1336) );
  NAND U1416 ( .A(n1337), .B(n1336), .Z(n1385) );
  NAND U1417 ( .A(b[7]), .B(a[23]), .Z(n1386) );
  XNOR U1418 ( .A(n1385), .B(n1386), .Z(n1388) );
  XOR U1419 ( .A(n1387), .B(n1388), .Z(n1394) );
  NANDN U1420 ( .A(n1338), .B(n42093), .Z(n1340) );
  XOR U1421 ( .A(n42134), .B(a[29]), .Z(n1379) );
  NANDN U1422 ( .A(n1379), .B(n42095), .Z(n1339) );
  NAND U1423 ( .A(n1340), .B(n1339), .Z(n1392) );
  NANDN U1424 ( .A(n1341), .B(n42231), .Z(n1343) );
  XOR U1425 ( .A(n164), .B(a[25]), .Z(n1382) );
  NANDN U1426 ( .A(n1382), .B(n42234), .Z(n1342) );
  AND U1427 ( .A(n1343), .B(n1342), .Z(n1391) );
  XNOR U1428 ( .A(n1392), .B(n1391), .Z(n1393) );
  XNOR U1429 ( .A(n1394), .B(n1393), .Z(n1398) );
  NANDN U1430 ( .A(n1345), .B(n1344), .Z(n1349) );
  NAND U1431 ( .A(n1347), .B(n1346), .Z(n1348) );
  AND U1432 ( .A(n1349), .B(n1348), .Z(n1397) );
  XOR U1433 ( .A(n1398), .B(n1397), .Z(n1399) );
  NANDN U1434 ( .A(n1351), .B(n1350), .Z(n1355) );
  NANDN U1435 ( .A(n1353), .B(n1352), .Z(n1354) );
  NAND U1436 ( .A(n1355), .B(n1354), .Z(n1400) );
  XOR U1437 ( .A(n1399), .B(n1400), .Z(n1367) );
  OR U1438 ( .A(n1357), .B(n1356), .Z(n1361) );
  NANDN U1439 ( .A(n1359), .B(n1358), .Z(n1360) );
  NAND U1440 ( .A(n1361), .B(n1360), .Z(n1368) );
  XNOR U1441 ( .A(n1367), .B(n1368), .Z(n1369) );
  XNOR U1442 ( .A(n1370), .B(n1369), .Z(n1403) );
  XNOR U1443 ( .A(n1403), .B(sreg[1047]), .Z(n1405) );
  NAND U1444 ( .A(n1362), .B(sreg[1046]), .Z(n1366) );
  OR U1445 ( .A(n1364), .B(n1363), .Z(n1365) );
  AND U1446 ( .A(n1366), .B(n1365), .Z(n1404) );
  XOR U1447 ( .A(n1405), .B(n1404), .Z(c[1047]) );
  NANDN U1448 ( .A(n1368), .B(n1367), .Z(n1372) );
  NAND U1449 ( .A(n1370), .B(n1369), .Z(n1371) );
  NAND U1450 ( .A(n1372), .B(n1371), .Z(n1411) );
  NAND U1451 ( .A(b[0]), .B(a[32]), .Z(n1373) );
  XNOR U1452 ( .A(b[1]), .B(n1373), .Z(n1375) );
  NAND U1453 ( .A(n19), .B(a[31]), .Z(n1374) );
  AND U1454 ( .A(n1375), .B(n1374), .Z(n1428) );
  XOR U1455 ( .A(a[28]), .B(n42197), .Z(n1417) );
  NANDN U1456 ( .A(n1417), .B(n42173), .Z(n1378) );
  NANDN U1457 ( .A(n1376), .B(n42172), .Z(n1377) );
  NAND U1458 ( .A(n1378), .B(n1377), .Z(n1426) );
  NAND U1459 ( .A(b[7]), .B(a[24]), .Z(n1427) );
  XNOR U1460 ( .A(n1426), .B(n1427), .Z(n1429) );
  XOR U1461 ( .A(n1428), .B(n1429), .Z(n1435) );
  NANDN U1462 ( .A(n1379), .B(n42093), .Z(n1381) );
  XOR U1463 ( .A(n42134), .B(a[30]), .Z(n1420) );
  NANDN U1464 ( .A(n1420), .B(n42095), .Z(n1380) );
  NAND U1465 ( .A(n1381), .B(n1380), .Z(n1433) );
  NANDN U1466 ( .A(n1382), .B(n42231), .Z(n1384) );
  XOR U1467 ( .A(n164), .B(a[26]), .Z(n1423) );
  NANDN U1468 ( .A(n1423), .B(n42234), .Z(n1383) );
  AND U1469 ( .A(n1384), .B(n1383), .Z(n1432) );
  XNOR U1470 ( .A(n1433), .B(n1432), .Z(n1434) );
  XNOR U1471 ( .A(n1435), .B(n1434), .Z(n1439) );
  NANDN U1472 ( .A(n1386), .B(n1385), .Z(n1390) );
  NAND U1473 ( .A(n1388), .B(n1387), .Z(n1389) );
  AND U1474 ( .A(n1390), .B(n1389), .Z(n1438) );
  XOR U1475 ( .A(n1439), .B(n1438), .Z(n1440) );
  NANDN U1476 ( .A(n1392), .B(n1391), .Z(n1396) );
  NANDN U1477 ( .A(n1394), .B(n1393), .Z(n1395) );
  NAND U1478 ( .A(n1396), .B(n1395), .Z(n1441) );
  XOR U1479 ( .A(n1440), .B(n1441), .Z(n1408) );
  OR U1480 ( .A(n1398), .B(n1397), .Z(n1402) );
  NANDN U1481 ( .A(n1400), .B(n1399), .Z(n1401) );
  NAND U1482 ( .A(n1402), .B(n1401), .Z(n1409) );
  XNOR U1483 ( .A(n1408), .B(n1409), .Z(n1410) );
  XNOR U1484 ( .A(n1411), .B(n1410), .Z(n1444) );
  XNOR U1485 ( .A(n1444), .B(sreg[1048]), .Z(n1446) );
  NAND U1486 ( .A(n1403), .B(sreg[1047]), .Z(n1407) );
  OR U1487 ( .A(n1405), .B(n1404), .Z(n1406) );
  AND U1488 ( .A(n1407), .B(n1406), .Z(n1445) );
  XOR U1489 ( .A(n1446), .B(n1445), .Z(c[1048]) );
  NANDN U1490 ( .A(n1409), .B(n1408), .Z(n1413) );
  NAND U1491 ( .A(n1411), .B(n1410), .Z(n1412) );
  NAND U1492 ( .A(n1413), .B(n1412), .Z(n1452) );
  NAND U1493 ( .A(b[0]), .B(a[33]), .Z(n1414) );
  XNOR U1494 ( .A(b[1]), .B(n1414), .Z(n1416) );
  NAND U1495 ( .A(n19), .B(a[32]), .Z(n1415) );
  AND U1496 ( .A(n1416), .B(n1415), .Z(n1469) );
  XOR U1497 ( .A(a[29]), .B(n42197), .Z(n1458) );
  NANDN U1498 ( .A(n1458), .B(n42173), .Z(n1419) );
  NANDN U1499 ( .A(n1417), .B(n42172), .Z(n1418) );
  NAND U1500 ( .A(n1419), .B(n1418), .Z(n1467) );
  NAND U1501 ( .A(b[7]), .B(a[25]), .Z(n1468) );
  XNOR U1502 ( .A(n1467), .B(n1468), .Z(n1470) );
  XOR U1503 ( .A(n1469), .B(n1470), .Z(n1476) );
  NANDN U1504 ( .A(n1420), .B(n42093), .Z(n1422) );
  XOR U1505 ( .A(n42134), .B(a[31]), .Z(n1461) );
  NANDN U1506 ( .A(n1461), .B(n42095), .Z(n1421) );
  NAND U1507 ( .A(n1422), .B(n1421), .Z(n1474) );
  NANDN U1508 ( .A(n1423), .B(n42231), .Z(n1425) );
  XOR U1509 ( .A(n164), .B(a[27]), .Z(n1464) );
  NANDN U1510 ( .A(n1464), .B(n42234), .Z(n1424) );
  AND U1511 ( .A(n1425), .B(n1424), .Z(n1473) );
  XNOR U1512 ( .A(n1474), .B(n1473), .Z(n1475) );
  XNOR U1513 ( .A(n1476), .B(n1475), .Z(n1480) );
  NANDN U1514 ( .A(n1427), .B(n1426), .Z(n1431) );
  NAND U1515 ( .A(n1429), .B(n1428), .Z(n1430) );
  AND U1516 ( .A(n1431), .B(n1430), .Z(n1479) );
  XOR U1517 ( .A(n1480), .B(n1479), .Z(n1481) );
  NANDN U1518 ( .A(n1433), .B(n1432), .Z(n1437) );
  NANDN U1519 ( .A(n1435), .B(n1434), .Z(n1436) );
  NAND U1520 ( .A(n1437), .B(n1436), .Z(n1482) );
  XOR U1521 ( .A(n1481), .B(n1482), .Z(n1449) );
  OR U1522 ( .A(n1439), .B(n1438), .Z(n1443) );
  NANDN U1523 ( .A(n1441), .B(n1440), .Z(n1442) );
  NAND U1524 ( .A(n1443), .B(n1442), .Z(n1450) );
  XNOR U1525 ( .A(n1449), .B(n1450), .Z(n1451) );
  XNOR U1526 ( .A(n1452), .B(n1451), .Z(n1485) );
  XNOR U1527 ( .A(n1485), .B(sreg[1049]), .Z(n1487) );
  NAND U1528 ( .A(n1444), .B(sreg[1048]), .Z(n1448) );
  OR U1529 ( .A(n1446), .B(n1445), .Z(n1447) );
  AND U1530 ( .A(n1448), .B(n1447), .Z(n1486) );
  XOR U1531 ( .A(n1487), .B(n1486), .Z(c[1049]) );
  NANDN U1532 ( .A(n1450), .B(n1449), .Z(n1454) );
  NAND U1533 ( .A(n1452), .B(n1451), .Z(n1453) );
  NAND U1534 ( .A(n1454), .B(n1453), .Z(n1493) );
  NAND U1535 ( .A(b[0]), .B(a[34]), .Z(n1455) );
  XNOR U1536 ( .A(b[1]), .B(n1455), .Z(n1457) );
  NAND U1537 ( .A(n19), .B(a[33]), .Z(n1456) );
  AND U1538 ( .A(n1457), .B(n1456), .Z(n1510) );
  XOR U1539 ( .A(a[30]), .B(n42197), .Z(n1499) );
  NANDN U1540 ( .A(n1499), .B(n42173), .Z(n1460) );
  NANDN U1541 ( .A(n1458), .B(n42172), .Z(n1459) );
  NAND U1542 ( .A(n1460), .B(n1459), .Z(n1508) );
  NAND U1543 ( .A(b[7]), .B(a[26]), .Z(n1509) );
  XNOR U1544 ( .A(n1508), .B(n1509), .Z(n1511) );
  XOR U1545 ( .A(n1510), .B(n1511), .Z(n1517) );
  NANDN U1546 ( .A(n1461), .B(n42093), .Z(n1463) );
  XOR U1547 ( .A(n42134), .B(a[32]), .Z(n1502) );
  NANDN U1548 ( .A(n1502), .B(n42095), .Z(n1462) );
  NAND U1549 ( .A(n1463), .B(n1462), .Z(n1515) );
  NANDN U1550 ( .A(n1464), .B(n42231), .Z(n1466) );
  XOR U1551 ( .A(n164), .B(a[28]), .Z(n1505) );
  NANDN U1552 ( .A(n1505), .B(n42234), .Z(n1465) );
  AND U1553 ( .A(n1466), .B(n1465), .Z(n1514) );
  XNOR U1554 ( .A(n1515), .B(n1514), .Z(n1516) );
  XNOR U1555 ( .A(n1517), .B(n1516), .Z(n1521) );
  NANDN U1556 ( .A(n1468), .B(n1467), .Z(n1472) );
  NAND U1557 ( .A(n1470), .B(n1469), .Z(n1471) );
  AND U1558 ( .A(n1472), .B(n1471), .Z(n1520) );
  XOR U1559 ( .A(n1521), .B(n1520), .Z(n1522) );
  NANDN U1560 ( .A(n1474), .B(n1473), .Z(n1478) );
  NANDN U1561 ( .A(n1476), .B(n1475), .Z(n1477) );
  NAND U1562 ( .A(n1478), .B(n1477), .Z(n1523) );
  XOR U1563 ( .A(n1522), .B(n1523), .Z(n1490) );
  OR U1564 ( .A(n1480), .B(n1479), .Z(n1484) );
  NANDN U1565 ( .A(n1482), .B(n1481), .Z(n1483) );
  NAND U1566 ( .A(n1484), .B(n1483), .Z(n1491) );
  XNOR U1567 ( .A(n1490), .B(n1491), .Z(n1492) );
  XNOR U1568 ( .A(n1493), .B(n1492), .Z(n1526) );
  XNOR U1569 ( .A(n1526), .B(sreg[1050]), .Z(n1528) );
  NAND U1570 ( .A(n1485), .B(sreg[1049]), .Z(n1489) );
  OR U1571 ( .A(n1487), .B(n1486), .Z(n1488) );
  AND U1572 ( .A(n1489), .B(n1488), .Z(n1527) );
  XOR U1573 ( .A(n1528), .B(n1527), .Z(c[1050]) );
  NANDN U1574 ( .A(n1491), .B(n1490), .Z(n1495) );
  NAND U1575 ( .A(n1493), .B(n1492), .Z(n1494) );
  NAND U1576 ( .A(n1495), .B(n1494), .Z(n1534) );
  NAND U1577 ( .A(b[0]), .B(a[35]), .Z(n1496) );
  XNOR U1578 ( .A(b[1]), .B(n1496), .Z(n1498) );
  NAND U1579 ( .A(n20), .B(a[34]), .Z(n1497) );
  AND U1580 ( .A(n1498), .B(n1497), .Z(n1551) );
  XOR U1581 ( .A(a[31]), .B(n42197), .Z(n1540) );
  NANDN U1582 ( .A(n1540), .B(n42173), .Z(n1501) );
  NANDN U1583 ( .A(n1499), .B(n42172), .Z(n1500) );
  NAND U1584 ( .A(n1501), .B(n1500), .Z(n1549) );
  NAND U1585 ( .A(b[7]), .B(a[27]), .Z(n1550) );
  XNOR U1586 ( .A(n1549), .B(n1550), .Z(n1552) );
  XOR U1587 ( .A(n1551), .B(n1552), .Z(n1558) );
  NANDN U1588 ( .A(n1502), .B(n42093), .Z(n1504) );
  XOR U1589 ( .A(n42134), .B(a[33]), .Z(n1543) );
  NANDN U1590 ( .A(n1543), .B(n42095), .Z(n1503) );
  NAND U1591 ( .A(n1504), .B(n1503), .Z(n1556) );
  NANDN U1592 ( .A(n1505), .B(n42231), .Z(n1507) );
  XOR U1593 ( .A(n164), .B(a[29]), .Z(n1546) );
  NANDN U1594 ( .A(n1546), .B(n42234), .Z(n1506) );
  AND U1595 ( .A(n1507), .B(n1506), .Z(n1555) );
  XNOR U1596 ( .A(n1556), .B(n1555), .Z(n1557) );
  XNOR U1597 ( .A(n1558), .B(n1557), .Z(n1562) );
  NANDN U1598 ( .A(n1509), .B(n1508), .Z(n1513) );
  NAND U1599 ( .A(n1511), .B(n1510), .Z(n1512) );
  AND U1600 ( .A(n1513), .B(n1512), .Z(n1561) );
  XOR U1601 ( .A(n1562), .B(n1561), .Z(n1563) );
  NANDN U1602 ( .A(n1515), .B(n1514), .Z(n1519) );
  NANDN U1603 ( .A(n1517), .B(n1516), .Z(n1518) );
  NAND U1604 ( .A(n1519), .B(n1518), .Z(n1564) );
  XOR U1605 ( .A(n1563), .B(n1564), .Z(n1531) );
  OR U1606 ( .A(n1521), .B(n1520), .Z(n1525) );
  NANDN U1607 ( .A(n1523), .B(n1522), .Z(n1524) );
  NAND U1608 ( .A(n1525), .B(n1524), .Z(n1532) );
  XNOR U1609 ( .A(n1531), .B(n1532), .Z(n1533) );
  XNOR U1610 ( .A(n1534), .B(n1533), .Z(n1567) );
  XNOR U1611 ( .A(n1567), .B(sreg[1051]), .Z(n1569) );
  NAND U1612 ( .A(n1526), .B(sreg[1050]), .Z(n1530) );
  OR U1613 ( .A(n1528), .B(n1527), .Z(n1529) );
  AND U1614 ( .A(n1530), .B(n1529), .Z(n1568) );
  XOR U1615 ( .A(n1569), .B(n1568), .Z(c[1051]) );
  NANDN U1616 ( .A(n1532), .B(n1531), .Z(n1536) );
  NAND U1617 ( .A(n1534), .B(n1533), .Z(n1535) );
  NAND U1618 ( .A(n1536), .B(n1535), .Z(n1575) );
  NAND U1619 ( .A(b[0]), .B(a[36]), .Z(n1537) );
  XNOR U1620 ( .A(b[1]), .B(n1537), .Z(n1539) );
  NAND U1621 ( .A(n20), .B(a[35]), .Z(n1538) );
  AND U1622 ( .A(n1539), .B(n1538), .Z(n1592) );
  XOR U1623 ( .A(a[32]), .B(n42197), .Z(n1581) );
  NANDN U1624 ( .A(n1581), .B(n42173), .Z(n1542) );
  NANDN U1625 ( .A(n1540), .B(n42172), .Z(n1541) );
  NAND U1626 ( .A(n1542), .B(n1541), .Z(n1590) );
  NAND U1627 ( .A(b[7]), .B(a[28]), .Z(n1591) );
  XNOR U1628 ( .A(n1590), .B(n1591), .Z(n1593) );
  XOR U1629 ( .A(n1592), .B(n1593), .Z(n1599) );
  NANDN U1630 ( .A(n1543), .B(n42093), .Z(n1545) );
  XOR U1631 ( .A(n42134), .B(a[34]), .Z(n1584) );
  NANDN U1632 ( .A(n1584), .B(n42095), .Z(n1544) );
  NAND U1633 ( .A(n1545), .B(n1544), .Z(n1597) );
  NANDN U1634 ( .A(n1546), .B(n42231), .Z(n1548) );
  XOR U1635 ( .A(n164), .B(a[30]), .Z(n1587) );
  NANDN U1636 ( .A(n1587), .B(n42234), .Z(n1547) );
  AND U1637 ( .A(n1548), .B(n1547), .Z(n1596) );
  XNOR U1638 ( .A(n1597), .B(n1596), .Z(n1598) );
  XNOR U1639 ( .A(n1599), .B(n1598), .Z(n1603) );
  NANDN U1640 ( .A(n1550), .B(n1549), .Z(n1554) );
  NAND U1641 ( .A(n1552), .B(n1551), .Z(n1553) );
  AND U1642 ( .A(n1554), .B(n1553), .Z(n1602) );
  XOR U1643 ( .A(n1603), .B(n1602), .Z(n1604) );
  NANDN U1644 ( .A(n1556), .B(n1555), .Z(n1560) );
  NANDN U1645 ( .A(n1558), .B(n1557), .Z(n1559) );
  NAND U1646 ( .A(n1560), .B(n1559), .Z(n1605) );
  XOR U1647 ( .A(n1604), .B(n1605), .Z(n1572) );
  OR U1648 ( .A(n1562), .B(n1561), .Z(n1566) );
  NANDN U1649 ( .A(n1564), .B(n1563), .Z(n1565) );
  NAND U1650 ( .A(n1566), .B(n1565), .Z(n1573) );
  XNOR U1651 ( .A(n1572), .B(n1573), .Z(n1574) );
  XNOR U1652 ( .A(n1575), .B(n1574), .Z(n1608) );
  XNOR U1653 ( .A(n1608), .B(sreg[1052]), .Z(n1610) );
  NAND U1654 ( .A(n1567), .B(sreg[1051]), .Z(n1571) );
  OR U1655 ( .A(n1569), .B(n1568), .Z(n1570) );
  AND U1656 ( .A(n1571), .B(n1570), .Z(n1609) );
  XOR U1657 ( .A(n1610), .B(n1609), .Z(c[1052]) );
  NANDN U1658 ( .A(n1573), .B(n1572), .Z(n1577) );
  NAND U1659 ( .A(n1575), .B(n1574), .Z(n1576) );
  NAND U1660 ( .A(n1577), .B(n1576), .Z(n1616) );
  NAND U1661 ( .A(b[0]), .B(a[37]), .Z(n1578) );
  XNOR U1662 ( .A(b[1]), .B(n1578), .Z(n1580) );
  NAND U1663 ( .A(n20), .B(a[36]), .Z(n1579) );
  AND U1664 ( .A(n1580), .B(n1579), .Z(n1633) );
  XOR U1665 ( .A(a[33]), .B(n42197), .Z(n1622) );
  NANDN U1666 ( .A(n1622), .B(n42173), .Z(n1583) );
  NANDN U1667 ( .A(n1581), .B(n42172), .Z(n1582) );
  NAND U1668 ( .A(n1583), .B(n1582), .Z(n1631) );
  NAND U1669 ( .A(b[7]), .B(a[29]), .Z(n1632) );
  XNOR U1670 ( .A(n1631), .B(n1632), .Z(n1634) );
  XOR U1671 ( .A(n1633), .B(n1634), .Z(n1640) );
  NANDN U1672 ( .A(n1584), .B(n42093), .Z(n1586) );
  XOR U1673 ( .A(n42134), .B(a[35]), .Z(n1625) );
  NANDN U1674 ( .A(n1625), .B(n42095), .Z(n1585) );
  NAND U1675 ( .A(n1586), .B(n1585), .Z(n1638) );
  NANDN U1676 ( .A(n1587), .B(n42231), .Z(n1589) );
  XOR U1677 ( .A(n164), .B(a[31]), .Z(n1628) );
  NANDN U1678 ( .A(n1628), .B(n42234), .Z(n1588) );
  AND U1679 ( .A(n1589), .B(n1588), .Z(n1637) );
  XNOR U1680 ( .A(n1638), .B(n1637), .Z(n1639) );
  XNOR U1681 ( .A(n1640), .B(n1639), .Z(n1644) );
  NANDN U1682 ( .A(n1591), .B(n1590), .Z(n1595) );
  NAND U1683 ( .A(n1593), .B(n1592), .Z(n1594) );
  AND U1684 ( .A(n1595), .B(n1594), .Z(n1643) );
  XOR U1685 ( .A(n1644), .B(n1643), .Z(n1645) );
  NANDN U1686 ( .A(n1597), .B(n1596), .Z(n1601) );
  NANDN U1687 ( .A(n1599), .B(n1598), .Z(n1600) );
  NAND U1688 ( .A(n1601), .B(n1600), .Z(n1646) );
  XOR U1689 ( .A(n1645), .B(n1646), .Z(n1613) );
  OR U1690 ( .A(n1603), .B(n1602), .Z(n1607) );
  NANDN U1691 ( .A(n1605), .B(n1604), .Z(n1606) );
  NAND U1692 ( .A(n1607), .B(n1606), .Z(n1614) );
  XNOR U1693 ( .A(n1613), .B(n1614), .Z(n1615) );
  XNOR U1694 ( .A(n1616), .B(n1615), .Z(n1649) );
  XNOR U1695 ( .A(n1649), .B(sreg[1053]), .Z(n1651) );
  NAND U1696 ( .A(n1608), .B(sreg[1052]), .Z(n1612) );
  OR U1697 ( .A(n1610), .B(n1609), .Z(n1611) );
  AND U1698 ( .A(n1612), .B(n1611), .Z(n1650) );
  XOR U1699 ( .A(n1651), .B(n1650), .Z(c[1053]) );
  NANDN U1700 ( .A(n1614), .B(n1613), .Z(n1618) );
  NAND U1701 ( .A(n1616), .B(n1615), .Z(n1617) );
  NAND U1702 ( .A(n1618), .B(n1617), .Z(n1657) );
  NAND U1703 ( .A(b[0]), .B(a[38]), .Z(n1619) );
  XNOR U1704 ( .A(b[1]), .B(n1619), .Z(n1621) );
  NAND U1705 ( .A(n20), .B(a[37]), .Z(n1620) );
  AND U1706 ( .A(n1621), .B(n1620), .Z(n1674) );
  XOR U1707 ( .A(a[34]), .B(n42197), .Z(n1663) );
  NANDN U1708 ( .A(n1663), .B(n42173), .Z(n1624) );
  NANDN U1709 ( .A(n1622), .B(n42172), .Z(n1623) );
  NAND U1710 ( .A(n1624), .B(n1623), .Z(n1672) );
  NAND U1711 ( .A(b[7]), .B(a[30]), .Z(n1673) );
  XNOR U1712 ( .A(n1672), .B(n1673), .Z(n1675) );
  XOR U1713 ( .A(n1674), .B(n1675), .Z(n1681) );
  NANDN U1714 ( .A(n1625), .B(n42093), .Z(n1627) );
  XOR U1715 ( .A(n42134), .B(a[36]), .Z(n1666) );
  NANDN U1716 ( .A(n1666), .B(n42095), .Z(n1626) );
  NAND U1717 ( .A(n1627), .B(n1626), .Z(n1679) );
  NANDN U1718 ( .A(n1628), .B(n42231), .Z(n1630) );
  XOR U1719 ( .A(n164), .B(a[32]), .Z(n1669) );
  NANDN U1720 ( .A(n1669), .B(n42234), .Z(n1629) );
  AND U1721 ( .A(n1630), .B(n1629), .Z(n1678) );
  XNOR U1722 ( .A(n1679), .B(n1678), .Z(n1680) );
  XNOR U1723 ( .A(n1681), .B(n1680), .Z(n1685) );
  NANDN U1724 ( .A(n1632), .B(n1631), .Z(n1636) );
  NAND U1725 ( .A(n1634), .B(n1633), .Z(n1635) );
  AND U1726 ( .A(n1636), .B(n1635), .Z(n1684) );
  XOR U1727 ( .A(n1685), .B(n1684), .Z(n1686) );
  NANDN U1728 ( .A(n1638), .B(n1637), .Z(n1642) );
  NANDN U1729 ( .A(n1640), .B(n1639), .Z(n1641) );
  NAND U1730 ( .A(n1642), .B(n1641), .Z(n1687) );
  XOR U1731 ( .A(n1686), .B(n1687), .Z(n1654) );
  OR U1732 ( .A(n1644), .B(n1643), .Z(n1648) );
  NANDN U1733 ( .A(n1646), .B(n1645), .Z(n1647) );
  NAND U1734 ( .A(n1648), .B(n1647), .Z(n1655) );
  XNOR U1735 ( .A(n1654), .B(n1655), .Z(n1656) );
  XNOR U1736 ( .A(n1657), .B(n1656), .Z(n1690) );
  XNOR U1737 ( .A(n1690), .B(sreg[1054]), .Z(n1692) );
  NAND U1738 ( .A(n1649), .B(sreg[1053]), .Z(n1653) );
  OR U1739 ( .A(n1651), .B(n1650), .Z(n1652) );
  AND U1740 ( .A(n1653), .B(n1652), .Z(n1691) );
  XOR U1741 ( .A(n1692), .B(n1691), .Z(c[1054]) );
  NANDN U1742 ( .A(n1655), .B(n1654), .Z(n1659) );
  NAND U1743 ( .A(n1657), .B(n1656), .Z(n1658) );
  NAND U1744 ( .A(n1659), .B(n1658), .Z(n1698) );
  NAND U1745 ( .A(b[0]), .B(a[39]), .Z(n1660) );
  XNOR U1746 ( .A(b[1]), .B(n1660), .Z(n1662) );
  NAND U1747 ( .A(n20), .B(a[38]), .Z(n1661) );
  AND U1748 ( .A(n1662), .B(n1661), .Z(n1715) );
  XOR U1749 ( .A(a[35]), .B(n42197), .Z(n1704) );
  NANDN U1750 ( .A(n1704), .B(n42173), .Z(n1665) );
  NANDN U1751 ( .A(n1663), .B(n42172), .Z(n1664) );
  NAND U1752 ( .A(n1665), .B(n1664), .Z(n1713) );
  NAND U1753 ( .A(b[7]), .B(a[31]), .Z(n1714) );
  XNOR U1754 ( .A(n1713), .B(n1714), .Z(n1716) );
  XOR U1755 ( .A(n1715), .B(n1716), .Z(n1722) );
  NANDN U1756 ( .A(n1666), .B(n42093), .Z(n1668) );
  XOR U1757 ( .A(n42134), .B(a[37]), .Z(n1707) );
  NANDN U1758 ( .A(n1707), .B(n42095), .Z(n1667) );
  NAND U1759 ( .A(n1668), .B(n1667), .Z(n1720) );
  NANDN U1760 ( .A(n1669), .B(n42231), .Z(n1671) );
  XOR U1761 ( .A(n164), .B(a[33]), .Z(n1710) );
  NANDN U1762 ( .A(n1710), .B(n42234), .Z(n1670) );
  AND U1763 ( .A(n1671), .B(n1670), .Z(n1719) );
  XNOR U1764 ( .A(n1720), .B(n1719), .Z(n1721) );
  XNOR U1765 ( .A(n1722), .B(n1721), .Z(n1726) );
  NANDN U1766 ( .A(n1673), .B(n1672), .Z(n1677) );
  NAND U1767 ( .A(n1675), .B(n1674), .Z(n1676) );
  AND U1768 ( .A(n1677), .B(n1676), .Z(n1725) );
  XOR U1769 ( .A(n1726), .B(n1725), .Z(n1727) );
  NANDN U1770 ( .A(n1679), .B(n1678), .Z(n1683) );
  NANDN U1771 ( .A(n1681), .B(n1680), .Z(n1682) );
  NAND U1772 ( .A(n1683), .B(n1682), .Z(n1728) );
  XOR U1773 ( .A(n1727), .B(n1728), .Z(n1695) );
  OR U1774 ( .A(n1685), .B(n1684), .Z(n1689) );
  NANDN U1775 ( .A(n1687), .B(n1686), .Z(n1688) );
  NAND U1776 ( .A(n1689), .B(n1688), .Z(n1696) );
  XNOR U1777 ( .A(n1695), .B(n1696), .Z(n1697) );
  XNOR U1778 ( .A(n1698), .B(n1697), .Z(n1731) );
  XNOR U1779 ( .A(n1731), .B(sreg[1055]), .Z(n1733) );
  NAND U1780 ( .A(n1690), .B(sreg[1054]), .Z(n1694) );
  OR U1781 ( .A(n1692), .B(n1691), .Z(n1693) );
  AND U1782 ( .A(n1694), .B(n1693), .Z(n1732) );
  XOR U1783 ( .A(n1733), .B(n1732), .Z(c[1055]) );
  NANDN U1784 ( .A(n1696), .B(n1695), .Z(n1700) );
  NAND U1785 ( .A(n1698), .B(n1697), .Z(n1699) );
  NAND U1786 ( .A(n1700), .B(n1699), .Z(n1739) );
  NAND U1787 ( .A(b[0]), .B(a[40]), .Z(n1701) );
  XNOR U1788 ( .A(b[1]), .B(n1701), .Z(n1703) );
  NAND U1789 ( .A(n20), .B(a[39]), .Z(n1702) );
  AND U1790 ( .A(n1703), .B(n1702), .Z(n1756) );
  XOR U1791 ( .A(a[36]), .B(n42197), .Z(n1745) );
  NANDN U1792 ( .A(n1745), .B(n42173), .Z(n1706) );
  NANDN U1793 ( .A(n1704), .B(n42172), .Z(n1705) );
  NAND U1794 ( .A(n1706), .B(n1705), .Z(n1754) );
  NAND U1795 ( .A(b[7]), .B(a[32]), .Z(n1755) );
  XNOR U1796 ( .A(n1754), .B(n1755), .Z(n1757) );
  XOR U1797 ( .A(n1756), .B(n1757), .Z(n1763) );
  NANDN U1798 ( .A(n1707), .B(n42093), .Z(n1709) );
  XOR U1799 ( .A(n42134), .B(a[38]), .Z(n1748) );
  NANDN U1800 ( .A(n1748), .B(n42095), .Z(n1708) );
  NAND U1801 ( .A(n1709), .B(n1708), .Z(n1761) );
  NANDN U1802 ( .A(n1710), .B(n42231), .Z(n1712) );
  XOR U1803 ( .A(n164), .B(a[34]), .Z(n1751) );
  NANDN U1804 ( .A(n1751), .B(n42234), .Z(n1711) );
  AND U1805 ( .A(n1712), .B(n1711), .Z(n1760) );
  XNOR U1806 ( .A(n1761), .B(n1760), .Z(n1762) );
  XNOR U1807 ( .A(n1763), .B(n1762), .Z(n1767) );
  NANDN U1808 ( .A(n1714), .B(n1713), .Z(n1718) );
  NAND U1809 ( .A(n1716), .B(n1715), .Z(n1717) );
  AND U1810 ( .A(n1718), .B(n1717), .Z(n1766) );
  XOR U1811 ( .A(n1767), .B(n1766), .Z(n1768) );
  NANDN U1812 ( .A(n1720), .B(n1719), .Z(n1724) );
  NANDN U1813 ( .A(n1722), .B(n1721), .Z(n1723) );
  NAND U1814 ( .A(n1724), .B(n1723), .Z(n1769) );
  XOR U1815 ( .A(n1768), .B(n1769), .Z(n1736) );
  OR U1816 ( .A(n1726), .B(n1725), .Z(n1730) );
  NANDN U1817 ( .A(n1728), .B(n1727), .Z(n1729) );
  NAND U1818 ( .A(n1730), .B(n1729), .Z(n1737) );
  XNOR U1819 ( .A(n1736), .B(n1737), .Z(n1738) );
  XNOR U1820 ( .A(n1739), .B(n1738), .Z(n1772) );
  XNOR U1821 ( .A(n1772), .B(sreg[1056]), .Z(n1774) );
  NAND U1822 ( .A(n1731), .B(sreg[1055]), .Z(n1735) );
  OR U1823 ( .A(n1733), .B(n1732), .Z(n1734) );
  AND U1824 ( .A(n1735), .B(n1734), .Z(n1773) );
  XOR U1825 ( .A(n1774), .B(n1773), .Z(c[1056]) );
  NANDN U1826 ( .A(n1737), .B(n1736), .Z(n1741) );
  NAND U1827 ( .A(n1739), .B(n1738), .Z(n1740) );
  NAND U1828 ( .A(n1741), .B(n1740), .Z(n1780) );
  NAND U1829 ( .A(b[0]), .B(a[41]), .Z(n1742) );
  XNOR U1830 ( .A(b[1]), .B(n1742), .Z(n1744) );
  NAND U1831 ( .A(n20), .B(a[40]), .Z(n1743) );
  AND U1832 ( .A(n1744), .B(n1743), .Z(n1797) );
  XOR U1833 ( .A(a[37]), .B(n42197), .Z(n1786) );
  NANDN U1834 ( .A(n1786), .B(n42173), .Z(n1747) );
  NANDN U1835 ( .A(n1745), .B(n42172), .Z(n1746) );
  NAND U1836 ( .A(n1747), .B(n1746), .Z(n1795) );
  NAND U1837 ( .A(b[7]), .B(a[33]), .Z(n1796) );
  XNOR U1838 ( .A(n1795), .B(n1796), .Z(n1798) );
  XOR U1839 ( .A(n1797), .B(n1798), .Z(n1804) );
  NANDN U1840 ( .A(n1748), .B(n42093), .Z(n1750) );
  XOR U1841 ( .A(n42134), .B(a[39]), .Z(n1789) );
  NANDN U1842 ( .A(n1789), .B(n42095), .Z(n1749) );
  NAND U1843 ( .A(n1750), .B(n1749), .Z(n1802) );
  NANDN U1844 ( .A(n1751), .B(n42231), .Z(n1753) );
  XOR U1845 ( .A(n165), .B(a[35]), .Z(n1792) );
  NANDN U1846 ( .A(n1792), .B(n42234), .Z(n1752) );
  AND U1847 ( .A(n1753), .B(n1752), .Z(n1801) );
  XNOR U1848 ( .A(n1802), .B(n1801), .Z(n1803) );
  XNOR U1849 ( .A(n1804), .B(n1803), .Z(n1808) );
  NANDN U1850 ( .A(n1755), .B(n1754), .Z(n1759) );
  NAND U1851 ( .A(n1757), .B(n1756), .Z(n1758) );
  AND U1852 ( .A(n1759), .B(n1758), .Z(n1807) );
  XOR U1853 ( .A(n1808), .B(n1807), .Z(n1809) );
  NANDN U1854 ( .A(n1761), .B(n1760), .Z(n1765) );
  NANDN U1855 ( .A(n1763), .B(n1762), .Z(n1764) );
  NAND U1856 ( .A(n1765), .B(n1764), .Z(n1810) );
  XOR U1857 ( .A(n1809), .B(n1810), .Z(n1777) );
  OR U1858 ( .A(n1767), .B(n1766), .Z(n1771) );
  NANDN U1859 ( .A(n1769), .B(n1768), .Z(n1770) );
  NAND U1860 ( .A(n1771), .B(n1770), .Z(n1778) );
  XNOR U1861 ( .A(n1777), .B(n1778), .Z(n1779) );
  XNOR U1862 ( .A(n1780), .B(n1779), .Z(n1813) );
  XNOR U1863 ( .A(n1813), .B(sreg[1057]), .Z(n1815) );
  NAND U1864 ( .A(n1772), .B(sreg[1056]), .Z(n1776) );
  OR U1865 ( .A(n1774), .B(n1773), .Z(n1775) );
  AND U1866 ( .A(n1776), .B(n1775), .Z(n1814) );
  XOR U1867 ( .A(n1815), .B(n1814), .Z(c[1057]) );
  NANDN U1868 ( .A(n1778), .B(n1777), .Z(n1782) );
  NAND U1869 ( .A(n1780), .B(n1779), .Z(n1781) );
  NAND U1870 ( .A(n1782), .B(n1781), .Z(n1821) );
  NAND U1871 ( .A(b[0]), .B(a[42]), .Z(n1783) );
  XNOR U1872 ( .A(b[1]), .B(n1783), .Z(n1785) );
  NAND U1873 ( .A(n21), .B(a[41]), .Z(n1784) );
  AND U1874 ( .A(n1785), .B(n1784), .Z(n1838) );
  XOR U1875 ( .A(a[38]), .B(n42197), .Z(n1827) );
  NANDN U1876 ( .A(n1827), .B(n42173), .Z(n1788) );
  NANDN U1877 ( .A(n1786), .B(n42172), .Z(n1787) );
  NAND U1878 ( .A(n1788), .B(n1787), .Z(n1836) );
  NAND U1879 ( .A(b[7]), .B(a[34]), .Z(n1837) );
  XNOR U1880 ( .A(n1836), .B(n1837), .Z(n1839) );
  XOR U1881 ( .A(n1838), .B(n1839), .Z(n1845) );
  NANDN U1882 ( .A(n1789), .B(n42093), .Z(n1791) );
  XOR U1883 ( .A(n42134), .B(a[40]), .Z(n1830) );
  NANDN U1884 ( .A(n1830), .B(n42095), .Z(n1790) );
  NAND U1885 ( .A(n1791), .B(n1790), .Z(n1843) );
  NANDN U1886 ( .A(n1792), .B(n42231), .Z(n1794) );
  XOR U1887 ( .A(n165), .B(a[36]), .Z(n1833) );
  NANDN U1888 ( .A(n1833), .B(n42234), .Z(n1793) );
  AND U1889 ( .A(n1794), .B(n1793), .Z(n1842) );
  XNOR U1890 ( .A(n1843), .B(n1842), .Z(n1844) );
  XNOR U1891 ( .A(n1845), .B(n1844), .Z(n1849) );
  NANDN U1892 ( .A(n1796), .B(n1795), .Z(n1800) );
  NAND U1893 ( .A(n1798), .B(n1797), .Z(n1799) );
  AND U1894 ( .A(n1800), .B(n1799), .Z(n1848) );
  XOR U1895 ( .A(n1849), .B(n1848), .Z(n1850) );
  NANDN U1896 ( .A(n1802), .B(n1801), .Z(n1806) );
  NANDN U1897 ( .A(n1804), .B(n1803), .Z(n1805) );
  NAND U1898 ( .A(n1806), .B(n1805), .Z(n1851) );
  XOR U1899 ( .A(n1850), .B(n1851), .Z(n1818) );
  OR U1900 ( .A(n1808), .B(n1807), .Z(n1812) );
  NANDN U1901 ( .A(n1810), .B(n1809), .Z(n1811) );
  NAND U1902 ( .A(n1812), .B(n1811), .Z(n1819) );
  XNOR U1903 ( .A(n1818), .B(n1819), .Z(n1820) );
  XNOR U1904 ( .A(n1821), .B(n1820), .Z(n1854) );
  XNOR U1905 ( .A(n1854), .B(sreg[1058]), .Z(n1856) );
  NAND U1906 ( .A(n1813), .B(sreg[1057]), .Z(n1817) );
  OR U1907 ( .A(n1815), .B(n1814), .Z(n1816) );
  AND U1908 ( .A(n1817), .B(n1816), .Z(n1855) );
  XOR U1909 ( .A(n1856), .B(n1855), .Z(c[1058]) );
  NANDN U1910 ( .A(n1819), .B(n1818), .Z(n1823) );
  NAND U1911 ( .A(n1821), .B(n1820), .Z(n1822) );
  NAND U1912 ( .A(n1823), .B(n1822), .Z(n1862) );
  NAND U1913 ( .A(b[0]), .B(a[43]), .Z(n1824) );
  XNOR U1914 ( .A(b[1]), .B(n1824), .Z(n1826) );
  NAND U1915 ( .A(n21), .B(a[42]), .Z(n1825) );
  AND U1916 ( .A(n1826), .B(n1825), .Z(n1879) );
  XOR U1917 ( .A(a[39]), .B(n42197), .Z(n1868) );
  NANDN U1918 ( .A(n1868), .B(n42173), .Z(n1829) );
  NANDN U1919 ( .A(n1827), .B(n42172), .Z(n1828) );
  NAND U1920 ( .A(n1829), .B(n1828), .Z(n1877) );
  NAND U1921 ( .A(b[7]), .B(a[35]), .Z(n1878) );
  XNOR U1922 ( .A(n1877), .B(n1878), .Z(n1880) );
  XOR U1923 ( .A(n1879), .B(n1880), .Z(n1886) );
  NANDN U1924 ( .A(n1830), .B(n42093), .Z(n1832) );
  XOR U1925 ( .A(n42134), .B(a[41]), .Z(n1871) );
  NANDN U1926 ( .A(n1871), .B(n42095), .Z(n1831) );
  NAND U1927 ( .A(n1832), .B(n1831), .Z(n1884) );
  NANDN U1928 ( .A(n1833), .B(n42231), .Z(n1835) );
  XOR U1929 ( .A(n165), .B(a[37]), .Z(n1874) );
  NANDN U1930 ( .A(n1874), .B(n42234), .Z(n1834) );
  AND U1931 ( .A(n1835), .B(n1834), .Z(n1883) );
  XNOR U1932 ( .A(n1884), .B(n1883), .Z(n1885) );
  XNOR U1933 ( .A(n1886), .B(n1885), .Z(n1890) );
  NANDN U1934 ( .A(n1837), .B(n1836), .Z(n1841) );
  NAND U1935 ( .A(n1839), .B(n1838), .Z(n1840) );
  AND U1936 ( .A(n1841), .B(n1840), .Z(n1889) );
  XOR U1937 ( .A(n1890), .B(n1889), .Z(n1891) );
  NANDN U1938 ( .A(n1843), .B(n1842), .Z(n1847) );
  NANDN U1939 ( .A(n1845), .B(n1844), .Z(n1846) );
  NAND U1940 ( .A(n1847), .B(n1846), .Z(n1892) );
  XOR U1941 ( .A(n1891), .B(n1892), .Z(n1859) );
  OR U1942 ( .A(n1849), .B(n1848), .Z(n1853) );
  NANDN U1943 ( .A(n1851), .B(n1850), .Z(n1852) );
  NAND U1944 ( .A(n1853), .B(n1852), .Z(n1860) );
  XNOR U1945 ( .A(n1859), .B(n1860), .Z(n1861) );
  XNOR U1946 ( .A(n1862), .B(n1861), .Z(n1895) );
  XNOR U1947 ( .A(n1895), .B(sreg[1059]), .Z(n1897) );
  NAND U1948 ( .A(n1854), .B(sreg[1058]), .Z(n1858) );
  OR U1949 ( .A(n1856), .B(n1855), .Z(n1857) );
  AND U1950 ( .A(n1858), .B(n1857), .Z(n1896) );
  XOR U1951 ( .A(n1897), .B(n1896), .Z(c[1059]) );
  NANDN U1952 ( .A(n1860), .B(n1859), .Z(n1864) );
  NAND U1953 ( .A(n1862), .B(n1861), .Z(n1863) );
  NAND U1954 ( .A(n1864), .B(n1863), .Z(n1903) );
  NAND U1955 ( .A(b[0]), .B(a[44]), .Z(n1865) );
  XNOR U1956 ( .A(b[1]), .B(n1865), .Z(n1867) );
  NAND U1957 ( .A(n21), .B(a[43]), .Z(n1866) );
  AND U1958 ( .A(n1867), .B(n1866), .Z(n1920) );
  XOR U1959 ( .A(a[40]), .B(n42197), .Z(n1909) );
  NANDN U1960 ( .A(n1909), .B(n42173), .Z(n1870) );
  NANDN U1961 ( .A(n1868), .B(n42172), .Z(n1869) );
  NAND U1962 ( .A(n1870), .B(n1869), .Z(n1918) );
  NAND U1963 ( .A(b[7]), .B(a[36]), .Z(n1919) );
  XNOR U1964 ( .A(n1918), .B(n1919), .Z(n1921) );
  XOR U1965 ( .A(n1920), .B(n1921), .Z(n1927) );
  NANDN U1966 ( .A(n1871), .B(n42093), .Z(n1873) );
  XOR U1967 ( .A(n42134), .B(a[42]), .Z(n1912) );
  NANDN U1968 ( .A(n1912), .B(n42095), .Z(n1872) );
  NAND U1969 ( .A(n1873), .B(n1872), .Z(n1925) );
  NANDN U1970 ( .A(n1874), .B(n42231), .Z(n1876) );
  XOR U1971 ( .A(n165), .B(a[38]), .Z(n1915) );
  NANDN U1972 ( .A(n1915), .B(n42234), .Z(n1875) );
  AND U1973 ( .A(n1876), .B(n1875), .Z(n1924) );
  XNOR U1974 ( .A(n1925), .B(n1924), .Z(n1926) );
  XNOR U1975 ( .A(n1927), .B(n1926), .Z(n1931) );
  NANDN U1976 ( .A(n1878), .B(n1877), .Z(n1882) );
  NAND U1977 ( .A(n1880), .B(n1879), .Z(n1881) );
  AND U1978 ( .A(n1882), .B(n1881), .Z(n1930) );
  XOR U1979 ( .A(n1931), .B(n1930), .Z(n1932) );
  NANDN U1980 ( .A(n1884), .B(n1883), .Z(n1888) );
  NANDN U1981 ( .A(n1886), .B(n1885), .Z(n1887) );
  NAND U1982 ( .A(n1888), .B(n1887), .Z(n1933) );
  XOR U1983 ( .A(n1932), .B(n1933), .Z(n1900) );
  OR U1984 ( .A(n1890), .B(n1889), .Z(n1894) );
  NANDN U1985 ( .A(n1892), .B(n1891), .Z(n1893) );
  NAND U1986 ( .A(n1894), .B(n1893), .Z(n1901) );
  XNOR U1987 ( .A(n1900), .B(n1901), .Z(n1902) );
  XNOR U1988 ( .A(n1903), .B(n1902), .Z(n1936) );
  XNOR U1989 ( .A(n1936), .B(sreg[1060]), .Z(n1938) );
  NAND U1990 ( .A(n1895), .B(sreg[1059]), .Z(n1899) );
  OR U1991 ( .A(n1897), .B(n1896), .Z(n1898) );
  AND U1992 ( .A(n1899), .B(n1898), .Z(n1937) );
  XOR U1993 ( .A(n1938), .B(n1937), .Z(c[1060]) );
  NANDN U1994 ( .A(n1901), .B(n1900), .Z(n1905) );
  NAND U1995 ( .A(n1903), .B(n1902), .Z(n1904) );
  NAND U1996 ( .A(n1905), .B(n1904), .Z(n1944) );
  NAND U1997 ( .A(b[0]), .B(a[45]), .Z(n1906) );
  XNOR U1998 ( .A(b[1]), .B(n1906), .Z(n1908) );
  NAND U1999 ( .A(n21), .B(a[44]), .Z(n1907) );
  AND U2000 ( .A(n1908), .B(n1907), .Z(n1961) );
  XOR U2001 ( .A(a[41]), .B(n42197), .Z(n1950) );
  NANDN U2002 ( .A(n1950), .B(n42173), .Z(n1911) );
  NANDN U2003 ( .A(n1909), .B(n42172), .Z(n1910) );
  NAND U2004 ( .A(n1911), .B(n1910), .Z(n1959) );
  NAND U2005 ( .A(b[7]), .B(a[37]), .Z(n1960) );
  XNOR U2006 ( .A(n1959), .B(n1960), .Z(n1962) );
  XOR U2007 ( .A(n1961), .B(n1962), .Z(n1968) );
  NANDN U2008 ( .A(n1912), .B(n42093), .Z(n1914) );
  XOR U2009 ( .A(n42134), .B(a[43]), .Z(n1953) );
  NANDN U2010 ( .A(n1953), .B(n42095), .Z(n1913) );
  NAND U2011 ( .A(n1914), .B(n1913), .Z(n1966) );
  NANDN U2012 ( .A(n1915), .B(n42231), .Z(n1917) );
  XOR U2013 ( .A(n165), .B(a[39]), .Z(n1956) );
  NANDN U2014 ( .A(n1956), .B(n42234), .Z(n1916) );
  AND U2015 ( .A(n1917), .B(n1916), .Z(n1965) );
  XNOR U2016 ( .A(n1966), .B(n1965), .Z(n1967) );
  XNOR U2017 ( .A(n1968), .B(n1967), .Z(n1972) );
  NANDN U2018 ( .A(n1919), .B(n1918), .Z(n1923) );
  NAND U2019 ( .A(n1921), .B(n1920), .Z(n1922) );
  AND U2020 ( .A(n1923), .B(n1922), .Z(n1971) );
  XOR U2021 ( .A(n1972), .B(n1971), .Z(n1973) );
  NANDN U2022 ( .A(n1925), .B(n1924), .Z(n1929) );
  NANDN U2023 ( .A(n1927), .B(n1926), .Z(n1928) );
  NAND U2024 ( .A(n1929), .B(n1928), .Z(n1974) );
  XOR U2025 ( .A(n1973), .B(n1974), .Z(n1941) );
  OR U2026 ( .A(n1931), .B(n1930), .Z(n1935) );
  NANDN U2027 ( .A(n1933), .B(n1932), .Z(n1934) );
  NAND U2028 ( .A(n1935), .B(n1934), .Z(n1942) );
  XNOR U2029 ( .A(n1941), .B(n1942), .Z(n1943) );
  XNOR U2030 ( .A(n1944), .B(n1943), .Z(n1977) );
  XNOR U2031 ( .A(n1977), .B(sreg[1061]), .Z(n1979) );
  NAND U2032 ( .A(n1936), .B(sreg[1060]), .Z(n1940) );
  OR U2033 ( .A(n1938), .B(n1937), .Z(n1939) );
  AND U2034 ( .A(n1940), .B(n1939), .Z(n1978) );
  XOR U2035 ( .A(n1979), .B(n1978), .Z(c[1061]) );
  NANDN U2036 ( .A(n1942), .B(n1941), .Z(n1946) );
  NAND U2037 ( .A(n1944), .B(n1943), .Z(n1945) );
  NAND U2038 ( .A(n1946), .B(n1945), .Z(n1985) );
  NAND U2039 ( .A(b[0]), .B(a[46]), .Z(n1947) );
  XNOR U2040 ( .A(b[1]), .B(n1947), .Z(n1949) );
  NAND U2041 ( .A(n21), .B(a[45]), .Z(n1948) );
  AND U2042 ( .A(n1949), .B(n1948), .Z(n2002) );
  XOR U2043 ( .A(a[42]), .B(n42197), .Z(n1991) );
  NANDN U2044 ( .A(n1991), .B(n42173), .Z(n1952) );
  NANDN U2045 ( .A(n1950), .B(n42172), .Z(n1951) );
  NAND U2046 ( .A(n1952), .B(n1951), .Z(n2000) );
  NAND U2047 ( .A(b[7]), .B(a[38]), .Z(n2001) );
  XNOR U2048 ( .A(n2000), .B(n2001), .Z(n2003) );
  XOR U2049 ( .A(n2002), .B(n2003), .Z(n2009) );
  NANDN U2050 ( .A(n1953), .B(n42093), .Z(n1955) );
  XOR U2051 ( .A(n42134), .B(a[44]), .Z(n1994) );
  NANDN U2052 ( .A(n1994), .B(n42095), .Z(n1954) );
  NAND U2053 ( .A(n1955), .B(n1954), .Z(n2007) );
  NANDN U2054 ( .A(n1956), .B(n42231), .Z(n1958) );
  XOR U2055 ( .A(n165), .B(a[40]), .Z(n1997) );
  NANDN U2056 ( .A(n1997), .B(n42234), .Z(n1957) );
  AND U2057 ( .A(n1958), .B(n1957), .Z(n2006) );
  XNOR U2058 ( .A(n2007), .B(n2006), .Z(n2008) );
  XNOR U2059 ( .A(n2009), .B(n2008), .Z(n2013) );
  NANDN U2060 ( .A(n1960), .B(n1959), .Z(n1964) );
  NAND U2061 ( .A(n1962), .B(n1961), .Z(n1963) );
  AND U2062 ( .A(n1964), .B(n1963), .Z(n2012) );
  XOR U2063 ( .A(n2013), .B(n2012), .Z(n2014) );
  NANDN U2064 ( .A(n1966), .B(n1965), .Z(n1970) );
  NANDN U2065 ( .A(n1968), .B(n1967), .Z(n1969) );
  NAND U2066 ( .A(n1970), .B(n1969), .Z(n2015) );
  XOR U2067 ( .A(n2014), .B(n2015), .Z(n1982) );
  OR U2068 ( .A(n1972), .B(n1971), .Z(n1976) );
  NANDN U2069 ( .A(n1974), .B(n1973), .Z(n1975) );
  NAND U2070 ( .A(n1976), .B(n1975), .Z(n1983) );
  XNOR U2071 ( .A(n1982), .B(n1983), .Z(n1984) );
  XNOR U2072 ( .A(n1985), .B(n1984), .Z(n2018) );
  XNOR U2073 ( .A(n2018), .B(sreg[1062]), .Z(n2020) );
  NAND U2074 ( .A(n1977), .B(sreg[1061]), .Z(n1981) );
  OR U2075 ( .A(n1979), .B(n1978), .Z(n1980) );
  AND U2076 ( .A(n1981), .B(n1980), .Z(n2019) );
  XOR U2077 ( .A(n2020), .B(n2019), .Z(c[1062]) );
  NANDN U2078 ( .A(n1983), .B(n1982), .Z(n1987) );
  NAND U2079 ( .A(n1985), .B(n1984), .Z(n1986) );
  NAND U2080 ( .A(n1987), .B(n1986), .Z(n2026) );
  NAND U2081 ( .A(b[0]), .B(a[47]), .Z(n1988) );
  XNOR U2082 ( .A(b[1]), .B(n1988), .Z(n1990) );
  NAND U2083 ( .A(n21), .B(a[46]), .Z(n1989) );
  AND U2084 ( .A(n1990), .B(n1989), .Z(n2043) );
  XOR U2085 ( .A(a[43]), .B(n42197), .Z(n2032) );
  NANDN U2086 ( .A(n2032), .B(n42173), .Z(n1993) );
  NANDN U2087 ( .A(n1991), .B(n42172), .Z(n1992) );
  NAND U2088 ( .A(n1993), .B(n1992), .Z(n2041) );
  NAND U2089 ( .A(b[7]), .B(a[39]), .Z(n2042) );
  XNOR U2090 ( .A(n2041), .B(n2042), .Z(n2044) );
  XOR U2091 ( .A(n2043), .B(n2044), .Z(n2050) );
  NANDN U2092 ( .A(n1994), .B(n42093), .Z(n1996) );
  XOR U2093 ( .A(n42134), .B(a[45]), .Z(n2035) );
  NANDN U2094 ( .A(n2035), .B(n42095), .Z(n1995) );
  NAND U2095 ( .A(n1996), .B(n1995), .Z(n2048) );
  NANDN U2096 ( .A(n1997), .B(n42231), .Z(n1999) );
  XOR U2097 ( .A(n165), .B(a[41]), .Z(n2038) );
  NANDN U2098 ( .A(n2038), .B(n42234), .Z(n1998) );
  AND U2099 ( .A(n1999), .B(n1998), .Z(n2047) );
  XNOR U2100 ( .A(n2048), .B(n2047), .Z(n2049) );
  XNOR U2101 ( .A(n2050), .B(n2049), .Z(n2054) );
  NANDN U2102 ( .A(n2001), .B(n2000), .Z(n2005) );
  NAND U2103 ( .A(n2003), .B(n2002), .Z(n2004) );
  AND U2104 ( .A(n2005), .B(n2004), .Z(n2053) );
  XOR U2105 ( .A(n2054), .B(n2053), .Z(n2055) );
  NANDN U2106 ( .A(n2007), .B(n2006), .Z(n2011) );
  NANDN U2107 ( .A(n2009), .B(n2008), .Z(n2010) );
  NAND U2108 ( .A(n2011), .B(n2010), .Z(n2056) );
  XOR U2109 ( .A(n2055), .B(n2056), .Z(n2023) );
  OR U2110 ( .A(n2013), .B(n2012), .Z(n2017) );
  NANDN U2111 ( .A(n2015), .B(n2014), .Z(n2016) );
  NAND U2112 ( .A(n2017), .B(n2016), .Z(n2024) );
  XNOR U2113 ( .A(n2023), .B(n2024), .Z(n2025) );
  XNOR U2114 ( .A(n2026), .B(n2025), .Z(n2059) );
  XNOR U2115 ( .A(n2059), .B(sreg[1063]), .Z(n2061) );
  NAND U2116 ( .A(n2018), .B(sreg[1062]), .Z(n2022) );
  OR U2117 ( .A(n2020), .B(n2019), .Z(n2021) );
  AND U2118 ( .A(n2022), .B(n2021), .Z(n2060) );
  XOR U2119 ( .A(n2061), .B(n2060), .Z(c[1063]) );
  NANDN U2120 ( .A(n2024), .B(n2023), .Z(n2028) );
  NAND U2121 ( .A(n2026), .B(n2025), .Z(n2027) );
  NAND U2122 ( .A(n2028), .B(n2027), .Z(n2067) );
  NAND U2123 ( .A(b[0]), .B(a[48]), .Z(n2029) );
  XNOR U2124 ( .A(b[1]), .B(n2029), .Z(n2031) );
  NAND U2125 ( .A(n21), .B(a[47]), .Z(n2030) );
  AND U2126 ( .A(n2031), .B(n2030), .Z(n2084) );
  XOR U2127 ( .A(a[44]), .B(n42197), .Z(n2073) );
  NANDN U2128 ( .A(n2073), .B(n42173), .Z(n2034) );
  NANDN U2129 ( .A(n2032), .B(n42172), .Z(n2033) );
  NAND U2130 ( .A(n2034), .B(n2033), .Z(n2082) );
  NAND U2131 ( .A(b[7]), .B(a[40]), .Z(n2083) );
  XNOR U2132 ( .A(n2082), .B(n2083), .Z(n2085) );
  XOR U2133 ( .A(n2084), .B(n2085), .Z(n2091) );
  NANDN U2134 ( .A(n2035), .B(n42093), .Z(n2037) );
  XOR U2135 ( .A(n42134), .B(a[46]), .Z(n2076) );
  NANDN U2136 ( .A(n2076), .B(n42095), .Z(n2036) );
  NAND U2137 ( .A(n2037), .B(n2036), .Z(n2089) );
  NANDN U2138 ( .A(n2038), .B(n42231), .Z(n2040) );
  XOR U2139 ( .A(n165), .B(a[42]), .Z(n2079) );
  NANDN U2140 ( .A(n2079), .B(n42234), .Z(n2039) );
  AND U2141 ( .A(n2040), .B(n2039), .Z(n2088) );
  XNOR U2142 ( .A(n2089), .B(n2088), .Z(n2090) );
  XNOR U2143 ( .A(n2091), .B(n2090), .Z(n2095) );
  NANDN U2144 ( .A(n2042), .B(n2041), .Z(n2046) );
  NAND U2145 ( .A(n2044), .B(n2043), .Z(n2045) );
  AND U2146 ( .A(n2046), .B(n2045), .Z(n2094) );
  XOR U2147 ( .A(n2095), .B(n2094), .Z(n2096) );
  NANDN U2148 ( .A(n2048), .B(n2047), .Z(n2052) );
  NANDN U2149 ( .A(n2050), .B(n2049), .Z(n2051) );
  NAND U2150 ( .A(n2052), .B(n2051), .Z(n2097) );
  XOR U2151 ( .A(n2096), .B(n2097), .Z(n2064) );
  OR U2152 ( .A(n2054), .B(n2053), .Z(n2058) );
  NANDN U2153 ( .A(n2056), .B(n2055), .Z(n2057) );
  NAND U2154 ( .A(n2058), .B(n2057), .Z(n2065) );
  XNOR U2155 ( .A(n2064), .B(n2065), .Z(n2066) );
  XNOR U2156 ( .A(n2067), .B(n2066), .Z(n2100) );
  XNOR U2157 ( .A(n2100), .B(sreg[1064]), .Z(n2102) );
  NAND U2158 ( .A(n2059), .B(sreg[1063]), .Z(n2063) );
  OR U2159 ( .A(n2061), .B(n2060), .Z(n2062) );
  AND U2160 ( .A(n2063), .B(n2062), .Z(n2101) );
  XOR U2161 ( .A(n2102), .B(n2101), .Z(c[1064]) );
  NANDN U2162 ( .A(n2065), .B(n2064), .Z(n2069) );
  NAND U2163 ( .A(n2067), .B(n2066), .Z(n2068) );
  NAND U2164 ( .A(n2069), .B(n2068), .Z(n2108) );
  NAND U2165 ( .A(b[0]), .B(a[49]), .Z(n2070) );
  XNOR U2166 ( .A(b[1]), .B(n2070), .Z(n2072) );
  NAND U2167 ( .A(n22), .B(a[48]), .Z(n2071) );
  AND U2168 ( .A(n2072), .B(n2071), .Z(n2125) );
  XOR U2169 ( .A(a[45]), .B(n42197), .Z(n2114) );
  NANDN U2170 ( .A(n2114), .B(n42173), .Z(n2075) );
  NANDN U2171 ( .A(n2073), .B(n42172), .Z(n2074) );
  NAND U2172 ( .A(n2075), .B(n2074), .Z(n2123) );
  NAND U2173 ( .A(b[7]), .B(a[41]), .Z(n2124) );
  XNOR U2174 ( .A(n2123), .B(n2124), .Z(n2126) );
  XOR U2175 ( .A(n2125), .B(n2126), .Z(n2132) );
  NANDN U2176 ( .A(n2076), .B(n42093), .Z(n2078) );
  XOR U2177 ( .A(n42134), .B(a[47]), .Z(n2117) );
  NANDN U2178 ( .A(n2117), .B(n42095), .Z(n2077) );
  NAND U2179 ( .A(n2078), .B(n2077), .Z(n2130) );
  NANDN U2180 ( .A(n2079), .B(n42231), .Z(n2081) );
  XOR U2181 ( .A(n165), .B(a[43]), .Z(n2120) );
  NANDN U2182 ( .A(n2120), .B(n42234), .Z(n2080) );
  AND U2183 ( .A(n2081), .B(n2080), .Z(n2129) );
  XNOR U2184 ( .A(n2130), .B(n2129), .Z(n2131) );
  XNOR U2185 ( .A(n2132), .B(n2131), .Z(n2136) );
  NANDN U2186 ( .A(n2083), .B(n2082), .Z(n2087) );
  NAND U2187 ( .A(n2085), .B(n2084), .Z(n2086) );
  AND U2188 ( .A(n2087), .B(n2086), .Z(n2135) );
  XOR U2189 ( .A(n2136), .B(n2135), .Z(n2137) );
  NANDN U2190 ( .A(n2089), .B(n2088), .Z(n2093) );
  NANDN U2191 ( .A(n2091), .B(n2090), .Z(n2092) );
  NAND U2192 ( .A(n2093), .B(n2092), .Z(n2138) );
  XOR U2193 ( .A(n2137), .B(n2138), .Z(n2105) );
  OR U2194 ( .A(n2095), .B(n2094), .Z(n2099) );
  NANDN U2195 ( .A(n2097), .B(n2096), .Z(n2098) );
  NAND U2196 ( .A(n2099), .B(n2098), .Z(n2106) );
  XNOR U2197 ( .A(n2105), .B(n2106), .Z(n2107) );
  XNOR U2198 ( .A(n2108), .B(n2107), .Z(n2141) );
  XNOR U2199 ( .A(n2141), .B(sreg[1065]), .Z(n2143) );
  NAND U2200 ( .A(n2100), .B(sreg[1064]), .Z(n2104) );
  OR U2201 ( .A(n2102), .B(n2101), .Z(n2103) );
  AND U2202 ( .A(n2104), .B(n2103), .Z(n2142) );
  XOR U2203 ( .A(n2143), .B(n2142), .Z(c[1065]) );
  NANDN U2204 ( .A(n2106), .B(n2105), .Z(n2110) );
  NAND U2205 ( .A(n2108), .B(n2107), .Z(n2109) );
  NAND U2206 ( .A(n2110), .B(n2109), .Z(n2149) );
  NAND U2207 ( .A(b[0]), .B(a[50]), .Z(n2111) );
  XNOR U2208 ( .A(b[1]), .B(n2111), .Z(n2113) );
  NAND U2209 ( .A(n22), .B(a[49]), .Z(n2112) );
  AND U2210 ( .A(n2113), .B(n2112), .Z(n2166) );
  XOR U2211 ( .A(a[46]), .B(n42197), .Z(n2155) );
  NANDN U2212 ( .A(n2155), .B(n42173), .Z(n2116) );
  NANDN U2213 ( .A(n2114), .B(n42172), .Z(n2115) );
  NAND U2214 ( .A(n2116), .B(n2115), .Z(n2164) );
  NAND U2215 ( .A(b[7]), .B(a[42]), .Z(n2165) );
  XNOR U2216 ( .A(n2164), .B(n2165), .Z(n2167) );
  XOR U2217 ( .A(n2166), .B(n2167), .Z(n2173) );
  NANDN U2218 ( .A(n2117), .B(n42093), .Z(n2119) );
  XOR U2219 ( .A(n42134), .B(a[48]), .Z(n2158) );
  NANDN U2220 ( .A(n2158), .B(n42095), .Z(n2118) );
  NAND U2221 ( .A(n2119), .B(n2118), .Z(n2171) );
  NANDN U2222 ( .A(n2120), .B(n42231), .Z(n2122) );
  XOR U2223 ( .A(n165), .B(a[44]), .Z(n2161) );
  NANDN U2224 ( .A(n2161), .B(n42234), .Z(n2121) );
  AND U2225 ( .A(n2122), .B(n2121), .Z(n2170) );
  XNOR U2226 ( .A(n2171), .B(n2170), .Z(n2172) );
  XNOR U2227 ( .A(n2173), .B(n2172), .Z(n2177) );
  NANDN U2228 ( .A(n2124), .B(n2123), .Z(n2128) );
  NAND U2229 ( .A(n2126), .B(n2125), .Z(n2127) );
  AND U2230 ( .A(n2128), .B(n2127), .Z(n2176) );
  XOR U2231 ( .A(n2177), .B(n2176), .Z(n2178) );
  NANDN U2232 ( .A(n2130), .B(n2129), .Z(n2134) );
  NANDN U2233 ( .A(n2132), .B(n2131), .Z(n2133) );
  NAND U2234 ( .A(n2134), .B(n2133), .Z(n2179) );
  XOR U2235 ( .A(n2178), .B(n2179), .Z(n2146) );
  OR U2236 ( .A(n2136), .B(n2135), .Z(n2140) );
  NANDN U2237 ( .A(n2138), .B(n2137), .Z(n2139) );
  NAND U2238 ( .A(n2140), .B(n2139), .Z(n2147) );
  XNOR U2239 ( .A(n2146), .B(n2147), .Z(n2148) );
  XNOR U2240 ( .A(n2149), .B(n2148), .Z(n2182) );
  XNOR U2241 ( .A(n2182), .B(sreg[1066]), .Z(n2184) );
  NAND U2242 ( .A(n2141), .B(sreg[1065]), .Z(n2145) );
  OR U2243 ( .A(n2143), .B(n2142), .Z(n2144) );
  AND U2244 ( .A(n2145), .B(n2144), .Z(n2183) );
  XOR U2245 ( .A(n2184), .B(n2183), .Z(c[1066]) );
  NANDN U2246 ( .A(n2147), .B(n2146), .Z(n2151) );
  NAND U2247 ( .A(n2149), .B(n2148), .Z(n2150) );
  NAND U2248 ( .A(n2151), .B(n2150), .Z(n2190) );
  NAND U2249 ( .A(b[0]), .B(a[51]), .Z(n2152) );
  XNOR U2250 ( .A(b[1]), .B(n2152), .Z(n2154) );
  NAND U2251 ( .A(n22), .B(a[50]), .Z(n2153) );
  AND U2252 ( .A(n2154), .B(n2153), .Z(n2207) );
  XOR U2253 ( .A(a[47]), .B(n42197), .Z(n2196) );
  NANDN U2254 ( .A(n2196), .B(n42173), .Z(n2157) );
  NANDN U2255 ( .A(n2155), .B(n42172), .Z(n2156) );
  NAND U2256 ( .A(n2157), .B(n2156), .Z(n2205) );
  NAND U2257 ( .A(b[7]), .B(a[43]), .Z(n2206) );
  XNOR U2258 ( .A(n2205), .B(n2206), .Z(n2208) );
  XOR U2259 ( .A(n2207), .B(n2208), .Z(n2214) );
  NANDN U2260 ( .A(n2158), .B(n42093), .Z(n2160) );
  XOR U2261 ( .A(n42134), .B(a[49]), .Z(n2199) );
  NANDN U2262 ( .A(n2199), .B(n42095), .Z(n2159) );
  NAND U2263 ( .A(n2160), .B(n2159), .Z(n2212) );
  NANDN U2264 ( .A(n2161), .B(n42231), .Z(n2163) );
  XOR U2265 ( .A(n165), .B(a[45]), .Z(n2202) );
  NANDN U2266 ( .A(n2202), .B(n42234), .Z(n2162) );
  AND U2267 ( .A(n2163), .B(n2162), .Z(n2211) );
  XNOR U2268 ( .A(n2212), .B(n2211), .Z(n2213) );
  XNOR U2269 ( .A(n2214), .B(n2213), .Z(n2218) );
  NANDN U2270 ( .A(n2165), .B(n2164), .Z(n2169) );
  NAND U2271 ( .A(n2167), .B(n2166), .Z(n2168) );
  AND U2272 ( .A(n2169), .B(n2168), .Z(n2217) );
  XOR U2273 ( .A(n2218), .B(n2217), .Z(n2219) );
  NANDN U2274 ( .A(n2171), .B(n2170), .Z(n2175) );
  NANDN U2275 ( .A(n2173), .B(n2172), .Z(n2174) );
  NAND U2276 ( .A(n2175), .B(n2174), .Z(n2220) );
  XOR U2277 ( .A(n2219), .B(n2220), .Z(n2187) );
  OR U2278 ( .A(n2177), .B(n2176), .Z(n2181) );
  NANDN U2279 ( .A(n2179), .B(n2178), .Z(n2180) );
  NAND U2280 ( .A(n2181), .B(n2180), .Z(n2188) );
  XNOR U2281 ( .A(n2187), .B(n2188), .Z(n2189) );
  XNOR U2282 ( .A(n2190), .B(n2189), .Z(n2223) );
  XNOR U2283 ( .A(n2223), .B(sreg[1067]), .Z(n2225) );
  NAND U2284 ( .A(n2182), .B(sreg[1066]), .Z(n2186) );
  OR U2285 ( .A(n2184), .B(n2183), .Z(n2185) );
  AND U2286 ( .A(n2186), .B(n2185), .Z(n2224) );
  XOR U2287 ( .A(n2225), .B(n2224), .Z(c[1067]) );
  NANDN U2288 ( .A(n2188), .B(n2187), .Z(n2192) );
  NAND U2289 ( .A(n2190), .B(n2189), .Z(n2191) );
  NAND U2290 ( .A(n2192), .B(n2191), .Z(n2231) );
  NAND U2291 ( .A(b[0]), .B(a[52]), .Z(n2193) );
  XNOR U2292 ( .A(b[1]), .B(n2193), .Z(n2195) );
  NAND U2293 ( .A(n22), .B(a[51]), .Z(n2194) );
  AND U2294 ( .A(n2195), .B(n2194), .Z(n2248) );
  XOR U2295 ( .A(a[48]), .B(n42197), .Z(n2237) );
  NANDN U2296 ( .A(n2237), .B(n42173), .Z(n2198) );
  NANDN U2297 ( .A(n2196), .B(n42172), .Z(n2197) );
  NAND U2298 ( .A(n2198), .B(n2197), .Z(n2246) );
  NAND U2299 ( .A(b[7]), .B(a[44]), .Z(n2247) );
  XNOR U2300 ( .A(n2246), .B(n2247), .Z(n2249) );
  XOR U2301 ( .A(n2248), .B(n2249), .Z(n2255) );
  NANDN U2302 ( .A(n2199), .B(n42093), .Z(n2201) );
  XOR U2303 ( .A(n42134), .B(a[50]), .Z(n2240) );
  NANDN U2304 ( .A(n2240), .B(n42095), .Z(n2200) );
  NAND U2305 ( .A(n2201), .B(n2200), .Z(n2253) );
  NANDN U2306 ( .A(n2202), .B(n42231), .Z(n2204) );
  XOR U2307 ( .A(n165), .B(a[46]), .Z(n2243) );
  NANDN U2308 ( .A(n2243), .B(n42234), .Z(n2203) );
  AND U2309 ( .A(n2204), .B(n2203), .Z(n2252) );
  XNOR U2310 ( .A(n2253), .B(n2252), .Z(n2254) );
  XNOR U2311 ( .A(n2255), .B(n2254), .Z(n2259) );
  NANDN U2312 ( .A(n2206), .B(n2205), .Z(n2210) );
  NAND U2313 ( .A(n2208), .B(n2207), .Z(n2209) );
  AND U2314 ( .A(n2210), .B(n2209), .Z(n2258) );
  XOR U2315 ( .A(n2259), .B(n2258), .Z(n2260) );
  NANDN U2316 ( .A(n2212), .B(n2211), .Z(n2216) );
  NANDN U2317 ( .A(n2214), .B(n2213), .Z(n2215) );
  NAND U2318 ( .A(n2216), .B(n2215), .Z(n2261) );
  XOR U2319 ( .A(n2260), .B(n2261), .Z(n2228) );
  OR U2320 ( .A(n2218), .B(n2217), .Z(n2222) );
  NANDN U2321 ( .A(n2220), .B(n2219), .Z(n2221) );
  NAND U2322 ( .A(n2222), .B(n2221), .Z(n2229) );
  XNOR U2323 ( .A(n2228), .B(n2229), .Z(n2230) );
  XNOR U2324 ( .A(n2231), .B(n2230), .Z(n2264) );
  XNOR U2325 ( .A(n2264), .B(sreg[1068]), .Z(n2266) );
  NAND U2326 ( .A(n2223), .B(sreg[1067]), .Z(n2227) );
  OR U2327 ( .A(n2225), .B(n2224), .Z(n2226) );
  AND U2328 ( .A(n2227), .B(n2226), .Z(n2265) );
  XOR U2329 ( .A(n2266), .B(n2265), .Z(c[1068]) );
  NANDN U2330 ( .A(n2229), .B(n2228), .Z(n2233) );
  NAND U2331 ( .A(n2231), .B(n2230), .Z(n2232) );
  NAND U2332 ( .A(n2233), .B(n2232), .Z(n2272) );
  NAND U2333 ( .A(b[0]), .B(a[53]), .Z(n2234) );
  XNOR U2334 ( .A(b[1]), .B(n2234), .Z(n2236) );
  NAND U2335 ( .A(n22), .B(a[52]), .Z(n2235) );
  AND U2336 ( .A(n2236), .B(n2235), .Z(n2289) );
  XOR U2337 ( .A(a[49]), .B(n42197), .Z(n2278) );
  NANDN U2338 ( .A(n2278), .B(n42173), .Z(n2239) );
  NANDN U2339 ( .A(n2237), .B(n42172), .Z(n2238) );
  NAND U2340 ( .A(n2239), .B(n2238), .Z(n2287) );
  NAND U2341 ( .A(b[7]), .B(a[45]), .Z(n2288) );
  XNOR U2342 ( .A(n2287), .B(n2288), .Z(n2290) );
  XOR U2343 ( .A(n2289), .B(n2290), .Z(n2296) );
  NANDN U2344 ( .A(n2240), .B(n42093), .Z(n2242) );
  XOR U2345 ( .A(n42134), .B(a[51]), .Z(n2281) );
  NANDN U2346 ( .A(n2281), .B(n42095), .Z(n2241) );
  NAND U2347 ( .A(n2242), .B(n2241), .Z(n2294) );
  NANDN U2348 ( .A(n2243), .B(n42231), .Z(n2245) );
  XOR U2349 ( .A(n166), .B(a[47]), .Z(n2284) );
  NANDN U2350 ( .A(n2284), .B(n42234), .Z(n2244) );
  AND U2351 ( .A(n2245), .B(n2244), .Z(n2293) );
  XNOR U2352 ( .A(n2294), .B(n2293), .Z(n2295) );
  XNOR U2353 ( .A(n2296), .B(n2295), .Z(n2300) );
  NANDN U2354 ( .A(n2247), .B(n2246), .Z(n2251) );
  NAND U2355 ( .A(n2249), .B(n2248), .Z(n2250) );
  AND U2356 ( .A(n2251), .B(n2250), .Z(n2299) );
  XOR U2357 ( .A(n2300), .B(n2299), .Z(n2301) );
  NANDN U2358 ( .A(n2253), .B(n2252), .Z(n2257) );
  NANDN U2359 ( .A(n2255), .B(n2254), .Z(n2256) );
  NAND U2360 ( .A(n2257), .B(n2256), .Z(n2302) );
  XOR U2361 ( .A(n2301), .B(n2302), .Z(n2269) );
  OR U2362 ( .A(n2259), .B(n2258), .Z(n2263) );
  NANDN U2363 ( .A(n2261), .B(n2260), .Z(n2262) );
  NAND U2364 ( .A(n2263), .B(n2262), .Z(n2270) );
  XNOR U2365 ( .A(n2269), .B(n2270), .Z(n2271) );
  XNOR U2366 ( .A(n2272), .B(n2271), .Z(n2305) );
  XNOR U2367 ( .A(n2305), .B(sreg[1069]), .Z(n2307) );
  NAND U2368 ( .A(n2264), .B(sreg[1068]), .Z(n2268) );
  OR U2369 ( .A(n2266), .B(n2265), .Z(n2267) );
  AND U2370 ( .A(n2268), .B(n2267), .Z(n2306) );
  XOR U2371 ( .A(n2307), .B(n2306), .Z(c[1069]) );
  NANDN U2372 ( .A(n2270), .B(n2269), .Z(n2274) );
  NAND U2373 ( .A(n2272), .B(n2271), .Z(n2273) );
  NAND U2374 ( .A(n2274), .B(n2273), .Z(n2313) );
  NAND U2375 ( .A(b[0]), .B(a[54]), .Z(n2275) );
  XNOR U2376 ( .A(b[1]), .B(n2275), .Z(n2277) );
  NAND U2377 ( .A(n22), .B(a[53]), .Z(n2276) );
  AND U2378 ( .A(n2277), .B(n2276), .Z(n2330) );
  XOR U2379 ( .A(a[50]), .B(n42197), .Z(n2319) );
  NANDN U2380 ( .A(n2319), .B(n42173), .Z(n2280) );
  NANDN U2381 ( .A(n2278), .B(n42172), .Z(n2279) );
  NAND U2382 ( .A(n2280), .B(n2279), .Z(n2328) );
  NAND U2383 ( .A(b[7]), .B(a[46]), .Z(n2329) );
  XNOR U2384 ( .A(n2328), .B(n2329), .Z(n2331) );
  XOR U2385 ( .A(n2330), .B(n2331), .Z(n2337) );
  NANDN U2386 ( .A(n2281), .B(n42093), .Z(n2283) );
  XOR U2387 ( .A(n42134), .B(a[52]), .Z(n2322) );
  NANDN U2388 ( .A(n2322), .B(n42095), .Z(n2282) );
  NAND U2389 ( .A(n2283), .B(n2282), .Z(n2335) );
  NANDN U2390 ( .A(n2284), .B(n42231), .Z(n2286) );
  XOR U2391 ( .A(n166), .B(a[48]), .Z(n2325) );
  NANDN U2392 ( .A(n2325), .B(n42234), .Z(n2285) );
  AND U2393 ( .A(n2286), .B(n2285), .Z(n2334) );
  XNOR U2394 ( .A(n2335), .B(n2334), .Z(n2336) );
  XNOR U2395 ( .A(n2337), .B(n2336), .Z(n2341) );
  NANDN U2396 ( .A(n2288), .B(n2287), .Z(n2292) );
  NAND U2397 ( .A(n2290), .B(n2289), .Z(n2291) );
  AND U2398 ( .A(n2292), .B(n2291), .Z(n2340) );
  XOR U2399 ( .A(n2341), .B(n2340), .Z(n2342) );
  NANDN U2400 ( .A(n2294), .B(n2293), .Z(n2298) );
  NANDN U2401 ( .A(n2296), .B(n2295), .Z(n2297) );
  NAND U2402 ( .A(n2298), .B(n2297), .Z(n2343) );
  XOR U2403 ( .A(n2342), .B(n2343), .Z(n2310) );
  OR U2404 ( .A(n2300), .B(n2299), .Z(n2304) );
  NANDN U2405 ( .A(n2302), .B(n2301), .Z(n2303) );
  NAND U2406 ( .A(n2304), .B(n2303), .Z(n2311) );
  XNOR U2407 ( .A(n2310), .B(n2311), .Z(n2312) );
  XNOR U2408 ( .A(n2313), .B(n2312), .Z(n2346) );
  XNOR U2409 ( .A(n2346), .B(sreg[1070]), .Z(n2348) );
  NAND U2410 ( .A(n2305), .B(sreg[1069]), .Z(n2309) );
  OR U2411 ( .A(n2307), .B(n2306), .Z(n2308) );
  AND U2412 ( .A(n2309), .B(n2308), .Z(n2347) );
  XOR U2413 ( .A(n2348), .B(n2347), .Z(c[1070]) );
  NANDN U2414 ( .A(n2311), .B(n2310), .Z(n2315) );
  NAND U2415 ( .A(n2313), .B(n2312), .Z(n2314) );
  NAND U2416 ( .A(n2315), .B(n2314), .Z(n2354) );
  NAND U2417 ( .A(b[0]), .B(a[55]), .Z(n2316) );
  XNOR U2418 ( .A(b[1]), .B(n2316), .Z(n2318) );
  NAND U2419 ( .A(n22), .B(a[54]), .Z(n2317) );
  AND U2420 ( .A(n2318), .B(n2317), .Z(n2371) );
  XOR U2421 ( .A(a[51]), .B(n42197), .Z(n2360) );
  NANDN U2422 ( .A(n2360), .B(n42173), .Z(n2321) );
  NANDN U2423 ( .A(n2319), .B(n42172), .Z(n2320) );
  NAND U2424 ( .A(n2321), .B(n2320), .Z(n2369) );
  NAND U2425 ( .A(b[7]), .B(a[47]), .Z(n2370) );
  XNOR U2426 ( .A(n2369), .B(n2370), .Z(n2372) );
  XOR U2427 ( .A(n2371), .B(n2372), .Z(n2378) );
  NANDN U2428 ( .A(n2322), .B(n42093), .Z(n2324) );
  XOR U2429 ( .A(n42134), .B(a[53]), .Z(n2363) );
  NANDN U2430 ( .A(n2363), .B(n42095), .Z(n2323) );
  NAND U2431 ( .A(n2324), .B(n2323), .Z(n2376) );
  NANDN U2432 ( .A(n2325), .B(n42231), .Z(n2327) );
  XOR U2433 ( .A(n166), .B(a[49]), .Z(n2366) );
  NANDN U2434 ( .A(n2366), .B(n42234), .Z(n2326) );
  AND U2435 ( .A(n2327), .B(n2326), .Z(n2375) );
  XNOR U2436 ( .A(n2376), .B(n2375), .Z(n2377) );
  XNOR U2437 ( .A(n2378), .B(n2377), .Z(n2382) );
  NANDN U2438 ( .A(n2329), .B(n2328), .Z(n2333) );
  NAND U2439 ( .A(n2331), .B(n2330), .Z(n2332) );
  AND U2440 ( .A(n2333), .B(n2332), .Z(n2381) );
  XOR U2441 ( .A(n2382), .B(n2381), .Z(n2383) );
  NANDN U2442 ( .A(n2335), .B(n2334), .Z(n2339) );
  NANDN U2443 ( .A(n2337), .B(n2336), .Z(n2338) );
  NAND U2444 ( .A(n2339), .B(n2338), .Z(n2384) );
  XOR U2445 ( .A(n2383), .B(n2384), .Z(n2351) );
  OR U2446 ( .A(n2341), .B(n2340), .Z(n2345) );
  NANDN U2447 ( .A(n2343), .B(n2342), .Z(n2344) );
  NAND U2448 ( .A(n2345), .B(n2344), .Z(n2352) );
  XNOR U2449 ( .A(n2351), .B(n2352), .Z(n2353) );
  XNOR U2450 ( .A(n2354), .B(n2353), .Z(n2387) );
  XNOR U2451 ( .A(n2387), .B(sreg[1071]), .Z(n2389) );
  NAND U2452 ( .A(n2346), .B(sreg[1070]), .Z(n2350) );
  OR U2453 ( .A(n2348), .B(n2347), .Z(n2349) );
  AND U2454 ( .A(n2350), .B(n2349), .Z(n2388) );
  XOR U2455 ( .A(n2389), .B(n2388), .Z(c[1071]) );
  NANDN U2456 ( .A(n2352), .B(n2351), .Z(n2356) );
  NAND U2457 ( .A(n2354), .B(n2353), .Z(n2355) );
  NAND U2458 ( .A(n2356), .B(n2355), .Z(n2395) );
  NAND U2459 ( .A(b[0]), .B(a[56]), .Z(n2357) );
  XNOR U2460 ( .A(b[1]), .B(n2357), .Z(n2359) );
  NAND U2461 ( .A(n23), .B(a[55]), .Z(n2358) );
  AND U2462 ( .A(n2359), .B(n2358), .Z(n2412) );
  XOR U2463 ( .A(a[52]), .B(n42197), .Z(n2401) );
  NANDN U2464 ( .A(n2401), .B(n42173), .Z(n2362) );
  NANDN U2465 ( .A(n2360), .B(n42172), .Z(n2361) );
  NAND U2466 ( .A(n2362), .B(n2361), .Z(n2410) );
  NAND U2467 ( .A(b[7]), .B(a[48]), .Z(n2411) );
  XNOR U2468 ( .A(n2410), .B(n2411), .Z(n2413) );
  XOR U2469 ( .A(n2412), .B(n2413), .Z(n2419) );
  NANDN U2470 ( .A(n2363), .B(n42093), .Z(n2365) );
  XOR U2471 ( .A(n42134), .B(a[54]), .Z(n2404) );
  NANDN U2472 ( .A(n2404), .B(n42095), .Z(n2364) );
  NAND U2473 ( .A(n2365), .B(n2364), .Z(n2417) );
  NANDN U2474 ( .A(n2366), .B(n42231), .Z(n2368) );
  XOR U2475 ( .A(n166), .B(a[50]), .Z(n2407) );
  NANDN U2476 ( .A(n2407), .B(n42234), .Z(n2367) );
  AND U2477 ( .A(n2368), .B(n2367), .Z(n2416) );
  XNOR U2478 ( .A(n2417), .B(n2416), .Z(n2418) );
  XNOR U2479 ( .A(n2419), .B(n2418), .Z(n2423) );
  NANDN U2480 ( .A(n2370), .B(n2369), .Z(n2374) );
  NAND U2481 ( .A(n2372), .B(n2371), .Z(n2373) );
  AND U2482 ( .A(n2374), .B(n2373), .Z(n2422) );
  XOR U2483 ( .A(n2423), .B(n2422), .Z(n2424) );
  NANDN U2484 ( .A(n2376), .B(n2375), .Z(n2380) );
  NANDN U2485 ( .A(n2378), .B(n2377), .Z(n2379) );
  NAND U2486 ( .A(n2380), .B(n2379), .Z(n2425) );
  XOR U2487 ( .A(n2424), .B(n2425), .Z(n2392) );
  OR U2488 ( .A(n2382), .B(n2381), .Z(n2386) );
  NANDN U2489 ( .A(n2384), .B(n2383), .Z(n2385) );
  NAND U2490 ( .A(n2386), .B(n2385), .Z(n2393) );
  XNOR U2491 ( .A(n2392), .B(n2393), .Z(n2394) );
  XNOR U2492 ( .A(n2395), .B(n2394), .Z(n2428) );
  XNOR U2493 ( .A(n2428), .B(sreg[1072]), .Z(n2430) );
  NAND U2494 ( .A(n2387), .B(sreg[1071]), .Z(n2391) );
  OR U2495 ( .A(n2389), .B(n2388), .Z(n2390) );
  AND U2496 ( .A(n2391), .B(n2390), .Z(n2429) );
  XOR U2497 ( .A(n2430), .B(n2429), .Z(c[1072]) );
  NANDN U2498 ( .A(n2393), .B(n2392), .Z(n2397) );
  NAND U2499 ( .A(n2395), .B(n2394), .Z(n2396) );
  NAND U2500 ( .A(n2397), .B(n2396), .Z(n2436) );
  NAND U2501 ( .A(b[0]), .B(a[57]), .Z(n2398) );
  XNOR U2502 ( .A(b[1]), .B(n2398), .Z(n2400) );
  NAND U2503 ( .A(n23), .B(a[56]), .Z(n2399) );
  AND U2504 ( .A(n2400), .B(n2399), .Z(n2453) );
  XOR U2505 ( .A(a[53]), .B(n42197), .Z(n2442) );
  NANDN U2506 ( .A(n2442), .B(n42173), .Z(n2403) );
  NANDN U2507 ( .A(n2401), .B(n42172), .Z(n2402) );
  NAND U2508 ( .A(n2403), .B(n2402), .Z(n2451) );
  NAND U2509 ( .A(b[7]), .B(a[49]), .Z(n2452) );
  XNOR U2510 ( .A(n2451), .B(n2452), .Z(n2454) );
  XOR U2511 ( .A(n2453), .B(n2454), .Z(n2460) );
  NANDN U2512 ( .A(n2404), .B(n42093), .Z(n2406) );
  XOR U2513 ( .A(n42134), .B(a[55]), .Z(n2445) );
  NANDN U2514 ( .A(n2445), .B(n42095), .Z(n2405) );
  NAND U2515 ( .A(n2406), .B(n2405), .Z(n2458) );
  NANDN U2516 ( .A(n2407), .B(n42231), .Z(n2409) );
  XOR U2517 ( .A(n166), .B(a[51]), .Z(n2448) );
  NANDN U2518 ( .A(n2448), .B(n42234), .Z(n2408) );
  AND U2519 ( .A(n2409), .B(n2408), .Z(n2457) );
  XNOR U2520 ( .A(n2458), .B(n2457), .Z(n2459) );
  XNOR U2521 ( .A(n2460), .B(n2459), .Z(n2464) );
  NANDN U2522 ( .A(n2411), .B(n2410), .Z(n2415) );
  NAND U2523 ( .A(n2413), .B(n2412), .Z(n2414) );
  AND U2524 ( .A(n2415), .B(n2414), .Z(n2463) );
  XOR U2525 ( .A(n2464), .B(n2463), .Z(n2465) );
  NANDN U2526 ( .A(n2417), .B(n2416), .Z(n2421) );
  NANDN U2527 ( .A(n2419), .B(n2418), .Z(n2420) );
  NAND U2528 ( .A(n2421), .B(n2420), .Z(n2466) );
  XOR U2529 ( .A(n2465), .B(n2466), .Z(n2433) );
  OR U2530 ( .A(n2423), .B(n2422), .Z(n2427) );
  NANDN U2531 ( .A(n2425), .B(n2424), .Z(n2426) );
  NAND U2532 ( .A(n2427), .B(n2426), .Z(n2434) );
  XNOR U2533 ( .A(n2433), .B(n2434), .Z(n2435) );
  XNOR U2534 ( .A(n2436), .B(n2435), .Z(n2469) );
  XNOR U2535 ( .A(n2469), .B(sreg[1073]), .Z(n2471) );
  NAND U2536 ( .A(n2428), .B(sreg[1072]), .Z(n2432) );
  OR U2537 ( .A(n2430), .B(n2429), .Z(n2431) );
  AND U2538 ( .A(n2432), .B(n2431), .Z(n2470) );
  XOR U2539 ( .A(n2471), .B(n2470), .Z(c[1073]) );
  NANDN U2540 ( .A(n2434), .B(n2433), .Z(n2438) );
  NAND U2541 ( .A(n2436), .B(n2435), .Z(n2437) );
  NAND U2542 ( .A(n2438), .B(n2437), .Z(n2477) );
  NAND U2543 ( .A(b[0]), .B(a[58]), .Z(n2439) );
  XNOR U2544 ( .A(b[1]), .B(n2439), .Z(n2441) );
  NAND U2545 ( .A(n23), .B(a[57]), .Z(n2440) );
  AND U2546 ( .A(n2441), .B(n2440), .Z(n2494) );
  XOR U2547 ( .A(a[54]), .B(n42197), .Z(n2483) );
  NANDN U2548 ( .A(n2483), .B(n42173), .Z(n2444) );
  NANDN U2549 ( .A(n2442), .B(n42172), .Z(n2443) );
  NAND U2550 ( .A(n2444), .B(n2443), .Z(n2492) );
  NAND U2551 ( .A(b[7]), .B(a[50]), .Z(n2493) );
  XNOR U2552 ( .A(n2492), .B(n2493), .Z(n2495) );
  XOR U2553 ( .A(n2494), .B(n2495), .Z(n2501) );
  NANDN U2554 ( .A(n2445), .B(n42093), .Z(n2447) );
  XOR U2555 ( .A(n42134), .B(a[56]), .Z(n2486) );
  NANDN U2556 ( .A(n2486), .B(n42095), .Z(n2446) );
  NAND U2557 ( .A(n2447), .B(n2446), .Z(n2499) );
  NANDN U2558 ( .A(n2448), .B(n42231), .Z(n2450) );
  XOR U2559 ( .A(n166), .B(a[52]), .Z(n2489) );
  NANDN U2560 ( .A(n2489), .B(n42234), .Z(n2449) );
  AND U2561 ( .A(n2450), .B(n2449), .Z(n2498) );
  XNOR U2562 ( .A(n2499), .B(n2498), .Z(n2500) );
  XNOR U2563 ( .A(n2501), .B(n2500), .Z(n2505) );
  NANDN U2564 ( .A(n2452), .B(n2451), .Z(n2456) );
  NAND U2565 ( .A(n2454), .B(n2453), .Z(n2455) );
  AND U2566 ( .A(n2456), .B(n2455), .Z(n2504) );
  XOR U2567 ( .A(n2505), .B(n2504), .Z(n2506) );
  NANDN U2568 ( .A(n2458), .B(n2457), .Z(n2462) );
  NANDN U2569 ( .A(n2460), .B(n2459), .Z(n2461) );
  NAND U2570 ( .A(n2462), .B(n2461), .Z(n2507) );
  XOR U2571 ( .A(n2506), .B(n2507), .Z(n2474) );
  OR U2572 ( .A(n2464), .B(n2463), .Z(n2468) );
  NANDN U2573 ( .A(n2466), .B(n2465), .Z(n2467) );
  NAND U2574 ( .A(n2468), .B(n2467), .Z(n2475) );
  XNOR U2575 ( .A(n2474), .B(n2475), .Z(n2476) );
  XNOR U2576 ( .A(n2477), .B(n2476), .Z(n2510) );
  XNOR U2577 ( .A(n2510), .B(sreg[1074]), .Z(n2512) );
  NAND U2578 ( .A(n2469), .B(sreg[1073]), .Z(n2473) );
  OR U2579 ( .A(n2471), .B(n2470), .Z(n2472) );
  AND U2580 ( .A(n2473), .B(n2472), .Z(n2511) );
  XOR U2581 ( .A(n2512), .B(n2511), .Z(c[1074]) );
  NANDN U2582 ( .A(n2475), .B(n2474), .Z(n2479) );
  NAND U2583 ( .A(n2477), .B(n2476), .Z(n2478) );
  NAND U2584 ( .A(n2479), .B(n2478), .Z(n2518) );
  NAND U2585 ( .A(b[0]), .B(a[59]), .Z(n2480) );
  XNOR U2586 ( .A(b[1]), .B(n2480), .Z(n2482) );
  NAND U2587 ( .A(n23), .B(a[58]), .Z(n2481) );
  AND U2588 ( .A(n2482), .B(n2481), .Z(n2535) );
  XOR U2589 ( .A(a[55]), .B(n42197), .Z(n2524) );
  NANDN U2590 ( .A(n2524), .B(n42173), .Z(n2485) );
  NANDN U2591 ( .A(n2483), .B(n42172), .Z(n2484) );
  NAND U2592 ( .A(n2485), .B(n2484), .Z(n2533) );
  NAND U2593 ( .A(b[7]), .B(a[51]), .Z(n2534) );
  XNOR U2594 ( .A(n2533), .B(n2534), .Z(n2536) );
  XOR U2595 ( .A(n2535), .B(n2536), .Z(n2542) );
  NANDN U2596 ( .A(n2486), .B(n42093), .Z(n2488) );
  XOR U2597 ( .A(n42134), .B(a[57]), .Z(n2527) );
  NANDN U2598 ( .A(n2527), .B(n42095), .Z(n2487) );
  NAND U2599 ( .A(n2488), .B(n2487), .Z(n2540) );
  NANDN U2600 ( .A(n2489), .B(n42231), .Z(n2491) );
  XOR U2601 ( .A(n166), .B(a[53]), .Z(n2530) );
  NANDN U2602 ( .A(n2530), .B(n42234), .Z(n2490) );
  AND U2603 ( .A(n2491), .B(n2490), .Z(n2539) );
  XNOR U2604 ( .A(n2540), .B(n2539), .Z(n2541) );
  XNOR U2605 ( .A(n2542), .B(n2541), .Z(n2546) );
  NANDN U2606 ( .A(n2493), .B(n2492), .Z(n2497) );
  NAND U2607 ( .A(n2495), .B(n2494), .Z(n2496) );
  AND U2608 ( .A(n2497), .B(n2496), .Z(n2545) );
  XOR U2609 ( .A(n2546), .B(n2545), .Z(n2547) );
  NANDN U2610 ( .A(n2499), .B(n2498), .Z(n2503) );
  NANDN U2611 ( .A(n2501), .B(n2500), .Z(n2502) );
  NAND U2612 ( .A(n2503), .B(n2502), .Z(n2548) );
  XOR U2613 ( .A(n2547), .B(n2548), .Z(n2515) );
  OR U2614 ( .A(n2505), .B(n2504), .Z(n2509) );
  NANDN U2615 ( .A(n2507), .B(n2506), .Z(n2508) );
  NAND U2616 ( .A(n2509), .B(n2508), .Z(n2516) );
  XNOR U2617 ( .A(n2515), .B(n2516), .Z(n2517) );
  XNOR U2618 ( .A(n2518), .B(n2517), .Z(n2551) );
  XNOR U2619 ( .A(n2551), .B(sreg[1075]), .Z(n2553) );
  NAND U2620 ( .A(n2510), .B(sreg[1074]), .Z(n2514) );
  OR U2621 ( .A(n2512), .B(n2511), .Z(n2513) );
  AND U2622 ( .A(n2514), .B(n2513), .Z(n2552) );
  XOR U2623 ( .A(n2553), .B(n2552), .Z(c[1075]) );
  NANDN U2624 ( .A(n2516), .B(n2515), .Z(n2520) );
  NAND U2625 ( .A(n2518), .B(n2517), .Z(n2519) );
  NAND U2626 ( .A(n2520), .B(n2519), .Z(n2559) );
  NAND U2627 ( .A(b[0]), .B(a[60]), .Z(n2521) );
  XNOR U2628 ( .A(b[1]), .B(n2521), .Z(n2523) );
  NAND U2629 ( .A(n23), .B(a[59]), .Z(n2522) );
  AND U2630 ( .A(n2523), .B(n2522), .Z(n2576) );
  XOR U2631 ( .A(a[56]), .B(n42197), .Z(n2565) );
  NANDN U2632 ( .A(n2565), .B(n42173), .Z(n2526) );
  NANDN U2633 ( .A(n2524), .B(n42172), .Z(n2525) );
  NAND U2634 ( .A(n2526), .B(n2525), .Z(n2574) );
  NAND U2635 ( .A(b[7]), .B(a[52]), .Z(n2575) );
  XNOR U2636 ( .A(n2574), .B(n2575), .Z(n2577) );
  XOR U2637 ( .A(n2576), .B(n2577), .Z(n2583) );
  NANDN U2638 ( .A(n2527), .B(n42093), .Z(n2529) );
  XOR U2639 ( .A(n42134), .B(a[58]), .Z(n2568) );
  NANDN U2640 ( .A(n2568), .B(n42095), .Z(n2528) );
  NAND U2641 ( .A(n2529), .B(n2528), .Z(n2581) );
  NANDN U2642 ( .A(n2530), .B(n42231), .Z(n2532) );
  XOR U2643 ( .A(n166), .B(a[54]), .Z(n2571) );
  NANDN U2644 ( .A(n2571), .B(n42234), .Z(n2531) );
  AND U2645 ( .A(n2532), .B(n2531), .Z(n2580) );
  XNOR U2646 ( .A(n2581), .B(n2580), .Z(n2582) );
  XNOR U2647 ( .A(n2583), .B(n2582), .Z(n2587) );
  NANDN U2648 ( .A(n2534), .B(n2533), .Z(n2538) );
  NAND U2649 ( .A(n2536), .B(n2535), .Z(n2537) );
  AND U2650 ( .A(n2538), .B(n2537), .Z(n2586) );
  XOR U2651 ( .A(n2587), .B(n2586), .Z(n2588) );
  NANDN U2652 ( .A(n2540), .B(n2539), .Z(n2544) );
  NANDN U2653 ( .A(n2542), .B(n2541), .Z(n2543) );
  NAND U2654 ( .A(n2544), .B(n2543), .Z(n2589) );
  XOR U2655 ( .A(n2588), .B(n2589), .Z(n2556) );
  OR U2656 ( .A(n2546), .B(n2545), .Z(n2550) );
  NANDN U2657 ( .A(n2548), .B(n2547), .Z(n2549) );
  NAND U2658 ( .A(n2550), .B(n2549), .Z(n2557) );
  XNOR U2659 ( .A(n2556), .B(n2557), .Z(n2558) );
  XNOR U2660 ( .A(n2559), .B(n2558), .Z(n2592) );
  XNOR U2661 ( .A(n2592), .B(sreg[1076]), .Z(n2594) );
  NAND U2662 ( .A(n2551), .B(sreg[1075]), .Z(n2555) );
  OR U2663 ( .A(n2553), .B(n2552), .Z(n2554) );
  AND U2664 ( .A(n2555), .B(n2554), .Z(n2593) );
  XOR U2665 ( .A(n2594), .B(n2593), .Z(c[1076]) );
  NANDN U2666 ( .A(n2557), .B(n2556), .Z(n2561) );
  NAND U2667 ( .A(n2559), .B(n2558), .Z(n2560) );
  NAND U2668 ( .A(n2561), .B(n2560), .Z(n2600) );
  NAND U2669 ( .A(b[0]), .B(a[61]), .Z(n2562) );
  XNOR U2670 ( .A(b[1]), .B(n2562), .Z(n2564) );
  NAND U2671 ( .A(n23), .B(a[60]), .Z(n2563) );
  AND U2672 ( .A(n2564), .B(n2563), .Z(n2617) );
  XOR U2673 ( .A(a[57]), .B(n42197), .Z(n2606) );
  NANDN U2674 ( .A(n2606), .B(n42173), .Z(n2567) );
  NANDN U2675 ( .A(n2565), .B(n42172), .Z(n2566) );
  NAND U2676 ( .A(n2567), .B(n2566), .Z(n2615) );
  NAND U2677 ( .A(b[7]), .B(a[53]), .Z(n2616) );
  XNOR U2678 ( .A(n2615), .B(n2616), .Z(n2618) );
  XOR U2679 ( .A(n2617), .B(n2618), .Z(n2624) );
  NANDN U2680 ( .A(n2568), .B(n42093), .Z(n2570) );
  XOR U2681 ( .A(n42134), .B(a[59]), .Z(n2609) );
  NANDN U2682 ( .A(n2609), .B(n42095), .Z(n2569) );
  NAND U2683 ( .A(n2570), .B(n2569), .Z(n2622) );
  NANDN U2684 ( .A(n2571), .B(n42231), .Z(n2573) );
  XOR U2685 ( .A(n166), .B(a[55]), .Z(n2612) );
  NANDN U2686 ( .A(n2612), .B(n42234), .Z(n2572) );
  AND U2687 ( .A(n2573), .B(n2572), .Z(n2621) );
  XNOR U2688 ( .A(n2622), .B(n2621), .Z(n2623) );
  XNOR U2689 ( .A(n2624), .B(n2623), .Z(n2628) );
  NANDN U2690 ( .A(n2575), .B(n2574), .Z(n2579) );
  NAND U2691 ( .A(n2577), .B(n2576), .Z(n2578) );
  AND U2692 ( .A(n2579), .B(n2578), .Z(n2627) );
  XOR U2693 ( .A(n2628), .B(n2627), .Z(n2629) );
  NANDN U2694 ( .A(n2581), .B(n2580), .Z(n2585) );
  NANDN U2695 ( .A(n2583), .B(n2582), .Z(n2584) );
  NAND U2696 ( .A(n2585), .B(n2584), .Z(n2630) );
  XOR U2697 ( .A(n2629), .B(n2630), .Z(n2597) );
  OR U2698 ( .A(n2587), .B(n2586), .Z(n2591) );
  NANDN U2699 ( .A(n2589), .B(n2588), .Z(n2590) );
  NAND U2700 ( .A(n2591), .B(n2590), .Z(n2598) );
  XNOR U2701 ( .A(n2597), .B(n2598), .Z(n2599) );
  XNOR U2702 ( .A(n2600), .B(n2599), .Z(n2633) );
  XNOR U2703 ( .A(n2633), .B(sreg[1077]), .Z(n2635) );
  NAND U2704 ( .A(n2592), .B(sreg[1076]), .Z(n2596) );
  OR U2705 ( .A(n2594), .B(n2593), .Z(n2595) );
  AND U2706 ( .A(n2596), .B(n2595), .Z(n2634) );
  XOR U2707 ( .A(n2635), .B(n2634), .Z(c[1077]) );
  NANDN U2708 ( .A(n2598), .B(n2597), .Z(n2602) );
  NAND U2709 ( .A(n2600), .B(n2599), .Z(n2601) );
  NAND U2710 ( .A(n2602), .B(n2601), .Z(n2641) );
  NAND U2711 ( .A(b[0]), .B(a[62]), .Z(n2603) );
  XNOR U2712 ( .A(b[1]), .B(n2603), .Z(n2605) );
  NAND U2713 ( .A(n23), .B(a[61]), .Z(n2604) );
  AND U2714 ( .A(n2605), .B(n2604), .Z(n2658) );
  XOR U2715 ( .A(a[58]), .B(n42197), .Z(n2647) );
  NANDN U2716 ( .A(n2647), .B(n42173), .Z(n2608) );
  NANDN U2717 ( .A(n2606), .B(n42172), .Z(n2607) );
  NAND U2718 ( .A(n2608), .B(n2607), .Z(n2656) );
  NAND U2719 ( .A(b[7]), .B(a[54]), .Z(n2657) );
  XNOR U2720 ( .A(n2656), .B(n2657), .Z(n2659) );
  XOR U2721 ( .A(n2658), .B(n2659), .Z(n2665) );
  NANDN U2722 ( .A(n2609), .B(n42093), .Z(n2611) );
  XOR U2723 ( .A(n42134), .B(a[60]), .Z(n2650) );
  NANDN U2724 ( .A(n2650), .B(n42095), .Z(n2610) );
  NAND U2725 ( .A(n2611), .B(n2610), .Z(n2663) );
  NANDN U2726 ( .A(n2612), .B(n42231), .Z(n2614) );
  XOR U2727 ( .A(n166), .B(a[56]), .Z(n2653) );
  NANDN U2728 ( .A(n2653), .B(n42234), .Z(n2613) );
  AND U2729 ( .A(n2614), .B(n2613), .Z(n2662) );
  XNOR U2730 ( .A(n2663), .B(n2662), .Z(n2664) );
  XNOR U2731 ( .A(n2665), .B(n2664), .Z(n2669) );
  NANDN U2732 ( .A(n2616), .B(n2615), .Z(n2620) );
  NAND U2733 ( .A(n2618), .B(n2617), .Z(n2619) );
  AND U2734 ( .A(n2620), .B(n2619), .Z(n2668) );
  XOR U2735 ( .A(n2669), .B(n2668), .Z(n2670) );
  NANDN U2736 ( .A(n2622), .B(n2621), .Z(n2626) );
  NANDN U2737 ( .A(n2624), .B(n2623), .Z(n2625) );
  NAND U2738 ( .A(n2626), .B(n2625), .Z(n2671) );
  XOR U2739 ( .A(n2670), .B(n2671), .Z(n2638) );
  OR U2740 ( .A(n2628), .B(n2627), .Z(n2632) );
  NANDN U2741 ( .A(n2630), .B(n2629), .Z(n2631) );
  NAND U2742 ( .A(n2632), .B(n2631), .Z(n2639) );
  XNOR U2743 ( .A(n2638), .B(n2639), .Z(n2640) );
  XNOR U2744 ( .A(n2641), .B(n2640), .Z(n2674) );
  XNOR U2745 ( .A(n2674), .B(sreg[1078]), .Z(n2676) );
  NAND U2746 ( .A(n2633), .B(sreg[1077]), .Z(n2637) );
  OR U2747 ( .A(n2635), .B(n2634), .Z(n2636) );
  AND U2748 ( .A(n2637), .B(n2636), .Z(n2675) );
  XOR U2749 ( .A(n2676), .B(n2675), .Z(c[1078]) );
  NANDN U2750 ( .A(n2639), .B(n2638), .Z(n2643) );
  NAND U2751 ( .A(n2641), .B(n2640), .Z(n2642) );
  NAND U2752 ( .A(n2643), .B(n2642), .Z(n2682) );
  NAND U2753 ( .A(b[0]), .B(a[63]), .Z(n2644) );
  XNOR U2754 ( .A(b[1]), .B(n2644), .Z(n2646) );
  NAND U2755 ( .A(n24), .B(a[62]), .Z(n2645) );
  AND U2756 ( .A(n2646), .B(n2645), .Z(n2699) );
  XOR U2757 ( .A(a[59]), .B(n42197), .Z(n2688) );
  NANDN U2758 ( .A(n2688), .B(n42173), .Z(n2649) );
  NANDN U2759 ( .A(n2647), .B(n42172), .Z(n2648) );
  NAND U2760 ( .A(n2649), .B(n2648), .Z(n2697) );
  NAND U2761 ( .A(b[7]), .B(a[55]), .Z(n2698) );
  XNOR U2762 ( .A(n2697), .B(n2698), .Z(n2700) );
  XOR U2763 ( .A(n2699), .B(n2700), .Z(n2706) );
  NANDN U2764 ( .A(n2650), .B(n42093), .Z(n2652) );
  XOR U2765 ( .A(n42134), .B(a[61]), .Z(n2691) );
  NANDN U2766 ( .A(n2691), .B(n42095), .Z(n2651) );
  NAND U2767 ( .A(n2652), .B(n2651), .Z(n2704) );
  NANDN U2768 ( .A(n2653), .B(n42231), .Z(n2655) );
  XOR U2769 ( .A(n166), .B(a[57]), .Z(n2694) );
  NANDN U2770 ( .A(n2694), .B(n42234), .Z(n2654) );
  AND U2771 ( .A(n2655), .B(n2654), .Z(n2703) );
  XNOR U2772 ( .A(n2704), .B(n2703), .Z(n2705) );
  XNOR U2773 ( .A(n2706), .B(n2705), .Z(n2710) );
  NANDN U2774 ( .A(n2657), .B(n2656), .Z(n2661) );
  NAND U2775 ( .A(n2659), .B(n2658), .Z(n2660) );
  AND U2776 ( .A(n2661), .B(n2660), .Z(n2709) );
  XOR U2777 ( .A(n2710), .B(n2709), .Z(n2711) );
  NANDN U2778 ( .A(n2663), .B(n2662), .Z(n2667) );
  NANDN U2779 ( .A(n2665), .B(n2664), .Z(n2666) );
  NAND U2780 ( .A(n2667), .B(n2666), .Z(n2712) );
  XOR U2781 ( .A(n2711), .B(n2712), .Z(n2679) );
  OR U2782 ( .A(n2669), .B(n2668), .Z(n2673) );
  NANDN U2783 ( .A(n2671), .B(n2670), .Z(n2672) );
  NAND U2784 ( .A(n2673), .B(n2672), .Z(n2680) );
  XNOR U2785 ( .A(n2679), .B(n2680), .Z(n2681) );
  XNOR U2786 ( .A(n2682), .B(n2681), .Z(n2715) );
  XNOR U2787 ( .A(n2715), .B(sreg[1079]), .Z(n2717) );
  NAND U2788 ( .A(n2674), .B(sreg[1078]), .Z(n2678) );
  OR U2789 ( .A(n2676), .B(n2675), .Z(n2677) );
  AND U2790 ( .A(n2678), .B(n2677), .Z(n2716) );
  XOR U2791 ( .A(n2717), .B(n2716), .Z(c[1079]) );
  NANDN U2792 ( .A(n2680), .B(n2679), .Z(n2684) );
  NAND U2793 ( .A(n2682), .B(n2681), .Z(n2683) );
  NAND U2794 ( .A(n2684), .B(n2683), .Z(n2723) );
  NAND U2795 ( .A(b[0]), .B(a[64]), .Z(n2685) );
  XNOR U2796 ( .A(b[1]), .B(n2685), .Z(n2687) );
  NAND U2797 ( .A(n24), .B(a[63]), .Z(n2686) );
  AND U2798 ( .A(n2687), .B(n2686), .Z(n2740) );
  XOR U2799 ( .A(a[60]), .B(n42197), .Z(n2729) );
  NANDN U2800 ( .A(n2729), .B(n42173), .Z(n2690) );
  NANDN U2801 ( .A(n2688), .B(n42172), .Z(n2689) );
  NAND U2802 ( .A(n2690), .B(n2689), .Z(n2738) );
  NAND U2803 ( .A(b[7]), .B(a[56]), .Z(n2739) );
  XNOR U2804 ( .A(n2738), .B(n2739), .Z(n2741) );
  XOR U2805 ( .A(n2740), .B(n2741), .Z(n2747) );
  NANDN U2806 ( .A(n2691), .B(n42093), .Z(n2693) );
  XOR U2807 ( .A(n42134), .B(a[62]), .Z(n2732) );
  NANDN U2808 ( .A(n2732), .B(n42095), .Z(n2692) );
  NAND U2809 ( .A(n2693), .B(n2692), .Z(n2745) );
  NANDN U2810 ( .A(n2694), .B(n42231), .Z(n2696) );
  XOR U2811 ( .A(n166), .B(a[58]), .Z(n2735) );
  NANDN U2812 ( .A(n2735), .B(n42234), .Z(n2695) );
  AND U2813 ( .A(n2696), .B(n2695), .Z(n2744) );
  XNOR U2814 ( .A(n2745), .B(n2744), .Z(n2746) );
  XNOR U2815 ( .A(n2747), .B(n2746), .Z(n2751) );
  NANDN U2816 ( .A(n2698), .B(n2697), .Z(n2702) );
  NAND U2817 ( .A(n2700), .B(n2699), .Z(n2701) );
  AND U2818 ( .A(n2702), .B(n2701), .Z(n2750) );
  XOR U2819 ( .A(n2751), .B(n2750), .Z(n2752) );
  NANDN U2820 ( .A(n2704), .B(n2703), .Z(n2708) );
  NANDN U2821 ( .A(n2706), .B(n2705), .Z(n2707) );
  NAND U2822 ( .A(n2708), .B(n2707), .Z(n2753) );
  XOR U2823 ( .A(n2752), .B(n2753), .Z(n2720) );
  OR U2824 ( .A(n2710), .B(n2709), .Z(n2714) );
  NANDN U2825 ( .A(n2712), .B(n2711), .Z(n2713) );
  NAND U2826 ( .A(n2714), .B(n2713), .Z(n2721) );
  XNOR U2827 ( .A(n2720), .B(n2721), .Z(n2722) );
  XNOR U2828 ( .A(n2723), .B(n2722), .Z(n2756) );
  XNOR U2829 ( .A(n2756), .B(sreg[1080]), .Z(n2758) );
  NAND U2830 ( .A(n2715), .B(sreg[1079]), .Z(n2719) );
  OR U2831 ( .A(n2717), .B(n2716), .Z(n2718) );
  AND U2832 ( .A(n2719), .B(n2718), .Z(n2757) );
  XOR U2833 ( .A(n2758), .B(n2757), .Z(c[1080]) );
  NANDN U2834 ( .A(n2721), .B(n2720), .Z(n2725) );
  NAND U2835 ( .A(n2723), .B(n2722), .Z(n2724) );
  NAND U2836 ( .A(n2725), .B(n2724), .Z(n2764) );
  NAND U2837 ( .A(b[0]), .B(a[65]), .Z(n2726) );
  XNOR U2838 ( .A(b[1]), .B(n2726), .Z(n2728) );
  NAND U2839 ( .A(n24), .B(a[64]), .Z(n2727) );
  AND U2840 ( .A(n2728), .B(n2727), .Z(n2781) );
  XOR U2841 ( .A(a[61]), .B(n42197), .Z(n2770) );
  NANDN U2842 ( .A(n2770), .B(n42173), .Z(n2731) );
  NANDN U2843 ( .A(n2729), .B(n42172), .Z(n2730) );
  NAND U2844 ( .A(n2731), .B(n2730), .Z(n2779) );
  NAND U2845 ( .A(b[7]), .B(a[57]), .Z(n2780) );
  XNOR U2846 ( .A(n2779), .B(n2780), .Z(n2782) );
  XOR U2847 ( .A(n2781), .B(n2782), .Z(n2788) );
  NANDN U2848 ( .A(n2732), .B(n42093), .Z(n2734) );
  XOR U2849 ( .A(n42134), .B(a[63]), .Z(n2773) );
  NANDN U2850 ( .A(n2773), .B(n42095), .Z(n2733) );
  NAND U2851 ( .A(n2734), .B(n2733), .Z(n2786) );
  NANDN U2852 ( .A(n2735), .B(n42231), .Z(n2737) );
  XOR U2853 ( .A(n167), .B(a[59]), .Z(n2776) );
  NANDN U2854 ( .A(n2776), .B(n42234), .Z(n2736) );
  AND U2855 ( .A(n2737), .B(n2736), .Z(n2785) );
  XNOR U2856 ( .A(n2786), .B(n2785), .Z(n2787) );
  XNOR U2857 ( .A(n2788), .B(n2787), .Z(n2792) );
  NANDN U2858 ( .A(n2739), .B(n2738), .Z(n2743) );
  NAND U2859 ( .A(n2741), .B(n2740), .Z(n2742) );
  AND U2860 ( .A(n2743), .B(n2742), .Z(n2791) );
  XOR U2861 ( .A(n2792), .B(n2791), .Z(n2793) );
  NANDN U2862 ( .A(n2745), .B(n2744), .Z(n2749) );
  NANDN U2863 ( .A(n2747), .B(n2746), .Z(n2748) );
  NAND U2864 ( .A(n2749), .B(n2748), .Z(n2794) );
  XOR U2865 ( .A(n2793), .B(n2794), .Z(n2761) );
  OR U2866 ( .A(n2751), .B(n2750), .Z(n2755) );
  NANDN U2867 ( .A(n2753), .B(n2752), .Z(n2754) );
  NAND U2868 ( .A(n2755), .B(n2754), .Z(n2762) );
  XNOR U2869 ( .A(n2761), .B(n2762), .Z(n2763) );
  XNOR U2870 ( .A(n2764), .B(n2763), .Z(n2797) );
  XNOR U2871 ( .A(n2797), .B(sreg[1081]), .Z(n2799) );
  NAND U2872 ( .A(n2756), .B(sreg[1080]), .Z(n2760) );
  OR U2873 ( .A(n2758), .B(n2757), .Z(n2759) );
  AND U2874 ( .A(n2760), .B(n2759), .Z(n2798) );
  XOR U2875 ( .A(n2799), .B(n2798), .Z(c[1081]) );
  NANDN U2876 ( .A(n2762), .B(n2761), .Z(n2766) );
  NAND U2877 ( .A(n2764), .B(n2763), .Z(n2765) );
  NAND U2878 ( .A(n2766), .B(n2765), .Z(n2805) );
  NAND U2879 ( .A(b[0]), .B(a[66]), .Z(n2767) );
  XNOR U2880 ( .A(b[1]), .B(n2767), .Z(n2769) );
  NAND U2881 ( .A(n24), .B(a[65]), .Z(n2768) );
  AND U2882 ( .A(n2769), .B(n2768), .Z(n2822) );
  XOR U2883 ( .A(a[62]), .B(n42197), .Z(n2811) );
  NANDN U2884 ( .A(n2811), .B(n42173), .Z(n2772) );
  NANDN U2885 ( .A(n2770), .B(n42172), .Z(n2771) );
  NAND U2886 ( .A(n2772), .B(n2771), .Z(n2820) );
  NAND U2887 ( .A(b[7]), .B(a[58]), .Z(n2821) );
  XNOR U2888 ( .A(n2820), .B(n2821), .Z(n2823) );
  XOR U2889 ( .A(n2822), .B(n2823), .Z(n2829) );
  NANDN U2890 ( .A(n2773), .B(n42093), .Z(n2775) );
  XOR U2891 ( .A(n42134), .B(a[64]), .Z(n2814) );
  NANDN U2892 ( .A(n2814), .B(n42095), .Z(n2774) );
  NAND U2893 ( .A(n2775), .B(n2774), .Z(n2827) );
  NANDN U2894 ( .A(n2776), .B(n42231), .Z(n2778) );
  XOR U2895 ( .A(n167), .B(a[60]), .Z(n2817) );
  NANDN U2896 ( .A(n2817), .B(n42234), .Z(n2777) );
  AND U2897 ( .A(n2778), .B(n2777), .Z(n2826) );
  XNOR U2898 ( .A(n2827), .B(n2826), .Z(n2828) );
  XNOR U2899 ( .A(n2829), .B(n2828), .Z(n2833) );
  NANDN U2900 ( .A(n2780), .B(n2779), .Z(n2784) );
  NAND U2901 ( .A(n2782), .B(n2781), .Z(n2783) );
  AND U2902 ( .A(n2784), .B(n2783), .Z(n2832) );
  XOR U2903 ( .A(n2833), .B(n2832), .Z(n2834) );
  NANDN U2904 ( .A(n2786), .B(n2785), .Z(n2790) );
  NANDN U2905 ( .A(n2788), .B(n2787), .Z(n2789) );
  NAND U2906 ( .A(n2790), .B(n2789), .Z(n2835) );
  XOR U2907 ( .A(n2834), .B(n2835), .Z(n2802) );
  OR U2908 ( .A(n2792), .B(n2791), .Z(n2796) );
  NANDN U2909 ( .A(n2794), .B(n2793), .Z(n2795) );
  NAND U2910 ( .A(n2796), .B(n2795), .Z(n2803) );
  XNOR U2911 ( .A(n2802), .B(n2803), .Z(n2804) );
  XNOR U2912 ( .A(n2805), .B(n2804), .Z(n2838) );
  XNOR U2913 ( .A(n2838), .B(sreg[1082]), .Z(n2840) );
  NAND U2914 ( .A(n2797), .B(sreg[1081]), .Z(n2801) );
  OR U2915 ( .A(n2799), .B(n2798), .Z(n2800) );
  AND U2916 ( .A(n2801), .B(n2800), .Z(n2839) );
  XOR U2917 ( .A(n2840), .B(n2839), .Z(c[1082]) );
  NANDN U2918 ( .A(n2803), .B(n2802), .Z(n2807) );
  NAND U2919 ( .A(n2805), .B(n2804), .Z(n2806) );
  NAND U2920 ( .A(n2807), .B(n2806), .Z(n2846) );
  NAND U2921 ( .A(b[0]), .B(a[67]), .Z(n2808) );
  XNOR U2922 ( .A(b[1]), .B(n2808), .Z(n2810) );
  NAND U2923 ( .A(n24), .B(a[66]), .Z(n2809) );
  AND U2924 ( .A(n2810), .B(n2809), .Z(n2863) );
  XOR U2925 ( .A(a[63]), .B(n42197), .Z(n2852) );
  NANDN U2926 ( .A(n2852), .B(n42173), .Z(n2813) );
  NANDN U2927 ( .A(n2811), .B(n42172), .Z(n2812) );
  NAND U2928 ( .A(n2813), .B(n2812), .Z(n2861) );
  NAND U2929 ( .A(b[7]), .B(a[59]), .Z(n2862) );
  XNOR U2930 ( .A(n2861), .B(n2862), .Z(n2864) );
  XOR U2931 ( .A(n2863), .B(n2864), .Z(n2870) );
  NANDN U2932 ( .A(n2814), .B(n42093), .Z(n2816) );
  XOR U2933 ( .A(n42134), .B(a[65]), .Z(n2855) );
  NANDN U2934 ( .A(n2855), .B(n42095), .Z(n2815) );
  NAND U2935 ( .A(n2816), .B(n2815), .Z(n2868) );
  NANDN U2936 ( .A(n2817), .B(n42231), .Z(n2819) );
  XOR U2937 ( .A(n167), .B(a[61]), .Z(n2858) );
  NANDN U2938 ( .A(n2858), .B(n42234), .Z(n2818) );
  AND U2939 ( .A(n2819), .B(n2818), .Z(n2867) );
  XNOR U2940 ( .A(n2868), .B(n2867), .Z(n2869) );
  XNOR U2941 ( .A(n2870), .B(n2869), .Z(n2874) );
  NANDN U2942 ( .A(n2821), .B(n2820), .Z(n2825) );
  NAND U2943 ( .A(n2823), .B(n2822), .Z(n2824) );
  AND U2944 ( .A(n2825), .B(n2824), .Z(n2873) );
  XOR U2945 ( .A(n2874), .B(n2873), .Z(n2875) );
  NANDN U2946 ( .A(n2827), .B(n2826), .Z(n2831) );
  NANDN U2947 ( .A(n2829), .B(n2828), .Z(n2830) );
  NAND U2948 ( .A(n2831), .B(n2830), .Z(n2876) );
  XOR U2949 ( .A(n2875), .B(n2876), .Z(n2843) );
  OR U2950 ( .A(n2833), .B(n2832), .Z(n2837) );
  NANDN U2951 ( .A(n2835), .B(n2834), .Z(n2836) );
  NAND U2952 ( .A(n2837), .B(n2836), .Z(n2844) );
  XNOR U2953 ( .A(n2843), .B(n2844), .Z(n2845) );
  XNOR U2954 ( .A(n2846), .B(n2845), .Z(n2879) );
  XNOR U2955 ( .A(n2879), .B(sreg[1083]), .Z(n2881) );
  NAND U2956 ( .A(n2838), .B(sreg[1082]), .Z(n2842) );
  OR U2957 ( .A(n2840), .B(n2839), .Z(n2841) );
  AND U2958 ( .A(n2842), .B(n2841), .Z(n2880) );
  XOR U2959 ( .A(n2881), .B(n2880), .Z(c[1083]) );
  NANDN U2960 ( .A(n2844), .B(n2843), .Z(n2848) );
  NAND U2961 ( .A(n2846), .B(n2845), .Z(n2847) );
  NAND U2962 ( .A(n2848), .B(n2847), .Z(n2887) );
  NAND U2963 ( .A(b[0]), .B(a[68]), .Z(n2849) );
  XNOR U2964 ( .A(b[1]), .B(n2849), .Z(n2851) );
  NAND U2965 ( .A(n24), .B(a[67]), .Z(n2850) );
  AND U2966 ( .A(n2851), .B(n2850), .Z(n2904) );
  XOR U2967 ( .A(a[64]), .B(n42197), .Z(n2893) );
  NANDN U2968 ( .A(n2893), .B(n42173), .Z(n2854) );
  NANDN U2969 ( .A(n2852), .B(n42172), .Z(n2853) );
  NAND U2970 ( .A(n2854), .B(n2853), .Z(n2902) );
  NAND U2971 ( .A(b[7]), .B(a[60]), .Z(n2903) );
  XNOR U2972 ( .A(n2902), .B(n2903), .Z(n2905) );
  XOR U2973 ( .A(n2904), .B(n2905), .Z(n2911) );
  NANDN U2974 ( .A(n2855), .B(n42093), .Z(n2857) );
  XOR U2975 ( .A(n42134), .B(a[66]), .Z(n2896) );
  NANDN U2976 ( .A(n2896), .B(n42095), .Z(n2856) );
  NAND U2977 ( .A(n2857), .B(n2856), .Z(n2909) );
  NANDN U2978 ( .A(n2858), .B(n42231), .Z(n2860) );
  XOR U2979 ( .A(n167), .B(a[62]), .Z(n2899) );
  NANDN U2980 ( .A(n2899), .B(n42234), .Z(n2859) );
  AND U2981 ( .A(n2860), .B(n2859), .Z(n2908) );
  XNOR U2982 ( .A(n2909), .B(n2908), .Z(n2910) );
  XNOR U2983 ( .A(n2911), .B(n2910), .Z(n2915) );
  NANDN U2984 ( .A(n2862), .B(n2861), .Z(n2866) );
  NAND U2985 ( .A(n2864), .B(n2863), .Z(n2865) );
  AND U2986 ( .A(n2866), .B(n2865), .Z(n2914) );
  XOR U2987 ( .A(n2915), .B(n2914), .Z(n2916) );
  NANDN U2988 ( .A(n2868), .B(n2867), .Z(n2872) );
  NANDN U2989 ( .A(n2870), .B(n2869), .Z(n2871) );
  NAND U2990 ( .A(n2872), .B(n2871), .Z(n2917) );
  XOR U2991 ( .A(n2916), .B(n2917), .Z(n2884) );
  OR U2992 ( .A(n2874), .B(n2873), .Z(n2878) );
  NANDN U2993 ( .A(n2876), .B(n2875), .Z(n2877) );
  NAND U2994 ( .A(n2878), .B(n2877), .Z(n2885) );
  XNOR U2995 ( .A(n2884), .B(n2885), .Z(n2886) );
  XNOR U2996 ( .A(n2887), .B(n2886), .Z(n2920) );
  XNOR U2997 ( .A(n2920), .B(sreg[1084]), .Z(n2922) );
  NAND U2998 ( .A(n2879), .B(sreg[1083]), .Z(n2883) );
  OR U2999 ( .A(n2881), .B(n2880), .Z(n2882) );
  AND U3000 ( .A(n2883), .B(n2882), .Z(n2921) );
  XOR U3001 ( .A(n2922), .B(n2921), .Z(c[1084]) );
  NANDN U3002 ( .A(n2885), .B(n2884), .Z(n2889) );
  NAND U3003 ( .A(n2887), .B(n2886), .Z(n2888) );
  NAND U3004 ( .A(n2889), .B(n2888), .Z(n2928) );
  NAND U3005 ( .A(b[0]), .B(a[69]), .Z(n2890) );
  XNOR U3006 ( .A(b[1]), .B(n2890), .Z(n2892) );
  NAND U3007 ( .A(n24), .B(a[68]), .Z(n2891) );
  AND U3008 ( .A(n2892), .B(n2891), .Z(n2945) );
  XOR U3009 ( .A(a[65]), .B(n42197), .Z(n2934) );
  NANDN U3010 ( .A(n2934), .B(n42173), .Z(n2895) );
  NANDN U3011 ( .A(n2893), .B(n42172), .Z(n2894) );
  NAND U3012 ( .A(n2895), .B(n2894), .Z(n2943) );
  NAND U3013 ( .A(b[7]), .B(a[61]), .Z(n2944) );
  XNOR U3014 ( .A(n2943), .B(n2944), .Z(n2946) );
  XOR U3015 ( .A(n2945), .B(n2946), .Z(n2952) );
  NANDN U3016 ( .A(n2896), .B(n42093), .Z(n2898) );
  XOR U3017 ( .A(n42134), .B(a[67]), .Z(n2937) );
  NANDN U3018 ( .A(n2937), .B(n42095), .Z(n2897) );
  NAND U3019 ( .A(n2898), .B(n2897), .Z(n2950) );
  NANDN U3020 ( .A(n2899), .B(n42231), .Z(n2901) );
  XOR U3021 ( .A(n167), .B(a[63]), .Z(n2940) );
  NANDN U3022 ( .A(n2940), .B(n42234), .Z(n2900) );
  AND U3023 ( .A(n2901), .B(n2900), .Z(n2949) );
  XNOR U3024 ( .A(n2950), .B(n2949), .Z(n2951) );
  XNOR U3025 ( .A(n2952), .B(n2951), .Z(n2956) );
  NANDN U3026 ( .A(n2903), .B(n2902), .Z(n2907) );
  NAND U3027 ( .A(n2905), .B(n2904), .Z(n2906) );
  AND U3028 ( .A(n2907), .B(n2906), .Z(n2955) );
  XOR U3029 ( .A(n2956), .B(n2955), .Z(n2957) );
  NANDN U3030 ( .A(n2909), .B(n2908), .Z(n2913) );
  NANDN U3031 ( .A(n2911), .B(n2910), .Z(n2912) );
  NAND U3032 ( .A(n2913), .B(n2912), .Z(n2958) );
  XOR U3033 ( .A(n2957), .B(n2958), .Z(n2925) );
  OR U3034 ( .A(n2915), .B(n2914), .Z(n2919) );
  NANDN U3035 ( .A(n2917), .B(n2916), .Z(n2918) );
  NAND U3036 ( .A(n2919), .B(n2918), .Z(n2926) );
  XNOR U3037 ( .A(n2925), .B(n2926), .Z(n2927) );
  XNOR U3038 ( .A(n2928), .B(n2927), .Z(n2961) );
  XNOR U3039 ( .A(n2961), .B(sreg[1085]), .Z(n2963) );
  NAND U3040 ( .A(n2920), .B(sreg[1084]), .Z(n2924) );
  OR U3041 ( .A(n2922), .B(n2921), .Z(n2923) );
  AND U3042 ( .A(n2924), .B(n2923), .Z(n2962) );
  XOR U3043 ( .A(n2963), .B(n2962), .Z(c[1085]) );
  NANDN U3044 ( .A(n2926), .B(n2925), .Z(n2930) );
  NAND U3045 ( .A(n2928), .B(n2927), .Z(n2929) );
  NAND U3046 ( .A(n2930), .B(n2929), .Z(n2969) );
  NAND U3047 ( .A(b[0]), .B(a[70]), .Z(n2931) );
  XNOR U3048 ( .A(b[1]), .B(n2931), .Z(n2933) );
  NAND U3049 ( .A(n25), .B(a[69]), .Z(n2932) );
  AND U3050 ( .A(n2933), .B(n2932), .Z(n2986) );
  XOR U3051 ( .A(a[66]), .B(n42197), .Z(n2975) );
  NANDN U3052 ( .A(n2975), .B(n42173), .Z(n2936) );
  NANDN U3053 ( .A(n2934), .B(n42172), .Z(n2935) );
  NAND U3054 ( .A(n2936), .B(n2935), .Z(n2984) );
  NAND U3055 ( .A(b[7]), .B(a[62]), .Z(n2985) );
  XNOR U3056 ( .A(n2984), .B(n2985), .Z(n2987) );
  XOR U3057 ( .A(n2986), .B(n2987), .Z(n2993) );
  NANDN U3058 ( .A(n2937), .B(n42093), .Z(n2939) );
  XOR U3059 ( .A(n42134), .B(a[68]), .Z(n2978) );
  NANDN U3060 ( .A(n2978), .B(n42095), .Z(n2938) );
  NAND U3061 ( .A(n2939), .B(n2938), .Z(n2991) );
  NANDN U3062 ( .A(n2940), .B(n42231), .Z(n2942) );
  XOR U3063 ( .A(n167), .B(a[64]), .Z(n2981) );
  NANDN U3064 ( .A(n2981), .B(n42234), .Z(n2941) );
  AND U3065 ( .A(n2942), .B(n2941), .Z(n2990) );
  XNOR U3066 ( .A(n2991), .B(n2990), .Z(n2992) );
  XNOR U3067 ( .A(n2993), .B(n2992), .Z(n2997) );
  NANDN U3068 ( .A(n2944), .B(n2943), .Z(n2948) );
  NAND U3069 ( .A(n2946), .B(n2945), .Z(n2947) );
  AND U3070 ( .A(n2948), .B(n2947), .Z(n2996) );
  XOR U3071 ( .A(n2997), .B(n2996), .Z(n2998) );
  NANDN U3072 ( .A(n2950), .B(n2949), .Z(n2954) );
  NANDN U3073 ( .A(n2952), .B(n2951), .Z(n2953) );
  NAND U3074 ( .A(n2954), .B(n2953), .Z(n2999) );
  XOR U3075 ( .A(n2998), .B(n2999), .Z(n2966) );
  OR U3076 ( .A(n2956), .B(n2955), .Z(n2960) );
  NANDN U3077 ( .A(n2958), .B(n2957), .Z(n2959) );
  NAND U3078 ( .A(n2960), .B(n2959), .Z(n2967) );
  XNOR U3079 ( .A(n2966), .B(n2967), .Z(n2968) );
  XNOR U3080 ( .A(n2969), .B(n2968), .Z(n3002) );
  XNOR U3081 ( .A(n3002), .B(sreg[1086]), .Z(n3004) );
  NAND U3082 ( .A(n2961), .B(sreg[1085]), .Z(n2965) );
  OR U3083 ( .A(n2963), .B(n2962), .Z(n2964) );
  AND U3084 ( .A(n2965), .B(n2964), .Z(n3003) );
  XOR U3085 ( .A(n3004), .B(n3003), .Z(c[1086]) );
  NANDN U3086 ( .A(n2967), .B(n2966), .Z(n2971) );
  NAND U3087 ( .A(n2969), .B(n2968), .Z(n2970) );
  NAND U3088 ( .A(n2971), .B(n2970), .Z(n3010) );
  NAND U3089 ( .A(b[0]), .B(a[71]), .Z(n2972) );
  XNOR U3090 ( .A(b[1]), .B(n2972), .Z(n2974) );
  NAND U3091 ( .A(n25), .B(a[70]), .Z(n2973) );
  AND U3092 ( .A(n2974), .B(n2973), .Z(n3027) );
  XOR U3093 ( .A(a[67]), .B(n42197), .Z(n3016) );
  NANDN U3094 ( .A(n3016), .B(n42173), .Z(n2977) );
  NANDN U3095 ( .A(n2975), .B(n42172), .Z(n2976) );
  NAND U3096 ( .A(n2977), .B(n2976), .Z(n3025) );
  NAND U3097 ( .A(b[7]), .B(a[63]), .Z(n3026) );
  XNOR U3098 ( .A(n3025), .B(n3026), .Z(n3028) );
  XOR U3099 ( .A(n3027), .B(n3028), .Z(n3034) );
  NANDN U3100 ( .A(n2978), .B(n42093), .Z(n2980) );
  XOR U3101 ( .A(n42134), .B(a[69]), .Z(n3019) );
  NANDN U3102 ( .A(n3019), .B(n42095), .Z(n2979) );
  NAND U3103 ( .A(n2980), .B(n2979), .Z(n3032) );
  NANDN U3104 ( .A(n2981), .B(n42231), .Z(n2983) );
  XOR U3105 ( .A(n167), .B(a[65]), .Z(n3022) );
  NANDN U3106 ( .A(n3022), .B(n42234), .Z(n2982) );
  AND U3107 ( .A(n2983), .B(n2982), .Z(n3031) );
  XNOR U3108 ( .A(n3032), .B(n3031), .Z(n3033) );
  XNOR U3109 ( .A(n3034), .B(n3033), .Z(n3038) );
  NANDN U3110 ( .A(n2985), .B(n2984), .Z(n2989) );
  NAND U3111 ( .A(n2987), .B(n2986), .Z(n2988) );
  AND U3112 ( .A(n2989), .B(n2988), .Z(n3037) );
  XOR U3113 ( .A(n3038), .B(n3037), .Z(n3039) );
  NANDN U3114 ( .A(n2991), .B(n2990), .Z(n2995) );
  NANDN U3115 ( .A(n2993), .B(n2992), .Z(n2994) );
  NAND U3116 ( .A(n2995), .B(n2994), .Z(n3040) );
  XOR U3117 ( .A(n3039), .B(n3040), .Z(n3007) );
  OR U3118 ( .A(n2997), .B(n2996), .Z(n3001) );
  NANDN U3119 ( .A(n2999), .B(n2998), .Z(n3000) );
  NAND U3120 ( .A(n3001), .B(n3000), .Z(n3008) );
  XNOR U3121 ( .A(n3007), .B(n3008), .Z(n3009) );
  XNOR U3122 ( .A(n3010), .B(n3009), .Z(n3043) );
  XNOR U3123 ( .A(n3043), .B(sreg[1087]), .Z(n3045) );
  NAND U3124 ( .A(n3002), .B(sreg[1086]), .Z(n3006) );
  OR U3125 ( .A(n3004), .B(n3003), .Z(n3005) );
  AND U3126 ( .A(n3006), .B(n3005), .Z(n3044) );
  XOR U3127 ( .A(n3045), .B(n3044), .Z(c[1087]) );
  NANDN U3128 ( .A(n3008), .B(n3007), .Z(n3012) );
  NAND U3129 ( .A(n3010), .B(n3009), .Z(n3011) );
  NAND U3130 ( .A(n3012), .B(n3011), .Z(n3051) );
  NAND U3131 ( .A(b[0]), .B(a[72]), .Z(n3013) );
  XNOR U3132 ( .A(b[1]), .B(n3013), .Z(n3015) );
  NAND U3133 ( .A(n25), .B(a[71]), .Z(n3014) );
  AND U3134 ( .A(n3015), .B(n3014), .Z(n3068) );
  XOR U3135 ( .A(a[68]), .B(n42197), .Z(n3057) );
  NANDN U3136 ( .A(n3057), .B(n42173), .Z(n3018) );
  NANDN U3137 ( .A(n3016), .B(n42172), .Z(n3017) );
  NAND U3138 ( .A(n3018), .B(n3017), .Z(n3066) );
  NAND U3139 ( .A(b[7]), .B(a[64]), .Z(n3067) );
  XNOR U3140 ( .A(n3066), .B(n3067), .Z(n3069) );
  XOR U3141 ( .A(n3068), .B(n3069), .Z(n3075) );
  NANDN U3142 ( .A(n3019), .B(n42093), .Z(n3021) );
  XOR U3143 ( .A(n42134), .B(a[70]), .Z(n3060) );
  NANDN U3144 ( .A(n3060), .B(n42095), .Z(n3020) );
  NAND U3145 ( .A(n3021), .B(n3020), .Z(n3073) );
  NANDN U3146 ( .A(n3022), .B(n42231), .Z(n3024) );
  XOR U3147 ( .A(n167), .B(a[66]), .Z(n3063) );
  NANDN U3148 ( .A(n3063), .B(n42234), .Z(n3023) );
  AND U3149 ( .A(n3024), .B(n3023), .Z(n3072) );
  XNOR U3150 ( .A(n3073), .B(n3072), .Z(n3074) );
  XNOR U3151 ( .A(n3075), .B(n3074), .Z(n3079) );
  NANDN U3152 ( .A(n3026), .B(n3025), .Z(n3030) );
  NAND U3153 ( .A(n3028), .B(n3027), .Z(n3029) );
  AND U3154 ( .A(n3030), .B(n3029), .Z(n3078) );
  XOR U3155 ( .A(n3079), .B(n3078), .Z(n3080) );
  NANDN U3156 ( .A(n3032), .B(n3031), .Z(n3036) );
  NANDN U3157 ( .A(n3034), .B(n3033), .Z(n3035) );
  NAND U3158 ( .A(n3036), .B(n3035), .Z(n3081) );
  XOR U3159 ( .A(n3080), .B(n3081), .Z(n3048) );
  OR U3160 ( .A(n3038), .B(n3037), .Z(n3042) );
  NANDN U3161 ( .A(n3040), .B(n3039), .Z(n3041) );
  NAND U3162 ( .A(n3042), .B(n3041), .Z(n3049) );
  XNOR U3163 ( .A(n3048), .B(n3049), .Z(n3050) );
  XNOR U3164 ( .A(n3051), .B(n3050), .Z(n3084) );
  XNOR U3165 ( .A(n3084), .B(sreg[1088]), .Z(n3086) );
  NAND U3166 ( .A(n3043), .B(sreg[1087]), .Z(n3047) );
  OR U3167 ( .A(n3045), .B(n3044), .Z(n3046) );
  AND U3168 ( .A(n3047), .B(n3046), .Z(n3085) );
  XOR U3169 ( .A(n3086), .B(n3085), .Z(c[1088]) );
  NANDN U3170 ( .A(n3049), .B(n3048), .Z(n3053) );
  NAND U3171 ( .A(n3051), .B(n3050), .Z(n3052) );
  NAND U3172 ( .A(n3053), .B(n3052), .Z(n3092) );
  NAND U3173 ( .A(b[0]), .B(a[73]), .Z(n3054) );
  XNOR U3174 ( .A(b[1]), .B(n3054), .Z(n3056) );
  NAND U3175 ( .A(n25), .B(a[72]), .Z(n3055) );
  AND U3176 ( .A(n3056), .B(n3055), .Z(n3109) );
  XOR U3177 ( .A(a[69]), .B(n42197), .Z(n3098) );
  NANDN U3178 ( .A(n3098), .B(n42173), .Z(n3059) );
  NANDN U3179 ( .A(n3057), .B(n42172), .Z(n3058) );
  NAND U3180 ( .A(n3059), .B(n3058), .Z(n3107) );
  NAND U3181 ( .A(b[7]), .B(a[65]), .Z(n3108) );
  XNOR U3182 ( .A(n3107), .B(n3108), .Z(n3110) );
  XOR U3183 ( .A(n3109), .B(n3110), .Z(n3116) );
  NANDN U3184 ( .A(n3060), .B(n42093), .Z(n3062) );
  XOR U3185 ( .A(n42134), .B(a[71]), .Z(n3101) );
  NANDN U3186 ( .A(n3101), .B(n42095), .Z(n3061) );
  NAND U3187 ( .A(n3062), .B(n3061), .Z(n3114) );
  NANDN U3188 ( .A(n3063), .B(n42231), .Z(n3065) );
  XOR U3189 ( .A(n167), .B(a[67]), .Z(n3104) );
  NANDN U3190 ( .A(n3104), .B(n42234), .Z(n3064) );
  AND U3191 ( .A(n3065), .B(n3064), .Z(n3113) );
  XNOR U3192 ( .A(n3114), .B(n3113), .Z(n3115) );
  XNOR U3193 ( .A(n3116), .B(n3115), .Z(n3120) );
  NANDN U3194 ( .A(n3067), .B(n3066), .Z(n3071) );
  NAND U3195 ( .A(n3069), .B(n3068), .Z(n3070) );
  AND U3196 ( .A(n3071), .B(n3070), .Z(n3119) );
  XOR U3197 ( .A(n3120), .B(n3119), .Z(n3121) );
  NANDN U3198 ( .A(n3073), .B(n3072), .Z(n3077) );
  NANDN U3199 ( .A(n3075), .B(n3074), .Z(n3076) );
  NAND U3200 ( .A(n3077), .B(n3076), .Z(n3122) );
  XOR U3201 ( .A(n3121), .B(n3122), .Z(n3089) );
  OR U3202 ( .A(n3079), .B(n3078), .Z(n3083) );
  NANDN U3203 ( .A(n3081), .B(n3080), .Z(n3082) );
  NAND U3204 ( .A(n3083), .B(n3082), .Z(n3090) );
  XNOR U3205 ( .A(n3089), .B(n3090), .Z(n3091) );
  XNOR U3206 ( .A(n3092), .B(n3091), .Z(n3125) );
  XNOR U3207 ( .A(n3125), .B(sreg[1089]), .Z(n3127) );
  NAND U3208 ( .A(n3084), .B(sreg[1088]), .Z(n3088) );
  OR U3209 ( .A(n3086), .B(n3085), .Z(n3087) );
  AND U3210 ( .A(n3088), .B(n3087), .Z(n3126) );
  XOR U3211 ( .A(n3127), .B(n3126), .Z(c[1089]) );
  NANDN U3212 ( .A(n3090), .B(n3089), .Z(n3094) );
  NAND U3213 ( .A(n3092), .B(n3091), .Z(n3093) );
  NAND U3214 ( .A(n3094), .B(n3093), .Z(n3133) );
  NAND U3215 ( .A(b[0]), .B(a[74]), .Z(n3095) );
  XNOR U3216 ( .A(b[1]), .B(n3095), .Z(n3097) );
  NAND U3217 ( .A(n25), .B(a[73]), .Z(n3096) );
  AND U3218 ( .A(n3097), .B(n3096), .Z(n3150) );
  XOR U3219 ( .A(a[70]), .B(n42197), .Z(n3139) );
  NANDN U3220 ( .A(n3139), .B(n42173), .Z(n3100) );
  NANDN U3221 ( .A(n3098), .B(n42172), .Z(n3099) );
  NAND U3222 ( .A(n3100), .B(n3099), .Z(n3148) );
  NAND U3223 ( .A(b[7]), .B(a[66]), .Z(n3149) );
  XNOR U3224 ( .A(n3148), .B(n3149), .Z(n3151) );
  XOR U3225 ( .A(n3150), .B(n3151), .Z(n3157) );
  NANDN U3226 ( .A(n3101), .B(n42093), .Z(n3103) );
  XOR U3227 ( .A(n42134), .B(a[72]), .Z(n3142) );
  NANDN U3228 ( .A(n3142), .B(n42095), .Z(n3102) );
  NAND U3229 ( .A(n3103), .B(n3102), .Z(n3155) );
  NANDN U3230 ( .A(n3104), .B(n42231), .Z(n3106) );
  XOR U3231 ( .A(n167), .B(a[68]), .Z(n3145) );
  NANDN U3232 ( .A(n3145), .B(n42234), .Z(n3105) );
  AND U3233 ( .A(n3106), .B(n3105), .Z(n3154) );
  XNOR U3234 ( .A(n3155), .B(n3154), .Z(n3156) );
  XNOR U3235 ( .A(n3157), .B(n3156), .Z(n3161) );
  NANDN U3236 ( .A(n3108), .B(n3107), .Z(n3112) );
  NAND U3237 ( .A(n3110), .B(n3109), .Z(n3111) );
  AND U3238 ( .A(n3112), .B(n3111), .Z(n3160) );
  XOR U3239 ( .A(n3161), .B(n3160), .Z(n3162) );
  NANDN U3240 ( .A(n3114), .B(n3113), .Z(n3118) );
  NANDN U3241 ( .A(n3116), .B(n3115), .Z(n3117) );
  NAND U3242 ( .A(n3118), .B(n3117), .Z(n3163) );
  XOR U3243 ( .A(n3162), .B(n3163), .Z(n3130) );
  OR U3244 ( .A(n3120), .B(n3119), .Z(n3124) );
  NANDN U3245 ( .A(n3122), .B(n3121), .Z(n3123) );
  NAND U3246 ( .A(n3124), .B(n3123), .Z(n3131) );
  XNOR U3247 ( .A(n3130), .B(n3131), .Z(n3132) );
  XNOR U3248 ( .A(n3133), .B(n3132), .Z(n3166) );
  XNOR U3249 ( .A(n3166), .B(sreg[1090]), .Z(n3168) );
  NAND U3250 ( .A(n3125), .B(sreg[1089]), .Z(n3129) );
  OR U3251 ( .A(n3127), .B(n3126), .Z(n3128) );
  AND U3252 ( .A(n3129), .B(n3128), .Z(n3167) );
  XOR U3253 ( .A(n3168), .B(n3167), .Z(c[1090]) );
  NANDN U3254 ( .A(n3131), .B(n3130), .Z(n3135) );
  NAND U3255 ( .A(n3133), .B(n3132), .Z(n3134) );
  NAND U3256 ( .A(n3135), .B(n3134), .Z(n3174) );
  NAND U3257 ( .A(b[0]), .B(a[75]), .Z(n3136) );
  XNOR U3258 ( .A(b[1]), .B(n3136), .Z(n3138) );
  NAND U3259 ( .A(n25), .B(a[74]), .Z(n3137) );
  AND U3260 ( .A(n3138), .B(n3137), .Z(n3191) );
  XOR U3261 ( .A(a[71]), .B(n42197), .Z(n3180) );
  NANDN U3262 ( .A(n3180), .B(n42173), .Z(n3141) );
  NANDN U3263 ( .A(n3139), .B(n42172), .Z(n3140) );
  NAND U3264 ( .A(n3141), .B(n3140), .Z(n3189) );
  NAND U3265 ( .A(b[7]), .B(a[67]), .Z(n3190) );
  XNOR U3266 ( .A(n3189), .B(n3190), .Z(n3192) );
  XOR U3267 ( .A(n3191), .B(n3192), .Z(n3198) );
  NANDN U3268 ( .A(n3142), .B(n42093), .Z(n3144) );
  XOR U3269 ( .A(n42134), .B(a[73]), .Z(n3183) );
  NANDN U3270 ( .A(n3183), .B(n42095), .Z(n3143) );
  NAND U3271 ( .A(n3144), .B(n3143), .Z(n3196) );
  NANDN U3272 ( .A(n3145), .B(n42231), .Z(n3147) );
  XOR U3273 ( .A(n167), .B(a[69]), .Z(n3186) );
  NANDN U3274 ( .A(n3186), .B(n42234), .Z(n3146) );
  AND U3275 ( .A(n3147), .B(n3146), .Z(n3195) );
  XNOR U3276 ( .A(n3196), .B(n3195), .Z(n3197) );
  XNOR U3277 ( .A(n3198), .B(n3197), .Z(n3202) );
  NANDN U3278 ( .A(n3149), .B(n3148), .Z(n3153) );
  NAND U3279 ( .A(n3151), .B(n3150), .Z(n3152) );
  AND U3280 ( .A(n3153), .B(n3152), .Z(n3201) );
  XOR U3281 ( .A(n3202), .B(n3201), .Z(n3203) );
  NANDN U3282 ( .A(n3155), .B(n3154), .Z(n3159) );
  NANDN U3283 ( .A(n3157), .B(n3156), .Z(n3158) );
  NAND U3284 ( .A(n3159), .B(n3158), .Z(n3204) );
  XOR U3285 ( .A(n3203), .B(n3204), .Z(n3171) );
  OR U3286 ( .A(n3161), .B(n3160), .Z(n3165) );
  NANDN U3287 ( .A(n3163), .B(n3162), .Z(n3164) );
  NAND U3288 ( .A(n3165), .B(n3164), .Z(n3172) );
  XNOR U3289 ( .A(n3171), .B(n3172), .Z(n3173) );
  XNOR U3290 ( .A(n3174), .B(n3173), .Z(n3207) );
  XNOR U3291 ( .A(n3207), .B(sreg[1091]), .Z(n3209) );
  NAND U3292 ( .A(n3166), .B(sreg[1090]), .Z(n3170) );
  OR U3293 ( .A(n3168), .B(n3167), .Z(n3169) );
  AND U3294 ( .A(n3170), .B(n3169), .Z(n3208) );
  XOR U3295 ( .A(n3209), .B(n3208), .Z(c[1091]) );
  NANDN U3296 ( .A(n3172), .B(n3171), .Z(n3176) );
  NAND U3297 ( .A(n3174), .B(n3173), .Z(n3175) );
  NAND U3298 ( .A(n3176), .B(n3175), .Z(n3215) );
  NAND U3299 ( .A(b[0]), .B(a[76]), .Z(n3177) );
  XNOR U3300 ( .A(b[1]), .B(n3177), .Z(n3179) );
  NAND U3301 ( .A(n25), .B(a[75]), .Z(n3178) );
  AND U3302 ( .A(n3179), .B(n3178), .Z(n3232) );
  XOR U3303 ( .A(a[72]), .B(n42197), .Z(n3221) );
  NANDN U3304 ( .A(n3221), .B(n42173), .Z(n3182) );
  NANDN U3305 ( .A(n3180), .B(n42172), .Z(n3181) );
  NAND U3306 ( .A(n3182), .B(n3181), .Z(n3230) );
  NAND U3307 ( .A(b[7]), .B(a[68]), .Z(n3231) );
  XNOR U3308 ( .A(n3230), .B(n3231), .Z(n3233) );
  XOR U3309 ( .A(n3232), .B(n3233), .Z(n3239) );
  NANDN U3310 ( .A(n3183), .B(n42093), .Z(n3185) );
  XOR U3311 ( .A(n42134), .B(a[74]), .Z(n3224) );
  NANDN U3312 ( .A(n3224), .B(n42095), .Z(n3184) );
  NAND U3313 ( .A(n3185), .B(n3184), .Z(n3237) );
  NANDN U3314 ( .A(n3186), .B(n42231), .Z(n3188) );
  XOR U3315 ( .A(n167), .B(a[70]), .Z(n3227) );
  NANDN U3316 ( .A(n3227), .B(n42234), .Z(n3187) );
  AND U3317 ( .A(n3188), .B(n3187), .Z(n3236) );
  XNOR U3318 ( .A(n3237), .B(n3236), .Z(n3238) );
  XNOR U3319 ( .A(n3239), .B(n3238), .Z(n3243) );
  NANDN U3320 ( .A(n3190), .B(n3189), .Z(n3194) );
  NAND U3321 ( .A(n3192), .B(n3191), .Z(n3193) );
  AND U3322 ( .A(n3194), .B(n3193), .Z(n3242) );
  XOR U3323 ( .A(n3243), .B(n3242), .Z(n3244) );
  NANDN U3324 ( .A(n3196), .B(n3195), .Z(n3200) );
  NANDN U3325 ( .A(n3198), .B(n3197), .Z(n3199) );
  NAND U3326 ( .A(n3200), .B(n3199), .Z(n3245) );
  XOR U3327 ( .A(n3244), .B(n3245), .Z(n3212) );
  OR U3328 ( .A(n3202), .B(n3201), .Z(n3206) );
  NANDN U3329 ( .A(n3204), .B(n3203), .Z(n3205) );
  NAND U3330 ( .A(n3206), .B(n3205), .Z(n3213) );
  XNOR U3331 ( .A(n3212), .B(n3213), .Z(n3214) );
  XNOR U3332 ( .A(n3215), .B(n3214), .Z(n3248) );
  XNOR U3333 ( .A(n3248), .B(sreg[1092]), .Z(n3250) );
  NAND U3334 ( .A(n3207), .B(sreg[1091]), .Z(n3211) );
  OR U3335 ( .A(n3209), .B(n3208), .Z(n3210) );
  AND U3336 ( .A(n3211), .B(n3210), .Z(n3249) );
  XOR U3337 ( .A(n3250), .B(n3249), .Z(c[1092]) );
  NANDN U3338 ( .A(n3213), .B(n3212), .Z(n3217) );
  NAND U3339 ( .A(n3215), .B(n3214), .Z(n3216) );
  NAND U3340 ( .A(n3217), .B(n3216), .Z(n3256) );
  NAND U3341 ( .A(b[0]), .B(a[77]), .Z(n3218) );
  XNOR U3342 ( .A(b[1]), .B(n3218), .Z(n3220) );
  NAND U3343 ( .A(n26), .B(a[76]), .Z(n3219) );
  AND U3344 ( .A(n3220), .B(n3219), .Z(n3273) );
  XOR U3345 ( .A(a[73]), .B(n42197), .Z(n3262) );
  NANDN U3346 ( .A(n3262), .B(n42173), .Z(n3223) );
  NANDN U3347 ( .A(n3221), .B(n42172), .Z(n3222) );
  NAND U3348 ( .A(n3223), .B(n3222), .Z(n3271) );
  NAND U3349 ( .A(b[7]), .B(a[69]), .Z(n3272) );
  XNOR U3350 ( .A(n3271), .B(n3272), .Z(n3274) );
  XOR U3351 ( .A(n3273), .B(n3274), .Z(n3280) );
  NANDN U3352 ( .A(n3224), .B(n42093), .Z(n3226) );
  XOR U3353 ( .A(n42134), .B(a[75]), .Z(n3265) );
  NANDN U3354 ( .A(n3265), .B(n42095), .Z(n3225) );
  NAND U3355 ( .A(n3226), .B(n3225), .Z(n3278) );
  NANDN U3356 ( .A(n3227), .B(n42231), .Z(n3229) );
  XOR U3357 ( .A(n168), .B(a[71]), .Z(n3268) );
  NANDN U3358 ( .A(n3268), .B(n42234), .Z(n3228) );
  AND U3359 ( .A(n3229), .B(n3228), .Z(n3277) );
  XNOR U3360 ( .A(n3278), .B(n3277), .Z(n3279) );
  XNOR U3361 ( .A(n3280), .B(n3279), .Z(n3284) );
  NANDN U3362 ( .A(n3231), .B(n3230), .Z(n3235) );
  NAND U3363 ( .A(n3233), .B(n3232), .Z(n3234) );
  AND U3364 ( .A(n3235), .B(n3234), .Z(n3283) );
  XOR U3365 ( .A(n3284), .B(n3283), .Z(n3285) );
  NANDN U3366 ( .A(n3237), .B(n3236), .Z(n3241) );
  NANDN U3367 ( .A(n3239), .B(n3238), .Z(n3240) );
  NAND U3368 ( .A(n3241), .B(n3240), .Z(n3286) );
  XOR U3369 ( .A(n3285), .B(n3286), .Z(n3253) );
  OR U3370 ( .A(n3243), .B(n3242), .Z(n3247) );
  NANDN U3371 ( .A(n3245), .B(n3244), .Z(n3246) );
  NAND U3372 ( .A(n3247), .B(n3246), .Z(n3254) );
  XNOR U3373 ( .A(n3253), .B(n3254), .Z(n3255) );
  XNOR U3374 ( .A(n3256), .B(n3255), .Z(n3289) );
  XNOR U3375 ( .A(n3289), .B(sreg[1093]), .Z(n3291) );
  NAND U3376 ( .A(n3248), .B(sreg[1092]), .Z(n3252) );
  OR U3377 ( .A(n3250), .B(n3249), .Z(n3251) );
  AND U3378 ( .A(n3252), .B(n3251), .Z(n3290) );
  XOR U3379 ( .A(n3291), .B(n3290), .Z(c[1093]) );
  NANDN U3380 ( .A(n3254), .B(n3253), .Z(n3258) );
  NAND U3381 ( .A(n3256), .B(n3255), .Z(n3257) );
  NAND U3382 ( .A(n3258), .B(n3257), .Z(n3297) );
  NAND U3383 ( .A(b[0]), .B(a[78]), .Z(n3259) );
  XNOR U3384 ( .A(b[1]), .B(n3259), .Z(n3261) );
  NAND U3385 ( .A(n26), .B(a[77]), .Z(n3260) );
  AND U3386 ( .A(n3261), .B(n3260), .Z(n3314) );
  XOR U3387 ( .A(a[74]), .B(n42197), .Z(n3303) );
  NANDN U3388 ( .A(n3303), .B(n42173), .Z(n3264) );
  NANDN U3389 ( .A(n3262), .B(n42172), .Z(n3263) );
  NAND U3390 ( .A(n3264), .B(n3263), .Z(n3312) );
  NAND U3391 ( .A(b[7]), .B(a[70]), .Z(n3313) );
  XNOR U3392 ( .A(n3312), .B(n3313), .Z(n3315) );
  XOR U3393 ( .A(n3314), .B(n3315), .Z(n3321) );
  NANDN U3394 ( .A(n3265), .B(n42093), .Z(n3267) );
  XOR U3395 ( .A(n42134), .B(a[76]), .Z(n3306) );
  NANDN U3396 ( .A(n3306), .B(n42095), .Z(n3266) );
  NAND U3397 ( .A(n3267), .B(n3266), .Z(n3319) );
  NANDN U3398 ( .A(n3268), .B(n42231), .Z(n3270) );
  XOR U3399 ( .A(n168), .B(a[72]), .Z(n3309) );
  NANDN U3400 ( .A(n3309), .B(n42234), .Z(n3269) );
  AND U3401 ( .A(n3270), .B(n3269), .Z(n3318) );
  XNOR U3402 ( .A(n3319), .B(n3318), .Z(n3320) );
  XNOR U3403 ( .A(n3321), .B(n3320), .Z(n3325) );
  NANDN U3404 ( .A(n3272), .B(n3271), .Z(n3276) );
  NAND U3405 ( .A(n3274), .B(n3273), .Z(n3275) );
  AND U3406 ( .A(n3276), .B(n3275), .Z(n3324) );
  XOR U3407 ( .A(n3325), .B(n3324), .Z(n3326) );
  NANDN U3408 ( .A(n3278), .B(n3277), .Z(n3282) );
  NANDN U3409 ( .A(n3280), .B(n3279), .Z(n3281) );
  NAND U3410 ( .A(n3282), .B(n3281), .Z(n3327) );
  XOR U3411 ( .A(n3326), .B(n3327), .Z(n3294) );
  OR U3412 ( .A(n3284), .B(n3283), .Z(n3288) );
  NANDN U3413 ( .A(n3286), .B(n3285), .Z(n3287) );
  NAND U3414 ( .A(n3288), .B(n3287), .Z(n3295) );
  XNOR U3415 ( .A(n3294), .B(n3295), .Z(n3296) );
  XNOR U3416 ( .A(n3297), .B(n3296), .Z(n3330) );
  XNOR U3417 ( .A(n3330), .B(sreg[1094]), .Z(n3332) );
  NAND U3418 ( .A(n3289), .B(sreg[1093]), .Z(n3293) );
  OR U3419 ( .A(n3291), .B(n3290), .Z(n3292) );
  AND U3420 ( .A(n3293), .B(n3292), .Z(n3331) );
  XOR U3421 ( .A(n3332), .B(n3331), .Z(c[1094]) );
  NANDN U3422 ( .A(n3295), .B(n3294), .Z(n3299) );
  NAND U3423 ( .A(n3297), .B(n3296), .Z(n3298) );
  NAND U3424 ( .A(n3299), .B(n3298), .Z(n3338) );
  NAND U3425 ( .A(b[0]), .B(a[79]), .Z(n3300) );
  XNOR U3426 ( .A(b[1]), .B(n3300), .Z(n3302) );
  NAND U3427 ( .A(n26), .B(a[78]), .Z(n3301) );
  AND U3428 ( .A(n3302), .B(n3301), .Z(n3355) );
  XOR U3429 ( .A(a[75]), .B(n42197), .Z(n3344) );
  NANDN U3430 ( .A(n3344), .B(n42173), .Z(n3305) );
  NANDN U3431 ( .A(n3303), .B(n42172), .Z(n3304) );
  NAND U3432 ( .A(n3305), .B(n3304), .Z(n3353) );
  NAND U3433 ( .A(b[7]), .B(a[71]), .Z(n3354) );
  XNOR U3434 ( .A(n3353), .B(n3354), .Z(n3356) );
  XOR U3435 ( .A(n3355), .B(n3356), .Z(n3362) );
  NANDN U3436 ( .A(n3306), .B(n42093), .Z(n3308) );
  XOR U3437 ( .A(n42134), .B(a[77]), .Z(n3347) );
  NANDN U3438 ( .A(n3347), .B(n42095), .Z(n3307) );
  NAND U3439 ( .A(n3308), .B(n3307), .Z(n3360) );
  NANDN U3440 ( .A(n3309), .B(n42231), .Z(n3311) );
  XOR U3441 ( .A(n168), .B(a[73]), .Z(n3350) );
  NANDN U3442 ( .A(n3350), .B(n42234), .Z(n3310) );
  AND U3443 ( .A(n3311), .B(n3310), .Z(n3359) );
  XNOR U3444 ( .A(n3360), .B(n3359), .Z(n3361) );
  XNOR U3445 ( .A(n3362), .B(n3361), .Z(n3366) );
  NANDN U3446 ( .A(n3313), .B(n3312), .Z(n3317) );
  NAND U3447 ( .A(n3315), .B(n3314), .Z(n3316) );
  AND U3448 ( .A(n3317), .B(n3316), .Z(n3365) );
  XOR U3449 ( .A(n3366), .B(n3365), .Z(n3367) );
  NANDN U3450 ( .A(n3319), .B(n3318), .Z(n3323) );
  NANDN U3451 ( .A(n3321), .B(n3320), .Z(n3322) );
  NAND U3452 ( .A(n3323), .B(n3322), .Z(n3368) );
  XOR U3453 ( .A(n3367), .B(n3368), .Z(n3335) );
  OR U3454 ( .A(n3325), .B(n3324), .Z(n3329) );
  NANDN U3455 ( .A(n3327), .B(n3326), .Z(n3328) );
  NAND U3456 ( .A(n3329), .B(n3328), .Z(n3336) );
  XNOR U3457 ( .A(n3335), .B(n3336), .Z(n3337) );
  XNOR U3458 ( .A(n3338), .B(n3337), .Z(n3371) );
  XNOR U3459 ( .A(n3371), .B(sreg[1095]), .Z(n3373) );
  NAND U3460 ( .A(n3330), .B(sreg[1094]), .Z(n3334) );
  OR U3461 ( .A(n3332), .B(n3331), .Z(n3333) );
  AND U3462 ( .A(n3334), .B(n3333), .Z(n3372) );
  XOR U3463 ( .A(n3373), .B(n3372), .Z(c[1095]) );
  NANDN U3464 ( .A(n3336), .B(n3335), .Z(n3340) );
  NAND U3465 ( .A(n3338), .B(n3337), .Z(n3339) );
  NAND U3466 ( .A(n3340), .B(n3339), .Z(n3379) );
  NAND U3467 ( .A(b[0]), .B(a[80]), .Z(n3341) );
  XNOR U3468 ( .A(b[1]), .B(n3341), .Z(n3343) );
  NAND U3469 ( .A(n26), .B(a[79]), .Z(n3342) );
  AND U3470 ( .A(n3343), .B(n3342), .Z(n3396) );
  XOR U3471 ( .A(a[76]), .B(n42197), .Z(n3385) );
  NANDN U3472 ( .A(n3385), .B(n42173), .Z(n3346) );
  NANDN U3473 ( .A(n3344), .B(n42172), .Z(n3345) );
  NAND U3474 ( .A(n3346), .B(n3345), .Z(n3394) );
  NAND U3475 ( .A(b[7]), .B(a[72]), .Z(n3395) );
  XNOR U3476 ( .A(n3394), .B(n3395), .Z(n3397) );
  XOR U3477 ( .A(n3396), .B(n3397), .Z(n3403) );
  NANDN U3478 ( .A(n3347), .B(n42093), .Z(n3349) );
  XOR U3479 ( .A(n42134), .B(a[78]), .Z(n3388) );
  NANDN U3480 ( .A(n3388), .B(n42095), .Z(n3348) );
  NAND U3481 ( .A(n3349), .B(n3348), .Z(n3401) );
  NANDN U3482 ( .A(n3350), .B(n42231), .Z(n3352) );
  XOR U3483 ( .A(n168), .B(a[74]), .Z(n3391) );
  NANDN U3484 ( .A(n3391), .B(n42234), .Z(n3351) );
  AND U3485 ( .A(n3352), .B(n3351), .Z(n3400) );
  XNOR U3486 ( .A(n3401), .B(n3400), .Z(n3402) );
  XNOR U3487 ( .A(n3403), .B(n3402), .Z(n3407) );
  NANDN U3488 ( .A(n3354), .B(n3353), .Z(n3358) );
  NAND U3489 ( .A(n3356), .B(n3355), .Z(n3357) );
  AND U3490 ( .A(n3358), .B(n3357), .Z(n3406) );
  XOR U3491 ( .A(n3407), .B(n3406), .Z(n3408) );
  NANDN U3492 ( .A(n3360), .B(n3359), .Z(n3364) );
  NANDN U3493 ( .A(n3362), .B(n3361), .Z(n3363) );
  NAND U3494 ( .A(n3364), .B(n3363), .Z(n3409) );
  XOR U3495 ( .A(n3408), .B(n3409), .Z(n3376) );
  OR U3496 ( .A(n3366), .B(n3365), .Z(n3370) );
  NANDN U3497 ( .A(n3368), .B(n3367), .Z(n3369) );
  NAND U3498 ( .A(n3370), .B(n3369), .Z(n3377) );
  XNOR U3499 ( .A(n3376), .B(n3377), .Z(n3378) );
  XNOR U3500 ( .A(n3379), .B(n3378), .Z(n3412) );
  XNOR U3501 ( .A(n3412), .B(sreg[1096]), .Z(n3414) );
  NAND U3502 ( .A(n3371), .B(sreg[1095]), .Z(n3375) );
  OR U3503 ( .A(n3373), .B(n3372), .Z(n3374) );
  AND U3504 ( .A(n3375), .B(n3374), .Z(n3413) );
  XOR U3505 ( .A(n3414), .B(n3413), .Z(c[1096]) );
  NANDN U3506 ( .A(n3377), .B(n3376), .Z(n3381) );
  NAND U3507 ( .A(n3379), .B(n3378), .Z(n3380) );
  NAND U3508 ( .A(n3381), .B(n3380), .Z(n3420) );
  NAND U3509 ( .A(b[0]), .B(a[81]), .Z(n3382) );
  XNOR U3510 ( .A(b[1]), .B(n3382), .Z(n3384) );
  NAND U3511 ( .A(n26), .B(a[80]), .Z(n3383) );
  AND U3512 ( .A(n3384), .B(n3383), .Z(n3437) );
  XOR U3513 ( .A(a[77]), .B(n42197), .Z(n3426) );
  NANDN U3514 ( .A(n3426), .B(n42173), .Z(n3387) );
  NANDN U3515 ( .A(n3385), .B(n42172), .Z(n3386) );
  NAND U3516 ( .A(n3387), .B(n3386), .Z(n3435) );
  NAND U3517 ( .A(b[7]), .B(a[73]), .Z(n3436) );
  XNOR U3518 ( .A(n3435), .B(n3436), .Z(n3438) );
  XOR U3519 ( .A(n3437), .B(n3438), .Z(n3444) );
  NANDN U3520 ( .A(n3388), .B(n42093), .Z(n3390) );
  XOR U3521 ( .A(n42134), .B(a[79]), .Z(n3429) );
  NANDN U3522 ( .A(n3429), .B(n42095), .Z(n3389) );
  NAND U3523 ( .A(n3390), .B(n3389), .Z(n3442) );
  NANDN U3524 ( .A(n3391), .B(n42231), .Z(n3393) );
  XOR U3525 ( .A(n168), .B(a[75]), .Z(n3432) );
  NANDN U3526 ( .A(n3432), .B(n42234), .Z(n3392) );
  AND U3527 ( .A(n3393), .B(n3392), .Z(n3441) );
  XNOR U3528 ( .A(n3442), .B(n3441), .Z(n3443) );
  XNOR U3529 ( .A(n3444), .B(n3443), .Z(n3448) );
  NANDN U3530 ( .A(n3395), .B(n3394), .Z(n3399) );
  NAND U3531 ( .A(n3397), .B(n3396), .Z(n3398) );
  AND U3532 ( .A(n3399), .B(n3398), .Z(n3447) );
  XOR U3533 ( .A(n3448), .B(n3447), .Z(n3449) );
  NANDN U3534 ( .A(n3401), .B(n3400), .Z(n3405) );
  NANDN U3535 ( .A(n3403), .B(n3402), .Z(n3404) );
  NAND U3536 ( .A(n3405), .B(n3404), .Z(n3450) );
  XOR U3537 ( .A(n3449), .B(n3450), .Z(n3417) );
  OR U3538 ( .A(n3407), .B(n3406), .Z(n3411) );
  NANDN U3539 ( .A(n3409), .B(n3408), .Z(n3410) );
  NAND U3540 ( .A(n3411), .B(n3410), .Z(n3418) );
  XNOR U3541 ( .A(n3417), .B(n3418), .Z(n3419) );
  XNOR U3542 ( .A(n3420), .B(n3419), .Z(n3453) );
  XNOR U3543 ( .A(n3453), .B(sreg[1097]), .Z(n3455) );
  NAND U3544 ( .A(n3412), .B(sreg[1096]), .Z(n3416) );
  OR U3545 ( .A(n3414), .B(n3413), .Z(n3415) );
  AND U3546 ( .A(n3416), .B(n3415), .Z(n3454) );
  XOR U3547 ( .A(n3455), .B(n3454), .Z(c[1097]) );
  NANDN U3548 ( .A(n3418), .B(n3417), .Z(n3422) );
  NAND U3549 ( .A(n3420), .B(n3419), .Z(n3421) );
  NAND U3550 ( .A(n3422), .B(n3421), .Z(n3461) );
  NAND U3551 ( .A(b[0]), .B(a[82]), .Z(n3423) );
  XNOR U3552 ( .A(b[1]), .B(n3423), .Z(n3425) );
  NAND U3553 ( .A(n26), .B(a[81]), .Z(n3424) );
  AND U3554 ( .A(n3425), .B(n3424), .Z(n3478) );
  XOR U3555 ( .A(a[78]), .B(n42197), .Z(n3467) );
  NANDN U3556 ( .A(n3467), .B(n42173), .Z(n3428) );
  NANDN U3557 ( .A(n3426), .B(n42172), .Z(n3427) );
  NAND U3558 ( .A(n3428), .B(n3427), .Z(n3476) );
  NAND U3559 ( .A(b[7]), .B(a[74]), .Z(n3477) );
  XNOR U3560 ( .A(n3476), .B(n3477), .Z(n3479) );
  XOR U3561 ( .A(n3478), .B(n3479), .Z(n3485) );
  NANDN U3562 ( .A(n3429), .B(n42093), .Z(n3431) );
  XOR U3563 ( .A(n42134), .B(a[80]), .Z(n3470) );
  NANDN U3564 ( .A(n3470), .B(n42095), .Z(n3430) );
  NAND U3565 ( .A(n3431), .B(n3430), .Z(n3483) );
  NANDN U3566 ( .A(n3432), .B(n42231), .Z(n3434) );
  XOR U3567 ( .A(n168), .B(a[76]), .Z(n3473) );
  NANDN U3568 ( .A(n3473), .B(n42234), .Z(n3433) );
  AND U3569 ( .A(n3434), .B(n3433), .Z(n3482) );
  XNOR U3570 ( .A(n3483), .B(n3482), .Z(n3484) );
  XNOR U3571 ( .A(n3485), .B(n3484), .Z(n3489) );
  NANDN U3572 ( .A(n3436), .B(n3435), .Z(n3440) );
  NAND U3573 ( .A(n3438), .B(n3437), .Z(n3439) );
  AND U3574 ( .A(n3440), .B(n3439), .Z(n3488) );
  XOR U3575 ( .A(n3489), .B(n3488), .Z(n3490) );
  NANDN U3576 ( .A(n3442), .B(n3441), .Z(n3446) );
  NANDN U3577 ( .A(n3444), .B(n3443), .Z(n3445) );
  NAND U3578 ( .A(n3446), .B(n3445), .Z(n3491) );
  XOR U3579 ( .A(n3490), .B(n3491), .Z(n3458) );
  OR U3580 ( .A(n3448), .B(n3447), .Z(n3452) );
  NANDN U3581 ( .A(n3450), .B(n3449), .Z(n3451) );
  NAND U3582 ( .A(n3452), .B(n3451), .Z(n3459) );
  XNOR U3583 ( .A(n3458), .B(n3459), .Z(n3460) );
  XNOR U3584 ( .A(n3461), .B(n3460), .Z(n3494) );
  XNOR U3585 ( .A(n3494), .B(sreg[1098]), .Z(n3496) );
  NAND U3586 ( .A(n3453), .B(sreg[1097]), .Z(n3457) );
  OR U3587 ( .A(n3455), .B(n3454), .Z(n3456) );
  AND U3588 ( .A(n3457), .B(n3456), .Z(n3495) );
  XOR U3589 ( .A(n3496), .B(n3495), .Z(c[1098]) );
  NANDN U3590 ( .A(n3459), .B(n3458), .Z(n3463) );
  NAND U3591 ( .A(n3461), .B(n3460), .Z(n3462) );
  NAND U3592 ( .A(n3463), .B(n3462), .Z(n3502) );
  NAND U3593 ( .A(b[0]), .B(a[83]), .Z(n3464) );
  XNOR U3594 ( .A(b[1]), .B(n3464), .Z(n3466) );
  NAND U3595 ( .A(n26), .B(a[82]), .Z(n3465) );
  AND U3596 ( .A(n3466), .B(n3465), .Z(n3519) );
  XOR U3597 ( .A(a[79]), .B(n42197), .Z(n3508) );
  NANDN U3598 ( .A(n3508), .B(n42173), .Z(n3469) );
  NANDN U3599 ( .A(n3467), .B(n42172), .Z(n3468) );
  NAND U3600 ( .A(n3469), .B(n3468), .Z(n3517) );
  NAND U3601 ( .A(b[7]), .B(a[75]), .Z(n3518) );
  XNOR U3602 ( .A(n3517), .B(n3518), .Z(n3520) );
  XOR U3603 ( .A(n3519), .B(n3520), .Z(n3526) );
  NANDN U3604 ( .A(n3470), .B(n42093), .Z(n3472) );
  XOR U3605 ( .A(n42134), .B(a[81]), .Z(n3511) );
  NANDN U3606 ( .A(n3511), .B(n42095), .Z(n3471) );
  NAND U3607 ( .A(n3472), .B(n3471), .Z(n3524) );
  NANDN U3608 ( .A(n3473), .B(n42231), .Z(n3475) );
  XOR U3609 ( .A(n168), .B(a[77]), .Z(n3514) );
  NANDN U3610 ( .A(n3514), .B(n42234), .Z(n3474) );
  AND U3611 ( .A(n3475), .B(n3474), .Z(n3523) );
  XNOR U3612 ( .A(n3524), .B(n3523), .Z(n3525) );
  XNOR U3613 ( .A(n3526), .B(n3525), .Z(n3530) );
  NANDN U3614 ( .A(n3477), .B(n3476), .Z(n3481) );
  NAND U3615 ( .A(n3479), .B(n3478), .Z(n3480) );
  AND U3616 ( .A(n3481), .B(n3480), .Z(n3529) );
  XOR U3617 ( .A(n3530), .B(n3529), .Z(n3531) );
  NANDN U3618 ( .A(n3483), .B(n3482), .Z(n3487) );
  NANDN U3619 ( .A(n3485), .B(n3484), .Z(n3486) );
  NAND U3620 ( .A(n3487), .B(n3486), .Z(n3532) );
  XOR U3621 ( .A(n3531), .B(n3532), .Z(n3499) );
  OR U3622 ( .A(n3489), .B(n3488), .Z(n3493) );
  NANDN U3623 ( .A(n3491), .B(n3490), .Z(n3492) );
  NAND U3624 ( .A(n3493), .B(n3492), .Z(n3500) );
  XNOR U3625 ( .A(n3499), .B(n3500), .Z(n3501) );
  XNOR U3626 ( .A(n3502), .B(n3501), .Z(n3535) );
  XNOR U3627 ( .A(n3535), .B(sreg[1099]), .Z(n3537) );
  NAND U3628 ( .A(n3494), .B(sreg[1098]), .Z(n3498) );
  OR U3629 ( .A(n3496), .B(n3495), .Z(n3497) );
  AND U3630 ( .A(n3498), .B(n3497), .Z(n3536) );
  XOR U3631 ( .A(n3537), .B(n3536), .Z(c[1099]) );
  NANDN U3632 ( .A(n3500), .B(n3499), .Z(n3504) );
  NAND U3633 ( .A(n3502), .B(n3501), .Z(n3503) );
  NAND U3634 ( .A(n3504), .B(n3503), .Z(n3543) );
  NAND U3635 ( .A(b[0]), .B(a[84]), .Z(n3505) );
  XNOR U3636 ( .A(b[1]), .B(n3505), .Z(n3507) );
  NAND U3637 ( .A(n27), .B(a[83]), .Z(n3506) );
  AND U3638 ( .A(n3507), .B(n3506), .Z(n3560) );
  XOR U3639 ( .A(a[80]), .B(n42197), .Z(n3549) );
  NANDN U3640 ( .A(n3549), .B(n42173), .Z(n3510) );
  NANDN U3641 ( .A(n3508), .B(n42172), .Z(n3509) );
  NAND U3642 ( .A(n3510), .B(n3509), .Z(n3558) );
  NAND U3643 ( .A(b[7]), .B(a[76]), .Z(n3559) );
  XNOR U3644 ( .A(n3558), .B(n3559), .Z(n3561) );
  XOR U3645 ( .A(n3560), .B(n3561), .Z(n3567) );
  NANDN U3646 ( .A(n3511), .B(n42093), .Z(n3513) );
  XOR U3647 ( .A(n42134), .B(a[82]), .Z(n3552) );
  NANDN U3648 ( .A(n3552), .B(n42095), .Z(n3512) );
  NAND U3649 ( .A(n3513), .B(n3512), .Z(n3565) );
  NANDN U3650 ( .A(n3514), .B(n42231), .Z(n3516) );
  XOR U3651 ( .A(n168), .B(a[78]), .Z(n3555) );
  NANDN U3652 ( .A(n3555), .B(n42234), .Z(n3515) );
  AND U3653 ( .A(n3516), .B(n3515), .Z(n3564) );
  XNOR U3654 ( .A(n3565), .B(n3564), .Z(n3566) );
  XNOR U3655 ( .A(n3567), .B(n3566), .Z(n3571) );
  NANDN U3656 ( .A(n3518), .B(n3517), .Z(n3522) );
  NAND U3657 ( .A(n3520), .B(n3519), .Z(n3521) );
  AND U3658 ( .A(n3522), .B(n3521), .Z(n3570) );
  XOR U3659 ( .A(n3571), .B(n3570), .Z(n3572) );
  NANDN U3660 ( .A(n3524), .B(n3523), .Z(n3528) );
  NANDN U3661 ( .A(n3526), .B(n3525), .Z(n3527) );
  NAND U3662 ( .A(n3528), .B(n3527), .Z(n3573) );
  XOR U3663 ( .A(n3572), .B(n3573), .Z(n3540) );
  OR U3664 ( .A(n3530), .B(n3529), .Z(n3534) );
  NANDN U3665 ( .A(n3532), .B(n3531), .Z(n3533) );
  NAND U3666 ( .A(n3534), .B(n3533), .Z(n3541) );
  XNOR U3667 ( .A(n3540), .B(n3541), .Z(n3542) );
  XNOR U3668 ( .A(n3543), .B(n3542), .Z(n3576) );
  XNOR U3669 ( .A(n3576), .B(sreg[1100]), .Z(n3578) );
  NAND U3670 ( .A(n3535), .B(sreg[1099]), .Z(n3539) );
  OR U3671 ( .A(n3537), .B(n3536), .Z(n3538) );
  AND U3672 ( .A(n3539), .B(n3538), .Z(n3577) );
  XOR U3673 ( .A(n3578), .B(n3577), .Z(c[1100]) );
  NANDN U3674 ( .A(n3541), .B(n3540), .Z(n3545) );
  NAND U3675 ( .A(n3543), .B(n3542), .Z(n3544) );
  NAND U3676 ( .A(n3545), .B(n3544), .Z(n3584) );
  NAND U3677 ( .A(b[0]), .B(a[85]), .Z(n3546) );
  XNOR U3678 ( .A(b[1]), .B(n3546), .Z(n3548) );
  NAND U3679 ( .A(n27), .B(a[84]), .Z(n3547) );
  AND U3680 ( .A(n3548), .B(n3547), .Z(n3601) );
  XOR U3681 ( .A(a[81]), .B(n42197), .Z(n3590) );
  NANDN U3682 ( .A(n3590), .B(n42173), .Z(n3551) );
  NANDN U3683 ( .A(n3549), .B(n42172), .Z(n3550) );
  NAND U3684 ( .A(n3551), .B(n3550), .Z(n3599) );
  NAND U3685 ( .A(b[7]), .B(a[77]), .Z(n3600) );
  XNOR U3686 ( .A(n3599), .B(n3600), .Z(n3602) );
  XOR U3687 ( .A(n3601), .B(n3602), .Z(n3608) );
  NANDN U3688 ( .A(n3552), .B(n42093), .Z(n3554) );
  XOR U3689 ( .A(n42134), .B(a[83]), .Z(n3593) );
  NANDN U3690 ( .A(n3593), .B(n42095), .Z(n3553) );
  NAND U3691 ( .A(n3554), .B(n3553), .Z(n3606) );
  NANDN U3692 ( .A(n3555), .B(n42231), .Z(n3557) );
  XOR U3693 ( .A(n168), .B(a[79]), .Z(n3596) );
  NANDN U3694 ( .A(n3596), .B(n42234), .Z(n3556) );
  AND U3695 ( .A(n3557), .B(n3556), .Z(n3605) );
  XNOR U3696 ( .A(n3606), .B(n3605), .Z(n3607) );
  XNOR U3697 ( .A(n3608), .B(n3607), .Z(n3612) );
  NANDN U3698 ( .A(n3559), .B(n3558), .Z(n3563) );
  NAND U3699 ( .A(n3561), .B(n3560), .Z(n3562) );
  AND U3700 ( .A(n3563), .B(n3562), .Z(n3611) );
  XOR U3701 ( .A(n3612), .B(n3611), .Z(n3613) );
  NANDN U3702 ( .A(n3565), .B(n3564), .Z(n3569) );
  NANDN U3703 ( .A(n3567), .B(n3566), .Z(n3568) );
  NAND U3704 ( .A(n3569), .B(n3568), .Z(n3614) );
  XOR U3705 ( .A(n3613), .B(n3614), .Z(n3581) );
  OR U3706 ( .A(n3571), .B(n3570), .Z(n3575) );
  NANDN U3707 ( .A(n3573), .B(n3572), .Z(n3574) );
  NAND U3708 ( .A(n3575), .B(n3574), .Z(n3582) );
  XNOR U3709 ( .A(n3581), .B(n3582), .Z(n3583) );
  XNOR U3710 ( .A(n3584), .B(n3583), .Z(n3617) );
  XNOR U3711 ( .A(n3617), .B(sreg[1101]), .Z(n3619) );
  NAND U3712 ( .A(n3576), .B(sreg[1100]), .Z(n3580) );
  OR U3713 ( .A(n3578), .B(n3577), .Z(n3579) );
  AND U3714 ( .A(n3580), .B(n3579), .Z(n3618) );
  XOR U3715 ( .A(n3619), .B(n3618), .Z(c[1101]) );
  NANDN U3716 ( .A(n3582), .B(n3581), .Z(n3586) );
  NAND U3717 ( .A(n3584), .B(n3583), .Z(n3585) );
  NAND U3718 ( .A(n3586), .B(n3585), .Z(n3625) );
  NAND U3719 ( .A(b[0]), .B(a[86]), .Z(n3587) );
  XNOR U3720 ( .A(b[1]), .B(n3587), .Z(n3589) );
  NAND U3721 ( .A(n27), .B(a[85]), .Z(n3588) );
  AND U3722 ( .A(n3589), .B(n3588), .Z(n3642) );
  XOR U3723 ( .A(a[82]), .B(n42197), .Z(n3631) );
  NANDN U3724 ( .A(n3631), .B(n42173), .Z(n3592) );
  NANDN U3725 ( .A(n3590), .B(n42172), .Z(n3591) );
  NAND U3726 ( .A(n3592), .B(n3591), .Z(n3640) );
  NAND U3727 ( .A(b[7]), .B(a[78]), .Z(n3641) );
  XNOR U3728 ( .A(n3640), .B(n3641), .Z(n3643) );
  XOR U3729 ( .A(n3642), .B(n3643), .Z(n3649) );
  NANDN U3730 ( .A(n3593), .B(n42093), .Z(n3595) );
  XOR U3731 ( .A(n42134), .B(a[84]), .Z(n3634) );
  NANDN U3732 ( .A(n3634), .B(n42095), .Z(n3594) );
  NAND U3733 ( .A(n3595), .B(n3594), .Z(n3647) );
  NANDN U3734 ( .A(n3596), .B(n42231), .Z(n3598) );
  XOR U3735 ( .A(n168), .B(a[80]), .Z(n3637) );
  NANDN U3736 ( .A(n3637), .B(n42234), .Z(n3597) );
  AND U3737 ( .A(n3598), .B(n3597), .Z(n3646) );
  XNOR U3738 ( .A(n3647), .B(n3646), .Z(n3648) );
  XNOR U3739 ( .A(n3649), .B(n3648), .Z(n3653) );
  NANDN U3740 ( .A(n3600), .B(n3599), .Z(n3604) );
  NAND U3741 ( .A(n3602), .B(n3601), .Z(n3603) );
  AND U3742 ( .A(n3604), .B(n3603), .Z(n3652) );
  XOR U3743 ( .A(n3653), .B(n3652), .Z(n3654) );
  NANDN U3744 ( .A(n3606), .B(n3605), .Z(n3610) );
  NANDN U3745 ( .A(n3608), .B(n3607), .Z(n3609) );
  NAND U3746 ( .A(n3610), .B(n3609), .Z(n3655) );
  XOR U3747 ( .A(n3654), .B(n3655), .Z(n3622) );
  OR U3748 ( .A(n3612), .B(n3611), .Z(n3616) );
  NANDN U3749 ( .A(n3614), .B(n3613), .Z(n3615) );
  NAND U3750 ( .A(n3616), .B(n3615), .Z(n3623) );
  XNOR U3751 ( .A(n3622), .B(n3623), .Z(n3624) );
  XNOR U3752 ( .A(n3625), .B(n3624), .Z(n3658) );
  XNOR U3753 ( .A(n3658), .B(sreg[1102]), .Z(n3660) );
  NAND U3754 ( .A(n3617), .B(sreg[1101]), .Z(n3621) );
  OR U3755 ( .A(n3619), .B(n3618), .Z(n3620) );
  AND U3756 ( .A(n3621), .B(n3620), .Z(n3659) );
  XOR U3757 ( .A(n3660), .B(n3659), .Z(c[1102]) );
  NANDN U3758 ( .A(n3623), .B(n3622), .Z(n3627) );
  NAND U3759 ( .A(n3625), .B(n3624), .Z(n3626) );
  NAND U3760 ( .A(n3627), .B(n3626), .Z(n3666) );
  NAND U3761 ( .A(b[0]), .B(a[87]), .Z(n3628) );
  XNOR U3762 ( .A(b[1]), .B(n3628), .Z(n3630) );
  NAND U3763 ( .A(n27), .B(a[86]), .Z(n3629) );
  AND U3764 ( .A(n3630), .B(n3629), .Z(n3683) );
  XOR U3765 ( .A(a[83]), .B(n42197), .Z(n3672) );
  NANDN U3766 ( .A(n3672), .B(n42173), .Z(n3633) );
  NANDN U3767 ( .A(n3631), .B(n42172), .Z(n3632) );
  NAND U3768 ( .A(n3633), .B(n3632), .Z(n3681) );
  NAND U3769 ( .A(b[7]), .B(a[79]), .Z(n3682) );
  XNOR U3770 ( .A(n3681), .B(n3682), .Z(n3684) );
  XOR U3771 ( .A(n3683), .B(n3684), .Z(n3690) );
  NANDN U3772 ( .A(n3634), .B(n42093), .Z(n3636) );
  XOR U3773 ( .A(n42134), .B(a[85]), .Z(n3675) );
  NANDN U3774 ( .A(n3675), .B(n42095), .Z(n3635) );
  NAND U3775 ( .A(n3636), .B(n3635), .Z(n3688) );
  NANDN U3776 ( .A(n3637), .B(n42231), .Z(n3639) );
  XOR U3777 ( .A(n168), .B(a[81]), .Z(n3678) );
  NANDN U3778 ( .A(n3678), .B(n42234), .Z(n3638) );
  AND U3779 ( .A(n3639), .B(n3638), .Z(n3687) );
  XNOR U3780 ( .A(n3688), .B(n3687), .Z(n3689) );
  XNOR U3781 ( .A(n3690), .B(n3689), .Z(n3694) );
  NANDN U3782 ( .A(n3641), .B(n3640), .Z(n3645) );
  NAND U3783 ( .A(n3643), .B(n3642), .Z(n3644) );
  AND U3784 ( .A(n3645), .B(n3644), .Z(n3693) );
  XOR U3785 ( .A(n3694), .B(n3693), .Z(n3695) );
  NANDN U3786 ( .A(n3647), .B(n3646), .Z(n3651) );
  NANDN U3787 ( .A(n3649), .B(n3648), .Z(n3650) );
  NAND U3788 ( .A(n3651), .B(n3650), .Z(n3696) );
  XOR U3789 ( .A(n3695), .B(n3696), .Z(n3663) );
  OR U3790 ( .A(n3653), .B(n3652), .Z(n3657) );
  NANDN U3791 ( .A(n3655), .B(n3654), .Z(n3656) );
  NAND U3792 ( .A(n3657), .B(n3656), .Z(n3664) );
  XNOR U3793 ( .A(n3663), .B(n3664), .Z(n3665) );
  XNOR U3794 ( .A(n3666), .B(n3665), .Z(n3699) );
  XNOR U3795 ( .A(n3699), .B(sreg[1103]), .Z(n3701) );
  NAND U3796 ( .A(n3658), .B(sreg[1102]), .Z(n3662) );
  OR U3797 ( .A(n3660), .B(n3659), .Z(n3661) );
  AND U3798 ( .A(n3662), .B(n3661), .Z(n3700) );
  XOR U3799 ( .A(n3701), .B(n3700), .Z(c[1103]) );
  NANDN U3800 ( .A(n3664), .B(n3663), .Z(n3668) );
  NAND U3801 ( .A(n3666), .B(n3665), .Z(n3667) );
  NAND U3802 ( .A(n3668), .B(n3667), .Z(n3707) );
  NAND U3803 ( .A(b[0]), .B(a[88]), .Z(n3669) );
  XNOR U3804 ( .A(b[1]), .B(n3669), .Z(n3671) );
  NAND U3805 ( .A(n27), .B(a[87]), .Z(n3670) );
  AND U3806 ( .A(n3671), .B(n3670), .Z(n3724) );
  XOR U3807 ( .A(a[84]), .B(n42197), .Z(n3713) );
  NANDN U3808 ( .A(n3713), .B(n42173), .Z(n3674) );
  NANDN U3809 ( .A(n3672), .B(n42172), .Z(n3673) );
  NAND U3810 ( .A(n3674), .B(n3673), .Z(n3722) );
  NAND U3811 ( .A(b[7]), .B(a[80]), .Z(n3723) );
  XNOR U3812 ( .A(n3722), .B(n3723), .Z(n3725) );
  XOR U3813 ( .A(n3724), .B(n3725), .Z(n3731) );
  NANDN U3814 ( .A(n3675), .B(n42093), .Z(n3677) );
  XOR U3815 ( .A(n42134), .B(a[86]), .Z(n3716) );
  NANDN U3816 ( .A(n3716), .B(n42095), .Z(n3676) );
  NAND U3817 ( .A(n3677), .B(n3676), .Z(n3729) );
  NANDN U3818 ( .A(n3678), .B(n42231), .Z(n3680) );
  XOR U3819 ( .A(n168), .B(a[82]), .Z(n3719) );
  NANDN U3820 ( .A(n3719), .B(n42234), .Z(n3679) );
  AND U3821 ( .A(n3680), .B(n3679), .Z(n3728) );
  XNOR U3822 ( .A(n3729), .B(n3728), .Z(n3730) );
  XNOR U3823 ( .A(n3731), .B(n3730), .Z(n3735) );
  NANDN U3824 ( .A(n3682), .B(n3681), .Z(n3686) );
  NAND U3825 ( .A(n3684), .B(n3683), .Z(n3685) );
  AND U3826 ( .A(n3686), .B(n3685), .Z(n3734) );
  XOR U3827 ( .A(n3735), .B(n3734), .Z(n3736) );
  NANDN U3828 ( .A(n3688), .B(n3687), .Z(n3692) );
  NANDN U3829 ( .A(n3690), .B(n3689), .Z(n3691) );
  NAND U3830 ( .A(n3692), .B(n3691), .Z(n3737) );
  XOR U3831 ( .A(n3736), .B(n3737), .Z(n3704) );
  OR U3832 ( .A(n3694), .B(n3693), .Z(n3698) );
  NANDN U3833 ( .A(n3696), .B(n3695), .Z(n3697) );
  NAND U3834 ( .A(n3698), .B(n3697), .Z(n3705) );
  XNOR U3835 ( .A(n3704), .B(n3705), .Z(n3706) );
  XNOR U3836 ( .A(n3707), .B(n3706), .Z(n3740) );
  XNOR U3837 ( .A(n3740), .B(sreg[1104]), .Z(n3742) );
  NAND U3838 ( .A(n3699), .B(sreg[1103]), .Z(n3703) );
  OR U3839 ( .A(n3701), .B(n3700), .Z(n3702) );
  AND U3840 ( .A(n3703), .B(n3702), .Z(n3741) );
  XOR U3841 ( .A(n3742), .B(n3741), .Z(c[1104]) );
  NANDN U3842 ( .A(n3705), .B(n3704), .Z(n3709) );
  NAND U3843 ( .A(n3707), .B(n3706), .Z(n3708) );
  NAND U3844 ( .A(n3709), .B(n3708), .Z(n3748) );
  NAND U3845 ( .A(b[0]), .B(a[89]), .Z(n3710) );
  XNOR U3846 ( .A(b[1]), .B(n3710), .Z(n3712) );
  NAND U3847 ( .A(n27), .B(a[88]), .Z(n3711) );
  AND U3848 ( .A(n3712), .B(n3711), .Z(n3765) );
  XOR U3849 ( .A(a[85]), .B(n42197), .Z(n3754) );
  NANDN U3850 ( .A(n3754), .B(n42173), .Z(n3715) );
  NANDN U3851 ( .A(n3713), .B(n42172), .Z(n3714) );
  NAND U3852 ( .A(n3715), .B(n3714), .Z(n3763) );
  NAND U3853 ( .A(b[7]), .B(a[81]), .Z(n3764) );
  XNOR U3854 ( .A(n3763), .B(n3764), .Z(n3766) );
  XOR U3855 ( .A(n3765), .B(n3766), .Z(n3772) );
  NANDN U3856 ( .A(n3716), .B(n42093), .Z(n3718) );
  XOR U3857 ( .A(n42134), .B(a[87]), .Z(n3757) );
  NANDN U3858 ( .A(n3757), .B(n42095), .Z(n3717) );
  NAND U3859 ( .A(n3718), .B(n3717), .Z(n3770) );
  NANDN U3860 ( .A(n3719), .B(n42231), .Z(n3721) );
  XOR U3861 ( .A(n169), .B(a[83]), .Z(n3760) );
  NANDN U3862 ( .A(n3760), .B(n42234), .Z(n3720) );
  AND U3863 ( .A(n3721), .B(n3720), .Z(n3769) );
  XNOR U3864 ( .A(n3770), .B(n3769), .Z(n3771) );
  XNOR U3865 ( .A(n3772), .B(n3771), .Z(n3776) );
  NANDN U3866 ( .A(n3723), .B(n3722), .Z(n3727) );
  NAND U3867 ( .A(n3725), .B(n3724), .Z(n3726) );
  AND U3868 ( .A(n3727), .B(n3726), .Z(n3775) );
  XOR U3869 ( .A(n3776), .B(n3775), .Z(n3777) );
  NANDN U3870 ( .A(n3729), .B(n3728), .Z(n3733) );
  NANDN U3871 ( .A(n3731), .B(n3730), .Z(n3732) );
  NAND U3872 ( .A(n3733), .B(n3732), .Z(n3778) );
  XOR U3873 ( .A(n3777), .B(n3778), .Z(n3745) );
  OR U3874 ( .A(n3735), .B(n3734), .Z(n3739) );
  NANDN U3875 ( .A(n3737), .B(n3736), .Z(n3738) );
  NAND U3876 ( .A(n3739), .B(n3738), .Z(n3746) );
  XNOR U3877 ( .A(n3745), .B(n3746), .Z(n3747) );
  XNOR U3878 ( .A(n3748), .B(n3747), .Z(n3781) );
  XNOR U3879 ( .A(n3781), .B(sreg[1105]), .Z(n3783) );
  NAND U3880 ( .A(n3740), .B(sreg[1104]), .Z(n3744) );
  OR U3881 ( .A(n3742), .B(n3741), .Z(n3743) );
  AND U3882 ( .A(n3744), .B(n3743), .Z(n3782) );
  XOR U3883 ( .A(n3783), .B(n3782), .Z(c[1105]) );
  NANDN U3884 ( .A(n3746), .B(n3745), .Z(n3750) );
  NAND U3885 ( .A(n3748), .B(n3747), .Z(n3749) );
  NAND U3886 ( .A(n3750), .B(n3749), .Z(n3789) );
  NAND U3887 ( .A(b[0]), .B(a[90]), .Z(n3751) );
  XNOR U3888 ( .A(b[1]), .B(n3751), .Z(n3753) );
  NAND U3889 ( .A(n27), .B(a[89]), .Z(n3752) );
  AND U3890 ( .A(n3753), .B(n3752), .Z(n3806) );
  XOR U3891 ( .A(a[86]), .B(n42197), .Z(n3795) );
  NANDN U3892 ( .A(n3795), .B(n42173), .Z(n3756) );
  NANDN U3893 ( .A(n3754), .B(n42172), .Z(n3755) );
  NAND U3894 ( .A(n3756), .B(n3755), .Z(n3804) );
  NAND U3895 ( .A(b[7]), .B(a[82]), .Z(n3805) );
  XNOR U3896 ( .A(n3804), .B(n3805), .Z(n3807) );
  XOR U3897 ( .A(n3806), .B(n3807), .Z(n3813) );
  NANDN U3898 ( .A(n3757), .B(n42093), .Z(n3759) );
  XOR U3899 ( .A(n42134), .B(a[88]), .Z(n3798) );
  NANDN U3900 ( .A(n3798), .B(n42095), .Z(n3758) );
  NAND U3901 ( .A(n3759), .B(n3758), .Z(n3811) );
  NANDN U3902 ( .A(n3760), .B(n42231), .Z(n3762) );
  XOR U3903 ( .A(n169), .B(a[84]), .Z(n3801) );
  NANDN U3904 ( .A(n3801), .B(n42234), .Z(n3761) );
  AND U3905 ( .A(n3762), .B(n3761), .Z(n3810) );
  XNOR U3906 ( .A(n3811), .B(n3810), .Z(n3812) );
  XNOR U3907 ( .A(n3813), .B(n3812), .Z(n3817) );
  NANDN U3908 ( .A(n3764), .B(n3763), .Z(n3768) );
  NAND U3909 ( .A(n3766), .B(n3765), .Z(n3767) );
  AND U3910 ( .A(n3768), .B(n3767), .Z(n3816) );
  XOR U3911 ( .A(n3817), .B(n3816), .Z(n3818) );
  NANDN U3912 ( .A(n3770), .B(n3769), .Z(n3774) );
  NANDN U3913 ( .A(n3772), .B(n3771), .Z(n3773) );
  NAND U3914 ( .A(n3774), .B(n3773), .Z(n3819) );
  XOR U3915 ( .A(n3818), .B(n3819), .Z(n3786) );
  OR U3916 ( .A(n3776), .B(n3775), .Z(n3780) );
  NANDN U3917 ( .A(n3778), .B(n3777), .Z(n3779) );
  NAND U3918 ( .A(n3780), .B(n3779), .Z(n3787) );
  XNOR U3919 ( .A(n3786), .B(n3787), .Z(n3788) );
  XNOR U3920 ( .A(n3789), .B(n3788), .Z(n3822) );
  XNOR U3921 ( .A(n3822), .B(sreg[1106]), .Z(n3824) );
  NAND U3922 ( .A(n3781), .B(sreg[1105]), .Z(n3785) );
  OR U3923 ( .A(n3783), .B(n3782), .Z(n3784) );
  AND U3924 ( .A(n3785), .B(n3784), .Z(n3823) );
  XOR U3925 ( .A(n3824), .B(n3823), .Z(c[1106]) );
  NANDN U3926 ( .A(n3787), .B(n3786), .Z(n3791) );
  NAND U3927 ( .A(n3789), .B(n3788), .Z(n3790) );
  NAND U3928 ( .A(n3791), .B(n3790), .Z(n3830) );
  NAND U3929 ( .A(b[0]), .B(a[91]), .Z(n3792) );
  XNOR U3930 ( .A(b[1]), .B(n3792), .Z(n3794) );
  NAND U3931 ( .A(n28), .B(a[90]), .Z(n3793) );
  AND U3932 ( .A(n3794), .B(n3793), .Z(n3847) );
  XOR U3933 ( .A(a[87]), .B(n42197), .Z(n3836) );
  NANDN U3934 ( .A(n3836), .B(n42173), .Z(n3797) );
  NANDN U3935 ( .A(n3795), .B(n42172), .Z(n3796) );
  NAND U3936 ( .A(n3797), .B(n3796), .Z(n3845) );
  NAND U3937 ( .A(b[7]), .B(a[83]), .Z(n3846) );
  XNOR U3938 ( .A(n3845), .B(n3846), .Z(n3848) );
  XOR U3939 ( .A(n3847), .B(n3848), .Z(n3854) );
  NANDN U3940 ( .A(n3798), .B(n42093), .Z(n3800) );
  XOR U3941 ( .A(n42134), .B(a[89]), .Z(n3839) );
  NANDN U3942 ( .A(n3839), .B(n42095), .Z(n3799) );
  NAND U3943 ( .A(n3800), .B(n3799), .Z(n3852) );
  NANDN U3944 ( .A(n3801), .B(n42231), .Z(n3803) );
  XOR U3945 ( .A(n169), .B(a[85]), .Z(n3842) );
  NANDN U3946 ( .A(n3842), .B(n42234), .Z(n3802) );
  AND U3947 ( .A(n3803), .B(n3802), .Z(n3851) );
  XNOR U3948 ( .A(n3852), .B(n3851), .Z(n3853) );
  XNOR U3949 ( .A(n3854), .B(n3853), .Z(n3858) );
  NANDN U3950 ( .A(n3805), .B(n3804), .Z(n3809) );
  NAND U3951 ( .A(n3807), .B(n3806), .Z(n3808) );
  AND U3952 ( .A(n3809), .B(n3808), .Z(n3857) );
  XOR U3953 ( .A(n3858), .B(n3857), .Z(n3859) );
  NANDN U3954 ( .A(n3811), .B(n3810), .Z(n3815) );
  NANDN U3955 ( .A(n3813), .B(n3812), .Z(n3814) );
  NAND U3956 ( .A(n3815), .B(n3814), .Z(n3860) );
  XOR U3957 ( .A(n3859), .B(n3860), .Z(n3827) );
  OR U3958 ( .A(n3817), .B(n3816), .Z(n3821) );
  NANDN U3959 ( .A(n3819), .B(n3818), .Z(n3820) );
  NAND U3960 ( .A(n3821), .B(n3820), .Z(n3828) );
  XNOR U3961 ( .A(n3827), .B(n3828), .Z(n3829) );
  XNOR U3962 ( .A(n3830), .B(n3829), .Z(n3863) );
  XNOR U3963 ( .A(n3863), .B(sreg[1107]), .Z(n3865) );
  NAND U3964 ( .A(n3822), .B(sreg[1106]), .Z(n3826) );
  OR U3965 ( .A(n3824), .B(n3823), .Z(n3825) );
  AND U3966 ( .A(n3826), .B(n3825), .Z(n3864) );
  XOR U3967 ( .A(n3865), .B(n3864), .Z(c[1107]) );
  NANDN U3968 ( .A(n3828), .B(n3827), .Z(n3832) );
  NAND U3969 ( .A(n3830), .B(n3829), .Z(n3831) );
  NAND U3970 ( .A(n3832), .B(n3831), .Z(n3871) );
  NAND U3971 ( .A(b[0]), .B(a[92]), .Z(n3833) );
  XNOR U3972 ( .A(b[1]), .B(n3833), .Z(n3835) );
  NAND U3973 ( .A(n28), .B(a[91]), .Z(n3834) );
  AND U3974 ( .A(n3835), .B(n3834), .Z(n3888) );
  XOR U3975 ( .A(a[88]), .B(n42197), .Z(n3877) );
  NANDN U3976 ( .A(n3877), .B(n42173), .Z(n3838) );
  NANDN U3977 ( .A(n3836), .B(n42172), .Z(n3837) );
  NAND U3978 ( .A(n3838), .B(n3837), .Z(n3886) );
  NAND U3979 ( .A(b[7]), .B(a[84]), .Z(n3887) );
  XNOR U3980 ( .A(n3886), .B(n3887), .Z(n3889) );
  XOR U3981 ( .A(n3888), .B(n3889), .Z(n3895) );
  NANDN U3982 ( .A(n3839), .B(n42093), .Z(n3841) );
  XOR U3983 ( .A(n42134), .B(a[90]), .Z(n3880) );
  NANDN U3984 ( .A(n3880), .B(n42095), .Z(n3840) );
  NAND U3985 ( .A(n3841), .B(n3840), .Z(n3893) );
  NANDN U3986 ( .A(n3842), .B(n42231), .Z(n3844) );
  XOR U3987 ( .A(n169), .B(a[86]), .Z(n3883) );
  NANDN U3988 ( .A(n3883), .B(n42234), .Z(n3843) );
  AND U3989 ( .A(n3844), .B(n3843), .Z(n3892) );
  XNOR U3990 ( .A(n3893), .B(n3892), .Z(n3894) );
  XNOR U3991 ( .A(n3895), .B(n3894), .Z(n3899) );
  NANDN U3992 ( .A(n3846), .B(n3845), .Z(n3850) );
  NAND U3993 ( .A(n3848), .B(n3847), .Z(n3849) );
  AND U3994 ( .A(n3850), .B(n3849), .Z(n3898) );
  XOR U3995 ( .A(n3899), .B(n3898), .Z(n3900) );
  NANDN U3996 ( .A(n3852), .B(n3851), .Z(n3856) );
  NANDN U3997 ( .A(n3854), .B(n3853), .Z(n3855) );
  NAND U3998 ( .A(n3856), .B(n3855), .Z(n3901) );
  XOR U3999 ( .A(n3900), .B(n3901), .Z(n3868) );
  OR U4000 ( .A(n3858), .B(n3857), .Z(n3862) );
  NANDN U4001 ( .A(n3860), .B(n3859), .Z(n3861) );
  NAND U4002 ( .A(n3862), .B(n3861), .Z(n3869) );
  XNOR U4003 ( .A(n3868), .B(n3869), .Z(n3870) );
  XNOR U4004 ( .A(n3871), .B(n3870), .Z(n3904) );
  XNOR U4005 ( .A(n3904), .B(sreg[1108]), .Z(n3906) );
  NAND U4006 ( .A(n3863), .B(sreg[1107]), .Z(n3867) );
  OR U4007 ( .A(n3865), .B(n3864), .Z(n3866) );
  AND U4008 ( .A(n3867), .B(n3866), .Z(n3905) );
  XOR U4009 ( .A(n3906), .B(n3905), .Z(c[1108]) );
  NANDN U4010 ( .A(n3869), .B(n3868), .Z(n3873) );
  NAND U4011 ( .A(n3871), .B(n3870), .Z(n3872) );
  NAND U4012 ( .A(n3873), .B(n3872), .Z(n3912) );
  NAND U4013 ( .A(b[0]), .B(a[93]), .Z(n3874) );
  XNOR U4014 ( .A(b[1]), .B(n3874), .Z(n3876) );
  NAND U4015 ( .A(n28), .B(a[92]), .Z(n3875) );
  AND U4016 ( .A(n3876), .B(n3875), .Z(n3929) );
  XOR U4017 ( .A(a[89]), .B(n42197), .Z(n3918) );
  NANDN U4018 ( .A(n3918), .B(n42173), .Z(n3879) );
  NANDN U4019 ( .A(n3877), .B(n42172), .Z(n3878) );
  NAND U4020 ( .A(n3879), .B(n3878), .Z(n3927) );
  NAND U4021 ( .A(b[7]), .B(a[85]), .Z(n3928) );
  XNOR U4022 ( .A(n3927), .B(n3928), .Z(n3930) );
  XOR U4023 ( .A(n3929), .B(n3930), .Z(n3936) );
  NANDN U4024 ( .A(n3880), .B(n42093), .Z(n3882) );
  XOR U4025 ( .A(n42134), .B(a[91]), .Z(n3921) );
  NANDN U4026 ( .A(n3921), .B(n42095), .Z(n3881) );
  NAND U4027 ( .A(n3882), .B(n3881), .Z(n3934) );
  NANDN U4028 ( .A(n3883), .B(n42231), .Z(n3885) );
  XOR U4029 ( .A(n169), .B(a[87]), .Z(n3924) );
  NANDN U4030 ( .A(n3924), .B(n42234), .Z(n3884) );
  AND U4031 ( .A(n3885), .B(n3884), .Z(n3933) );
  XNOR U4032 ( .A(n3934), .B(n3933), .Z(n3935) );
  XNOR U4033 ( .A(n3936), .B(n3935), .Z(n3940) );
  NANDN U4034 ( .A(n3887), .B(n3886), .Z(n3891) );
  NAND U4035 ( .A(n3889), .B(n3888), .Z(n3890) );
  AND U4036 ( .A(n3891), .B(n3890), .Z(n3939) );
  XOR U4037 ( .A(n3940), .B(n3939), .Z(n3941) );
  NANDN U4038 ( .A(n3893), .B(n3892), .Z(n3897) );
  NANDN U4039 ( .A(n3895), .B(n3894), .Z(n3896) );
  NAND U4040 ( .A(n3897), .B(n3896), .Z(n3942) );
  XOR U4041 ( .A(n3941), .B(n3942), .Z(n3909) );
  OR U4042 ( .A(n3899), .B(n3898), .Z(n3903) );
  NANDN U4043 ( .A(n3901), .B(n3900), .Z(n3902) );
  NAND U4044 ( .A(n3903), .B(n3902), .Z(n3910) );
  XNOR U4045 ( .A(n3909), .B(n3910), .Z(n3911) );
  XNOR U4046 ( .A(n3912), .B(n3911), .Z(n3945) );
  XNOR U4047 ( .A(n3945), .B(sreg[1109]), .Z(n3947) );
  NAND U4048 ( .A(n3904), .B(sreg[1108]), .Z(n3908) );
  OR U4049 ( .A(n3906), .B(n3905), .Z(n3907) );
  AND U4050 ( .A(n3908), .B(n3907), .Z(n3946) );
  XOR U4051 ( .A(n3947), .B(n3946), .Z(c[1109]) );
  NANDN U4052 ( .A(n3910), .B(n3909), .Z(n3914) );
  NAND U4053 ( .A(n3912), .B(n3911), .Z(n3913) );
  NAND U4054 ( .A(n3914), .B(n3913), .Z(n3953) );
  NAND U4055 ( .A(b[0]), .B(a[94]), .Z(n3915) );
  XNOR U4056 ( .A(b[1]), .B(n3915), .Z(n3917) );
  NAND U4057 ( .A(n28), .B(a[93]), .Z(n3916) );
  AND U4058 ( .A(n3917), .B(n3916), .Z(n3970) );
  XOR U4059 ( .A(a[90]), .B(n42197), .Z(n3959) );
  NANDN U4060 ( .A(n3959), .B(n42173), .Z(n3920) );
  NANDN U4061 ( .A(n3918), .B(n42172), .Z(n3919) );
  NAND U4062 ( .A(n3920), .B(n3919), .Z(n3968) );
  NAND U4063 ( .A(b[7]), .B(a[86]), .Z(n3969) );
  XNOR U4064 ( .A(n3968), .B(n3969), .Z(n3971) );
  XOR U4065 ( .A(n3970), .B(n3971), .Z(n3977) );
  NANDN U4066 ( .A(n3921), .B(n42093), .Z(n3923) );
  XOR U4067 ( .A(n42134), .B(a[92]), .Z(n3962) );
  NANDN U4068 ( .A(n3962), .B(n42095), .Z(n3922) );
  NAND U4069 ( .A(n3923), .B(n3922), .Z(n3975) );
  NANDN U4070 ( .A(n3924), .B(n42231), .Z(n3926) );
  XOR U4071 ( .A(n169), .B(a[88]), .Z(n3965) );
  NANDN U4072 ( .A(n3965), .B(n42234), .Z(n3925) );
  AND U4073 ( .A(n3926), .B(n3925), .Z(n3974) );
  XNOR U4074 ( .A(n3975), .B(n3974), .Z(n3976) );
  XNOR U4075 ( .A(n3977), .B(n3976), .Z(n3981) );
  NANDN U4076 ( .A(n3928), .B(n3927), .Z(n3932) );
  NAND U4077 ( .A(n3930), .B(n3929), .Z(n3931) );
  AND U4078 ( .A(n3932), .B(n3931), .Z(n3980) );
  XOR U4079 ( .A(n3981), .B(n3980), .Z(n3982) );
  NANDN U4080 ( .A(n3934), .B(n3933), .Z(n3938) );
  NANDN U4081 ( .A(n3936), .B(n3935), .Z(n3937) );
  NAND U4082 ( .A(n3938), .B(n3937), .Z(n3983) );
  XOR U4083 ( .A(n3982), .B(n3983), .Z(n3950) );
  OR U4084 ( .A(n3940), .B(n3939), .Z(n3944) );
  NANDN U4085 ( .A(n3942), .B(n3941), .Z(n3943) );
  NAND U4086 ( .A(n3944), .B(n3943), .Z(n3951) );
  XNOR U4087 ( .A(n3950), .B(n3951), .Z(n3952) );
  XNOR U4088 ( .A(n3953), .B(n3952), .Z(n3986) );
  XNOR U4089 ( .A(n3986), .B(sreg[1110]), .Z(n3988) );
  NAND U4090 ( .A(n3945), .B(sreg[1109]), .Z(n3949) );
  OR U4091 ( .A(n3947), .B(n3946), .Z(n3948) );
  AND U4092 ( .A(n3949), .B(n3948), .Z(n3987) );
  XOR U4093 ( .A(n3988), .B(n3987), .Z(c[1110]) );
  NANDN U4094 ( .A(n3951), .B(n3950), .Z(n3955) );
  NAND U4095 ( .A(n3953), .B(n3952), .Z(n3954) );
  NAND U4096 ( .A(n3955), .B(n3954), .Z(n3994) );
  NAND U4097 ( .A(b[0]), .B(a[95]), .Z(n3956) );
  XNOR U4098 ( .A(b[1]), .B(n3956), .Z(n3958) );
  NAND U4099 ( .A(n28), .B(a[94]), .Z(n3957) );
  AND U4100 ( .A(n3958), .B(n3957), .Z(n4011) );
  XOR U4101 ( .A(a[91]), .B(n42197), .Z(n4000) );
  NANDN U4102 ( .A(n4000), .B(n42173), .Z(n3961) );
  NANDN U4103 ( .A(n3959), .B(n42172), .Z(n3960) );
  NAND U4104 ( .A(n3961), .B(n3960), .Z(n4009) );
  NAND U4105 ( .A(b[7]), .B(a[87]), .Z(n4010) );
  XNOR U4106 ( .A(n4009), .B(n4010), .Z(n4012) );
  XOR U4107 ( .A(n4011), .B(n4012), .Z(n4018) );
  NANDN U4108 ( .A(n3962), .B(n42093), .Z(n3964) );
  XOR U4109 ( .A(n42134), .B(a[93]), .Z(n4003) );
  NANDN U4110 ( .A(n4003), .B(n42095), .Z(n3963) );
  NAND U4111 ( .A(n3964), .B(n3963), .Z(n4016) );
  NANDN U4112 ( .A(n3965), .B(n42231), .Z(n3967) );
  XOR U4113 ( .A(n169), .B(a[89]), .Z(n4006) );
  NANDN U4114 ( .A(n4006), .B(n42234), .Z(n3966) );
  AND U4115 ( .A(n3967), .B(n3966), .Z(n4015) );
  XNOR U4116 ( .A(n4016), .B(n4015), .Z(n4017) );
  XNOR U4117 ( .A(n4018), .B(n4017), .Z(n4022) );
  NANDN U4118 ( .A(n3969), .B(n3968), .Z(n3973) );
  NAND U4119 ( .A(n3971), .B(n3970), .Z(n3972) );
  AND U4120 ( .A(n3973), .B(n3972), .Z(n4021) );
  XOR U4121 ( .A(n4022), .B(n4021), .Z(n4023) );
  NANDN U4122 ( .A(n3975), .B(n3974), .Z(n3979) );
  NANDN U4123 ( .A(n3977), .B(n3976), .Z(n3978) );
  NAND U4124 ( .A(n3979), .B(n3978), .Z(n4024) );
  XOR U4125 ( .A(n4023), .B(n4024), .Z(n3991) );
  OR U4126 ( .A(n3981), .B(n3980), .Z(n3985) );
  NANDN U4127 ( .A(n3983), .B(n3982), .Z(n3984) );
  NAND U4128 ( .A(n3985), .B(n3984), .Z(n3992) );
  XNOR U4129 ( .A(n3991), .B(n3992), .Z(n3993) );
  XNOR U4130 ( .A(n3994), .B(n3993), .Z(n4027) );
  XNOR U4131 ( .A(n4027), .B(sreg[1111]), .Z(n4029) );
  NAND U4132 ( .A(n3986), .B(sreg[1110]), .Z(n3990) );
  OR U4133 ( .A(n3988), .B(n3987), .Z(n3989) );
  AND U4134 ( .A(n3990), .B(n3989), .Z(n4028) );
  XOR U4135 ( .A(n4029), .B(n4028), .Z(c[1111]) );
  NANDN U4136 ( .A(n3992), .B(n3991), .Z(n3996) );
  NAND U4137 ( .A(n3994), .B(n3993), .Z(n3995) );
  NAND U4138 ( .A(n3996), .B(n3995), .Z(n4035) );
  NAND U4139 ( .A(b[0]), .B(a[96]), .Z(n3997) );
  XNOR U4140 ( .A(b[1]), .B(n3997), .Z(n3999) );
  NAND U4141 ( .A(n28), .B(a[95]), .Z(n3998) );
  AND U4142 ( .A(n3999), .B(n3998), .Z(n4052) );
  XOR U4143 ( .A(a[92]), .B(n42197), .Z(n4041) );
  NANDN U4144 ( .A(n4041), .B(n42173), .Z(n4002) );
  NANDN U4145 ( .A(n4000), .B(n42172), .Z(n4001) );
  NAND U4146 ( .A(n4002), .B(n4001), .Z(n4050) );
  NAND U4147 ( .A(b[7]), .B(a[88]), .Z(n4051) );
  XNOR U4148 ( .A(n4050), .B(n4051), .Z(n4053) );
  XOR U4149 ( .A(n4052), .B(n4053), .Z(n4059) );
  NANDN U4150 ( .A(n4003), .B(n42093), .Z(n4005) );
  XOR U4151 ( .A(n42134), .B(a[94]), .Z(n4044) );
  NANDN U4152 ( .A(n4044), .B(n42095), .Z(n4004) );
  NAND U4153 ( .A(n4005), .B(n4004), .Z(n4057) );
  NANDN U4154 ( .A(n4006), .B(n42231), .Z(n4008) );
  XOR U4155 ( .A(n169), .B(a[90]), .Z(n4047) );
  NANDN U4156 ( .A(n4047), .B(n42234), .Z(n4007) );
  AND U4157 ( .A(n4008), .B(n4007), .Z(n4056) );
  XNOR U4158 ( .A(n4057), .B(n4056), .Z(n4058) );
  XNOR U4159 ( .A(n4059), .B(n4058), .Z(n4063) );
  NANDN U4160 ( .A(n4010), .B(n4009), .Z(n4014) );
  NAND U4161 ( .A(n4012), .B(n4011), .Z(n4013) );
  AND U4162 ( .A(n4014), .B(n4013), .Z(n4062) );
  XOR U4163 ( .A(n4063), .B(n4062), .Z(n4064) );
  NANDN U4164 ( .A(n4016), .B(n4015), .Z(n4020) );
  NANDN U4165 ( .A(n4018), .B(n4017), .Z(n4019) );
  NAND U4166 ( .A(n4020), .B(n4019), .Z(n4065) );
  XOR U4167 ( .A(n4064), .B(n4065), .Z(n4032) );
  OR U4168 ( .A(n4022), .B(n4021), .Z(n4026) );
  NANDN U4169 ( .A(n4024), .B(n4023), .Z(n4025) );
  NAND U4170 ( .A(n4026), .B(n4025), .Z(n4033) );
  XNOR U4171 ( .A(n4032), .B(n4033), .Z(n4034) );
  XNOR U4172 ( .A(n4035), .B(n4034), .Z(n4068) );
  XNOR U4173 ( .A(n4068), .B(sreg[1112]), .Z(n4070) );
  NAND U4174 ( .A(n4027), .B(sreg[1111]), .Z(n4031) );
  OR U4175 ( .A(n4029), .B(n4028), .Z(n4030) );
  AND U4176 ( .A(n4031), .B(n4030), .Z(n4069) );
  XOR U4177 ( .A(n4070), .B(n4069), .Z(c[1112]) );
  NANDN U4178 ( .A(n4033), .B(n4032), .Z(n4037) );
  NAND U4179 ( .A(n4035), .B(n4034), .Z(n4036) );
  NAND U4180 ( .A(n4037), .B(n4036), .Z(n4076) );
  NAND U4181 ( .A(b[0]), .B(a[97]), .Z(n4038) );
  XNOR U4182 ( .A(b[1]), .B(n4038), .Z(n4040) );
  NAND U4183 ( .A(n28), .B(a[96]), .Z(n4039) );
  AND U4184 ( .A(n4040), .B(n4039), .Z(n4093) );
  XOR U4185 ( .A(a[93]), .B(n42197), .Z(n4082) );
  NANDN U4186 ( .A(n4082), .B(n42173), .Z(n4043) );
  NANDN U4187 ( .A(n4041), .B(n42172), .Z(n4042) );
  NAND U4188 ( .A(n4043), .B(n4042), .Z(n4091) );
  NAND U4189 ( .A(b[7]), .B(a[89]), .Z(n4092) );
  XNOR U4190 ( .A(n4091), .B(n4092), .Z(n4094) );
  XOR U4191 ( .A(n4093), .B(n4094), .Z(n4100) );
  NANDN U4192 ( .A(n4044), .B(n42093), .Z(n4046) );
  XOR U4193 ( .A(n42134), .B(a[95]), .Z(n4085) );
  NANDN U4194 ( .A(n4085), .B(n42095), .Z(n4045) );
  NAND U4195 ( .A(n4046), .B(n4045), .Z(n4098) );
  NANDN U4196 ( .A(n4047), .B(n42231), .Z(n4049) );
  XOR U4197 ( .A(n169), .B(a[91]), .Z(n4088) );
  NANDN U4198 ( .A(n4088), .B(n42234), .Z(n4048) );
  AND U4199 ( .A(n4049), .B(n4048), .Z(n4097) );
  XNOR U4200 ( .A(n4098), .B(n4097), .Z(n4099) );
  XNOR U4201 ( .A(n4100), .B(n4099), .Z(n4104) );
  NANDN U4202 ( .A(n4051), .B(n4050), .Z(n4055) );
  NAND U4203 ( .A(n4053), .B(n4052), .Z(n4054) );
  AND U4204 ( .A(n4055), .B(n4054), .Z(n4103) );
  XOR U4205 ( .A(n4104), .B(n4103), .Z(n4105) );
  NANDN U4206 ( .A(n4057), .B(n4056), .Z(n4061) );
  NANDN U4207 ( .A(n4059), .B(n4058), .Z(n4060) );
  NAND U4208 ( .A(n4061), .B(n4060), .Z(n4106) );
  XOR U4209 ( .A(n4105), .B(n4106), .Z(n4073) );
  OR U4210 ( .A(n4063), .B(n4062), .Z(n4067) );
  NANDN U4211 ( .A(n4065), .B(n4064), .Z(n4066) );
  NAND U4212 ( .A(n4067), .B(n4066), .Z(n4074) );
  XNOR U4213 ( .A(n4073), .B(n4074), .Z(n4075) );
  XNOR U4214 ( .A(n4076), .B(n4075), .Z(n4109) );
  XNOR U4215 ( .A(n4109), .B(sreg[1113]), .Z(n4111) );
  NAND U4216 ( .A(n4068), .B(sreg[1112]), .Z(n4072) );
  OR U4217 ( .A(n4070), .B(n4069), .Z(n4071) );
  AND U4218 ( .A(n4072), .B(n4071), .Z(n4110) );
  XOR U4219 ( .A(n4111), .B(n4110), .Z(c[1113]) );
  NANDN U4220 ( .A(n4074), .B(n4073), .Z(n4078) );
  NAND U4221 ( .A(n4076), .B(n4075), .Z(n4077) );
  NAND U4222 ( .A(n4078), .B(n4077), .Z(n4117) );
  NAND U4223 ( .A(b[0]), .B(a[98]), .Z(n4079) );
  XNOR U4224 ( .A(b[1]), .B(n4079), .Z(n4081) );
  NAND U4225 ( .A(n29), .B(a[97]), .Z(n4080) );
  AND U4226 ( .A(n4081), .B(n4080), .Z(n4134) );
  XOR U4227 ( .A(a[94]), .B(n42197), .Z(n4123) );
  NANDN U4228 ( .A(n4123), .B(n42173), .Z(n4084) );
  NANDN U4229 ( .A(n4082), .B(n42172), .Z(n4083) );
  NAND U4230 ( .A(n4084), .B(n4083), .Z(n4132) );
  NAND U4231 ( .A(b[7]), .B(a[90]), .Z(n4133) );
  XNOR U4232 ( .A(n4132), .B(n4133), .Z(n4135) );
  XOR U4233 ( .A(n4134), .B(n4135), .Z(n4141) );
  NANDN U4234 ( .A(n4085), .B(n42093), .Z(n4087) );
  XOR U4235 ( .A(n42134), .B(a[96]), .Z(n4126) );
  NANDN U4236 ( .A(n4126), .B(n42095), .Z(n4086) );
  NAND U4237 ( .A(n4087), .B(n4086), .Z(n4139) );
  NANDN U4238 ( .A(n4088), .B(n42231), .Z(n4090) );
  XOR U4239 ( .A(n169), .B(a[92]), .Z(n4129) );
  NANDN U4240 ( .A(n4129), .B(n42234), .Z(n4089) );
  AND U4241 ( .A(n4090), .B(n4089), .Z(n4138) );
  XNOR U4242 ( .A(n4139), .B(n4138), .Z(n4140) );
  XNOR U4243 ( .A(n4141), .B(n4140), .Z(n4145) );
  NANDN U4244 ( .A(n4092), .B(n4091), .Z(n4096) );
  NAND U4245 ( .A(n4094), .B(n4093), .Z(n4095) );
  AND U4246 ( .A(n4096), .B(n4095), .Z(n4144) );
  XOR U4247 ( .A(n4145), .B(n4144), .Z(n4146) );
  NANDN U4248 ( .A(n4098), .B(n4097), .Z(n4102) );
  NANDN U4249 ( .A(n4100), .B(n4099), .Z(n4101) );
  NAND U4250 ( .A(n4102), .B(n4101), .Z(n4147) );
  XOR U4251 ( .A(n4146), .B(n4147), .Z(n4114) );
  OR U4252 ( .A(n4104), .B(n4103), .Z(n4108) );
  NANDN U4253 ( .A(n4106), .B(n4105), .Z(n4107) );
  NAND U4254 ( .A(n4108), .B(n4107), .Z(n4115) );
  XNOR U4255 ( .A(n4114), .B(n4115), .Z(n4116) );
  XNOR U4256 ( .A(n4117), .B(n4116), .Z(n4150) );
  XNOR U4257 ( .A(n4150), .B(sreg[1114]), .Z(n4152) );
  NAND U4258 ( .A(n4109), .B(sreg[1113]), .Z(n4113) );
  OR U4259 ( .A(n4111), .B(n4110), .Z(n4112) );
  AND U4260 ( .A(n4113), .B(n4112), .Z(n4151) );
  XOR U4261 ( .A(n4152), .B(n4151), .Z(c[1114]) );
  NANDN U4262 ( .A(n4115), .B(n4114), .Z(n4119) );
  NAND U4263 ( .A(n4117), .B(n4116), .Z(n4118) );
  NAND U4264 ( .A(n4119), .B(n4118), .Z(n4158) );
  NAND U4265 ( .A(b[0]), .B(a[99]), .Z(n4120) );
  XNOR U4266 ( .A(b[1]), .B(n4120), .Z(n4122) );
  NAND U4267 ( .A(n29), .B(a[98]), .Z(n4121) );
  AND U4268 ( .A(n4122), .B(n4121), .Z(n4175) );
  XOR U4269 ( .A(a[95]), .B(n42197), .Z(n4164) );
  NANDN U4270 ( .A(n4164), .B(n42173), .Z(n4125) );
  NANDN U4271 ( .A(n4123), .B(n42172), .Z(n4124) );
  NAND U4272 ( .A(n4125), .B(n4124), .Z(n4173) );
  NAND U4273 ( .A(b[7]), .B(a[91]), .Z(n4174) );
  XNOR U4274 ( .A(n4173), .B(n4174), .Z(n4176) );
  XOR U4275 ( .A(n4175), .B(n4176), .Z(n4182) );
  NANDN U4276 ( .A(n4126), .B(n42093), .Z(n4128) );
  XOR U4277 ( .A(n42134), .B(a[97]), .Z(n4167) );
  NANDN U4278 ( .A(n4167), .B(n42095), .Z(n4127) );
  NAND U4279 ( .A(n4128), .B(n4127), .Z(n4180) );
  NANDN U4280 ( .A(n4129), .B(n42231), .Z(n4131) );
  XOR U4281 ( .A(n169), .B(a[93]), .Z(n4170) );
  NANDN U4282 ( .A(n4170), .B(n42234), .Z(n4130) );
  AND U4283 ( .A(n4131), .B(n4130), .Z(n4179) );
  XNOR U4284 ( .A(n4180), .B(n4179), .Z(n4181) );
  XNOR U4285 ( .A(n4182), .B(n4181), .Z(n4186) );
  NANDN U4286 ( .A(n4133), .B(n4132), .Z(n4137) );
  NAND U4287 ( .A(n4135), .B(n4134), .Z(n4136) );
  AND U4288 ( .A(n4137), .B(n4136), .Z(n4185) );
  XOR U4289 ( .A(n4186), .B(n4185), .Z(n4187) );
  NANDN U4290 ( .A(n4139), .B(n4138), .Z(n4143) );
  NANDN U4291 ( .A(n4141), .B(n4140), .Z(n4142) );
  NAND U4292 ( .A(n4143), .B(n4142), .Z(n4188) );
  XOR U4293 ( .A(n4187), .B(n4188), .Z(n4155) );
  OR U4294 ( .A(n4145), .B(n4144), .Z(n4149) );
  NANDN U4295 ( .A(n4147), .B(n4146), .Z(n4148) );
  NAND U4296 ( .A(n4149), .B(n4148), .Z(n4156) );
  XNOR U4297 ( .A(n4155), .B(n4156), .Z(n4157) );
  XNOR U4298 ( .A(n4158), .B(n4157), .Z(n4191) );
  XNOR U4299 ( .A(n4191), .B(sreg[1115]), .Z(n4193) );
  NAND U4300 ( .A(n4150), .B(sreg[1114]), .Z(n4154) );
  OR U4301 ( .A(n4152), .B(n4151), .Z(n4153) );
  AND U4302 ( .A(n4154), .B(n4153), .Z(n4192) );
  XOR U4303 ( .A(n4193), .B(n4192), .Z(c[1115]) );
  NANDN U4304 ( .A(n4156), .B(n4155), .Z(n4160) );
  NAND U4305 ( .A(n4158), .B(n4157), .Z(n4159) );
  NAND U4306 ( .A(n4160), .B(n4159), .Z(n4199) );
  NAND U4307 ( .A(b[0]), .B(a[100]), .Z(n4161) );
  XNOR U4308 ( .A(b[1]), .B(n4161), .Z(n4163) );
  NAND U4309 ( .A(n29), .B(a[99]), .Z(n4162) );
  AND U4310 ( .A(n4163), .B(n4162), .Z(n4216) );
  XOR U4311 ( .A(a[96]), .B(n42197), .Z(n4205) );
  NANDN U4312 ( .A(n4205), .B(n42173), .Z(n4166) );
  NANDN U4313 ( .A(n4164), .B(n42172), .Z(n4165) );
  NAND U4314 ( .A(n4166), .B(n4165), .Z(n4214) );
  NAND U4315 ( .A(b[7]), .B(a[92]), .Z(n4215) );
  XNOR U4316 ( .A(n4214), .B(n4215), .Z(n4217) );
  XOR U4317 ( .A(n4216), .B(n4217), .Z(n4223) );
  NANDN U4318 ( .A(n4167), .B(n42093), .Z(n4169) );
  XOR U4319 ( .A(n42134), .B(a[98]), .Z(n4208) );
  NANDN U4320 ( .A(n4208), .B(n42095), .Z(n4168) );
  NAND U4321 ( .A(n4169), .B(n4168), .Z(n4221) );
  NANDN U4322 ( .A(n4170), .B(n42231), .Z(n4172) );
  XOR U4323 ( .A(n169), .B(a[94]), .Z(n4211) );
  NANDN U4324 ( .A(n4211), .B(n42234), .Z(n4171) );
  AND U4325 ( .A(n4172), .B(n4171), .Z(n4220) );
  XNOR U4326 ( .A(n4221), .B(n4220), .Z(n4222) );
  XNOR U4327 ( .A(n4223), .B(n4222), .Z(n4227) );
  NANDN U4328 ( .A(n4174), .B(n4173), .Z(n4178) );
  NAND U4329 ( .A(n4176), .B(n4175), .Z(n4177) );
  AND U4330 ( .A(n4178), .B(n4177), .Z(n4226) );
  XOR U4331 ( .A(n4227), .B(n4226), .Z(n4228) );
  NANDN U4332 ( .A(n4180), .B(n4179), .Z(n4184) );
  NANDN U4333 ( .A(n4182), .B(n4181), .Z(n4183) );
  NAND U4334 ( .A(n4184), .B(n4183), .Z(n4229) );
  XOR U4335 ( .A(n4228), .B(n4229), .Z(n4196) );
  OR U4336 ( .A(n4186), .B(n4185), .Z(n4190) );
  NANDN U4337 ( .A(n4188), .B(n4187), .Z(n4189) );
  NAND U4338 ( .A(n4190), .B(n4189), .Z(n4197) );
  XNOR U4339 ( .A(n4196), .B(n4197), .Z(n4198) );
  XNOR U4340 ( .A(n4199), .B(n4198), .Z(n4232) );
  XNOR U4341 ( .A(n4232), .B(sreg[1116]), .Z(n4234) );
  NAND U4342 ( .A(n4191), .B(sreg[1115]), .Z(n4195) );
  OR U4343 ( .A(n4193), .B(n4192), .Z(n4194) );
  AND U4344 ( .A(n4195), .B(n4194), .Z(n4233) );
  XOR U4345 ( .A(n4234), .B(n4233), .Z(c[1116]) );
  NANDN U4346 ( .A(n4197), .B(n4196), .Z(n4201) );
  NAND U4347 ( .A(n4199), .B(n4198), .Z(n4200) );
  NAND U4348 ( .A(n4201), .B(n4200), .Z(n4240) );
  NAND U4349 ( .A(b[0]), .B(a[101]), .Z(n4202) );
  XNOR U4350 ( .A(b[1]), .B(n4202), .Z(n4204) );
  NAND U4351 ( .A(n29), .B(a[100]), .Z(n4203) );
  AND U4352 ( .A(n4204), .B(n4203), .Z(n4257) );
  XOR U4353 ( .A(a[97]), .B(n42197), .Z(n4246) );
  NANDN U4354 ( .A(n4246), .B(n42173), .Z(n4207) );
  NANDN U4355 ( .A(n4205), .B(n42172), .Z(n4206) );
  NAND U4356 ( .A(n4207), .B(n4206), .Z(n4255) );
  NAND U4357 ( .A(b[7]), .B(a[93]), .Z(n4256) );
  XNOR U4358 ( .A(n4255), .B(n4256), .Z(n4258) );
  XOR U4359 ( .A(n4257), .B(n4258), .Z(n4264) );
  NANDN U4360 ( .A(n4208), .B(n42093), .Z(n4210) );
  XOR U4361 ( .A(n42134), .B(a[99]), .Z(n4249) );
  NANDN U4362 ( .A(n4249), .B(n42095), .Z(n4209) );
  NAND U4363 ( .A(n4210), .B(n4209), .Z(n4262) );
  NANDN U4364 ( .A(n4211), .B(n42231), .Z(n4213) );
  XOR U4365 ( .A(n170), .B(a[95]), .Z(n4252) );
  NANDN U4366 ( .A(n4252), .B(n42234), .Z(n4212) );
  AND U4367 ( .A(n4213), .B(n4212), .Z(n4261) );
  XNOR U4368 ( .A(n4262), .B(n4261), .Z(n4263) );
  XNOR U4369 ( .A(n4264), .B(n4263), .Z(n4268) );
  NANDN U4370 ( .A(n4215), .B(n4214), .Z(n4219) );
  NAND U4371 ( .A(n4217), .B(n4216), .Z(n4218) );
  AND U4372 ( .A(n4219), .B(n4218), .Z(n4267) );
  XOR U4373 ( .A(n4268), .B(n4267), .Z(n4269) );
  NANDN U4374 ( .A(n4221), .B(n4220), .Z(n4225) );
  NANDN U4375 ( .A(n4223), .B(n4222), .Z(n4224) );
  NAND U4376 ( .A(n4225), .B(n4224), .Z(n4270) );
  XOR U4377 ( .A(n4269), .B(n4270), .Z(n4237) );
  OR U4378 ( .A(n4227), .B(n4226), .Z(n4231) );
  NANDN U4379 ( .A(n4229), .B(n4228), .Z(n4230) );
  NAND U4380 ( .A(n4231), .B(n4230), .Z(n4238) );
  XNOR U4381 ( .A(n4237), .B(n4238), .Z(n4239) );
  XNOR U4382 ( .A(n4240), .B(n4239), .Z(n4273) );
  XNOR U4383 ( .A(n4273), .B(sreg[1117]), .Z(n4275) );
  NAND U4384 ( .A(n4232), .B(sreg[1116]), .Z(n4236) );
  OR U4385 ( .A(n4234), .B(n4233), .Z(n4235) );
  AND U4386 ( .A(n4236), .B(n4235), .Z(n4274) );
  XOR U4387 ( .A(n4275), .B(n4274), .Z(c[1117]) );
  NANDN U4388 ( .A(n4238), .B(n4237), .Z(n4242) );
  NAND U4389 ( .A(n4240), .B(n4239), .Z(n4241) );
  NAND U4390 ( .A(n4242), .B(n4241), .Z(n4281) );
  NAND U4391 ( .A(b[0]), .B(a[102]), .Z(n4243) );
  XNOR U4392 ( .A(b[1]), .B(n4243), .Z(n4245) );
  NAND U4393 ( .A(n29), .B(a[101]), .Z(n4244) );
  AND U4394 ( .A(n4245), .B(n4244), .Z(n4298) );
  XOR U4395 ( .A(a[98]), .B(n42197), .Z(n4287) );
  NANDN U4396 ( .A(n4287), .B(n42173), .Z(n4248) );
  NANDN U4397 ( .A(n4246), .B(n42172), .Z(n4247) );
  NAND U4398 ( .A(n4248), .B(n4247), .Z(n4296) );
  NAND U4399 ( .A(b[7]), .B(a[94]), .Z(n4297) );
  XNOR U4400 ( .A(n4296), .B(n4297), .Z(n4299) );
  XOR U4401 ( .A(n4298), .B(n4299), .Z(n4305) );
  NANDN U4402 ( .A(n4249), .B(n42093), .Z(n4251) );
  XOR U4403 ( .A(n42134), .B(a[100]), .Z(n4290) );
  NANDN U4404 ( .A(n4290), .B(n42095), .Z(n4250) );
  NAND U4405 ( .A(n4251), .B(n4250), .Z(n4303) );
  NANDN U4406 ( .A(n4252), .B(n42231), .Z(n4254) );
  XOR U4407 ( .A(n170), .B(a[96]), .Z(n4293) );
  NANDN U4408 ( .A(n4293), .B(n42234), .Z(n4253) );
  AND U4409 ( .A(n4254), .B(n4253), .Z(n4302) );
  XNOR U4410 ( .A(n4303), .B(n4302), .Z(n4304) );
  XNOR U4411 ( .A(n4305), .B(n4304), .Z(n4309) );
  NANDN U4412 ( .A(n4256), .B(n4255), .Z(n4260) );
  NAND U4413 ( .A(n4258), .B(n4257), .Z(n4259) );
  AND U4414 ( .A(n4260), .B(n4259), .Z(n4308) );
  XOR U4415 ( .A(n4309), .B(n4308), .Z(n4310) );
  NANDN U4416 ( .A(n4262), .B(n4261), .Z(n4266) );
  NANDN U4417 ( .A(n4264), .B(n4263), .Z(n4265) );
  NAND U4418 ( .A(n4266), .B(n4265), .Z(n4311) );
  XOR U4419 ( .A(n4310), .B(n4311), .Z(n4278) );
  OR U4420 ( .A(n4268), .B(n4267), .Z(n4272) );
  NANDN U4421 ( .A(n4270), .B(n4269), .Z(n4271) );
  NAND U4422 ( .A(n4272), .B(n4271), .Z(n4279) );
  XNOR U4423 ( .A(n4278), .B(n4279), .Z(n4280) );
  XNOR U4424 ( .A(n4281), .B(n4280), .Z(n4314) );
  XNOR U4425 ( .A(n4314), .B(sreg[1118]), .Z(n4316) );
  NAND U4426 ( .A(n4273), .B(sreg[1117]), .Z(n4277) );
  OR U4427 ( .A(n4275), .B(n4274), .Z(n4276) );
  AND U4428 ( .A(n4277), .B(n4276), .Z(n4315) );
  XOR U4429 ( .A(n4316), .B(n4315), .Z(c[1118]) );
  NANDN U4430 ( .A(n4279), .B(n4278), .Z(n4283) );
  NAND U4431 ( .A(n4281), .B(n4280), .Z(n4282) );
  NAND U4432 ( .A(n4283), .B(n4282), .Z(n4322) );
  NAND U4433 ( .A(b[0]), .B(a[103]), .Z(n4284) );
  XNOR U4434 ( .A(b[1]), .B(n4284), .Z(n4286) );
  NAND U4435 ( .A(n29), .B(a[102]), .Z(n4285) );
  AND U4436 ( .A(n4286), .B(n4285), .Z(n4339) );
  XOR U4437 ( .A(a[99]), .B(n42197), .Z(n4328) );
  NANDN U4438 ( .A(n4328), .B(n42173), .Z(n4289) );
  NANDN U4439 ( .A(n4287), .B(n42172), .Z(n4288) );
  NAND U4440 ( .A(n4289), .B(n4288), .Z(n4337) );
  NAND U4441 ( .A(b[7]), .B(a[95]), .Z(n4338) );
  XNOR U4442 ( .A(n4337), .B(n4338), .Z(n4340) );
  XOR U4443 ( .A(n4339), .B(n4340), .Z(n4346) );
  NANDN U4444 ( .A(n4290), .B(n42093), .Z(n4292) );
  XOR U4445 ( .A(n42134), .B(a[101]), .Z(n4331) );
  NANDN U4446 ( .A(n4331), .B(n42095), .Z(n4291) );
  NAND U4447 ( .A(n4292), .B(n4291), .Z(n4344) );
  NANDN U4448 ( .A(n4293), .B(n42231), .Z(n4295) );
  XOR U4449 ( .A(n170), .B(a[97]), .Z(n4334) );
  NANDN U4450 ( .A(n4334), .B(n42234), .Z(n4294) );
  AND U4451 ( .A(n4295), .B(n4294), .Z(n4343) );
  XNOR U4452 ( .A(n4344), .B(n4343), .Z(n4345) );
  XNOR U4453 ( .A(n4346), .B(n4345), .Z(n4350) );
  NANDN U4454 ( .A(n4297), .B(n4296), .Z(n4301) );
  NAND U4455 ( .A(n4299), .B(n4298), .Z(n4300) );
  AND U4456 ( .A(n4301), .B(n4300), .Z(n4349) );
  XOR U4457 ( .A(n4350), .B(n4349), .Z(n4351) );
  NANDN U4458 ( .A(n4303), .B(n4302), .Z(n4307) );
  NANDN U4459 ( .A(n4305), .B(n4304), .Z(n4306) );
  NAND U4460 ( .A(n4307), .B(n4306), .Z(n4352) );
  XOR U4461 ( .A(n4351), .B(n4352), .Z(n4319) );
  OR U4462 ( .A(n4309), .B(n4308), .Z(n4313) );
  NANDN U4463 ( .A(n4311), .B(n4310), .Z(n4312) );
  NAND U4464 ( .A(n4313), .B(n4312), .Z(n4320) );
  XNOR U4465 ( .A(n4319), .B(n4320), .Z(n4321) );
  XNOR U4466 ( .A(n4322), .B(n4321), .Z(n4355) );
  XNOR U4467 ( .A(n4355), .B(sreg[1119]), .Z(n4357) );
  NAND U4468 ( .A(n4314), .B(sreg[1118]), .Z(n4318) );
  OR U4469 ( .A(n4316), .B(n4315), .Z(n4317) );
  AND U4470 ( .A(n4318), .B(n4317), .Z(n4356) );
  XOR U4471 ( .A(n4357), .B(n4356), .Z(c[1119]) );
  NANDN U4472 ( .A(n4320), .B(n4319), .Z(n4324) );
  NAND U4473 ( .A(n4322), .B(n4321), .Z(n4323) );
  NAND U4474 ( .A(n4324), .B(n4323), .Z(n4363) );
  NAND U4475 ( .A(b[0]), .B(a[104]), .Z(n4325) );
  XNOR U4476 ( .A(b[1]), .B(n4325), .Z(n4327) );
  NAND U4477 ( .A(n29), .B(a[103]), .Z(n4326) );
  AND U4478 ( .A(n4327), .B(n4326), .Z(n4380) );
  XOR U4479 ( .A(a[100]), .B(n42197), .Z(n4369) );
  NANDN U4480 ( .A(n4369), .B(n42173), .Z(n4330) );
  NANDN U4481 ( .A(n4328), .B(n42172), .Z(n4329) );
  NAND U4482 ( .A(n4330), .B(n4329), .Z(n4378) );
  NAND U4483 ( .A(b[7]), .B(a[96]), .Z(n4379) );
  XNOR U4484 ( .A(n4378), .B(n4379), .Z(n4381) );
  XOR U4485 ( .A(n4380), .B(n4381), .Z(n4387) );
  NANDN U4486 ( .A(n4331), .B(n42093), .Z(n4333) );
  XOR U4487 ( .A(n42134), .B(a[102]), .Z(n4372) );
  NANDN U4488 ( .A(n4372), .B(n42095), .Z(n4332) );
  NAND U4489 ( .A(n4333), .B(n4332), .Z(n4385) );
  NANDN U4490 ( .A(n4334), .B(n42231), .Z(n4336) );
  XOR U4491 ( .A(n170), .B(a[98]), .Z(n4375) );
  NANDN U4492 ( .A(n4375), .B(n42234), .Z(n4335) );
  AND U4493 ( .A(n4336), .B(n4335), .Z(n4384) );
  XNOR U4494 ( .A(n4385), .B(n4384), .Z(n4386) );
  XNOR U4495 ( .A(n4387), .B(n4386), .Z(n4391) );
  NANDN U4496 ( .A(n4338), .B(n4337), .Z(n4342) );
  NAND U4497 ( .A(n4340), .B(n4339), .Z(n4341) );
  AND U4498 ( .A(n4342), .B(n4341), .Z(n4390) );
  XOR U4499 ( .A(n4391), .B(n4390), .Z(n4392) );
  NANDN U4500 ( .A(n4344), .B(n4343), .Z(n4348) );
  NANDN U4501 ( .A(n4346), .B(n4345), .Z(n4347) );
  NAND U4502 ( .A(n4348), .B(n4347), .Z(n4393) );
  XOR U4503 ( .A(n4392), .B(n4393), .Z(n4360) );
  OR U4504 ( .A(n4350), .B(n4349), .Z(n4354) );
  NANDN U4505 ( .A(n4352), .B(n4351), .Z(n4353) );
  NAND U4506 ( .A(n4354), .B(n4353), .Z(n4361) );
  XNOR U4507 ( .A(n4360), .B(n4361), .Z(n4362) );
  XNOR U4508 ( .A(n4363), .B(n4362), .Z(n4396) );
  XNOR U4509 ( .A(n4396), .B(sreg[1120]), .Z(n4398) );
  NAND U4510 ( .A(n4355), .B(sreg[1119]), .Z(n4359) );
  OR U4511 ( .A(n4357), .B(n4356), .Z(n4358) );
  AND U4512 ( .A(n4359), .B(n4358), .Z(n4397) );
  XOR U4513 ( .A(n4398), .B(n4397), .Z(c[1120]) );
  NANDN U4514 ( .A(n4361), .B(n4360), .Z(n4365) );
  NAND U4515 ( .A(n4363), .B(n4362), .Z(n4364) );
  NAND U4516 ( .A(n4365), .B(n4364), .Z(n4404) );
  NAND U4517 ( .A(b[0]), .B(a[105]), .Z(n4366) );
  XNOR U4518 ( .A(b[1]), .B(n4366), .Z(n4368) );
  NAND U4519 ( .A(n30), .B(a[104]), .Z(n4367) );
  AND U4520 ( .A(n4368), .B(n4367), .Z(n4421) );
  XOR U4521 ( .A(a[101]), .B(n42197), .Z(n4410) );
  NANDN U4522 ( .A(n4410), .B(n42173), .Z(n4371) );
  NANDN U4523 ( .A(n4369), .B(n42172), .Z(n4370) );
  NAND U4524 ( .A(n4371), .B(n4370), .Z(n4419) );
  NAND U4525 ( .A(b[7]), .B(a[97]), .Z(n4420) );
  XNOR U4526 ( .A(n4419), .B(n4420), .Z(n4422) );
  XOR U4527 ( .A(n4421), .B(n4422), .Z(n4428) );
  NANDN U4528 ( .A(n4372), .B(n42093), .Z(n4374) );
  XOR U4529 ( .A(n42134), .B(a[103]), .Z(n4413) );
  NANDN U4530 ( .A(n4413), .B(n42095), .Z(n4373) );
  NAND U4531 ( .A(n4374), .B(n4373), .Z(n4426) );
  NANDN U4532 ( .A(n4375), .B(n42231), .Z(n4377) );
  XOR U4533 ( .A(n170), .B(a[99]), .Z(n4416) );
  NANDN U4534 ( .A(n4416), .B(n42234), .Z(n4376) );
  AND U4535 ( .A(n4377), .B(n4376), .Z(n4425) );
  XNOR U4536 ( .A(n4426), .B(n4425), .Z(n4427) );
  XNOR U4537 ( .A(n4428), .B(n4427), .Z(n4432) );
  NANDN U4538 ( .A(n4379), .B(n4378), .Z(n4383) );
  NAND U4539 ( .A(n4381), .B(n4380), .Z(n4382) );
  AND U4540 ( .A(n4383), .B(n4382), .Z(n4431) );
  XOR U4541 ( .A(n4432), .B(n4431), .Z(n4433) );
  NANDN U4542 ( .A(n4385), .B(n4384), .Z(n4389) );
  NANDN U4543 ( .A(n4387), .B(n4386), .Z(n4388) );
  NAND U4544 ( .A(n4389), .B(n4388), .Z(n4434) );
  XOR U4545 ( .A(n4433), .B(n4434), .Z(n4401) );
  OR U4546 ( .A(n4391), .B(n4390), .Z(n4395) );
  NANDN U4547 ( .A(n4393), .B(n4392), .Z(n4394) );
  NAND U4548 ( .A(n4395), .B(n4394), .Z(n4402) );
  XNOR U4549 ( .A(n4401), .B(n4402), .Z(n4403) );
  XNOR U4550 ( .A(n4404), .B(n4403), .Z(n4437) );
  XNOR U4551 ( .A(n4437), .B(sreg[1121]), .Z(n4439) );
  NAND U4552 ( .A(n4396), .B(sreg[1120]), .Z(n4400) );
  OR U4553 ( .A(n4398), .B(n4397), .Z(n4399) );
  AND U4554 ( .A(n4400), .B(n4399), .Z(n4438) );
  XOR U4555 ( .A(n4439), .B(n4438), .Z(c[1121]) );
  NANDN U4556 ( .A(n4402), .B(n4401), .Z(n4406) );
  NAND U4557 ( .A(n4404), .B(n4403), .Z(n4405) );
  NAND U4558 ( .A(n4406), .B(n4405), .Z(n4445) );
  NAND U4559 ( .A(b[0]), .B(a[106]), .Z(n4407) );
  XNOR U4560 ( .A(b[1]), .B(n4407), .Z(n4409) );
  NAND U4561 ( .A(n30), .B(a[105]), .Z(n4408) );
  AND U4562 ( .A(n4409), .B(n4408), .Z(n4462) );
  XOR U4563 ( .A(a[102]), .B(n42197), .Z(n4451) );
  NANDN U4564 ( .A(n4451), .B(n42173), .Z(n4412) );
  NANDN U4565 ( .A(n4410), .B(n42172), .Z(n4411) );
  NAND U4566 ( .A(n4412), .B(n4411), .Z(n4460) );
  NAND U4567 ( .A(b[7]), .B(a[98]), .Z(n4461) );
  XNOR U4568 ( .A(n4460), .B(n4461), .Z(n4463) );
  XOR U4569 ( .A(n4462), .B(n4463), .Z(n4469) );
  NANDN U4570 ( .A(n4413), .B(n42093), .Z(n4415) );
  XOR U4571 ( .A(n42134), .B(a[104]), .Z(n4454) );
  NANDN U4572 ( .A(n4454), .B(n42095), .Z(n4414) );
  NAND U4573 ( .A(n4415), .B(n4414), .Z(n4467) );
  NANDN U4574 ( .A(n4416), .B(n42231), .Z(n4418) );
  XOR U4575 ( .A(n170), .B(a[100]), .Z(n4457) );
  NANDN U4576 ( .A(n4457), .B(n42234), .Z(n4417) );
  AND U4577 ( .A(n4418), .B(n4417), .Z(n4466) );
  XNOR U4578 ( .A(n4467), .B(n4466), .Z(n4468) );
  XNOR U4579 ( .A(n4469), .B(n4468), .Z(n4473) );
  NANDN U4580 ( .A(n4420), .B(n4419), .Z(n4424) );
  NAND U4581 ( .A(n4422), .B(n4421), .Z(n4423) );
  AND U4582 ( .A(n4424), .B(n4423), .Z(n4472) );
  XOR U4583 ( .A(n4473), .B(n4472), .Z(n4474) );
  NANDN U4584 ( .A(n4426), .B(n4425), .Z(n4430) );
  NANDN U4585 ( .A(n4428), .B(n4427), .Z(n4429) );
  NAND U4586 ( .A(n4430), .B(n4429), .Z(n4475) );
  XOR U4587 ( .A(n4474), .B(n4475), .Z(n4442) );
  OR U4588 ( .A(n4432), .B(n4431), .Z(n4436) );
  NANDN U4589 ( .A(n4434), .B(n4433), .Z(n4435) );
  NAND U4590 ( .A(n4436), .B(n4435), .Z(n4443) );
  XNOR U4591 ( .A(n4442), .B(n4443), .Z(n4444) );
  XNOR U4592 ( .A(n4445), .B(n4444), .Z(n4478) );
  XNOR U4593 ( .A(n4478), .B(sreg[1122]), .Z(n4480) );
  NAND U4594 ( .A(n4437), .B(sreg[1121]), .Z(n4441) );
  OR U4595 ( .A(n4439), .B(n4438), .Z(n4440) );
  AND U4596 ( .A(n4441), .B(n4440), .Z(n4479) );
  XOR U4597 ( .A(n4480), .B(n4479), .Z(c[1122]) );
  NANDN U4598 ( .A(n4443), .B(n4442), .Z(n4447) );
  NAND U4599 ( .A(n4445), .B(n4444), .Z(n4446) );
  NAND U4600 ( .A(n4447), .B(n4446), .Z(n4486) );
  NAND U4601 ( .A(b[0]), .B(a[107]), .Z(n4448) );
  XNOR U4602 ( .A(b[1]), .B(n4448), .Z(n4450) );
  NAND U4603 ( .A(n30), .B(a[106]), .Z(n4449) );
  AND U4604 ( .A(n4450), .B(n4449), .Z(n4503) );
  XOR U4605 ( .A(a[103]), .B(n42197), .Z(n4492) );
  NANDN U4606 ( .A(n4492), .B(n42173), .Z(n4453) );
  NANDN U4607 ( .A(n4451), .B(n42172), .Z(n4452) );
  NAND U4608 ( .A(n4453), .B(n4452), .Z(n4501) );
  NAND U4609 ( .A(b[7]), .B(a[99]), .Z(n4502) );
  XNOR U4610 ( .A(n4501), .B(n4502), .Z(n4504) );
  XOR U4611 ( .A(n4503), .B(n4504), .Z(n4510) );
  NANDN U4612 ( .A(n4454), .B(n42093), .Z(n4456) );
  XOR U4613 ( .A(n42134), .B(a[105]), .Z(n4495) );
  NANDN U4614 ( .A(n4495), .B(n42095), .Z(n4455) );
  NAND U4615 ( .A(n4456), .B(n4455), .Z(n4508) );
  NANDN U4616 ( .A(n4457), .B(n42231), .Z(n4459) );
  XOR U4617 ( .A(n170), .B(a[101]), .Z(n4498) );
  NANDN U4618 ( .A(n4498), .B(n42234), .Z(n4458) );
  AND U4619 ( .A(n4459), .B(n4458), .Z(n4507) );
  XNOR U4620 ( .A(n4508), .B(n4507), .Z(n4509) );
  XNOR U4621 ( .A(n4510), .B(n4509), .Z(n4514) );
  NANDN U4622 ( .A(n4461), .B(n4460), .Z(n4465) );
  NAND U4623 ( .A(n4463), .B(n4462), .Z(n4464) );
  AND U4624 ( .A(n4465), .B(n4464), .Z(n4513) );
  XOR U4625 ( .A(n4514), .B(n4513), .Z(n4515) );
  NANDN U4626 ( .A(n4467), .B(n4466), .Z(n4471) );
  NANDN U4627 ( .A(n4469), .B(n4468), .Z(n4470) );
  NAND U4628 ( .A(n4471), .B(n4470), .Z(n4516) );
  XOR U4629 ( .A(n4515), .B(n4516), .Z(n4483) );
  OR U4630 ( .A(n4473), .B(n4472), .Z(n4477) );
  NANDN U4631 ( .A(n4475), .B(n4474), .Z(n4476) );
  NAND U4632 ( .A(n4477), .B(n4476), .Z(n4484) );
  XNOR U4633 ( .A(n4483), .B(n4484), .Z(n4485) );
  XNOR U4634 ( .A(n4486), .B(n4485), .Z(n4519) );
  XNOR U4635 ( .A(n4519), .B(sreg[1123]), .Z(n4521) );
  NAND U4636 ( .A(n4478), .B(sreg[1122]), .Z(n4482) );
  OR U4637 ( .A(n4480), .B(n4479), .Z(n4481) );
  AND U4638 ( .A(n4482), .B(n4481), .Z(n4520) );
  XOR U4639 ( .A(n4521), .B(n4520), .Z(c[1123]) );
  NANDN U4640 ( .A(n4484), .B(n4483), .Z(n4488) );
  NAND U4641 ( .A(n4486), .B(n4485), .Z(n4487) );
  NAND U4642 ( .A(n4488), .B(n4487), .Z(n4527) );
  NAND U4643 ( .A(b[0]), .B(a[108]), .Z(n4489) );
  XNOR U4644 ( .A(b[1]), .B(n4489), .Z(n4491) );
  NAND U4645 ( .A(n30), .B(a[107]), .Z(n4490) );
  AND U4646 ( .A(n4491), .B(n4490), .Z(n4544) );
  XOR U4647 ( .A(a[104]), .B(n42197), .Z(n4533) );
  NANDN U4648 ( .A(n4533), .B(n42173), .Z(n4494) );
  NANDN U4649 ( .A(n4492), .B(n42172), .Z(n4493) );
  NAND U4650 ( .A(n4494), .B(n4493), .Z(n4542) );
  NAND U4651 ( .A(b[7]), .B(a[100]), .Z(n4543) );
  XNOR U4652 ( .A(n4542), .B(n4543), .Z(n4545) );
  XOR U4653 ( .A(n4544), .B(n4545), .Z(n4551) );
  NANDN U4654 ( .A(n4495), .B(n42093), .Z(n4497) );
  XOR U4655 ( .A(n42134), .B(a[106]), .Z(n4536) );
  NANDN U4656 ( .A(n4536), .B(n42095), .Z(n4496) );
  NAND U4657 ( .A(n4497), .B(n4496), .Z(n4549) );
  NANDN U4658 ( .A(n4498), .B(n42231), .Z(n4500) );
  XOR U4659 ( .A(n170), .B(a[102]), .Z(n4539) );
  NANDN U4660 ( .A(n4539), .B(n42234), .Z(n4499) );
  AND U4661 ( .A(n4500), .B(n4499), .Z(n4548) );
  XNOR U4662 ( .A(n4549), .B(n4548), .Z(n4550) );
  XNOR U4663 ( .A(n4551), .B(n4550), .Z(n4555) );
  NANDN U4664 ( .A(n4502), .B(n4501), .Z(n4506) );
  NAND U4665 ( .A(n4504), .B(n4503), .Z(n4505) );
  AND U4666 ( .A(n4506), .B(n4505), .Z(n4554) );
  XOR U4667 ( .A(n4555), .B(n4554), .Z(n4556) );
  NANDN U4668 ( .A(n4508), .B(n4507), .Z(n4512) );
  NANDN U4669 ( .A(n4510), .B(n4509), .Z(n4511) );
  NAND U4670 ( .A(n4512), .B(n4511), .Z(n4557) );
  XOR U4671 ( .A(n4556), .B(n4557), .Z(n4524) );
  OR U4672 ( .A(n4514), .B(n4513), .Z(n4518) );
  NANDN U4673 ( .A(n4516), .B(n4515), .Z(n4517) );
  NAND U4674 ( .A(n4518), .B(n4517), .Z(n4525) );
  XNOR U4675 ( .A(n4524), .B(n4525), .Z(n4526) );
  XNOR U4676 ( .A(n4527), .B(n4526), .Z(n4560) );
  XNOR U4677 ( .A(n4560), .B(sreg[1124]), .Z(n4562) );
  NAND U4678 ( .A(n4519), .B(sreg[1123]), .Z(n4523) );
  OR U4679 ( .A(n4521), .B(n4520), .Z(n4522) );
  AND U4680 ( .A(n4523), .B(n4522), .Z(n4561) );
  XOR U4681 ( .A(n4562), .B(n4561), .Z(c[1124]) );
  NANDN U4682 ( .A(n4525), .B(n4524), .Z(n4529) );
  NAND U4683 ( .A(n4527), .B(n4526), .Z(n4528) );
  NAND U4684 ( .A(n4529), .B(n4528), .Z(n4568) );
  NAND U4685 ( .A(b[0]), .B(a[109]), .Z(n4530) );
  XNOR U4686 ( .A(b[1]), .B(n4530), .Z(n4532) );
  NAND U4687 ( .A(n30), .B(a[108]), .Z(n4531) );
  AND U4688 ( .A(n4532), .B(n4531), .Z(n4585) );
  XOR U4689 ( .A(a[105]), .B(n42197), .Z(n4574) );
  NANDN U4690 ( .A(n4574), .B(n42173), .Z(n4535) );
  NANDN U4691 ( .A(n4533), .B(n42172), .Z(n4534) );
  NAND U4692 ( .A(n4535), .B(n4534), .Z(n4583) );
  NAND U4693 ( .A(b[7]), .B(a[101]), .Z(n4584) );
  XNOR U4694 ( .A(n4583), .B(n4584), .Z(n4586) );
  XOR U4695 ( .A(n4585), .B(n4586), .Z(n4592) );
  NANDN U4696 ( .A(n4536), .B(n42093), .Z(n4538) );
  XOR U4697 ( .A(n42134), .B(a[107]), .Z(n4577) );
  NANDN U4698 ( .A(n4577), .B(n42095), .Z(n4537) );
  NAND U4699 ( .A(n4538), .B(n4537), .Z(n4590) );
  NANDN U4700 ( .A(n4539), .B(n42231), .Z(n4541) );
  XOR U4701 ( .A(n170), .B(a[103]), .Z(n4580) );
  NANDN U4702 ( .A(n4580), .B(n42234), .Z(n4540) );
  AND U4703 ( .A(n4541), .B(n4540), .Z(n4589) );
  XNOR U4704 ( .A(n4590), .B(n4589), .Z(n4591) );
  XNOR U4705 ( .A(n4592), .B(n4591), .Z(n4596) );
  NANDN U4706 ( .A(n4543), .B(n4542), .Z(n4547) );
  NAND U4707 ( .A(n4545), .B(n4544), .Z(n4546) );
  AND U4708 ( .A(n4547), .B(n4546), .Z(n4595) );
  XOR U4709 ( .A(n4596), .B(n4595), .Z(n4597) );
  NANDN U4710 ( .A(n4549), .B(n4548), .Z(n4553) );
  NANDN U4711 ( .A(n4551), .B(n4550), .Z(n4552) );
  NAND U4712 ( .A(n4553), .B(n4552), .Z(n4598) );
  XOR U4713 ( .A(n4597), .B(n4598), .Z(n4565) );
  OR U4714 ( .A(n4555), .B(n4554), .Z(n4559) );
  NANDN U4715 ( .A(n4557), .B(n4556), .Z(n4558) );
  NAND U4716 ( .A(n4559), .B(n4558), .Z(n4566) );
  XNOR U4717 ( .A(n4565), .B(n4566), .Z(n4567) );
  XNOR U4718 ( .A(n4568), .B(n4567), .Z(n4601) );
  XNOR U4719 ( .A(n4601), .B(sreg[1125]), .Z(n4603) );
  NAND U4720 ( .A(n4560), .B(sreg[1124]), .Z(n4564) );
  OR U4721 ( .A(n4562), .B(n4561), .Z(n4563) );
  AND U4722 ( .A(n4564), .B(n4563), .Z(n4602) );
  XOR U4723 ( .A(n4603), .B(n4602), .Z(c[1125]) );
  NANDN U4724 ( .A(n4566), .B(n4565), .Z(n4570) );
  NAND U4725 ( .A(n4568), .B(n4567), .Z(n4569) );
  NAND U4726 ( .A(n4570), .B(n4569), .Z(n4609) );
  NAND U4727 ( .A(b[0]), .B(a[110]), .Z(n4571) );
  XNOR U4728 ( .A(b[1]), .B(n4571), .Z(n4573) );
  NAND U4729 ( .A(n30), .B(a[109]), .Z(n4572) );
  AND U4730 ( .A(n4573), .B(n4572), .Z(n4626) );
  XOR U4731 ( .A(a[106]), .B(n42197), .Z(n4615) );
  NANDN U4732 ( .A(n4615), .B(n42173), .Z(n4576) );
  NANDN U4733 ( .A(n4574), .B(n42172), .Z(n4575) );
  NAND U4734 ( .A(n4576), .B(n4575), .Z(n4624) );
  NAND U4735 ( .A(b[7]), .B(a[102]), .Z(n4625) );
  XNOR U4736 ( .A(n4624), .B(n4625), .Z(n4627) );
  XOR U4737 ( .A(n4626), .B(n4627), .Z(n4633) );
  NANDN U4738 ( .A(n4577), .B(n42093), .Z(n4579) );
  XOR U4739 ( .A(n42134), .B(a[108]), .Z(n4618) );
  NANDN U4740 ( .A(n4618), .B(n42095), .Z(n4578) );
  NAND U4741 ( .A(n4579), .B(n4578), .Z(n4631) );
  NANDN U4742 ( .A(n4580), .B(n42231), .Z(n4582) );
  XOR U4743 ( .A(n170), .B(a[104]), .Z(n4621) );
  NANDN U4744 ( .A(n4621), .B(n42234), .Z(n4581) );
  AND U4745 ( .A(n4582), .B(n4581), .Z(n4630) );
  XNOR U4746 ( .A(n4631), .B(n4630), .Z(n4632) );
  XNOR U4747 ( .A(n4633), .B(n4632), .Z(n4637) );
  NANDN U4748 ( .A(n4584), .B(n4583), .Z(n4588) );
  NAND U4749 ( .A(n4586), .B(n4585), .Z(n4587) );
  AND U4750 ( .A(n4588), .B(n4587), .Z(n4636) );
  XOR U4751 ( .A(n4637), .B(n4636), .Z(n4638) );
  NANDN U4752 ( .A(n4590), .B(n4589), .Z(n4594) );
  NANDN U4753 ( .A(n4592), .B(n4591), .Z(n4593) );
  NAND U4754 ( .A(n4594), .B(n4593), .Z(n4639) );
  XOR U4755 ( .A(n4638), .B(n4639), .Z(n4606) );
  OR U4756 ( .A(n4596), .B(n4595), .Z(n4600) );
  NANDN U4757 ( .A(n4598), .B(n4597), .Z(n4599) );
  NAND U4758 ( .A(n4600), .B(n4599), .Z(n4607) );
  XNOR U4759 ( .A(n4606), .B(n4607), .Z(n4608) );
  XNOR U4760 ( .A(n4609), .B(n4608), .Z(n4642) );
  XNOR U4761 ( .A(n4642), .B(sreg[1126]), .Z(n4644) );
  NAND U4762 ( .A(n4601), .B(sreg[1125]), .Z(n4605) );
  OR U4763 ( .A(n4603), .B(n4602), .Z(n4604) );
  AND U4764 ( .A(n4605), .B(n4604), .Z(n4643) );
  XOR U4765 ( .A(n4644), .B(n4643), .Z(c[1126]) );
  NANDN U4766 ( .A(n4607), .B(n4606), .Z(n4611) );
  NAND U4767 ( .A(n4609), .B(n4608), .Z(n4610) );
  NAND U4768 ( .A(n4611), .B(n4610), .Z(n4650) );
  NAND U4769 ( .A(b[0]), .B(a[111]), .Z(n4612) );
  XNOR U4770 ( .A(b[1]), .B(n4612), .Z(n4614) );
  NAND U4771 ( .A(n30), .B(a[110]), .Z(n4613) );
  AND U4772 ( .A(n4614), .B(n4613), .Z(n4667) );
  XOR U4773 ( .A(a[107]), .B(n42197), .Z(n4656) );
  NANDN U4774 ( .A(n4656), .B(n42173), .Z(n4617) );
  NANDN U4775 ( .A(n4615), .B(n42172), .Z(n4616) );
  NAND U4776 ( .A(n4617), .B(n4616), .Z(n4665) );
  NAND U4777 ( .A(b[7]), .B(a[103]), .Z(n4666) );
  XNOR U4778 ( .A(n4665), .B(n4666), .Z(n4668) );
  XOR U4779 ( .A(n4667), .B(n4668), .Z(n4674) );
  NANDN U4780 ( .A(n4618), .B(n42093), .Z(n4620) );
  XOR U4781 ( .A(n42134), .B(a[109]), .Z(n4659) );
  NANDN U4782 ( .A(n4659), .B(n42095), .Z(n4619) );
  NAND U4783 ( .A(n4620), .B(n4619), .Z(n4672) );
  NANDN U4784 ( .A(n4621), .B(n42231), .Z(n4623) );
  XOR U4785 ( .A(n170), .B(a[105]), .Z(n4662) );
  NANDN U4786 ( .A(n4662), .B(n42234), .Z(n4622) );
  AND U4787 ( .A(n4623), .B(n4622), .Z(n4671) );
  XNOR U4788 ( .A(n4672), .B(n4671), .Z(n4673) );
  XNOR U4789 ( .A(n4674), .B(n4673), .Z(n4678) );
  NANDN U4790 ( .A(n4625), .B(n4624), .Z(n4629) );
  NAND U4791 ( .A(n4627), .B(n4626), .Z(n4628) );
  AND U4792 ( .A(n4629), .B(n4628), .Z(n4677) );
  XOR U4793 ( .A(n4678), .B(n4677), .Z(n4679) );
  NANDN U4794 ( .A(n4631), .B(n4630), .Z(n4635) );
  NANDN U4795 ( .A(n4633), .B(n4632), .Z(n4634) );
  NAND U4796 ( .A(n4635), .B(n4634), .Z(n4680) );
  XOR U4797 ( .A(n4679), .B(n4680), .Z(n4647) );
  OR U4798 ( .A(n4637), .B(n4636), .Z(n4641) );
  NANDN U4799 ( .A(n4639), .B(n4638), .Z(n4640) );
  NAND U4800 ( .A(n4641), .B(n4640), .Z(n4648) );
  XNOR U4801 ( .A(n4647), .B(n4648), .Z(n4649) );
  XNOR U4802 ( .A(n4650), .B(n4649), .Z(n4683) );
  XNOR U4803 ( .A(n4683), .B(sreg[1127]), .Z(n4685) );
  NAND U4804 ( .A(n4642), .B(sreg[1126]), .Z(n4646) );
  OR U4805 ( .A(n4644), .B(n4643), .Z(n4645) );
  AND U4806 ( .A(n4646), .B(n4645), .Z(n4684) );
  XOR U4807 ( .A(n4685), .B(n4684), .Z(c[1127]) );
  NANDN U4808 ( .A(n4648), .B(n4647), .Z(n4652) );
  NAND U4809 ( .A(n4650), .B(n4649), .Z(n4651) );
  NAND U4810 ( .A(n4652), .B(n4651), .Z(n4691) );
  NAND U4811 ( .A(b[0]), .B(a[112]), .Z(n4653) );
  XNOR U4812 ( .A(b[1]), .B(n4653), .Z(n4655) );
  NAND U4813 ( .A(n31), .B(a[111]), .Z(n4654) );
  AND U4814 ( .A(n4655), .B(n4654), .Z(n4708) );
  XOR U4815 ( .A(a[108]), .B(n42197), .Z(n4697) );
  NANDN U4816 ( .A(n4697), .B(n42173), .Z(n4658) );
  NANDN U4817 ( .A(n4656), .B(n42172), .Z(n4657) );
  NAND U4818 ( .A(n4658), .B(n4657), .Z(n4706) );
  NAND U4819 ( .A(b[7]), .B(a[104]), .Z(n4707) );
  XNOR U4820 ( .A(n4706), .B(n4707), .Z(n4709) );
  XOR U4821 ( .A(n4708), .B(n4709), .Z(n4715) );
  NANDN U4822 ( .A(n4659), .B(n42093), .Z(n4661) );
  XOR U4823 ( .A(n42134), .B(a[110]), .Z(n4700) );
  NANDN U4824 ( .A(n4700), .B(n42095), .Z(n4660) );
  NAND U4825 ( .A(n4661), .B(n4660), .Z(n4713) );
  NANDN U4826 ( .A(n4662), .B(n42231), .Z(n4664) );
  XOR U4827 ( .A(n170), .B(a[106]), .Z(n4703) );
  NANDN U4828 ( .A(n4703), .B(n42234), .Z(n4663) );
  AND U4829 ( .A(n4664), .B(n4663), .Z(n4712) );
  XNOR U4830 ( .A(n4713), .B(n4712), .Z(n4714) );
  XNOR U4831 ( .A(n4715), .B(n4714), .Z(n4719) );
  NANDN U4832 ( .A(n4666), .B(n4665), .Z(n4670) );
  NAND U4833 ( .A(n4668), .B(n4667), .Z(n4669) );
  AND U4834 ( .A(n4670), .B(n4669), .Z(n4718) );
  XOR U4835 ( .A(n4719), .B(n4718), .Z(n4720) );
  NANDN U4836 ( .A(n4672), .B(n4671), .Z(n4676) );
  NANDN U4837 ( .A(n4674), .B(n4673), .Z(n4675) );
  NAND U4838 ( .A(n4676), .B(n4675), .Z(n4721) );
  XOR U4839 ( .A(n4720), .B(n4721), .Z(n4688) );
  OR U4840 ( .A(n4678), .B(n4677), .Z(n4682) );
  NANDN U4841 ( .A(n4680), .B(n4679), .Z(n4681) );
  NAND U4842 ( .A(n4682), .B(n4681), .Z(n4689) );
  XNOR U4843 ( .A(n4688), .B(n4689), .Z(n4690) );
  XNOR U4844 ( .A(n4691), .B(n4690), .Z(n4724) );
  XNOR U4845 ( .A(n4724), .B(sreg[1128]), .Z(n4726) );
  NAND U4846 ( .A(n4683), .B(sreg[1127]), .Z(n4687) );
  OR U4847 ( .A(n4685), .B(n4684), .Z(n4686) );
  AND U4848 ( .A(n4687), .B(n4686), .Z(n4725) );
  XOR U4849 ( .A(n4726), .B(n4725), .Z(c[1128]) );
  NANDN U4850 ( .A(n4689), .B(n4688), .Z(n4693) );
  NAND U4851 ( .A(n4691), .B(n4690), .Z(n4692) );
  NAND U4852 ( .A(n4693), .B(n4692), .Z(n4732) );
  NAND U4853 ( .A(b[0]), .B(a[113]), .Z(n4694) );
  XNOR U4854 ( .A(b[1]), .B(n4694), .Z(n4696) );
  NAND U4855 ( .A(n31), .B(a[112]), .Z(n4695) );
  AND U4856 ( .A(n4696), .B(n4695), .Z(n4749) );
  XOR U4857 ( .A(a[109]), .B(n42197), .Z(n4738) );
  NANDN U4858 ( .A(n4738), .B(n42173), .Z(n4699) );
  NANDN U4859 ( .A(n4697), .B(n42172), .Z(n4698) );
  NAND U4860 ( .A(n4699), .B(n4698), .Z(n4747) );
  NAND U4861 ( .A(b[7]), .B(a[105]), .Z(n4748) );
  XNOR U4862 ( .A(n4747), .B(n4748), .Z(n4750) );
  XOR U4863 ( .A(n4749), .B(n4750), .Z(n4756) );
  NANDN U4864 ( .A(n4700), .B(n42093), .Z(n4702) );
  XOR U4865 ( .A(n42134), .B(a[111]), .Z(n4741) );
  NANDN U4866 ( .A(n4741), .B(n42095), .Z(n4701) );
  NAND U4867 ( .A(n4702), .B(n4701), .Z(n4754) );
  NANDN U4868 ( .A(n4703), .B(n42231), .Z(n4705) );
  XOR U4869 ( .A(n171), .B(a[107]), .Z(n4744) );
  NANDN U4870 ( .A(n4744), .B(n42234), .Z(n4704) );
  AND U4871 ( .A(n4705), .B(n4704), .Z(n4753) );
  XNOR U4872 ( .A(n4754), .B(n4753), .Z(n4755) );
  XNOR U4873 ( .A(n4756), .B(n4755), .Z(n4760) );
  NANDN U4874 ( .A(n4707), .B(n4706), .Z(n4711) );
  NAND U4875 ( .A(n4709), .B(n4708), .Z(n4710) );
  AND U4876 ( .A(n4711), .B(n4710), .Z(n4759) );
  XOR U4877 ( .A(n4760), .B(n4759), .Z(n4761) );
  NANDN U4878 ( .A(n4713), .B(n4712), .Z(n4717) );
  NANDN U4879 ( .A(n4715), .B(n4714), .Z(n4716) );
  NAND U4880 ( .A(n4717), .B(n4716), .Z(n4762) );
  XOR U4881 ( .A(n4761), .B(n4762), .Z(n4729) );
  OR U4882 ( .A(n4719), .B(n4718), .Z(n4723) );
  NANDN U4883 ( .A(n4721), .B(n4720), .Z(n4722) );
  NAND U4884 ( .A(n4723), .B(n4722), .Z(n4730) );
  XNOR U4885 ( .A(n4729), .B(n4730), .Z(n4731) );
  XNOR U4886 ( .A(n4732), .B(n4731), .Z(n4765) );
  XNOR U4887 ( .A(n4765), .B(sreg[1129]), .Z(n4767) );
  NAND U4888 ( .A(n4724), .B(sreg[1128]), .Z(n4728) );
  OR U4889 ( .A(n4726), .B(n4725), .Z(n4727) );
  AND U4890 ( .A(n4728), .B(n4727), .Z(n4766) );
  XOR U4891 ( .A(n4767), .B(n4766), .Z(c[1129]) );
  NANDN U4892 ( .A(n4730), .B(n4729), .Z(n4734) );
  NAND U4893 ( .A(n4732), .B(n4731), .Z(n4733) );
  NAND U4894 ( .A(n4734), .B(n4733), .Z(n4773) );
  NAND U4895 ( .A(b[0]), .B(a[114]), .Z(n4735) );
  XNOR U4896 ( .A(b[1]), .B(n4735), .Z(n4737) );
  NAND U4897 ( .A(n31), .B(a[113]), .Z(n4736) );
  AND U4898 ( .A(n4737), .B(n4736), .Z(n4790) );
  XOR U4899 ( .A(a[110]), .B(n42197), .Z(n4779) );
  NANDN U4900 ( .A(n4779), .B(n42173), .Z(n4740) );
  NANDN U4901 ( .A(n4738), .B(n42172), .Z(n4739) );
  NAND U4902 ( .A(n4740), .B(n4739), .Z(n4788) );
  NAND U4903 ( .A(b[7]), .B(a[106]), .Z(n4789) );
  XNOR U4904 ( .A(n4788), .B(n4789), .Z(n4791) );
  XOR U4905 ( .A(n4790), .B(n4791), .Z(n4797) );
  NANDN U4906 ( .A(n4741), .B(n42093), .Z(n4743) );
  XOR U4907 ( .A(n42134), .B(a[112]), .Z(n4782) );
  NANDN U4908 ( .A(n4782), .B(n42095), .Z(n4742) );
  NAND U4909 ( .A(n4743), .B(n4742), .Z(n4795) );
  NANDN U4910 ( .A(n4744), .B(n42231), .Z(n4746) );
  XOR U4911 ( .A(n171), .B(a[108]), .Z(n4785) );
  NANDN U4912 ( .A(n4785), .B(n42234), .Z(n4745) );
  AND U4913 ( .A(n4746), .B(n4745), .Z(n4794) );
  XNOR U4914 ( .A(n4795), .B(n4794), .Z(n4796) );
  XNOR U4915 ( .A(n4797), .B(n4796), .Z(n4801) );
  NANDN U4916 ( .A(n4748), .B(n4747), .Z(n4752) );
  NAND U4917 ( .A(n4750), .B(n4749), .Z(n4751) );
  AND U4918 ( .A(n4752), .B(n4751), .Z(n4800) );
  XOR U4919 ( .A(n4801), .B(n4800), .Z(n4802) );
  NANDN U4920 ( .A(n4754), .B(n4753), .Z(n4758) );
  NANDN U4921 ( .A(n4756), .B(n4755), .Z(n4757) );
  NAND U4922 ( .A(n4758), .B(n4757), .Z(n4803) );
  XOR U4923 ( .A(n4802), .B(n4803), .Z(n4770) );
  OR U4924 ( .A(n4760), .B(n4759), .Z(n4764) );
  NANDN U4925 ( .A(n4762), .B(n4761), .Z(n4763) );
  NAND U4926 ( .A(n4764), .B(n4763), .Z(n4771) );
  XNOR U4927 ( .A(n4770), .B(n4771), .Z(n4772) );
  XNOR U4928 ( .A(n4773), .B(n4772), .Z(n4806) );
  XNOR U4929 ( .A(n4806), .B(sreg[1130]), .Z(n4808) );
  NAND U4930 ( .A(n4765), .B(sreg[1129]), .Z(n4769) );
  OR U4931 ( .A(n4767), .B(n4766), .Z(n4768) );
  AND U4932 ( .A(n4769), .B(n4768), .Z(n4807) );
  XOR U4933 ( .A(n4808), .B(n4807), .Z(c[1130]) );
  NANDN U4934 ( .A(n4771), .B(n4770), .Z(n4775) );
  NAND U4935 ( .A(n4773), .B(n4772), .Z(n4774) );
  NAND U4936 ( .A(n4775), .B(n4774), .Z(n4814) );
  NAND U4937 ( .A(b[0]), .B(a[115]), .Z(n4776) );
  XNOR U4938 ( .A(b[1]), .B(n4776), .Z(n4778) );
  NAND U4939 ( .A(n31), .B(a[114]), .Z(n4777) );
  AND U4940 ( .A(n4778), .B(n4777), .Z(n4831) );
  XOR U4941 ( .A(a[111]), .B(n42197), .Z(n4820) );
  NANDN U4942 ( .A(n4820), .B(n42173), .Z(n4781) );
  NANDN U4943 ( .A(n4779), .B(n42172), .Z(n4780) );
  NAND U4944 ( .A(n4781), .B(n4780), .Z(n4829) );
  NAND U4945 ( .A(b[7]), .B(a[107]), .Z(n4830) );
  XNOR U4946 ( .A(n4829), .B(n4830), .Z(n4832) );
  XOR U4947 ( .A(n4831), .B(n4832), .Z(n4838) );
  NANDN U4948 ( .A(n4782), .B(n42093), .Z(n4784) );
  XOR U4949 ( .A(n42134), .B(a[113]), .Z(n4823) );
  NANDN U4950 ( .A(n4823), .B(n42095), .Z(n4783) );
  NAND U4951 ( .A(n4784), .B(n4783), .Z(n4836) );
  NANDN U4952 ( .A(n4785), .B(n42231), .Z(n4787) );
  XOR U4953 ( .A(n171), .B(a[109]), .Z(n4826) );
  NANDN U4954 ( .A(n4826), .B(n42234), .Z(n4786) );
  AND U4955 ( .A(n4787), .B(n4786), .Z(n4835) );
  XNOR U4956 ( .A(n4836), .B(n4835), .Z(n4837) );
  XNOR U4957 ( .A(n4838), .B(n4837), .Z(n4842) );
  NANDN U4958 ( .A(n4789), .B(n4788), .Z(n4793) );
  NAND U4959 ( .A(n4791), .B(n4790), .Z(n4792) );
  AND U4960 ( .A(n4793), .B(n4792), .Z(n4841) );
  XOR U4961 ( .A(n4842), .B(n4841), .Z(n4843) );
  NANDN U4962 ( .A(n4795), .B(n4794), .Z(n4799) );
  NANDN U4963 ( .A(n4797), .B(n4796), .Z(n4798) );
  NAND U4964 ( .A(n4799), .B(n4798), .Z(n4844) );
  XOR U4965 ( .A(n4843), .B(n4844), .Z(n4811) );
  OR U4966 ( .A(n4801), .B(n4800), .Z(n4805) );
  NANDN U4967 ( .A(n4803), .B(n4802), .Z(n4804) );
  NAND U4968 ( .A(n4805), .B(n4804), .Z(n4812) );
  XNOR U4969 ( .A(n4811), .B(n4812), .Z(n4813) );
  XNOR U4970 ( .A(n4814), .B(n4813), .Z(n4847) );
  XNOR U4971 ( .A(n4847), .B(sreg[1131]), .Z(n4849) );
  NAND U4972 ( .A(n4806), .B(sreg[1130]), .Z(n4810) );
  OR U4973 ( .A(n4808), .B(n4807), .Z(n4809) );
  AND U4974 ( .A(n4810), .B(n4809), .Z(n4848) );
  XOR U4975 ( .A(n4849), .B(n4848), .Z(c[1131]) );
  NANDN U4976 ( .A(n4812), .B(n4811), .Z(n4816) );
  NAND U4977 ( .A(n4814), .B(n4813), .Z(n4815) );
  NAND U4978 ( .A(n4816), .B(n4815), .Z(n4855) );
  NAND U4979 ( .A(b[0]), .B(a[116]), .Z(n4817) );
  XNOR U4980 ( .A(b[1]), .B(n4817), .Z(n4819) );
  NAND U4981 ( .A(n31), .B(a[115]), .Z(n4818) );
  AND U4982 ( .A(n4819), .B(n4818), .Z(n4872) );
  XOR U4983 ( .A(a[112]), .B(n42197), .Z(n4861) );
  NANDN U4984 ( .A(n4861), .B(n42173), .Z(n4822) );
  NANDN U4985 ( .A(n4820), .B(n42172), .Z(n4821) );
  NAND U4986 ( .A(n4822), .B(n4821), .Z(n4870) );
  NAND U4987 ( .A(b[7]), .B(a[108]), .Z(n4871) );
  XNOR U4988 ( .A(n4870), .B(n4871), .Z(n4873) );
  XOR U4989 ( .A(n4872), .B(n4873), .Z(n4879) );
  NANDN U4990 ( .A(n4823), .B(n42093), .Z(n4825) );
  XOR U4991 ( .A(n42134), .B(a[114]), .Z(n4864) );
  NANDN U4992 ( .A(n4864), .B(n42095), .Z(n4824) );
  NAND U4993 ( .A(n4825), .B(n4824), .Z(n4877) );
  NANDN U4994 ( .A(n4826), .B(n42231), .Z(n4828) );
  XOR U4995 ( .A(n171), .B(a[110]), .Z(n4867) );
  NANDN U4996 ( .A(n4867), .B(n42234), .Z(n4827) );
  AND U4997 ( .A(n4828), .B(n4827), .Z(n4876) );
  XNOR U4998 ( .A(n4877), .B(n4876), .Z(n4878) );
  XNOR U4999 ( .A(n4879), .B(n4878), .Z(n4883) );
  NANDN U5000 ( .A(n4830), .B(n4829), .Z(n4834) );
  NAND U5001 ( .A(n4832), .B(n4831), .Z(n4833) );
  AND U5002 ( .A(n4834), .B(n4833), .Z(n4882) );
  XOR U5003 ( .A(n4883), .B(n4882), .Z(n4884) );
  NANDN U5004 ( .A(n4836), .B(n4835), .Z(n4840) );
  NANDN U5005 ( .A(n4838), .B(n4837), .Z(n4839) );
  NAND U5006 ( .A(n4840), .B(n4839), .Z(n4885) );
  XOR U5007 ( .A(n4884), .B(n4885), .Z(n4852) );
  OR U5008 ( .A(n4842), .B(n4841), .Z(n4846) );
  NANDN U5009 ( .A(n4844), .B(n4843), .Z(n4845) );
  NAND U5010 ( .A(n4846), .B(n4845), .Z(n4853) );
  XNOR U5011 ( .A(n4852), .B(n4853), .Z(n4854) );
  XNOR U5012 ( .A(n4855), .B(n4854), .Z(n4888) );
  XNOR U5013 ( .A(n4888), .B(sreg[1132]), .Z(n4890) );
  NAND U5014 ( .A(n4847), .B(sreg[1131]), .Z(n4851) );
  OR U5015 ( .A(n4849), .B(n4848), .Z(n4850) );
  AND U5016 ( .A(n4851), .B(n4850), .Z(n4889) );
  XOR U5017 ( .A(n4890), .B(n4889), .Z(c[1132]) );
  NANDN U5018 ( .A(n4853), .B(n4852), .Z(n4857) );
  NAND U5019 ( .A(n4855), .B(n4854), .Z(n4856) );
  NAND U5020 ( .A(n4857), .B(n4856), .Z(n4896) );
  NAND U5021 ( .A(b[0]), .B(a[117]), .Z(n4858) );
  XNOR U5022 ( .A(b[1]), .B(n4858), .Z(n4860) );
  NAND U5023 ( .A(n31), .B(a[116]), .Z(n4859) );
  AND U5024 ( .A(n4860), .B(n4859), .Z(n4913) );
  XOR U5025 ( .A(a[113]), .B(n42197), .Z(n4902) );
  NANDN U5026 ( .A(n4902), .B(n42173), .Z(n4863) );
  NANDN U5027 ( .A(n4861), .B(n42172), .Z(n4862) );
  NAND U5028 ( .A(n4863), .B(n4862), .Z(n4911) );
  NAND U5029 ( .A(b[7]), .B(a[109]), .Z(n4912) );
  XNOR U5030 ( .A(n4911), .B(n4912), .Z(n4914) );
  XOR U5031 ( .A(n4913), .B(n4914), .Z(n4920) );
  NANDN U5032 ( .A(n4864), .B(n42093), .Z(n4866) );
  XOR U5033 ( .A(n42134), .B(a[115]), .Z(n4905) );
  NANDN U5034 ( .A(n4905), .B(n42095), .Z(n4865) );
  NAND U5035 ( .A(n4866), .B(n4865), .Z(n4918) );
  NANDN U5036 ( .A(n4867), .B(n42231), .Z(n4869) );
  XOR U5037 ( .A(n171), .B(a[111]), .Z(n4908) );
  NANDN U5038 ( .A(n4908), .B(n42234), .Z(n4868) );
  AND U5039 ( .A(n4869), .B(n4868), .Z(n4917) );
  XNOR U5040 ( .A(n4918), .B(n4917), .Z(n4919) );
  XNOR U5041 ( .A(n4920), .B(n4919), .Z(n4924) );
  NANDN U5042 ( .A(n4871), .B(n4870), .Z(n4875) );
  NAND U5043 ( .A(n4873), .B(n4872), .Z(n4874) );
  AND U5044 ( .A(n4875), .B(n4874), .Z(n4923) );
  XOR U5045 ( .A(n4924), .B(n4923), .Z(n4925) );
  NANDN U5046 ( .A(n4877), .B(n4876), .Z(n4881) );
  NANDN U5047 ( .A(n4879), .B(n4878), .Z(n4880) );
  NAND U5048 ( .A(n4881), .B(n4880), .Z(n4926) );
  XOR U5049 ( .A(n4925), .B(n4926), .Z(n4893) );
  OR U5050 ( .A(n4883), .B(n4882), .Z(n4887) );
  NANDN U5051 ( .A(n4885), .B(n4884), .Z(n4886) );
  NAND U5052 ( .A(n4887), .B(n4886), .Z(n4894) );
  XNOR U5053 ( .A(n4893), .B(n4894), .Z(n4895) );
  XNOR U5054 ( .A(n4896), .B(n4895), .Z(n4929) );
  XNOR U5055 ( .A(n4929), .B(sreg[1133]), .Z(n4931) );
  NAND U5056 ( .A(n4888), .B(sreg[1132]), .Z(n4892) );
  OR U5057 ( .A(n4890), .B(n4889), .Z(n4891) );
  AND U5058 ( .A(n4892), .B(n4891), .Z(n4930) );
  XOR U5059 ( .A(n4931), .B(n4930), .Z(c[1133]) );
  NANDN U5060 ( .A(n4894), .B(n4893), .Z(n4898) );
  NAND U5061 ( .A(n4896), .B(n4895), .Z(n4897) );
  NAND U5062 ( .A(n4898), .B(n4897), .Z(n4937) );
  NAND U5063 ( .A(b[0]), .B(a[118]), .Z(n4899) );
  XNOR U5064 ( .A(b[1]), .B(n4899), .Z(n4901) );
  NAND U5065 ( .A(n31), .B(a[117]), .Z(n4900) );
  AND U5066 ( .A(n4901), .B(n4900), .Z(n4954) );
  XOR U5067 ( .A(a[114]), .B(n42197), .Z(n4943) );
  NANDN U5068 ( .A(n4943), .B(n42173), .Z(n4904) );
  NANDN U5069 ( .A(n4902), .B(n42172), .Z(n4903) );
  NAND U5070 ( .A(n4904), .B(n4903), .Z(n4952) );
  NAND U5071 ( .A(b[7]), .B(a[110]), .Z(n4953) );
  XNOR U5072 ( .A(n4952), .B(n4953), .Z(n4955) );
  XOR U5073 ( .A(n4954), .B(n4955), .Z(n4961) );
  NANDN U5074 ( .A(n4905), .B(n42093), .Z(n4907) );
  XOR U5075 ( .A(n42134), .B(a[116]), .Z(n4946) );
  NANDN U5076 ( .A(n4946), .B(n42095), .Z(n4906) );
  NAND U5077 ( .A(n4907), .B(n4906), .Z(n4959) );
  NANDN U5078 ( .A(n4908), .B(n42231), .Z(n4910) );
  XOR U5079 ( .A(n171), .B(a[112]), .Z(n4949) );
  NANDN U5080 ( .A(n4949), .B(n42234), .Z(n4909) );
  AND U5081 ( .A(n4910), .B(n4909), .Z(n4958) );
  XNOR U5082 ( .A(n4959), .B(n4958), .Z(n4960) );
  XNOR U5083 ( .A(n4961), .B(n4960), .Z(n4965) );
  NANDN U5084 ( .A(n4912), .B(n4911), .Z(n4916) );
  NAND U5085 ( .A(n4914), .B(n4913), .Z(n4915) );
  AND U5086 ( .A(n4916), .B(n4915), .Z(n4964) );
  XOR U5087 ( .A(n4965), .B(n4964), .Z(n4966) );
  NANDN U5088 ( .A(n4918), .B(n4917), .Z(n4922) );
  NANDN U5089 ( .A(n4920), .B(n4919), .Z(n4921) );
  NAND U5090 ( .A(n4922), .B(n4921), .Z(n4967) );
  XOR U5091 ( .A(n4966), .B(n4967), .Z(n4934) );
  OR U5092 ( .A(n4924), .B(n4923), .Z(n4928) );
  NANDN U5093 ( .A(n4926), .B(n4925), .Z(n4927) );
  NAND U5094 ( .A(n4928), .B(n4927), .Z(n4935) );
  XNOR U5095 ( .A(n4934), .B(n4935), .Z(n4936) );
  XNOR U5096 ( .A(n4937), .B(n4936), .Z(n4970) );
  XNOR U5097 ( .A(n4970), .B(sreg[1134]), .Z(n4972) );
  NAND U5098 ( .A(n4929), .B(sreg[1133]), .Z(n4933) );
  OR U5099 ( .A(n4931), .B(n4930), .Z(n4932) );
  AND U5100 ( .A(n4933), .B(n4932), .Z(n4971) );
  XOR U5101 ( .A(n4972), .B(n4971), .Z(c[1134]) );
  NANDN U5102 ( .A(n4935), .B(n4934), .Z(n4939) );
  NAND U5103 ( .A(n4937), .B(n4936), .Z(n4938) );
  NAND U5104 ( .A(n4939), .B(n4938), .Z(n4978) );
  NAND U5105 ( .A(b[0]), .B(a[119]), .Z(n4940) );
  XNOR U5106 ( .A(b[1]), .B(n4940), .Z(n4942) );
  NAND U5107 ( .A(n32), .B(a[118]), .Z(n4941) );
  AND U5108 ( .A(n4942), .B(n4941), .Z(n4995) );
  XOR U5109 ( .A(a[115]), .B(n42197), .Z(n4984) );
  NANDN U5110 ( .A(n4984), .B(n42173), .Z(n4945) );
  NANDN U5111 ( .A(n4943), .B(n42172), .Z(n4944) );
  NAND U5112 ( .A(n4945), .B(n4944), .Z(n4993) );
  NAND U5113 ( .A(b[7]), .B(a[111]), .Z(n4994) );
  XNOR U5114 ( .A(n4993), .B(n4994), .Z(n4996) );
  XOR U5115 ( .A(n4995), .B(n4996), .Z(n5002) );
  NANDN U5116 ( .A(n4946), .B(n42093), .Z(n4948) );
  XOR U5117 ( .A(n42134), .B(a[117]), .Z(n4987) );
  NANDN U5118 ( .A(n4987), .B(n42095), .Z(n4947) );
  NAND U5119 ( .A(n4948), .B(n4947), .Z(n5000) );
  NANDN U5120 ( .A(n4949), .B(n42231), .Z(n4951) );
  XOR U5121 ( .A(n171), .B(a[113]), .Z(n4990) );
  NANDN U5122 ( .A(n4990), .B(n42234), .Z(n4950) );
  AND U5123 ( .A(n4951), .B(n4950), .Z(n4999) );
  XNOR U5124 ( .A(n5000), .B(n4999), .Z(n5001) );
  XNOR U5125 ( .A(n5002), .B(n5001), .Z(n5006) );
  NANDN U5126 ( .A(n4953), .B(n4952), .Z(n4957) );
  NAND U5127 ( .A(n4955), .B(n4954), .Z(n4956) );
  AND U5128 ( .A(n4957), .B(n4956), .Z(n5005) );
  XOR U5129 ( .A(n5006), .B(n5005), .Z(n5007) );
  NANDN U5130 ( .A(n4959), .B(n4958), .Z(n4963) );
  NANDN U5131 ( .A(n4961), .B(n4960), .Z(n4962) );
  NAND U5132 ( .A(n4963), .B(n4962), .Z(n5008) );
  XOR U5133 ( .A(n5007), .B(n5008), .Z(n4975) );
  OR U5134 ( .A(n4965), .B(n4964), .Z(n4969) );
  NANDN U5135 ( .A(n4967), .B(n4966), .Z(n4968) );
  NAND U5136 ( .A(n4969), .B(n4968), .Z(n4976) );
  XNOR U5137 ( .A(n4975), .B(n4976), .Z(n4977) );
  XNOR U5138 ( .A(n4978), .B(n4977), .Z(n5011) );
  XNOR U5139 ( .A(n5011), .B(sreg[1135]), .Z(n5013) );
  NAND U5140 ( .A(n4970), .B(sreg[1134]), .Z(n4974) );
  OR U5141 ( .A(n4972), .B(n4971), .Z(n4973) );
  AND U5142 ( .A(n4974), .B(n4973), .Z(n5012) );
  XOR U5143 ( .A(n5013), .B(n5012), .Z(c[1135]) );
  NANDN U5144 ( .A(n4976), .B(n4975), .Z(n4980) );
  NAND U5145 ( .A(n4978), .B(n4977), .Z(n4979) );
  NAND U5146 ( .A(n4980), .B(n4979), .Z(n5019) );
  NAND U5147 ( .A(b[0]), .B(a[120]), .Z(n4981) );
  XNOR U5148 ( .A(b[1]), .B(n4981), .Z(n4983) );
  NAND U5149 ( .A(n32), .B(a[119]), .Z(n4982) );
  AND U5150 ( .A(n4983), .B(n4982), .Z(n5036) );
  XOR U5151 ( .A(a[116]), .B(n42197), .Z(n5025) );
  NANDN U5152 ( .A(n5025), .B(n42173), .Z(n4986) );
  NANDN U5153 ( .A(n4984), .B(n42172), .Z(n4985) );
  NAND U5154 ( .A(n4986), .B(n4985), .Z(n5034) );
  NAND U5155 ( .A(b[7]), .B(a[112]), .Z(n5035) );
  XNOR U5156 ( .A(n5034), .B(n5035), .Z(n5037) );
  XOR U5157 ( .A(n5036), .B(n5037), .Z(n5043) );
  NANDN U5158 ( .A(n4987), .B(n42093), .Z(n4989) );
  XOR U5159 ( .A(n42134), .B(a[118]), .Z(n5028) );
  NANDN U5160 ( .A(n5028), .B(n42095), .Z(n4988) );
  NAND U5161 ( .A(n4989), .B(n4988), .Z(n5041) );
  NANDN U5162 ( .A(n4990), .B(n42231), .Z(n4992) );
  XOR U5163 ( .A(n171), .B(a[114]), .Z(n5031) );
  NANDN U5164 ( .A(n5031), .B(n42234), .Z(n4991) );
  AND U5165 ( .A(n4992), .B(n4991), .Z(n5040) );
  XNOR U5166 ( .A(n5041), .B(n5040), .Z(n5042) );
  XNOR U5167 ( .A(n5043), .B(n5042), .Z(n5047) );
  NANDN U5168 ( .A(n4994), .B(n4993), .Z(n4998) );
  NAND U5169 ( .A(n4996), .B(n4995), .Z(n4997) );
  AND U5170 ( .A(n4998), .B(n4997), .Z(n5046) );
  XOR U5171 ( .A(n5047), .B(n5046), .Z(n5048) );
  NANDN U5172 ( .A(n5000), .B(n4999), .Z(n5004) );
  NANDN U5173 ( .A(n5002), .B(n5001), .Z(n5003) );
  NAND U5174 ( .A(n5004), .B(n5003), .Z(n5049) );
  XOR U5175 ( .A(n5048), .B(n5049), .Z(n5016) );
  OR U5176 ( .A(n5006), .B(n5005), .Z(n5010) );
  NANDN U5177 ( .A(n5008), .B(n5007), .Z(n5009) );
  NAND U5178 ( .A(n5010), .B(n5009), .Z(n5017) );
  XNOR U5179 ( .A(n5016), .B(n5017), .Z(n5018) );
  XNOR U5180 ( .A(n5019), .B(n5018), .Z(n5052) );
  XNOR U5181 ( .A(n5052), .B(sreg[1136]), .Z(n5054) );
  NAND U5182 ( .A(n5011), .B(sreg[1135]), .Z(n5015) );
  OR U5183 ( .A(n5013), .B(n5012), .Z(n5014) );
  AND U5184 ( .A(n5015), .B(n5014), .Z(n5053) );
  XOR U5185 ( .A(n5054), .B(n5053), .Z(c[1136]) );
  NANDN U5186 ( .A(n5017), .B(n5016), .Z(n5021) );
  NAND U5187 ( .A(n5019), .B(n5018), .Z(n5020) );
  NAND U5188 ( .A(n5021), .B(n5020), .Z(n5060) );
  NAND U5189 ( .A(b[0]), .B(a[121]), .Z(n5022) );
  XNOR U5190 ( .A(b[1]), .B(n5022), .Z(n5024) );
  NAND U5191 ( .A(n32), .B(a[120]), .Z(n5023) );
  AND U5192 ( .A(n5024), .B(n5023), .Z(n5077) );
  XOR U5193 ( .A(a[117]), .B(n42197), .Z(n5066) );
  NANDN U5194 ( .A(n5066), .B(n42173), .Z(n5027) );
  NANDN U5195 ( .A(n5025), .B(n42172), .Z(n5026) );
  NAND U5196 ( .A(n5027), .B(n5026), .Z(n5075) );
  NAND U5197 ( .A(b[7]), .B(a[113]), .Z(n5076) );
  XNOR U5198 ( .A(n5075), .B(n5076), .Z(n5078) );
  XOR U5199 ( .A(n5077), .B(n5078), .Z(n5084) );
  NANDN U5200 ( .A(n5028), .B(n42093), .Z(n5030) );
  XOR U5201 ( .A(n42134), .B(a[119]), .Z(n5069) );
  NANDN U5202 ( .A(n5069), .B(n42095), .Z(n5029) );
  NAND U5203 ( .A(n5030), .B(n5029), .Z(n5082) );
  NANDN U5204 ( .A(n5031), .B(n42231), .Z(n5033) );
  XOR U5205 ( .A(n171), .B(a[115]), .Z(n5072) );
  NANDN U5206 ( .A(n5072), .B(n42234), .Z(n5032) );
  AND U5207 ( .A(n5033), .B(n5032), .Z(n5081) );
  XNOR U5208 ( .A(n5082), .B(n5081), .Z(n5083) );
  XNOR U5209 ( .A(n5084), .B(n5083), .Z(n5088) );
  NANDN U5210 ( .A(n5035), .B(n5034), .Z(n5039) );
  NAND U5211 ( .A(n5037), .B(n5036), .Z(n5038) );
  AND U5212 ( .A(n5039), .B(n5038), .Z(n5087) );
  XOR U5213 ( .A(n5088), .B(n5087), .Z(n5089) );
  NANDN U5214 ( .A(n5041), .B(n5040), .Z(n5045) );
  NANDN U5215 ( .A(n5043), .B(n5042), .Z(n5044) );
  NAND U5216 ( .A(n5045), .B(n5044), .Z(n5090) );
  XOR U5217 ( .A(n5089), .B(n5090), .Z(n5057) );
  OR U5218 ( .A(n5047), .B(n5046), .Z(n5051) );
  NANDN U5219 ( .A(n5049), .B(n5048), .Z(n5050) );
  NAND U5220 ( .A(n5051), .B(n5050), .Z(n5058) );
  XNOR U5221 ( .A(n5057), .B(n5058), .Z(n5059) );
  XNOR U5222 ( .A(n5060), .B(n5059), .Z(n5093) );
  XNOR U5223 ( .A(n5093), .B(sreg[1137]), .Z(n5095) );
  NAND U5224 ( .A(n5052), .B(sreg[1136]), .Z(n5056) );
  OR U5225 ( .A(n5054), .B(n5053), .Z(n5055) );
  AND U5226 ( .A(n5056), .B(n5055), .Z(n5094) );
  XOR U5227 ( .A(n5095), .B(n5094), .Z(c[1137]) );
  NANDN U5228 ( .A(n5058), .B(n5057), .Z(n5062) );
  NAND U5229 ( .A(n5060), .B(n5059), .Z(n5061) );
  NAND U5230 ( .A(n5062), .B(n5061), .Z(n5101) );
  NAND U5231 ( .A(b[0]), .B(a[122]), .Z(n5063) );
  XNOR U5232 ( .A(b[1]), .B(n5063), .Z(n5065) );
  NAND U5233 ( .A(n32), .B(a[121]), .Z(n5064) );
  AND U5234 ( .A(n5065), .B(n5064), .Z(n5118) );
  XOR U5235 ( .A(a[118]), .B(n42197), .Z(n5107) );
  NANDN U5236 ( .A(n5107), .B(n42173), .Z(n5068) );
  NANDN U5237 ( .A(n5066), .B(n42172), .Z(n5067) );
  NAND U5238 ( .A(n5068), .B(n5067), .Z(n5116) );
  NAND U5239 ( .A(b[7]), .B(a[114]), .Z(n5117) );
  XNOR U5240 ( .A(n5116), .B(n5117), .Z(n5119) );
  XOR U5241 ( .A(n5118), .B(n5119), .Z(n5125) );
  NANDN U5242 ( .A(n5069), .B(n42093), .Z(n5071) );
  XOR U5243 ( .A(n42134), .B(a[120]), .Z(n5110) );
  NANDN U5244 ( .A(n5110), .B(n42095), .Z(n5070) );
  NAND U5245 ( .A(n5071), .B(n5070), .Z(n5123) );
  NANDN U5246 ( .A(n5072), .B(n42231), .Z(n5074) );
  XOR U5247 ( .A(n171), .B(a[116]), .Z(n5113) );
  NANDN U5248 ( .A(n5113), .B(n42234), .Z(n5073) );
  AND U5249 ( .A(n5074), .B(n5073), .Z(n5122) );
  XNOR U5250 ( .A(n5123), .B(n5122), .Z(n5124) );
  XNOR U5251 ( .A(n5125), .B(n5124), .Z(n5129) );
  NANDN U5252 ( .A(n5076), .B(n5075), .Z(n5080) );
  NAND U5253 ( .A(n5078), .B(n5077), .Z(n5079) );
  AND U5254 ( .A(n5080), .B(n5079), .Z(n5128) );
  XOR U5255 ( .A(n5129), .B(n5128), .Z(n5130) );
  NANDN U5256 ( .A(n5082), .B(n5081), .Z(n5086) );
  NANDN U5257 ( .A(n5084), .B(n5083), .Z(n5085) );
  NAND U5258 ( .A(n5086), .B(n5085), .Z(n5131) );
  XOR U5259 ( .A(n5130), .B(n5131), .Z(n5098) );
  OR U5260 ( .A(n5088), .B(n5087), .Z(n5092) );
  NANDN U5261 ( .A(n5090), .B(n5089), .Z(n5091) );
  NAND U5262 ( .A(n5092), .B(n5091), .Z(n5099) );
  XNOR U5263 ( .A(n5098), .B(n5099), .Z(n5100) );
  XNOR U5264 ( .A(n5101), .B(n5100), .Z(n5134) );
  XNOR U5265 ( .A(n5134), .B(sreg[1138]), .Z(n5136) );
  NAND U5266 ( .A(n5093), .B(sreg[1137]), .Z(n5097) );
  OR U5267 ( .A(n5095), .B(n5094), .Z(n5096) );
  AND U5268 ( .A(n5097), .B(n5096), .Z(n5135) );
  XOR U5269 ( .A(n5136), .B(n5135), .Z(c[1138]) );
  NANDN U5270 ( .A(n5099), .B(n5098), .Z(n5103) );
  NAND U5271 ( .A(n5101), .B(n5100), .Z(n5102) );
  NAND U5272 ( .A(n5103), .B(n5102), .Z(n5142) );
  NAND U5273 ( .A(b[0]), .B(a[123]), .Z(n5104) );
  XNOR U5274 ( .A(b[1]), .B(n5104), .Z(n5106) );
  NAND U5275 ( .A(n32), .B(a[122]), .Z(n5105) );
  AND U5276 ( .A(n5106), .B(n5105), .Z(n5159) );
  XOR U5277 ( .A(a[119]), .B(n42197), .Z(n5148) );
  NANDN U5278 ( .A(n5148), .B(n42173), .Z(n5109) );
  NANDN U5279 ( .A(n5107), .B(n42172), .Z(n5108) );
  NAND U5280 ( .A(n5109), .B(n5108), .Z(n5157) );
  NAND U5281 ( .A(b[7]), .B(a[115]), .Z(n5158) );
  XNOR U5282 ( .A(n5157), .B(n5158), .Z(n5160) );
  XOR U5283 ( .A(n5159), .B(n5160), .Z(n5166) );
  NANDN U5284 ( .A(n5110), .B(n42093), .Z(n5112) );
  XOR U5285 ( .A(n42134), .B(a[121]), .Z(n5151) );
  NANDN U5286 ( .A(n5151), .B(n42095), .Z(n5111) );
  NAND U5287 ( .A(n5112), .B(n5111), .Z(n5164) );
  NANDN U5288 ( .A(n5113), .B(n42231), .Z(n5115) );
  XOR U5289 ( .A(n171), .B(a[117]), .Z(n5154) );
  NANDN U5290 ( .A(n5154), .B(n42234), .Z(n5114) );
  AND U5291 ( .A(n5115), .B(n5114), .Z(n5163) );
  XNOR U5292 ( .A(n5164), .B(n5163), .Z(n5165) );
  XNOR U5293 ( .A(n5166), .B(n5165), .Z(n5170) );
  NANDN U5294 ( .A(n5117), .B(n5116), .Z(n5121) );
  NAND U5295 ( .A(n5119), .B(n5118), .Z(n5120) );
  AND U5296 ( .A(n5121), .B(n5120), .Z(n5169) );
  XOR U5297 ( .A(n5170), .B(n5169), .Z(n5171) );
  NANDN U5298 ( .A(n5123), .B(n5122), .Z(n5127) );
  NANDN U5299 ( .A(n5125), .B(n5124), .Z(n5126) );
  NAND U5300 ( .A(n5127), .B(n5126), .Z(n5172) );
  XOR U5301 ( .A(n5171), .B(n5172), .Z(n5139) );
  OR U5302 ( .A(n5129), .B(n5128), .Z(n5133) );
  NANDN U5303 ( .A(n5131), .B(n5130), .Z(n5132) );
  NAND U5304 ( .A(n5133), .B(n5132), .Z(n5140) );
  XNOR U5305 ( .A(n5139), .B(n5140), .Z(n5141) );
  XNOR U5306 ( .A(n5142), .B(n5141), .Z(n5175) );
  XNOR U5307 ( .A(n5175), .B(sreg[1139]), .Z(n5177) );
  NAND U5308 ( .A(n5134), .B(sreg[1138]), .Z(n5138) );
  OR U5309 ( .A(n5136), .B(n5135), .Z(n5137) );
  AND U5310 ( .A(n5138), .B(n5137), .Z(n5176) );
  XOR U5311 ( .A(n5177), .B(n5176), .Z(c[1139]) );
  NANDN U5312 ( .A(n5140), .B(n5139), .Z(n5144) );
  NAND U5313 ( .A(n5142), .B(n5141), .Z(n5143) );
  NAND U5314 ( .A(n5144), .B(n5143), .Z(n5183) );
  NAND U5315 ( .A(b[0]), .B(a[124]), .Z(n5145) );
  XNOR U5316 ( .A(b[1]), .B(n5145), .Z(n5147) );
  NAND U5317 ( .A(n32), .B(a[123]), .Z(n5146) );
  AND U5318 ( .A(n5147), .B(n5146), .Z(n5200) );
  XOR U5319 ( .A(a[120]), .B(n42197), .Z(n5189) );
  NANDN U5320 ( .A(n5189), .B(n42173), .Z(n5150) );
  NANDN U5321 ( .A(n5148), .B(n42172), .Z(n5149) );
  NAND U5322 ( .A(n5150), .B(n5149), .Z(n5198) );
  NAND U5323 ( .A(b[7]), .B(a[116]), .Z(n5199) );
  XNOR U5324 ( .A(n5198), .B(n5199), .Z(n5201) );
  XOR U5325 ( .A(n5200), .B(n5201), .Z(n5207) );
  NANDN U5326 ( .A(n5151), .B(n42093), .Z(n5153) );
  XOR U5327 ( .A(n42134), .B(a[122]), .Z(n5192) );
  NANDN U5328 ( .A(n5192), .B(n42095), .Z(n5152) );
  NAND U5329 ( .A(n5153), .B(n5152), .Z(n5205) );
  NANDN U5330 ( .A(n5154), .B(n42231), .Z(n5156) );
  XOR U5331 ( .A(n171), .B(a[118]), .Z(n5195) );
  NANDN U5332 ( .A(n5195), .B(n42234), .Z(n5155) );
  AND U5333 ( .A(n5156), .B(n5155), .Z(n5204) );
  XNOR U5334 ( .A(n5205), .B(n5204), .Z(n5206) );
  XNOR U5335 ( .A(n5207), .B(n5206), .Z(n5211) );
  NANDN U5336 ( .A(n5158), .B(n5157), .Z(n5162) );
  NAND U5337 ( .A(n5160), .B(n5159), .Z(n5161) );
  AND U5338 ( .A(n5162), .B(n5161), .Z(n5210) );
  XOR U5339 ( .A(n5211), .B(n5210), .Z(n5212) );
  NANDN U5340 ( .A(n5164), .B(n5163), .Z(n5168) );
  NANDN U5341 ( .A(n5166), .B(n5165), .Z(n5167) );
  NAND U5342 ( .A(n5168), .B(n5167), .Z(n5213) );
  XOR U5343 ( .A(n5212), .B(n5213), .Z(n5180) );
  OR U5344 ( .A(n5170), .B(n5169), .Z(n5174) );
  NANDN U5345 ( .A(n5172), .B(n5171), .Z(n5173) );
  NAND U5346 ( .A(n5174), .B(n5173), .Z(n5181) );
  XNOR U5347 ( .A(n5180), .B(n5181), .Z(n5182) );
  XNOR U5348 ( .A(n5183), .B(n5182), .Z(n5216) );
  XNOR U5349 ( .A(n5216), .B(sreg[1140]), .Z(n5218) );
  NAND U5350 ( .A(n5175), .B(sreg[1139]), .Z(n5179) );
  OR U5351 ( .A(n5177), .B(n5176), .Z(n5178) );
  AND U5352 ( .A(n5179), .B(n5178), .Z(n5217) );
  XOR U5353 ( .A(n5218), .B(n5217), .Z(c[1140]) );
  NANDN U5354 ( .A(n5181), .B(n5180), .Z(n5185) );
  NAND U5355 ( .A(n5183), .B(n5182), .Z(n5184) );
  NAND U5356 ( .A(n5185), .B(n5184), .Z(n5224) );
  NAND U5357 ( .A(b[0]), .B(a[125]), .Z(n5186) );
  XNOR U5358 ( .A(b[1]), .B(n5186), .Z(n5188) );
  NAND U5359 ( .A(n32), .B(a[124]), .Z(n5187) );
  AND U5360 ( .A(n5188), .B(n5187), .Z(n5241) );
  XOR U5361 ( .A(a[121]), .B(n42197), .Z(n5230) );
  NANDN U5362 ( .A(n5230), .B(n42173), .Z(n5191) );
  NANDN U5363 ( .A(n5189), .B(n42172), .Z(n5190) );
  NAND U5364 ( .A(n5191), .B(n5190), .Z(n5239) );
  NAND U5365 ( .A(b[7]), .B(a[117]), .Z(n5240) );
  XNOR U5366 ( .A(n5239), .B(n5240), .Z(n5242) );
  XOR U5367 ( .A(n5241), .B(n5242), .Z(n5248) );
  NANDN U5368 ( .A(n5192), .B(n42093), .Z(n5194) );
  XOR U5369 ( .A(n42134), .B(a[123]), .Z(n5233) );
  NANDN U5370 ( .A(n5233), .B(n42095), .Z(n5193) );
  NAND U5371 ( .A(n5194), .B(n5193), .Z(n5246) );
  NANDN U5372 ( .A(n5195), .B(n42231), .Z(n5197) );
  XOR U5373 ( .A(n172), .B(a[119]), .Z(n5236) );
  NANDN U5374 ( .A(n5236), .B(n42234), .Z(n5196) );
  AND U5375 ( .A(n5197), .B(n5196), .Z(n5245) );
  XNOR U5376 ( .A(n5246), .B(n5245), .Z(n5247) );
  XNOR U5377 ( .A(n5248), .B(n5247), .Z(n5252) );
  NANDN U5378 ( .A(n5199), .B(n5198), .Z(n5203) );
  NAND U5379 ( .A(n5201), .B(n5200), .Z(n5202) );
  AND U5380 ( .A(n5203), .B(n5202), .Z(n5251) );
  XOR U5381 ( .A(n5252), .B(n5251), .Z(n5253) );
  NANDN U5382 ( .A(n5205), .B(n5204), .Z(n5209) );
  NANDN U5383 ( .A(n5207), .B(n5206), .Z(n5208) );
  NAND U5384 ( .A(n5209), .B(n5208), .Z(n5254) );
  XOR U5385 ( .A(n5253), .B(n5254), .Z(n5221) );
  OR U5386 ( .A(n5211), .B(n5210), .Z(n5215) );
  NANDN U5387 ( .A(n5213), .B(n5212), .Z(n5214) );
  NAND U5388 ( .A(n5215), .B(n5214), .Z(n5222) );
  XNOR U5389 ( .A(n5221), .B(n5222), .Z(n5223) );
  XNOR U5390 ( .A(n5224), .B(n5223), .Z(n5257) );
  XNOR U5391 ( .A(n5257), .B(sreg[1141]), .Z(n5259) );
  NAND U5392 ( .A(n5216), .B(sreg[1140]), .Z(n5220) );
  OR U5393 ( .A(n5218), .B(n5217), .Z(n5219) );
  AND U5394 ( .A(n5220), .B(n5219), .Z(n5258) );
  XOR U5395 ( .A(n5259), .B(n5258), .Z(c[1141]) );
  NANDN U5396 ( .A(n5222), .B(n5221), .Z(n5226) );
  NAND U5397 ( .A(n5224), .B(n5223), .Z(n5225) );
  NAND U5398 ( .A(n5226), .B(n5225), .Z(n5265) );
  NAND U5399 ( .A(b[0]), .B(a[126]), .Z(n5227) );
  XNOR U5400 ( .A(b[1]), .B(n5227), .Z(n5229) );
  NAND U5401 ( .A(n33), .B(a[125]), .Z(n5228) );
  AND U5402 ( .A(n5229), .B(n5228), .Z(n5282) );
  XOR U5403 ( .A(a[122]), .B(n42197), .Z(n5271) );
  NANDN U5404 ( .A(n5271), .B(n42173), .Z(n5232) );
  NANDN U5405 ( .A(n5230), .B(n42172), .Z(n5231) );
  NAND U5406 ( .A(n5232), .B(n5231), .Z(n5280) );
  NAND U5407 ( .A(b[7]), .B(a[118]), .Z(n5281) );
  XNOR U5408 ( .A(n5280), .B(n5281), .Z(n5283) );
  XOR U5409 ( .A(n5282), .B(n5283), .Z(n5289) );
  NANDN U5410 ( .A(n5233), .B(n42093), .Z(n5235) );
  XOR U5411 ( .A(n42134), .B(a[124]), .Z(n5274) );
  NANDN U5412 ( .A(n5274), .B(n42095), .Z(n5234) );
  NAND U5413 ( .A(n5235), .B(n5234), .Z(n5287) );
  NANDN U5414 ( .A(n5236), .B(n42231), .Z(n5238) );
  XOR U5415 ( .A(n172), .B(a[120]), .Z(n5277) );
  NANDN U5416 ( .A(n5277), .B(n42234), .Z(n5237) );
  AND U5417 ( .A(n5238), .B(n5237), .Z(n5286) );
  XNOR U5418 ( .A(n5287), .B(n5286), .Z(n5288) );
  XNOR U5419 ( .A(n5289), .B(n5288), .Z(n5293) );
  NANDN U5420 ( .A(n5240), .B(n5239), .Z(n5244) );
  NAND U5421 ( .A(n5242), .B(n5241), .Z(n5243) );
  AND U5422 ( .A(n5244), .B(n5243), .Z(n5292) );
  XOR U5423 ( .A(n5293), .B(n5292), .Z(n5294) );
  NANDN U5424 ( .A(n5246), .B(n5245), .Z(n5250) );
  NANDN U5425 ( .A(n5248), .B(n5247), .Z(n5249) );
  NAND U5426 ( .A(n5250), .B(n5249), .Z(n5295) );
  XOR U5427 ( .A(n5294), .B(n5295), .Z(n5262) );
  OR U5428 ( .A(n5252), .B(n5251), .Z(n5256) );
  NANDN U5429 ( .A(n5254), .B(n5253), .Z(n5255) );
  NAND U5430 ( .A(n5256), .B(n5255), .Z(n5263) );
  XNOR U5431 ( .A(n5262), .B(n5263), .Z(n5264) );
  XNOR U5432 ( .A(n5265), .B(n5264), .Z(n5298) );
  XNOR U5433 ( .A(n5298), .B(sreg[1142]), .Z(n5300) );
  NAND U5434 ( .A(n5257), .B(sreg[1141]), .Z(n5261) );
  OR U5435 ( .A(n5259), .B(n5258), .Z(n5260) );
  AND U5436 ( .A(n5261), .B(n5260), .Z(n5299) );
  XOR U5437 ( .A(n5300), .B(n5299), .Z(c[1142]) );
  NANDN U5438 ( .A(n5263), .B(n5262), .Z(n5267) );
  NAND U5439 ( .A(n5265), .B(n5264), .Z(n5266) );
  NAND U5440 ( .A(n5267), .B(n5266), .Z(n5306) );
  NAND U5441 ( .A(b[0]), .B(a[127]), .Z(n5268) );
  XNOR U5442 ( .A(b[1]), .B(n5268), .Z(n5270) );
  NAND U5443 ( .A(n33), .B(a[126]), .Z(n5269) );
  AND U5444 ( .A(n5270), .B(n5269), .Z(n5323) );
  XOR U5445 ( .A(a[123]), .B(n42197), .Z(n5312) );
  NANDN U5446 ( .A(n5312), .B(n42173), .Z(n5273) );
  NANDN U5447 ( .A(n5271), .B(n42172), .Z(n5272) );
  NAND U5448 ( .A(n5273), .B(n5272), .Z(n5321) );
  NAND U5449 ( .A(b[7]), .B(a[119]), .Z(n5322) );
  XNOR U5450 ( .A(n5321), .B(n5322), .Z(n5324) );
  XOR U5451 ( .A(n5323), .B(n5324), .Z(n5330) );
  NANDN U5452 ( .A(n5274), .B(n42093), .Z(n5276) );
  XOR U5453 ( .A(n42134), .B(a[125]), .Z(n5315) );
  NANDN U5454 ( .A(n5315), .B(n42095), .Z(n5275) );
  NAND U5455 ( .A(n5276), .B(n5275), .Z(n5328) );
  NANDN U5456 ( .A(n5277), .B(n42231), .Z(n5279) );
  XOR U5457 ( .A(n172), .B(a[121]), .Z(n5318) );
  NANDN U5458 ( .A(n5318), .B(n42234), .Z(n5278) );
  AND U5459 ( .A(n5279), .B(n5278), .Z(n5327) );
  XNOR U5460 ( .A(n5328), .B(n5327), .Z(n5329) );
  XNOR U5461 ( .A(n5330), .B(n5329), .Z(n5334) );
  NANDN U5462 ( .A(n5281), .B(n5280), .Z(n5285) );
  NAND U5463 ( .A(n5283), .B(n5282), .Z(n5284) );
  AND U5464 ( .A(n5285), .B(n5284), .Z(n5333) );
  XOR U5465 ( .A(n5334), .B(n5333), .Z(n5335) );
  NANDN U5466 ( .A(n5287), .B(n5286), .Z(n5291) );
  NANDN U5467 ( .A(n5289), .B(n5288), .Z(n5290) );
  NAND U5468 ( .A(n5291), .B(n5290), .Z(n5336) );
  XOR U5469 ( .A(n5335), .B(n5336), .Z(n5303) );
  OR U5470 ( .A(n5293), .B(n5292), .Z(n5297) );
  NANDN U5471 ( .A(n5295), .B(n5294), .Z(n5296) );
  NAND U5472 ( .A(n5297), .B(n5296), .Z(n5304) );
  XNOR U5473 ( .A(n5303), .B(n5304), .Z(n5305) );
  XNOR U5474 ( .A(n5306), .B(n5305), .Z(n5339) );
  XNOR U5475 ( .A(n5339), .B(sreg[1143]), .Z(n5341) );
  NAND U5476 ( .A(n5298), .B(sreg[1142]), .Z(n5302) );
  OR U5477 ( .A(n5300), .B(n5299), .Z(n5301) );
  AND U5478 ( .A(n5302), .B(n5301), .Z(n5340) );
  XOR U5479 ( .A(n5341), .B(n5340), .Z(c[1143]) );
  NANDN U5480 ( .A(n5304), .B(n5303), .Z(n5308) );
  NAND U5481 ( .A(n5306), .B(n5305), .Z(n5307) );
  NAND U5482 ( .A(n5308), .B(n5307), .Z(n5347) );
  NAND U5483 ( .A(b[0]), .B(a[128]), .Z(n5309) );
  XNOR U5484 ( .A(b[1]), .B(n5309), .Z(n5311) );
  NAND U5485 ( .A(n33), .B(a[127]), .Z(n5310) );
  AND U5486 ( .A(n5311), .B(n5310), .Z(n5364) );
  XOR U5487 ( .A(a[124]), .B(n42197), .Z(n5353) );
  NANDN U5488 ( .A(n5353), .B(n42173), .Z(n5314) );
  NANDN U5489 ( .A(n5312), .B(n42172), .Z(n5313) );
  NAND U5490 ( .A(n5314), .B(n5313), .Z(n5362) );
  NAND U5491 ( .A(b[7]), .B(a[120]), .Z(n5363) );
  XNOR U5492 ( .A(n5362), .B(n5363), .Z(n5365) );
  XOR U5493 ( .A(n5364), .B(n5365), .Z(n5371) );
  NANDN U5494 ( .A(n5315), .B(n42093), .Z(n5317) );
  XOR U5495 ( .A(n42134), .B(a[126]), .Z(n5356) );
  NANDN U5496 ( .A(n5356), .B(n42095), .Z(n5316) );
  NAND U5497 ( .A(n5317), .B(n5316), .Z(n5369) );
  NANDN U5498 ( .A(n5318), .B(n42231), .Z(n5320) );
  XOR U5499 ( .A(n172), .B(a[122]), .Z(n5359) );
  NANDN U5500 ( .A(n5359), .B(n42234), .Z(n5319) );
  AND U5501 ( .A(n5320), .B(n5319), .Z(n5368) );
  XNOR U5502 ( .A(n5369), .B(n5368), .Z(n5370) );
  XNOR U5503 ( .A(n5371), .B(n5370), .Z(n5375) );
  NANDN U5504 ( .A(n5322), .B(n5321), .Z(n5326) );
  NAND U5505 ( .A(n5324), .B(n5323), .Z(n5325) );
  AND U5506 ( .A(n5326), .B(n5325), .Z(n5374) );
  XOR U5507 ( .A(n5375), .B(n5374), .Z(n5376) );
  NANDN U5508 ( .A(n5328), .B(n5327), .Z(n5332) );
  NANDN U5509 ( .A(n5330), .B(n5329), .Z(n5331) );
  NAND U5510 ( .A(n5332), .B(n5331), .Z(n5377) );
  XOR U5511 ( .A(n5376), .B(n5377), .Z(n5344) );
  OR U5512 ( .A(n5334), .B(n5333), .Z(n5338) );
  NANDN U5513 ( .A(n5336), .B(n5335), .Z(n5337) );
  NAND U5514 ( .A(n5338), .B(n5337), .Z(n5345) );
  XNOR U5515 ( .A(n5344), .B(n5345), .Z(n5346) );
  XNOR U5516 ( .A(n5347), .B(n5346), .Z(n5380) );
  XNOR U5517 ( .A(n5380), .B(sreg[1144]), .Z(n5382) );
  NAND U5518 ( .A(n5339), .B(sreg[1143]), .Z(n5343) );
  OR U5519 ( .A(n5341), .B(n5340), .Z(n5342) );
  AND U5520 ( .A(n5343), .B(n5342), .Z(n5381) );
  XOR U5521 ( .A(n5382), .B(n5381), .Z(c[1144]) );
  NANDN U5522 ( .A(n5345), .B(n5344), .Z(n5349) );
  NAND U5523 ( .A(n5347), .B(n5346), .Z(n5348) );
  NAND U5524 ( .A(n5349), .B(n5348), .Z(n5388) );
  NAND U5525 ( .A(b[0]), .B(a[129]), .Z(n5350) );
  XNOR U5526 ( .A(b[1]), .B(n5350), .Z(n5352) );
  NAND U5527 ( .A(n33), .B(a[128]), .Z(n5351) );
  AND U5528 ( .A(n5352), .B(n5351), .Z(n5405) );
  XOR U5529 ( .A(a[125]), .B(n42197), .Z(n5394) );
  NANDN U5530 ( .A(n5394), .B(n42173), .Z(n5355) );
  NANDN U5531 ( .A(n5353), .B(n42172), .Z(n5354) );
  NAND U5532 ( .A(n5355), .B(n5354), .Z(n5403) );
  NAND U5533 ( .A(b[7]), .B(a[121]), .Z(n5404) );
  XNOR U5534 ( .A(n5403), .B(n5404), .Z(n5406) );
  XOR U5535 ( .A(n5405), .B(n5406), .Z(n5412) );
  NANDN U5536 ( .A(n5356), .B(n42093), .Z(n5358) );
  XOR U5537 ( .A(n42134), .B(a[127]), .Z(n5397) );
  NANDN U5538 ( .A(n5397), .B(n42095), .Z(n5357) );
  NAND U5539 ( .A(n5358), .B(n5357), .Z(n5410) );
  NANDN U5540 ( .A(n5359), .B(n42231), .Z(n5361) );
  XOR U5541 ( .A(n172), .B(a[123]), .Z(n5400) );
  NANDN U5542 ( .A(n5400), .B(n42234), .Z(n5360) );
  AND U5543 ( .A(n5361), .B(n5360), .Z(n5409) );
  XNOR U5544 ( .A(n5410), .B(n5409), .Z(n5411) );
  XNOR U5545 ( .A(n5412), .B(n5411), .Z(n5416) );
  NANDN U5546 ( .A(n5363), .B(n5362), .Z(n5367) );
  NAND U5547 ( .A(n5365), .B(n5364), .Z(n5366) );
  AND U5548 ( .A(n5367), .B(n5366), .Z(n5415) );
  XOR U5549 ( .A(n5416), .B(n5415), .Z(n5417) );
  NANDN U5550 ( .A(n5369), .B(n5368), .Z(n5373) );
  NANDN U5551 ( .A(n5371), .B(n5370), .Z(n5372) );
  NAND U5552 ( .A(n5373), .B(n5372), .Z(n5418) );
  XOR U5553 ( .A(n5417), .B(n5418), .Z(n5385) );
  OR U5554 ( .A(n5375), .B(n5374), .Z(n5379) );
  NANDN U5555 ( .A(n5377), .B(n5376), .Z(n5378) );
  NAND U5556 ( .A(n5379), .B(n5378), .Z(n5386) );
  XNOR U5557 ( .A(n5385), .B(n5386), .Z(n5387) );
  XNOR U5558 ( .A(n5388), .B(n5387), .Z(n5421) );
  XNOR U5559 ( .A(n5421), .B(sreg[1145]), .Z(n5423) );
  NAND U5560 ( .A(n5380), .B(sreg[1144]), .Z(n5384) );
  OR U5561 ( .A(n5382), .B(n5381), .Z(n5383) );
  AND U5562 ( .A(n5384), .B(n5383), .Z(n5422) );
  XOR U5563 ( .A(n5423), .B(n5422), .Z(c[1145]) );
  NANDN U5564 ( .A(n5386), .B(n5385), .Z(n5390) );
  NAND U5565 ( .A(n5388), .B(n5387), .Z(n5389) );
  NAND U5566 ( .A(n5390), .B(n5389), .Z(n5429) );
  NAND U5567 ( .A(b[0]), .B(a[130]), .Z(n5391) );
  XNOR U5568 ( .A(b[1]), .B(n5391), .Z(n5393) );
  NAND U5569 ( .A(n33), .B(a[129]), .Z(n5392) );
  AND U5570 ( .A(n5393), .B(n5392), .Z(n5446) );
  XOR U5571 ( .A(a[126]), .B(n42197), .Z(n5435) );
  NANDN U5572 ( .A(n5435), .B(n42173), .Z(n5396) );
  NANDN U5573 ( .A(n5394), .B(n42172), .Z(n5395) );
  NAND U5574 ( .A(n5396), .B(n5395), .Z(n5444) );
  NAND U5575 ( .A(b[7]), .B(a[122]), .Z(n5445) );
  XNOR U5576 ( .A(n5444), .B(n5445), .Z(n5447) );
  XOR U5577 ( .A(n5446), .B(n5447), .Z(n5453) );
  NANDN U5578 ( .A(n5397), .B(n42093), .Z(n5399) );
  XOR U5579 ( .A(n42134), .B(a[128]), .Z(n5438) );
  NANDN U5580 ( .A(n5438), .B(n42095), .Z(n5398) );
  NAND U5581 ( .A(n5399), .B(n5398), .Z(n5451) );
  NANDN U5582 ( .A(n5400), .B(n42231), .Z(n5402) );
  XOR U5583 ( .A(n172), .B(a[124]), .Z(n5441) );
  NANDN U5584 ( .A(n5441), .B(n42234), .Z(n5401) );
  AND U5585 ( .A(n5402), .B(n5401), .Z(n5450) );
  XNOR U5586 ( .A(n5451), .B(n5450), .Z(n5452) );
  XNOR U5587 ( .A(n5453), .B(n5452), .Z(n5457) );
  NANDN U5588 ( .A(n5404), .B(n5403), .Z(n5408) );
  NAND U5589 ( .A(n5406), .B(n5405), .Z(n5407) );
  AND U5590 ( .A(n5408), .B(n5407), .Z(n5456) );
  XOR U5591 ( .A(n5457), .B(n5456), .Z(n5458) );
  NANDN U5592 ( .A(n5410), .B(n5409), .Z(n5414) );
  NANDN U5593 ( .A(n5412), .B(n5411), .Z(n5413) );
  NAND U5594 ( .A(n5414), .B(n5413), .Z(n5459) );
  XOR U5595 ( .A(n5458), .B(n5459), .Z(n5426) );
  OR U5596 ( .A(n5416), .B(n5415), .Z(n5420) );
  NANDN U5597 ( .A(n5418), .B(n5417), .Z(n5419) );
  NAND U5598 ( .A(n5420), .B(n5419), .Z(n5427) );
  XNOR U5599 ( .A(n5426), .B(n5427), .Z(n5428) );
  XNOR U5600 ( .A(n5429), .B(n5428), .Z(n5462) );
  XNOR U5601 ( .A(n5462), .B(sreg[1146]), .Z(n5464) );
  NAND U5602 ( .A(n5421), .B(sreg[1145]), .Z(n5425) );
  OR U5603 ( .A(n5423), .B(n5422), .Z(n5424) );
  AND U5604 ( .A(n5425), .B(n5424), .Z(n5463) );
  XOR U5605 ( .A(n5464), .B(n5463), .Z(c[1146]) );
  NANDN U5606 ( .A(n5427), .B(n5426), .Z(n5431) );
  NAND U5607 ( .A(n5429), .B(n5428), .Z(n5430) );
  NAND U5608 ( .A(n5431), .B(n5430), .Z(n5470) );
  NAND U5609 ( .A(b[0]), .B(a[131]), .Z(n5432) );
  XNOR U5610 ( .A(b[1]), .B(n5432), .Z(n5434) );
  NAND U5611 ( .A(n33), .B(a[130]), .Z(n5433) );
  AND U5612 ( .A(n5434), .B(n5433), .Z(n5487) );
  XOR U5613 ( .A(a[127]), .B(n42197), .Z(n5476) );
  NANDN U5614 ( .A(n5476), .B(n42173), .Z(n5437) );
  NANDN U5615 ( .A(n5435), .B(n42172), .Z(n5436) );
  NAND U5616 ( .A(n5437), .B(n5436), .Z(n5485) );
  NAND U5617 ( .A(b[7]), .B(a[123]), .Z(n5486) );
  XNOR U5618 ( .A(n5485), .B(n5486), .Z(n5488) );
  XOR U5619 ( .A(n5487), .B(n5488), .Z(n5494) );
  NANDN U5620 ( .A(n5438), .B(n42093), .Z(n5440) );
  XOR U5621 ( .A(n42134), .B(a[129]), .Z(n5479) );
  NANDN U5622 ( .A(n5479), .B(n42095), .Z(n5439) );
  NAND U5623 ( .A(n5440), .B(n5439), .Z(n5492) );
  NANDN U5624 ( .A(n5441), .B(n42231), .Z(n5443) );
  XOR U5625 ( .A(n172), .B(a[125]), .Z(n5482) );
  NANDN U5626 ( .A(n5482), .B(n42234), .Z(n5442) );
  AND U5627 ( .A(n5443), .B(n5442), .Z(n5491) );
  XNOR U5628 ( .A(n5492), .B(n5491), .Z(n5493) );
  XNOR U5629 ( .A(n5494), .B(n5493), .Z(n5498) );
  NANDN U5630 ( .A(n5445), .B(n5444), .Z(n5449) );
  NAND U5631 ( .A(n5447), .B(n5446), .Z(n5448) );
  AND U5632 ( .A(n5449), .B(n5448), .Z(n5497) );
  XOR U5633 ( .A(n5498), .B(n5497), .Z(n5499) );
  NANDN U5634 ( .A(n5451), .B(n5450), .Z(n5455) );
  NANDN U5635 ( .A(n5453), .B(n5452), .Z(n5454) );
  NAND U5636 ( .A(n5455), .B(n5454), .Z(n5500) );
  XOR U5637 ( .A(n5499), .B(n5500), .Z(n5467) );
  OR U5638 ( .A(n5457), .B(n5456), .Z(n5461) );
  NANDN U5639 ( .A(n5459), .B(n5458), .Z(n5460) );
  NAND U5640 ( .A(n5461), .B(n5460), .Z(n5468) );
  XNOR U5641 ( .A(n5467), .B(n5468), .Z(n5469) );
  XNOR U5642 ( .A(n5470), .B(n5469), .Z(n5503) );
  XNOR U5643 ( .A(n5503), .B(sreg[1147]), .Z(n5505) );
  NAND U5644 ( .A(n5462), .B(sreg[1146]), .Z(n5466) );
  OR U5645 ( .A(n5464), .B(n5463), .Z(n5465) );
  AND U5646 ( .A(n5466), .B(n5465), .Z(n5504) );
  XOR U5647 ( .A(n5505), .B(n5504), .Z(c[1147]) );
  NANDN U5648 ( .A(n5468), .B(n5467), .Z(n5472) );
  NAND U5649 ( .A(n5470), .B(n5469), .Z(n5471) );
  NAND U5650 ( .A(n5472), .B(n5471), .Z(n5511) );
  NAND U5651 ( .A(b[0]), .B(a[132]), .Z(n5473) );
  XNOR U5652 ( .A(b[1]), .B(n5473), .Z(n5475) );
  NAND U5653 ( .A(n33), .B(a[131]), .Z(n5474) );
  AND U5654 ( .A(n5475), .B(n5474), .Z(n5528) );
  XOR U5655 ( .A(a[128]), .B(n42197), .Z(n5517) );
  NANDN U5656 ( .A(n5517), .B(n42173), .Z(n5478) );
  NANDN U5657 ( .A(n5476), .B(n42172), .Z(n5477) );
  NAND U5658 ( .A(n5478), .B(n5477), .Z(n5526) );
  NAND U5659 ( .A(b[7]), .B(a[124]), .Z(n5527) );
  XNOR U5660 ( .A(n5526), .B(n5527), .Z(n5529) );
  XOR U5661 ( .A(n5528), .B(n5529), .Z(n5535) );
  NANDN U5662 ( .A(n5479), .B(n42093), .Z(n5481) );
  XOR U5663 ( .A(n42134), .B(a[130]), .Z(n5520) );
  NANDN U5664 ( .A(n5520), .B(n42095), .Z(n5480) );
  NAND U5665 ( .A(n5481), .B(n5480), .Z(n5533) );
  NANDN U5666 ( .A(n5482), .B(n42231), .Z(n5484) );
  XOR U5667 ( .A(n172), .B(a[126]), .Z(n5523) );
  NANDN U5668 ( .A(n5523), .B(n42234), .Z(n5483) );
  AND U5669 ( .A(n5484), .B(n5483), .Z(n5532) );
  XNOR U5670 ( .A(n5533), .B(n5532), .Z(n5534) );
  XNOR U5671 ( .A(n5535), .B(n5534), .Z(n5539) );
  NANDN U5672 ( .A(n5486), .B(n5485), .Z(n5490) );
  NAND U5673 ( .A(n5488), .B(n5487), .Z(n5489) );
  AND U5674 ( .A(n5490), .B(n5489), .Z(n5538) );
  XOR U5675 ( .A(n5539), .B(n5538), .Z(n5540) );
  NANDN U5676 ( .A(n5492), .B(n5491), .Z(n5496) );
  NANDN U5677 ( .A(n5494), .B(n5493), .Z(n5495) );
  NAND U5678 ( .A(n5496), .B(n5495), .Z(n5541) );
  XOR U5679 ( .A(n5540), .B(n5541), .Z(n5508) );
  OR U5680 ( .A(n5498), .B(n5497), .Z(n5502) );
  NANDN U5681 ( .A(n5500), .B(n5499), .Z(n5501) );
  NAND U5682 ( .A(n5502), .B(n5501), .Z(n5509) );
  XNOR U5683 ( .A(n5508), .B(n5509), .Z(n5510) );
  XNOR U5684 ( .A(n5511), .B(n5510), .Z(n5544) );
  XNOR U5685 ( .A(n5544), .B(sreg[1148]), .Z(n5546) );
  NAND U5686 ( .A(n5503), .B(sreg[1147]), .Z(n5507) );
  OR U5687 ( .A(n5505), .B(n5504), .Z(n5506) );
  AND U5688 ( .A(n5507), .B(n5506), .Z(n5545) );
  XOR U5689 ( .A(n5546), .B(n5545), .Z(c[1148]) );
  NANDN U5690 ( .A(n5509), .B(n5508), .Z(n5513) );
  NAND U5691 ( .A(n5511), .B(n5510), .Z(n5512) );
  NAND U5692 ( .A(n5513), .B(n5512), .Z(n5552) );
  NAND U5693 ( .A(b[0]), .B(a[133]), .Z(n5514) );
  XNOR U5694 ( .A(b[1]), .B(n5514), .Z(n5516) );
  NAND U5695 ( .A(n34), .B(a[132]), .Z(n5515) );
  AND U5696 ( .A(n5516), .B(n5515), .Z(n5569) );
  XOR U5697 ( .A(a[129]), .B(n42197), .Z(n5558) );
  NANDN U5698 ( .A(n5558), .B(n42173), .Z(n5519) );
  NANDN U5699 ( .A(n5517), .B(n42172), .Z(n5518) );
  NAND U5700 ( .A(n5519), .B(n5518), .Z(n5567) );
  NAND U5701 ( .A(b[7]), .B(a[125]), .Z(n5568) );
  XNOR U5702 ( .A(n5567), .B(n5568), .Z(n5570) );
  XOR U5703 ( .A(n5569), .B(n5570), .Z(n5576) );
  NANDN U5704 ( .A(n5520), .B(n42093), .Z(n5522) );
  XOR U5705 ( .A(n42134), .B(a[131]), .Z(n5561) );
  NANDN U5706 ( .A(n5561), .B(n42095), .Z(n5521) );
  NAND U5707 ( .A(n5522), .B(n5521), .Z(n5574) );
  NANDN U5708 ( .A(n5523), .B(n42231), .Z(n5525) );
  XOR U5709 ( .A(n172), .B(a[127]), .Z(n5564) );
  NANDN U5710 ( .A(n5564), .B(n42234), .Z(n5524) );
  AND U5711 ( .A(n5525), .B(n5524), .Z(n5573) );
  XNOR U5712 ( .A(n5574), .B(n5573), .Z(n5575) );
  XNOR U5713 ( .A(n5576), .B(n5575), .Z(n5580) );
  NANDN U5714 ( .A(n5527), .B(n5526), .Z(n5531) );
  NAND U5715 ( .A(n5529), .B(n5528), .Z(n5530) );
  AND U5716 ( .A(n5531), .B(n5530), .Z(n5579) );
  XOR U5717 ( .A(n5580), .B(n5579), .Z(n5581) );
  NANDN U5718 ( .A(n5533), .B(n5532), .Z(n5537) );
  NANDN U5719 ( .A(n5535), .B(n5534), .Z(n5536) );
  NAND U5720 ( .A(n5537), .B(n5536), .Z(n5582) );
  XOR U5721 ( .A(n5581), .B(n5582), .Z(n5549) );
  OR U5722 ( .A(n5539), .B(n5538), .Z(n5543) );
  NANDN U5723 ( .A(n5541), .B(n5540), .Z(n5542) );
  NAND U5724 ( .A(n5543), .B(n5542), .Z(n5550) );
  XNOR U5725 ( .A(n5549), .B(n5550), .Z(n5551) );
  XNOR U5726 ( .A(n5552), .B(n5551), .Z(n5585) );
  XNOR U5727 ( .A(n5585), .B(sreg[1149]), .Z(n5587) );
  NAND U5728 ( .A(n5544), .B(sreg[1148]), .Z(n5548) );
  OR U5729 ( .A(n5546), .B(n5545), .Z(n5547) );
  AND U5730 ( .A(n5548), .B(n5547), .Z(n5586) );
  XOR U5731 ( .A(n5587), .B(n5586), .Z(c[1149]) );
  NANDN U5732 ( .A(n5550), .B(n5549), .Z(n5554) );
  NAND U5733 ( .A(n5552), .B(n5551), .Z(n5553) );
  NAND U5734 ( .A(n5554), .B(n5553), .Z(n5593) );
  NAND U5735 ( .A(b[0]), .B(a[134]), .Z(n5555) );
  XNOR U5736 ( .A(b[1]), .B(n5555), .Z(n5557) );
  NAND U5737 ( .A(n34), .B(a[133]), .Z(n5556) );
  AND U5738 ( .A(n5557), .B(n5556), .Z(n5610) );
  XOR U5739 ( .A(a[130]), .B(n42197), .Z(n5599) );
  NANDN U5740 ( .A(n5599), .B(n42173), .Z(n5560) );
  NANDN U5741 ( .A(n5558), .B(n42172), .Z(n5559) );
  NAND U5742 ( .A(n5560), .B(n5559), .Z(n5608) );
  NAND U5743 ( .A(b[7]), .B(a[126]), .Z(n5609) );
  XNOR U5744 ( .A(n5608), .B(n5609), .Z(n5611) );
  XOR U5745 ( .A(n5610), .B(n5611), .Z(n5617) );
  NANDN U5746 ( .A(n5561), .B(n42093), .Z(n5563) );
  XOR U5747 ( .A(n42134), .B(a[132]), .Z(n5602) );
  NANDN U5748 ( .A(n5602), .B(n42095), .Z(n5562) );
  NAND U5749 ( .A(n5563), .B(n5562), .Z(n5615) );
  NANDN U5750 ( .A(n5564), .B(n42231), .Z(n5566) );
  XOR U5751 ( .A(n172), .B(a[128]), .Z(n5605) );
  NANDN U5752 ( .A(n5605), .B(n42234), .Z(n5565) );
  AND U5753 ( .A(n5566), .B(n5565), .Z(n5614) );
  XNOR U5754 ( .A(n5615), .B(n5614), .Z(n5616) );
  XNOR U5755 ( .A(n5617), .B(n5616), .Z(n5621) );
  NANDN U5756 ( .A(n5568), .B(n5567), .Z(n5572) );
  NAND U5757 ( .A(n5570), .B(n5569), .Z(n5571) );
  AND U5758 ( .A(n5572), .B(n5571), .Z(n5620) );
  XOR U5759 ( .A(n5621), .B(n5620), .Z(n5622) );
  NANDN U5760 ( .A(n5574), .B(n5573), .Z(n5578) );
  NANDN U5761 ( .A(n5576), .B(n5575), .Z(n5577) );
  NAND U5762 ( .A(n5578), .B(n5577), .Z(n5623) );
  XOR U5763 ( .A(n5622), .B(n5623), .Z(n5590) );
  OR U5764 ( .A(n5580), .B(n5579), .Z(n5584) );
  NANDN U5765 ( .A(n5582), .B(n5581), .Z(n5583) );
  NAND U5766 ( .A(n5584), .B(n5583), .Z(n5591) );
  XNOR U5767 ( .A(n5590), .B(n5591), .Z(n5592) );
  XNOR U5768 ( .A(n5593), .B(n5592), .Z(n5626) );
  XNOR U5769 ( .A(n5626), .B(sreg[1150]), .Z(n5628) );
  NAND U5770 ( .A(n5585), .B(sreg[1149]), .Z(n5589) );
  OR U5771 ( .A(n5587), .B(n5586), .Z(n5588) );
  AND U5772 ( .A(n5589), .B(n5588), .Z(n5627) );
  XOR U5773 ( .A(n5628), .B(n5627), .Z(c[1150]) );
  NANDN U5774 ( .A(n5591), .B(n5590), .Z(n5595) );
  NAND U5775 ( .A(n5593), .B(n5592), .Z(n5594) );
  NAND U5776 ( .A(n5595), .B(n5594), .Z(n5634) );
  NAND U5777 ( .A(b[0]), .B(a[135]), .Z(n5596) );
  XNOR U5778 ( .A(b[1]), .B(n5596), .Z(n5598) );
  NAND U5779 ( .A(n34), .B(a[134]), .Z(n5597) );
  AND U5780 ( .A(n5598), .B(n5597), .Z(n5651) );
  XOR U5781 ( .A(a[131]), .B(n42197), .Z(n5640) );
  NANDN U5782 ( .A(n5640), .B(n42173), .Z(n5601) );
  NANDN U5783 ( .A(n5599), .B(n42172), .Z(n5600) );
  NAND U5784 ( .A(n5601), .B(n5600), .Z(n5649) );
  NAND U5785 ( .A(b[7]), .B(a[127]), .Z(n5650) );
  XNOR U5786 ( .A(n5649), .B(n5650), .Z(n5652) );
  XOR U5787 ( .A(n5651), .B(n5652), .Z(n5658) );
  NANDN U5788 ( .A(n5602), .B(n42093), .Z(n5604) );
  XOR U5789 ( .A(n42134), .B(a[133]), .Z(n5643) );
  NANDN U5790 ( .A(n5643), .B(n42095), .Z(n5603) );
  NAND U5791 ( .A(n5604), .B(n5603), .Z(n5656) );
  NANDN U5792 ( .A(n5605), .B(n42231), .Z(n5607) );
  XOR U5793 ( .A(n172), .B(a[129]), .Z(n5646) );
  NANDN U5794 ( .A(n5646), .B(n42234), .Z(n5606) );
  AND U5795 ( .A(n5607), .B(n5606), .Z(n5655) );
  XNOR U5796 ( .A(n5656), .B(n5655), .Z(n5657) );
  XNOR U5797 ( .A(n5658), .B(n5657), .Z(n5662) );
  NANDN U5798 ( .A(n5609), .B(n5608), .Z(n5613) );
  NAND U5799 ( .A(n5611), .B(n5610), .Z(n5612) );
  AND U5800 ( .A(n5613), .B(n5612), .Z(n5661) );
  XOR U5801 ( .A(n5662), .B(n5661), .Z(n5663) );
  NANDN U5802 ( .A(n5615), .B(n5614), .Z(n5619) );
  NANDN U5803 ( .A(n5617), .B(n5616), .Z(n5618) );
  NAND U5804 ( .A(n5619), .B(n5618), .Z(n5664) );
  XOR U5805 ( .A(n5663), .B(n5664), .Z(n5631) );
  OR U5806 ( .A(n5621), .B(n5620), .Z(n5625) );
  NANDN U5807 ( .A(n5623), .B(n5622), .Z(n5624) );
  NAND U5808 ( .A(n5625), .B(n5624), .Z(n5632) );
  XNOR U5809 ( .A(n5631), .B(n5632), .Z(n5633) );
  XNOR U5810 ( .A(n5634), .B(n5633), .Z(n5667) );
  XNOR U5811 ( .A(n5667), .B(sreg[1151]), .Z(n5669) );
  NAND U5812 ( .A(n5626), .B(sreg[1150]), .Z(n5630) );
  OR U5813 ( .A(n5628), .B(n5627), .Z(n5629) );
  AND U5814 ( .A(n5630), .B(n5629), .Z(n5668) );
  XOR U5815 ( .A(n5669), .B(n5668), .Z(c[1151]) );
  NANDN U5816 ( .A(n5632), .B(n5631), .Z(n5636) );
  NAND U5817 ( .A(n5634), .B(n5633), .Z(n5635) );
  NAND U5818 ( .A(n5636), .B(n5635), .Z(n5675) );
  NAND U5819 ( .A(b[0]), .B(a[136]), .Z(n5637) );
  XNOR U5820 ( .A(b[1]), .B(n5637), .Z(n5639) );
  NAND U5821 ( .A(n34), .B(a[135]), .Z(n5638) );
  AND U5822 ( .A(n5639), .B(n5638), .Z(n5692) );
  XOR U5823 ( .A(a[132]), .B(n42197), .Z(n5681) );
  NANDN U5824 ( .A(n5681), .B(n42173), .Z(n5642) );
  NANDN U5825 ( .A(n5640), .B(n42172), .Z(n5641) );
  NAND U5826 ( .A(n5642), .B(n5641), .Z(n5690) );
  NAND U5827 ( .A(b[7]), .B(a[128]), .Z(n5691) );
  XNOR U5828 ( .A(n5690), .B(n5691), .Z(n5693) );
  XOR U5829 ( .A(n5692), .B(n5693), .Z(n5699) );
  NANDN U5830 ( .A(n5643), .B(n42093), .Z(n5645) );
  XOR U5831 ( .A(n42134), .B(a[134]), .Z(n5684) );
  NANDN U5832 ( .A(n5684), .B(n42095), .Z(n5644) );
  NAND U5833 ( .A(n5645), .B(n5644), .Z(n5697) );
  NANDN U5834 ( .A(n5646), .B(n42231), .Z(n5648) );
  XOR U5835 ( .A(n172), .B(a[130]), .Z(n5687) );
  NANDN U5836 ( .A(n5687), .B(n42234), .Z(n5647) );
  AND U5837 ( .A(n5648), .B(n5647), .Z(n5696) );
  XNOR U5838 ( .A(n5697), .B(n5696), .Z(n5698) );
  XNOR U5839 ( .A(n5699), .B(n5698), .Z(n5703) );
  NANDN U5840 ( .A(n5650), .B(n5649), .Z(n5654) );
  NAND U5841 ( .A(n5652), .B(n5651), .Z(n5653) );
  AND U5842 ( .A(n5654), .B(n5653), .Z(n5702) );
  XOR U5843 ( .A(n5703), .B(n5702), .Z(n5704) );
  NANDN U5844 ( .A(n5656), .B(n5655), .Z(n5660) );
  NANDN U5845 ( .A(n5658), .B(n5657), .Z(n5659) );
  NAND U5846 ( .A(n5660), .B(n5659), .Z(n5705) );
  XOR U5847 ( .A(n5704), .B(n5705), .Z(n5672) );
  OR U5848 ( .A(n5662), .B(n5661), .Z(n5666) );
  NANDN U5849 ( .A(n5664), .B(n5663), .Z(n5665) );
  NAND U5850 ( .A(n5666), .B(n5665), .Z(n5673) );
  XNOR U5851 ( .A(n5672), .B(n5673), .Z(n5674) );
  XNOR U5852 ( .A(n5675), .B(n5674), .Z(n5708) );
  XNOR U5853 ( .A(n5708), .B(sreg[1152]), .Z(n5710) );
  NAND U5854 ( .A(n5667), .B(sreg[1151]), .Z(n5671) );
  OR U5855 ( .A(n5669), .B(n5668), .Z(n5670) );
  AND U5856 ( .A(n5671), .B(n5670), .Z(n5709) );
  XOR U5857 ( .A(n5710), .B(n5709), .Z(c[1152]) );
  NANDN U5858 ( .A(n5673), .B(n5672), .Z(n5677) );
  NAND U5859 ( .A(n5675), .B(n5674), .Z(n5676) );
  NAND U5860 ( .A(n5677), .B(n5676), .Z(n5716) );
  NAND U5861 ( .A(b[0]), .B(a[137]), .Z(n5678) );
  XNOR U5862 ( .A(b[1]), .B(n5678), .Z(n5680) );
  NAND U5863 ( .A(n34), .B(a[136]), .Z(n5679) );
  AND U5864 ( .A(n5680), .B(n5679), .Z(n5733) );
  XOR U5865 ( .A(a[133]), .B(n42197), .Z(n5722) );
  NANDN U5866 ( .A(n5722), .B(n42173), .Z(n5683) );
  NANDN U5867 ( .A(n5681), .B(n42172), .Z(n5682) );
  NAND U5868 ( .A(n5683), .B(n5682), .Z(n5731) );
  NAND U5869 ( .A(b[7]), .B(a[129]), .Z(n5732) );
  XNOR U5870 ( .A(n5731), .B(n5732), .Z(n5734) );
  XOR U5871 ( .A(n5733), .B(n5734), .Z(n5740) );
  NANDN U5872 ( .A(n5684), .B(n42093), .Z(n5686) );
  XOR U5873 ( .A(n42134), .B(a[135]), .Z(n5725) );
  NANDN U5874 ( .A(n5725), .B(n42095), .Z(n5685) );
  NAND U5875 ( .A(n5686), .B(n5685), .Z(n5738) );
  NANDN U5876 ( .A(n5687), .B(n42231), .Z(n5689) );
  XOR U5877 ( .A(n173), .B(a[131]), .Z(n5728) );
  NANDN U5878 ( .A(n5728), .B(n42234), .Z(n5688) );
  AND U5879 ( .A(n5689), .B(n5688), .Z(n5737) );
  XNOR U5880 ( .A(n5738), .B(n5737), .Z(n5739) );
  XNOR U5881 ( .A(n5740), .B(n5739), .Z(n5744) );
  NANDN U5882 ( .A(n5691), .B(n5690), .Z(n5695) );
  NAND U5883 ( .A(n5693), .B(n5692), .Z(n5694) );
  AND U5884 ( .A(n5695), .B(n5694), .Z(n5743) );
  XOR U5885 ( .A(n5744), .B(n5743), .Z(n5745) );
  NANDN U5886 ( .A(n5697), .B(n5696), .Z(n5701) );
  NANDN U5887 ( .A(n5699), .B(n5698), .Z(n5700) );
  NAND U5888 ( .A(n5701), .B(n5700), .Z(n5746) );
  XOR U5889 ( .A(n5745), .B(n5746), .Z(n5713) );
  OR U5890 ( .A(n5703), .B(n5702), .Z(n5707) );
  NANDN U5891 ( .A(n5705), .B(n5704), .Z(n5706) );
  NAND U5892 ( .A(n5707), .B(n5706), .Z(n5714) );
  XNOR U5893 ( .A(n5713), .B(n5714), .Z(n5715) );
  XNOR U5894 ( .A(n5716), .B(n5715), .Z(n5749) );
  XNOR U5895 ( .A(n5749), .B(sreg[1153]), .Z(n5751) );
  NAND U5896 ( .A(n5708), .B(sreg[1152]), .Z(n5712) );
  OR U5897 ( .A(n5710), .B(n5709), .Z(n5711) );
  AND U5898 ( .A(n5712), .B(n5711), .Z(n5750) );
  XOR U5899 ( .A(n5751), .B(n5750), .Z(c[1153]) );
  NANDN U5900 ( .A(n5714), .B(n5713), .Z(n5718) );
  NAND U5901 ( .A(n5716), .B(n5715), .Z(n5717) );
  NAND U5902 ( .A(n5718), .B(n5717), .Z(n5757) );
  NAND U5903 ( .A(b[0]), .B(a[138]), .Z(n5719) );
  XNOR U5904 ( .A(b[1]), .B(n5719), .Z(n5721) );
  NAND U5905 ( .A(n34), .B(a[137]), .Z(n5720) );
  AND U5906 ( .A(n5721), .B(n5720), .Z(n5774) );
  XOR U5907 ( .A(a[134]), .B(n42197), .Z(n5763) );
  NANDN U5908 ( .A(n5763), .B(n42173), .Z(n5724) );
  NANDN U5909 ( .A(n5722), .B(n42172), .Z(n5723) );
  NAND U5910 ( .A(n5724), .B(n5723), .Z(n5772) );
  NAND U5911 ( .A(b[7]), .B(a[130]), .Z(n5773) );
  XNOR U5912 ( .A(n5772), .B(n5773), .Z(n5775) );
  XOR U5913 ( .A(n5774), .B(n5775), .Z(n5781) );
  NANDN U5914 ( .A(n5725), .B(n42093), .Z(n5727) );
  XOR U5915 ( .A(n42134), .B(a[136]), .Z(n5766) );
  NANDN U5916 ( .A(n5766), .B(n42095), .Z(n5726) );
  NAND U5917 ( .A(n5727), .B(n5726), .Z(n5779) );
  NANDN U5918 ( .A(n5728), .B(n42231), .Z(n5730) );
  XOR U5919 ( .A(n173), .B(a[132]), .Z(n5769) );
  NANDN U5920 ( .A(n5769), .B(n42234), .Z(n5729) );
  AND U5921 ( .A(n5730), .B(n5729), .Z(n5778) );
  XNOR U5922 ( .A(n5779), .B(n5778), .Z(n5780) );
  XNOR U5923 ( .A(n5781), .B(n5780), .Z(n5785) );
  NANDN U5924 ( .A(n5732), .B(n5731), .Z(n5736) );
  NAND U5925 ( .A(n5734), .B(n5733), .Z(n5735) );
  AND U5926 ( .A(n5736), .B(n5735), .Z(n5784) );
  XOR U5927 ( .A(n5785), .B(n5784), .Z(n5786) );
  NANDN U5928 ( .A(n5738), .B(n5737), .Z(n5742) );
  NANDN U5929 ( .A(n5740), .B(n5739), .Z(n5741) );
  NAND U5930 ( .A(n5742), .B(n5741), .Z(n5787) );
  XOR U5931 ( .A(n5786), .B(n5787), .Z(n5754) );
  OR U5932 ( .A(n5744), .B(n5743), .Z(n5748) );
  NANDN U5933 ( .A(n5746), .B(n5745), .Z(n5747) );
  NAND U5934 ( .A(n5748), .B(n5747), .Z(n5755) );
  XNOR U5935 ( .A(n5754), .B(n5755), .Z(n5756) );
  XNOR U5936 ( .A(n5757), .B(n5756), .Z(n5790) );
  XNOR U5937 ( .A(n5790), .B(sreg[1154]), .Z(n5792) );
  NAND U5938 ( .A(n5749), .B(sreg[1153]), .Z(n5753) );
  OR U5939 ( .A(n5751), .B(n5750), .Z(n5752) );
  AND U5940 ( .A(n5753), .B(n5752), .Z(n5791) );
  XOR U5941 ( .A(n5792), .B(n5791), .Z(c[1154]) );
  NANDN U5942 ( .A(n5755), .B(n5754), .Z(n5759) );
  NAND U5943 ( .A(n5757), .B(n5756), .Z(n5758) );
  NAND U5944 ( .A(n5759), .B(n5758), .Z(n5798) );
  NAND U5945 ( .A(b[0]), .B(a[139]), .Z(n5760) );
  XNOR U5946 ( .A(b[1]), .B(n5760), .Z(n5762) );
  NAND U5947 ( .A(n34), .B(a[138]), .Z(n5761) );
  AND U5948 ( .A(n5762), .B(n5761), .Z(n5815) );
  XOR U5949 ( .A(a[135]), .B(n42197), .Z(n5804) );
  NANDN U5950 ( .A(n5804), .B(n42173), .Z(n5765) );
  NANDN U5951 ( .A(n5763), .B(n42172), .Z(n5764) );
  NAND U5952 ( .A(n5765), .B(n5764), .Z(n5813) );
  NAND U5953 ( .A(b[7]), .B(a[131]), .Z(n5814) );
  XNOR U5954 ( .A(n5813), .B(n5814), .Z(n5816) );
  XOR U5955 ( .A(n5815), .B(n5816), .Z(n5822) );
  NANDN U5956 ( .A(n5766), .B(n42093), .Z(n5768) );
  XOR U5957 ( .A(n42134), .B(a[137]), .Z(n5807) );
  NANDN U5958 ( .A(n5807), .B(n42095), .Z(n5767) );
  NAND U5959 ( .A(n5768), .B(n5767), .Z(n5820) );
  NANDN U5960 ( .A(n5769), .B(n42231), .Z(n5771) );
  XOR U5961 ( .A(n173), .B(a[133]), .Z(n5810) );
  NANDN U5962 ( .A(n5810), .B(n42234), .Z(n5770) );
  AND U5963 ( .A(n5771), .B(n5770), .Z(n5819) );
  XNOR U5964 ( .A(n5820), .B(n5819), .Z(n5821) );
  XNOR U5965 ( .A(n5822), .B(n5821), .Z(n5826) );
  NANDN U5966 ( .A(n5773), .B(n5772), .Z(n5777) );
  NAND U5967 ( .A(n5775), .B(n5774), .Z(n5776) );
  AND U5968 ( .A(n5777), .B(n5776), .Z(n5825) );
  XOR U5969 ( .A(n5826), .B(n5825), .Z(n5827) );
  NANDN U5970 ( .A(n5779), .B(n5778), .Z(n5783) );
  NANDN U5971 ( .A(n5781), .B(n5780), .Z(n5782) );
  NAND U5972 ( .A(n5783), .B(n5782), .Z(n5828) );
  XOR U5973 ( .A(n5827), .B(n5828), .Z(n5795) );
  OR U5974 ( .A(n5785), .B(n5784), .Z(n5789) );
  NANDN U5975 ( .A(n5787), .B(n5786), .Z(n5788) );
  NAND U5976 ( .A(n5789), .B(n5788), .Z(n5796) );
  XNOR U5977 ( .A(n5795), .B(n5796), .Z(n5797) );
  XNOR U5978 ( .A(n5798), .B(n5797), .Z(n5831) );
  XNOR U5979 ( .A(n5831), .B(sreg[1155]), .Z(n5833) );
  NAND U5980 ( .A(n5790), .B(sreg[1154]), .Z(n5794) );
  OR U5981 ( .A(n5792), .B(n5791), .Z(n5793) );
  AND U5982 ( .A(n5794), .B(n5793), .Z(n5832) );
  XOR U5983 ( .A(n5833), .B(n5832), .Z(c[1155]) );
  NANDN U5984 ( .A(n5796), .B(n5795), .Z(n5800) );
  NAND U5985 ( .A(n5798), .B(n5797), .Z(n5799) );
  NAND U5986 ( .A(n5800), .B(n5799), .Z(n5839) );
  NAND U5987 ( .A(b[0]), .B(a[140]), .Z(n5801) );
  XNOR U5988 ( .A(b[1]), .B(n5801), .Z(n5803) );
  NAND U5989 ( .A(n35), .B(a[139]), .Z(n5802) );
  AND U5990 ( .A(n5803), .B(n5802), .Z(n5856) );
  XOR U5991 ( .A(a[136]), .B(n42197), .Z(n5845) );
  NANDN U5992 ( .A(n5845), .B(n42173), .Z(n5806) );
  NANDN U5993 ( .A(n5804), .B(n42172), .Z(n5805) );
  NAND U5994 ( .A(n5806), .B(n5805), .Z(n5854) );
  NAND U5995 ( .A(b[7]), .B(a[132]), .Z(n5855) );
  XNOR U5996 ( .A(n5854), .B(n5855), .Z(n5857) );
  XOR U5997 ( .A(n5856), .B(n5857), .Z(n5863) );
  NANDN U5998 ( .A(n5807), .B(n42093), .Z(n5809) );
  XOR U5999 ( .A(n42134), .B(a[138]), .Z(n5848) );
  NANDN U6000 ( .A(n5848), .B(n42095), .Z(n5808) );
  NAND U6001 ( .A(n5809), .B(n5808), .Z(n5861) );
  NANDN U6002 ( .A(n5810), .B(n42231), .Z(n5812) );
  XOR U6003 ( .A(n173), .B(a[134]), .Z(n5851) );
  NANDN U6004 ( .A(n5851), .B(n42234), .Z(n5811) );
  AND U6005 ( .A(n5812), .B(n5811), .Z(n5860) );
  XNOR U6006 ( .A(n5861), .B(n5860), .Z(n5862) );
  XNOR U6007 ( .A(n5863), .B(n5862), .Z(n5867) );
  NANDN U6008 ( .A(n5814), .B(n5813), .Z(n5818) );
  NAND U6009 ( .A(n5816), .B(n5815), .Z(n5817) );
  AND U6010 ( .A(n5818), .B(n5817), .Z(n5866) );
  XOR U6011 ( .A(n5867), .B(n5866), .Z(n5868) );
  NANDN U6012 ( .A(n5820), .B(n5819), .Z(n5824) );
  NANDN U6013 ( .A(n5822), .B(n5821), .Z(n5823) );
  NAND U6014 ( .A(n5824), .B(n5823), .Z(n5869) );
  XOR U6015 ( .A(n5868), .B(n5869), .Z(n5836) );
  OR U6016 ( .A(n5826), .B(n5825), .Z(n5830) );
  NANDN U6017 ( .A(n5828), .B(n5827), .Z(n5829) );
  NAND U6018 ( .A(n5830), .B(n5829), .Z(n5837) );
  XNOR U6019 ( .A(n5836), .B(n5837), .Z(n5838) );
  XNOR U6020 ( .A(n5839), .B(n5838), .Z(n5872) );
  XNOR U6021 ( .A(n5872), .B(sreg[1156]), .Z(n5874) );
  NAND U6022 ( .A(n5831), .B(sreg[1155]), .Z(n5835) );
  OR U6023 ( .A(n5833), .B(n5832), .Z(n5834) );
  AND U6024 ( .A(n5835), .B(n5834), .Z(n5873) );
  XOR U6025 ( .A(n5874), .B(n5873), .Z(c[1156]) );
  NANDN U6026 ( .A(n5837), .B(n5836), .Z(n5841) );
  NAND U6027 ( .A(n5839), .B(n5838), .Z(n5840) );
  NAND U6028 ( .A(n5841), .B(n5840), .Z(n5880) );
  NAND U6029 ( .A(b[0]), .B(a[141]), .Z(n5842) );
  XNOR U6030 ( .A(b[1]), .B(n5842), .Z(n5844) );
  NAND U6031 ( .A(n35), .B(a[140]), .Z(n5843) );
  AND U6032 ( .A(n5844), .B(n5843), .Z(n5897) );
  XOR U6033 ( .A(a[137]), .B(n42197), .Z(n5886) );
  NANDN U6034 ( .A(n5886), .B(n42173), .Z(n5847) );
  NANDN U6035 ( .A(n5845), .B(n42172), .Z(n5846) );
  NAND U6036 ( .A(n5847), .B(n5846), .Z(n5895) );
  NAND U6037 ( .A(b[7]), .B(a[133]), .Z(n5896) );
  XNOR U6038 ( .A(n5895), .B(n5896), .Z(n5898) );
  XOR U6039 ( .A(n5897), .B(n5898), .Z(n5904) );
  NANDN U6040 ( .A(n5848), .B(n42093), .Z(n5850) );
  XOR U6041 ( .A(n42134), .B(a[139]), .Z(n5889) );
  NANDN U6042 ( .A(n5889), .B(n42095), .Z(n5849) );
  NAND U6043 ( .A(n5850), .B(n5849), .Z(n5902) );
  NANDN U6044 ( .A(n5851), .B(n42231), .Z(n5853) );
  XOR U6045 ( .A(n173), .B(a[135]), .Z(n5892) );
  NANDN U6046 ( .A(n5892), .B(n42234), .Z(n5852) );
  AND U6047 ( .A(n5853), .B(n5852), .Z(n5901) );
  XNOR U6048 ( .A(n5902), .B(n5901), .Z(n5903) );
  XNOR U6049 ( .A(n5904), .B(n5903), .Z(n5908) );
  NANDN U6050 ( .A(n5855), .B(n5854), .Z(n5859) );
  NAND U6051 ( .A(n5857), .B(n5856), .Z(n5858) );
  AND U6052 ( .A(n5859), .B(n5858), .Z(n5907) );
  XOR U6053 ( .A(n5908), .B(n5907), .Z(n5909) );
  NANDN U6054 ( .A(n5861), .B(n5860), .Z(n5865) );
  NANDN U6055 ( .A(n5863), .B(n5862), .Z(n5864) );
  NAND U6056 ( .A(n5865), .B(n5864), .Z(n5910) );
  XOR U6057 ( .A(n5909), .B(n5910), .Z(n5877) );
  OR U6058 ( .A(n5867), .B(n5866), .Z(n5871) );
  NANDN U6059 ( .A(n5869), .B(n5868), .Z(n5870) );
  NAND U6060 ( .A(n5871), .B(n5870), .Z(n5878) );
  XNOR U6061 ( .A(n5877), .B(n5878), .Z(n5879) );
  XNOR U6062 ( .A(n5880), .B(n5879), .Z(n5913) );
  XNOR U6063 ( .A(n5913), .B(sreg[1157]), .Z(n5915) );
  NAND U6064 ( .A(n5872), .B(sreg[1156]), .Z(n5876) );
  OR U6065 ( .A(n5874), .B(n5873), .Z(n5875) );
  AND U6066 ( .A(n5876), .B(n5875), .Z(n5914) );
  XOR U6067 ( .A(n5915), .B(n5914), .Z(c[1157]) );
  NANDN U6068 ( .A(n5878), .B(n5877), .Z(n5882) );
  NAND U6069 ( .A(n5880), .B(n5879), .Z(n5881) );
  NAND U6070 ( .A(n5882), .B(n5881), .Z(n5921) );
  NAND U6071 ( .A(b[0]), .B(a[142]), .Z(n5883) );
  XNOR U6072 ( .A(b[1]), .B(n5883), .Z(n5885) );
  NAND U6073 ( .A(n35), .B(a[141]), .Z(n5884) );
  AND U6074 ( .A(n5885), .B(n5884), .Z(n5938) );
  XOR U6075 ( .A(a[138]), .B(n42197), .Z(n5927) );
  NANDN U6076 ( .A(n5927), .B(n42173), .Z(n5888) );
  NANDN U6077 ( .A(n5886), .B(n42172), .Z(n5887) );
  NAND U6078 ( .A(n5888), .B(n5887), .Z(n5936) );
  NAND U6079 ( .A(b[7]), .B(a[134]), .Z(n5937) );
  XNOR U6080 ( .A(n5936), .B(n5937), .Z(n5939) );
  XOR U6081 ( .A(n5938), .B(n5939), .Z(n5945) );
  NANDN U6082 ( .A(n5889), .B(n42093), .Z(n5891) );
  XOR U6083 ( .A(n42134), .B(a[140]), .Z(n5930) );
  NANDN U6084 ( .A(n5930), .B(n42095), .Z(n5890) );
  NAND U6085 ( .A(n5891), .B(n5890), .Z(n5943) );
  NANDN U6086 ( .A(n5892), .B(n42231), .Z(n5894) );
  XOR U6087 ( .A(n173), .B(a[136]), .Z(n5933) );
  NANDN U6088 ( .A(n5933), .B(n42234), .Z(n5893) );
  AND U6089 ( .A(n5894), .B(n5893), .Z(n5942) );
  XNOR U6090 ( .A(n5943), .B(n5942), .Z(n5944) );
  XNOR U6091 ( .A(n5945), .B(n5944), .Z(n5949) );
  NANDN U6092 ( .A(n5896), .B(n5895), .Z(n5900) );
  NAND U6093 ( .A(n5898), .B(n5897), .Z(n5899) );
  AND U6094 ( .A(n5900), .B(n5899), .Z(n5948) );
  XOR U6095 ( .A(n5949), .B(n5948), .Z(n5950) );
  NANDN U6096 ( .A(n5902), .B(n5901), .Z(n5906) );
  NANDN U6097 ( .A(n5904), .B(n5903), .Z(n5905) );
  NAND U6098 ( .A(n5906), .B(n5905), .Z(n5951) );
  XOR U6099 ( .A(n5950), .B(n5951), .Z(n5918) );
  OR U6100 ( .A(n5908), .B(n5907), .Z(n5912) );
  NANDN U6101 ( .A(n5910), .B(n5909), .Z(n5911) );
  NAND U6102 ( .A(n5912), .B(n5911), .Z(n5919) );
  XNOR U6103 ( .A(n5918), .B(n5919), .Z(n5920) );
  XNOR U6104 ( .A(n5921), .B(n5920), .Z(n5954) );
  XNOR U6105 ( .A(n5954), .B(sreg[1158]), .Z(n5956) );
  NAND U6106 ( .A(n5913), .B(sreg[1157]), .Z(n5917) );
  OR U6107 ( .A(n5915), .B(n5914), .Z(n5916) );
  AND U6108 ( .A(n5917), .B(n5916), .Z(n5955) );
  XOR U6109 ( .A(n5956), .B(n5955), .Z(c[1158]) );
  NANDN U6110 ( .A(n5919), .B(n5918), .Z(n5923) );
  NAND U6111 ( .A(n5921), .B(n5920), .Z(n5922) );
  NAND U6112 ( .A(n5923), .B(n5922), .Z(n5962) );
  NAND U6113 ( .A(b[0]), .B(a[143]), .Z(n5924) );
  XNOR U6114 ( .A(b[1]), .B(n5924), .Z(n5926) );
  NAND U6115 ( .A(n35), .B(a[142]), .Z(n5925) );
  AND U6116 ( .A(n5926), .B(n5925), .Z(n5979) );
  XOR U6117 ( .A(a[139]), .B(n42197), .Z(n5968) );
  NANDN U6118 ( .A(n5968), .B(n42173), .Z(n5929) );
  NANDN U6119 ( .A(n5927), .B(n42172), .Z(n5928) );
  NAND U6120 ( .A(n5929), .B(n5928), .Z(n5977) );
  NAND U6121 ( .A(b[7]), .B(a[135]), .Z(n5978) );
  XNOR U6122 ( .A(n5977), .B(n5978), .Z(n5980) );
  XOR U6123 ( .A(n5979), .B(n5980), .Z(n5986) );
  NANDN U6124 ( .A(n5930), .B(n42093), .Z(n5932) );
  XOR U6125 ( .A(n42134), .B(a[141]), .Z(n5971) );
  NANDN U6126 ( .A(n5971), .B(n42095), .Z(n5931) );
  NAND U6127 ( .A(n5932), .B(n5931), .Z(n5984) );
  NANDN U6128 ( .A(n5933), .B(n42231), .Z(n5935) );
  XOR U6129 ( .A(n173), .B(a[137]), .Z(n5974) );
  NANDN U6130 ( .A(n5974), .B(n42234), .Z(n5934) );
  AND U6131 ( .A(n5935), .B(n5934), .Z(n5983) );
  XNOR U6132 ( .A(n5984), .B(n5983), .Z(n5985) );
  XNOR U6133 ( .A(n5986), .B(n5985), .Z(n5990) );
  NANDN U6134 ( .A(n5937), .B(n5936), .Z(n5941) );
  NAND U6135 ( .A(n5939), .B(n5938), .Z(n5940) );
  AND U6136 ( .A(n5941), .B(n5940), .Z(n5989) );
  XOR U6137 ( .A(n5990), .B(n5989), .Z(n5991) );
  NANDN U6138 ( .A(n5943), .B(n5942), .Z(n5947) );
  NANDN U6139 ( .A(n5945), .B(n5944), .Z(n5946) );
  NAND U6140 ( .A(n5947), .B(n5946), .Z(n5992) );
  XOR U6141 ( .A(n5991), .B(n5992), .Z(n5959) );
  OR U6142 ( .A(n5949), .B(n5948), .Z(n5953) );
  NANDN U6143 ( .A(n5951), .B(n5950), .Z(n5952) );
  NAND U6144 ( .A(n5953), .B(n5952), .Z(n5960) );
  XNOR U6145 ( .A(n5959), .B(n5960), .Z(n5961) );
  XNOR U6146 ( .A(n5962), .B(n5961), .Z(n5995) );
  XNOR U6147 ( .A(n5995), .B(sreg[1159]), .Z(n5997) );
  NAND U6148 ( .A(n5954), .B(sreg[1158]), .Z(n5958) );
  OR U6149 ( .A(n5956), .B(n5955), .Z(n5957) );
  AND U6150 ( .A(n5958), .B(n5957), .Z(n5996) );
  XOR U6151 ( .A(n5997), .B(n5996), .Z(c[1159]) );
  NANDN U6152 ( .A(n5960), .B(n5959), .Z(n5964) );
  NAND U6153 ( .A(n5962), .B(n5961), .Z(n5963) );
  NAND U6154 ( .A(n5964), .B(n5963), .Z(n6003) );
  NAND U6155 ( .A(b[0]), .B(a[144]), .Z(n5965) );
  XNOR U6156 ( .A(b[1]), .B(n5965), .Z(n5967) );
  NAND U6157 ( .A(n35), .B(a[143]), .Z(n5966) );
  AND U6158 ( .A(n5967), .B(n5966), .Z(n6020) );
  XOR U6159 ( .A(a[140]), .B(n42197), .Z(n6009) );
  NANDN U6160 ( .A(n6009), .B(n42173), .Z(n5970) );
  NANDN U6161 ( .A(n5968), .B(n42172), .Z(n5969) );
  NAND U6162 ( .A(n5970), .B(n5969), .Z(n6018) );
  NAND U6163 ( .A(b[7]), .B(a[136]), .Z(n6019) );
  XNOR U6164 ( .A(n6018), .B(n6019), .Z(n6021) );
  XOR U6165 ( .A(n6020), .B(n6021), .Z(n6027) );
  NANDN U6166 ( .A(n5971), .B(n42093), .Z(n5973) );
  XOR U6167 ( .A(n42134), .B(a[142]), .Z(n6012) );
  NANDN U6168 ( .A(n6012), .B(n42095), .Z(n5972) );
  NAND U6169 ( .A(n5973), .B(n5972), .Z(n6025) );
  NANDN U6170 ( .A(n5974), .B(n42231), .Z(n5976) );
  XOR U6171 ( .A(n173), .B(a[138]), .Z(n6015) );
  NANDN U6172 ( .A(n6015), .B(n42234), .Z(n5975) );
  AND U6173 ( .A(n5976), .B(n5975), .Z(n6024) );
  XNOR U6174 ( .A(n6025), .B(n6024), .Z(n6026) );
  XNOR U6175 ( .A(n6027), .B(n6026), .Z(n6031) );
  NANDN U6176 ( .A(n5978), .B(n5977), .Z(n5982) );
  NAND U6177 ( .A(n5980), .B(n5979), .Z(n5981) );
  AND U6178 ( .A(n5982), .B(n5981), .Z(n6030) );
  XOR U6179 ( .A(n6031), .B(n6030), .Z(n6032) );
  NANDN U6180 ( .A(n5984), .B(n5983), .Z(n5988) );
  NANDN U6181 ( .A(n5986), .B(n5985), .Z(n5987) );
  NAND U6182 ( .A(n5988), .B(n5987), .Z(n6033) );
  XOR U6183 ( .A(n6032), .B(n6033), .Z(n6000) );
  OR U6184 ( .A(n5990), .B(n5989), .Z(n5994) );
  NANDN U6185 ( .A(n5992), .B(n5991), .Z(n5993) );
  NAND U6186 ( .A(n5994), .B(n5993), .Z(n6001) );
  XNOR U6187 ( .A(n6000), .B(n6001), .Z(n6002) );
  XNOR U6188 ( .A(n6003), .B(n6002), .Z(n6036) );
  XNOR U6189 ( .A(n6036), .B(sreg[1160]), .Z(n6038) );
  NAND U6190 ( .A(n5995), .B(sreg[1159]), .Z(n5999) );
  OR U6191 ( .A(n5997), .B(n5996), .Z(n5998) );
  AND U6192 ( .A(n5999), .B(n5998), .Z(n6037) );
  XOR U6193 ( .A(n6038), .B(n6037), .Z(c[1160]) );
  NANDN U6194 ( .A(n6001), .B(n6000), .Z(n6005) );
  NAND U6195 ( .A(n6003), .B(n6002), .Z(n6004) );
  NAND U6196 ( .A(n6005), .B(n6004), .Z(n6044) );
  NAND U6197 ( .A(b[0]), .B(a[145]), .Z(n6006) );
  XNOR U6198 ( .A(b[1]), .B(n6006), .Z(n6008) );
  NAND U6199 ( .A(n35), .B(a[144]), .Z(n6007) );
  AND U6200 ( .A(n6008), .B(n6007), .Z(n6061) );
  XOR U6201 ( .A(a[141]), .B(n42197), .Z(n6050) );
  NANDN U6202 ( .A(n6050), .B(n42173), .Z(n6011) );
  NANDN U6203 ( .A(n6009), .B(n42172), .Z(n6010) );
  NAND U6204 ( .A(n6011), .B(n6010), .Z(n6059) );
  NAND U6205 ( .A(b[7]), .B(a[137]), .Z(n6060) );
  XNOR U6206 ( .A(n6059), .B(n6060), .Z(n6062) );
  XOR U6207 ( .A(n6061), .B(n6062), .Z(n6068) );
  NANDN U6208 ( .A(n6012), .B(n42093), .Z(n6014) );
  XOR U6209 ( .A(n42134), .B(a[143]), .Z(n6053) );
  NANDN U6210 ( .A(n6053), .B(n42095), .Z(n6013) );
  NAND U6211 ( .A(n6014), .B(n6013), .Z(n6066) );
  NANDN U6212 ( .A(n6015), .B(n42231), .Z(n6017) );
  XOR U6213 ( .A(n173), .B(a[139]), .Z(n6056) );
  NANDN U6214 ( .A(n6056), .B(n42234), .Z(n6016) );
  AND U6215 ( .A(n6017), .B(n6016), .Z(n6065) );
  XNOR U6216 ( .A(n6066), .B(n6065), .Z(n6067) );
  XNOR U6217 ( .A(n6068), .B(n6067), .Z(n6072) );
  NANDN U6218 ( .A(n6019), .B(n6018), .Z(n6023) );
  NAND U6219 ( .A(n6021), .B(n6020), .Z(n6022) );
  AND U6220 ( .A(n6023), .B(n6022), .Z(n6071) );
  XOR U6221 ( .A(n6072), .B(n6071), .Z(n6073) );
  NANDN U6222 ( .A(n6025), .B(n6024), .Z(n6029) );
  NANDN U6223 ( .A(n6027), .B(n6026), .Z(n6028) );
  NAND U6224 ( .A(n6029), .B(n6028), .Z(n6074) );
  XOR U6225 ( .A(n6073), .B(n6074), .Z(n6041) );
  OR U6226 ( .A(n6031), .B(n6030), .Z(n6035) );
  NANDN U6227 ( .A(n6033), .B(n6032), .Z(n6034) );
  NAND U6228 ( .A(n6035), .B(n6034), .Z(n6042) );
  XNOR U6229 ( .A(n6041), .B(n6042), .Z(n6043) );
  XNOR U6230 ( .A(n6044), .B(n6043), .Z(n6077) );
  XNOR U6231 ( .A(n6077), .B(sreg[1161]), .Z(n6079) );
  NAND U6232 ( .A(n6036), .B(sreg[1160]), .Z(n6040) );
  OR U6233 ( .A(n6038), .B(n6037), .Z(n6039) );
  AND U6234 ( .A(n6040), .B(n6039), .Z(n6078) );
  XOR U6235 ( .A(n6079), .B(n6078), .Z(c[1161]) );
  NANDN U6236 ( .A(n6042), .B(n6041), .Z(n6046) );
  NAND U6237 ( .A(n6044), .B(n6043), .Z(n6045) );
  NAND U6238 ( .A(n6046), .B(n6045), .Z(n6085) );
  NAND U6239 ( .A(b[0]), .B(a[146]), .Z(n6047) );
  XNOR U6240 ( .A(b[1]), .B(n6047), .Z(n6049) );
  NAND U6241 ( .A(n35), .B(a[145]), .Z(n6048) );
  AND U6242 ( .A(n6049), .B(n6048), .Z(n6102) );
  XOR U6243 ( .A(a[142]), .B(n42197), .Z(n6091) );
  NANDN U6244 ( .A(n6091), .B(n42173), .Z(n6052) );
  NANDN U6245 ( .A(n6050), .B(n42172), .Z(n6051) );
  NAND U6246 ( .A(n6052), .B(n6051), .Z(n6100) );
  NAND U6247 ( .A(b[7]), .B(a[138]), .Z(n6101) );
  XNOR U6248 ( .A(n6100), .B(n6101), .Z(n6103) );
  XOR U6249 ( .A(n6102), .B(n6103), .Z(n6109) );
  NANDN U6250 ( .A(n6053), .B(n42093), .Z(n6055) );
  XOR U6251 ( .A(n42134), .B(a[144]), .Z(n6094) );
  NANDN U6252 ( .A(n6094), .B(n42095), .Z(n6054) );
  NAND U6253 ( .A(n6055), .B(n6054), .Z(n6107) );
  NANDN U6254 ( .A(n6056), .B(n42231), .Z(n6058) );
  XOR U6255 ( .A(n173), .B(a[140]), .Z(n6097) );
  NANDN U6256 ( .A(n6097), .B(n42234), .Z(n6057) );
  AND U6257 ( .A(n6058), .B(n6057), .Z(n6106) );
  XNOR U6258 ( .A(n6107), .B(n6106), .Z(n6108) );
  XNOR U6259 ( .A(n6109), .B(n6108), .Z(n6113) );
  NANDN U6260 ( .A(n6060), .B(n6059), .Z(n6064) );
  NAND U6261 ( .A(n6062), .B(n6061), .Z(n6063) );
  AND U6262 ( .A(n6064), .B(n6063), .Z(n6112) );
  XOR U6263 ( .A(n6113), .B(n6112), .Z(n6114) );
  NANDN U6264 ( .A(n6066), .B(n6065), .Z(n6070) );
  NANDN U6265 ( .A(n6068), .B(n6067), .Z(n6069) );
  NAND U6266 ( .A(n6070), .B(n6069), .Z(n6115) );
  XOR U6267 ( .A(n6114), .B(n6115), .Z(n6082) );
  OR U6268 ( .A(n6072), .B(n6071), .Z(n6076) );
  NANDN U6269 ( .A(n6074), .B(n6073), .Z(n6075) );
  NAND U6270 ( .A(n6076), .B(n6075), .Z(n6083) );
  XNOR U6271 ( .A(n6082), .B(n6083), .Z(n6084) );
  XNOR U6272 ( .A(n6085), .B(n6084), .Z(n6118) );
  XNOR U6273 ( .A(n6118), .B(sreg[1162]), .Z(n6120) );
  NAND U6274 ( .A(n6077), .B(sreg[1161]), .Z(n6081) );
  OR U6275 ( .A(n6079), .B(n6078), .Z(n6080) );
  AND U6276 ( .A(n6081), .B(n6080), .Z(n6119) );
  XOR U6277 ( .A(n6120), .B(n6119), .Z(c[1162]) );
  NANDN U6278 ( .A(n6083), .B(n6082), .Z(n6087) );
  NAND U6279 ( .A(n6085), .B(n6084), .Z(n6086) );
  NAND U6280 ( .A(n6087), .B(n6086), .Z(n6126) );
  NAND U6281 ( .A(b[0]), .B(a[147]), .Z(n6088) );
  XNOR U6282 ( .A(b[1]), .B(n6088), .Z(n6090) );
  NAND U6283 ( .A(n36), .B(a[146]), .Z(n6089) );
  AND U6284 ( .A(n6090), .B(n6089), .Z(n6143) );
  XOR U6285 ( .A(a[143]), .B(n42197), .Z(n6132) );
  NANDN U6286 ( .A(n6132), .B(n42173), .Z(n6093) );
  NANDN U6287 ( .A(n6091), .B(n42172), .Z(n6092) );
  NAND U6288 ( .A(n6093), .B(n6092), .Z(n6141) );
  NAND U6289 ( .A(b[7]), .B(a[139]), .Z(n6142) );
  XNOR U6290 ( .A(n6141), .B(n6142), .Z(n6144) );
  XOR U6291 ( .A(n6143), .B(n6144), .Z(n6150) );
  NANDN U6292 ( .A(n6094), .B(n42093), .Z(n6096) );
  XOR U6293 ( .A(n42134), .B(a[145]), .Z(n6135) );
  NANDN U6294 ( .A(n6135), .B(n42095), .Z(n6095) );
  NAND U6295 ( .A(n6096), .B(n6095), .Z(n6148) );
  NANDN U6296 ( .A(n6097), .B(n42231), .Z(n6099) );
  XOR U6297 ( .A(n173), .B(a[141]), .Z(n6138) );
  NANDN U6298 ( .A(n6138), .B(n42234), .Z(n6098) );
  AND U6299 ( .A(n6099), .B(n6098), .Z(n6147) );
  XNOR U6300 ( .A(n6148), .B(n6147), .Z(n6149) );
  XNOR U6301 ( .A(n6150), .B(n6149), .Z(n6154) );
  NANDN U6302 ( .A(n6101), .B(n6100), .Z(n6105) );
  NAND U6303 ( .A(n6103), .B(n6102), .Z(n6104) );
  AND U6304 ( .A(n6105), .B(n6104), .Z(n6153) );
  XOR U6305 ( .A(n6154), .B(n6153), .Z(n6155) );
  NANDN U6306 ( .A(n6107), .B(n6106), .Z(n6111) );
  NANDN U6307 ( .A(n6109), .B(n6108), .Z(n6110) );
  NAND U6308 ( .A(n6111), .B(n6110), .Z(n6156) );
  XOR U6309 ( .A(n6155), .B(n6156), .Z(n6123) );
  OR U6310 ( .A(n6113), .B(n6112), .Z(n6117) );
  NANDN U6311 ( .A(n6115), .B(n6114), .Z(n6116) );
  NAND U6312 ( .A(n6117), .B(n6116), .Z(n6124) );
  XNOR U6313 ( .A(n6123), .B(n6124), .Z(n6125) );
  XNOR U6314 ( .A(n6126), .B(n6125), .Z(n6159) );
  XNOR U6315 ( .A(n6159), .B(sreg[1163]), .Z(n6161) );
  NAND U6316 ( .A(n6118), .B(sreg[1162]), .Z(n6122) );
  OR U6317 ( .A(n6120), .B(n6119), .Z(n6121) );
  AND U6318 ( .A(n6122), .B(n6121), .Z(n6160) );
  XOR U6319 ( .A(n6161), .B(n6160), .Z(c[1163]) );
  NANDN U6320 ( .A(n6124), .B(n6123), .Z(n6128) );
  NAND U6321 ( .A(n6126), .B(n6125), .Z(n6127) );
  NAND U6322 ( .A(n6128), .B(n6127), .Z(n6167) );
  NAND U6323 ( .A(b[0]), .B(a[148]), .Z(n6129) );
  XNOR U6324 ( .A(b[1]), .B(n6129), .Z(n6131) );
  NAND U6325 ( .A(n36), .B(a[147]), .Z(n6130) );
  AND U6326 ( .A(n6131), .B(n6130), .Z(n6184) );
  XOR U6327 ( .A(a[144]), .B(n42197), .Z(n6173) );
  NANDN U6328 ( .A(n6173), .B(n42173), .Z(n6134) );
  NANDN U6329 ( .A(n6132), .B(n42172), .Z(n6133) );
  NAND U6330 ( .A(n6134), .B(n6133), .Z(n6182) );
  NAND U6331 ( .A(b[7]), .B(a[140]), .Z(n6183) );
  XNOR U6332 ( .A(n6182), .B(n6183), .Z(n6185) );
  XOR U6333 ( .A(n6184), .B(n6185), .Z(n6191) );
  NANDN U6334 ( .A(n6135), .B(n42093), .Z(n6137) );
  XOR U6335 ( .A(n42134), .B(a[146]), .Z(n6176) );
  NANDN U6336 ( .A(n6176), .B(n42095), .Z(n6136) );
  NAND U6337 ( .A(n6137), .B(n6136), .Z(n6189) );
  NANDN U6338 ( .A(n6138), .B(n42231), .Z(n6140) );
  XOR U6339 ( .A(n173), .B(a[142]), .Z(n6179) );
  NANDN U6340 ( .A(n6179), .B(n42234), .Z(n6139) );
  AND U6341 ( .A(n6140), .B(n6139), .Z(n6188) );
  XNOR U6342 ( .A(n6189), .B(n6188), .Z(n6190) );
  XNOR U6343 ( .A(n6191), .B(n6190), .Z(n6195) );
  NANDN U6344 ( .A(n6142), .B(n6141), .Z(n6146) );
  NAND U6345 ( .A(n6144), .B(n6143), .Z(n6145) );
  AND U6346 ( .A(n6146), .B(n6145), .Z(n6194) );
  XOR U6347 ( .A(n6195), .B(n6194), .Z(n6196) );
  NANDN U6348 ( .A(n6148), .B(n6147), .Z(n6152) );
  NANDN U6349 ( .A(n6150), .B(n6149), .Z(n6151) );
  NAND U6350 ( .A(n6152), .B(n6151), .Z(n6197) );
  XOR U6351 ( .A(n6196), .B(n6197), .Z(n6164) );
  OR U6352 ( .A(n6154), .B(n6153), .Z(n6158) );
  NANDN U6353 ( .A(n6156), .B(n6155), .Z(n6157) );
  NAND U6354 ( .A(n6158), .B(n6157), .Z(n6165) );
  XNOR U6355 ( .A(n6164), .B(n6165), .Z(n6166) );
  XNOR U6356 ( .A(n6167), .B(n6166), .Z(n6200) );
  XNOR U6357 ( .A(n6200), .B(sreg[1164]), .Z(n6202) );
  NAND U6358 ( .A(n6159), .B(sreg[1163]), .Z(n6163) );
  OR U6359 ( .A(n6161), .B(n6160), .Z(n6162) );
  AND U6360 ( .A(n6163), .B(n6162), .Z(n6201) );
  XOR U6361 ( .A(n6202), .B(n6201), .Z(c[1164]) );
  NANDN U6362 ( .A(n6165), .B(n6164), .Z(n6169) );
  NAND U6363 ( .A(n6167), .B(n6166), .Z(n6168) );
  NAND U6364 ( .A(n6169), .B(n6168), .Z(n6208) );
  NAND U6365 ( .A(b[0]), .B(a[149]), .Z(n6170) );
  XNOR U6366 ( .A(b[1]), .B(n6170), .Z(n6172) );
  NAND U6367 ( .A(n36), .B(a[148]), .Z(n6171) );
  AND U6368 ( .A(n6172), .B(n6171), .Z(n6225) );
  XOR U6369 ( .A(a[145]), .B(n42197), .Z(n6214) );
  NANDN U6370 ( .A(n6214), .B(n42173), .Z(n6175) );
  NANDN U6371 ( .A(n6173), .B(n42172), .Z(n6174) );
  NAND U6372 ( .A(n6175), .B(n6174), .Z(n6223) );
  NAND U6373 ( .A(b[7]), .B(a[141]), .Z(n6224) );
  XNOR U6374 ( .A(n6223), .B(n6224), .Z(n6226) );
  XOR U6375 ( .A(n6225), .B(n6226), .Z(n6232) );
  NANDN U6376 ( .A(n6176), .B(n42093), .Z(n6178) );
  XOR U6377 ( .A(n42134), .B(a[147]), .Z(n6217) );
  NANDN U6378 ( .A(n6217), .B(n42095), .Z(n6177) );
  NAND U6379 ( .A(n6178), .B(n6177), .Z(n6230) );
  NANDN U6380 ( .A(n6179), .B(n42231), .Z(n6181) );
  XOR U6381 ( .A(n174), .B(a[143]), .Z(n6220) );
  NANDN U6382 ( .A(n6220), .B(n42234), .Z(n6180) );
  AND U6383 ( .A(n6181), .B(n6180), .Z(n6229) );
  XNOR U6384 ( .A(n6230), .B(n6229), .Z(n6231) );
  XNOR U6385 ( .A(n6232), .B(n6231), .Z(n6236) );
  NANDN U6386 ( .A(n6183), .B(n6182), .Z(n6187) );
  NAND U6387 ( .A(n6185), .B(n6184), .Z(n6186) );
  AND U6388 ( .A(n6187), .B(n6186), .Z(n6235) );
  XOR U6389 ( .A(n6236), .B(n6235), .Z(n6237) );
  NANDN U6390 ( .A(n6189), .B(n6188), .Z(n6193) );
  NANDN U6391 ( .A(n6191), .B(n6190), .Z(n6192) );
  NAND U6392 ( .A(n6193), .B(n6192), .Z(n6238) );
  XOR U6393 ( .A(n6237), .B(n6238), .Z(n6205) );
  OR U6394 ( .A(n6195), .B(n6194), .Z(n6199) );
  NANDN U6395 ( .A(n6197), .B(n6196), .Z(n6198) );
  NAND U6396 ( .A(n6199), .B(n6198), .Z(n6206) );
  XNOR U6397 ( .A(n6205), .B(n6206), .Z(n6207) );
  XNOR U6398 ( .A(n6208), .B(n6207), .Z(n6241) );
  XNOR U6399 ( .A(n6241), .B(sreg[1165]), .Z(n6243) );
  NAND U6400 ( .A(n6200), .B(sreg[1164]), .Z(n6204) );
  OR U6401 ( .A(n6202), .B(n6201), .Z(n6203) );
  AND U6402 ( .A(n6204), .B(n6203), .Z(n6242) );
  XOR U6403 ( .A(n6243), .B(n6242), .Z(c[1165]) );
  NANDN U6404 ( .A(n6206), .B(n6205), .Z(n6210) );
  NAND U6405 ( .A(n6208), .B(n6207), .Z(n6209) );
  NAND U6406 ( .A(n6210), .B(n6209), .Z(n6249) );
  NAND U6407 ( .A(b[0]), .B(a[150]), .Z(n6211) );
  XNOR U6408 ( .A(b[1]), .B(n6211), .Z(n6213) );
  NAND U6409 ( .A(n36), .B(a[149]), .Z(n6212) );
  AND U6410 ( .A(n6213), .B(n6212), .Z(n6266) );
  XOR U6411 ( .A(a[146]), .B(n42197), .Z(n6255) );
  NANDN U6412 ( .A(n6255), .B(n42173), .Z(n6216) );
  NANDN U6413 ( .A(n6214), .B(n42172), .Z(n6215) );
  NAND U6414 ( .A(n6216), .B(n6215), .Z(n6264) );
  NAND U6415 ( .A(b[7]), .B(a[142]), .Z(n6265) );
  XNOR U6416 ( .A(n6264), .B(n6265), .Z(n6267) );
  XOR U6417 ( .A(n6266), .B(n6267), .Z(n6273) );
  NANDN U6418 ( .A(n6217), .B(n42093), .Z(n6219) );
  XOR U6419 ( .A(n42134), .B(a[148]), .Z(n6258) );
  NANDN U6420 ( .A(n6258), .B(n42095), .Z(n6218) );
  NAND U6421 ( .A(n6219), .B(n6218), .Z(n6271) );
  NANDN U6422 ( .A(n6220), .B(n42231), .Z(n6222) );
  XOR U6423 ( .A(n174), .B(a[144]), .Z(n6261) );
  NANDN U6424 ( .A(n6261), .B(n42234), .Z(n6221) );
  AND U6425 ( .A(n6222), .B(n6221), .Z(n6270) );
  XNOR U6426 ( .A(n6271), .B(n6270), .Z(n6272) );
  XNOR U6427 ( .A(n6273), .B(n6272), .Z(n6277) );
  NANDN U6428 ( .A(n6224), .B(n6223), .Z(n6228) );
  NAND U6429 ( .A(n6226), .B(n6225), .Z(n6227) );
  AND U6430 ( .A(n6228), .B(n6227), .Z(n6276) );
  XOR U6431 ( .A(n6277), .B(n6276), .Z(n6278) );
  NANDN U6432 ( .A(n6230), .B(n6229), .Z(n6234) );
  NANDN U6433 ( .A(n6232), .B(n6231), .Z(n6233) );
  NAND U6434 ( .A(n6234), .B(n6233), .Z(n6279) );
  XOR U6435 ( .A(n6278), .B(n6279), .Z(n6246) );
  OR U6436 ( .A(n6236), .B(n6235), .Z(n6240) );
  NANDN U6437 ( .A(n6238), .B(n6237), .Z(n6239) );
  NAND U6438 ( .A(n6240), .B(n6239), .Z(n6247) );
  XNOR U6439 ( .A(n6246), .B(n6247), .Z(n6248) );
  XNOR U6440 ( .A(n6249), .B(n6248), .Z(n6282) );
  XNOR U6441 ( .A(n6282), .B(sreg[1166]), .Z(n6284) );
  NAND U6442 ( .A(n6241), .B(sreg[1165]), .Z(n6245) );
  OR U6443 ( .A(n6243), .B(n6242), .Z(n6244) );
  AND U6444 ( .A(n6245), .B(n6244), .Z(n6283) );
  XOR U6445 ( .A(n6284), .B(n6283), .Z(c[1166]) );
  NANDN U6446 ( .A(n6247), .B(n6246), .Z(n6251) );
  NAND U6447 ( .A(n6249), .B(n6248), .Z(n6250) );
  NAND U6448 ( .A(n6251), .B(n6250), .Z(n6290) );
  NAND U6449 ( .A(b[0]), .B(a[151]), .Z(n6252) );
  XNOR U6450 ( .A(b[1]), .B(n6252), .Z(n6254) );
  NAND U6451 ( .A(n36), .B(a[150]), .Z(n6253) );
  AND U6452 ( .A(n6254), .B(n6253), .Z(n6307) );
  XOR U6453 ( .A(a[147]), .B(n42197), .Z(n6296) );
  NANDN U6454 ( .A(n6296), .B(n42173), .Z(n6257) );
  NANDN U6455 ( .A(n6255), .B(n42172), .Z(n6256) );
  NAND U6456 ( .A(n6257), .B(n6256), .Z(n6305) );
  NAND U6457 ( .A(b[7]), .B(a[143]), .Z(n6306) );
  XNOR U6458 ( .A(n6305), .B(n6306), .Z(n6308) );
  XOR U6459 ( .A(n6307), .B(n6308), .Z(n6314) );
  NANDN U6460 ( .A(n6258), .B(n42093), .Z(n6260) );
  XOR U6461 ( .A(n42134), .B(a[149]), .Z(n6299) );
  NANDN U6462 ( .A(n6299), .B(n42095), .Z(n6259) );
  NAND U6463 ( .A(n6260), .B(n6259), .Z(n6312) );
  NANDN U6464 ( .A(n6261), .B(n42231), .Z(n6263) );
  XOR U6465 ( .A(n174), .B(a[145]), .Z(n6302) );
  NANDN U6466 ( .A(n6302), .B(n42234), .Z(n6262) );
  AND U6467 ( .A(n6263), .B(n6262), .Z(n6311) );
  XNOR U6468 ( .A(n6312), .B(n6311), .Z(n6313) );
  XNOR U6469 ( .A(n6314), .B(n6313), .Z(n6318) );
  NANDN U6470 ( .A(n6265), .B(n6264), .Z(n6269) );
  NAND U6471 ( .A(n6267), .B(n6266), .Z(n6268) );
  AND U6472 ( .A(n6269), .B(n6268), .Z(n6317) );
  XOR U6473 ( .A(n6318), .B(n6317), .Z(n6319) );
  NANDN U6474 ( .A(n6271), .B(n6270), .Z(n6275) );
  NANDN U6475 ( .A(n6273), .B(n6272), .Z(n6274) );
  NAND U6476 ( .A(n6275), .B(n6274), .Z(n6320) );
  XOR U6477 ( .A(n6319), .B(n6320), .Z(n6287) );
  OR U6478 ( .A(n6277), .B(n6276), .Z(n6281) );
  NANDN U6479 ( .A(n6279), .B(n6278), .Z(n6280) );
  NAND U6480 ( .A(n6281), .B(n6280), .Z(n6288) );
  XNOR U6481 ( .A(n6287), .B(n6288), .Z(n6289) );
  XNOR U6482 ( .A(n6290), .B(n6289), .Z(n6323) );
  XNOR U6483 ( .A(n6323), .B(sreg[1167]), .Z(n6325) );
  NAND U6484 ( .A(n6282), .B(sreg[1166]), .Z(n6286) );
  OR U6485 ( .A(n6284), .B(n6283), .Z(n6285) );
  AND U6486 ( .A(n6286), .B(n6285), .Z(n6324) );
  XOR U6487 ( .A(n6325), .B(n6324), .Z(c[1167]) );
  NANDN U6488 ( .A(n6288), .B(n6287), .Z(n6292) );
  NAND U6489 ( .A(n6290), .B(n6289), .Z(n6291) );
  NAND U6490 ( .A(n6292), .B(n6291), .Z(n6331) );
  NAND U6491 ( .A(b[0]), .B(a[152]), .Z(n6293) );
  XNOR U6492 ( .A(b[1]), .B(n6293), .Z(n6295) );
  NAND U6493 ( .A(n36), .B(a[151]), .Z(n6294) );
  AND U6494 ( .A(n6295), .B(n6294), .Z(n6348) );
  XOR U6495 ( .A(a[148]), .B(n42197), .Z(n6337) );
  NANDN U6496 ( .A(n6337), .B(n42173), .Z(n6298) );
  NANDN U6497 ( .A(n6296), .B(n42172), .Z(n6297) );
  NAND U6498 ( .A(n6298), .B(n6297), .Z(n6346) );
  NAND U6499 ( .A(b[7]), .B(a[144]), .Z(n6347) );
  XNOR U6500 ( .A(n6346), .B(n6347), .Z(n6349) );
  XOR U6501 ( .A(n6348), .B(n6349), .Z(n6355) );
  NANDN U6502 ( .A(n6299), .B(n42093), .Z(n6301) );
  XOR U6503 ( .A(n42134), .B(a[150]), .Z(n6340) );
  NANDN U6504 ( .A(n6340), .B(n42095), .Z(n6300) );
  NAND U6505 ( .A(n6301), .B(n6300), .Z(n6353) );
  NANDN U6506 ( .A(n6302), .B(n42231), .Z(n6304) );
  XOR U6507 ( .A(n174), .B(a[146]), .Z(n6343) );
  NANDN U6508 ( .A(n6343), .B(n42234), .Z(n6303) );
  AND U6509 ( .A(n6304), .B(n6303), .Z(n6352) );
  XNOR U6510 ( .A(n6353), .B(n6352), .Z(n6354) );
  XNOR U6511 ( .A(n6355), .B(n6354), .Z(n6359) );
  NANDN U6512 ( .A(n6306), .B(n6305), .Z(n6310) );
  NAND U6513 ( .A(n6308), .B(n6307), .Z(n6309) );
  AND U6514 ( .A(n6310), .B(n6309), .Z(n6358) );
  XOR U6515 ( .A(n6359), .B(n6358), .Z(n6360) );
  NANDN U6516 ( .A(n6312), .B(n6311), .Z(n6316) );
  NANDN U6517 ( .A(n6314), .B(n6313), .Z(n6315) );
  NAND U6518 ( .A(n6316), .B(n6315), .Z(n6361) );
  XOR U6519 ( .A(n6360), .B(n6361), .Z(n6328) );
  OR U6520 ( .A(n6318), .B(n6317), .Z(n6322) );
  NANDN U6521 ( .A(n6320), .B(n6319), .Z(n6321) );
  NAND U6522 ( .A(n6322), .B(n6321), .Z(n6329) );
  XNOR U6523 ( .A(n6328), .B(n6329), .Z(n6330) );
  XNOR U6524 ( .A(n6331), .B(n6330), .Z(n6364) );
  XNOR U6525 ( .A(n6364), .B(sreg[1168]), .Z(n6366) );
  NAND U6526 ( .A(n6323), .B(sreg[1167]), .Z(n6327) );
  OR U6527 ( .A(n6325), .B(n6324), .Z(n6326) );
  AND U6528 ( .A(n6327), .B(n6326), .Z(n6365) );
  XOR U6529 ( .A(n6366), .B(n6365), .Z(c[1168]) );
  NANDN U6530 ( .A(n6329), .B(n6328), .Z(n6333) );
  NAND U6531 ( .A(n6331), .B(n6330), .Z(n6332) );
  NAND U6532 ( .A(n6333), .B(n6332), .Z(n6372) );
  NAND U6533 ( .A(b[0]), .B(a[153]), .Z(n6334) );
  XNOR U6534 ( .A(b[1]), .B(n6334), .Z(n6336) );
  NAND U6535 ( .A(n36), .B(a[152]), .Z(n6335) );
  AND U6536 ( .A(n6336), .B(n6335), .Z(n6389) );
  XOR U6537 ( .A(a[149]), .B(n42197), .Z(n6378) );
  NANDN U6538 ( .A(n6378), .B(n42173), .Z(n6339) );
  NANDN U6539 ( .A(n6337), .B(n42172), .Z(n6338) );
  NAND U6540 ( .A(n6339), .B(n6338), .Z(n6387) );
  NAND U6541 ( .A(b[7]), .B(a[145]), .Z(n6388) );
  XNOR U6542 ( .A(n6387), .B(n6388), .Z(n6390) );
  XOR U6543 ( .A(n6389), .B(n6390), .Z(n6396) );
  NANDN U6544 ( .A(n6340), .B(n42093), .Z(n6342) );
  XOR U6545 ( .A(n42134), .B(a[151]), .Z(n6381) );
  NANDN U6546 ( .A(n6381), .B(n42095), .Z(n6341) );
  NAND U6547 ( .A(n6342), .B(n6341), .Z(n6394) );
  NANDN U6548 ( .A(n6343), .B(n42231), .Z(n6345) );
  XOR U6549 ( .A(n174), .B(a[147]), .Z(n6384) );
  NANDN U6550 ( .A(n6384), .B(n42234), .Z(n6344) );
  AND U6551 ( .A(n6345), .B(n6344), .Z(n6393) );
  XNOR U6552 ( .A(n6394), .B(n6393), .Z(n6395) );
  XNOR U6553 ( .A(n6396), .B(n6395), .Z(n6400) );
  NANDN U6554 ( .A(n6347), .B(n6346), .Z(n6351) );
  NAND U6555 ( .A(n6349), .B(n6348), .Z(n6350) );
  AND U6556 ( .A(n6351), .B(n6350), .Z(n6399) );
  XOR U6557 ( .A(n6400), .B(n6399), .Z(n6401) );
  NANDN U6558 ( .A(n6353), .B(n6352), .Z(n6357) );
  NANDN U6559 ( .A(n6355), .B(n6354), .Z(n6356) );
  NAND U6560 ( .A(n6357), .B(n6356), .Z(n6402) );
  XOR U6561 ( .A(n6401), .B(n6402), .Z(n6369) );
  OR U6562 ( .A(n6359), .B(n6358), .Z(n6363) );
  NANDN U6563 ( .A(n6361), .B(n6360), .Z(n6362) );
  NAND U6564 ( .A(n6363), .B(n6362), .Z(n6370) );
  XNOR U6565 ( .A(n6369), .B(n6370), .Z(n6371) );
  XNOR U6566 ( .A(n6372), .B(n6371), .Z(n6405) );
  XNOR U6567 ( .A(n6405), .B(sreg[1169]), .Z(n6407) );
  NAND U6568 ( .A(n6364), .B(sreg[1168]), .Z(n6368) );
  OR U6569 ( .A(n6366), .B(n6365), .Z(n6367) );
  AND U6570 ( .A(n6368), .B(n6367), .Z(n6406) );
  XOR U6571 ( .A(n6407), .B(n6406), .Z(c[1169]) );
  NANDN U6572 ( .A(n6370), .B(n6369), .Z(n6374) );
  NAND U6573 ( .A(n6372), .B(n6371), .Z(n6373) );
  NAND U6574 ( .A(n6374), .B(n6373), .Z(n6413) );
  NAND U6575 ( .A(b[0]), .B(a[154]), .Z(n6375) );
  XNOR U6576 ( .A(b[1]), .B(n6375), .Z(n6377) );
  NAND U6577 ( .A(n37), .B(a[153]), .Z(n6376) );
  AND U6578 ( .A(n6377), .B(n6376), .Z(n6430) );
  XOR U6579 ( .A(a[150]), .B(n42197), .Z(n6419) );
  NANDN U6580 ( .A(n6419), .B(n42173), .Z(n6380) );
  NANDN U6581 ( .A(n6378), .B(n42172), .Z(n6379) );
  NAND U6582 ( .A(n6380), .B(n6379), .Z(n6428) );
  NAND U6583 ( .A(b[7]), .B(a[146]), .Z(n6429) );
  XNOR U6584 ( .A(n6428), .B(n6429), .Z(n6431) );
  XOR U6585 ( .A(n6430), .B(n6431), .Z(n6437) );
  NANDN U6586 ( .A(n6381), .B(n42093), .Z(n6383) );
  XOR U6587 ( .A(n42134), .B(a[152]), .Z(n6422) );
  NANDN U6588 ( .A(n6422), .B(n42095), .Z(n6382) );
  NAND U6589 ( .A(n6383), .B(n6382), .Z(n6435) );
  NANDN U6590 ( .A(n6384), .B(n42231), .Z(n6386) );
  XOR U6591 ( .A(n174), .B(a[148]), .Z(n6425) );
  NANDN U6592 ( .A(n6425), .B(n42234), .Z(n6385) );
  AND U6593 ( .A(n6386), .B(n6385), .Z(n6434) );
  XNOR U6594 ( .A(n6435), .B(n6434), .Z(n6436) );
  XNOR U6595 ( .A(n6437), .B(n6436), .Z(n6441) );
  NANDN U6596 ( .A(n6388), .B(n6387), .Z(n6392) );
  NAND U6597 ( .A(n6390), .B(n6389), .Z(n6391) );
  AND U6598 ( .A(n6392), .B(n6391), .Z(n6440) );
  XOR U6599 ( .A(n6441), .B(n6440), .Z(n6442) );
  NANDN U6600 ( .A(n6394), .B(n6393), .Z(n6398) );
  NANDN U6601 ( .A(n6396), .B(n6395), .Z(n6397) );
  NAND U6602 ( .A(n6398), .B(n6397), .Z(n6443) );
  XOR U6603 ( .A(n6442), .B(n6443), .Z(n6410) );
  OR U6604 ( .A(n6400), .B(n6399), .Z(n6404) );
  NANDN U6605 ( .A(n6402), .B(n6401), .Z(n6403) );
  NAND U6606 ( .A(n6404), .B(n6403), .Z(n6411) );
  XNOR U6607 ( .A(n6410), .B(n6411), .Z(n6412) );
  XNOR U6608 ( .A(n6413), .B(n6412), .Z(n6446) );
  XNOR U6609 ( .A(n6446), .B(sreg[1170]), .Z(n6448) );
  NAND U6610 ( .A(n6405), .B(sreg[1169]), .Z(n6409) );
  OR U6611 ( .A(n6407), .B(n6406), .Z(n6408) );
  AND U6612 ( .A(n6409), .B(n6408), .Z(n6447) );
  XOR U6613 ( .A(n6448), .B(n6447), .Z(c[1170]) );
  NANDN U6614 ( .A(n6411), .B(n6410), .Z(n6415) );
  NAND U6615 ( .A(n6413), .B(n6412), .Z(n6414) );
  NAND U6616 ( .A(n6415), .B(n6414), .Z(n6454) );
  NAND U6617 ( .A(b[0]), .B(a[155]), .Z(n6416) );
  XNOR U6618 ( .A(b[1]), .B(n6416), .Z(n6418) );
  NAND U6619 ( .A(n37), .B(a[154]), .Z(n6417) );
  AND U6620 ( .A(n6418), .B(n6417), .Z(n6471) );
  XOR U6621 ( .A(a[151]), .B(n42197), .Z(n6460) );
  NANDN U6622 ( .A(n6460), .B(n42173), .Z(n6421) );
  NANDN U6623 ( .A(n6419), .B(n42172), .Z(n6420) );
  NAND U6624 ( .A(n6421), .B(n6420), .Z(n6469) );
  NAND U6625 ( .A(b[7]), .B(a[147]), .Z(n6470) );
  XNOR U6626 ( .A(n6469), .B(n6470), .Z(n6472) );
  XOR U6627 ( .A(n6471), .B(n6472), .Z(n6478) );
  NANDN U6628 ( .A(n6422), .B(n42093), .Z(n6424) );
  XOR U6629 ( .A(n42134), .B(a[153]), .Z(n6463) );
  NANDN U6630 ( .A(n6463), .B(n42095), .Z(n6423) );
  NAND U6631 ( .A(n6424), .B(n6423), .Z(n6476) );
  NANDN U6632 ( .A(n6425), .B(n42231), .Z(n6427) );
  XOR U6633 ( .A(n174), .B(a[149]), .Z(n6466) );
  NANDN U6634 ( .A(n6466), .B(n42234), .Z(n6426) );
  AND U6635 ( .A(n6427), .B(n6426), .Z(n6475) );
  XNOR U6636 ( .A(n6476), .B(n6475), .Z(n6477) );
  XNOR U6637 ( .A(n6478), .B(n6477), .Z(n6482) );
  NANDN U6638 ( .A(n6429), .B(n6428), .Z(n6433) );
  NAND U6639 ( .A(n6431), .B(n6430), .Z(n6432) );
  AND U6640 ( .A(n6433), .B(n6432), .Z(n6481) );
  XOR U6641 ( .A(n6482), .B(n6481), .Z(n6483) );
  NANDN U6642 ( .A(n6435), .B(n6434), .Z(n6439) );
  NANDN U6643 ( .A(n6437), .B(n6436), .Z(n6438) );
  NAND U6644 ( .A(n6439), .B(n6438), .Z(n6484) );
  XOR U6645 ( .A(n6483), .B(n6484), .Z(n6451) );
  OR U6646 ( .A(n6441), .B(n6440), .Z(n6445) );
  NANDN U6647 ( .A(n6443), .B(n6442), .Z(n6444) );
  NAND U6648 ( .A(n6445), .B(n6444), .Z(n6452) );
  XNOR U6649 ( .A(n6451), .B(n6452), .Z(n6453) );
  XNOR U6650 ( .A(n6454), .B(n6453), .Z(n6487) );
  XNOR U6651 ( .A(n6487), .B(sreg[1171]), .Z(n6489) );
  NAND U6652 ( .A(n6446), .B(sreg[1170]), .Z(n6450) );
  OR U6653 ( .A(n6448), .B(n6447), .Z(n6449) );
  AND U6654 ( .A(n6450), .B(n6449), .Z(n6488) );
  XOR U6655 ( .A(n6489), .B(n6488), .Z(c[1171]) );
  NANDN U6656 ( .A(n6452), .B(n6451), .Z(n6456) );
  NAND U6657 ( .A(n6454), .B(n6453), .Z(n6455) );
  NAND U6658 ( .A(n6456), .B(n6455), .Z(n6495) );
  NAND U6659 ( .A(b[0]), .B(a[156]), .Z(n6457) );
  XNOR U6660 ( .A(b[1]), .B(n6457), .Z(n6459) );
  NAND U6661 ( .A(n37), .B(a[155]), .Z(n6458) );
  AND U6662 ( .A(n6459), .B(n6458), .Z(n6512) );
  XOR U6663 ( .A(a[152]), .B(n42197), .Z(n6501) );
  NANDN U6664 ( .A(n6501), .B(n42173), .Z(n6462) );
  NANDN U6665 ( .A(n6460), .B(n42172), .Z(n6461) );
  NAND U6666 ( .A(n6462), .B(n6461), .Z(n6510) );
  NAND U6667 ( .A(b[7]), .B(a[148]), .Z(n6511) );
  XNOR U6668 ( .A(n6510), .B(n6511), .Z(n6513) );
  XOR U6669 ( .A(n6512), .B(n6513), .Z(n6519) );
  NANDN U6670 ( .A(n6463), .B(n42093), .Z(n6465) );
  XOR U6671 ( .A(n42134), .B(a[154]), .Z(n6504) );
  NANDN U6672 ( .A(n6504), .B(n42095), .Z(n6464) );
  NAND U6673 ( .A(n6465), .B(n6464), .Z(n6517) );
  NANDN U6674 ( .A(n6466), .B(n42231), .Z(n6468) );
  XOR U6675 ( .A(n174), .B(a[150]), .Z(n6507) );
  NANDN U6676 ( .A(n6507), .B(n42234), .Z(n6467) );
  AND U6677 ( .A(n6468), .B(n6467), .Z(n6516) );
  XNOR U6678 ( .A(n6517), .B(n6516), .Z(n6518) );
  XNOR U6679 ( .A(n6519), .B(n6518), .Z(n6523) );
  NANDN U6680 ( .A(n6470), .B(n6469), .Z(n6474) );
  NAND U6681 ( .A(n6472), .B(n6471), .Z(n6473) );
  AND U6682 ( .A(n6474), .B(n6473), .Z(n6522) );
  XOR U6683 ( .A(n6523), .B(n6522), .Z(n6524) );
  NANDN U6684 ( .A(n6476), .B(n6475), .Z(n6480) );
  NANDN U6685 ( .A(n6478), .B(n6477), .Z(n6479) );
  NAND U6686 ( .A(n6480), .B(n6479), .Z(n6525) );
  XOR U6687 ( .A(n6524), .B(n6525), .Z(n6492) );
  OR U6688 ( .A(n6482), .B(n6481), .Z(n6486) );
  NANDN U6689 ( .A(n6484), .B(n6483), .Z(n6485) );
  NAND U6690 ( .A(n6486), .B(n6485), .Z(n6493) );
  XNOR U6691 ( .A(n6492), .B(n6493), .Z(n6494) );
  XNOR U6692 ( .A(n6495), .B(n6494), .Z(n6528) );
  XNOR U6693 ( .A(n6528), .B(sreg[1172]), .Z(n6530) );
  NAND U6694 ( .A(n6487), .B(sreg[1171]), .Z(n6491) );
  OR U6695 ( .A(n6489), .B(n6488), .Z(n6490) );
  AND U6696 ( .A(n6491), .B(n6490), .Z(n6529) );
  XOR U6697 ( .A(n6530), .B(n6529), .Z(c[1172]) );
  NANDN U6698 ( .A(n6493), .B(n6492), .Z(n6497) );
  NAND U6699 ( .A(n6495), .B(n6494), .Z(n6496) );
  NAND U6700 ( .A(n6497), .B(n6496), .Z(n6536) );
  NAND U6701 ( .A(b[0]), .B(a[157]), .Z(n6498) );
  XNOR U6702 ( .A(b[1]), .B(n6498), .Z(n6500) );
  NAND U6703 ( .A(n37), .B(a[156]), .Z(n6499) );
  AND U6704 ( .A(n6500), .B(n6499), .Z(n6553) );
  XOR U6705 ( .A(a[153]), .B(n42197), .Z(n6542) );
  NANDN U6706 ( .A(n6542), .B(n42173), .Z(n6503) );
  NANDN U6707 ( .A(n6501), .B(n42172), .Z(n6502) );
  NAND U6708 ( .A(n6503), .B(n6502), .Z(n6551) );
  NAND U6709 ( .A(b[7]), .B(a[149]), .Z(n6552) );
  XNOR U6710 ( .A(n6551), .B(n6552), .Z(n6554) );
  XOR U6711 ( .A(n6553), .B(n6554), .Z(n6560) );
  NANDN U6712 ( .A(n6504), .B(n42093), .Z(n6506) );
  XOR U6713 ( .A(n42134), .B(a[155]), .Z(n6545) );
  NANDN U6714 ( .A(n6545), .B(n42095), .Z(n6505) );
  NAND U6715 ( .A(n6506), .B(n6505), .Z(n6558) );
  NANDN U6716 ( .A(n6507), .B(n42231), .Z(n6509) );
  XOR U6717 ( .A(n174), .B(a[151]), .Z(n6548) );
  NANDN U6718 ( .A(n6548), .B(n42234), .Z(n6508) );
  AND U6719 ( .A(n6509), .B(n6508), .Z(n6557) );
  XNOR U6720 ( .A(n6558), .B(n6557), .Z(n6559) );
  XNOR U6721 ( .A(n6560), .B(n6559), .Z(n6564) );
  NANDN U6722 ( .A(n6511), .B(n6510), .Z(n6515) );
  NAND U6723 ( .A(n6513), .B(n6512), .Z(n6514) );
  AND U6724 ( .A(n6515), .B(n6514), .Z(n6563) );
  XOR U6725 ( .A(n6564), .B(n6563), .Z(n6565) );
  NANDN U6726 ( .A(n6517), .B(n6516), .Z(n6521) );
  NANDN U6727 ( .A(n6519), .B(n6518), .Z(n6520) );
  NAND U6728 ( .A(n6521), .B(n6520), .Z(n6566) );
  XOR U6729 ( .A(n6565), .B(n6566), .Z(n6533) );
  OR U6730 ( .A(n6523), .B(n6522), .Z(n6527) );
  NANDN U6731 ( .A(n6525), .B(n6524), .Z(n6526) );
  NAND U6732 ( .A(n6527), .B(n6526), .Z(n6534) );
  XNOR U6733 ( .A(n6533), .B(n6534), .Z(n6535) );
  XNOR U6734 ( .A(n6536), .B(n6535), .Z(n6569) );
  XNOR U6735 ( .A(n6569), .B(sreg[1173]), .Z(n6571) );
  NAND U6736 ( .A(n6528), .B(sreg[1172]), .Z(n6532) );
  OR U6737 ( .A(n6530), .B(n6529), .Z(n6531) );
  AND U6738 ( .A(n6532), .B(n6531), .Z(n6570) );
  XOR U6739 ( .A(n6571), .B(n6570), .Z(c[1173]) );
  NANDN U6740 ( .A(n6534), .B(n6533), .Z(n6538) );
  NAND U6741 ( .A(n6536), .B(n6535), .Z(n6537) );
  NAND U6742 ( .A(n6538), .B(n6537), .Z(n6577) );
  NAND U6743 ( .A(b[0]), .B(a[158]), .Z(n6539) );
  XNOR U6744 ( .A(b[1]), .B(n6539), .Z(n6541) );
  NAND U6745 ( .A(n37), .B(a[157]), .Z(n6540) );
  AND U6746 ( .A(n6541), .B(n6540), .Z(n6594) );
  XOR U6747 ( .A(a[154]), .B(n42197), .Z(n6583) );
  NANDN U6748 ( .A(n6583), .B(n42173), .Z(n6544) );
  NANDN U6749 ( .A(n6542), .B(n42172), .Z(n6543) );
  NAND U6750 ( .A(n6544), .B(n6543), .Z(n6592) );
  NAND U6751 ( .A(b[7]), .B(a[150]), .Z(n6593) );
  XNOR U6752 ( .A(n6592), .B(n6593), .Z(n6595) );
  XOR U6753 ( .A(n6594), .B(n6595), .Z(n6601) );
  NANDN U6754 ( .A(n6545), .B(n42093), .Z(n6547) );
  XOR U6755 ( .A(n42134), .B(a[156]), .Z(n6586) );
  NANDN U6756 ( .A(n6586), .B(n42095), .Z(n6546) );
  NAND U6757 ( .A(n6547), .B(n6546), .Z(n6599) );
  NANDN U6758 ( .A(n6548), .B(n42231), .Z(n6550) );
  XOR U6759 ( .A(n174), .B(a[152]), .Z(n6589) );
  NANDN U6760 ( .A(n6589), .B(n42234), .Z(n6549) );
  AND U6761 ( .A(n6550), .B(n6549), .Z(n6598) );
  XNOR U6762 ( .A(n6599), .B(n6598), .Z(n6600) );
  XNOR U6763 ( .A(n6601), .B(n6600), .Z(n6605) );
  NANDN U6764 ( .A(n6552), .B(n6551), .Z(n6556) );
  NAND U6765 ( .A(n6554), .B(n6553), .Z(n6555) );
  AND U6766 ( .A(n6556), .B(n6555), .Z(n6604) );
  XOR U6767 ( .A(n6605), .B(n6604), .Z(n6606) );
  NANDN U6768 ( .A(n6558), .B(n6557), .Z(n6562) );
  NANDN U6769 ( .A(n6560), .B(n6559), .Z(n6561) );
  NAND U6770 ( .A(n6562), .B(n6561), .Z(n6607) );
  XOR U6771 ( .A(n6606), .B(n6607), .Z(n6574) );
  OR U6772 ( .A(n6564), .B(n6563), .Z(n6568) );
  NANDN U6773 ( .A(n6566), .B(n6565), .Z(n6567) );
  NAND U6774 ( .A(n6568), .B(n6567), .Z(n6575) );
  XNOR U6775 ( .A(n6574), .B(n6575), .Z(n6576) );
  XNOR U6776 ( .A(n6577), .B(n6576), .Z(n6610) );
  XNOR U6777 ( .A(n6610), .B(sreg[1174]), .Z(n6612) );
  NAND U6778 ( .A(n6569), .B(sreg[1173]), .Z(n6573) );
  OR U6779 ( .A(n6571), .B(n6570), .Z(n6572) );
  AND U6780 ( .A(n6573), .B(n6572), .Z(n6611) );
  XOR U6781 ( .A(n6612), .B(n6611), .Z(c[1174]) );
  NANDN U6782 ( .A(n6575), .B(n6574), .Z(n6579) );
  NAND U6783 ( .A(n6577), .B(n6576), .Z(n6578) );
  NAND U6784 ( .A(n6579), .B(n6578), .Z(n6618) );
  NAND U6785 ( .A(b[0]), .B(a[159]), .Z(n6580) );
  XNOR U6786 ( .A(b[1]), .B(n6580), .Z(n6582) );
  NAND U6787 ( .A(n37), .B(a[158]), .Z(n6581) );
  AND U6788 ( .A(n6582), .B(n6581), .Z(n6635) );
  XOR U6789 ( .A(a[155]), .B(n42197), .Z(n6624) );
  NANDN U6790 ( .A(n6624), .B(n42173), .Z(n6585) );
  NANDN U6791 ( .A(n6583), .B(n42172), .Z(n6584) );
  NAND U6792 ( .A(n6585), .B(n6584), .Z(n6633) );
  NAND U6793 ( .A(b[7]), .B(a[151]), .Z(n6634) );
  XNOR U6794 ( .A(n6633), .B(n6634), .Z(n6636) );
  XOR U6795 ( .A(n6635), .B(n6636), .Z(n6642) );
  NANDN U6796 ( .A(n6586), .B(n42093), .Z(n6588) );
  XOR U6797 ( .A(n42134), .B(a[157]), .Z(n6627) );
  NANDN U6798 ( .A(n6627), .B(n42095), .Z(n6587) );
  NAND U6799 ( .A(n6588), .B(n6587), .Z(n6640) );
  NANDN U6800 ( .A(n6589), .B(n42231), .Z(n6591) );
  XOR U6801 ( .A(n174), .B(a[153]), .Z(n6630) );
  NANDN U6802 ( .A(n6630), .B(n42234), .Z(n6590) );
  AND U6803 ( .A(n6591), .B(n6590), .Z(n6639) );
  XNOR U6804 ( .A(n6640), .B(n6639), .Z(n6641) );
  XNOR U6805 ( .A(n6642), .B(n6641), .Z(n6646) );
  NANDN U6806 ( .A(n6593), .B(n6592), .Z(n6597) );
  NAND U6807 ( .A(n6595), .B(n6594), .Z(n6596) );
  AND U6808 ( .A(n6597), .B(n6596), .Z(n6645) );
  XOR U6809 ( .A(n6646), .B(n6645), .Z(n6647) );
  NANDN U6810 ( .A(n6599), .B(n6598), .Z(n6603) );
  NANDN U6811 ( .A(n6601), .B(n6600), .Z(n6602) );
  NAND U6812 ( .A(n6603), .B(n6602), .Z(n6648) );
  XOR U6813 ( .A(n6647), .B(n6648), .Z(n6615) );
  OR U6814 ( .A(n6605), .B(n6604), .Z(n6609) );
  NANDN U6815 ( .A(n6607), .B(n6606), .Z(n6608) );
  NAND U6816 ( .A(n6609), .B(n6608), .Z(n6616) );
  XNOR U6817 ( .A(n6615), .B(n6616), .Z(n6617) );
  XNOR U6818 ( .A(n6618), .B(n6617), .Z(n6651) );
  XNOR U6819 ( .A(n6651), .B(sreg[1175]), .Z(n6653) );
  NAND U6820 ( .A(n6610), .B(sreg[1174]), .Z(n6614) );
  OR U6821 ( .A(n6612), .B(n6611), .Z(n6613) );
  AND U6822 ( .A(n6614), .B(n6613), .Z(n6652) );
  XOR U6823 ( .A(n6653), .B(n6652), .Z(c[1175]) );
  NANDN U6824 ( .A(n6616), .B(n6615), .Z(n6620) );
  NAND U6825 ( .A(n6618), .B(n6617), .Z(n6619) );
  NAND U6826 ( .A(n6620), .B(n6619), .Z(n6659) );
  NAND U6827 ( .A(b[0]), .B(a[160]), .Z(n6621) );
  XNOR U6828 ( .A(b[1]), .B(n6621), .Z(n6623) );
  NAND U6829 ( .A(n37), .B(a[159]), .Z(n6622) );
  AND U6830 ( .A(n6623), .B(n6622), .Z(n6676) );
  XOR U6831 ( .A(a[156]), .B(n42197), .Z(n6665) );
  NANDN U6832 ( .A(n6665), .B(n42173), .Z(n6626) );
  NANDN U6833 ( .A(n6624), .B(n42172), .Z(n6625) );
  NAND U6834 ( .A(n6626), .B(n6625), .Z(n6674) );
  NAND U6835 ( .A(b[7]), .B(a[152]), .Z(n6675) );
  XNOR U6836 ( .A(n6674), .B(n6675), .Z(n6677) );
  XOR U6837 ( .A(n6676), .B(n6677), .Z(n6683) );
  NANDN U6838 ( .A(n6627), .B(n42093), .Z(n6629) );
  XOR U6839 ( .A(n42134), .B(a[158]), .Z(n6668) );
  NANDN U6840 ( .A(n6668), .B(n42095), .Z(n6628) );
  NAND U6841 ( .A(n6629), .B(n6628), .Z(n6681) );
  NANDN U6842 ( .A(n6630), .B(n42231), .Z(n6632) );
  XOR U6843 ( .A(n174), .B(a[154]), .Z(n6671) );
  NANDN U6844 ( .A(n6671), .B(n42234), .Z(n6631) );
  AND U6845 ( .A(n6632), .B(n6631), .Z(n6680) );
  XNOR U6846 ( .A(n6681), .B(n6680), .Z(n6682) );
  XNOR U6847 ( .A(n6683), .B(n6682), .Z(n6687) );
  NANDN U6848 ( .A(n6634), .B(n6633), .Z(n6638) );
  NAND U6849 ( .A(n6636), .B(n6635), .Z(n6637) );
  AND U6850 ( .A(n6638), .B(n6637), .Z(n6686) );
  XOR U6851 ( .A(n6687), .B(n6686), .Z(n6688) );
  NANDN U6852 ( .A(n6640), .B(n6639), .Z(n6644) );
  NANDN U6853 ( .A(n6642), .B(n6641), .Z(n6643) );
  NAND U6854 ( .A(n6644), .B(n6643), .Z(n6689) );
  XOR U6855 ( .A(n6688), .B(n6689), .Z(n6656) );
  OR U6856 ( .A(n6646), .B(n6645), .Z(n6650) );
  NANDN U6857 ( .A(n6648), .B(n6647), .Z(n6649) );
  NAND U6858 ( .A(n6650), .B(n6649), .Z(n6657) );
  XNOR U6859 ( .A(n6656), .B(n6657), .Z(n6658) );
  XNOR U6860 ( .A(n6659), .B(n6658), .Z(n6692) );
  XNOR U6861 ( .A(n6692), .B(sreg[1176]), .Z(n6694) );
  NAND U6862 ( .A(n6651), .B(sreg[1175]), .Z(n6655) );
  OR U6863 ( .A(n6653), .B(n6652), .Z(n6654) );
  AND U6864 ( .A(n6655), .B(n6654), .Z(n6693) );
  XOR U6865 ( .A(n6694), .B(n6693), .Z(c[1176]) );
  NANDN U6866 ( .A(n6657), .B(n6656), .Z(n6661) );
  NAND U6867 ( .A(n6659), .B(n6658), .Z(n6660) );
  NAND U6868 ( .A(n6661), .B(n6660), .Z(n6700) );
  NAND U6869 ( .A(b[0]), .B(a[161]), .Z(n6662) );
  XNOR U6870 ( .A(b[1]), .B(n6662), .Z(n6664) );
  NAND U6871 ( .A(n38), .B(a[160]), .Z(n6663) );
  AND U6872 ( .A(n6664), .B(n6663), .Z(n6717) );
  XOR U6873 ( .A(a[157]), .B(n42197), .Z(n6706) );
  NANDN U6874 ( .A(n6706), .B(n42173), .Z(n6667) );
  NANDN U6875 ( .A(n6665), .B(n42172), .Z(n6666) );
  NAND U6876 ( .A(n6667), .B(n6666), .Z(n6715) );
  NAND U6877 ( .A(b[7]), .B(a[153]), .Z(n6716) );
  XNOR U6878 ( .A(n6715), .B(n6716), .Z(n6718) );
  XOR U6879 ( .A(n6717), .B(n6718), .Z(n6724) );
  NANDN U6880 ( .A(n6668), .B(n42093), .Z(n6670) );
  XOR U6881 ( .A(n42134), .B(a[159]), .Z(n6709) );
  NANDN U6882 ( .A(n6709), .B(n42095), .Z(n6669) );
  NAND U6883 ( .A(n6670), .B(n6669), .Z(n6722) );
  NANDN U6884 ( .A(n6671), .B(n42231), .Z(n6673) );
  XOR U6885 ( .A(n175), .B(a[155]), .Z(n6712) );
  NANDN U6886 ( .A(n6712), .B(n42234), .Z(n6672) );
  AND U6887 ( .A(n6673), .B(n6672), .Z(n6721) );
  XNOR U6888 ( .A(n6722), .B(n6721), .Z(n6723) );
  XNOR U6889 ( .A(n6724), .B(n6723), .Z(n6728) );
  NANDN U6890 ( .A(n6675), .B(n6674), .Z(n6679) );
  NAND U6891 ( .A(n6677), .B(n6676), .Z(n6678) );
  AND U6892 ( .A(n6679), .B(n6678), .Z(n6727) );
  XOR U6893 ( .A(n6728), .B(n6727), .Z(n6729) );
  NANDN U6894 ( .A(n6681), .B(n6680), .Z(n6685) );
  NANDN U6895 ( .A(n6683), .B(n6682), .Z(n6684) );
  NAND U6896 ( .A(n6685), .B(n6684), .Z(n6730) );
  XOR U6897 ( .A(n6729), .B(n6730), .Z(n6697) );
  OR U6898 ( .A(n6687), .B(n6686), .Z(n6691) );
  NANDN U6899 ( .A(n6689), .B(n6688), .Z(n6690) );
  NAND U6900 ( .A(n6691), .B(n6690), .Z(n6698) );
  XNOR U6901 ( .A(n6697), .B(n6698), .Z(n6699) );
  XNOR U6902 ( .A(n6700), .B(n6699), .Z(n6733) );
  XNOR U6903 ( .A(n6733), .B(sreg[1177]), .Z(n6735) );
  NAND U6904 ( .A(n6692), .B(sreg[1176]), .Z(n6696) );
  OR U6905 ( .A(n6694), .B(n6693), .Z(n6695) );
  AND U6906 ( .A(n6696), .B(n6695), .Z(n6734) );
  XOR U6907 ( .A(n6735), .B(n6734), .Z(c[1177]) );
  NANDN U6908 ( .A(n6698), .B(n6697), .Z(n6702) );
  NAND U6909 ( .A(n6700), .B(n6699), .Z(n6701) );
  NAND U6910 ( .A(n6702), .B(n6701), .Z(n6741) );
  NAND U6911 ( .A(b[0]), .B(a[162]), .Z(n6703) );
  XNOR U6912 ( .A(b[1]), .B(n6703), .Z(n6705) );
  NAND U6913 ( .A(n38), .B(a[161]), .Z(n6704) );
  AND U6914 ( .A(n6705), .B(n6704), .Z(n6758) );
  XOR U6915 ( .A(a[158]), .B(n42197), .Z(n6747) );
  NANDN U6916 ( .A(n6747), .B(n42173), .Z(n6708) );
  NANDN U6917 ( .A(n6706), .B(n42172), .Z(n6707) );
  NAND U6918 ( .A(n6708), .B(n6707), .Z(n6756) );
  NAND U6919 ( .A(b[7]), .B(a[154]), .Z(n6757) );
  XNOR U6920 ( .A(n6756), .B(n6757), .Z(n6759) );
  XOR U6921 ( .A(n6758), .B(n6759), .Z(n6765) );
  NANDN U6922 ( .A(n6709), .B(n42093), .Z(n6711) );
  XOR U6923 ( .A(n42134), .B(a[160]), .Z(n6750) );
  NANDN U6924 ( .A(n6750), .B(n42095), .Z(n6710) );
  NAND U6925 ( .A(n6711), .B(n6710), .Z(n6763) );
  NANDN U6926 ( .A(n6712), .B(n42231), .Z(n6714) );
  XOR U6927 ( .A(n175), .B(a[156]), .Z(n6753) );
  NANDN U6928 ( .A(n6753), .B(n42234), .Z(n6713) );
  AND U6929 ( .A(n6714), .B(n6713), .Z(n6762) );
  XNOR U6930 ( .A(n6763), .B(n6762), .Z(n6764) );
  XNOR U6931 ( .A(n6765), .B(n6764), .Z(n6769) );
  NANDN U6932 ( .A(n6716), .B(n6715), .Z(n6720) );
  NAND U6933 ( .A(n6718), .B(n6717), .Z(n6719) );
  AND U6934 ( .A(n6720), .B(n6719), .Z(n6768) );
  XOR U6935 ( .A(n6769), .B(n6768), .Z(n6770) );
  NANDN U6936 ( .A(n6722), .B(n6721), .Z(n6726) );
  NANDN U6937 ( .A(n6724), .B(n6723), .Z(n6725) );
  NAND U6938 ( .A(n6726), .B(n6725), .Z(n6771) );
  XOR U6939 ( .A(n6770), .B(n6771), .Z(n6738) );
  OR U6940 ( .A(n6728), .B(n6727), .Z(n6732) );
  NANDN U6941 ( .A(n6730), .B(n6729), .Z(n6731) );
  NAND U6942 ( .A(n6732), .B(n6731), .Z(n6739) );
  XNOR U6943 ( .A(n6738), .B(n6739), .Z(n6740) );
  XNOR U6944 ( .A(n6741), .B(n6740), .Z(n6774) );
  XNOR U6945 ( .A(n6774), .B(sreg[1178]), .Z(n6776) );
  NAND U6946 ( .A(n6733), .B(sreg[1177]), .Z(n6737) );
  OR U6947 ( .A(n6735), .B(n6734), .Z(n6736) );
  AND U6948 ( .A(n6737), .B(n6736), .Z(n6775) );
  XOR U6949 ( .A(n6776), .B(n6775), .Z(c[1178]) );
  NANDN U6950 ( .A(n6739), .B(n6738), .Z(n6743) );
  NAND U6951 ( .A(n6741), .B(n6740), .Z(n6742) );
  NAND U6952 ( .A(n6743), .B(n6742), .Z(n6782) );
  NAND U6953 ( .A(b[0]), .B(a[163]), .Z(n6744) );
  XNOR U6954 ( .A(b[1]), .B(n6744), .Z(n6746) );
  NAND U6955 ( .A(n38), .B(a[162]), .Z(n6745) );
  AND U6956 ( .A(n6746), .B(n6745), .Z(n6799) );
  XOR U6957 ( .A(a[159]), .B(n42197), .Z(n6788) );
  NANDN U6958 ( .A(n6788), .B(n42173), .Z(n6749) );
  NANDN U6959 ( .A(n6747), .B(n42172), .Z(n6748) );
  NAND U6960 ( .A(n6749), .B(n6748), .Z(n6797) );
  NAND U6961 ( .A(b[7]), .B(a[155]), .Z(n6798) );
  XNOR U6962 ( .A(n6797), .B(n6798), .Z(n6800) );
  XOR U6963 ( .A(n6799), .B(n6800), .Z(n6806) );
  NANDN U6964 ( .A(n6750), .B(n42093), .Z(n6752) );
  XOR U6965 ( .A(n42134), .B(a[161]), .Z(n6791) );
  NANDN U6966 ( .A(n6791), .B(n42095), .Z(n6751) );
  NAND U6967 ( .A(n6752), .B(n6751), .Z(n6804) );
  NANDN U6968 ( .A(n6753), .B(n42231), .Z(n6755) );
  XOR U6969 ( .A(n175), .B(a[157]), .Z(n6794) );
  NANDN U6970 ( .A(n6794), .B(n42234), .Z(n6754) );
  AND U6971 ( .A(n6755), .B(n6754), .Z(n6803) );
  XNOR U6972 ( .A(n6804), .B(n6803), .Z(n6805) );
  XNOR U6973 ( .A(n6806), .B(n6805), .Z(n6810) );
  NANDN U6974 ( .A(n6757), .B(n6756), .Z(n6761) );
  NAND U6975 ( .A(n6759), .B(n6758), .Z(n6760) );
  AND U6976 ( .A(n6761), .B(n6760), .Z(n6809) );
  XOR U6977 ( .A(n6810), .B(n6809), .Z(n6811) );
  NANDN U6978 ( .A(n6763), .B(n6762), .Z(n6767) );
  NANDN U6979 ( .A(n6765), .B(n6764), .Z(n6766) );
  NAND U6980 ( .A(n6767), .B(n6766), .Z(n6812) );
  XOR U6981 ( .A(n6811), .B(n6812), .Z(n6779) );
  OR U6982 ( .A(n6769), .B(n6768), .Z(n6773) );
  NANDN U6983 ( .A(n6771), .B(n6770), .Z(n6772) );
  NAND U6984 ( .A(n6773), .B(n6772), .Z(n6780) );
  XNOR U6985 ( .A(n6779), .B(n6780), .Z(n6781) );
  XNOR U6986 ( .A(n6782), .B(n6781), .Z(n6815) );
  XNOR U6987 ( .A(n6815), .B(sreg[1179]), .Z(n6817) );
  NAND U6988 ( .A(n6774), .B(sreg[1178]), .Z(n6778) );
  OR U6989 ( .A(n6776), .B(n6775), .Z(n6777) );
  AND U6990 ( .A(n6778), .B(n6777), .Z(n6816) );
  XOR U6991 ( .A(n6817), .B(n6816), .Z(c[1179]) );
  NANDN U6992 ( .A(n6780), .B(n6779), .Z(n6784) );
  NAND U6993 ( .A(n6782), .B(n6781), .Z(n6783) );
  NAND U6994 ( .A(n6784), .B(n6783), .Z(n6823) );
  NAND U6995 ( .A(b[0]), .B(a[164]), .Z(n6785) );
  XNOR U6996 ( .A(b[1]), .B(n6785), .Z(n6787) );
  NAND U6997 ( .A(n38), .B(a[163]), .Z(n6786) );
  AND U6998 ( .A(n6787), .B(n6786), .Z(n6840) );
  XOR U6999 ( .A(a[160]), .B(n42197), .Z(n6829) );
  NANDN U7000 ( .A(n6829), .B(n42173), .Z(n6790) );
  NANDN U7001 ( .A(n6788), .B(n42172), .Z(n6789) );
  NAND U7002 ( .A(n6790), .B(n6789), .Z(n6838) );
  NAND U7003 ( .A(b[7]), .B(a[156]), .Z(n6839) );
  XNOR U7004 ( .A(n6838), .B(n6839), .Z(n6841) );
  XOR U7005 ( .A(n6840), .B(n6841), .Z(n6847) );
  NANDN U7006 ( .A(n6791), .B(n42093), .Z(n6793) );
  XOR U7007 ( .A(n42134), .B(a[162]), .Z(n6832) );
  NANDN U7008 ( .A(n6832), .B(n42095), .Z(n6792) );
  NAND U7009 ( .A(n6793), .B(n6792), .Z(n6845) );
  NANDN U7010 ( .A(n6794), .B(n42231), .Z(n6796) );
  XOR U7011 ( .A(n175), .B(a[158]), .Z(n6835) );
  NANDN U7012 ( .A(n6835), .B(n42234), .Z(n6795) );
  AND U7013 ( .A(n6796), .B(n6795), .Z(n6844) );
  XNOR U7014 ( .A(n6845), .B(n6844), .Z(n6846) );
  XNOR U7015 ( .A(n6847), .B(n6846), .Z(n6851) );
  NANDN U7016 ( .A(n6798), .B(n6797), .Z(n6802) );
  NAND U7017 ( .A(n6800), .B(n6799), .Z(n6801) );
  AND U7018 ( .A(n6802), .B(n6801), .Z(n6850) );
  XOR U7019 ( .A(n6851), .B(n6850), .Z(n6852) );
  NANDN U7020 ( .A(n6804), .B(n6803), .Z(n6808) );
  NANDN U7021 ( .A(n6806), .B(n6805), .Z(n6807) );
  NAND U7022 ( .A(n6808), .B(n6807), .Z(n6853) );
  XOR U7023 ( .A(n6852), .B(n6853), .Z(n6820) );
  OR U7024 ( .A(n6810), .B(n6809), .Z(n6814) );
  NANDN U7025 ( .A(n6812), .B(n6811), .Z(n6813) );
  NAND U7026 ( .A(n6814), .B(n6813), .Z(n6821) );
  XNOR U7027 ( .A(n6820), .B(n6821), .Z(n6822) );
  XNOR U7028 ( .A(n6823), .B(n6822), .Z(n6856) );
  XNOR U7029 ( .A(n6856), .B(sreg[1180]), .Z(n6858) );
  NAND U7030 ( .A(n6815), .B(sreg[1179]), .Z(n6819) );
  OR U7031 ( .A(n6817), .B(n6816), .Z(n6818) );
  AND U7032 ( .A(n6819), .B(n6818), .Z(n6857) );
  XOR U7033 ( .A(n6858), .B(n6857), .Z(c[1180]) );
  NANDN U7034 ( .A(n6821), .B(n6820), .Z(n6825) );
  NAND U7035 ( .A(n6823), .B(n6822), .Z(n6824) );
  NAND U7036 ( .A(n6825), .B(n6824), .Z(n6864) );
  NAND U7037 ( .A(b[0]), .B(a[165]), .Z(n6826) );
  XNOR U7038 ( .A(b[1]), .B(n6826), .Z(n6828) );
  NAND U7039 ( .A(n38), .B(a[164]), .Z(n6827) );
  AND U7040 ( .A(n6828), .B(n6827), .Z(n6881) );
  XOR U7041 ( .A(a[161]), .B(n42197), .Z(n6870) );
  NANDN U7042 ( .A(n6870), .B(n42173), .Z(n6831) );
  NANDN U7043 ( .A(n6829), .B(n42172), .Z(n6830) );
  NAND U7044 ( .A(n6831), .B(n6830), .Z(n6879) );
  NAND U7045 ( .A(b[7]), .B(a[157]), .Z(n6880) );
  XNOR U7046 ( .A(n6879), .B(n6880), .Z(n6882) );
  XOR U7047 ( .A(n6881), .B(n6882), .Z(n6888) );
  NANDN U7048 ( .A(n6832), .B(n42093), .Z(n6834) );
  XOR U7049 ( .A(n42134), .B(a[163]), .Z(n6873) );
  NANDN U7050 ( .A(n6873), .B(n42095), .Z(n6833) );
  NAND U7051 ( .A(n6834), .B(n6833), .Z(n6886) );
  NANDN U7052 ( .A(n6835), .B(n42231), .Z(n6837) );
  XOR U7053 ( .A(n175), .B(a[159]), .Z(n6876) );
  NANDN U7054 ( .A(n6876), .B(n42234), .Z(n6836) );
  AND U7055 ( .A(n6837), .B(n6836), .Z(n6885) );
  XNOR U7056 ( .A(n6886), .B(n6885), .Z(n6887) );
  XNOR U7057 ( .A(n6888), .B(n6887), .Z(n6892) );
  NANDN U7058 ( .A(n6839), .B(n6838), .Z(n6843) );
  NAND U7059 ( .A(n6841), .B(n6840), .Z(n6842) );
  AND U7060 ( .A(n6843), .B(n6842), .Z(n6891) );
  XOR U7061 ( .A(n6892), .B(n6891), .Z(n6893) );
  NANDN U7062 ( .A(n6845), .B(n6844), .Z(n6849) );
  NANDN U7063 ( .A(n6847), .B(n6846), .Z(n6848) );
  NAND U7064 ( .A(n6849), .B(n6848), .Z(n6894) );
  XOR U7065 ( .A(n6893), .B(n6894), .Z(n6861) );
  OR U7066 ( .A(n6851), .B(n6850), .Z(n6855) );
  NANDN U7067 ( .A(n6853), .B(n6852), .Z(n6854) );
  NAND U7068 ( .A(n6855), .B(n6854), .Z(n6862) );
  XNOR U7069 ( .A(n6861), .B(n6862), .Z(n6863) );
  XNOR U7070 ( .A(n6864), .B(n6863), .Z(n6897) );
  XNOR U7071 ( .A(n6897), .B(sreg[1181]), .Z(n6899) );
  NAND U7072 ( .A(n6856), .B(sreg[1180]), .Z(n6860) );
  OR U7073 ( .A(n6858), .B(n6857), .Z(n6859) );
  AND U7074 ( .A(n6860), .B(n6859), .Z(n6898) );
  XOR U7075 ( .A(n6899), .B(n6898), .Z(c[1181]) );
  NANDN U7076 ( .A(n6862), .B(n6861), .Z(n6866) );
  NAND U7077 ( .A(n6864), .B(n6863), .Z(n6865) );
  NAND U7078 ( .A(n6866), .B(n6865), .Z(n6905) );
  NAND U7079 ( .A(b[0]), .B(a[166]), .Z(n6867) );
  XNOR U7080 ( .A(b[1]), .B(n6867), .Z(n6869) );
  NAND U7081 ( .A(n38), .B(a[165]), .Z(n6868) );
  AND U7082 ( .A(n6869), .B(n6868), .Z(n6922) );
  XOR U7083 ( .A(a[162]), .B(n42197), .Z(n6911) );
  NANDN U7084 ( .A(n6911), .B(n42173), .Z(n6872) );
  NANDN U7085 ( .A(n6870), .B(n42172), .Z(n6871) );
  NAND U7086 ( .A(n6872), .B(n6871), .Z(n6920) );
  NAND U7087 ( .A(b[7]), .B(a[158]), .Z(n6921) );
  XNOR U7088 ( .A(n6920), .B(n6921), .Z(n6923) );
  XOR U7089 ( .A(n6922), .B(n6923), .Z(n6929) );
  NANDN U7090 ( .A(n6873), .B(n42093), .Z(n6875) );
  XOR U7091 ( .A(n42134), .B(a[164]), .Z(n6914) );
  NANDN U7092 ( .A(n6914), .B(n42095), .Z(n6874) );
  NAND U7093 ( .A(n6875), .B(n6874), .Z(n6927) );
  NANDN U7094 ( .A(n6876), .B(n42231), .Z(n6878) );
  XOR U7095 ( .A(n175), .B(a[160]), .Z(n6917) );
  NANDN U7096 ( .A(n6917), .B(n42234), .Z(n6877) );
  AND U7097 ( .A(n6878), .B(n6877), .Z(n6926) );
  XNOR U7098 ( .A(n6927), .B(n6926), .Z(n6928) );
  XNOR U7099 ( .A(n6929), .B(n6928), .Z(n6933) );
  NANDN U7100 ( .A(n6880), .B(n6879), .Z(n6884) );
  NAND U7101 ( .A(n6882), .B(n6881), .Z(n6883) );
  AND U7102 ( .A(n6884), .B(n6883), .Z(n6932) );
  XOR U7103 ( .A(n6933), .B(n6932), .Z(n6934) );
  NANDN U7104 ( .A(n6886), .B(n6885), .Z(n6890) );
  NANDN U7105 ( .A(n6888), .B(n6887), .Z(n6889) );
  NAND U7106 ( .A(n6890), .B(n6889), .Z(n6935) );
  XOR U7107 ( .A(n6934), .B(n6935), .Z(n6902) );
  OR U7108 ( .A(n6892), .B(n6891), .Z(n6896) );
  NANDN U7109 ( .A(n6894), .B(n6893), .Z(n6895) );
  NAND U7110 ( .A(n6896), .B(n6895), .Z(n6903) );
  XNOR U7111 ( .A(n6902), .B(n6903), .Z(n6904) );
  XNOR U7112 ( .A(n6905), .B(n6904), .Z(n6938) );
  XNOR U7113 ( .A(n6938), .B(sreg[1182]), .Z(n6940) );
  NAND U7114 ( .A(n6897), .B(sreg[1181]), .Z(n6901) );
  OR U7115 ( .A(n6899), .B(n6898), .Z(n6900) );
  AND U7116 ( .A(n6901), .B(n6900), .Z(n6939) );
  XOR U7117 ( .A(n6940), .B(n6939), .Z(c[1182]) );
  NANDN U7118 ( .A(n6903), .B(n6902), .Z(n6907) );
  NAND U7119 ( .A(n6905), .B(n6904), .Z(n6906) );
  NAND U7120 ( .A(n6907), .B(n6906), .Z(n6946) );
  NAND U7121 ( .A(b[0]), .B(a[167]), .Z(n6908) );
  XNOR U7122 ( .A(b[1]), .B(n6908), .Z(n6910) );
  NAND U7123 ( .A(n38), .B(a[166]), .Z(n6909) );
  AND U7124 ( .A(n6910), .B(n6909), .Z(n6963) );
  XOR U7125 ( .A(a[163]), .B(n42197), .Z(n6952) );
  NANDN U7126 ( .A(n6952), .B(n42173), .Z(n6913) );
  NANDN U7127 ( .A(n6911), .B(n42172), .Z(n6912) );
  NAND U7128 ( .A(n6913), .B(n6912), .Z(n6961) );
  NAND U7129 ( .A(b[7]), .B(a[159]), .Z(n6962) );
  XNOR U7130 ( .A(n6961), .B(n6962), .Z(n6964) );
  XOR U7131 ( .A(n6963), .B(n6964), .Z(n6970) );
  NANDN U7132 ( .A(n6914), .B(n42093), .Z(n6916) );
  XOR U7133 ( .A(n42134), .B(a[165]), .Z(n6955) );
  NANDN U7134 ( .A(n6955), .B(n42095), .Z(n6915) );
  NAND U7135 ( .A(n6916), .B(n6915), .Z(n6968) );
  NANDN U7136 ( .A(n6917), .B(n42231), .Z(n6919) );
  XOR U7137 ( .A(n175), .B(a[161]), .Z(n6958) );
  NANDN U7138 ( .A(n6958), .B(n42234), .Z(n6918) );
  AND U7139 ( .A(n6919), .B(n6918), .Z(n6967) );
  XNOR U7140 ( .A(n6968), .B(n6967), .Z(n6969) );
  XNOR U7141 ( .A(n6970), .B(n6969), .Z(n6974) );
  NANDN U7142 ( .A(n6921), .B(n6920), .Z(n6925) );
  NAND U7143 ( .A(n6923), .B(n6922), .Z(n6924) );
  AND U7144 ( .A(n6925), .B(n6924), .Z(n6973) );
  XOR U7145 ( .A(n6974), .B(n6973), .Z(n6975) );
  NANDN U7146 ( .A(n6927), .B(n6926), .Z(n6931) );
  NANDN U7147 ( .A(n6929), .B(n6928), .Z(n6930) );
  NAND U7148 ( .A(n6931), .B(n6930), .Z(n6976) );
  XOR U7149 ( .A(n6975), .B(n6976), .Z(n6943) );
  OR U7150 ( .A(n6933), .B(n6932), .Z(n6937) );
  NANDN U7151 ( .A(n6935), .B(n6934), .Z(n6936) );
  NAND U7152 ( .A(n6937), .B(n6936), .Z(n6944) );
  XNOR U7153 ( .A(n6943), .B(n6944), .Z(n6945) );
  XNOR U7154 ( .A(n6946), .B(n6945), .Z(n6979) );
  XNOR U7155 ( .A(n6979), .B(sreg[1183]), .Z(n6981) );
  NAND U7156 ( .A(n6938), .B(sreg[1182]), .Z(n6942) );
  OR U7157 ( .A(n6940), .B(n6939), .Z(n6941) );
  AND U7158 ( .A(n6942), .B(n6941), .Z(n6980) );
  XOR U7159 ( .A(n6981), .B(n6980), .Z(c[1183]) );
  NANDN U7160 ( .A(n6944), .B(n6943), .Z(n6948) );
  NAND U7161 ( .A(n6946), .B(n6945), .Z(n6947) );
  NAND U7162 ( .A(n6948), .B(n6947), .Z(n6987) );
  NAND U7163 ( .A(b[0]), .B(a[168]), .Z(n6949) );
  XNOR U7164 ( .A(b[1]), .B(n6949), .Z(n6951) );
  NAND U7165 ( .A(n39), .B(a[167]), .Z(n6950) );
  AND U7166 ( .A(n6951), .B(n6950), .Z(n7004) );
  XOR U7167 ( .A(a[164]), .B(n42197), .Z(n6993) );
  NANDN U7168 ( .A(n6993), .B(n42173), .Z(n6954) );
  NANDN U7169 ( .A(n6952), .B(n42172), .Z(n6953) );
  NAND U7170 ( .A(n6954), .B(n6953), .Z(n7002) );
  NAND U7171 ( .A(b[7]), .B(a[160]), .Z(n7003) );
  XNOR U7172 ( .A(n7002), .B(n7003), .Z(n7005) );
  XOR U7173 ( .A(n7004), .B(n7005), .Z(n7011) );
  NANDN U7174 ( .A(n6955), .B(n42093), .Z(n6957) );
  XOR U7175 ( .A(n42134), .B(a[166]), .Z(n6996) );
  NANDN U7176 ( .A(n6996), .B(n42095), .Z(n6956) );
  NAND U7177 ( .A(n6957), .B(n6956), .Z(n7009) );
  NANDN U7178 ( .A(n6958), .B(n42231), .Z(n6960) );
  XOR U7179 ( .A(n175), .B(a[162]), .Z(n6999) );
  NANDN U7180 ( .A(n6999), .B(n42234), .Z(n6959) );
  AND U7181 ( .A(n6960), .B(n6959), .Z(n7008) );
  XNOR U7182 ( .A(n7009), .B(n7008), .Z(n7010) );
  XNOR U7183 ( .A(n7011), .B(n7010), .Z(n7015) );
  NANDN U7184 ( .A(n6962), .B(n6961), .Z(n6966) );
  NAND U7185 ( .A(n6964), .B(n6963), .Z(n6965) );
  AND U7186 ( .A(n6966), .B(n6965), .Z(n7014) );
  XOR U7187 ( .A(n7015), .B(n7014), .Z(n7016) );
  NANDN U7188 ( .A(n6968), .B(n6967), .Z(n6972) );
  NANDN U7189 ( .A(n6970), .B(n6969), .Z(n6971) );
  NAND U7190 ( .A(n6972), .B(n6971), .Z(n7017) );
  XOR U7191 ( .A(n7016), .B(n7017), .Z(n6984) );
  OR U7192 ( .A(n6974), .B(n6973), .Z(n6978) );
  NANDN U7193 ( .A(n6976), .B(n6975), .Z(n6977) );
  NAND U7194 ( .A(n6978), .B(n6977), .Z(n6985) );
  XNOR U7195 ( .A(n6984), .B(n6985), .Z(n6986) );
  XNOR U7196 ( .A(n6987), .B(n6986), .Z(n7020) );
  XNOR U7197 ( .A(n7020), .B(sreg[1184]), .Z(n7022) );
  NAND U7198 ( .A(n6979), .B(sreg[1183]), .Z(n6983) );
  OR U7199 ( .A(n6981), .B(n6980), .Z(n6982) );
  AND U7200 ( .A(n6983), .B(n6982), .Z(n7021) );
  XOR U7201 ( .A(n7022), .B(n7021), .Z(c[1184]) );
  NANDN U7202 ( .A(n6985), .B(n6984), .Z(n6989) );
  NAND U7203 ( .A(n6987), .B(n6986), .Z(n6988) );
  NAND U7204 ( .A(n6989), .B(n6988), .Z(n7028) );
  NAND U7205 ( .A(b[0]), .B(a[169]), .Z(n6990) );
  XNOR U7206 ( .A(b[1]), .B(n6990), .Z(n6992) );
  NAND U7207 ( .A(n39), .B(a[168]), .Z(n6991) );
  AND U7208 ( .A(n6992), .B(n6991), .Z(n7045) );
  XOR U7209 ( .A(a[165]), .B(n42197), .Z(n7034) );
  NANDN U7210 ( .A(n7034), .B(n42173), .Z(n6995) );
  NANDN U7211 ( .A(n6993), .B(n42172), .Z(n6994) );
  NAND U7212 ( .A(n6995), .B(n6994), .Z(n7043) );
  NAND U7213 ( .A(b[7]), .B(a[161]), .Z(n7044) );
  XNOR U7214 ( .A(n7043), .B(n7044), .Z(n7046) );
  XOR U7215 ( .A(n7045), .B(n7046), .Z(n7052) );
  NANDN U7216 ( .A(n6996), .B(n42093), .Z(n6998) );
  XOR U7217 ( .A(n42134), .B(a[167]), .Z(n7037) );
  NANDN U7218 ( .A(n7037), .B(n42095), .Z(n6997) );
  NAND U7219 ( .A(n6998), .B(n6997), .Z(n7050) );
  NANDN U7220 ( .A(n6999), .B(n42231), .Z(n7001) );
  XOR U7221 ( .A(n175), .B(a[163]), .Z(n7040) );
  NANDN U7222 ( .A(n7040), .B(n42234), .Z(n7000) );
  AND U7223 ( .A(n7001), .B(n7000), .Z(n7049) );
  XNOR U7224 ( .A(n7050), .B(n7049), .Z(n7051) );
  XNOR U7225 ( .A(n7052), .B(n7051), .Z(n7056) );
  NANDN U7226 ( .A(n7003), .B(n7002), .Z(n7007) );
  NAND U7227 ( .A(n7005), .B(n7004), .Z(n7006) );
  AND U7228 ( .A(n7007), .B(n7006), .Z(n7055) );
  XOR U7229 ( .A(n7056), .B(n7055), .Z(n7057) );
  NANDN U7230 ( .A(n7009), .B(n7008), .Z(n7013) );
  NANDN U7231 ( .A(n7011), .B(n7010), .Z(n7012) );
  NAND U7232 ( .A(n7013), .B(n7012), .Z(n7058) );
  XOR U7233 ( .A(n7057), .B(n7058), .Z(n7025) );
  OR U7234 ( .A(n7015), .B(n7014), .Z(n7019) );
  NANDN U7235 ( .A(n7017), .B(n7016), .Z(n7018) );
  NAND U7236 ( .A(n7019), .B(n7018), .Z(n7026) );
  XNOR U7237 ( .A(n7025), .B(n7026), .Z(n7027) );
  XNOR U7238 ( .A(n7028), .B(n7027), .Z(n7061) );
  XNOR U7239 ( .A(n7061), .B(sreg[1185]), .Z(n7063) );
  NAND U7240 ( .A(n7020), .B(sreg[1184]), .Z(n7024) );
  OR U7241 ( .A(n7022), .B(n7021), .Z(n7023) );
  AND U7242 ( .A(n7024), .B(n7023), .Z(n7062) );
  XOR U7243 ( .A(n7063), .B(n7062), .Z(c[1185]) );
  NANDN U7244 ( .A(n7026), .B(n7025), .Z(n7030) );
  NAND U7245 ( .A(n7028), .B(n7027), .Z(n7029) );
  NAND U7246 ( .A(n7030), .B(n7029), .Z(n7069) );
  NAND U7247 ( .A(b[0]), .B(a[170]), .Z(n7031) );
  XNOR U7248 ( .A(b[1]), .B(n7031), .Z(n7033) );
  NAND U7249 ( .A(n39), .B(a[169]), .Z(n7032) );
  AND U7250 ( .A(n7033), .B(n7032), .Z(n7086) );
  XOR U7251 ( .A(a[166]), .B(n42197), .Z(n7075) );
  NANDN U7252 ( .A(n7075), .B(n42173), .Z(n7036) );
  NANDN U7253 ( .A(n7034), .B(n42172), .Z(n7035) );
  NAND U7254 ( .A(n7036), .B(n7035), .Z(n7084) );
  NAND U7255 ( .A(b[7]), .B(a[162]), .Z(n7085) );
  XNOR U7256 ( .A(n7084), .B(n7085), .Z(n7087) );
  XOR U7257 ( .A(n7086), .B(n7087), .Z(n7093) );
  NANDN U7258 ( .A(n7037), .B(n42093), .Z(n7039) );
  XOR U7259 ( .A(n42134), .B(a[168]), .Z(n7078) );
  NANDN U7260 ( .A(n7078), .B(n42095), .Z(n7038) );
  NAND U7261 ( .A(n7039), .B(n7038), .Z(n7091) );
  NANDN U7262 ( .A(n7040), .B(n42231), .Z(n7042) );
  XOR U7263 ( .A(n175), .B(a[164]), .Z(n7081) );
  NANDN U7264 ( .A(n7081), .B(n42234), .Z(n7041) );
  AND U7265 ( .A(n7042), .B(n7041), .Z(n7090) );
  XNOR U7266 ( .A(n7091), .B(n7090), .Z(n7092) );
  XNOR U7267 ( .A(n7093), .B(n7092), .Z(n7097) );
  NANDN U7268 ( .A(n7044), .B(n7043), .Z(n7048) );
  NAND U7269 ( .A(n7046), .B(n7045), .Z(n7047) );
  AND U7270 ( .A(n7048), .B(n7047), .Z(n7096) );
  XOR U7271 ( .A(n7097), .B(n7096), .Z(n7098) );
  NANDN U7272 ( .A(n7050), .B(n7049), .Z(n7054) );
  NANDN U7273 ( .A(n7052), .B(n7051), .Z(n7053) );
  NAND U7274 ( .A(n7054), .B(n7053), .Z(n7099) );
  XOR U7275 ( .A(n7098), .B(n7099), .Z(n7066) );
  OR U7276 ( .A(n7056), .B(n7055), .Z(n7060) );
  NANDN U7277 ( .A(n7058), .B(n7057), .Z(n7059) );
  NAND U7278 ( .A(n7060), .B(n7059), .Z(n7067) );
  XNOR U7279 ( .A(n7066), .B(n7067), .Z(n7068) );
  XNOR U7280 ( .A(n7069), .B(n7068), .Z(n7102) );
  XNOR U7281 ( .A(n7102), .B(sreg[1186]), .Z(n7104) );
  NAND U7282 ( .A(n7061), .B(sreg[1185]), .Z(n7065) );
  OR U7283 ( .A(n7063), .B(n7062), .Z(n7064) );
  AND U7284 ( .A(n7065), .B(n7064), .Z(n7103) );
  XOR U7285 ( .A(n7104), .B(n7103), .Z(c[1186]) );
  NANDN U7286 ( .A(n7067), .B(n7066), .Z(n7071) );
  NAND U7287 ( .A(n7069), .B(n7068), .Z(n7070) );
  NAND U7288 ( .A(n7071), .B(n7070), .Z(n7110) );
  NAND U7289 ( .A(b[0]), .B(a[171]), .Z(n7072) );
  XNOR U7290 ( .A(b[1]), .B(n7072), .Z(n7074) );
  NAND U7291 ( .A(n39), .B(a[170]), .Z(n7073) );
  AND U7292 ( .A(n7074), .B(n7073), .Z(n7127) );
  XOR U7293 ( .A(a[167]), .B(n42197), .Z(n7116) );
  NANDN U7294 ( .A(n7116), .B(n42173), .Z(n7077) );
  NANDN U7295 ( .A(n7075), .B(n42172), .Z(n7076) );
  NAND U7296 ( .A(n7077), .B(n7076), .Z(n7125) );
  NAND U7297 ( .A(b[7]), .B(a[163]), .Z(n7126) );
  XNOR U7298 ( .A(n7125), .B(n7126), .Z(n7128) );
  XOR U7299 ( .A(n7127), .B(n7128), .Z(n7134) );
  NANDN U7300 ( .A(n7078), .B(n42093), .Z(n7080) );
  XOR U7301 ( .A(n42134), .B(a[169]), .Z(n7119) );
  NANDN U7302 ( .A(n7119), .B(n42095), .Z(n7079) );
  NAND U7303 ( .A(n7080), .B(n7079), .Z(n7132) );
  NANDN U7304 ( .A(n7081), .B(n42231), .Z(n7083) );
  XOR U7305 ( .A(n175), .B(a[165]), .Z(n7122) );
  NANDN U7306 ( .A(n7122), .B(n42234), .Z(n7082) );
  AND U7307 ( .A(n7083), .B(n7082), .Z(n7131) );
  XNOR U7308 ( .A(n7132), .B(n7131), .Z(n7133) );
  XNOR U7309 ( .A(n7134), .B(n7133), .Z(n7138) );
  NANDN U7310 ( .A(n7085), .B(n7084), .Z(n7089) );
  NAND U7311 ( .A(n7087), .B(n7086), .Z(n7088) );
  AND U7312 ( .A(n7089), .B(n7088), .Z(n7137) );
  XOR U7313 ( .A(n7138), .B(n7137), .Z(n7139) );
  NANDN U7314 ( .A(n7091), .B(n7090), .Z(n7095) );
  NANDN U7315 ( .A(n7093), .B(n7092), .Z(n7094) );
  NAND U7316 ( .A(n7095), .B(n7094), .Z(n7140) );
  XOR U7317 ( .A(n7139), .B(n7140), .Z(n7107) );
  OR U7318 ( .A(n7097), .B(n7096), .Z(n7101) );
  NANDN U7319 ( .A(n7099), .B(n7098), .Z(n7100) );
  NAND U7320 ( .A(n7101), .B(n7100), .Z(n7108) );
  XNOR U7321 ( .A(n7107), .B(n7108), .Z(n7109) );
  XNOR U7322 ( .A(n7110), .B(n7109), .Z(n7143) );
  XNOR U7323 ( .A(n7143), .B(sreg[1187]), .Z(n7145) );
  NAND U7324 ( .A(n7102), .B(sreg[1186]), .Z(n7106) );
  OR U7325 ( .A(n7104), .B(n7103), .Z(n7105) );
  AND U7326 ( .A(n7106), .B(n7105), .Z(n7144) );
  XOR U7327 ( .A(n7145), .B(n7144), .Z(c[1187]) );
  NANDN U7328 ( .A(n7108), .B(n7107), .Z(n7112) );
  NAND U7329 ( .A(n7110), .B(n7109), .Z(n7111) );
  NAND U7330 ( .A(n7112), .B(n7111), .Z(n7151) );
  NAND U7331 ( .A(b[0]), .B(a[172]), .Z(n7113) );
  XNOR U7332 ( .A(b[1]), .B(n7113), .Z(n7115) );
  NAND U7333 ( .A(n39), .B(a[171]), .Z(n7114) );
  AND U7334 ( .A(n7115), .B(n7114), .Z(n7168) );
  XOR U7335 ( .A(a[168]), .B(n42197), .Z(n7157) );
  NANDN U7336 ( .A(n7157), .B(n42173), .Z(n7118) );
  NANDN U7337 ( .A(n7116), .B(n42172), .Z(n7117) );
  NAND U7338 ( .A(n7118), .B(n7117), .Z(n7166) );
  NAND U7339 ( .A(b[7]), .B(a[164]), .Z(n7167) );
  XNOR U7340 ( .A(n7166), .B(n7167), .Z(n7169) );
  XOR U7341 ( .A(n7168), .B(n7169), .Z(n7175) );
  NANDN U7342 ( .A(n7119), .B(n42093), .Z(n7121) );
  XOR U7343 ( .A(n42134), .B(a[170]), .Z(n7160) );
  NANDN U7344 ( .A(n7160), .B(n42095), .Z(n7120) );
  NAND U7345 ( .A(n7121), .B(n7120), .Z(n7173) );
  NANDN U7346 ( .A(n7122), .B(n42231), .Z(n7124) );
  XOR U7347 ( .A(n175), .B(a[166]), .Z(n7163) );
  NANDN U7348 ( .A(n7163), .B(n42234), .Z(n7123) );
  AND U7349 ( .A(n7124), .B(n7123), .Z(n7172) );
  XNOR U7350 ( .A(n7173), .B(n7172), .Z(n7174) );
  XNOR U7351 ( .A(n7175), .B(n7174), .Z(n7179) );
  NANDN U7352 ( .A(n7126), .B(n7125), .Z(n7130) );
  NAND U7353 ( .A(n7128), .B(n7127), .Z(n7129) );
  AND U7354 ( .A(n7130), .B(n7129), .Z(n7178) );
  XOR U7355 ( .A(n7179), .B(n7178), .Z(n7180) );
  NANDN U7356 ( .A(n7132), .B(n7131), .Z(n7136) );
  NANDN U7357 ( .A(n7134), .B(n7133), .Z(n7135) );
  NAND U7358 ( .A(n7136), .B(n7135), .Z(n7181) );
  XOR U7359 ( .A(n7180), .B(n7181), .Z(n7148) );
  OR U7360 ( .A(n7138), .B(n7137), .Z(n7142) );
  NANDN U7361 ( .A(n7140), .B(n7139), .Z(n7141) );
  NAND U7362 ( .A(n7142), .B(n7141), .Z(n7149) );
  XNOR U7363 ( .A(n7148), .B(n7149), .Z(n7150) );
  XNOR U7364 ( .A(n7151), .B(n7150), .Z(n7184) );
  XNOR U7365 ( .A(n7184), .B(sreg[1188]), .Z(n7186) );
  NAND U7366 ( .A(n7143), .B(sreg[1187]), .Z(n7147) );
  OR U7367 ( .A(n7145), .B(n7144), .Z(n7146) );
  AND U7368 ( .A(n7147), .B(n7146), .Z(n7185) );
  XOR U7369 ( .A(n7186), .B(n7185), .Z(c[1188]) );
  NANDN U7370 ( .A(n7149), .B(n7148), .Z(n7153) );
  NAND U7371 ( .A(n7151), .B(n7150), .Z(n7152) );
  NAND U7372 ( .A(n7153), .B(n7152), .Z(n7192) );
  NAND U7373 ( .A(b[0]), .B(a[173]), .Z(n7154) );
  XNOR U7374 ( .A(b[1]), .B(n7154), .Z(n7156) );
  NAND U7375 ( .A(n39), .B(a[172]), .Z(n7155) );
  AND U7376 ( .A(n7156), .B(n7155), .Z(n7209) );
  XOR U7377 ( .A(a[169]), .B(n42197), .Z(n7198) );
  NANDN U7378 ( .A(n7198), .B(n42173), .Z(n7159) );
  NANDN U7379 ( .A(n7157), .B(n42172), .Z(n7158) );
  NAND U7380 ( .A(n7159), .B(n7158), .Z(n7207) );
  NAND U7381 ( .A(b[7]), .B(a[165]), .Z(n7208) );
  XNOR U7382 ( .A(n7207), .B(n7208), .Z(n7210) );
  XOR U7383 ( .A(n7209), .B(n7210), .Z(n7216) );
  NANDN U7384 ( .A(n7160), .B(n42093), .Z(n7162) );
  XOR U7385 ( .A(n42134), .B(a[171]), .Z(n7201) );
  NANDN U7386 ( .A(n7201), .B(n42095), .Z(n7161) );
  NAND U7387 ( .A(n7162), .B(n7161), .Z(n7214) );
  NANDN U7388 ( .A(n7163), .B(n42231), .Z(n7165) );
  XOR U7389 ( .A(n176), .B(a[167]), .Z(n7204) );
  NANDN U7390 ( .A(n7204), .B(n42234), .Z(n7164) );
  AND U7391 ( .A(n7165), .B(n7164), .Z(n7213) );
  XNOR U7392 ( .A(n7214), .B(n7213), .Z(n7215) );
  XNOR U7393 ( .A(n7216), .B(n7215), .Z(n7220) );
  NANDN U7394 ( .A(n7167), .B(n7166), .Z(n7171) );
  NAND U7395 ( .A(n7169), .B(n7168), .Z(n7170) );
  AND U7396 ( .A(n7171), .B(n7170), .Z(n7219) );
  XOR U7397 ( .A(n7220), .B(n7219), .Z(n7221) );
  NANDN U7398 ( .A(n7173), .B(n7172), .Z(n7177) );
  NANDN U7399 ( .A(n7175), .B(n7174), .Z(n7176) );
  NAND U7400 ( .A(n7177), .B(n7176), .Z(n7222) );
  XOR U7401 ( .A(n7221), .B(n7222), .Z(n7189) );
  OR U7402 ( .A(n7179), .B(n7178), .Z(n7183) );
  NANDN U7403 ( .A(n7181), .B(n7180), .Z(n7182) );
  NAND U7404 ( .A(n7183), .B(n7182), .Z(n7190) );
  XNOR U7405 ( .A(n7189), .B(n7190), .Z(n7191) );
  XNOR U7406 ( .A(n7192), .B(n7191), .Z(n7225) );
  XNOR U7407 ( .A(n7225), .B(sreg[1189]), .Z(n7227) );
  NAND U7408 ( .A(n7184), .B(sreg[1188]), .Z(n7188) );
  OR U7409 ( .A(n7186), .B(n7185), .Z(n7187) );
  AND U7410 ( .A(n7188), .B(n7187), .Z(n7226) );
  XOR U7411 ( .A(n7227), .B(n7226), .Z(c[1189]) );
  NANDN U7412 ( .A(n7190), .B(n7189), .Z(n7194) );
  NAND U7413 ( .A(n7192), .B(n7191), .Z(n7193) );
  NAND U7414 ( .A(n7194), .B(n7193), .Z(n7233) );
  NAND U7415 ( .A(b[0]), .B(a[174]), .Z(n7195) );
  XNOR U7416 ( .A(b[1]), .B(n7195), .Z(n7197) );
  NAND U7417 ( .A(n39), .B(a[173]), .Z(n7196) );
  AND U7418 ( .A(n7197), .B(n7196), .Z(n7250) );
  XOR U7419 ( .A(a[170]), .B(n42197), .Z(n7239) );
  NANDN U7420 ( .A(n7239), .B(n42173), .Z(n7200) );
  NANDN U7421 ( .A(n7198), .B(n42172), .Z(n7199) );
  NAND U7422 ( .A(n7200), .B(n7199), .Z(n7248) );
  NAND U7423 ( .A(b[7]), .B(a[166]), .Z(n7249) );
  XNOR U7424 ( .A(n7248), .B(n7249), .Z(n7251) );
  XOR U7425 ( .A(n7250), .B(n7251), .Z(n7257) );
  NANDN U7426 ( .A(n7201), .B(n42093), .Z(n7203) );
  XOR U7427 ( .A(n42134), .B(a[172]), .Z(n7242) );
  NANDN U7428 ( .A(n7242), .B(n42095), .Z(n7202) );
  NAND U7429 ( .A(n7203), .B(n7202), .Z(n7255) );
  NANDN U7430 ( .A(n7204), .B(n42231), .Z(n7206) );
  XOR U7431 ( .A(n176), .B(a[168]), .Z(n7245) );
  NANDN U7432 ( .A(n7245), .B(n42234), .Z(n7205) );
  AND U7433 ( .A(n7206), .B(n7205), .Z(n7254) );
  XNOR U7434 ( .A(n7255), .B(n7254), .Z(n7256) );
  XNOR U7435 ( .A(n7257), .B(n7256), .Z(n7261) );
  NANDN U7436 ( .A(n7208), .B(n7207), .Z(n7212) );
  NAND U7437 ( .A(n7210), .B(n7209), .Z(n7211) );
  AND U7438 ( .A(n7212), .B(n7211), .Z(n7260) );
  XOR U7439 ( .A(n7261), .B(n7260), .Z(n7262) );
  NANDN U7440 ( .A(n7214), .B(n7213), .Z(n7218) );
  NANDN U7441 ( .A(n7216), .B(n7215), .Z(n7217) );
  NAND U7442 ( .A(n7218), .B(n7217), .Z(n7263) );
  XOR U7443 ( .A(n7262), .B(n7263), .Z(n7230) );
  OR U7444 ( .A(n7220), .B(n7219), .Z(n7224) );
  NANDN U7445 ( .A(n7222), .B(n7221), .Z(n7223) );
  NAND U7446 ( .A(n7224), .B(n7223), .Z(n7231) );
  XNOR U7447 ( .A(n7230), .B(n7231), .Z(n7232) );
  XNOR U7448 ( .A(n7233), .B(n7232), .Z(n7266) );
  XNOR U7449 ( .A(n7266), .B(sreg[1190]), .Z(n7268) );
  NAND U7450 ( .A(n7225), .B(sreg[1189]), .Z(n7229) );
  OR U7451 ( .A(n7227), .B(n7226), .Z(n7228) );
  AND U7452 ( .A(n7229), .B(n7228), .Z(n7267) );
  XOR U7453 ( .A(n7268), .B(n7267), .Z(c[1190]) );
  NANDN U7454 ( .A(n7231), .B(n7230), .Z(n7235) );
  NAND U7455 ( .A(n7233), .B(n7232), .Z(n7234) );
  NAND U7456 ( .A(n7235), .B(n7234), .Z(n7274) );
  NAND U7457 ( .A(b[0]), .B(a[175]), .Z(n7236) );
  XNOR U7458 ( .A(b[1]), .B(n7236), .Z(n7238) );
  NAND U7459 ( .A(n40), .B(a[174]), .Z(n7237) );
  AND U7460 ( .A(n7238), .B(n7237), .Z(n7291) );
  XOR U7461 ( .A(a[171]), .B(n42197), .Z(n7280) );
  NANDN U7462 ( .A(n7280), .B(n42173), .Z(n7241) );
  NANDN U7463 ( .A(n7239), .B(n42172), .Z(n7240) );
  NAND U7464 ( .A(n7241), .B(n7240), .Z(n7289) );
  NAND U7465 ( .A(b[7]), .B(a[167]), .Z(n7290) );
  XNOR U7466 ( .A(n7289), .B(n7290), .Z(n7292) );
  XOR U7467 ( .A(n7291), .B(n7292), .Z(n7298) );
  NANDN U7468 ( .A(n7242), .B(n42093), .Z(n7244) );
  XOR U7469 ( .A(n42134), .B(a[173]), .Z(n7283) );
  NANDN U7470 ( .A(n7283), .B(n42095), .Z(n7243) );
  NAND U7471 ( .A(n7244), .B(n7243), .Z(n7296) );
  NANDN U7472 ( .A(n7245), .B(n42231), .Z(n7247) );
  XOR U7473 ( .A(n176), .B(a[169]), .Z(n7286) );
  NANDN U7474 ( .A(n7286), .B(n42234), .Z(n7246) );
  AND U7475 ( .A(n7247), .B(n7246), .Z(n7295) );
  XNOR U7476 ( .A(n7296), .B(n7295), .Z(n7297) );
  XNOR U7477 ( .A(n7298), .B(n7297), .Z(n7302) );
  NANDN U7478 ( .A(n7249), .B(n7248), .Z(n7253) );
  NAND U7479 ( .A(n7251), .B(n7250), .Z(n7252) );
  AND U7480 ( .A(n7253), .B(n7252), .Z(n7301) );
  XOR U7481 ( .A(n7302), .B(n7301), .Z(n7303) );
  NANDN U7482 ( .A(n7255), .B(n7254), .Z(n7259) );
  NANDN U7483 ( .A(n7257), .B(n7256), .Z(n7258) );
  NAND U7484 ( .A(n7259), .B(n7258), .Z(n7304) );
  XOR U7485 ( .A(n7303), .B(n7304), .Z(n7271) );
  OR U7486 ( .A(n7261), .B(n7260), .Z(n7265) );
  NANDN U7487 ( .A(n7263), .B(n7262), .Z(n7264) );
  NAND U7488 ( .A(n7265), .B(n7264), .Z(n7272) );
  XNOR U7489 ( .A(n7271), .B(n7272), .Z(n7273) );
  XNOR U7490 ( .A(n7274), .B(n7273), .Z(n7307) );
  XNOR U7491 ( .A(n7307), .B(sreg[1191]), .Z(n7309) );
  NAND U7492 ( .A(n7266), .B(sreg[1190]), .Z(n7270) );
  OR U7493 ( .A(n7268), .B(n7267), .Z(n7269) );
  AND U7494 ( .A(n7270), .B(n7269), .Z(n7308) );
  XOR U7495 ( .A(n7309), .B(n7308), .Z(c[1191]) );
  NANDN U7496 ( .A(n7272), .B(n7271), .Z(n7276) );
  NAND U7497 ( .A(n7274), .B(n7273), .Z(n7275) );
  NAND U7498 ( .A(n7276), .B(n7275), .Z(n7315) );
  NAND U7499 ( .A(b[0]), .B(a[176]), .Z(n7277) );
  XNOR U7500 ( .A(b[1]), .B(n7277), .Z(n7279) );
  NAND U7501 ( .A(n40), .B(a[175]), .Z(n7278) );
  AND U7502 ( .A(n7279), .B(n7278), .Z(n7332) );
  XOR U7503 ( .A(a[172]), .B(n42197), .Z(n7321) );
  NANDN U7504 ( .A(n7321), .B(n42173), .Z(n7282) );
  NANDN U7505 ( .A(n7280), .B(n42172), .Z(n7281) );
  NAND U7506 ( .A(n7282), .B(n7281), .Z(n7330) );
  NAND U7507 ( .A(b[7]), .B(a[168]), .Z(n7331) );
  XNOR U7508 ( .A(n7330), .B(n7331), .Z(n7333) );
  XOR U7509 ( .A(n7332), .B(n7333), .Z(n7339) );
  NANDN U7510 ( .A(n7283), .B(n42093), .Z(n7285) );
  XOR U7511 ( .A(n42134), .B(a[174]), .Z(n7324) );
  NANDN U7512 ( .A(n7324), .B(n42095), .Z(n7284) );
  NAND U7513 ( .A(n7285), .B(n7284), .Z(n7337) );
  NANDN U7514 ( .A(n7286), .B(n42231), .Z(n7288) );
  XOR U7515 ( .A(n176), .B(a[170]), .Z(n7327) );
  NANDN U7516 ( .A(n7327), .B(n42234), .Z(n7287) );
  AND U7517 ( .A(n7288), .B(n7287), .Z(n7336) );
  XNOR U7518 ( .A(n7337), .B(n7336), .Z(n7338) );
  XNOR U7519 ( .A(n7339), .B(n7338), .Z(n7343) );
  NANDN U7520 ( .A(n7290), .B(n7289), .Z(n7294) );
  NAND U7521 ( .A(n7292), .B(n7291), .Z(n7293) );
  AND U7522 ( .A(n7294), .B(n7293), .Z(n7342) );
  XOR U7523 ( .A(n7343), .B(n7342), .Z(n7344) );
  NANDN U7524 ( .A(n7296), .B(n7295), .Z(n7300) );
  NANDN U7525 ( .A(n7298), .B(n7297), .Z(n7299) );
  NAND U7526 ( .A(n7300), .B(n7299), .Z(n7345) );
  XOR U7527 ( .A(n7344), .B(n7345), .Z(n7312) );
  OR U7528 ( .A(n7302), .B(n7301), .Z(n7306) );
  NANDN U7529 ( .A(n7304), .B(n7303), .Z(n7305) );
  NAND U7530 ( .A(n7306), .B(n7305), .Z(n7313) );
  XNOR U7531 ( .A(n7312), .B(n7313), .Z(n7314) );
  XNOR U7532 ( .A(n7315), .B(n7314), .Z(n7348) );
  XNOR U7533 ( .A(n7348), .B(sreg[1192]), .Z(n7350) );
  NAND U7534 ( .A(n7307), .B(sreg[1191]), .Z(n7311) );
  OR U7535 ( .A(n7309), .B(n7308), .Z(n7310) );
  AND U7536 ( .A(n7311), .B(n7310), .Z(n7349) );
  XOR U7537 ( .A(n7350), .B(n7349), .Z(c[1192]) );
  NANDN U7538 ( .A(n7313), .B(n7312), .Z(n7317) );
  NAND U7539 ( .A(n7315), .B(n7314), .Z(n7316) );
  NAND U7540 ( .A(n7317), .B(n7316), .Z(n7356) );
  NAND U7541 ( .A(b[0]), .B(a[177]), .Z(n7318) );
  XNOR U7542 ( .A(b[1]), .B(n7318), .Z(n7320) );
  NAND U7543 ( .A(n40), .B(a[176]), .Z(n7319) );
  AND U7544 ( .A(n7320), .B(n7319), .Z(n7373) );
  XOR U7545 ( .A(a[173]), .B(n42197), .Z(n7362) );
  NANDN U7546 ( .A(n7362), .B(n42173), .Z(n7323) );
  NANDN U7547 ( .A(n7321), .B(n42172), .Z(n7322) );
  NAND U7548 ( .A(n7323), .B(n7322), .Z(n7371) );
  NAND U7549 ( .A(b[7]), .B(a[169]), .Z(n7372) );
  XNOR U7550 ( .A(n7371), .B(n7372), .Z(n7374) );
  XOR U7551 ( .A(n7373), .B(n7374), .Z(n7380) );
  NANDN U7552 ( .A(n7324), .B(n42093), .Z(n7326) );
  XOR U7553 ( .A(n42134), .B(a[175]), .Z(n7365) );
  NANDN U7554 ( .A(n7365), .B(n42095), .Z(n7325) );
  NAND U7555 ( .A(n7326), .B(n7325), .Z(n7378) );
  NANDN U7556 ( .A(n7327), .B(n42231), .Z(n7329) );
  XOR U7557 ( .A(n176), .B(a[171]), .Z(n7368) );
  NANDN U7558 ( .A(n7368), .B(n42234), .Z(n7328) );
  AND U7559 ( .A(n7329), .B(n7328), .Z(n7377) );
  XNOR U7560 ( .A(n7378), .B(n7377), .Z(n7379) );
  XNOR U7561 ( .A(n7380), .B(n7379), .Z(n7384) );
  NANDN U7562 ( .A(n7331), .B(n7330), .Z(n7335) );
  NAND U7563 ( .A(n7333), .B(n7332), .Z(n7334) );
  AND U7564 ( .A(n7335), .B(n7334), .Z(n7383) );
  XOR U7565 ( .A(n7384), .B(n7383), .Z(n7385) );
  NANDN U7566 ( .A(n7337), .B(n7336), .Z(n7341) );
  NANDN U7567 ( .A(n7339), .B(n7338), .Z(n7340) );
  NAND U7568 ( .A(n7341), .B(n7340), .Z(n7386) );
  XOR U7569 ( .A(n7385), .B(n7386), .Z(n7353) );
  OR U7570 ( .A(n7343), .B(n7342), .Z(n7347) );
  NANDN U7571 ( .A(n7345), .B(n7344), .Z(n7346) );
  NAND U7572 ( .A(n7347), .B(n7346), .Z(n7354) );
  XNOR U7573 ( .A(n7353), .B(n7354), .Z(n7355) );
  XNOR U7574 ( .A(n7356), .B(n7355), .Z(n7389) );
  XNOR U7575 ( .A(n7389), .B(sreg[1193]), .Z(n7391) );
  NAND U7576 ( .A(n7348), .B(sreg[1192]), .Z(n7352) );
  OR U7577 ( .A(n7350), .B(n7349), .Z(n7351) );
  AND U7578 ( .A(n7352), .B(n7351), .Z(n7390) );
  XOR U7579 ( .A(n7391), .B(n7390), .Z(c[1193]) );
  NANDN U7580 ( .A(n7354), .B(n7353), .Z(n7358) );
  NAND U7581 ( .A(n7356), .B(n7355), .Z(n7357) );
  NAND U7582 ( .A(n7358), .B(n7357), .Z(n7397) );
  NAND U7583 ( .A(b[0]), .B(a[178]), .Z(n7359) );
  XNOR U7584 ( .A(b[1]), .B(n7359), .Z(n7361) );
  NAND U7585 ( .A(n40), .B(a[177]), .Z(n7360) );
  AND U7586 ( .A(n7361), .B(n7360), .Z(n7414) );
  XOR U7587 ( .A(a[174]), .B(n42197), .Z(n7403) );
  NANDN U7588 ( .A(n7403), .B(n42173), .Z(n7364) );
  NANDN U7589 ( .A(n7362), .B(n42172), .Z(n7363) );
  NAND U7590 ( .A(n7364), .B(n7363), .Z(n7412) );
  NAND U7591 ( .A(b[7]), .B(a[170]), .Z(n7413) );
  XNOR U7592 ( .A(n7412), .B(n7413), .Z(n7415) );
  XOR U7593 ( .A(n7414), .B(n7415), .Z(n7421) );
  NANDN U7594 ( .A(n7365), .B(n42093), .Z(n7367) );
  XOR U7595 ( .A(n42134), .B(a[176]), .Z(n7406) );
  NANDN U7596 ( .A(n7406), .B(n42095), .Z(n7366) );
  NAND U7597 ( .A(n7367), .B(n7366), .Z(n7419) );
  NANDN U7598 ( .A(n7368), .B(n42231), .Z(n7370) );
  XOR U7599 ( .A(n176), .B(a[172]), .Z(n7409) );
  NANDN U7600 ( .A(n7409), .B(n42234), .Z(n7369) );
  AND U7601 ( .A(n7370), .B(n7369), .Z(n7418) );
  XNOR U7602 ( .A(n7419), .B(n7418), .Z(n7420) );
  XNOR U7603 ( .A(n7421), .B(n7420), .Z(n7425) );
  NANDN U7604 ( .A(n7372), .B(n7371), .Z(n7376) );
  NAND U7605 ( .A(n7374), .B(n7373), .Z(n7375) );
  AND U7606 ( .A(n7376), .B(n7375), .Z(n7424) );
  XOR U7607 ( .A(n7425), .B(n7424), .Z(n7426) );
  NANDN U7608 ( .A(n7378), .B(n7377), .Z(n7382) );
  NANDN U7609 ( .A(n7380), .B(n7379), .Z(n7381) );
  NAND U7610 ( .A(n7382), .B(n7381), .Z(n7427) );
  XOR U7611 ( .A(n7426), .B(n7427), .Z(n7394) );
  OR U7612 ( .A(n7384), .B(n7383), .Z(n7388) );
  NANDN U7613 ( .A(n7386), .B(n7385), .Z(n7387) );
  NAND U7614 ( .A(n7388), .B(n7387), .Z(n7395) );
  XNOR U7615 ( .A(n7394), .B(n7395), .Z(n7396) );
  XNOR U7616 ( .A(n7397), .B(n7396), .Z(n7430) );
  XNOR U7617 ( .A(n7430), .B(sreg[1194]), .Z(n7432) );
  NAND U7618 ( .A(n7389), .B(sreg[1193]), .Z(n7393) );
  OR U7619 ( .A(n7391), .B(n7390), .Z(n7392) );
  AND U7620 ( .A(n7393), .B(n7392), .Z(n7431) );
  XOR U7621 ( .A(n7432), .B(n7431), .Z(c[1194]) );
  NANDN U7622 ( .A(n7395), .B(n7394), .Z(n7399) );
  NAND U7623 ( .A(n7397), .B(n7396), .Z(n7398) );
  NAND U7624 ( .A(n7399), .B(n7398), .Z(n7438) );
  NAND U7625 ( .A(b[0]), .B(a[179]), .Z(n7400) );
  XNOR U7626 ( .A(b[1]), .B(n7400), .Z(n7402) );
  NAND U7627 ( .A(n40), .B(a[178]), .Z(n7401) );
  AND U7628 ( .A(n7402), .B(n7401), .Z(n7455) );
  XOR U7629 ( .A(a[175]), .B(n42197), .Z(n7444) );
  NANDN U7630 ( .A(n7444), .B(n42173), .Z(n7405) );
  NANDN U7631 ( .A(n7403), .B(n42172), .Z(n7404) );
  NAND U7632 ( .A(n7405), .B(n7404), .Z(n7453) );
  NAND U7633 ( .A(b[7]), .B(a[171]), .Z(n7454) );
  XNOR U7634 ( .A(n7453), .B(n7454), .Z(n7456) );
  XOR U7635 ( .A(n7455), .B(n7456), .Z(n7462) );
  NANDN U7636 ( .A(n7406), .B(n42093), .Z(n7408) );
  XOR U7637 ( .A(n42134), .B(a[177]), .Z(n7447) );
  NANDN U7638 ( .A(n7447), .B(n42095), .Z(n7407) );
  NAND U7639 ( .A(n7408), .B(n7407), .Z(n7460) );
  NANDN U7640 ( .A(n7409), .B(n42231), .Z(n7411) );
  XOR U7641 ( .A(n176), .B(a[173]), .Z(n7450) );
  NANDN U7642 ( .A(n7450), .B(n42234), .Z(n7410) );
  AND U7643 ( .A(n7411), .B(n7410), .Z(n7459) );
  XNOR U7644 ( .A(n7460), .B(n7459), .Z(n7461) );
  XNOR U7645 ( .A(n7462), .B(n7461), .Z(n7466) );
  NANDN U7646 ( .A(n7413), .B(n7412), .Z(n7417) );
  NAND U7647 ( .A(n7415), .B(n7414), .Z(n7416) );
  AND U7648 ( .A(n7417), .B(n7416), .Z(n7465) );
  XOR U7649 ( .A(n7466), .B(n7465), .Z(n7467) );
  NANDN U7650 ( .A(n7419), .B(n7418), .Z(n7423) );
  NANDN U7651 ( .A(n7421), .B(n7420), .Z(n7422) );
  NAND U7652 ( .A(n7423), .B(n7422), .Z(n7468) );
  XOR U7653 ( .A(n7467), .B(n7468), .Z(n7435) );
  OR U7654 ( .A(n7425), .B(n7424), .Z(n7429) );
  NANDN U7655 ( .A(n7427), .B(n7426), .Z(n7428) );
  NAND U7656 ( .A(n7429), .B(n7428), .Z(n7436) );
  XNOR U7657 ( .A(n7435), .B(n7436), .Z(n7437) );
  XNOR U7658 ( .A(n7438), .B(n7437), .Z(n7471) );
  XNOR U7659 ( .A(n7471), .B(sreg[1195]), .Z(n7473) );
  NAND U7660 ( .A(n7430), .B(sreg[1194]), .Z(n7434) );
  OR U7661 ( .A(n7432), .B(n7431), .Z(n7433) );
  AND U7662 ( .A(n7434), .B(n7433), .Z(n7472) );
  XOR U7663 ( .A(n7473), .B(n7472), .Z(c[1195]) );
  NANDN U7664 ( .A(n7436), .B(n7435), .Z(n7440) );
  NAND U7665 ( .A(n7438), .B(n7437), .Z(n7439) );
  NAND U7666 ( .A(n7440), .B(n7439), .Z(n7479) );
  NAND U7667 ( .A(b[0]), .B(a[180]), .Z(n7441) );
  XNOR U7668 ( .A(b[1]), .B(n7441), .Z(n7443) );
  NAND U7669 ( .A(n40), .B(a[179]), .Z(n7442) );
  AND U7670 ( .A(n7443), .B(n7442), .Z(n7496) );
  XOR U7671 ( .A(a[176]), .B(n42197), .Z(n7485) );
  NANDN U7672 ( .A(n7485), .B(n42173), .Z(n7446) );
  NANDN U7673 ( .A(n7444), .B(n42172), .Z(n7445) );
  NAND U7674 ( .A(n7446), .B(n7445), .Z(n7494) );
  NAND U7675 ( .A(b[7]), .B(a[172]), .Z(n7495) );
  XNOR U7676 ( .A(n7494), .B(n7495), .Z(n7497) );
  XOR U7677 ( .A(n7496), .B(n7497), .Z(n7503) );
  NANDN U7678 ( .A(n7447), .B(n42093), .Z(n7449) );
  XOR U7679 ( .A(n42134), .B(a[178]), .Z(n7488) );
  NANDN U7680 ( .A(n7488), .B(n42095), .Z(n7448) );
  NAND U7681 ( .A(n7449), .B(n7448), .Z(n7501) );
  NANDN U7682 ( .A(n7450), .B(n42231), .Z(n7452) );
  XOR U7683 ( .A(n176), .B(a[174]), .Z(n7491) );
  NANDN U7684 ( .A(n7491), .B(n42234), .Z(n7451) );
  AND U7685 ( .A(n7452), .B(n7451), .Z(n7500) );
  XNOR U7686 ( .A(n7501), .B(n7500), .Z(n7502) );
  XNOR U7687 ( .A(n7503), .B(n7502), .Z(n7507) );
  NANDN U7688 ( .A(n7454), .B(n7453), .Z(n7458) );
  NAND U7689 ( .A(n7456), .B(n7455), .Z(n7457) );
  AND U7690 ( .A(n7458), .B(n7457), .Z(n7506) );
  XOR U7691 ( .A(n7507), .B(n7506), .Z(n7508) );
  NANDN U7692 ( .A(n7460), .B(n7459), .Z(n7464) );
  NANDN U7693 ( .A(n7462), .B(n7461), .Z(n7463) );
  NAND U7694 ( .A(n7464), .B(n7463), .Z(n7509) );
  XOR U7695 ( .A(n7508), .B(n7509), .Z(n7476) );
  OR U7696 ( .A(n7466), .B(n7465), .Z(n7470) );
  NANDN U7697 ( .A(n7468), .B(n7467), .Z(n7469) );
  NAND U7698 ( .A(n7470), .B(n7469), .Z(n7477) );
  XNOR U7699 ( .A(n7476), .B(n7477), .Z(n7478) );
  XNOR U7700 ( .A(n7479), .B(n7478), .Z(n7512) );
  XNOR U7701 ( .A(n7512), .B(sreg[1196]), .Z(n7514) );
  NAND U7702 ( .A(n7471), .B(sreg[1195]), .Z(n7475) );
  OR U7703 ( .A(n7473), .B(n7472), .Z(n7474) );
  AND U7704 ( .A(n7475), .B(n7474), .Z(n7513) );
  XOR U7705 ( .A(n7514), .B(n7513), .Z(c[1196]) );
  NANDN U7706 ( .A(n7477), .B(n7476), .Z(n7481) );
  NAND U7707 ( .A(n7479), .B(n7478), .Z(n7480) );
  NAND U7708 ( .A(n7481), .B(n7480), .Z(n7520) );
  NAND U7709 ( .A(b[0]), .B(a[181]), .Z(n7482) );
  XNOR U7710 ( .A(b[1]), .B(n7482), .Z(n7484) );
  NAND U7711 ( .A(n40), .B(a[180]), .Z(n7483) );
  AND U7712 ( .A(n7484), .B(n7483), .Z(n7537) );
  XOR U7713 ( .A(a[177]), .B(n42197), .Z(n7526) );
  NANDN U7714 ( .A(n7526), .B(n42173), .Z(n7487) );
  NANDN U7715 ( .A(n7485), .B(n42172), .Z(n7486) );
  NAND U7716 ( .A(n7487), .B(n7486), .Z(n7535) );
  NAND U7717 ( .A(b[7]), .B(a[173]), .Z(n7536) );
  XNOR U7718 ( .A(n7535), .B(n7536), .Z(n7538) );
  XOR U7719 ( .A(n7537), .B(n7538), .Z(n7544) );
  NANDN U7720 ( .A(n7488), .B(n42093), .Z(n7490) );
  XOR U7721 ( .A(n42134), .B(a[179]), .Z(n7529) );
  NANDN U7722 ( .A(n7529), .B(n42095), .Z(n7489) );
  NAND U7723 ( .A(n7490), .B(n7489), .Z(n7542) );
  NANDN U7724 ( .A(n7491), .B(n42231), .Z(n7493) );
  XOR U7725 ( .A(n176), .B(a[175]), .Z(n7532) );
  NANDN U7726 ( .A(n7532), .B(n42234), .Z(n7492) );
  AND U7727 ( .A(n7493), .B(n7492), .Z(n7541) );
  XNOR U7728 ( .A(n7542), .B(n7541), .Z(n7543) );
  XNOR U7729 ( .A(n7544), .B(n7543), .Z(n7548) );
  NANDN U7730 ( .A(n7495), .B(n7494), .Z(n7499) );
  NAND U7731 ( .A(n7497), .B(n7496), .Z(n7498) );
  AND U7732 ( .A(n7499), .B(n7498), .Z(n7547) );
  XOR U7733 ( .A(n7548), .B(n7547), .Z(n7549) );
  NANDN U7734 ( .A(n7501), .B(n7500), .Z(n7505) );
  NANDN U7735 ( .A(n7503), .B(n7502), .Z(n7504) );
  NAND U7736 ( .A(n7505), .B(n7504), .Z(n7550) );
  XOR U7737 ( .A(n7549), .B(n7550), .Z(n7517) );
  OR U7738 ( .A(n7507), .B(n7506), .Z(n7511) );
  NANDN U7739 ( .A(n7509), .B(n7508), .Z(n7510) );
  NAND U7740 ( .A(n7511), .B(n7510), .Z(n7518) );
  XNOR U7741 ( .A(n7517), .B(n7518), .Z(n7519) );
  XNOR U7742 ( .A(n7520), .B(n7519), .Z(n7553) );
  XNOR U7743 ( .A(n7553), .B(sreg[1197]), .Z(n7555) );
  NAND U7744 ( .A(n7512), .B(sreg[1196]), .Z(n7516) );
  OR U7745 ( .A(n7514), .B(n7513), .Z(n7515) );
  AND U7746 ( .A(n7516), .B(n7515), .Z(n7554) );
  XOR U7747 ( .A(n7555), .B(n7554), .Z(c[1197]) );
  NANDN U7748 ( .A(n7518), .B(n7517), .Z(n7522) );
  NAND U7749 ( .A(n7520), .B(n7519), .Z(n7521) );
  NAND U7750 ( .A(n7522), .B(n7521), .Z(n7561) );
  NAND U7751 ( .A(b[0]), .B(a[182]), .Z(n7523) );
  XNOR U7752 ( .A(b[1]), .B(n7523), .Z(n7525) );
  NAND U7753 ( .A(n41), .B(a[181]), .Z(n7524) );
  AND U7754 ( .A(n7525), .B(n7524), .Z(n7578) );
  XOR U7755 ( .A(a[178]), .B(n42197), .Z(n7567) );
  NANDN U7756 ( .A(n7567), .B(n42173), .Z(n7528) );
  NANDN U7757 ( .A(n7526), .B(n42172), .Z(n7527) );
  NAND U7758 ( .A(n7528), .B(n7527), .Z(n7576) );
  NAND U7759 ( .A(b[7]), .B(a[174]), .Z(n7577) );
  XNOR U7760 ( .A(n7576), .B(n7577), .Z(n7579) );
  XOR U7761 ( .A(n7578), .B(n7579), .Z(n7585) );
  NANDN U7762 ( .A(n7529), .B(n42093), .Z(n7531) );
  XOR U7763 ( .A(n42134), .B(a[180]), .Z(n7570) );
  NANDN U7764 ( .A(n7570), .B(n42095), .Z(n7530) );
  NAND U7765 ( .A(n7531), .B(n7530), .Z(n7583) );
  NANDN U7766 ( .A(n7532), .B(n42231), .Z(n7534) );
  XOR U7767 ( .A(n176), .B(a[176]), .Z(n7573) );
  NANDN U7768 ( .A(n7573), .B(n42234), .Z(n7533) );
  AND U7769 ( .A(n7534), .B(n7533), .Z(n7582) );
  XNOR U7770 ( .A(n7583), .B(n7582), .Z(n7584) );
  XNOR U7771 ( .A(n7585), .B(n7584), .Z(n7589) );
  NANDN U7772 ( .A(n7536), .B(n7535), .Z(n7540) );
  NAND U7773 ( .A(n7538), .B(n7537), .Z(n7539) );
  AND U7774 ( .A(n7540), .B(n7539), .Z(n7588) );
  XOR U7775 ( .A(n7589), .B(n7588), .Z(n7590) );
  NANDN U7776 ( .A(n7542), .B(n7541), .Z(n7546) );
  NANDN U7777 ( .A(n7544), .B(n7543), .Z(n7545) );
  NAND U7778 ( .A(n7546), .B(n7545), .Z(n7591) );
  XOR U7779 ( .A(n7590), .B(n7591), .Z(n7558) );
  OR U7780 ( .A(n7548), .B(n7547), .Z(n7552) );
  NANDN U7781 ( .A(n7550), .B(n7549), .Z(n7551) );
  NAND U7782 ( .A(n7552), .B(n7551), .Z(n7559) );
  XNOR U7783 ( .A(n7558), .B(n7559), .Z(n7560) );
  XNOR U7784 ( .A(n7561), .B(n7560), .Z(n7594) );
  XNOR U7785 ( .A(n7594), .B(sreg[1198]), .Z(n7596) );
  NAND U7786 ( .A(n7553), .B(sreg[1197]), .Z(n7557) );
  OR U7787 ( .A(n7555), .B(n7554), .Z(n7556) );
  AND U7788 ( .A(n7557), .B(n7556), .Z(n7595) );
  XOR U7789 ( .A(n7596), .B(n7595), .Z(c[1198]) );
  NANDN U7790 ( .A(n7559), .B(n7558), .Z(n7563) );
  NAND U7791 ( .A(n7561), .B(n7560), .Z(n7562) );
  NAND U7792 ( .A(n7563), .B(n7562), .Z(n7602) );
  NAND U7793 ( .A(b[0]), .B(a[183]), .Z(n7564) );
  XNOR U7794 ( .A(b[1]), .B(n7564), .Z(n7566) );
  NAND U7795 ( .A(n41), .B(a[182]), .Z(n7565) );
  AND U7796 ( .A(n7566), .B(n7565), .Z(n7619) );
  XOR U7797 ( .A(a[179]), .B(n42197), .Z(n7608) );
  NANDN U7798 ( .A(n7608), .B(n42173), .Z(n7569) );
  NANDN U7799 ( .A(n7567), .B(n42172), .Z(n7568) );
  NAND U7800 ( .A(n7569), .B(n7568), .Z(n7617) );
  NAND U7801 ( .A(b[7]), .B(a[175]), .Z(n7618) );
  XNOR U7802 ( .A(n7617), .B(n7618), .Z(n7620) );
  XOR U7803 ( .A(n7619), .B(n7620), .Z(n7626) );
  NANDN U7804 ( .A(n7570), .B(n42093), .Z(n7572) );
  XOR U7805 ( .A(n42134), .B(a[181]), .Z(n7611) );
  NANDN U7806 ( .A(n7611), .B(n42095), .Z(n7571) );
  NAND U7807 ( .A(n7572), .B(n7571), .Z(n7624) );
  NANDN U7808 ( .A(n7573), .B(n42231), .Z(n7575) );
  XOR U7809 ( .A(n176), .B(a[177]), .Z(n7614) );
  NANDN U7810 ( .A(n7614), .B(n42234), .Z(n7574) );
  AND U7811 ( .A(n7575), .B(n7574), .Z(n7623) );
  XNOR U7812 ( .A(n7624), .B(n7623), .Z(n7625) );
  XNOR U7813 ( .A(n7626), .B(n7625), .Z(n7630) );
  NANDN U7814 ( .A(n7577), .B(n7576), .Z(n7581) );
  NAND U7815 ( .A(n7579), .B(n7578), .Z(n7580) );
  AND U7816 ( .A(n7581), .B(n7580), .Z(n7629) );
  XOR U7817 ( .A(n7630), .B(n7629), .Z(n7631) );
  NANDN U7818 ( .A(n7583), .B(n7582), .Z(n7587) );
  NANDN U7819 ( .A(n7585), .B(n7584), .Z(n7586) );
  NAND U7820 ( .A(n7587), .B(n7586), .Z(n7632) );
  XOR U7821 ( .A(n7631), .B(n7632), .Z(n7599) );
  OR U7822 ( .A(n7589), .B(n7588), .Z(n7593) );
  NANDN U7823 ( .A(n7591), .B(n7590), .Z(n7592) );
  NAND U7824 ( .A(n7593), .B(n7592), .Z(n7600) );
  XNOR U7825 ( .A(n7599), .B(n7600), .Z(n7601) );
  XNOR U7826 ( .A(n7602), .B(n7601), .Z(n7635) );
  XNOR U7827 ( .A(n7635), .B(sreg[1199]), .Z(n7637) );
  NAND U7828 ( .A(n7594), .B(sreg[1198]), .Z(n7598) );
  OR U7829 ( .A(n7596), .B(n7595), .Z(n7597) );
  AND U7830 ( .A(n7598), .B(n7597), .Z(n7636) );
  XOR U7831 ( .A(n7637), .B(n7636), .Z(c[1199]) );
  NANDN U7832 ( .A(n7600), .B(n7599), .Z(n7604) );
  NAND U7833 ( .A(n7602), .B(n7601), .Z(n7603) );
  NAND U7834 ( .A(n7604), .B(n7603), .Z(n7643) );
  NAND U7835 ( .A(b[0]), .B(a[184]), .Z(n7605) );
  XNOR U7836 ( .A(b[1]), .B(n7605), .Z(n7607) );
  NAND U7837 ( .A(n41), .B(a[183]), .Z(n7606) );
  AND U7838 ( .A(n7607), .B(n7606), .Z(n7660) );
  XOR U7839 ( .A(a[180]), .B(n42197), .Z(n7649) );
  NANDN U7840 ( .A(n7649), .B(n42173), .Z(n7610) );
  NANDN U7841 ( .A(n7608), .B(n42172), .Z(n7609) );
  NAND U7842 ( .A(n7610), .B(n7609), .Z(n7658) );
  NAND U7843 ( .A(b[7]), .B(a[176]), .Z(n7659) );
  XNOR U7844 ( .A(n7658), .B(n7659), .Z(n7661) );
  XOR U7845 ( .A(n7660), .B(n7661), .Z(n7667) );
  NANDN U7846 ( .A(n7611), .B(n42093), .Z(n7613) );
  XOR U7847 ( .A(n42134), .B(a[182]), .Z(n7652) );
  NANDN U7848 ( .A(n7652), .B(n42095), .Z(n7612) );
  NAND U7849 ( .A(n7613), .B(n7612), .Z(n7665) );
  NANDN U7850 ( .A(n7614), .B(n42231), .Z(n7616) );
  XOR U7851 ( .A(n176), .B(a[178]), .Z(n7655) );
  NANDN U7852 ( .A(n7655), .B(n42234), .Z(n7615) );
  AND U7853 ( .A(n7616), .B(n7615), .Z(n7664) );
  XNOR U7854 ( .A(n7665), .B(n7664), .Z(n7666) );
  XNOR U7855 ( .A(n7667), .B(n7666), .Z(n7671) );
  NANDN U7856 ( .A(n7618), .B(n7617), .Z(n7622) );
  NAND U7857 ( .A(n7620), .B(n7619), .Z(n7621) );
  AND U7858 ( .A(n7622), .B(n7621), .Z(n7670) );
  XOR U7859 ( .A(n7671), .B(n7670), .Z(n7672) );
  NANDN U7860 ( .A(n7624), .B(n7623), .Z(n7628) );
  NANDN U7861 ( .A(n7626), .B(n7625), .Z(n7627) );
  NAND U7862 ( .A(n7628), .B(n7627), .Z(n7673) );
  XOR U7863 ( .A(n7672), .B(n7673), .Z(n7640) );
  OR U7864 ( .A(n7630), .B(n7629), .Z(n7634) );
  NANDN U7865 ( .A(n7632), .B(n7631), .Z(n7633) );
  NAND U7866 ( .A(n7634), .B(n7633), .Z(n7641) );
  XNOR U7867 ( .A(n7640), .B(n7641), .Z(n7642) );
  XNOR U7868 ( .A(n7643), .B(n7642), .Z(n7676) );
  XNOR U7869 ( .A(n7676), .B(sreg[1200]), .Z(n7678) );
  NAND U7870 ( .A(n7635), .B(sreg[1199]), .Z(n7639) );
  OR U7871 ( .A(n7637), .B(n7636), .Z(n7638) );
  AND U7872 ( .A(n7639), .B(n7638), .Z(n7677) );
  XOR U7873 ( .A(n7678), .B(n7677), .Z(c[1200]) );
  NANDN U7874 ( .A(n7641), .B(n7640), .Z(n7645) );
  NAND U7875 ( .A(n7643), .B(n7642), .Z(n7644) );
  NAND U7876 ( .A(n7645), .B(n7644), .Z(n7684) );
  NAND U7877 ( .A(b[0]), .B(a[185]), .Z(n7646) );
  XNOR U7878 ( .A(b[1]), .B(n7646), .Z(n7648) );
  NAND U7879 ( .A(n41), .B(a[184]), .Z(n7647) );
  AND U7880 ( .A(n7648), .B(n7647), .Z(n7701) );
  XOR U7881 ( .A(a[181]), .B(n42197), .Z(n7690) );
  NANDN U7882 ( .A(n7690), .B(n42173), .Z(n7651) );
  NANDN U7883 ( .A(n7649), .B(n42172), .Z(n7650) );
  NAND U7884 ( .A(n7651), .B(n7650), .Z(n7699) );
  NAND U7885 ( .A(b[7]), .B(a[177]), .Z(n7700) );
  XNOR U7886 ( .A(n7699), .B(n7700), .Z(n7702) );
  XOR U7887 ( .A(n7701), .B(n7702), .Z(n7708) );
  NANDN U7888 ( .A(n7652), .B(n42093), .Z(n7654) );
  XOR U7889 ( .A(n42134), .B(a[183]), .Z(n7693) );
  NANDN U7890 ( .A(n7693), .B(n42095), .Z(n7653) );
  NAND U7891 ( .A(n7654), .B(n7653), .Z(n7706) );
  NANDN U7892 ( .A(n7655), .B(n42231), .Z(n7657) );
  XOR U7893 ( .A(n177), .B(a[179]), .Z(n7696) );
  NANDN U7894 ( .A(n7696), .B(n42234), .Z(n7656) );
  AND U7895 ( .A(n7657), .B(n7656), .Z(n7705) );
  XNOR U7896 ( .A(n7706), .B(n7705), .Z(n7707) );
  XNOR U7897 ( .A(n7708), .B(n7707), .Z(n7712) );
  NANDN U7898 ( .A(n7659), .B(n7658), .Z(n7663) );
  NAND U7899 ( .A(n7661), .B(n7660), .Z(n7662) );
  AND U7900 ( .A(n7663), .B(n7662), .Z(n7711) );
  XOR U7901 ( .A(n7712), .B(n7711), .Z(n7713) );
  NANDN U7902 ( .A(n7665), .B(n7664), .Z(n7669) );
  NANDN U7903 ( .A(n7667), .B(n7666), .Z(n7668) );
  NAND U7904 ( .A(n7669), .B(n7668), .Z(n7714) );
  XOR U7905 ( .A(n7713), .B(n7714), .Z(n7681) );
  OR U7906 ( .A(n7671), .B(n7670), .Z(n7675) );
  NANDN U7907 ( .A(n7673), .B(n7672), .Z(n7674) );
  NAND U7908 ( .A(n7675), .B(n7674), .Z(n7682) );
  XNOR U7909 ( .A(n7681), .B(n7682), .Z(n7683) );
  XNOR U7910 ( .A(n7684), .B(n7683), .Z(n7717) );
  XNOR U7911 ( .A(n7717), .B(sreg[1201]), .Z(n7719) );
  NAND U7912 ( .A(n7676), .B(sreg[1200]), .Z(n7680) );
  OR U7913 ( .A(n7678), .B(n7677), .Z(n7679) );
  AND U7914 ( .A(n7680), .B(n7679), .Z(n7718) );
  XOR U7915 ( .A(n7719), .B(n7718), .Z(c[1201]) );
  NANDN U7916 ( .A(n7682), .B(n7681), .Z(n7686) );
  NAND U7917 ( .A(n7684), .B(n7683), .Z(n7685) );
  NAND U7918 ( .A(n7686), .B(n7685), .Z(n7725) );
  NAND U7919 ( .A(b[0]), .B(a[186]), .Z(n7687) );
  XNOR U7920 ( .A(b[1]), .B(n7687), .Z(n7689) );
  NAND U7921 ( .A(n41), .B(a[185]), .Z(n7688) );
  AND U7922 ( .A(n7689), .B(n7688), .Z(n7742) );
  XOR U7923 ( .A(a[182]), .B(n42197), .Z(n7731) );
  NANDN U7924 ( .A(n7731), .B(n42173), .Z(n7692) );
  NANDN U7925 ( .A(n7690), .B(n42172), .Z(n7691) );
  NAND U7926 ( .A(n7692), .B(n7691), .Z(n7740) );
  NAND U7927 ( .A(b[7]), .B(a[178]), .Z(n7741) );
  XNOR U7928 ( .A(n7740), .B(n7741), .Z(n7743) );
  XOR U7929 ( .A(n7742), .B(n7743), .Z(n7749) );
  NANDN U7930 ( .A(n7693), .B(n42093), .Z(n7695) );
  XOR U7931 ( .A(n42134), .B(a[184]), .Z(n7734) );
  NANDN U7932 ( .A(n7734), .B(n42095), .Z(n7694) );
  NAND U7933 ( .A(n7695), .B(n7694), .Z(n7747) );
  NANDN U7934 ( .A(n7696), .B(n42231), .Z(n7698) );
  XOR U7935 ( .A(n177), .B(a[180]), .Z(n7737) );
  NANDN U7936 ( .A(n7737), .B(n42234), .Z(n7697) );
  AND U7937 ( .A(n7698), .B(n7697), .Z(n7746) );
  XNOR U7938 ( .A(n7747), .B(n7746), .Z(n7748) );
  XNOR U7939 ( .A(n7749), .B(n7748), .Z(n7753) );
  NANDN U7940 ( .A(n7700), .B(n7699), .Z(n7704) );
  NAND U7941 ( .A(n7702), .B(n7701), .Z(n7703) );
  AND U7942 ( .A(n7704), .B(n7703), .Z(n7752) );
  XOR U7943 ( .A(n7753), .B(n7752), .Z(n7754) );
  NANDN U7944 ( .A(n7706), .B(n7705), .Z(n7710) );
  NANDN U7945 ( .A(n7708), .B(n7707), .Z(n7709) );
  NAND U7946 ( .A(n7710), .B(n7709), .Z(n7755) );
  XOR U7947 ( .A(n7754), .B(n7755), .Z(n7722) );
  OR U7948 ( .A(n7712), .B(n7711), .Z(n7716) );
  NANDN U7949 ( .A(n7714), .B(n7713), .Z(n7715) );
  NAND U7950 ( .A(n7716), .B(n7715), .Z(n7723) );
  XNOR U7951 ( .A(n7722), .B(n7723), .Z(n7724) );
  XNOR U7952 ( .A(n7725), .B(n7724), .Z(n7758) );
  XNOR U7953 ( .A(n7758), .B(sreg[1202]), .Z(n7760) );
  NAND U7954 ( .A(n7717), .B(sreg[1201]), .Z(n7721) );
  OR U7955 ( .A(n7719), .B(n7718), .Z(n7720) );
  AND U7956 ( .A(n7721), .B(n7720), .Z(n7759) );
  XOR U7957 ( .A(n7760), .B(n7759), .Z(c[1202]) );
  NANDN U7958 ( .A(n7723), .B(n7722), .Z(n7727) );
  NAND U7959 ( .A(n7725), .B(n7724), .Z(n7726) );
  NAND U7960 ( .A(n7727), .B(n7726), .Z(n7766) );
  NAND U7961 ( .A(b[0]), .B(a[187]), .Z(n7728) );
  XNOR U7962 ( .A(b[1]), .B(n7728), .Z(n7730) );
  NAND U7963 ( .A(n41), .B(a[186]), .Z(n7729) );
  AND U7964 ( .A(n7730), .B(n7729), .Z(n7783) );
  XOR U7965 ( .A(a[183]), .B(n42197), .Z(n7772) );
  NANDN U7966 ( .A(n7772), .B(n42173), .Z(n7733) );
  NANDN U7967 ( .A(n7731), .B(n42172), .Z(n7732) );
  NAND U7968 ( .A(n7733), .B(n7732), .Z(n7781) );
  NAND U7969 ( .A(b[7]), .B(a[179]), .Z(n7782) );
  XNOR U7970 ( .A(n7781), .B(n7782), .Z(n7784) );
  XOR U7971 ( .A(n7783), .B(n7784), .Z(n7790) );
  NANDN U7972 ( .A(n7734), .B(n42093), .Z(n7736) );
  XOR U7973 ( .A(n42134), .B(a[185]), .Z(n7775) );
  NANDN U7974 ( .A(n7775), .B(n42095), .Z(n7735) );
  NAND U7975 ( .A(n7736), .B(n7735), .Z(n7788) );
  NANDN U7976 ( .A(n7737), .B(n42231), .Z(n7739) );
  XOR U7977 ( .A(n177), .B(a[181]), .Z(n7778) );
  NANDN U7978 ( .A(n7778), .B(n42234), .Z(n7738) );
  AND U7979 ( .A(n7739), .B(n7738), .Z(n7787) );
  XNOR U7980 ( .A(n7788), .B(n7787), .Z(n7789) );
  XNOR U7981 ( .A(n7790), .B(n7789), .Z(n7794) );
  NANDN U7982 ( .A(n7741), .B(n7740), .Z(n7745) );
  NAND U7983 ( .A(n7743), .B(n7742), .Z(n7744) );
  AND U7984 ( .A(n7745), .B(n7744), .Z(n7793) );
  XOR U7985 ( .A(n7794), .B(n7793), .Z(n7795) );
  NANDN U7986 ( .A(n7747), .B(n7746), .Z(n7751) );
  NANDN U7987 ( .A(n7749), .B(n7748), .Z(n7750) );
  NAND U7988 ( .A(n7751), .B(n7750), .Z(n7796) );
  XOR U7989 ( .A(n7795), .B(n7796), .Z(n7763) );
  OR U7990 ( .A(n7753), .B(n7752), .Z(n7757) );
  NANDN U7991 ( .A(n7755), .B(n7754), .Z(n7756) );
  NAND U7992 ( .A(n7757), .B(n7756), .Z(n7764) );
  XNOR U7993 ( .A(n7763), .B(n7764), .Z(n7765) );
  XNOR U7994 ( .A(n7766), .B(n7765), .Z(n7799) );
  XNOR U7995 ( .A(n7799), .B(sreg[1203]), .Z(n7801) );
  NAND U7996 ( .A(n7758), .B(sreg[1202]), .Z(n7762) );
  OR U7997 ( .A(n7760), .B(n7759), .Z(n7761) );
  AND U7998 ( .A(n7762), .B(n7761), .Z(n7800) );
  XOR U7999 ( .A(n7801), .B(n7800), .Z(c[1203]) );
  NANDN U8000 ( .A(n7764), .B(n7763), .Z(n7768) );
  NAND U8001 ( .A(n7766), .B(n7765), .Z(n7767) );
  NAND U8002 ( .A(n7768), .B(n7767), .Z(n7807) );
  NAND U8003 ( .A(b[0]), .B(a[188]), .Z(n7769) );
  XNOR U8004 ( .A(b[1]), .B(n7769), .Z(n7771) );
  NAND U8005 ( .A(n41), .B(a[187]), .Z(n7770) );
  AND U8006 ( .A(n7771), .B(n7770), .Z(n7824) );
  XOR U8007 ( .A(a[184]), .B(n42197), .Z(n7813) );
  NANDN U8008 ( .A(n7813), .B(n42173), .Z(n7774) );
  NANDN U8009 ( .A(n7772), .B(n42172), .Z(n7773) );
  NAND U8010 ( .A(n7774), .B(n7773), .Z(n7822) );
  NAND U8011 ( .A(b[7]), .B(a[180]), .Z(n7823) );
  XNOR U8012 ( .A(n7822), .B(n7823), .Z(n7825) );
  XOR U8013 ( .A(n7824), .B(n7825), .Z(n7831) );
  NANDN U8014 ( .A(n7775), .B(n42093), .Z(n7777) );
  XOR U8015 ( .A(n42134), .B(a[186]), .Z(n7816) );
  NANDN U8016 ( .A(n7816), .B(n42095), .Z(n7776) );
  NAND U8017 ( .A(n7777), .B(n7776), .Z(n7829) );
  NANDN U8018 ( .A(n7778), .B(n42231), .Z(n7780) );
  XOR U8019 ( .A(n177), .B(a[182]), .Z(n7819) );
  NANDN U8020 ( .A(n7819), .B(n42234), .Z(n7779) );
  AND U8021 ( .A(n7780), .B(n7779), .Z(n7828) );
  XNOR U8022 ( .A(n7829), .B(n7828), .Z(n7830) );
  XNOR U8023 ( .A(n7831), .B(n7830), .Z(n7835) );
  NANDN U8024 ( .A(n7782), .B(n7781), .Z(n7786) );
  NAND U8025 ( .A(n7784), .B(n7783), .Z(n7785) );
  AND U8026 ( .A(n7786), .B(n7785), .Z(n7834) );
  XOR U8027 ( .A(n7835), .B(n7834), .Z(n7836) );
  NANDN U8028 ( .A(n7788), .B(n7787), .Z(n7792) );
  NANDN U8029 ( .A(n7790), .B(n7789), .Z(n7791) );
  NAND U8030 ( .A(n7792), .B(n7791), .Z(n7837) );
  XOR U8031 ( .A(n7836), .B(n7837), .Z(n7804) );
  OR U8032 ( .A(n7794), .B(n7793), .Z(n7798) );
  NANDN U8033 ( .A(n7796), .B(n7795), .Z(n7797) );
  NAND U8034 ( .A(n7798), .B(n7797), .Z(n7805) );
  XNOR U8035 ( .A(n7804), .B(n7805), .Z(n7806) );
  XNOR U8036 ( .A(n7807), .B(n7806), .Z(n7840) );
  XNOR U8037 ( .A(n7840), .B(sreg[1204]), .Z(n7842) );
  NAND U8038 ( .A(n7799), .B(sreg[1203]), .Z(n7803) );
  OR U8039 ( .A(n7801), .B(n7800), .Z(n7802) );
  AND U8040 ( .A(n7803), .B(n7802), .Z(n7841) );
  XOR U8041 ( .A(n7842), .B(n7841), .Z(c[1204]) );
  NANDN U8042 ( .A(n7805), .B(n7804), .Z(n7809) );
  NAND U8043 ( .A(n7807), .B(n7806), .Z(n7808) );
  NAND U8044 ( .A(n7809), .B(n7808), .Z(n7848) );
  NAND U8045 ( .A(b[0]), .B(a[189]), .Z(n7810) );
  XNOR U8046 ( .A(b[1]), .B(n7810), .Z(n7812) );
  NAND U8047 ( .A(n42), .B(a[188]), .Z(n7811) );
  AND U8048 ( .A(n7812), .B(n7811), .Z(n7865) );
  XOR U8049 ( .A(a[185]), .B(n42197), .Z(n7854) );
  NANDN U8050 ( .A(n7854), .B(n42173), .Z(n7815) );
  NANDN U8051 ( .A(n7813), .B(n42172), .Z(n7814) );
  NAND U8052 ( .A(n7815), .B(n7814), .Z(n7863) );
  NAND U8053 ( .A(b[7]), .B(a[181]), .Z(n7864) );
  XNOR U8054 ( .A(n7863), .B(n7864), .Z(n7866) );
  XOR U8055 ( .A(n7865), .B(n7866), .Z(n7872) );
  NANDN U8056 ( .A(n7816), .B(n42093), .Z(n7818) );
  XOR U8057 ( .A(n42134), .B(a[187]), .Z(n7857) );
  NANDN U8058 ( .A(n7857), .B(n42095), .Z(n7817) );
  NAND U8059 ( .A(n7818), .B(n7817), .Z(n7870) );
  NANDN U8060 ( .A(n7819), .B(n42231), .Z(n7821) );
  XOR U8061 ( .A(n177), .B(a[183]), .Z(n7860) );
  NANDN U8062 ( .A(n7860), .B(n42234), .Z(n7820) );
  AND U8063 ( .A(n7821), .B(n7820), .Z(n7869) );
  XNOR U8064 ( .A(n7870), .B(n7869), .Z(n7871) );
  XNOR U8065 ( .A(n7872), .B(n7871), .Z(n7876) );
  NANDN U8066 ( .A(n7823), .B(n7822), .Z(n7827) );
  NAND U8067 ( .A(n7825), .B(n7824), .Z(n7826) );
  AND U8068 ( .A(n7827), .B(n7826), .Z(n7875) );
  XOR U8069 ( .A(n7876), .B(n7875), .Z(n7877) );
  NANDN U8070 ( .A(n7829), .B(n7828), .Z(n7833) );
  NANDN U8071 ( .A(n7831), .B(n7830), .Z(n7832) );
  NAND U8072 ( .A(n7833), .B(n7832), .Z(n7878) );
  XOR U8073 ( .A(n7877), .B(n7878), .Z(n7845) );
  OR U8074 ( .A(n7835), .B(n7834), .Z(n7839) );
  NANDN U8075 ( .A(n7837), .B(n7836), .Z(n7838) );
  NAND U8076 ( .A(n7839), .B(n7838), .Z(n7846) );
  XNOR U8077 ( .A(n7845), .B(n7846), .Z(n7847) );
  XNOR U8078 ( .A(n7848), .B(n7847), .Z(n7881) );
  XNOR U8079 ( .A(n7881), .B(sreg[1205]), .Z(n7883) );
  NAND U8080 ( .A(n7840), .B(sreg[1204]), .Z(n7844) );
  OR U8081 ( .A(n7842), .B(n7841), .Z(n7843) );
  AND U8082 ( .A(n7844), .B(n7843), .Z(n7882) );
  XOR U8083 ( .A(n7883), .B(n7882), .Z(c[1205]) );
  NANDN U8084 ( .A(n7846), .B(n7845), .Z(n7850) );
  NAND U8085 ( .A(n7848), .B(n7847), .Z(n7849) );
  NAND U8086 ( .A(n7850), .B(n7849), .Z(n7889) );
  NAND U8087 ( .A(b[0]), .B(a[190]), .Z(n7851) );
  XNOR U8088 ( .A(b[1]), .B(n7851), .Z(n7853) );
  NAND U8089 ( .A(n42), .B(a[189]), .Z(n7852) );
  AND U8090 ( .A(n7853), .B(n7852), .Z(n7906) );
  XOR U8091 ( .A(a[186]), .B(n42197), .Z(n7895) );
  NANDN U8092 ( .A(n7895), .B(n42173), .Z(n7856) );
  NANDN U8093 ( .A(n7854), .B(n42172), .Z(n7855) );
  NAND U8094 ( .A(n7856), .B(n7855), .Z(n7904) );
  NAND U8095 ( .A(b[7]), .B(a[182]), .Z(n7905) );
  XNOR U8096 ( .A(n7904), .B(n7905), .Z(n7907) );
  XOR U8097 ( .A(n7906), .B(n7907), .Z(n7913) );
  NANDN U8098 ( .A(n7857), .B(n42093), .Z(n7859) );
  XOR U8099 ( .A(n42134), .B(a[188]), .Z(n7898) );
  NANDN U8100 ( .A(n7898), .B(n42095), .Z(n7858) );
  NAND U8101 ( .A(n7859), .B(n7858), .Z(n7911) );
  NANDN U8102 ( .A(n7860), .B(n42231), .Z(n7862) );
  XOR U8103 ( .A(n177), .B(a[184]), .Z(n7901) );
  NANDN U8104 ( .A(n7901), .B(n42234), .Z(n7861) );
  AND U8105 ( .A(n7862), .B(n7861), .Z(n7910) );
  XNOR U8106 ( .A(n7911), .B(n7910), .Z(n7912) );
  XNOR U8107 ( .A(n7913), .B(n7912), .Z(n7917) );
  NANDN U8108 ( .A(n7864), .B(n7863), .Z(n7868) );
  NAND U8109 ( .A(n7866), .B(n7865), .Z(n7867) );
  AND U8110 ( .A(n7868), .B(n7867), .Z(n7916) );
  XOR U8111 ( .A(n7917), .B(n7916), .Z(n7918) );
  NANDN U8112 ( .A(n7870), .B(n7869), .Z(n7874) );
  NANDN U8113 ( .A(n7872), .B(n7871), .Z(n7873) );
  NAND U8114 ( .A(n7874), .B(n7873), .Z(n7919) );
  XOR U8115 ( .A(n7918), .B(n7919), .Z(n7886) );
  OR U8116 ( .A(n7876), .B(n7875), .Z(n7880) );
  NANDN U8117 ( .A(n7878), .B(n7877), .Z(n7879) );
  NAND U8118 ( .A(n7880), .B(n7879), .Z(n7887) );
  XNOR U8119 ( .A(n7886), .B(n7887), .Z(n7888) );
  XNOR U8120 ( .A(n7889), .B(n7888), .Z(n7922) );
  XNOR U8121 ( .A(n7922), .B(sreg[1206]), .Z(n7924) );
  NAND U8122 ( .A(n7881), .B(sreg[1205]), .Z(n7885) );
  OR U8123 ( .A(n7883), .B(n7882), .Z(n7884) );
  AND U8124 ( .A(n7885), .B(n7884), .Z(n7923) );
  XOR U8125 ( .A(n7924), .B(n7923), .Z(c[1206]) );
  NANDN U8126 ( .A(n7887), .B(n7886), .Z(n7891) );
  NAND U8127 ( .A(n7889), .B(n7888), .Z(n7890) );
  NAND U8128 ( .A(n7891), .B(n7890), .Z(n7930) );
  NAND U8129 ( .A(b[0]), .B(a[191]), .Z(n7892) );
  XNOR U8130 ( .A(b[1]), .B(n7892), .Z(n7894) );
  NAND U8131 ( .A(n42), .B(a[190]), .Z(n7893) );
  AND U8132 ( .A(n7894), .B(n7893), .Z(n7947) );
  XOR U8133 ( .A(a[187]), .B(n42197), .Z(n7936) );
  NANDN U8134 ( .A(n7936), .B(n42173), .Z(n7897) );
  NANDN U8135 ( .A(n7895), .B(n42172), .Z(n7896) );
  NAND U8136 ( .A(n7897), .B(n7896), .Z(n7945) );
  NAND U8137 ( .A(b[7]), .B(a[183]), .Z(n7946) );
  XNOR U8138 ( .A(n7945), .B(n7946), .Z(n7948) );
  XOR U8139 ( .A(n7947), .B(n7948), .Z(n7954) );
  NANDN U8140 ( .A(n7898), .B(n42093), .Z(n7900) );
  XOR U8141 ( .A(n42134), .B(a[189]), .Z(n7939) );
  NANDN U8142 ( .A(n7939), .B(n42095), .Z(n7899) );
  NAND U8143 ( .A(n7900), .B(n7899), .Z(n7952) );
  NANDN U8144 ( .A(n7901), .B(n42231), .Z(n7903) );
  XOR U8145 ( .A(n177), .B(a[185]), .Z(n7942) );
  NANDN U8146 ( .A(n7942), .B(n42234), .Z(n7902) );
  AND U8147 ( .A(n7903), .B(n7902), .Z(n7951) );
  XNOR U8148 ( .A(n7952), .B(n7951), .Z(n7953) );
  XNOR U8149 ( .A(n7954), .B(n7953), .Z(n7958) );
  NANDN U8150 ( .A(n7905), .B(n7904), .Z(n7909) );
  NAND U8151 ( .A(n7907), .B(n7906), .Z(n7908) );
  AND U8152 ( .A(n7909), .B(n7908), .Z(n7957) );
  XOR U8153 ( .A(n7958), .B(n7957), .Z(n7959) );
  NANDN U8154 ( .A(n7911), .B(n7910), .Z(n7915) );
  NANDN U8155 ( .A(n7913), .B(n7912), .Z(n7914) );
  NAND U8156 ( .A(n7915), .B(n7914), .Z(n7960) );
  XOR U8157 ( .A(n7959), .B(n7960), .Z(n7927) );
  OR U8158 ( .A(n7917), .B(n7916), .Z(n7921) );
  NANDN U8159 ( .A(n7919), .B(n7918), .Z(n7920) );
  NAND U8160 ( .A(n7921), .B(n7920), .Z(n7928) );
  XNOR U8161 ( .A(n7927), .B(n7928), .Z(n7929) );
  XNOR U8162 ( .A(n7930), .B(n7929), .Z(n7963) );
  XNOR U8163 ( .A(n7963), .B(sreg[1207]), .Z(n7965) );
  NAND U8164 ( .A(n7922), .B(sreg[1206]), .Z(n7926) );
  OR U8165 ( .A(n7924), .B(n7923), .Z(n7925) );
  AND U8166 ( .A(n7926), .B(n7925), .Z(n7964) );
  XOR U8167 ( .A(n7965), .B(n7964), .Z(c[1207]) );
  NANDN U8168 ( .A(n7928), .B(n7927), .Z(n7932) );
  NAND U8169 ( .A(n7930), .B(n7929), .Z(n7931) );
  NAND U8170 ( .A(n7932), .B(n7931), .Z(n7971) );
  NAND U8171 ( .A(b[0]), .B(a[192]), .Z(n7933) );
  XNOR U8172 ( .A(b[1]), .B(n7933), .Z(n7935) );
  NAND U8173 ( .A(n42), .B(a[191]), .Z(n7934) );
  AND U8174 ( .A(n7935), .B(n7934), .Z(n7988) );
  XOR U8175 ( .A(a[188]), .B(n42197), .Z(n7977) );
  NANDN U8176 ( .A(n7977), .B(n42173), .Z(n7938) );
  NANDN U8177 ( .A(n7936), .B(n42172), .Z(n7937) );
  NAND U8178 ( .A(n7938), .B(n7937), .Z(n7986) );
  NAND U8179 ( .A(b[7]), .B(a[184]), .Z(n7987) );
  XNOR U8180 ( .A(n7986), .B(n7987), .Z(n7989) );
  XOR U8181 ( .A(n7988), .B(n7989), .Z(n7995) );
  NANDN U8182 ( .A(n7939), .B(n42093), .Z(n7941) );
  XOR U8183 ( .A(n42134), .B(a[190]), .Z(n7980) );
  NANDN U8184 ( .A(n7980), .B(n42095), .Z(n7940) );
  NAND U8185 ( .A(n7941), .B(n7940), .Z(n7993) );
  NANDN U8186 ( .A(n7942), .B(n42231), .Z(n7944) );
  XOR U8187 ( .A(n177), .B(a[186]), .Z(n7983) );
  NANDN U8188 ( .A(n7983), .B(n42234), .Z(n7943) );
  AND U8189 ( .A(n7944), .B(n7943), .Z(n7992) );
  XNOR U8190 ( .A(n7993), .B(n7992), .Z(n7994) );
  XNOR U8191 ( .A(n7995), .B(n7994), .Z(n7999) );
  NANDN U8192 ( .A(n7946), .B(n7945), .Z(n7950) );
  NAND U8193 ( .A(n7948), .B(n7947), .Z(n7949) );
  AND U8194 ( .A(n7950), .B(n7949), .Z(n7998) );
  XOR U8195 ( .A(n7999), .B(n7998), .Z(n8000) );
  NANDN U8196 ( .A(n7952), .B(n7951), .Z(n7956) );
  NANDN U8197 ( .A(n7954), .B(n7953), .Z(n7955) );
  NAND U8198 ( .A(n7956), .B(n7955), .Z(n8001) );
  XOR U8199 ( .A(n8000), .B(n8001), .Z(n7968) );
  OR U8200 ( .A(n7958), .B(n7957), .Z(n7962) );
  NANDN U8201 ( .A(n7960), .B(n7959), .Z(n7961) );
  NAND U8202 ( .A(n7962), .B(n7961), .Z(n7969) );
  XNOR U8203 ( .A(n7968), .B(n7969), .Z(n7970) );
  XNOR U8204 ( .A(n7971), .B(n7970), .Z(n8004) );
  XNOR U8205 ( .A(n8004), .B(sreg[1208]), .Z(n8006) );
  NAND U8206 ( .A(n7963), .B(sreg[1207]), .Z(n7967) );
  OR U8207 ( .A(n7965), .B(n7964), .Z(n7966) );
  AND U8208 ( .A(n7967), .B(n7966), .Z(n8005) );
  XOR U8209 ( .A(n8006), .B(n8005), .Z(c[1208]) );
  NANDN U8210 ( .A(n7969), .B(n7968), .Z(n7973) );
  NAND U8211 ( .A(n7971), .B(n7970), .Z(n7972) );
  NAND U8212 ( .A(n7973), .B(n7972), .Z(n8012) );
  NAND U8213 ( .A(b[0]), .B(a[193]), .Z(n7974) );
  XNOR U8214 ( .A(b[1]), .B(n7974), .Z(n7976) );
  NAND U8215 ( .A(n42), .B(a[192]), .Z(n7975) );
  AND U8216 ( .A(n7976), .B(n7975), .Z(n8029) );
  XOR U8217 ( .A(a[189]), .B(n42197), .Z(n8018) );
  NANDN U8218 ( .A(n8018), .B(n42173), .Z(n7979) );
  NANDN U8219 ( .A(n7977), .B(n42172), .Z(n7978) );
  NAND U8220 ( .A(n7979), .B(n7978), .Z(n8027) );
  NAND U8221 ( .A(b[7]), .B(a[185]), .Z(n8028) );
  XNOR U8222 ( .A(n8027), .B(n8028), .Z(n8030) );
  XOR U8223 ( .A(n8029), .B(n8030), .Z(n8036) );
  NANDN U8224 ( .A(n7980), .B(n42093), .Z(n7982) );
  XOR U8225 ( .A(n42134), .B(a[191]), .Z(n8021) );
  NANDN U8226 ( .A(n8021), .B(n42095), .Z(n7981) );
  NAND U8227 ( .A(n7982), .B(n7981), .Z(n8034) );
  NANDN U8228 ( .A(n7983), .B(n42231), .Z(n7985) );
  XOR U8229 ( .A(n177), .B(a[187]), .Z(n8024) );
  NANDN U8230 ( .A(n8024), .B(n42234), .Z(n7984) );
  AND U8231 ( .A(n7985), .B(n7984), .Z(n8033) );
  XNOR U8232 ( .A(n8034), .B(n8033), .Z(n8035) );
  XNOR U8233 ( .A(n8036), .B(n8035), .Z(n8040) );
  NANDN U8234 ( .A(n7987), .B(n7986), .Z(n7991) );
  NAND U8235 ( .A(n7989), .B(n7988), .Z(n7990) );
  AND U8236 ( .A(n7991), .B(n7990), .Z(n8039) );
  XOR U8237 ( .A(n8040), .B(n8039), .Z(n8041) );
  NANDN U8238 ( .A(n7993), .B(n7992), .Z(n7997) );
  NANDN U8239 ( .A(n7995), .B(n7994), .Z(n7996) );
  NAND U8240 ( .A(n7997), .B(n7996), .Z(n8042) );
  XOR U8241 ( .A(n8041), .B(n8042), .Z(n8009) );
  OR U8242 ( .A(n7999), .B(n7998), .Z(n8003) );
  NANDN U8243 ( .A(n8001), .B(n8000), .Z(n8002) );
  NAND U8244 ( .A(n8003), .B(n8002), .Z(n8010) );
  XNOR U8245 ( .A(n8009), .B(n8010), .Z(n8011) );
  XNOR U8246 ( .A(n8012), .B(n8011), .Z(n8045) );
  XNOR U8247 ( .A(n8045), .B(sreg[1209]), .Z(n8047) );
  NAND U8248 ( .A(n8004), .B(sreg[1208]), .Z(n8008) );
  OR U8249 ( .A(n8006), .B(n8005), .Z(n8007) );
  AND U8250 ( .A(n8008), .B(n8007), .Z(n8046) );
  XOR U8251 ( .A(n8047), .B(n8046), .Z(c[1209]) );
  NANDN U8252 ( .A(n8010), .B(n8009), .Z(n8014) );
  NAND U8253 ( .A(n8012), .B(n8011), .Z(n8013) );
  NAND U8254 ( .A(n8014), .B(n8013), .Z(n8053) );
  NAND U8255 ( .A(b[0]), .B(a[194]), .Z(n8015) );
  XNOR U8256 ( .A(b[1]), .B(n8015), .Z(n8017) );
  NAND U8257 ( .A(n42), .B(a[193]), .Z(n8016) );
  AND U8258 ( .A(n8017), .B(n8016), .Z(n8070) );
  XOR U8259 ( .A(a[190]), .B(n42197), .Z(n8059) );
  NANDN U8260 ( .A(n8059), .B(n42173), .Z(n8020) );
  NANDN U8261 ( .A(n8018), .B(n42172), .Z(n8019) );
  NAND U8262 ( .A(n8020), .B(n8019), .Z(n8068) );
  NAND U8263 ( .A(b[7]), .B(a[186]), .Z(n8069) );
  XNOR U8264 ( .A(n8068), .B(n8069), .Z(n8071) );
  XOR U8265 ( .A(n8070), .B(n8071), .Z(n8077) );
  NANDN U8266 ( .A(n8021), .B(n42093), .Z(n8023) );
  XOR U8267 ( .A(n42134), .B(a[192]), .Z(n8062) );
  NANDN U8268 ( .A(n8062), .B(n42095), .Z(n8022) );
  NAND U8269 ( .A(n8023), .B(n8022), .Z(n8075) );
  NANDN U8270 ( .A(n8024), .B(n42231), .Z(n8026) );
  XOR U8271 ( .A(n177), .B(a[188]), .Z(n8065) );
  NANDN U8272 ( .A(n8065), .B(n42234), .Z(n8025) );
  AND U8273 ( .A(n8026), .B(n8025), .Z(n8074) );
  XNOR U8274 ( .A(n8075), .B(n8074), .Z(n8076) );
  XNOR U8275 ( .A(n8077), .B(n8076), .Z(n8081) );
  NANDN U8276 ( .A(n8028), .B(n8027), .Z(n8032) );
  NAND U8277 ( .A(n8030), .B(n8029), .Z(n8031) );
  AND U8278 ( .A(n8032), .B(n8031), .Z(n8080) );
  XOR U8279 ( .A(n8081), .B(n8080), .Z(n8082) );
  NANDN U8280 ( .A(n8034), .B(n8033), .Z(n8038) );
  NANDN U8281 ( .A(n8036), .B(n8035), .Z(n8037) );
  NAND U8282 ( .A(n8038), .B(n8037), .Z(n8083) );
  XOR U8283 ( .A(n8082), .B(n8083), .Z(n8050) );
  OR U8284 ( .A(n8040), .B(n8039), .Z(n8044) );
  NANDN U8285 ( .A(n8042), .B(n8041), .Z(n8043) );
  NAND U8286 ( .A(n8044), .B(n8043), .Z(n8051) );
  XNOR U8287 ( .A(n8050), .B(n8051), .Z(n8052) );
  XNOR U8288 ( .A(n8053), .B(n8052), .Z(n8086) );
  XNOR U8289 ( .A(n8086), .B(sreg[1210]), .Z(n8088) );
  NAND U8290 ( .A(n8045), .B(sreg[1209]), .Z(n8049) );
  OR U8291 ( .A(n8047), .B(n8046), .Z(n8048) );
  AND U8292 ( .A(n8049), .B(n8048), .Z(n8087) );
  XOR U8293 ( .A(n8088), .B(n8087), .Z(c[1210]) );
  NANDN U8294 ( .A(n8051), .B(n8050), .Z(n8055) );
  NAND U8295 ( .A(n8053), .B(n8052), .Z(n8054) );
  NAND U8296 ( .A(n8055), .B(n8054), .Z(n8094) );
  NAND U8297 ( .A(b[0]), .B(a[195]), .Z(n8056) );
  XNOR U8298 ( .A(b[1]), .B(n8056), .Z(n8058) );
  NAND U8299 ( .A(n42), .B(a[194]), .Z(n8057) );
  AND U8300 ( .A(n8058), .B(n8057), .Z(n8111) );
  XOR U8301 ( .A(a[191]), .B(n42197), .Z(n8100) );
  NANDN U8302 ( .A(n8100), .B(n42173), .Z(n8061) );
  NANDN U8303 ( .A(n8059), .B(n42172), .Z(n8060) );
  NAND U8304 ( .A(n8061), .B(n8060), .Z(n8109) );
  NAND U8305 ( .A(b[7]), .B(a[187]), .Z(n8110) );
  XNOR U8306 ( .A(n8109), .B(n8110), .Z(n8112) );
  XOR U8307 ( .A(n8111), .B(n8112), .Z(n8118) );
  NANDN U8308 ( .A(n8062), .B(n42093), .Z(n8064) );
  XOR U8309 ( .A(n42134), .B(a[193]), .Z(n8103) );
  NANDN U8310 ( .A(n8103), .B(n42095), .Z(n8063) );
  NAND U8311 ( .A(n8064), .B(n8063), .Z(n8116) );
  NANDN U8312 ( .A(n8065), .B(n42231), .Z(n8067) );
  XOR U8313 ( .A(n177), .B(a[189]), .Z(n8106) );
  NANDN U8314 ( .A(n8106), .B(n42234), .Z(n8066) );
  AND U8315 ( .A(n8067), .B(n8066), .Z(n8115) );
  XNOR U8316 ( .A(n8116), .B(n8115), .Z(n8117) );
  XNOR U8317 ( .A(n8118), .B(n8117), .Z(n8122) );
  NANDN U8318 ( .A(n8069), .B(n8068), .Z(n8073) );
  NAND U8319 ( .A(n8071), .B(n8070), .Z(n8072) );
  AND U8320 ( .A(n8073), .B(n8072), .Z(n8121) );
  XOR U8321 ( .A(n8122), .B(n8121), .Z(n8123) );
  NANDN U8322 ( .A(n8075), .B(n8074), .Z(n8079) );
  NANDN U8323 ( .A(n8077), .B(n8076), .Z(n8078) );
  NAND U8324 ( .A(n8079), .B(n8078), .Z(n8124) );
  XOR U8325 ( .A(n8123), .B(n8124), .Z(n8091) );
  OR U8326 ( .A(n8081), .B(n8080), .Z(n8085) );
  NANDN U8327 ( .A(n8083), .B(n8082), .Z(n8084) );
  NAND U8328 ( .A(n8085), .B(n8084), .Z(n8092) );
  XNOR U8329 ( .A(n8091), .B(n8092), .Z(n8093) );
  XNOR U8330 ( .A(n8094), .B(n8093), .Z(n8127) );
  XNOR U8331 ( .A(n8127), .B(sreg[1211]), .Z(n8129) );
  NAND U8332 ( .A(n8086), .B(sreg[1210]), .Z(n8090) );
  OR U8333 ( .A(n8088), .B(n8087), .Z(n8089) );
  AND U8334 ( .A(n8090), .B(n8089), .Z(n8128) );
  XOR U8335 ( .A(n8129), .B(n8128), .Z(c[1211]) );
  NANDN U8336 ( .A(n8092), .B(n8091), .Z(n8096) );
  NAND U8337 ( .A(n8094), .B(n8093), .Z(n8095) );
  NAND U8338 ( .A(n8096), .B(n8095), .Z(n8135) );
  NAND U8339 ( .A(b[0]), .B(a[196]), .Z(n8097) );
  XNOR U8340 ( .A(b[1]), .B(n8097), .Z(n8099) );
  NAND U8341 ( .A(n43), .B(a[195]), .Z(n8098) );
  AND U8342 ( .A(n8099), .B(n8098), .Z(n8152) );
  XOR U8343 ( .A(a[192]), .B(n42197), .Z(n8141) );
  NANDN U8344 ( .A(n8141), .B(n42173), .Z(n8102) );
  NANDN U8345 ( .A(n8100), .B(n42172), .Z(n8101) );
  NAND U8346 ( .A(n8102), .B(n8101), .Z(n8150) );
  NAND U8347 ( .A(b[7]), .B(a[188]), .Z(n8151) );
  XNOR U8348 ( .A(n8150), .B(n8151), .Z(n8153) );
  XOR U8349 ( .A(n8152), .B(n8153), .Z(n8159) );
  NANDN U8350 ( .A(n8103), .B(n42093), .Z(n8105) );
  XOR U8351 ( .A(n42134), .B(a[194]), .Z(n8144) );
  NANDN U8352 ( .A(n8144), .B(n42095), .Z(n8104) );
  NAND U8353 ( .A(n8105), .B(n8104), .Z(n8157) );
  NANDN U8354 ( .A(n8106), .B(n42231), .Z(n8108) );
  XOR U8355 ( .A(n177), .B(a[190]), .Z(n8147) );
  NANDN U8356 ( .A(n8147), .B(n42234), .Z(n8107) );
  AND U8357 ( .A(n8108), .B(n8107), .Z(n8156) );
  XNOR U8358 ( .A(n8157), .B(n8156), .Z(n8158) );
  XNOR U8359 ( .A(n8159), .B(n8158), .Z(n8163) );
  NANDN U8360 ( .A(n8110), .B(n8109), .Z(n8114) );
  NAND U8361 ( .A(n8112), .B(n8111), .Z(n8113) );
  AND U8362 ( .A(n8114), .B(n8113), .Z(n8162) );
  XOR U8363 ( .A(n8163), .B(n8162), .Z(n8164) );
  NANDN U8364 ( .A(n8116), .B(n8115), .Z(n8120) );
  NANDN U8365 ( .A(n8118), .B(n8117), .Z(n8119) );
  NAND U8366 ( .A(n8120), .B(n8119), .Z(n8165) );
  XOR U8367 ( .A(n8164), .B(n8165), .Z(n8132) );
  OR U8368 ( .A(n8122), .B(n8121), .Z(n8126) );
  NANDN U8369 ( .A(n8124), .B(n8123), .Z(n8125) );
  NAND U8370 ( .A(n8126), .B(n8125), .Z(n8133) );
  XNOR U8371 ( .A(n8132), .B(n8133), .Z(n8134) );
  XNOR U8372 ( .A(n8135), .B(n8134), .Z(n8168) );
  XNOR U8373 ( .A(n8168), .B(sreg[1212]), .Z(n8170) );
  NAND U8374 ( .A(n8127), .B(sreg[1211]), .Z(n8131) );
  OR U8375 ( .A(n8129), .B(n8128), .Z(n8130) );
  AND U8376 ( .A(n8131), .B(n8130), .Z(n8169) );
  XOR U8377 ( .A(n8170), .B(n8169), .Z(c[1212]) );
  NANDN U8378 ( .A(n8133), .B(n8132), .Z(n8137) );
  NAND U8379 ( .A(n8135), .B(n8134), .Z(n8136) );
  NAND U8380 ( .A(n8137), .B(n8136), .Z(n8176) );
  NAND U8381 ( .A(b[0]), .B(a[197]), .Z(n8138) );
  XNOR U8382 ( .A(b[1]), .B(n8138), .Z(n8140) );
  NAND U8383 ( .A(n43), .B(a[196]), .Z(n8139) );
  AND U8384 ( .A(n8140), .B(n8139), .Z(n8193) );
  XOR U8385 ( .A(a[193]), .B(n42197), .Z(n8182) );
  NANDN U8386 ( .A(n8182), .B(n42173), .Z(n8143) );
  NANDN U8387 ( .A(n8141), .B(n42172), .Z(n8142) );
  NAND U8388 ( .A(n8143), .B(n8142), .Z(n8191) );
  NAND U8389 ( .A(b[7]), .B(a[189]), .Z(n8192) );
  XNOR U8390 ( .A(n8191), .B(n8192), .Z(n8194) );
  XOR U8391 ( .A(n8193), .B(n8194), .Z(n8200) );
  NANDN U8392 ( .A(n8144), .B(n42093), .Z(n8146) );
  XOR U8393 ( .A(n42134), .B(a[195]), .Z(n8185) );
  NANDN U8394 ( .A(n8185), .B(n42095), .Z(n8145) );
  NAND U8395 ( .A(n8146), .B(n8145), .Z(n8198) );
  NANDN U8396 ( .A(n8147), .B(n42231), .Z(n8149) );
  XOR U8397 ( .A(n178), .B(a[191]), .Z(n8188) );
  NANDN U8398 ( .A(n8188), .B(n42234), .Z(n8148) );
  AND U8399 ( .A(n8149), .B(n8148), .Z(n8197) );
  XNOR U8400 ( .A(n8198), .B(n8197), .Z(n8199) );
  XNOR U8401 ( .A(n8200), .B(n8199), .Z(n8204) );
  NANDN U8402 ( .A(n8151), .B(n8150), .Z(n8155) );
  NAND U8403 ( .A(n8153), .B(n8152), .Z(n8154) );
  AND U8404 ( .A(n8155), .B(n8154), .Z(n8203) );
  XOR U8405 ( .A(n8204), .B(n8203), .Z(n8205) );
  NANDN U8406 ( .A(n8157), .B(n8156), .Z(n8161) );
  NANDN U8407 ( .A(n8159), .B(n8158), .Z(n8160) );
  NAND U8408 ( .A(n8161), .B(n8160), .Z(n8206) );
  XOR U8409 ( .A(n8205), .B(n8206), .Z(n8173) );
  OR U8410 ( .A(n8163), .B(n8162), .Z(n8167) );
  NANDN U8411 ( .A(n8165), .B(n8164), .Z(n8166) );
  NAND U8412 ( .A(n8167), .B(n8166), .Z(n8174) );
  XNOR U8413 ( .A(n8173), .B(n8174), .Z(n8175) );
  XNOR U8414 ( .A(n8176), .B(n8175), .Z(n8209) );
  XNOR U8415 ( .A(n8209), .B(sreg[1213]), .Z(n8211) );
  NAND U8416 ( .A(n8168), .B(sreg[1212]), .Z(n8172) );
  OR U8417 ( .A(n8170), .B(n8169), .Z(n8171) );
  AND U8418 ( .A(n8172), .B(n8171), .Z(n8210) );
  XOR U8419 ( .A(n8211), .B(n8210), .Z(c[1213]) );
  NANDN U8420 ( .A(n8174), .B(n8173), .Z(n8178) );
  NAND U8421 ( .A(n8176), .B(n8175), .Z(n8177) );
  NAND U8422 ( .A(n8178), .B(n8177), .Z(n8217) );
  NAND U8423 ( .A(b[0]), .B(a[198]), .Z(n8179) );
  XNOR U8424 ( .A(b[1]), .B(n8179), .Z(n8181) );
  NAND U8425 ( .A(n43), .B(a[197]), .Z(n8180) );
  AND U8426 ( .A(n8181), .B(n8180), .Z(n8234) );
  XOR U8427 ( .A(a[194]), .B(n42197), .Z(n8223) );
  NANDN U8428 ( .A(n8223), .B(n42173), .Z(n8184) );
  NANDN U8429 ( .A(n8182), .B(n42172), .Z(n8183) );
  NAND U8430 ( .A(n8184), .B(n8183), .Z(n8232) );
  NAND U8431 ( .A(b[7]), .B(a[190]), .Z(n8233) );
  XNOR U8432 ( .A(n8232), .B(n8233), .Z(n8235) );
  XOR U8433 ( .A(n8234), .B(n8235), .Z(n8241) );
  NANDN U8434 ( .A(n8185), .B(n42093), .Z(n8187) );
  XOR U8435 ( .A(n42134), .B(a[196]), .Z(n8226) );
  NANDN U8436 ( .A(n8226), .B(n42095), .Z(n8186) );
  NAND U8437 ( .A(n8187), .B(n8186), .Z(n8239) );
  NANDN U8438 ( .A(n8188), .B(n42231), .Z(n8190) );
  XOR U8439 ( .A(n178), .B(a[192]), .Z(n8229) );
  NANDN U8440 ( .A(n8229), .B(n42234), .Z(n8189) );
  AND U8441 ( .A(n8190), .B(n8189), .Z(n8238) );
  XNOR U8442 ( .A(n8239), .B(n8238), .Z(n8240) );
  XNOR U8443 ( .A(n8241), .B(n8240), .Z(n8245) );
  NANDN U8444 ( .A(n8192), .B(n8191), .Z(n8196) );
  NAND U8445 ( .A(n8194), .B(n8193), .Z(n8195) );
  AND U8446 ( .A(n8196), .B(n8195), .Z(n8244) );
  XOR U8447 ( .A(n8245), .B(n8244), .Z(n8246) );
  NANDN U8448 ( .A(n8198), .B(n8197), .Z(n8202) );
  NANDN U8449 ( .A(n8200), .B(n8199), .Z(n8201) );
  NAND U8450 ( .A(n8202), .B(n8201), .Z(n8247) );
  XOR U8451 ( .A(n8246), .B(n8247), .Z(n8214) );
  OR U8452 ( .A(n8204), .B(n8203), .Z(n8208) );
  NANDN U8453 ( .A(n8206), .B(n8205), .Z(n8207) );
  NAND U8454 ( .A(n8208), .B(n8207), .Z(n8215) );
  XNOR U8455 ( .A(n8214), .B(n8215), .Z(n8216) );
  XNOR U8456 ( .A(n8217), .B(n8216), .Z(n8250) );
  XNOR U8457 ( .A(n8250), .B(sreg[1214]), .Z(n8252) );
  NAND U8458 ( .A(n8209), .B(sreg[1213]), .Z(n8213) );
  OR U8459 ( .A(n8211), .B(n8210), .Z(n8212) );
  AND U8460 ( .A(n8213), .B(n8212), .Z(n8251) );
  XOR U8461 ( .A(n8252), .B(n8251), .Z(c[1214]) );
  NANDN U8462 ( .A(n8215), .B(n8214), .Z(n8219) );
  NAND U8463 ( .A(n8217), .B(n8216), .Z(n8218) );
  NAND U8464 ( .A(n8219), .B(n8218), .Z(n8258) );
  NAND U8465 ( .A(b[0]), .B(a[199]), .Z(n8220) );
  XNOR U8466 ( .A(b[1]), .B(n8220), .Z(n8222) );
  NAND U8467 ( .A(n43), .B(a[198]), .Z(n8221) );
  AND U8468 ( .A(n8222), .B(n8221), .Z(n8275) );
  XOR U8469 ( .A(a[195]), .B(n42197), .Z(n8264) );
  NANDN U8470 ( .A(n8264), .B(n42173), .Z(n8225) );
  NANDN U8471 ( .A(n8223), .B(n42172), .Z(n8224) );
  NAND U8472 ( .A(n8225), .B(n8224), .Z(n8273) );
  NAND U8473 ( .A(b[7]), .B(a[191]), .Z(n8274) );
  XNOR U8474 ( .A(n8273), .B(n8274), .Z(n8276) );
  XOR U8475 ( .A(n8275), .B(n8276), .Z(n8282) );
  NANDN U8476 ( .A(n8226), .B(n42093), .Z(n8228) );
  XOR U8477 ( .A(n42134), .B(a[197]), .Z(n8267) );
  NANDN U8478 ( .A(n8267), .B(n42095), .Z(n8227) );
  NAND U8479 ( .A(n8228), .B(n8227), .Z(n8280) );
  NANDN U8480 ( .A(n8229), .B(n42231), .Z(n8231) );
  XOR U8481 ( .A(n178), .B(a[193]), .Z(n8270) );
  NANDN U8482 ( .A(n8270), .B(n42234), .Z(n8230) );
  AND U8483 ( .A(n8231), .B(n8230), .Z(n8279) );
  XNOR U8484 ( .A(n8280), .B(n8279), .Z(n8281) );
  XNOR U8485 ( .A(n8282), .B(n8281), .Z(n8286) );
  NANDN U8486 ( .A(n8233), .B(n8232), .Z(n8237) );
  NAND U8487 ( .A(n8235), .B(n8234), .Z(n8236) );
  AND U8488 ( .A(n8237), .B(n8236), .Z(n8285) );
  XOR U8489 ( .A(n8286), .B(n8285), .Z(n8287) );
  NANDN U8490 ( .A(n8239), .B(n8238), .Z(n8243) );
  NANDN U8491 ( .A(n8241), .B(n8240), .Z(n8242) );
  NAND U8492 ( .A(n8243), .B(n8242), .Z(n8288) );
  XOR U8493 ( .A(n8287), .B(n8288), .Z(n8255) );
  OR U8494 ( .A(n8245), .B(n8244), .Z(n8249) );
  NANDN U8495 ( .A(n8247), .B(n8246), .Z(n8248) );
  NAND U8496 ( .A(n8249), .B(n8248), .Z(n8256) );
  XNOR U8497 ( .A(n8255), .B(n8256), .Z(n8257) );
  XNOR U8498 ( .A(n8258), .B(n8257), .Z(n8291) );
  XNOR U8499 ( .A(n8291), .B(sreg[1215]), .Z(n8293) );
  NAND U8500 ( .A(n8250), .B(sreg[1214]), .Z(n8254) );
  OR U8501 ( .A(n8252), .B(n8251), .Z(n8253) );
  AND U8502 ( .A(n8254), .B(n8253), .Z(n8292) );
  XOR U8503 ( .A(n8293), .B(n8292), .Z(c[1215]) );
  NANDN U8504 ( .A(n8256), .B(n8255), .Z(n8260) );
  NAND U8505 ( .A(n8258), .B(n8257), .Z(n8259) );
  NAND U8506 ( .A(n8260), .B(n8259), .Z(n8299) );
  NAND U8507 ( .A(b[0]), .B(a[200]), .Z(n8261) );
  XNOR U8508 ( .A(b[1]), .B(n8261), .Z(n8263) );
  NAND U8509 ( .A(n43), .B(a[199]), .Z(n8262) );
  AND U8510 ( .A(n8263), .B(n8262), .Z(n8316) );
  XOR U8511 ( .A(a[196]), .B(n42197), .Z(n8305) );
  NANDN U8512 ( .A(n8305), .B(n42173), .Z(n8266) );
  NANDN U8513 ( .A(n8264), .B(n42172), .Z(n8265) );
  NAND U8514 ( .A(n8266), .B(n8265), .Z(n8314) );
  NAND U8515 ( .A(b[7]), .B(a[192]), .Z(n8315) );
  XNOR U8516 ( .A(n8314), .B(n8315), .Z(n8317) );
  XOR U8517 ( .A(n8316), .B(n8317), .Z(n8323) );
  NANDN U8518 ( .A(n8267), .B(n42093), .Z(n8269) );
  XOR U8519 ( .A(n42134), .B(a[198]), .Z(n8308) );
  NANDN U8520 ( .A(n8308), .B(n42095), .Z(n8268) );
  NAND U8521 ( .A(n8269), .B(n8268), .Z(n8321) );
  NANDN U8522 ( .A(n8270), .B(n42231), .Z(n8272) );
  XOR U8523 ( .A(n178), .B(a[194]), .Z(n8311) );
  NANDN U8524 ( .A(n8311), .B(n42234), .Z(n8271) );
  AND U8525 ( .A(n8272), .B(n8271), .Z(n8320) );
  XNOR U8526 ( .A(n8321), .B(n8320), .Z(n8322) );
  XNOR U8527 ( .A(n8323), .B(n8322), .Z(n8327) );
  NANDN U8528 ( .A(n8274), .B(n8273), .Z(n8278) );
  NAND U8529 ( .A(n8276), .B(n8275), .Z(n8277) );
  AND U8530 ( .A(n8278), .B(n8277), .Z(n8326) );
  XOR U8531 ( .A(n8327), .B(n8326), .Z(n8328) );
  NANDN U8532 ( .A(n8280), .B(n8279), .Z(n8284) );
  NANDN U8533 ( .A(n8282), .B(n8281), .Z(n8283) );
  NAND U8534 ( .A(n8284), .B(n8283), .Z(n8329) );
  XOR U8535 ( .A(n8328), .B(n8329), .Z(n8296) );
  OR U8536 ( .A(n8286), .B(n8285), .Z(n8290) );
  NANDN U8537 ( .A(n8288), .B(n8287), .Z(n8289) );
  NAND U8538 ( .A(n8290), .B(n8289), .Z(n8297) );
  XNOR U8539 ( .A(n8296), .B(n8297), .Z(n8298) );
  XNOR U8540 ( .A(n8299), .B(n8298), .Z(n8332) );
  XNOR U8541 ( .A(n8332), .B(sreg[1216]), .Z(n8334) );
  NAND U8542 ( .A(n8291), .B(sreg[1215]), .Z(n8295) );
  OR U8543 ( .A(n8293), .B(n8292), .Z(n8294) );
  AND U8544 ( .A(n8295), .B(n8294), .Z(n8333) );
  XOR U8545 ( .A(n8334), .B(n8333), .Z(c[1216]) );
  NANDN U8546 ( .A(n8297), .B(n8296), .Z(n8301) );
  NAND U8547 ( .A(n8299), .B(n8298), .Z(n8300) );
  NAND U8548 ( .A(n8301), .B(n8300), .Z(n8340) );
  NAND U8549 ( .A(b[0]), .B(a[201]), .Z(n8302) );
  XNOR U8550 ( .A(b[1]), .B(n8302), .Z(n8304) );
  NAND U8551 ( .A(n43), .B(a[200]), .Z(n8303) );
  AND U8552 ( .A(n8304), .B(n8303), .Z(n8357) );
  XOR U8553 ( .A(a[197]), .B(n42197), .Z(n8346) );
  NANDN U8554 ( .A(n8346), .B(n42173), .Z(n8307) );
  NANDN U8555 ( .A(n8305), .B(n42172), .Z(n8306) );
  NAND U8556 ( .A(n8307), .B(n8306), .Z(n8355) );
  NAND U8557 ( .A(b[7]), .B(a[193]), .Z(n8356) );
  XNOR U8558 ( .A(n8355), .B(n8356), .Z(n8358) );
  XOR U8559 ( .A(n8357), .B(n8358), .Z(n8364) );
  NANDN U8560 ( .A(n8308), .B(n42093), .Z(n8310) );
  XOR U8561 ( .A(n42134), .B(a[199]), .Z(n8349) );
  NANDN U8562 ( .A(n8349), .B(n42095), .Z(n8309) );
  NAND U8563 ( .A(n8310), .B(n8309), .Z(n8362) );
  NANDN U8564 ( .A(n8311), .B(n42231), .Z(n8313) );
  XOR U8565 ( .A(n178), .B(a[195]), .Z(n8352) );
  NANDN U8566 ( .A(n8352), .B(n42234), .Z(n8312) );
  AND U8567 ( .A(n8313), .B(n8312), .Z(n8361) );
  XNOR U8568 ( .A(n8362), .B(n8361), .Z(n8363) );
  XNOR U8569 ( .A(n8364), .B(n8363), .Z(n8368) );
  NANDN U8570 ( .A(n8315), .B(n8314), .Z(n8319) );
  NAND U8571 ( .A(n8317), .B(n8316), .Z(n8318) );
  AND U8572 ( .A(n8319), .B(n8318), .Z(n8367) );
  XOR U8573 ( .A(n8368), .B(n8367), .Z(n8369) );
  NANDN U8574 ( .A(n8321), .B(n8320), .Z(n8325) );
  NANDN U8575 ( .A(n8323), .B(n8322), .Z(n8324) );
  NAND U8576 ( .A(n8325), .B(n8324), .Z(n8370) );
  XOR U8577 ( .A(n8369), .B(n8370), .Z(n8337) );
  OR U8578 ( .A(n8327), .B(n8326), .Z(n8331) );
  NANDN U8579 ( .A(n8329), .B(n8328), .Z(n8330) );
  NAND U8580 ( .A(n8331), .B(n8330), .Z(n8338) );
  XNOR U8581 ( .A(n8337), .B(n8338), .Z(n8339) );
  XNOR U8582 ( .A(n8340), .B(n8339), .Z(n8373) );
  XNOR U8583 ( .A(n8373), .B(sreg[1217]), .Z(n8375) );
  NAND U8584 ( .A(n8332), .B(sreg[1216]), .Z(n8336) );
  OR U8585 ( .A(n8334), .B(n8333), .Z(n8335) );
  AND U8586 ( .A(n8336), .B(n8335), .Z(n8374) );
  XOR U8587 ( .A(n8375), .B(n8374), .Z(c[1217]) );
  NANDN U8588 ( .A(n8338), .B(n8337), .Z(n8342) );
  NAND U8589 ( .A(n8340), .B(n8339), .Z(n8341) );
  NAND U8590 ( .A(n8342), .B(n8341), .Z(n8381) );
  NAND U8591 ( .A(b[0]), .B(a[202]), .Z(n8343) );
  XNOR U8592 ( .A(b[1]), .B(n8343), .Z(n8345) );
  NAND U8593 ( .A(n43), .B(a[201]), .Z(n8344) );
  AND U8594 ( .A(n8345), .B(n8344), .Z(n8398) );
  XOR U8595 ( .A(a[198]), .B(n42197), .Z(n8387) );
  NANDN U8596 ( .A(n8387), .B(n42173), .Z(n8348) );
  NANDN U8597 ( .A(n8346), .B(n42172), .Z(n8347) );
  NAND U8598 ( .A(n8348), .B(n8347), .Z(n8396) );
  NAND U8599 ( .A(b[7]), .B(a[194]), .Z(n8397) );
  XNOR U8600 ( .A(n8396), .B(n8397), .Z(n8399) );
  XOR U8601 ( .A(n8398), .B(n8399), .Z(n8405) );
  NANDN U8602 ( .A(n8349), .B(n42093), .Z(n8351) );
  XOR U8603 ( .A(n42134), .B(a[200]), .Z(n8390) );
  NANDN U8604 ( .A(n8390), .B(n42095), .Z(n8350) );
  NAND U8605 ( .A(n8351), .B(n8350), .Z(n8403) );
  NANDN U8606 ( .A(n8352), .B(n42231), .Z(n8354) );
  XOR U8607 ( .A(n178), .B(a[196]), .Z(n8393) );
  NANDN U8608 ( .A(n8393), .B(n42234), .Z(n8353) );
  AND U8609 ( .A(n8354), .B(n8353), .Z(n8402) );
  XNOR U8610 ( .A(n8403), .B(n8402), .Z(n8404) );
  XNOR U8611 ( .A(n8405), .B(n8404), .Z(n8409) );
  NANDN U8612 ( .A(n8356), .B(n8355), .Z(n8360) );
  NAND U8613 ( .A(n8358), .B(n8357), .Z(n8359) );
  AND U8614 ( .A(n8360), .B(n8359), .Z(n8408) );
  XOR U8615 ( .A(n8409), .B(n8408), .Z(n8410) );
  NANDN U8616 ( .A(n8362), .B(n8361), .Z(n8366) );
  NANDN U8617 ( .A(n8364), .B(n8363), .Z(n8365) );
  NAND U8618 ( .A(n8366), .B(n8365), .Z(n8411) );
  XOR U8619 ( .A(n8410), .B(n8411), .Z(n8378) );
  OR U8620 ( .A(n8368), .B(n8367), .Z(n8372) );
  NANDN U8621 ( .A(n8370), .B(n8369), .Z(n8371) );
  NAND U8622 ( .A(n8372), .B(n8371), .Z(n8379) );
  XNOR U8623 ( .A(n8378), .B(n8379), .Z(n8380) );
  XNOR U8624 ( .A(n8381), .B(n8380), .Z(n8414) );
  XNOR U8625 ( .A(n8414), .B(sreg[1218]), .Z(n8416) );
  NAND U8626 ( .A(n8373), .B(sreg[1217]), .Z(n8377) );
  OR U8627 ( .A(n8375), .B(n8374), .Z(n8376) );
  AND U8628 ( .A(n8377), .B(n8376), .Z(n8415) );
  XOR U8629 ( .A(n8416), .B(n8415), .Z(c[1218]) );
  NANDN U8630 ( .A(n8379), .B(n8378), .Z(n8383) );
  NAND U8631 ( .A(n8381), .B(n8380), .Z(n8382) );
  NAND U8632 ( .A(n8383), .B(n8382), .Z(n8422) );
  NAND U8633 ( .A(b[0]), .B(a[203]), .Z(n8384) );
  XNOR U8634 ( .A(b[1]), .B(n8384), .Z(n8386) );
  NAND U8635 ( .A(n44), .B(a[202]), .Z(n8385) );
  AND U8636 ( .A(n8386), .B(n8385), .Z(n8439) );
  XOR U8637 ( .A(a[199]), .B(n42197), .Z(n8428) );
  NANDN U8638 ( .A(n8428), .B(n42173), .Z(n8389) );
  NANDN U8639 ( .A(n8387), .B(n42172), .Z(n8388) );
  NAND U8640 ( .A(n8389), .B(n8388), .Z(n8437) );
  NAND U8641 ( .A(b[7]), .B(a[195]), .Z(n8438) );
  XNOR U8642 ( .A(n8437), .B(n8438), .Z(n8440) );
  XOR U8643 ( .A(n8439), .B(n8440), .Z(n8446) );
  NANDN U8644 ( .A(n8390), .B(n42093), .Z(n8392) );
  XOR U8645 ( .A(n42134), .B(a[201]), .Z(n8431) );
  NANDN U8646 ( .A(n8431), .B(n42095), .Z(n8391) );
  NAND U8647 ( .A(n8392), .B(n8391), .Z(n8444) );
  NANDN U8648 ( .A(n8393), .B(n42231), .Z(n8395) );
  XOR U8649 ( .A(n178), .B(a[197]), .Z(n8434) );
  NANDN U8650 ( .A(n8434), .B(n42234), .Z(n8394) );
  AND U8651 ( .A(n8395), .B(n8394), .Z(n8443) );
  XNOR U8652 ( .A(n8444), .B(n8443), .Z(n8445) );
  XNOR U8653 ( .A(n8446), .B(n8445), .Z(n8450) );
  NANDN U8654 ( .A(n8397), .B(n8396), .Z(n8401) );
  NAND U8655 ( .A(n8399), .B(n8398), .Z(n8400) );
  AND U8656 ( .A(n8401), .B(n8400), .Z(n8449) );
  XOR U8657 ( .A(n8450), .B(n8449), .Z(n8451) );
  NANDN U8658 ( .A(n8403), .B(n8402), .Z(n8407) );
  NANDN U8659 ( .A(n8405), .B(n8404), .Z(n8406) );
  NAND U8660 ( .A(n8407), .B(n8406), .Z(n8452) );
  XOR U8661 ( .A(n8451), .B(n8452), .Z(n8419) );
  OR U8662 ( .A(n8409), .B(n8408), .Z(n8413) );
  NANDN U8663 ( .A(n8411), .B(n8410), .Z(n8412) );
  NAND U8664 ( .A(n8413), .B(n8412), .Z(n8420) );
  XNOR U8665 ( .A(n8419), .B(n8420), .Z(n8421) );
  XNOR U8666 ( .A(n8422), .B(n8421), .Z(n8455) );
  XNOR U8667 ( .A(n8455), .B(sreg[1219]), .Z(n8457) );
  NAND U8668 ( .A(n8414), .B(sreg[1218]), .Z(n8418) );
  OR U8669 ( .A(n8416), .B(n8415), .Z(n8417) );
  AND U8670 ( .A(n8418), .B(n8417), .Z(n8456) );
  XOR U8671 ( .A(n8457), .B(n8456), .Z(c[1219]) );
  NANDN U8672 ( .A(n8420), .B(n8419), .Z(n8424) );
  NAND U8673 ( .A(n8422), .B(n8421), .Z(n8423) );
  NAND U8674 ( .A(n8424), .B(n8423), .Z(n8463) );
  NAND U8675 ( .A(b[0]), .B(a[204]), .Z(n8425) );
  XNOR U8676 ( .A(b[1]), .B(n8425), .Z(n8427) );
  NAND U8677 ( .A(n44), .B(a[203]), .Z(n8426) );
  AND U8678 ( .A(n8427), .B(n8426), .Z(n8480) );
  XOR U8679 ( .A(a[200]), .B(n42197), .Z(n8469) );
  NANDN U8680 ( .A(n8469), .B(n42173), .Z(n8430) );
  NANDN U8681 ( .A(n8428), .B(n42172), .Z(n8429) );
  NAND U8682 ( .A(n8430), .B(n8429), .Z(n8478) );
  NAND U8683 ( .A(b[7]), .B(a[196]), .Z(n8479) );
  XNOR U8684 ( .A(n8478), .B(n8479), .Z(n8481) );
  XOR U8685 ( .A(n8480), .B(n8481), .Z(n8487) );
  NANDN U8686 ( .A(n8431), .B(n42093), .Z(n8433) );
  XOR U8687 ( .A(n42134), .B(a[202]), .Z(n8472) );
  NANDN U8688 ( .A(n8472), .B(n42095), .Z(n8432) );
  NAND U8689 ( .A(n8433), .B(n8432), .Z(n8485) );
  NANDN U8690 ( .A(n8434), .B(n42231), .Z(n8436) );
  XOR U8691 ( .A(n178), .B(a[198]), .Z(n8475) );
  NANDN U8692 ( .A(n8475), .B(n42234), .Z(n8435) );
  AND U8693 ( .A(n8436), .B(n8435), .Z(n8484) );
  XNOR U8694 ( .A(n8485), .B(n8484), .Z(n8486) );
  XNOR U8695 ( .A(n8487), .B(n8486), .Z(n8491) );
  NANDN U8696 ( .A(n8438), .B(n8437), .Z(n8442) );
  NAND U8697 ( .A(n8440), .B(n8439), .Z(n8441) );
  AND U8698 ( .A(n8442), .B(n8441), .Z(n8490) );
  XOR U8699 ( .A(n8491), .B(n8490), .Z(n8492) );
  NANDN U8700 ( .A(n8444), .B(n8443), .Z(n8448) );
  NANDN U8701 ( .A(n8446), .B(n8445), .Z(n8447) );
  NAND U8702 ( .A(n8448), .B(n8447), .Z(n8493) );
  XOR U8703 ( .A(n8492), .B(n8493), .Z(n8460) );
  OR U8704 ( .A(n8450), .B(n8449), .Z(n8454) );
  NANDN U8705 ( .A(n8452), .B(n8451), .Z(n8453) );
  NAND U8706 ( .A(n8454), .B(n8453), .Z(n8461) );
  XNOR U8707 ( .A(n8460), .B(n8461), .Z(n8462) );
  XNOR U8708 ( .A(n8463), .B(n8462), .Z(n8496) );
  XNOR U8709 ( .A(n8496), .B(sreg[1220]), .Z(n8498) );
  NAND U8710 ( .A(n8455), .B(sreg[1219]), .Z(n8459) );
  OR U8711 ( .A(n8457), .B(n8456), .Z(n8458) );
  AND U8712 ( .A(n8459), .B(n8458), .Z(n8497) );
  XOR U8713 ( .A(n8498), .B(n8497), .Z(c[1220]) );
  NANDN U8714 ( .A(n8461), .B(n8460), .Z(n8465) );
  NAND U8715 ( .A(n8463), .B(n8462), .Z(n8464) );
  NAND U8716 ( .A(n8465), .B(n8464), .Z(n8504) );
  NAND U8717 ( .A(b[0]), .B(a[205]), .Z(n8466) );
  XNOR U8718 ( .A(b[1]), .B(n8466), .Z(n8468) );
  NAND U8719 ( .A(n44), .B(a[204]), .Z(n8467) );
  AND U8720 ( .A(n8468), .B(n8467), .Z(n8521) );
  XOR U8721 ( .A(a[201]), .B(n42197), .Z(n8510) );
  NANDN U8722 ( .A(n8510), .B(n42173), .Z(n8471) );
  NANDN U8723 ( .A(n8469), .B(n42172), .Z(n8470) );
  NAND U8724 ( .A(n8471), .B(n8470), .Z(n8519) );
  NAND U8725 ( .A(b[7]), .B(a[197]), .Z(n8520) );
  XNOR U8726 ( .A(n8519), .B(n8520), .Z(n8522) );
  XOR U8727 ( .A(n8521), .B(n8522), .Z(n8528) );
  NANDN U8728 ( .A(n8472), .B(n42093), .Z(n8474) );
  XOR U8729 ( .A(n42134), .B(a[203]), .Z(n8513) );
  NANDN U8730 ( .A(n8513), .B(n42095), .Z(n8473) );
  NAND U8731 ( .A(n8474), .B(n8473), .Z(n8526) );
  NANDN U8732 ( .A(n8475), .B(n42231), .Z(n8477) );
  XOR U8733 ( .A(n178), .B(a[199]), .Z(n8516) );
  NANDN U8734 ( .A(n8516), .B(n42234), .Z(n8476) );
  AND U8735 ( .A(n8477), .B(n8476), .Z(n8525) );
  XNOR U8736 ( .A(n8526), .B(n8525), .Z(n8527) );
  XNOR U8737 ( .A(n8528), .B(n8527), .Z(n8532) );
  NANDN U8738 ( .A(n8479), .B(n8478), .Z(n8483) );
  NAND U8739 ( .A(n8481), .B(n8480), .Z(n8482) );
  AND U8740 ( .A(n8483), .B(n8482), .Z(n8531) );
  XOR U8741 ( .A(n8532), .B(n8531), .Z(n8533) );
  NANDN U8742 ( .A(n8485), .B(n8484), .Z(n8489) );
  NANDN U8743 ( .A(n8487), .B(n8486), .Z(n8488) );
  NAND U8744 ( .A(n8489), .B(n8488), .Z(n8534) );
  XOR U8745 ( .A(n8533), .B(n8534), .Z(n8501) );
  OR U8746 ( .A(n8491), .B(n8490), .Z(n8495) );
  NANDN U8747 ( .A(n8493), .B(n8492), .Z(n8494) );
  NAND U8748 ( .A(n8495), .B(n8494), .Z(n8502) );
  XNOR U8749 ( .A(n8501), .B(n8502), .Z(n8503) );
  XNOR U8750 ( .A(n8504), .B(n8503), .Z(n8537) );
  XNOR U8751 ( .A(n8537), .B(sreg[1221]), .Z(n8539) );
  NAND U8752 ( .A(n8496), .B(sreg[1220]), .Z(n8500) );
  OR U8753 ( .A(n8498), .B(n8497), .Z(n8499) );
  AND U8754 ( .A(n8500), .B(n8499), .Z(n8538) );
  XOR U8755 ( .A(n8539), .B(n8538), .Z(c[1221]) );
  NANDN U8756 ( .A(n8502), .B(n8501), .Z(n8506) );
  NAND U8757 ( .A(n8504), .B(n8503), .Z(n8505) );
  NAND U8758 ( .A(n8506), .B(n8505), .Z(n8545) );
  NAND U8759 ( .A(b[0]), .B(a[206]), .Z(n8507) );
  XNOR U8760 ( .A(b[1]), .B(n8507), .Z(n8509) );
  NAND U8761 ( .A(n44), .B(a[205]), .Z(n8508) );
  AND U8762 ( .A(n8509), .B(n8508), .Z(n8562) );
  XOR U8763 ( .A(a[202]), .B(n42197), .Z(n8551) );
  NANDN U8764 ( .A(n8551), .B(n42173), .Z(n8512) );
  NANDN U8765 ( .A(n8510), .B(n42172), .Z(n8511) );
  NAND U8766 ( .A(n8512), .B(n8511), .Z(n8560) );
  NAND U8767 ( .A(b[7]), .B(a[198]), .Z(n8561) );
  XNOR U8768 ( .A(n8560), .B(n8561), .Z(n8563) );
  XOR U8769 ( .A(n8562), .B(n8563), .Z(n8569) );
  NANDN U8770 ( .A(n8513), .B(n42093), .Z(n8515) );
  XOR U8771 ( .A(n42134), .B(a[204]), .Z(n8554) );
  NANDN U8772 ( .A(n8554), .B(n42095), .Z(n8514) );
  NAND U8773 ( .A(n8515), .B(n8514), .Z(n8567) );
  NANDN U8774 ( .A(n8516), .B(n42231), .Z(n8518) );
  XOR U8775 ( .A(n178), .B(a[200]), .Z(n8557) );
  NANDN U8776 ( .A(n8557), .B(n42234), .Z(n8517) );
  AND U8777 ( .A(n8518), .B(n8517), .Z(n8566) );
  XNOR U8778 ( .A(n8567), .B(n8566), .Z(n8568) );
  XNOR U8779 ( .A(n8569), .B(n8568), .Z(n8573) );
  NANDN U8780 ( .A(n8520), .B(n8519), .Z(n8524) );
  NAND U8781 ( .A(n8522), .B(n8521), .Z(n8523) );
  AND U8782 ( .A(n8524), .B(n8523), .Z(n8572) );
  XOR U8783 ( .A(n8573), .B(n8572), .Z(n8574) );
  NANDN U8784 ( .A(n8526), .B(n8525), .Z(n8530) );
  NANDN U8785 ( .A(n8528), .B(n8527), .Z(n8529) );
  NAND U8786 ( .A(n8530), .B(n8529), .Z(n8575) );
  XOR U8787 ( .A(n8574), .B(n8575), .Z(n8542) );
  OR U8788 ( .A(n8532), .B(n8531), .Z(n8536) );
  NANDN U8789 ( .A(n8534), .B(n8533), .Z(n8535) );
  NAND U8790 ( .A(n8536), .B(n8535), .Z(n8543) );
  XNOR U8791 ( .A(n8542), .B(n8543), .Z(n8544) );
  XNOR U8792 ( .A(n8545), .B(n8544), .Z(n8578) );
  XNOR U8793 ( .A(n8578), .B(sreg[1222]), .Z(n8580) );
  NAND U8794 ( .A(n8537), .B(sreg[1221]), .Z(n8541) );
  OR U8795 ( .A(n8539), .B(n8538), .Z(n8540) );
  AND U8796 ( .A(n8541), .B(n8540), .Z(n8579) );
  XOR U8797 ( .A(n8580), .B(n8579), .Z(c[1222]) );
  NANDN U8798 ( .A(n8543), .B(n8542), .Z(n8547) );
  NAND U8799 ( .A(n8545), .B(n8544), .Z(n8546) );
  NAND U8800 ( .A(n8547), .B(n8546), .Z(n8586) );
  NAND U8801 ( .A(b[0]), .B(a[207]), .Z(n8548) );
  XNOR U8802 ( .A(b[1]), .B(n8548), .Z(n8550) );
  NAND U8803 ( .A(n44), .B(a[206]), .Z(n8549) );
  AND U8804 ( .A(n8550), .B(n8549), .Z(n8603) );
  XOR U8805 ( .A(a[203]), .B(n42197), .Z(n8592) );
  NANDN U8806 ( .A(n8592), .B(n42173), .Z(n8553) );
  NANDN U8807 ( .A(n8551), .B(n42172), .Z(n8552) );
  NAND U8808 ( .A(n8553), .B(n8552), .Z(n8601) );
  NAND U8809 ( .A(b[7]), .B(a[199]), .Z(n8602) );
  XNOR U8810 ( .A(n8601), .B(n8602), .Z(n8604) );
  XOR U8811 ( .A(n8603), .B(n8604), .Z(n8610) );
  NANDN U8812 ( .A(n8554), .B(n42093), .Z(n8556) );
  XOR U8813 ( .A(n42134), .B(a[205]), .Z(n8595) );
  NANDN U8814 ( .A(n8595), .B(n42095), .Z(n8555) );
  NAND U8815 ( .A(n8556), .B(n8555), .Z(n8608) );
  NANDN U8816 ( .A(n8557), .B(n42231), .Z(n8559) );
  XOR U8817 ( .A(n178), .B(a[201]), .Z(n8598) );
  NANDN U8818 ( .A(n8598), .B(n42234), .Z(n8558) );
  AND U8819 ( .A(n8559), .B(n8558), .Z(n8607) );
  XNOR U8820 ( .A(n8608), .B(n8607), .Z(n8609) );
  XNOR U8821 ( .A(n8610), .B(n8609), .Z(n8614) );
  NANDN U8822 ( .A(n8561), .B(n8560), .Z(n8565) );
  NAND U8823 ( .A(n8563), .B(n8562), .Z(n8564) );
  AND U8824 ( .A(n8565), .B(n8564), .Z(n8613) );
  XOR U8825 ( .A(n8614), .B(n8613), .Z(n8615) );
  NANDN U8826 ( .A(n8567), .B(n8566), .Z(n8571) );
  NANDN U8827 ( .A(n8569), .B(n8568), .Z(n8570) );
  NAND U8828 ( .A(n8571), .B(n8570), .Z(n8616) );
  XOR U8829 ( .A(n8615), .B(n8616), .Z(n8583) );
  OR U8830 ( .A(n8573), .B(n8572), .Z(n8577) );
  NANDN U8831 ( .A(n8575), .B(n8574), .Z(n8576) );
  NAND U8832 ( .A(n8577), .B(n8576), .Z(n8584) );
  XNOR U8833 ( .A(n8583), .B(n8584), .Z(n8585) );
  XNOR U8834 ( .A(n8586), .B(n8585), .Z(n8619) );
  XNOR U8835 ( .A(n8619), .B(sreg[1223]), .Z(n8621) );
  NAND U8836 ( .A(n8578), .B(sreg[1222]), .Z(n8582) );
  OR U8837 ( .A(n8580), .B(n8579), .Z(n8581) );
  AND U8838 ( .A(n8582), .B(n8581), .Z(n8620) );
  XOR U8839 ( .A(n8621), .B(n8620), .Z(c[1223]) );
  NANDN U8840 ( .A(n8584), .B(n8583), .Z(n8588) );
  NAND U8841 ( .A(n8586), .B(n8585), .Z(n8587) );
  NAND U8842 ( .A(n8588), .B(n8587), .Z(n8627) );
  NAND U8843 ( .A(b[0]), .B(a[208]), .Z(n8589) );
  XNOR U8844 ( .A(b[1]), .B(n8589), .Z(n8591) );
  NAND U8845 ( .A(n44), .B(a[207]), .Z(n8590) );
  AND U8846 ( .A(n8591), .B(n8590), .Z(n8644) );
  XOR U8847 ( .A(a[204]), .B(n42197), .Z(n8633) );
  NANDN U8848 ( .A(n8633), .B(n42173), .Z(n8594) );
  NANDN U8849 ( .A(n8592), .B(n42172), .Z(n8593) );
  NAND U8850 ( .A(n8594), .B(n8593), .Z(n8642) );
  NAND U8851 ( .A(b[7]), .B(a[200]), .Z(n8643) );
  XNOR U8852 ( .A(n8642), .B(n8643), .Z(n8645) );
  XOR U8853 ( .A(n8644), .B(n8645), .Z(n8651) );
  NANDN U8854 ( .A(n8595), .B(n42093), .Z(n8597) );
  XOR U8855 ( .A(n42134), .B(a[206]), .Z(n8636) );
  NANDN U8856 ( .A(n8636), .B(n42095), .Z(n8596) );
  NAND U8857 ( .A(n8597), .B(n8596), .Z(n8649) );
  NANDN U8858 ( .A(n8598), .B(n42231), .Z(n8600) );
  XOR U8859 ( .A(n178), .B(a[202]), .Z(n8639) );
  NANDN U8860 ( .A(n8639), .B(n42234), .Z(n8599) );
  AND U8861 ( .A(n8600), .B(n8599), .Z(n8648) );
  XNOR U8862 ( .A(n8649), .B(n8648), .Z(n8650) );
  XNOR U8863 ( .A(n8651), .B(n8650), .Z(n8655) );
  NANDN U8864 ( .A(n8602), .B(n8601), .Z(n8606) );
  NAND U8865 ( .A(n8604), .B(n8603), .Z(n8605) );
  AND U8866 ( .A(n8606), .B(n8605), .Z(n8654) );
  XOR U8867 ( .A(n8655), .B(n8654), .Z(n8656) );
  NANDN U8868 ( .A(n8608), .B(n8607), .Z(n8612) );
  NANDN U8869 ( .A(n8610), .B(n8609), .Z(n8611) );
  NAND U8870 ( .A(n8612), .B(n8611), .Z(n8657) );
  XOR U8871 ( .A(n8656), .B(n8657), .Z(n8624) );
  OR U8872 ( .A(n8614), .B(n8613), .Z(n8618) );
  NANDN U8873 ( .A(n8616), .B(n8615), .Z(n8617) );
  NAND U8874 ( .A(n8618), .B(n8617), .Z(n8625) );
  XNOR U8875 ( .A(n8624), .B(n8625), .Z(n8626) );
  XNOR U8876 ( .A(n8627), .B(n8626), .Z(n8660) );
  XNOR U8877 ( .A(n8660), .B(sreg[1224]), .Z(n8662) );
  NAND U8878 ( .A(n8619), .B(sreg[1223]), .Z(n8623) );
  OR U8879 ( .A(n8621), .B(n8620), .Z(n8622) );
  AND U8880 ( .A(n8623), .B(n8622), .Z(n8661) );
  XOR U8881 ( .A(n8662), .B(n8661), .Z(c[1224]) );
  NANDN U8882 ( .A(n8625), .B(n8624), .Z(n8629) );
  NAND U8883 ( .A(n8627), .B(n8626), .Z(n8628) );
  NAND U8884 ( .A(n8629), .B(n8628), .Z(n8668) );
  NAND U8885 ( .A(b[0]), .B(a[209]), .Z(n8630) );
  XNOR U8886 ( .A(b[1]), .B(n8630), .Z(n8632) );
  NAND U8887 ( .A(n44), .B(a[208]), .Z(n8631) );
  AND U8888 ( .A(n8632), .B(n8631), .Z(n8685) );
  XOR U8889 ( .A(a[205]), .B(n42197), .Z(n8674) );
  NANDN U8890 ( .A(n8674), .B(n42173), .Z(n8635) );
  NANDN U8891 ( .A(n8633), .B(n42172), .Z(n8634) );
  NAND U8892 ( .A(n8635), .B(n8634), .Z(n8683) );
  NAND U8893 ( .A(b[7]), .B(a[201]), .Z(n8684) );
  XNOR U8894 ( .A(n8683), .B(n8684), .Z(n8686) );
  XOR U8895 ( .A(n8685), .B(n8686), .Z(n8692) );
  NANDN U8896 ( .A(n8636), .B(n42093), .Z(n8638) );
  XOR U8897 ( .A(n42134), .B(a[207]), .Z(n8677) );
  NANDN U8898 ( .A(n8677), .B(n42095), .Z(n8637) );
  NAND U8899 ( .A(n8638), .B(n8637), .Z(n8690) );
  NANDN U8900 ( .A(n8639), .B(n42231), .Z(n8641) );
  XOR U8901 ( .A(n179), .B(a[203]), .Z(n8680) );
  NANDN U8902 ( .A(n8680), .B(n42234), .Z(n8640) );
  AND U8903 ( .A(n8641), .B(n8640), .Z(n8689) );
  XNOR U8904 ( .A(n8690), .B(n8689), .Z(n8691) );
  XNOR U8905 ( .A(n8692), .B(n8691), .Z(n8696) );
  NANDN U8906 ( .A(n8643), .B(n8642), .Z(n8647) );
  NAND U8907 ( .A(n8645), .B(n8644), .Z(n8646) );
  AND U8908 ( .A(n8647), .B(n8646), .Z(n8695) );
  XOR U8909 ( .A(n8696), .B(n8695), .Z(n8697) );
  NANDN U8910 ( .A(n8649), .B(n8648), .Z(n8653) );
  NANDN U8911 ( .A(n8651), .B(n8650), .Z(n8652) );
  NAND U8912 ( .A(n8653), .B(n8652), .Z(n8698) );
  XOR U8913 ( .A(n8697), .B(n8698), .Z(n8665) );
  OR U8914 ( .A(n8655), .B(n8654), .Z(n8659) );
  NANDN U8915 ( .A(n8657), .B(n8656), .Z(n8658) );
  NAND U8916 ( .A(n8659), .B(n8658), .Z(n8666) );
  XNOR U8917 ( .A(n8665), .B(n8666), .Z(n8667) );
  XNOR U8918 ( .A(n8668), .B(n8667), .Z(n8701) );
  XNOR U8919 ( .A(n8701), .B(sreg[1225]), .Z(n8703) );
  NAND U8920 ( .A(n8660), .B(sreg[1224]), .Z(n8664) );
  OR U8921 ( .A(n8662), .B(n8661), .Z(n8663) );
  AND U8922 ( .A(n8664), .B(n8663), .Z(n8702) );
  XOR U8923 ( .A(n8703), .B(n8702), .Z(c[1225]) );
  NANDN U8924 ( .A(n8666), .B(n8665), .Z(n8670) );
  NAND U8925 ( .A(n8668), .B(n8667), .Z(n8669) );
  NAND U8926 ( .A(n8670), .B(n8669), .Z(n8709) );
  NAND U8927 ( .A(b[0]), .B(a[210]), .Z(n8671) );
  XNOR U8928 ( .A(b[1]), .B(n8671), .Z(n8673) );
  NAND U8929 ( .A(n45), .B(a[209]), .Z(n8672) );
  AND U8930 ( .A(n8673), .B(n8672), .Z(n8726) );
  XOR U8931 ( .A(a[206]), .B(n42197), .Z(n8715) );
  NANDN U8932 ( .A(n8715), .B(n42173), .Z(n8676) );
  NANDN U8933 ( .A(n8674), .B(n42172), .Z(n8675) );
  NAND U8934 ( .A(n8676), .B(n8675), .Z(n8724) );
  NAND U8935 ( .A(b[7]), .B(a[202]), .Z(n8725) );
  XNOR U8936 ( .A(n8724), .B(n8725), .Z(n8727) );
  XOR U8937 ( .A(n8726), .B(n8727), .Z(n8733) );
  NANDN U8938 ( .A(n8677), .B(n42093), .Z(n8679) );
  XOR U8939 ( .A(n42134), .B(a[208]), .Z(n8718) );
  NANDN U8940 ( .A(n8718), .B(n42095), .Z(n8678) );
  NAND U8941 ( .A(n8679), .B(n8678), .Z(n8731) );
  NANDN U8942 ( .A(n8680), .B(n42231), .Z(n8682) );
  XOR U8943 ( .A(n179), .B(a[204]), .Z(n8721) );
  NANDN U8944 ( .A(n8721), .B(n42234), .Z(n8681) );
  AND U8945 ( .A(n8682), .B(n8681), .Z(n8730) );
  XNOR U8946 ( .A(n8731), .B(n8730), .Z(n8732) );
  XNOR U8947 ( .A(n8733), .B(n8732), .Z(n8737) );
  NANDN U8948 ( .A(n8684), .B(n8683), .Z(n8688) );
  NAND U8949 ( .A(n8686), .B(n8685), .Z(n8687) );
  AND U8950 ( .A(n8688), .B(n8687), .Z(n8736) );
  XOR U8951 ( .A(n8737), .B(n8736), .Z(n8738) );
  NANDN U8952 ( .A(n8690), .B(n8689), .Z(n8694) );
  NANDN U8953 ( .A(n8692), .B(n8691), .Z(n8693) );
  NAND U8954 ( .A(n8694), .B(n8693), .Z(n8739) );
  XOR U8955 ( .A(n8738), .B(n8739), .Z(n8706) );
  OR U8956 ( .A(n8696), .B(n8695), .Z(n8700) );
  NANDN U8957 ( .A(n8698), .B(n8697), .Z(n8699) );
  NAND U8958 ( .A(n8700), .B(n8699), .Z(n8707) );
  XNOR U8959 ( .A(n8706), .B(n8707), .Z(n8708) );
  XNOR U8960 ( .A(n8709), .B(n8708), .Z(n8742) );
  XNOR U8961 ( .A(n8742), .B(sreg[1226]), .Z(n8744) );
  NAND U8962 ( .A(n8701), .B(sreg[1225]), .Z(n8705) );
  OR U8963 ( .A(n8703), .B(n8702), .Z(n8704) );
  AND U8964 ( .A(n8705), .B(n8704), .Z(n8743) );
  XOR U8965 ( .A(n8744), .B(n8743), .Z(c[1226]) );
  NANDN U8966 ( .A(n8707), .B(n8706), .Z(n8711) );
  NAND U8967 ( .A(n8709), .B(n8708), .Z(n8710) );
  NAND U8968 ( .A(n8711), .B(n8710), .Z(n8750) );
  NAND U8969 ( .A(b[0]), .B(a[211]), .Z(n8712) );
  XNOR U8970 ( .A(b[1]), .B(n8712), .Z(n8714) );
  NAND U8971 ( .A(n45), .B(a[210]), .Z(n8713) );
  AND U8972 ( .A(n8714), .B(n8713), .Z(n8767) );
  XOR U8973 ( .A(a[207]), .B(n42197), .Z(n8756) );
  NANDN U8974 ( .A(n8756), .B(n42173), .Z(n8717) );
  NANDN U8975 ( .A(n8715), .B(n42172), .Z(n8716) );
  NAND U8976 ( .A(n8717), .B(n8716), .Z(n8765) );
  NAND U8977 ( .A(b[7]), .B(a[203]), .Z(n8766) );
  XNOR U8978 ( .A(n8765), .B(n8766), .Z(n8768) );
  XOR U8979 ( .A(n8767), .B(n8768), .Z(n8774) );
  NANDN U8980 ( .A(n8718), .B(n42093), .Z(n8720) );
  XOR U8981 ( .A(n42134), .B(a[209]), .Z(n8759) );
  NANDN U8982 ( .A(n8759), .B(n42095), .Z(n8719) );
  NAND U8983 ( .A(n8720), .B(n8719), .Z(n8772) );
  NANDN U8984 ( .A(n8721), .B(n42231), .Z(n8723) );
  XOR U8985 ( .A(n179), .B(a[205]), .Z(n8762) );
  NANDN U8986 ( .A(n8762), .B(n42234), .Z(n8722) );
  AND U8987 ( .A(n8723), .B(n8722), .Z(n8771) );
  XNOR U8988 ( .A(n8772), .B(n8771), .Z(n8773) );
  XNOR U8989 ( .A(n8774), .B(n8773), .Z(n8778) );
  NANDN U8990 ( .A(n8725), .B(n8724), .Z(n8729) );
  NAND U8991 ( .A(n8727), .B(n8726), .Z(n8728) );
  AND U8992 ( .A(n8729), .B(n8728), .Z(n8777) );
  XOR U8993 ( .A(n8778), .B(n8777), .Z(n8779) );
  NANDN U8994 ( .A(n8731), .B(n8730), .Z(n8735) );
  NANDN U8995 ( .A(n8733), .B(n8732), .Z(n8734) );
  NAND U8996 ( .A(n8735), .B(n8734), .Z(n8780) );
  XOR U8997 ( .A(n8779), .B(n8780), .Z(n8747) );
  OR U8998 ( .A(n8737), .B(n8736), .Z(n8741) );
  NANDN U8999 ( .A(n8739), .B(n8738), .Z(n8740) );
  NAND U9000 ( .A(n8741), .B(n8740), .Z(n8748) );
  XNOR U9001 ( .A(n8747), .B(n8748), .Z(n8749) );
  XNOR U9002 ( .A(n8750), .B(n8749), .Z(n8783) );
  XNOR U9003 ( .A(n8783), .B(sreg[1227]), .Z(n8785) );
  NAND U9004 ( .A(n8742), .B(sreg[1226]), .Z(n8746) );
  OR U9005 ( .A(n8744), .B(n8743), .Z(n8745) );
  AND U9006 ( .A(n8746), .B(n8745), .Z(n8784) );
  XOR U9007 ( .A(n8785), .B(n8784), .Z(c[1227]) );
  NANDN U9008 ( .A(n8748), .B(n8747), .Z(n8752) );
  NAND U9009 ( .A(n8750), .B(n8749), .Z(n8751) );
  NAND U9010 ( .A(n8752), .B(n8751), .Z(n8791) );
  NAND U9011 ( .A(b[0]), .B(a[212]), .Z(n8753) );
  XNOR U9012 ( .A(b[1]), .B(n8753), .Z(n8755) );
  NAND U9013 ( .A(n45), .B(a[211]), .Z(n8754) );
  AND U9014 ( .A(n8755), .B(n8754), .Z(n8808) );
  XOR U9015 ( .A(a[208]), .B(n42197), .Z(n8797) );
  NANDN U9016 ( .A(n8797), .B(n42173), .Z(n8758) );
  NANDN U9017 ( .A(n8756), .B(n42172), .Z(n8757) );
  NAND U9018 ( .A(n8758), .B(n8757), .Z(n8806) );
  NAND U9019 ( .A(b[7]), .B(a[204]), .Z(n8807) );
  XNOR U9020 ( .A(n8806), .B(n8807), .Z(n8809) );
  XOR U9021 ( .A(n8808), .B(n8809), .Z(n8815) );
  NANDN U9022 ( .A(n8759), .B(n42093), .Z(n8761) );
  XOR U9023 ( .A(n42134), .B(a[210]), .Z(n8800) );
  NANDN U9024 ( .A(n8800), .B(n42095), .Z(n8760) );
  NAND U9025 ( .A(n8761), .B(n8760), .Z(n8813) );
  NANDN U9026 ( .A(n8762), .B(n42231), .Z(n8764) );
  XOR U9027 ( .A(n179), .B(a[206]), .Z(n8803) );
  NANDN U9028 ( .A(n8803), .B(n42234), .Z(n8763) );
  AND U9029 ( .A(n8764), .B(n8763), .Z(n8812) );
  XNOR U9030 ( .A(n8813), .B(n8812), .Z(n8814) );
  XNOR U9031 ( .A(n8815), .B(n8814), .Z(n8819) );
  NANDN U9032 ( .A(n8766), .B(n8765), .Z(n8770) );
  NAND U9033 ( .A(n8768), .B(n8767), .Z(n8769) );
  AND U9034 ( .A(n8770), .B(n8769), .Z(n8818) );
  XOR U9035 ( .A(n8819), .B(n8818), .Z(n8820) );
  NANDN U9036 ( .A(n8772), .B(n8771), .Z(n8776) );
  NANDN U9037 ( .A(n8774), .B(n8773), .Z(n8775) );
  NAND U9038 ( .A(n8776), .B(n8775), .Z(n8821) );
  XOR U9039 ( .A(n8820), .B(n8821), .Z(n8788) );
  OR U9040 ( .A(n8778), .B(n8777), .Z(n8782) );
  NANDN U9041 ( .A(n8780), .B(n8779), .Z(n8781) );
  NAND U9042 ( .A(n8782), .B(n8781), .Z(n8789) );
  XNOR U9043 ( .A(n8788), .B(n8789), .Z(n8790) );
  XNOR U9044 ( .A(n8791), .B(n8790), .Z(n8824) );
  XNOR U9045 ( .A(n8824), .B(sreg[1228]), .Z(n8826) );
  NAND U9046 ( .A(n8783), .B(sreg[1227]), .Z(n8787) );
  OR U9047 ( .A(n8785), .B(n8784), .Z(n8786) );
  AND U9048 ( .A(n8787), .B(n8786), .Z(n8825) );
  XOR U9049 ( .A(n8826), .B(n8825), .Z(c[1228]) );
  NANDN U9050 ( .A(n8789), .B(n8788), .Z(n8793) );
  NAND U9051 ( .A(n8791), .B(n8790), .Z(n8792) );
  NAND U9052 ( .A(n8793), .B(n8792), .Z(n8832) );
  NAND U9053 ( .A(b[0]), .B(a[213]), .Z(n8794) );
  XNOR U9054 ( .A(b[1]), .B(n8794), .Z(n8796) );
  NAND U9055 ( .A(n45), .B(a[212]), .Z(n8795) );
  AND U9056 ( .A(n8796), .B(n8795), .Z(n8849) );
  XOR U9057 ( .A(a[209]), .B(n42197), .Z(n8838) );
  NANDN U9058 ( .A(n8838), .B(n42173), .Z(n8799) );
  NANDN U9059 ( .A(n8797), .B(n42172), .Z(n8798) );
  NAND U9060 ( .A(n8799), .B(n8798), .Z(n8847) );
  NAND U9061 ( .A(b[7]), .B(a[205]), .Z(n8848) );
  XNOR U9062 ( .A(n8847), .B(n8848), .Z(n8850) );
  XOR U9063 ( .A(n8849), .B(n8850), .Z(n8856) );
  NANDN U9064 ( .A(n8800), .B(n42093), .Z(n8802) );
  XOR U9065 ( .A(n42134), .B(a[211]), .Z(n8841) );
  NANDN U9066 ( .A(n8841), .B(n42095), .Z(n8801) );
  NAND U9067 ( .A(n8802), .B(n8801), .Z(n8854) );
  NANDN U9068 ( .A(n8803), .B(n42231), .Z(n8805) );
  XOR U9069 ( .A(n179), .B(a[207]), .Z(n8844) );
  NANDN U9070 ( .A(n8844), .B(n42234), .Z(n8804) );
  AND U9071 ( .A(n8805), .B(n8804), .Z(n8853) );
  XNOR U9072 ( .A(n8854), .B(n8853), .Z(n8855) );
  XNOR U9073 ( .A(n8856), .B(n8855), .Z(n8860) );
  NANDN U9074 ( .A(n8807), .B(n8806), .Z(n8811) );
  NAND U9075 ( .A(n8809), .B(n8808), .Z(n8810) );
  AND U9076 ( .A(n8811), .B(n8810), .Z(n8859) );
  XOR U9077 ( .A(n8860), .B(n8859), .Z(n8861) );
  NANDN U9078 ( .A(n8813), .B(n8812), .Z(n8817) );
  NANDN U9079 ( .A(n8815), .B(n8814), .Z(n8816) );
  NAND U9080 ( .A(n8817), .B(n8816), .Z(n8862) );
  XOR U9081 ( .A(n8861), .B(n8862), .Z(n8829) );
  OR U9082 ( .A(n8819), .B(n8818), .Z(n8823) );
  NANDN U9083 ( .A(n8821), .B(n8820), .Z(n8822) );
  NAND U9084 ( .A(n8823), .B(n8822), .Z(n8830) );
  XNOR U9085 ( .A(n8829), .B(n8830), .Z(n8831) );
  XNOR U9086 ( .A(n8832), .B(n8831), .Z(n8865) );
  XNOR U9087 ( .A(n8865), .B(sreg[1229]), .Z(n8867) );
  NAND U9088 ( .A(n8824), .B(sreg[1228]), .Z(n8828) );
  OR U9089 ( .A(n8826), .B(n8825), .Z(n8827) );
  AND U9090 ( .A(n8828), .B(n8827), .Z(n8866) );
  XOR U9091 ( .A(n8867), .B(n8866), .Z(c[1229]) );
  NANDN U9092 ( .A(n8830), .B(n8829), .Z(n8834) );
  NAND U9093 ( .A(n8832), .B(n8831), .Z(n8833) );
  NAND U9094 ( .A(n8834), .B(n8833), .Z(n8873) );
  NAND U9095 ( .A(b[0]), .B(a[214]), .Z(n8835) );
  XNOR U9096 ( .A(b[1]), .B(n8835), .Z(n8837) );
  NAND U9097 ( .A(n45), .B(a[213]), .Z(n8836) );
  AND U9098 ( .A(n8837), .B(n8836), .Z(n8890) );
  XOR U9099 ( .A(a[210]), .B(n42197), .Z(n8879) );
  NANDN U9100 ( .A(n8879), .B(n42173), .Z(n8840) );
  NANDN U9101 ( .A(n8838), .B(n42172), .Z(n8839) );
  NAND U9102 ( .A(n8840), .B(n8839), .Z(n8888) );
  NAND U9103 ( .A(b[7]), .B(a[206]), .Z(n8889) );
  XNOR U9104 ( .A(n8888), .B(n8889), .Z(n8891) );
  XOR U9105 ( .A(n8890), .B(n8891), .Z(n8897) );
  NANDN U9106 ( .A(n8841), .B(n42093), .Z(n8843) );
  XOR U9107 ( .A(n42134), .B(a[212]), .Z(n8882) );
  NANDN U9108 ( .A(n8882), .B(n42095), .Z(n8842) );
  NAND U9109 ( .A(n8843), .B(n8842), .Z(n8895) );
  NANDN U9110 ( .A(n8844), .B(n42231), .Z(n8846) );
  XOR U9111 ( .A(n179), .B(a[208]), .Z(n8885) );
  NANDN U9112 ( .A(n8885), .B(n42234), .Z(n8845) );
  AND U9113 ( .A(n8846), .B(n8845), .Z(n8894) );
  XNOR U9114 ( .A(n8895), .B(n8894), .Z(n8896) );
  XNOR U9115 ( .A(n8897), .B(n8896), .Z(n8901) );
  NANDN U9116 ( .A(n8848), .B(n8847), .Z(n8852) );
  NAND U9117 ( .A(n8850), .B(n8849), .Z(n8851) );
  AND U9118 ( .A(n8852), .B(n8851), .Z(n8900) );
  XOR U9119 ( .A(n8901), .B(n8900), .Z(n8902) );
  NANDN U9120 ( .A(n8854), .B(n8853), .Z(n8858) );
  NANDN U9121 ( .A(n8856), .B(n8855), .Z(n8857) );
  NAND U9122 ( .A(n8858), .B(n8857), .Z(n8903) );
  XOR U9123 ( .A(n8902), .B(n8903), .Z(n8870) );
  OR U9124 ( .A(n8860), .B(n8859), .Z(n8864) );
  NANDN U9125 ( .A(n8862), .B(n8861), .Z(n8863) );
  NAND U9126 ( .A(n8864), .B(n8863), .Z(n8871) );
  XNOR U9127 ( .A(n8870), .B(n8871), .Z(n8872) );
  XNOR U9128 ( .A(n8873), .B(n8872), .Z(n8906) );
  XNOR U9129 ( .A(n8906), .B(sreg[1230]), .Z(n8908) );
  NAND U9130 ( .A(n8865), .B(sreg[1229]), .Z(n8869) );
  OR U9131 ( .A(n8867), .B(n8866), .Z(n8868) );
  AND U9132 ( .A(n8869), .B(n8868), .Z(n8907) );
  XOR U9133 ( .A(n8908), .B(n8907), .Z(c[1230]) );
  NANDN U9134 ( .A(n8871), .B(n8870), .Z(n8875) );
  NAND U9135 ( .A(n8873), .B(n8872), .Z(n8874) );
  NAND U9136 ( .A(n8875), .B(n8874), .Z(n8914) );
  NAND U9137 ( .A(b[0]), .B(a[215]), .Z(n8876) );
  XNOR U9138 ( .A(b[1]), .B(n8876), .Z(n8878) );
  NAND U9139 ( .A(n45), .B(a[214]), .Z(n8877) );
  AND U9140 ( .A(n8878), .B(n8877), .Z(n8931) );
  XOR U9141 ( .A(a[211]), .B(n42197), .Z(n8920) );
  NANDN U9142 ( .A(n8920), .B(n42173), .Z(n8881) );
  NANDN U9143 ( .A(n8879), .B(n42172), .Z(n8880) );
  NAND U9144 ( .A(n8881), .B(n8880), .Z(n8929) );
  NAND U9145 ( .A(b[7]), .B(a[207]), .Z(n8930) );
  XNOR U9146 ( .A(n8929), .B(n8930), .Z(n8932) );
  XOR U9147 ( .A(n8931), .B(n8932), .Z(n8938) );
  NANDN U9148 ( .A(n8882), .B(n42093), .Z(n8884) );
  XOR U9149 ( .A(n42134), .B(a[213]), .Z(n8923) );
  NANDN U9150 ( .A(n8923), .B(n42095), .Z(n8883) );
  NAND U9151 ( .A(n8884), .B(n8883), .Z(n8936) );
  NANDN U9152 ( .A(n8885), .B(n42231), .Z(n8887) );
  XOR U9153 ( .A(n179), .B(a[209]), .Z(n8926) );
  NANDN U9154 ( .A(n8926), .B(n42234), .Z(n8886) );
  AND U9155 ( .A(n8887), .B(n8886), .Z(n8935) );
  XNOR U9156 ( .A(n8936), .B(n8935), .Z(n8937) );
  XNOR U9157 ( .A(n8938), .B(n8937), .Z(n8942) );
  NANDN U9158 ( .A(n8889), .B(n8888), .Z(n8893) );
  NAND U9159 ( .A(n8891), .B(n8890), .Z(n8892) );
  AND U9160 ( .A(n8893), .B(n8892), .Z(n8941) );
  XOR U9161 ( .A(n8942), .B(n8941), .Z(n8943) );
  NANDN U9162 ( .A(n8895), .B(n8894), .Z(n8899) );
  NANDN U9163 ( .A(n8897), .B(n8896), .Z(n8898) );
  NAND U9164 ( .A(n8899), .B(n8898), .Z(n8944) );
  XOR U9165 ( .A(n8943), .B(n8944), .Z(n8911) );
  OR U9166 ( .A(n8901), .B(n8900), .Z(n8905) );
  NANDN U9167 ( .A(n8903), .B(n8902), .Z(n8904) );
  NAND U9168 ( .A(n8905), .B(n8904), .Z(n8912) );
  XNOR U9169 ( .A(n8911), .B(n8912), .Z(n8913) );
  XNOR U9170 ( .A(n8914), .B(n8913), .Z(n8947) );
  XNOR U9171 ( .A(n8947), .B(sreg[1231]), .Z(n8949) );
  NAND U9172 ( .A(n8906), .B(sreg[1230]), .Z(n8910) );
  OR U9173 ( .A(n8908), .B(n8907), .Z(n8909) );
  AND U9174 ( .A(n8910), .B(n8909), .Z(n8948) );
  XOR U9175 ( .A(n8949), .B(n8948), .Z(c[1231]) );
  NANDN U9176 ( .A(n8912), .B(n8911), .Z(n8916) );
  NAND U9177 ( .A(n8914), .B(n8913), .Z(n8915) );
  NAND U9178 ( .A(n8916), .B(n8915), .Z(n8955) );
  NAND U9179 ( .A(b[0]), .B(a[216]), .Z(n8917) );
  XNOR U9180 ( .A(b[1]), .B(n8917), .Z(n8919) );
  NAND U9181 ( .A(n45), .B(a[215]), .Z(n8918) );
  AND U9182 ( .A(n8919), .B(n8918), .Z(n8972) );
  XOR U9183 ( .A(a[212]), .B(n42197), .Z(n8961) );
  NANDN U9184 ( .A(n8961), .B(n42173), .Z(n8922) );
  NANDN U9185 ( .A(n8920), .B(n42172), .Z(n8921) );
  NAND U9186 ( .A(n8922), .B(n8921), .Z(n8970) );
  NAND U9187 ( .A(b[7]), .B(a[208]), .Z(n8971) );
  XNOR U9188 ( .A(n8970), .B(n8971), .Z(n8973) );
  XOR U9189 ( .A(n8972), .B(n8973), .Z(n8979) );
  NANDN U9190 ( .A(n8923), .B(n42093), .Z(n8925) );
  XOR U9191 ( .A(n42134), .B(a[214]), .Z(n8964) );
  NANDN U9192 ( .A(n8964), .B(n42095), .Z(n8924) );
  NAND U9193 ( .A(n8925), .B(n8924), .Z(n8977) );
  NANDN U9194 ( .A(n8926), .B(n42231), .Z(n8928) );
  XOR U9195 ( .A(n179), .B(a[210]), .Z(n8967) );
  NANDN U9196 ( .A(n8967), .B(n42234), .Z(n8927) );
  AND U9197 ( .A(n8928), .B(n8927), .Z(n8976) );
  XNOR U9198 ( .A(n8977), .B(n8976), .Z(n8978) );
  XNOR U9199 ( .A(n8979), .B(n8978), .Z(n8983) );
  NANDN U9200 ( .A(n8930), .B(n8929), .Z(n8934) );
  NAND U9201 ( .A(n8932), .B(n8931), .Z(n8933) );
  AND U9202 ( .A(n8934), .B(n8933), .Z(n8982) );
  XOR U9203 ( .A(n8983), .B(n8982), .Z(n8984) );
  NANDN U9204 ( .A(n8936), .B(n8935), .Z(n8940) );
  NANDN U9205 ( .A(n8938), .B(n8937), .Z(n8939) );
  NAND U9206 ( .A(n8940), .B(n8939), .Z(n8985) );
  XOR U9207 ( .A(n8984), .B(n8985), .Z(n8952) );
  OR U9208 ( .A(n8942), .B(n8941), .Z(n8946) );
  NANDN U9209 ( .A(n8944), .B(n8943), .Z(n8945) );
  NAND U9210 ( .A(n8946), .B(n8945), .Z(n8953) );
  XNOR U9211 ( .A(n8952), .B(n8953), .Z(n8954) );
  XNOR U9212 ( .A(n8955), .B(n8954), .Z(n8988) );
  XNOR U9213 ( .A(n8988), .B(sreg[1232]), .Z(n8990) );
  NAND U9214 ( .A(n8947), .B(sreg[1231]), .Z(n8951) );
  OR U9215 ( .A(n8949), .B(n8948), .Z(n8950) );
  AND U9216 ( .A(n8951), .B(n8950), .Z(n8989) );
  XOR U9217 ( .A(n8990), .B(n8989), .Z(c[1232]) );
  NANDN U9218 ( .A(n8953), .B(n8952), .Z(n8957) );
  NAND U9219 ( .A(n8955), .B(n8954), .Z(n8956) );
  NAND U9220 ( .A(n8957), .B(n8956), .Z(n8996) );
  NAND U9221 ( .A(b[0]), .B(a[217]), .Z(n8958) );
  XNOR U9222 ( .A(b[1]), .B(n8958), .Z(n8960) );
  NAND U9223 ( .A(n46), .B(a[216]), .Z(n8959) );
  AND U9224 ( .A(n8960), .B(n8959), .Z(n9013) );
  XOR U9225 ( .A(a[213]), .B(n42197), .Z(n9002) );
  NANDN U9226 ( .A(n9002), .B(n42173), .Z(n8963) );
  NANDN U9227 ( .A(n8961), .B(n42172), .Z(n8962) );
  NAND U9228 ( .A(n8963), .B(n8962), .Z(n9011) );
  NAND U9229 ( .A(b[7]), .B(a[209]), .Z(n9012) );
  XNOR U9230 ( .A(n9011), .B(n9012), .Z(n9014) );
  XOR U9231 ( .A(n9013), .B(n9014), .Z(n9020) );
  NANDN U9232 ( .A(n8964), .B(n42093), .Z(n8966) );
  XOR U9233 ( .A(n42134), .B(a[215]), .Z(n9005) );
  NANDN U9234 ( .A(n9005), .B(n42095), .Z(n8965) );
  NAND U9235 ( .A(n8966), .B(n8965), .Z(n9018) );
  NANDN U9236 ( .A(n8967), .B(n42231), .Z(n8969) );
  XOR U9237 ( .A(n179), .B(a[211]), .Z(n9008) );
  NANDN U9238 ( .A(n9008), .B(n42234), .Z(n8968) );
  AND U9239 ( .A(n8969), .B(n8968), .Z(n9017) );
  XNOR U9240 ( .A(n9018), .B(n9017), .Z(n9019) );
  XNOR U9241 ( .A(n9020), .B(n9019), .Z(n9024) );
  NANDN U9242 ( .A(n8971), .B(n8970), .Z(n8975) );
  NAND U9243 ( .A(n8973), .B(n8972), .Z(n8974) );
  AND U9244 ( .A(n8975), .B(n8974), .Z(n9023) );
  XOR U9245 ( .A(n9024), .B(n9023), .Z(n9025) );
  NANDN U9246 ( .A(n8977), .B(n8976), .Z(n8981) );
  NANDN U9247 ( .A(n8979), .B(n8978), .Z(n8980) );
  NAND U9248 ( .A(n8981), .B(n8980), .Z(n9026) );
  XOR U9249 ( .A(n9025), .B(n9026), .Z(n8993) );
  OR U9250 ( .A(n8983), .B(n8982), .Z(n8987) );
  NANDN U9251 ( .A(n8985), .B(n8984), .Z(n8986) );
  NAND U9252 ( .A(n8987), .B(n8986), .Z(n8994) );
  XNOR U9253 ( .A(n8993), .B(n8994), .Z(n8995) );
  XNOR U9254 ( .A(n8996), .B(n8995), .Z(n9029) );
  XNOR U9255 ( .A(n9029), .B(sreg[1233]), .Z(n9031) );
  NAND U9256 ( .A(n8988), .B(sreg[1232]), .Z(n8992) );
  OR U9257 ( .A(n8990), .B(n8989), .Z(n8991) );
  AND U9258 ( .A(n8992), .B(n8991), .Z(n9030) );
  XOR U9259 ( .A(n9031), .B(n9030), .Z(c[1233]) );
  NANDN U9260 ( .A(n8994), .B(n8993), .Z(n8998) );
  NAND U9261 ( .A(n8996), .B(n8995), .Z(n8997) );
  NAND U9262 ( .A(n8998), .B(n8997), .Z(n9037) );
  NAND U9263 ( .A(b[0]), .B(a[218]), .Z(n8999) );
  XNOR U9264 ( .A(b[1]), .B(n8999), .Z(n9001) );
  NAND U9265 ( .A(n46), .B(a[217]), .Z(n9000) );
  AND U9266 ( .A(n9001), .B(n9000), .Z(n9054) );
  XOR U9267 ( .A(a[214]), .B(n42197), .Z(n9043) );
  NANDN U9268 ( .A(n9043), .B(n42173), .Z(n9004) );
  NANDN U9269 ( .A(n9002), .B(n42172), .Z(n9003) );
  NAND U9270 ( .A(n9004), .B(n9003), .Z(n9052) );
  NAND U9271 ( .A(b[7]), .B(a[210]), .Z(n9053) );
  XNOR U9272 ( .A(n9052), .B(n9053), .Z(n9055) );
  XOR U9273 ( .A(n9054), .B(n9055), .Z(n9061) );
  NANDN U9274 ( .A(n9005), .B(n42093), .Z(n9007) );
  XOR U9275 ( .A(n42134), .B(a[216]), .Z(n9046) );
  NANDN U9276 ( .A(n9046), .B(n42095), .Z(n9006) );
  NAND U9277 ( .A(n9007), .B(n9006), .Z(n9059) );
  NANDN U9278 ( .A(n9008), .B(n42231), .Z(n9010) );
  XOR U9279 ( .A(n179), .B(a[212]), .Z(n9049) );
  NANDN U9280 ( .A(n9049), .B(n42234), .Z(n9009) );
  AND U9281 ( .A(n9010), .B(n9009), .Z(n9058) );
  XNOR U9282 ( .A(n9059), .B(n9058), .Z(n9060) );
  XNOR U9283 ( .A(n9061), .B(n9060), .Z(n9065) );
  NANDN U9284 ( .A(n9012), .B(n9011), .Z(n9016) );
  NAND U9285 ( .A(n9014), .B(n9013), .Z(n9015) );
  AND U9286 ( .A(n9016), .B(n9015), .Z(n9064) );
  XOR U9287 ( .A(n9065), .B(n9064), .Z(n9066) );
  NANDN U9288 ( .A(n9018), .B(n9017), .Z(n9022) );
  NANDN U9289 ( .A(n9020), .B(n9019), .Z(n9021) );
  NAND U9290 ( .A(n9022), .B(n9021), .Z(n9067) );
  XOR U9291 ( .A(n9066), .B(n9067), .Z(n9034) );
  OR U9292 ( .A(n9024), .B(n9023), .Z(n9028) );
  NANDN U9293 ( .A(n9026), .B(n9025), .Z(n9027) );
  NAND U9294 ( .A(n9028), .B(n9027), .Z(n9035) );
  XNOR U9295 ( .A(n9034), .B(n9035), .Z(n9036) );
  XNOR U9296 ( .A(n9037), .B(n9036), .Z(n9070) );
  XNOR U9297 ( .A(n9070), .B(sreg[1234]), .Z(n9072) );
  NAND U9298 ( .A(n9029), .B(sreg[1233]), .Z(n9033) );
  OR U9299 ( .A(n9031), .B(n9030), .Z(n9032) );
  AND U9300 ( .A(n9033), .B(n9032), .Z(n9071) );
  XOR U9301 ( .A(n9072), .B(n9071), .Z(c[1234]) );
  NANDN U9302 ( .A(n9035), .B(n9034), .Z(n9039) );
  NAND U9303 ( .A(n9037), .B(n9036), .Z(n9038) );
  NAND U9304 ( .A(n9039), .B(n9038), .Z(n9078) );
  NAND U9305 ( .A(b[0]), .B(a[219]), .Z(n9040) );
  XNOR U9306 ( .A(b[1]), .B(n9040), .Z(n9042) );
  NAND U9307 ( .A(n46), .B(a[218]), .Z(n9041) );
  AND U9308 ( .A(n9042), .B(n9041), .Z(n9095) );
  XOR U9309 ( .A(a[215]), .B(n42197), .Z(n9084) );
  NANDN U9310 ( .A(n9084), .B(n42173), .Z(n9045) );
  NANDN U9311 ( .A(n9043), .B(n42172), .Z(n9044) );
  NAND U9312 ( .A(n9045), .B(n9044), .Z(n9093) );
  NAND U9313 ( .A(b[7]), .B(a[211]), .Z(n9094) );
  XNOR U9314 ( .A(n9093), .B(n9094), .Z(n9096) );
  XOR U9315 ( .A(n9095), .B(n9096), .Z(n9102) );
  NANDN U9316 ( .A(n9046), .B(n42093), .Z(n9048) );
  XOR U9317 ( .A(n42134), .B(a[217]), .Z(n9087) );
  NANDN U9318 ( .A(n9087), .B(n42095), .Z(n9047) );
  NAND U9319 ( .A(n9048), .B(n9047), .Z(n9100) );
  NANDN U9320 ( .A(n9049), .B(n42231), .Z(n9051) );
  XOR U9321 ( .A(n179), .B(a[213]), .Z(n9090) );
  NANDN U9322 ( .A(n9090), .B(n42234), .Z(n9050) );
  AND U9323 ( .A(n9051), .B(n9050), .Z(n9099) );
  XNOR U9324 ( .A(n9100), .B(n9099), .Z(n9101) );
  XNOR U9325 ( .A(n9102), .B(n9101), .Z(n9106) );
  NANDN U9326 ( .A(n9053), .B(n9052), .Z(n9057) );
  NAND U9327 ( .A(n9055), .B(n9054), .Z(n9056) );
  AND U9328 ( .A(n9057), .B(n9056), .Z(n9105) );
  XOR U9329 ( .A(n9106), .B(n9105), .Z(n9107) );
  NANDN U9330 ( .A(n9059), .B(n9058), .Z(n9063) );
  NANDN U9331 ( .A(n9061), .B(n9060), .Z(n9062) );
  NAND U9332 ( .A(n9063), .B(n9062), .Z(n9108) );
  XOR U9333 ( .A(n9107), .B(n9108), .Z(n9075) );
  OR U9334 ( .A(n9065), .B(n9064), .Z(n9069) );
  NANDN U9335 ( .A(n9067), .B(n9066), .Z(n9068) );
  NAND U9336 ( .A(n9069), .B(n9068), .Z(n9076) );
  XNOR U9337 ( .A(n9075), .B(n9076), .Z(n9077) );
  XNOR U9338 ( .A(n9078), .B(n9077), .Z(n9111) );
  XNOR U9339 ( .A(n9111), .B(sreg[1235]), .Z(n9113) );
  NAND U9340 ( .A(n9070), .B(sreg[1234]), .Z(n9074) );
  OR U9341 ( .A(n9072), .B(n9071), .Z(n9073) );
  AND U9342 ( .A(n9074), .B(n9073), .Z(n9112) );
  XOR U9343 ( .A(n9113), .B(n9112), .Z(c[1235]) );
  NANDN U9344 ( .A(n9076), .B(n9075), .Z(n9080) );
  NAND U9345 ( .A(n9078), .B(n9077), .Z(n9079) );
  NAND U9346 ( .A(n9080), .B(n9079), .Z(n9119) );
  NAND U9347 ( .A(b[0]), .B(a[220]), .Z(n9081) );
  XNOR U9348 ( .A(b[1]), .B(n9081), .Z(n9083) );
  NAND U9349 ( .A(n46), .B(a[219]), .Z(n9082) );
  AND U9350 ( .A(n9083), .B(n9082), .Z(n9136) );
  XOR U9351 ( .A(a[216]), .B(n42197), .Z(n9125) );
  NANDN U9352 ( .A(n9125), .B(n42173), .Z(n9086) );
  NANDN U9353 ( .A(n9084), .B(n42172), .Z(n9085) );
  NAND U9354 ( .A(n9086), .B(n9085), .Z(n9134) );
  NAND U9355 ( .A(b[7]), .B(a[212]), .Z(n9135) );
  XNOR U9356 ( .A(n9134), .B(n9135), .Z(n9137) );
  XOR U9357 ( .A(n9136), .B(n9137), .Z(n9143) );
  NANDN U9358 ( .A(n9087), .B(n42093), .Z(n9089) );
  XOR U9359 ( .A(n42134), .B(a[218]), .Z(n9128) );
  NANDN U9360 ( .A(n9128), .B(n42095), .Z(n9088) );
  NAND U9361 ( .A(n9089), .B(n9088), .Z(n9141) );
  NANDN U9362 ( .A(n9090), .B(n42231), .Z(n9092) );
  XOR U9363 ( .A(n179), .B(a[214]), .Z(n9131) );
  NANDN U9364 ( .A(n9131), .B(n42234), .Z(n9091) );
  AND U9365 ( .A(n9092), .B(n9091), .Z(n9140) );
  XNOR U9366 ( .A(n9141), .B(n9140), .Z(n9142) );
  XNOR U9367 ( .A(n9143), .B(n9142), .Z(n9147) );
  NANDN U9368 ( .A(n9094), .B(n9093), .Z(n9098) );
  NAND U9369 ( .A(n9096), .B(n9095), .Z(n9097) );
  AND U9370 ( .A(n9098), .B(n9097), .Z(n9146) );
  XOR U9371 ( .A(n9147), .B(n9146), .Z(n9148) );
  NANDN U9372 ( .A(n9100), .B(n9099), .Z(n9104) );
  NANDN U9373 ( .A(n9102), .B(n9101), .Z(n9103) );
  NAND U9374 ( .A(n9104), .B(n9103), .Z(n9149) );
  XOR U9375 ( .A(n9148), .B(n9149), .Z(n9116) );
  OR U9376 ( .A(n9106), .B(n9105), .Z(n9110) );
  NANDN U9377 ( .A(n9108), .B(n9107), .Z(n9109) );
  NAND U9378 ( .A(n9110), .B(n9109), .Z(n9117) );
  XNOR U9379 ( .A(n9116), .B(n9117), .Z(n9118) );
  XNOR U9380 ( .A(n9119), .B(n9118), .Z(n9152) );
  XNOR U9381 ( .A(n9152), .B(sreg[1236]), .Z(n9154) );
  NAND U9382 ( .A(n9111), .B(sreg[1235]), .Z(n9115) );
  OR U9383 ( .A(n9113), .B(n9112), .Z(n9114) );
  AND U9384 ( .A(n9115), .B(n9114), .Z(n9153) );
  XOR U9385 ( .A(n9154), .B(n9153), .Z(c[1236]) );
  NANDN U9386 ( .A(n9117), .B(n9116), .Z(n9121) );
  NAND U9387 ( .A(n9119), .B(n9118), .Z(n9120) );
  NAND U9388 ( .A(n9121), .B(n9120), .Z(n9160) );
  NAND U9389 ( .A(b[0]), .B(a[221]), .Z(n9122) );
  XNOR U9390 ( .A(b[1]), .B(n9122), .Z(n9124) );
  NAND U9391 ( .A(n46), .B(a[220]), .Z(n9123) );
  AND U9392 ( .A(n9124), .B(n9123), .Z(n9177) );
  XOR U9393 ( .A(a[217]), .B(n42197), .Z(n9166) );
  NANDN U9394 ( .A(n9166), .B(n42173), .Z(n9127) );
  NANDN U9395 ( .A(n9125), .B(n42172), .Z(n9126) );
  NAND U9396 ( .A(n9127), .B(n9126), .Z(n9175) );
  NAND U9397 ( .A(b[7]), .B(a[213]), .Z(n9176) );
  XNOR U9398 ( .A(n9175), .B(n9176), .Z(n9178) );
  XOR U9399 ( .A(n9177), .B(n9178), .Z(n9184) );
  NANDN U9400 ( .A(n9128), .B(n42093), .Z(n9130) );
  XOR U9401 ( .A(n42134), .B(a[219]), .Z(n9169) );
  NANDN U9402 ( .A(n9169), .B(n42095), .Z(n9129) );
  NAND U9403 ( .A(n9130), .B(n9129), .Z(n9182) );
  NANDN U9404 ( .A(n9131), .B(n42231), .Z(n9133) );
  XOR U9405 ( .A(n180), .B(a[215]), .Z(n9172) );
  NANDN U9406 ( .A(n9172), .B(n42234), .Z(n9132) );
  AND U9407 ( .A(n9133), .B(n9132), .Z(n9181) );
  XNOR U9408 ( .A(n9182), .B(n9181), .Z(n9183) );
  XNOR U9409 ( .A(n9184), .B(n9183), .Z(n9188) );
  NANDN U9410 ( .A(n9135), .B(n9134), .Z(n9139) );
  NAND U9411 ( .A(n9137), .B(n9136), .Z(n9138) );
  AND U9412 ( .A(n9139), .B(n9138), .Z(n9187) );
  XOR U9413 ( .A(n9188), .B(n9187), .Z(n9189) );
  NANDN U9414 ( .A(n9141), .B(n9140), .Z(n9145) );
  NANDN U9415 ( .A(n9143), .B(n9142), .Z(n9144) );
  NAND U9416 ( .A(n9145), .B(n9144), .Z(n9190) );
  XOR U9417 ( .A(n9189), .B(n9190), .Z(n9157) );
  OR U9418 ( .A(n9147), .B(n9146), .Z(n9151) );
  NANDN U9419 ( .A(n9149), .B(n9148), .Z(n9150) );
  NAND U9420 ( .A(n9151), .B(n9150), .Z(n9158) );
  XNOR U9421 ( .A(n9157), .B(n9158), .Z(n9159) );
  XNOR U9422 ( .A(n9160), .B(n9159), .Z(n9193) );
  XNOR U9423 ( .A(n9193), .B(sreg[1237]), .Z(n9195) );
  NAND U9424 ( .A(n9152), .B(sreg[1236]), .Z(n9156) );
  OR U9425 ( .A(n9154), .B(n9153), .Z(n9155) );
  AND U9426 ( .A(n9156), .B(n9155), .Z(n9194) );
  XOR U9427 ( .A(n9195), .B(n9194), .Z(c[1237]) );
  NANDN U9428 ( .A(n9158), .B(n9157), .Z(n9162) );
  NAND U9429 ( .A(n9160), .B(n9159), .Z(n9161) );
  NAND U9430 ( .A(n9162), .B(n9161), .Z(n9201) );
  NAND U9431 ( .A(b[0]), .B(a[222]), .Z(n9163) );
  XNOR U9432 ( .A(b[1]), .B(n9163), .Z(n9165) );
  NAND U9433 ( .A(n46), .B(a[221]), .Z(n9164) );
  AND U9434 ( .A(n9165), .B(n9164), .Z(n9218) );
  XOR U9435 ( .A(a[218]), .B(n42197), .Z(n9207) );
  NANDN U9436 ( .A(n9207), .B(n42173), .Z(n9168) );
  NANDN U9437 ( .A(n9166), .B(n42172), .Z(n9167) );
  NAND U9438 ( .A(n9168), .B(n9167), .Z(n9216) );
  NAND U9439 ( .A(b[7]), .B(a[214]), .Z(n9217) );
  XNOR U9440 ( .A(n9216), .B(n9217), .Z(n9219) );
  XOR U9441 ( .A(n9218), .B(n9219), .Z(n9225) );
  NANDN U9442 ( .A(n9169), .B(n42093), .Z(n9171) );
  XOR U9443 ( .A(n42134), .B(a[220]), .Z(n9210) );
  NANDN U9444 ( .A(n9210), .B(n42095), .Z(n9170) );
  NAND U9445 ( .A(n9171), .B(n9170), .Z(n9223) );
  NANDN U9446 ( .A(n9172), .B(n42231), .Z(n9174) );
  XOR U9447 ( .A(n180), .B(a[216]), .Z(n9213) );
  NANDN U9448 ( .A(n9213), .B(n42234), .Z(n9173) );
  AND U9449 ( .A(n9174), .B(n9173), .Z(n9222) );
  XNOR U9450 ( .A(n9223), .B(n9222), .Z(n9224) );
  XNOR U9451 ( .A(n9225), .B(n9224), .Z(n9229) );
  NANDN U9452 ( .A(n9176), .B(n9175), .Z(n9180) );
  NAND U9453 ( .A(n9178), .B(n9177), .Z(n9179) );
  AND U9454 ( .A(n9180), .B(n9179), .Z(n9228) );
  XOR U9455 ( .A(n9229), .B(n9228), .Z(n9230) );
  NANDN U9456 ( .A(n9182), .B(n9181), .Z(n9186) );
  NANDN U9457 ( .A(n9184), .B(n9183), .Z(n9185) );
  NAND U9458 ( .A(n9186), .B(n9185), .Z(n9231) );
  XOR U9459 ( .A(n9230), .B(n9231), .Z(n9198) );
  OR U9460 ( .A(n9188), .B(n9187), .Z(n9192) );
  NANDN U9461 ( .A(n9190), .B(n9189), .Z(n9191) );
  NAND U9462 ( .A(n9192), .B(n9191), .Z(n9199) );
  XNOR U9463 ( .A(n9198), .B(n9199), .Z(n9200) );
  XNOR U9464 ( .A(n9201), .B(n9200), .Z(n9234) );
  XNOR U9465 ( .A(n9234), .B(sreg[1238]), .Z(n9236) );
  NAND U9466 ( .A(n9193), .B(sreg[1237]), .Z(n9197) );
  OR U9467 ( .A(n9195), .B(n9194), .Z(n9196) );
  AND U9468 ( .A(n9197), .B(n9196), .Z(n9235) );
  XOR U9469 ( .A(n9236), .B(n9235), .Z(c[1238]) );
  NANDN U9470 ( .A(n9199), .B(n9198), .Z(n9203) );
  NAND U9471 ( .A(n9201), .B(n9200), .Z(n9202) );
  NAND U9472 ( .A(n9203), .B(n9202), .Z(n9242) );
  NAND U9473 ( .A(b[0]), .B(a[223]), .Z(n9204) );
  XNOR U9474 ( .A(b[1]), .B(n9204), .Z(n9206) );
  NAND U9475 ( .A(n46), .B(a[222]), .Z(n9205) );
  AND U9476 ( .A(n9206), .B(n9205), .Z(n9259) );
  XOR U9477 ( .A(a[219]), .B(n42197), .Z(n9248) );
  NANDN U9478 ( .A(n9248), .B(n42173), .Z(n9209) );
  NANDN U9479 ( .A(n9207), .B(n42172), .Z(n9208) );
  NAND U9480 ( .A(n9209), .B(n9208), .Z(n9257) );
  NAND U9481 ( .A(b[7]), .B(a[215]), .Z(n9258) );
  XNOR U9482 ( .A(n9257), .B(n9258), .Z(n9260) );
  XOR U9483 ( .A(n9259), .B(n9260), .Z(n9266) );
  NANDN U9484 ( .A(n9210), .B(n42093), .Z(n9212) );
  XOR U9485 ( .A(n42134), .B(a[221]), .Z(n9251) );
  NANDN U9486 ( .A(n9251), .B(n42095), .Z(n9211) );
  NAND U9487 ( .A(n9212), .B(n9211), .Z(n9264) );
  NANDN U9488 ( .A(n9213), .B(n42231), .Z(n9215) );
  XOR U9489 ( .A(n180), .B(a[217]), .Z(n9254) );
  NANDN U9490 ( .A(n9254), .B(n42234), .Z(n9214) );
  AND U9491 ( .A(n9215), .B(n9214), .Z(n9263) );
  XNOR U9492 ( .A(n9264), .B(n9263), .Z(n9265) );
  XNOR U9493 ( .A(n9266), .B(n9265), .Z(n9270) );
  NANDN U9494 ( .A(n9217), .B(n9216), .Z(n9221) );
  NAND U9495 ( .A(n9219), .B(n9218), .Z(n9220) );
  AND U9496 ( .A(n9221), .B(n9220), .Z(n9269) );
  XOR U9497 ( .A(n9270), .B(n9269), .Z(n9271) );
  NANDN U9498 ( .A(n9223), .B(n9222), .Z(n9227) );
  NANDN U9499 ( .A(n9225), .B(n9224), .Z(n9226) );
  NAND U9500 ( .A(n9227), .B(n9226), .Z(n9272) );
  XOR U9501 ( .A(n9271), .B(n9272), .Z(n9239) );
  OR U9502 ( .A(n9229), .B(n9228), .Z(n9233) );
  NANDN U9503 ( .A(n9231), .B(n9230), .Z(n9232) );
  NAND U9504 ( .A(n9233), .B(n9232), .Z(n9240) );
  XNOR U9505 ( .A(n9239), .B(n9240), .Z(n9241) );
  XNOR U9506 ( .A(n9242), .B(n9241), .Z(n9275) );
  XNOR U9507 ( .A(n9275), .B(sreg[1239]), .Z(n9277) );
  NAND U9508 ( .A(n9234), .B(sreg[1238]), .Z(n9238) );
  OR U9509 ( .A(n9236), .B(n9235), .Z(n9237) );
  AND U9510 ( .A(n9238), .B(n9237), .Z(n9276) );
  XOR U9511 ( .A(n9277), .B(n9276), .Z(c[1239]) );
  NANDN U9512 ( .A(n9240), .B(n9239), .Z(n9244) );
  NAND U9513 ( .A(n9242), .B(n9241), .Z(n9243) );
  NAND U9514 ( .A(n9244), .B(n9243), .Z(n9283) );
  NAND U9515 ( .A(b[0]), .B(a[224]), .Z(n9245) );
  XNOR U9516 ( .A(b[1]), .B(n9245), .Z(n9247) );
  NAND U9517 ( .A(n47), .B(a[223]), .Z(n9246) );
  AND U9518 ( .A(n9247), .B(n9246), .Z(n9300) );
  XOR U9519 ( .A(a[220]), .B(n42197), .Z(n9289) );
  NANDN U9520 ( .A(n9289), .B(n42173), .Z(n9250) );
  NANDN U9521 ( .A(n9248), .B(n42172), .Z(n9249) );
  NAND U9522 ( .A(n9250), .B(n9249), .Z(n9298) );
  NAND U9523 ( .A(b[7]), .B(a[216]), .Z(n9299) );
  XNOR U9524 ( .A(n9298), .B(n9299), .Z(n9301) );
  XOR U9525 ( .A(n9300), .B(n9301), .Z(n9307) );
  NANDN U9526 ( .A(n9251), .B(n42093), .Z(n9253) );
  XOR U9527 ( .A(n42134), .B(a[222]), .Z(n9292) );
  NANDN U9528 ( .A(n9292), .B(n42095), .Z(n9252) );
  NAND U9529 ( .A(n9253), .B(n9252), .Z(n9305) );
  NANDN U9530 ( .A(n9254), .B(n42231), .Z(n9256) );
  XOR U9531 ( .A(n180), .B(a[218]), .Z(n9295) );
  NANDN U9532 ( .A(n9295), .B(n42234), .Z(n9255) );
  AND U9533 ( .A(n9256), .B(n9255), .Z(n9304) );
  XNOR U9534 ( .A(n9305), .B(n9304), .Z(n9306) );
  XNOR U9535 ( .A(n9307), .B(n9306), .Z(n9311) );
  NANDN U9536 ( .A(n9258), .B(n9257), .Z(n9262) );
  NAND U9537 ( .A(n9260), .B(n9259), .Z(n9261) );
  AND U9538 ( .A(n9262), .B(n9261), .Z(n9310) );
  XOR U9539 ( .A(n9311), .B(n9310), .Z(n9312) );
  NANDN U9540 ( .A(n9264), .B(n9263), .Z(n9268) );
  NANDN U9541 ( .A(n9266), .B(n9265), .Z(n9267) );
  NAND U9542 ( .A(n9268), .B(n9267), .Z(n9313) );
  XOR U9543 ( .A(n9312), .B(n9313), .Z(n9280) );
  OR U9544 ( .A(n9270), .B(n9269), .Z(n9274) );
  NANDN U9545 ( .A(n9272), .B(n9271), .Z(n9273) );
  NAND U9546 ( .A(n9274), .B(n9273), .Z(n9281) );
  XNOR U9547 ( .A(n9280), .B(n9281), .Z(n9282) );
  XNOR U9548 ( .A(n9283), .B(n9282), .Z(n9316) );
  XNOR U9549 ( .A(n9316), .B(sreg[1240]), .Z(n9318) );
  NAND U9550 ( .A(n9275), .B(sreg[1239]), .Z(n9279) );
  OR U9551 ( .A(n9277), .B(n9276), .Z(n9278) );
  AND U9552 ( .A(n9279), .B(n9278), .Z(n9317) );
  XOR U9553 ( .A(n9318), .B(n9317), .Z(c[1240]) );
  NANDN U9554 ( .A(n9281), .B(n9280), .Z(n9285) );
  NAND U9555 ( .A(n9283), .B(n9282), .Z(n9284) );
  NAND U9556 ( .A(n9285), .B(n9284), .Z(n9324) );
  NAND U9557 ( .A(b[0]), .B(a[225]), .Z(n9286) );
  XNOR U9558 ( .A(b[1]), .B(n9286), .Z(n9288) );
  NAND U9559 ( .A(n47), .B(a[224]), .Z(n9287) );
  AND U9560 ( .A(n9288), .B(n9287), .Z(n9341) );
  XOR U9561 ( .A(a[221]), .B(n42197), .Z(n9330) );
  NANDN U9562 ( .A(n9330), .B(n42173), .Z(n9291) );
  NANDN U9563 ( .A(n9289), .B(n42172), .Z(n9290) );
  NAND U9564 ( .A(n9291), .B(n9290), .Z(n9339) );
  NAND U9565 ( .A(b[7]), .B(a[217]), .Z(n9340) );
  XNOR U9566 ( .A(n9339), .B(n9340), .Z(n9342) );
  XOR U9567 ( .A(n9341), .B(n9342), .Z(n9348) );
  NANDN U9568 ( .A(n9292), .B(n42093), .Z(n9294) );
  XOR U9569 ( .A(n42134), .B(a[223]), .Z(n9333) );
  NANDN U9570 ( .A(n9333), .B(n42095), .Z(n9293) );
  NAND U9571 ( .A(n9294), .B(n9293), .Z(n9346) );
  NANDN U9572 ( .A(n9295), .B(n42231), .Z(n9297) );
  XOR U9573 ( .A(n180), .B(a[219]), .Z(n9336) );
  NANDN U9574 ( .A(n9336), .B(n42234), .Z(n9296) );
  AND U9575 ( .A(n9297), .B(n9296), .Z(n9345) );
  XNOR U9576 ( .A(n9346), .B(n9345), .Z(n9347) );
  XNOR U9577 ( .A(n9348), .B(n9347), .Z(n9352) );
  NANDN U9578 ( .A(n9299), .B(n9298), .Z(n9303) );
  NAND U9579 ( .A(n9301), .B(n9300), .Z(n9302) );
  AND U9580 ( .A(n9303), .B(n9302), .Z(n9351) );
  XOR U9581 ( .A(n9352), .B(n9351), .Z(n9353) );
  NANDN U9582 ( .A(n9305), .B(n9304), .Z(n9309) );
  NANDN U9583 ( .A(n9307), .B(n9306), .Z(n9308) );
  NAND U9584 ( .A(n9309), .B(n9308), .Z(n9354) );
  XOR U9585 ( .A(n9353), .B(n9354), .Z(n9321) );
  OR U9586 ( .A(n9311), .B(n9310), .Z(n9315) );
  NANDN U9587 ( .A(n9313), .B(n9312), .Z(n9314) );
  NAND U9588 ( .A(n9315), .B(n9314), .Z(n9322) );
  XNOR U9589 ( .A(n9321), .B(n9322), .Z(n9323) );
  XNOR U9590 ( .A(n9324), .B(n9323), .Z(n9357) );
  XNOR U9591 ( .A(n9357), .B(sreg[1241]), .Z(n9359) );
  NAND U9592 ( .A(n9316), .B(sreg[1240]), .Z(n9320) );
  OR U9593 ( .A(n9318), .B(n9317), .Z(n9319) );
  AND U9594 ( .A(n9320), .B(n9319), .Z(n9358) );
  XOR U9595 ( .A(n9359), .B(n9358), .Z(c[1241]) );
  NANDN U9596 ( .A(n9322), .B(n9321), .Z(n9326) );
  NAND U9597 ( .A(n9324), .B(n9323), .Z(n9325) );
  NAND U9598 ( .A(n9326), .B(n9325), .Z(n9365) );
  NAND U9599 ( .A(b[0]), .B(a[226]), .Z(n9327) );
  XNOR U9600 ( .A(b[1]), .B(n9327), .Z(n9329) );
  NAND U9601 ( .A(n47), .B(a[225]), .Z(n9328) );
  AND U9602 ( .A(n9329), .B(n9328), .Z(n9382) );
  XOR U9603 ( .A(a[222]), .B(n42197), .Z(n9371) );
  NANDN U9604 ( .A(n9371), .B(n42173), .Z(n9332) );
  NANDN U9605 ( .A(n9330), .B(n42172), .Z(n9331) );
  NAND U9606 ( .A(n9332), .B(n9331), .Z(n9380) );
  NAND U9607 ( .A(b[7]), .B(a[218]), .Z(n9381) );
  XNOR U9608 ( .A(n9380), .B(n9381), .Z(n9383) );
  XOR U9609 ( .A(n9382), .B(n9383), .Z(n9389) );
  NANDN U9610 ( .A(n9333), .B(n42093), .Z(n9335) );
  XOR U9611 ( .A(n42134), .B(a[224]), .Z(n9374) );
  NANDN U9612 ( .A(n9374), .B(n42095), .Z(n9334) );
  NAND U9613 ( .A(n9335), .B(n9334), .Z(n9387) );
  NANDN U9614 ( .A(n9336), .B(n42231), .Z(n9338) );
  XOR U9615 ( .A(n180), .B(a[220]), .Z(n9377) );
  NANDN U9616 ( .A(n9377), .B(n42234), .Z(n9337) );
  AND U9617 ( .A(n9338), .B(n9337), .Z(n9386) );
  XNOR U9618 ( .A(n9387), .B(n9386), .Z(n9388) );
  XNOR U9619 ( .A(n9389), .B(n9388), .Z(n9393) );
  NANDN U9620 ( .A(n9340), .B(n9339), .Z(n9344) );
  NAND U9621 ( .A(n9342), .B(n9341), .Z(n9343) );
  AND U9622 ( .A(n9344), .B(n9343), .Z(n9392) );
  XOR U9623 ( .A(n9393), .B(n9392), .Z(n9394) );
  NANDN U9624 ( .A(n9346), .B(n9345), .Z(n9350) );
  NANDN U9625 ( .A(n9348), .B(n9347), .Z(n9349) );
  NAND U9626 ( .A(n9350), .B(n9349), .Z(n9395) );
  XOR U9627 ( .A(n9394), .B(n9395), .Z(n9362) );
  OR U9628 ( .A(n9352), .B(n9351), .Z(n9356) );
  NANDN U9629 ( .A(n9354), .B(n9353), .Z(n9355) );
  NAND U9630 ( .A(n9356), .B(n9355), .Z(n9363) );
  XNOR U9631 ( .A(n9362), .B(n9363), .Z(n9364) );
  XNOR U9632 ( .A(n9365), .B(n9364), .Z(n9398) );
  XNOR U9633 ( .A(n9398), .B(sreg[1242]), .Z(n9400) );
  NAND U9634 ( .A(n9357), .B(sreg[1241]), .Z(n9361) );
  OR U9635 ( .A(n9359), .B(n9358), .Z(n9360) );
  AND U9636 ( .A(n9361), .B(n9360), .Z(n9399) );
  XOR U9637 ( .A(n9400), .B(n9399), .Z(c[1242]) );
  NANDN U9638 ( .A(n9363), .B(n9362), .Z(n9367) );
  NAND U9639 ( .A(n9365), .B(n9364), .Z(n9366) );
  NAND U9640 ( .A(n9367), .B(n9366), .Z(n9406) );
  NAND U9641 ( .A(b[0]), .B(a[227]), .Z(n9368) );
  XNOR U9642 ( .A(b[1]), .B(n9368), .Z(n9370) );
  NAND U9643 ( .A(n47), .B(a[226]), .Z(n9369) );
  AND U9644 ( .A(n9370), .B(n9369), .Z(n9423) );
  XOR U9645 ( .A(a[223]), .B(n42197), .Z(n9412) );
  NANDN U9646 ( .A(n9412), .B(n42173), .Z(n9373) );
  NANDN U9647 ( .A(n9371), .B(n42172), .Z(n9372) );
  NAND U9648 ( .A(n9373), .B(n9372), .Z(n9421) );
  NAND U9649 ( .A(b[7]), .B(a[219]), .Z(n9422) );
  XNOR U9650 ( .A(n9421), .B(n9422), .Z(n9424) );
  XOR U9651 ( .A(n9423), .B(n9424), .Z(n9430) );
  NANDN U9652 ( .A(n9374), .B(n42093), .Z(n9376) );
  XOR U9653 ( .A(n42134), .B(a[225]), .Z(n9415) );
  NANDN U9654 ( .A(n9415), .B(n42095), .Z(n9375) );
  NAND U9655 ( .A(n9376), .B(n9375), .Z(n9428) );
  NANDN U9656 ( .A(n9377), .B(n42231), .Z(n9379) );
  XOR U9657 ( .A(n180), .B(a[221]), .Z(n9418) );
  NANDN U9658 ( .A(n9418), .B(n42234), .Z(n9378) );
  AND U9659 ( .A(n9379), .B(n9378), .Z(n9427) );
  XNOR U9660 ( .A(n9428), .B(n9427), .Z(n9429) );
  XNOR U9661 ( .A(n9430), .B(n9429), .Z(n9434) );
  NANDN U9662 ( .A(n9381), .B(n9380), .Z(n9385) );
  NAND U9663 ( .A(n9383), .B(n9382), .Z(n9384) );
  AND U9664 ( .A(n9385), .B(n9384), .Z(n9433) );
  XOR U9665 ( .A(n9434), .B(n9433), .Z(n9435) );
  NANDN U9666 ( .A(n9387), .B(n9386), .Z(n9391) );
  NANDN U9667 ( .A(n9389), .B(n9388), .Z(n9390) );
  NAND U9668 ( .A(n9391), .B(n9390), .Z(n9436) );
  XOR U9669 ( .A(n9435), .B(n9436), .Z(n9403) );
  OR U9670 ( .A(n9393), .B(n9392), .Z(n9397) );
  NANDN U9671 ( .A(n9395), .B(n9394), .Z(n9396) );
  NAND U9672 ( .A(n9397), .B(n9396), .Z(n9404) );
  XNOR U9673 ( .A(n9403), .B(n9404), .Z(n9405) );
  XNOR U9674 ( .A(n9406), .B(n9405), .Z(n9439) );
  XNOR U9675 ( .A(n9439), .B(sreg[1243]), .Z(n9441) );
  NAND U9676 ( .A(n9398), .B(sreg[1242]), .Z(n9402) );
  OR U9677 ( .A(n9400), .B(n9399), .Z(n9401) );
  AND U9678 ( .A(n9402), .B(n9401), .Z(n9440) );
  XOR U9679 ( .A(n9441), .B(n9440), .Z(c[1243]) );
  NANDN U9680 ( .A(n9404), .B(n9403), .Z(n9408) );
  NAND U9681 ( .A(n9406), .B(n9405), .Z(n9407) );
  NAND U9682 ( .A(n9408), .B(n9407), .Z(n9447) );
  NAND U9683 ( .A(b[0]), .B(a[228]), .Z(n9409) );
  XNOR U9684 ( .A(b[1]), .B(n9409), .Z(n9411) );
  NAND U9685 ( .A(n47), .B(a[227]), .Z(n9410) );
  AND U9686 ( .A(n9411), .B(n9410), .Z(n9464) );
  XOR U9687 ( .A(a[224]), .B(n42197), .Z(n9453) );
  NANDN U9688 ( .A(n9453), .B(n42173), .Z(n9414) );
  NANDN U9689 ( .A(n9412), .B(n42172), .Z(n9413) );
  NAND U9690 ( .A(n9414), .B(n9413), .Z(n9462) );
  NAND U9691 ( .A(b[7]), .B(a[220]), .Z(n9463) );
  XNOR U9692 ( .A(n9462), .B(n9463), .Z(n9465) );
  XOR U9693 ( .A(n9464), .B(n9465), .Z(n9471) );
  NANDN U9694 ( .A(n9415), .B(n42093), .Z(n9417) );
  XOR U9695 ( .A(n42134), .B(a[226]), .Z(n9456) );
  NANDN U9696 ( .A(n9456), .B(n42095), .Z(n9416) );
  NAND U9697 ( .A(n9417), .B(n9416), .Z(n9469) );
  NANDN U9698 ( .A(n9418), .B(n42231), .Z(n9420) );
  XOR U9699 ( .A(n180), .B(a[222]), .Z(n9459) );
  NANDN U9700 ( .A(n9459), .B(n42234), .Z(n9419) );
  AND U9701 ( .A(n9420), .B(n9419), .Z(n9468) );
  XNOR U9702 ( .A(n9469), .B(n9468), .Z(n9470) );
  XNOR U9703 ( .A(n9471), .B(n9470), .Z(n9475) );
  NANDN U9704 ( .A(n9422), .B(n9421), .Z(n9426) );
  NAND U9705 ( .A(n9424), .B(n9423), .Z(n9425) );
  AND U9706 ( .A(n9426), .B(n9425), .Z(n9474) );
  XOR U9707 ( .A(n9475), .B(n9474), .Z(n9476) );
  NANDN U9708 ( .A(n9428), .B(n9427), .Z(n9432) );
  NANDN U9709 ( .A(n9430), .B(n9429), .Z(n9431) );
  NAND U9710 ( .A(n9432), .B(n9431), .Z(n9477) );
  XOR U9711 ( .A(n9476), .B(n9477), .Z(n9444) );
  OR U9712 ( .A(n9434), .B(n9433), .Z(n9438) );
  NANDN U9713 ( .A(n9436), .B(n9435), .Z(n9437) );
  NAND U9714 ( .A(n9438), .B(n9437), .Z(n9445) );
  XNOR U9715 ( .A(n9444), .B(n9445), .Z(n9446) );
  XNOR U9716 ( .A(n9447), .B(n9446), .Z(n9480) );
  XNOR U9717 ( .A(n9480), .B(sreg[1244]), .Z(n9482) );
  NAND U9718 ( .A(n9439), .B(sreg[1243]), .Z(n9443) );
  OR U9719 ( .A(n9441), .B(n9440), .Z(n9442) );
  AND U9720 ( .A(n9443), .B(n9442), .Z(n9481) );
  XOR U9721 ( .A(n9482), .B(n9481), .Z(c[1244]) );
  NANDN U9722 ( .A(n9445), .B(n9444), .Z(n9449) );
  NAND U9723 ( .A(n9447), .B(n9446), .Z(n9448) );
  NAND U9724 ( .A(n9449), .B(n9448), .Z(n9488) );
  NAND U9725 ( .A(b[0]), .B(a[229]), .Z(n9450) );
  XNOR U9726 ( .A(b[1]), .B(n9450), .Z(n9452) );
  NAND U9727 ( .A(n47), .B(a[228]), .Z(n9451) );
  AND U9728 ( .A(n9452), .B(n9451), .Z(n9505) );
  XOR U9729 ( .A(a[225]), .B(n42197), .Z(n9494) );
  NANDN U9730 ( .A(n9494), .B(n42173), .Z(n9455) );
  NANDN U9731 ( .A(n9453), .B(n42172), .Z(n9454) );
  NAND U9732 ( .A(n9455), .B(n9454), .Z(n9503) );
  NAND U9733 ( .A(b[7]), .B(a[221]), .Z(n9504) );
  XNOR U9734 ( .A(n9503), .B(n9504), .Z(n9506) );
  XOR U9735 ( .A(n9505), .B(n9506), .Z(n9512) );
  NANDN U9736 ( .A(n9456), .B(n42093), .Z(n9458) );
  XOR U9737 ( .A(n42134), .B(a[227]), .Z(n9497) );
  NANDN U9738 ( .A(n9497), .B(n42095), .Z(n9457) );
  NAND U9739 ( .A(n9458), .B(n9457), .Z(n9510) );
  NANDN U9740 ( .A(n9459), .B(n42231), .Z(n9461) );
  XOR U9741 ( .A(n180), .B(a[223]), .Z(n9500) );
  NANDN U9742 ( .A(n9500), .B(n42234), .Z(n9460) );
  AND U9743 ( .A(n9461), .B(n9460), .Z(n9509) );
  XNOR U9744 ( .A(n9510), .B(n9509), .Z(n9511) );
  XNOR U9745 ( .A(n9512), .B(n9511), .Z(n9516) );
  NANDN U9746 ( .A(n9463), .B(n9462), .Z(n9467) );
  NAND U9747 ( .A(n9465), .B(n9464), .Z(n9466) );
  AND U9748 ( .A(n9467), .B(n9466), .Z(n9515) );
  XOR U9749 ( .A(n9516), .B(n9515), .Z(n9517) );
  NANDN U9750 ( .A(n9469), .B(n9468), .Z(n9473) );
  NANDN U9751 ( .A(n9471), .B(n9470), .Z(n9472) );
  NAND U9752 ( .A(n9473), .B(n9472), .Z(n9518) );
  XOR U9753 ( .A(n9517), .B(n9518), .Z(n9485) );
  OR U9754 ( .A(n9475), .B(n9474), .Z(n9479) );
  NANDN U9755 ( .A(n9477), .B(n9476), .Z(n9478) );
  NAND U9756 ( .A(n9479), .B(n9478), .Z(n9486) );
  XNOR U9757 ( .A(n9485), .B(n9486), .Z(n9487) );
  XNOR U9758 ( .A(n9488), .B(n9487), .Z(n9521) );
  XNOR U9759 ( .A(n9521), .B(sreg[1245]), .Z(n9523) );
  NAND U9760 ( .A(n9480), .B(sreg[1244]), .Z(n9484) );
  OR U9761 ( .A(n9482), .B(n9481), .Z(n9483) );
  AND U9762 ( .A(n9484), .B(n9483), .Z(n9522) );
  XOR U9763 ( .A(n9523), .B(n9522), .Z(c[1245]) );
  NANDN U9764 ( .A(n9486), .B(n9485), .Z(n9490) );
  NAND U9765 ( .A(n9488), .B(n9487), .Z(n9489) );
  NAND U9766 ( .A(n9490), .B(n9489), .Z(n9529) );
  NAND U9767 ( .A(b[0]), .B(a[230]), .Z(n9491) );
  XNOR U9768 ( .A(b[1]), .B(n9491), .Z(n9493) );
  NAND U9769 ( .A(n47), .B(a[229]), .Z(n9492) );
  AND U9770 ( .A(n9493), .B(n9492), .Z(n9546) );
  XOR U9771 ( .A(a[226]), .B(n42197), .Z(n9535) );
  NANDN U9772 ( .A(n9535), .B(n42173), .Z(n9496) );
  NANDN U9773 ( .A(n9494), .B(n42172), .Z(n9495) );
  NAND U9774 ( .A(n9496), .B(n9495), .Z(n9544) );
  NAND U9775 ( .A(b[7]), .B(a[222]), .Z(n9545) );
  XNOR U9776 ( .A(n9544), .B(n9545), .Z(n9547) );
  XOR U9777 ( .A(n9546), .B(n9547), .Z(n9553) );
  NANDN U9778 ( .A(n9497), .B(n42093), .Z(n9499) );
  XOR U9779 ( .A(n42134), .B(a[228]), .Z(n9538) );
  NANDN U9780 ( .A(n9538), .B(n42095), .Z(n9498) );
  NAND U9781 ( .A(n9499), .B(n9498), .Z(n9551) );
  NANDN U9782 ( .A(n9500), .B(n42231), .Z(n9502) );
  XOR U9783 ( .A(n180), .B(a[224]), .Z(n9541) );
  NANDN U9784 ( .A(n9541), .B(n42234), .Z(n9501) );
  AND U9785 ( .A(n9502), .B(n9501), .Z(n9550) );
  XNOR U9786 ( .A(n9551), .B(n9550), .Z(n9552) );
  XNOR U9787 ( .A(n9553), .B(n9552), .Z(n9557) );
  NANDN U9788 ( .A(n9504), .B(n9503), .Z(n9508) );
  NAND U9789 ( .A(n9506), .B(n9505), .Z(n9507) );
  AND U9790 ( .A(n9508), .B(n9507), .Z(n9556) );
  XOR U9791 ( .A(n9557), .B(n9556), .Z(n9558) );
  NANDN U9792 ( .A(n9510), .B(n9509), .Z(n9514) );
  NANDN U9793 ( .A(n9512), .B(n9511), .Z(n9513) );
  NAND U9794 ( .A(n9514), .B(n9513), .Z(n9559) );
  XOR U9795 ( .A(n9558), .B(n9559), .Z(n9526) );
  OR U9796 ( .A(n9516), .B(n9515), .Z(n9520) );
  NANDN U9797 ( .A(n9518), .B(n9517), .Z(n9519) );
  NAND U9798 ( .A(n9520), .B(n9519), .Z(n9527) );
  XNOR U9799 ( .A(n9526), .B(n9527), .Z(n9528) );
  XNOR U9800 ( .A(n9529), .B(n9528), .Z(n9562) );
  XNOR U9801 ( .A(n9562), .B(sreg[1246]), .Z(n9564) );
  NAND U9802 ( .A(n9521), .B(sreg[1245]), .Z(n9525) );
  OR U9803 ( .A(n9523), .B(n9522), .Z(n9524) );
  AND U9804 ( .A(n9525), .B(n9524), .Z(n9563) );
  XOR U9805 ( .A(n9564), .B(n9563), .Z(c[1246]) );
  NANDN U9806 ( .A(n9527), .B(n9526), .Z(n9531) );
  NAND U9807 ( .A(n9529), .B(n9528), .Z(n9530) );
  NAND U9808 ( .A(n9531), .B(n9530), .Z(n9570) );
  NAND U9809 ( .A(b[0]), .B(a[231]), .Z(n9532) );
  XNOR U9810 ( .A(b[1]), .B(n9532), .Z(n9534) );
  NAND U9811 ( .A(n48), .B(a[230]), .Z(n9533) );
  AND U9812 ( .A(n9534), .B(n9533), .Z(n9587) );
  XOR U9813 ( .A(a[227]), .B(n42197), .Z(n9576) );
  NANDN U9814 ( .A(n9576), .B(n42173), .Z(n9537) );
  NANDN U9815 ( .A(n9535), .B(n42172), .Z(n9536) );
  NAND U9816 ( .A(n9537), .B(n9536), .Z(n9585) );
  NAND U9817 ( .A(b[7]), .B(a[223]), .Z(n9586) );
  XNOR U9818 ( .A(n9585), .B(n9586), .Z(n9588) );
  XOR U9819 ( .A(n9587), .B(n9588), .Z(n9594) );
  NANDN U9820 ( .A(n9538), .B(n42093), .Z(n9540) );
  XOR U9821 ( .A(n42134), .B(a[229]), .Z(n9579) );
  NANDN U9822 ( .A(n9579), .B(n42095), .Z(n9539) );
  NAND U9823 ( .A(n9540), .B(n9539), .Z(n9592) );
  NANDN U9824 ( .A(n9541), .B(n42231), .Z(n9543) );
  XOR U9825 ( .A(n180), .B(a[225]), .Z(n9582) );
  NANDN U9826 ( .A(n9582), .B(n42234), .Z(n9542) );
  AND U9827 ( .A(n9543), .B(n9542), .Z(n9591) );
  XNOR U9828 ( .A(n9592), .B(n9591), .Z(n9593) );
  XNOR U9829 ( .A(n9594), .B(n9593), .Z(n9598) );
  NANDN U9830 ( .A(n9545), .B(n9544), .Z(n9549) );
  NAND U9831 ( .A(n9547), .B(n9546), .Z(n9548) );
  AND U9832 ( .A(n9549), .B(n9548), .Z(n9597) );
  XOR U9833 ( .A(n9598), .B(n9597), .Z(n9599) );
  NANDN U9834 ( .A(n9551), .B(n9550), .Z(n9555) );
  NANDN U9835 ( .A(n9553), .B(n9552), .Z(n9554) );
  NAND U9836 ( .A(n9555), .B(n9554), .Z(n9600) );
  XOR U9837 ( .A(n9599), .B(n9600), .Z(n9567) );
  OR U9838 ( .A(n9557), .B(n9556), .Z(n9561) );
  NANDN U9839 ( .A(n9559), .B(n9558), .Z(n9560) );
  NAND U9840 ( .A(n9561), .B(n9560), .Z(n9568) );
  XNOR U9841 ( .A(n9567), .B(n9568), .Z(n9569) );
  XNOR U9842 ( .A(n9570), .B(n9569), .Z(n9603) );
  XNOR U9843 ( .A(n9603), .B(sreg[1247]), .Z(n9605) );
  NAND U9844 ( .A(n9562), .B(sreg[1246]), .Z(n9566) );
  OR U9845 ( .A(n9564), .B(n9563), .Z(n9565) );
  AND U9846 ( .A(n9566), .B(n9565), .Z(n9604) );
  XOR U9847 ( .A(n9605), .B(n9604), .Z(c[1247]) );
  NANDN U9848 ( .A(n9568), .B(n9567), .Z(n9572) );
  NAND U9849 ( .A(n9570), .B(n9569), .Z(n9571) );
  NAND U9850 ( .A(n9572), .B(n9571), .Z(n9611) );
  NAND U9851 ( .A(b[0]), .B(a[232]), .Z(n9573) );
  XNOR U9852 ( .A(b[1]), .B(n9573), .Z(n9575) );
  NAND U9853 ( .A(n48), .B(a[231]), .Z(n9574) );
  AND U9854 ( .A(n9575), .B(n9574), .Z(n9628) );
  XOR U9855 ( .A(a[228]), .B(n42197), .Z(n9617) );
  NANDN U9856 ( .A(n9617), .B(n42173), .Z(n9578) );
  NANDN U9857 ( .A(n9576), .B(n42172), .Z(n9577) );
  NAND U9858 ( .A(n9578), .B(n9577), .Z(n9626) );
  NAND U9859 ( .A(b[7]), .B(a[224]), .Z(n9627) );
  XNOR U9860 ( .A(n9626), .B(n9627), .Z(n9629) );
  XOR U9861 ( .A(n9628), .B(n9629), .Z(n9635) );
  NANDN U9862 ( .A(n9579), .B(n42093), .Z(n9581) );
  XOR U9863 ( .A(n42134), .B(a[230]), .Z(n9620) );
  NANDN U9864 ( .A(n9620), .B(n42095), .Z(n9580) );
  NAND U9865 ( .A(n9581), .B(n9580), .Z(n9633) );
  NANDN U9866 ( .A(n9582), .B(n42231), .Z(n9584) );
  XOR U9867 ( .A(n180), .B(a[226]), .Z(n9623) );
  NANDN U9868 ( .A(n9623), .B(n42234), .Z(n9583) );
  AND U9869 ( .A(n9584), .B(n9583), .Z(n9632) );
  XNOR U9870 ( .A(n9633), .B(n9632), .Z(n9634) );
  XNOR U9871 ( .A(n9635), .B(n9634), .Z(n9639) );
  NANDN U9872 ( .A(n9586), .B(n9585), .Z(n9590) );
  NAND U9873 ( .A(n9588), .B(n9587), .Z(n9589) );
  AND U9874 ( .A(n9590), .B(n9589), .Z(n9638) );
  XOR U9875 ( .A(n9639), .B(n9638), .Z(n9640) );
  NANDN U9876 ( .A(n9592), .B(n9591), .Z(n9596) );
  NANDN U9877 ( .A(n9594), .B(n9593), .Z(n9595) );
  NAND U9878 ( .A(n9596), .B(n9595), .Z(n9641) );
  XOR U9879 ( .A(n9640), .B(n9641), .Z(n9608) );
  OR U9880 ( .A(n9598), .B(n9597), .Z(n9602) );
  NANDN U9881 ( .A(n9600), .B(n9599), .Z(n9601) );
  NAND U9882 ( .A(n9602), .B(n9601), .Z(n9609) );
  XNOR U9883 ( .A(n9608), .B(n9609), .Z(n9610) );
  XNOR U9884 ( .A(n9611), .B(n9610), .Z(n9644) );
  XNOR U9885 ( .A(n9644), .B(sreg[1248]), .Z(n9646) );
  NAND U9886 ( .A(n9603), .B(sreg[1247]), .Z(n9607) );
  OR U9887 ( .A(n9605), .B(n9604), .Z(n9606) );
  AND U9888 ( .A(n9607), .B(n9606), .Z(n9645) );
  XOR U9889 ( .A(n9646), .B(n9645), .Z(c[1248]) );
  NANDN U9890 ( .A(n9609), .B(n9608), .Z(n9613) );
  NAND U9891 ( .A(n9611), .B(n9610), .Z(n9612) );
  NAND U9892 ( .A(n9613), .B(n9612), .Z(n9652) );
  NAND U9893 ( .A(b[0]), .B(a[233]), .Z(n9614) );
  XNOR U9894 ( .A(b[1]), .B(n9614), .Z(n9616) );
  NAND U9895 ( .A(n48), .B(a[232]), .Z(n9615) );
  AND U9896 ( .A(n9616), .B(n9615), .Z(n9669) );
  XOR U9897 ( .A(a[229]), .B(n42197), .Z(n9658) );
  NANDN U9898 ( .A(n9658), .B(n42173), .Z(n9619) );
  NANDN U9899 ( .A(n9617), .B(n42172), .Z(n9618) );
  NAND U9900 ( .A(n9619), .B(n9618), .Z(n9667) );
  NAND U9901 ( .A(b[7]), .B(a[225]), .Z(n9668) );
  XNOR U9902 ( .A(n9667), .B(n9668), .Z(n9670) );
  XOR U9903 ( .A(n9669), .B(n9670), .Z(n9676) );
  NANDN U9904 ( .A(n9620), .B(n42093), .Z(n9622) );
  XOR U9905 ( .A(n42134), .B(a[231]), .Z(n9661) );
  NANDN U9906 ( .A(n9661), .B(n42095), .Z(n9621) );
  NAND U9907 ( .A(n9622), .B(n9621), .Z(n9674) );
  NANDN U9908 ( .A(n9623), .B(n42231), .Z(n9625) );
  XOR U9909 ( .A(n181), .B(a[227]), .Z(n9664) );
  NANDN U9910 ( .A(n9664), .B(n42234), .Z(n9624) );
  AND U9911 ( .A(n9625), .B(n9624), .Z(n9673) );
  XNOR U9912 ( .A(n9674), .B(n9673), .Z(n9675) );
  XNOR U9913 ( .A(n9676), .B(n9675), .Z(n9680) );
  NANDN U9914 ( .A(n9627), .B(n9626), .Z(n9631) );
  NAND U9915 ( .A(n9629), .B(n9628), .Z(n9630) );
  AND U9916 ( .A(n9631), .B(n9630), .Z(n9679) );
  XOR U9917 ( .A(n9680), .B(n9679), .Z(n9681) );
  NANDN U9918 ( .A(n9633), .B(n9632), .Z(n9637) );
  NANDN U9919 ( .A(n9635), .B(n9634), .Z(n9636) );
  NAND U9920 ( .A(n9637), .B(n9636), .Z(n9682) );
  XOR U9921 ( .A(n9681), .B(n9682), .Z(n9649) );
  OR U9922 ( .A(n9639), .B(n9638), .Z(n9643) );
  NANDN U9923 ( .A(n9641), .B(n9640), .Z(n9642) );
  NAND U9924 ( .A(n9643), .B(n9642), .Z(n9650) );
  XNOR U9925 ( .A(n9649), .B(n9650), .Z(n9651) );
  XNOR U9926 ( .A(n9652), .B(n9651), .Z(n9685) );
  XNOR U9927 ( .A(n9685), .B(sreg[1249]), .Z(n9687) );
  NAND U9928 ( .A(n9644), .B(sreg[1248]), .Z(n9648) );
  OR U9929 ( .A(n9646), .B(n9645), .Z(n9647) );
  AND U9930 ( .A(n9648), .B(n9647), .Z(n9686) );
  XOR U9931 ( .A(n9687), .B(n9686), .Z(c[1249]) );
  NANDN U9932 ( .A(n9650), .B(n9649), .Z(n9654) );
  NAND U9933 ( .A(n9652), .B(n9651), .Z(n9653) );
  NAND U9934 ( .A(n9654), .B(n9653), .Z(n9693) );
  NAND U9935 ( .A(b[0]), .B(a[234]), .Z(n9655) );
  XNOR U9936 ( .A(b[1]), .B(n9655), .Z(n9657) );
  NAND U9937 ( .A(n48), .B(a[233]), .Z(n9656) );
  AND U9938 ( .A(n9657), .B(n9656), .Z(n9710) );
  XOR U9939 ( .A(a[230]), .B(n42197), .Z(n9699) );
  NANDN U9940 ( .A(n9699), .B(n42173), .Z(n9660) );
  NANDN U9941 ( .A(n9658), .B(n42172), .Z(n9659) );
  NAND U9942 ( .A(n9660), .B(n9659), .Z(n9708) );
  NAND U9943 ( .A(b[7]), .B(a[226]), .Z(n9709) );
  XNOR U9944 ( .A(n9708), .B(n9709), .Z(n9711) );
  XOR U9945 ( .A(n9710), .B(n9711), .Z(n9717) );
  NANDN U9946 ( .A(n9661), .B(n42093), .Z(n9663) );
  XOR U9947 ( .A(n42134), .B(a[232]), .Z(n9702) );
  NANDN U9948 ( .A(n9702), .B(n42095), .Z(n9662) );
  NAND U9949 ( .A(n9663), .B(n9662), .Z(n9715) );
  NANDN U9950 ( .A(n9664), .B(n42231), .Z(n9666) );
  XOR U9951 ( .A(n181), .B(a[228]), .Z(n9705) );
  NANDN U9952 ( .A(n9705), .B(n42234), .Z(n9665) );
  AND U9953 ( .A(n9666), .B(n9665), .Z(n9714) );
  XNOR U9954 ( .A(n9715), .B(n9714), .Z(n9716) );
  XNOR U9955 ( .A(n9717), .B(n9716), .Z(n9721) );
  NANDN U9956 ( .A(n9668), .B(n9667), .Z(n9672) );
  NAND U9957 ( .A(n9670), .B(n9669), .Z(n9671) );
  AND U9958 ( .A(n9672), .B(n9671), .Z(n9720) );
  XOR U9959 ( .A(n9721), .B(n9720), .Z(n9722) );
  NANDN U9960 ( .A(n9674), .B(n9673), .Z(n9678) );
  NANDN U9961 ( .A(n9676), .B(n9675), .Z(n9677) );
  NAND U9962 ( .A(n9678), .B(n9677), .Z(n9723) );
  XOR U9963 ( .A(n9722), .B(n9723), .Z(n9690) );
  OR U9964 ( .A(n9680), .B(n9679), .Z(n9684) );
  NANDN U9965 ( .A(n9682), .B(n9681), .Z(n9683) );
  NAND U9966 ( .A(n9684), .B(n9683), .Z(n9691) );
  XNOR U9967 ( .A(n9690), .B(n9691), .Z(n9692) );
  XNOR U9968 ( .A(n9693), .B(n9692), .Z(n9726) );
  XNOR U9969 ( .A(n9726), .B(sreg[1250]), .Z(n9728) );
  NAND U9970 ( .A(n9685), .B(sreg[1249]), .Z(n9689) );
  OR U9971 ( .A(n9687), .B(n9686), .Z(n9688) );
  AND U9972 ( .A(n9689), .B(n9688), .Z(n9727) );
  XOR U9973 ( .A(n9728), .B(n9727), .Z(c[1250]) );
  NANDN U9974 ( .A(n9691), .B(n9690), .Z(n9695) );
  NAND U9975 ( .A(n9693), .B(n9692), .Z(n9694) );
  NAND U9976 ( .A(n9695), .B(n9694), .Z(n9734) );
  NAND U9977 ( .A(b[0]), .B(a[235]), .Z(n9696) );
  XNOR U9978 ( .A(b[1]), .B(n9696), .Z(n9698) );
  NAND U9979 ( .A(n48), .B(a[234]), .Z(n9697) );
  AND U9980 ( .A(n9698), .B(n9697), .Z(n9751) );
  XOR U9981 ( .A(a[231]), .B(n42197), .Z(n9740) );
  NANDN U9982 ( .A(n9740), .B(n42173), .Z(n9701) );
  NANDN U9983 ( .A(n9699), .B(n42172), .Z(n9700) );
  NAND U9984 ( .A(n9701), .B(n9700), .Z(n9749) );
  NAND U9985 ( .A(b[7]), .B(a[227]), .Z(n9750) );
  XNOR U9986 ( .A(n9749), .B(n9750), .Z(n9752) );
  XOR U9987 ( .A(n9751), .B(n9752), .Z(n9758) );
  NANDN U9988 ( .A(n9702), .B(n42093), .Z(n9704) );
  XOR U9989 ( .A(n42134), .B(a[233]), .Z(n9743) );
  NANDN U9990 ( .A(n9743), .B(n42095), .Z(n9703) );
  NAND U9991 ( .A(n9704), .B(n9703), .Z(n9756) );
  NANDN U9992 ( .A(n9705), .B(n42231), .Z(n9707) );
  XOR U9993 ( .A(n181), .B(a[229]), .Z(n9746) );
  NANDN U9994 ( .A(n9746), .B(n42234), .Z(n9706) );
  AND U9995 ( .A(n9707), .B(n9706), .Z(n9755) );
  XNOR U9996 ( .A(n9756), .B(n9755), .Z(n9757) );
  XNOR U9997 ( .A(n9758), .B(n9757), .Z(n9762) );
  NANDN U9998 ( .A(n9709), .B(n9708), .Z(n9713) );
  NAND U9999 ( .A(n9711), .B(n9710), .Z(n9712) );
  AND U10000 ( .A(n9713), .B(n9712), .Z(n9761) );
  XOR U10001 ( .A(n9762), .B(n9761), .Z(n9763) );
  NANDN U10002 ( .A(n9715), .B(n9714), .Z(n9719) );
  NANDN U10003 ( .A(n9717), .B(n9716), .Z(n9718) );
  NAND U10004 ( .A(n9719), .B(n9718), .Z(n9764) );
  XOR U10005 ( .A(n9763), .B(n9764), .Z(n9731) );
  OR U10006 ( .A(n9721), .B(n9720), .Z(n9725) );
  NANDN U10007 ( .A(n9723), .B(n9722), .Z(n9724) );
  NAND U10008 ( .A(n9725), .B(n9724), .Z(n9732) );
  XNOR U10009 ( .A(n9731), .B(n9732), .Z(n9733) );
  XNOR U10010 ( .A(n9734), .B(n9733), .Z(n9767) );
  XNOR U10011 ( .A(n9767), .B(sreg[1251]), .Z(n9769) );
  NAND U10012 ( .A(n9726), .B(sreg[1250]), .Z(n9730) );
  OR U10013 ( .A(n9728), .B(n9727), .Z(n9729) );
  AND U10014 ( .A(n9730), .B(n9729), .Z(n9768) );
  XOR U10015 ( .A(n9769), .B(n9768), .Z(c[1251]) );
  NANDN U10016 ( .A(n9732), .B(n9731), .Z(n9736) );
  NAND U10017 ( .A(n9734), .B(n9733), .Z(n9735) );
  NAND U10018 ( .A(n9736), .B(n9735), .Z(n9775) );
  NAND U10019 ( .A(b[0]), .B(a[236]), .Z(n9737) );
  XNOR U10020 ( .A(b[1]), .B(n9737), .Z(n9739) );
  NAND U10021 ( .A(n48), .B(a[235]), .Z(n9738) );
  AND U10022 ( .A(n9739), .B(n9738), .Z(n9792) );
  XOR U10023 ( .A(a[232]), .B(n42197), .Z(n9781) );
  NANDN U10024 ( .A(n9781), .B(n42173), .Z(n9742) );
  NANDN U10025 ( .A(n9740), .B(n42172), .Z(n9741) );
  NAND U10026 ( .A(n9742), .B(n9741), .Z(n9790) );
  NAND U10027 ( .A(b[7]), .B(a[228]), .Z(n9791) );
  XNOR U10028 ( .A(n9790), .B(n9791), .Z(n9793) );
  XOR U10029 ( .A(n9792), .B(n9793), .Z(n9799) );
  NANDN U10030 ( .A(n9743), .B(n42093), .Z(n9745) );
  XOR U10031 ( .A(n42134), .B(a[234]), .Z(n9784) );
  NANDN U10032 ( .A(n9784), .B(n42095), .Z(n9744) );
  NAND U10033 ( .A(n9745), .B(n9744), .Z(n9797) );
  NANDN U10034 ( .A(n9746), .B(n42231), .Z(n9748) );
  XOR U10035 ( .A(n181), .B(a[230]), .Z(n9787) );
  NANDN U10036 ( .A(n9787), .B(n42234), .Z(n9747) );
  AND U10037 ( .A(n9748), .B(n9747), .Z(n9796) );
  XNOR U10038 ( .A(n9797), .B(n9796), .Z(n9798) );
  XNOR U10039 ( .A(n9799), .B(n9798), .Z(n9803) );
  NANDN U10040 ( .A(n9750), .B(n9749), .Z(n9754) );
  NAND U10041 ( .A(n9752), .B(n9751), .Z(n9753) );
  AND U10042 ( .A(n9754), .B(n9753), .Z(n9802) );
  XOR U10043 ( .A(n9803), .B(n9802), .Z(n9804) );
  NANDN U10044 ( .A(n9756), .B(n9755), .Z(n9760) );
  NANDN U10045 ( .A(n9758), .B(n9757), .Z(n9759) );
  NAND U10046 ( .A(n9760), .B(n9759), .Z(n9805) );
  XOR U10047 ( .A(n9804), .B(n9805), .Z(n9772) );
  OR U10048 ( .A(n9762), .B(n9761), .Z(n9766) );
  NANDN U10049 ( .A(n9764), .B(n9763), .Z(n9765) );
  NAND U10050 ( .A(n9766), .B(n9765), .Z(n9773) );
  XNOR U10051 ( .A(n9772), .B(n9773), .Z(n9774) );
  XNOR U10052 ( .A(n9775), .B(n9774), .Z(n9808) );
  XNOR U10053 ( .A(n9808), .B(sreg[1252]), .Z(n9810) );
  NAND U10054 ( .A(n9767), .B(sreg[1251]), .Z(n9771) );
  OR U10055 ( .A(n9769), .B(n9768), .Z(n9770) );
  AND U10056 ( .A(n9771), .B(n9770), .Z(n9809) );
  XOR U10057 ( .A(n9810), .B(n9809), .Z(c[1252]) );
  NANDN U10058 ( .A(n9773), .B(n9772), .Z(n9777) );
  NAND U10059 ( .A(n9775), .B(n9774), .Z(n9776) );
  NAND U10060 ( .A(n9777), .B(n9776), .Z(n9816) );
  NAND U10061 ( .A(b[0]), .B(a[237]), .Z(n9778) );
  XNOR U10062 ( .A(b[1]), .B(n9778), .Z(n9780) );
  NAND U10063 ( .A(n48), .B(a[236]), .Z(n9779) );
  AND U10064 ( .A(n9780), .B(n9779), .Z(n9833) );
  XOR U10065 ( .A(a[233]), .B(n42197), .Z(n9822) );
  NANDN U10066 ( .A(n9822), .B(n42173), .Z(n9783) );
  NANDN U10067 ( .A(n9781), .B(n42172), .Z(n9782) );
  NAND U10068 ( .A(n9783), .B(n9782), .Z(n9831) );
  NAND U10069 ( .A(b[7]), .B(a[229]), .Z(n9832) );
  XNOR U10070 ( .A(n9831), .B(n9832), .Z(n9834) );
  XOR U10071 ( .A(n9833), .B(n9834), .Z(n9840) );
  NANDN U10072 ( .A(n9784), .B(n42093), .Z(n9786) );
  XOR U10073 ( .A(n42134), .B(a[235]), .Z(n9825) );
  NANDN U10074 ( .A(n9825), .B(n42095), .Z(n9785) );
  NAND U10075 ( .A(n9786), .B(n9785), .Z(n9838) );
  NANDN U10076 ( .A(n9787), .B(n42231), .Z(n9789) );
  XOR U10077 ( .A(n181), .B(a[231]), .Z(n9828) );
  NANDN U10078 ( .A(n9828), .B(n42234), .Z(n9788) );
  AND U10079 ( .A(n9789), .B(n9788), .Z(n9837) );
  XNOR U10080 ( .A(n9838), .B(n9837), .Z(n9839) );
  XNOR U10081 ( .A(n9840), .B(n9839), .Z(n9844) );
  NANDN U10082 ( .A(n9791), .B(n9790), .Z(n9795) );
  NAND U10083 ( .A(n9793), .B(n9792), .Z(n9794) );
  AND U10084 ( .A(n9795), .B(n9794), .Z(n9843) );
  XOR U10085 ( .A(n9844), .B(n9843), .Z(n9845) );
  NANDN U10086 ( .A(n9797), .B(n9796), .Z(n9801) );
  NANDN U10087 ( .A(n9799), .B(n9798), .Z(n9800) );
  NAND U10088 ( .A(n9801), .B(n9800), .Z(n9846) );
  XOR U10089 ( .A(n9845), .B(n9846), .Z(n9813) );
  OR U10090 ( .A(n9803), .B(n9802), .Z(n9807) );
  NANDN U10091 ( .A(n9805), .B(n9804), .Z(n9806) );
  NAND U10092 ( .A(n9807), .B(n9806), .Z(n9814) );
  XNOR U10093 ( .A(n9813), .B(n9814), .Z(n9815) );
  XNOR U10094 ( .A(n9816), .B(n9815), .Z(n9849) );
  XNOR U10095 ( .A(n9849), .B(sreg[1253]), .Z(n9851) );
  NAND U10096 ( .A(n9808), .B(sreg[1252]), .Z(n9812) );
  OR U10097 ( .A(n9810), .B(n9809), .Z(n9811) );
  AND U10098 ( .A(n9812), .B(n9811), .Z(n9850) );
  XOR U10099 ( .A(n9851), .B(n9850), .Z(c[1253]) );
  NANDN U10100 ( .A(n9814), .B(n9813), .Z(n9818) );
  NAND U10101 ( .A(n9816), .B(n9815), .Z(n9817) );
  NAND U10102 ( .A(n9818), .B(n9817), .Z(n9857) );
  NAND U10103 ( .A(b[0]), .B(a[238]), .Z(n9819) );
  XNOR U10104 ( .A(b[1]), .B(n9819), .Z(n9821) );
  NAND U10105 ( .A(n49), .B(a[237]), .Z(n9820) );
  AND U10106 ( .A(n9821), .B(n9820), .Z(n9874) );
  XOR U10107 ( .A(a[234]), .B(n42197), .Z(n9863) );
  NANDN U10108 ( .A(n9863), .B(n42173), .Z(n9824) );
  NANDN U10109 ( .A(n9822), .B(n42172), .Z(n9823) );
  NAND U10110 ( .A(n9824), .B(n9823), .Z(n9872) );
  NAND U10111 ( .A(b[7]), .B(a[230]), .Z(n9873) );
  XNOR U10112 ( .A(n9872), .B(n9873), .Z(n9875) );
  XOR U10113 ( .A(n9874), .B(n9875), .Z(n9881) );
  NANDN U10114 ( .A(n9825), .B(n42093), .Z(n9827) );
  XOR U10115 ( .A(n42134), .B(a[236]), .Z(n9866) );
  NANDN U10116 ( .A(n9866), .B(n42095), .Z(n9826) );
  NAND U10117 ( .A(n9827), .B(n9826), .Z(n9879) );
  NANDN U10118 ( .A(n9828), .B(n42231), .Z(n9830) );
  XOR U10119 ( .A(n181), .B(a[232]), .Z(n9869) );
  NANDN U10120 ( .A(n9869), .B(n42234), .Z(n9829) );
  AND U10121 ( .A(n9830), .B(n9829), .Z(n9878) );
  XNOR U10122 ( .A(n9879), .B(n9878), .Z(n9880) );
  XNOR U10123 ( .A(n9881), .B(n9880), .Z(n9885) );
  NANDN U10124 ( .A(n9832), .B(n9831), .Z(n9836) );
  NAND U10125 ( .A(n9834), .B(n9833), .Z(n9835) );
  AND U10126 ( .A(n9836), .B(n9835), .Z(n9884) );
  XOR U10127 ( .A(n9885), .B(n9884), .Z(n9886) );
  NANDN U10128 ( .A(n9838), .B(n9837), .Z(n9842) );
  NANDN U10129 ( .A(n9840), .B(n9839), .Z(n9841) );
  NAND U10130 ( .A(n9842), .B(n9841), .Z(n9887) );
  XOR U10131 ( .A(n9886), .B(n9887), .Z(n9854) );
  OR U10132 ( .A(n9844), .B(n9843), .Z(n9848) );
  NANDN U10133 ( .A(n9846), .B(n9845), .Z(n9847) );
  NAND U10134 ( .A(n9848), .B(n9847), .Z(n9855) );
  XNOR U10135 ( .A(n9854), .B(n9855), .Z(n9856) );
  XNOR U10136 ( .A(n9857), .B(n9856), .Z(n9890) );
  XNOR U10137 ( .A(n9890), .B(sreg[1254]), .Z(n9892) );
  NAND U10138 ( .A(n9849), .B(sreg[1253]), .Z(n9853) );
  OR U10139 ( .A(n9851), .B(n9850), .Z(n9852) );
  AND U10140 ( .A(n9853), .B(n9852), .Z(n9891) );
  XOR U10141 ( .A(n9892), .B(n9891), .Z(c[1254]) );
  NANDN U10142 ( .A(n9855), .B(n9854), .Z(n9859) );
  NAND U10143 ( .A(n9857), .B(n9856), .Z(n9858) );
  NAND U10144 ( .A(n9859), .B(n9858), .Z(n9898) );
  NAND U10145 ( .A(b[0]), .B(a[239]), .Z(n9860) );
  XNOR U10146 ( .A(b[1]), .B(n9860), .Z(n9862) );
  NAND U10147 ( .A(n49), .B(a[238]), .Z(n9861) );
  AND U10148 ( .A(n9862), .B(n9861), .Z(n9915) );
  XOR U10149 ( .A(a[235]), .B(n42197), .Z(n9904) );
  NANDN U10150 ( .A(n9904), .B(n42173), .Z(n9865) );
  NANDN U10151 ( .A(n9863), .B(n42172), .Z(n9864) );
  NAND U10152 ( .A(n9865), .B(n9864), .Z(n9913) );
  NAND U10153 ( .A(b[7]), .B(a[231]), .Z(n9914) );
  XNOR U10154 ( .A(n9913), .B(n9914), .Z(n9916) );
  XOR U10155 ( .A(n9915), .B(n9916), .Z(n9922) );
  NANDN U10156 ( .A(n9866), .B(n42093), .Z(n9868) );
  XOR U10157 ( .A(n42134), .B(a[237]), .Z(n9907) );
  NANDN U10158 ( .A(n9907), .B(n42095), .Z(n9867) );
  NAND U10159 ( .A(n9868), .B(n9867), .Z(n9920) );
  NANDN U10160 ( .A(n9869), .B(n42231), .Z(n9871) );
  XOR U10161 ( .A(n181), .B(a[233]), .Z(n9910) );
  NANDN U10162 ( .A(n9910), .B(n42234), .Z(n9870) );
  AND U10163 ( .A(n9871), .B(n9870), .Z(n9919) );
  XNOR U10164 ( .A(n9920), .B(n9919), .Z(n9921) );
  XNOR U10165 ( .A(n9922), .B(n9921), .Z(n9926) );
  NANDN U10166 ( .A(n9873), .B(n9872), .Z(n9877) );
  NAND U10167 ( .A(n9875), .B(n9874), .Z(n9876) );
  AND U10168 ( .A(n9877), .B(n9876), .Z(n9925) );
  XOR U10169 ( .A(n9926), .B(n9925), .Z(n9927) );
  NANDN U10170 ( .A(n9879), .B(n9878), .Z(n9883) );
  NANDN U10171 ( .A(n9881), .B(n9880), .Z(n9882) );
  NAND U10172 ( .A(n9883), .B(n9882), .Z(n9928) );
  XOR U10173 ( .A(n9927), .B(n9928), .Z(n9895) );
  OR U10174 ( .A(n9885), .B(n9884), .Z(n9889) );
  NANDN U10175 ( .A(n9887), .B(n9886), .Z(n9888) );
  NAND U10176 ( .A(n9889), .B(n9888), .Z(n9896) );
  XNOR U10177 ( .A(n9895), .B(n9896), .Z(n9897) );
  XNOR U10178 ( .A(n9898), .B(n9897), .Z(n9931) );
  XNOR U10179 ( .A(n9931), .B(sreg[1255]), .Z(n9933) );
  NAND U10180 ( .A(n9890), .B(sreg[1254]), .Z(n9894) );
  OR U10181 ( .A(n9892), .B(n9891), .Z(n9893) );
  AND U10182 ( .A(n9894), .B(n9893), .Z(n9932) );
  XOR U10183 ( .A(n9933), .B(n9932), .Z(c[1255]) );
  NANDN U10184 ( .A(n9896), .B(n9895), .Z(n9900) );
  NAND U10185 ( .A(n9898), .B(n9897), .Z(n9899) );
  NAND U10186 ( .A(n9900), .B(n9899), .Z(n9939) );
  NAND U10187 ( .A(b[0]), .B(a[240]), .Z(n9901) );
  XNOR U10188 ( .A(b[1]), .B(n9901), .Z(n9903) );
  NAND U10189 ( .A(n49), .B(a[239]), .Z(n9902) );
  AND U10190 ( .A(n9903), .B(n9902), .Z(n9956) );
  XOR U10191 ( .A(a[236]), .B(n42197), .Z(n9945) );
  NANDN U10192 ( .A(n9945), .B(n42173), .Z(n9906) );
  NANDN U10193 ( .A(n9904), .B(n42172), .Z(n9905) );
  NAND U10194 ( .A(n9906), .B(n9905), .Z(n9954) );
  NAND U10195 ( .A(b[7]), .B(a[232]), .Z(n9955) );
  XNOR U10196 ( .A(n9954), .B(n9955), .Z(n9957) );
  XOR U10197 ( .A(n9956), .B(n9957), .Z(n9963) );
  NANDN U10198 ( .A(n9907), .B(n42093), .Z(n9909) );
  XOR U10199 ( .A(n42134), .B(a[238]), .Z(n9948) );
  NANDN U10200 ( .A(n9948), .B(n42095), .Z(n9908) );
  NAND U10201 ( .A(n9909), .B(n9908), .Z(n9961) );
  NANDN U10202 ( .A(n9910), .B(n42231), .Z(n9912) );
  XOR U10203 ( .A(n181), .B(a[234]), .Z(n9951) );
  NANDN U10204 ( .A(n9951), .B(n42234), .Z(n9911) );
  AND U10205 ( .A(n9912), .B(n9911), .Z(n9960) );
  XNOR U10206 ( .A(n9961), .B(n9960), .Z(n9962) );
  XNOR U10207 ( .A(n9963), .B(n9962), .Z(n9967) );
  NANDN U10208 ( .A(n9914), .B(n9913), .Z(n9918) );
  NAND U10209 ( .A(n9916), .B(n9915), .Z(n9917) );
  AND U10210 ( .A(n9918), .B(n9917), .Z(n9966) );
  XOR U10211 ( .A(n9967), .B(n9966), .Z(n9968) );
  NANDN U10212 ( .A(n9920), .B(n9919), .Z(n9924) );
  NANDN U10213 ( .A(n9922), .B(n9921), .Z(n9923) );
  NAND U10214 ( .A(n9924), .B(n9923), .Z(n9969) );
  XOR U10215 ( .A(n9968), .B(n9969), .Z(n9936) );
  OR U10216 ( .A(n9926), .B(n9925), .Z(n9930) );
  NANDN U10217 ( .A(n9928), .B(n9927), .Z(n9929) );
  NAND U10218 ( .A(n9930), .B(n9929), .Z(n9937) );
  XNOR U10219 ( .A(n9936), .B(n9937), .Z(n9938) );
  XNOR U10220 ( .A(n9939), .B(n9938), .Z(n9972) );
  XNOR U10221 ( .A(n9972), .B(sreg[1256]), .Z(n9974) );
  NAND U10222 ( .A(n9931), .B(sreg[1255]), .Z(n9935) );
  OR U10223 ( .A(n9933), .B(n9932), .Z(n9934) );
  AND U10224 ( .A(n9935), .B(n9934), .Z(n9973) );
  XOR U10225 ( .A(n9974), .B(n9973), .Z(c[1256]) );
  NANDN U10226 ( .A(n9937), .B(n9936), .Z(n9941) );
  NAND U10227 ( .A(n9939), .B(n9938), .Z(n9940) );
  NAND U10228 ( .A(n9941), .B(n9940), .Z(n9980) );
  NAND U10229 ( .A(b[0]), .B(a[241]), .Z(n9942) );
  XNOR U10230 ( .A(b[1]), .B(n9942), .Z(n9944) );
  NAND U10231 ( .A(n49), .B(a[240]), .Z(n9943) );
  AND U10232 ( .A(n9944), .B(n9943), .Z(n9997) );
  XOR U10233 ( .A(a[237]), .B(n42197), .Z(n9986) );
  NANDN U10234 ( .A(n9986), .B(n42173), .Z(n9947) );
  NANDN U10235 ( .A(n9945), .B(n42172), .Z(n9946) );
  NAND U10236 ( .A(n9947), .B(n9946), .Z(n9995) );
  NAND U10237 ( .A(b[7]), .B(a[233]), .Z(n9996) );
  XNOR U10238 ( .A(n9995), .B(n9996), .Z(n9998) );
  XOR U10239 ( .A(n9997), .B(n9998), .Z(n10004) );
  NANDN U10240 ( .A(n9948), .B(n42093), .Z(n9950) );
  XOR U10241 ( .A(n42134), .B(a[239]), .Z(n9989) );
  NANDN U10242 ( .A(n9989), .B(n42095), .Z(n9949) );
  NAND U10243 ( .A(n9950), .B(n9949), .Z(n10002) );
  NANDN U10244 ( .A(n9951), .B(n42231), .Z(n9953) );
  XOR U10245 ( .A(n181), .B(a[235]), .Z(n9992) );
  NANDN U10246 ( .A(n9992), .B(n42234), .Z(n9952) );
  AND U10247 ( .A(n9953), .B(n9952), .Z(n10001) );
  XNOR U10248 ( .A(n10002), .B(n10001), .Z(n10003) );
  XNOR U10249 ( .A(n10004), .B(n10003), .Z(n10008) );
  NANDN U10250 ( .A(n9955), .B(n9954), .Z(n9959) );
  NAND U10251 ( .A(n9957), .B(n9956), .Z(n9958) );
  AND U10252 ( .A(n9959), .B(n9958), .Z(n10007) );
  XOR U10253 ( .A(n10008), .B(n10007), .Z(n10009) );
  NANDN U10254 ( .A(n9961), .B(n9960), .Z(n9965) );
  NANDN U10255 ( .A(n9963), .B(n9962), .Z(n9964) );
  NAND U10256 ( .A(n9965), .B(n9964), .Z(n10010) );
  XOR U10257 ( .A(n10009), .B(n10010), .Z(n9977) );
  OR U10258 ( .A(n9967), .B(n9966), .Z(n9971) );
  NANDN U10259 ( .A(n9969), .B(n9968), .Z(n9970) );
  NAND U10260 ( .A(n9971), .B(n9970), .Z(n9978) );
  XNOR U10261 ( .A(n9977), .B(n9978), .Z(n9979) );
  XNOR U10262 ( .A(n9980), .B(n9979), .Z(n10013) );
  XNOR U10263 ( .A(n10013), .B(sreg[1257]), .Z(n10015) );
  NAND U10264 ( .A(n9972), .B(sreg[1256]), .Z(n9976) );
  OR U10265 ( .A(n9974), .B(n9973), .Z(n9975) );
  AND U10266 ( .A(n9976), .B(n9975), .Z(n10014) );
  XOR U10267 ( .A(n10015), .B(n10014), .Z(c[1257]) );
  NANDN U10268 ( .A(n9978), .B(n9977), .Z(n9982) );
  NAND U10269 ( .A(n9980), .B(n9979), .Z(n9981) );
  NAND U10270 ( .A(n9982), .B(n9981), .Z(n10021) );
  NAND U10271 ( .A(b[0]), .B(a[242]), .Z(n9983) );
  XNOR U10272 ( .A(b[1]), .B(n9983), .Z(n9985) );
  NAND U10273 ( .A(n49), .B(a[241]), .Z(n9984) );
  AND U10274 ( .A(n9985), .B(n9984), .Z(n10038) );
  XOR U10275 ( .A(a[238]), .B(n42197), .Z(n10027) );
  NANDN U10276 ( .A(n10027), .B(n42173), .Z(n9988) );
  NANDN U10277 ( .A(n9986), .B(n42172), .Z(n9987) );
  NAND U10278 ( .A(n9988), .B(n9987), .Z(n10036) );
  NAND U10279 ( .A(b[7]), .B(a[234]), .Z(n10037) );
  XNOR U10280 ( .A(n10036), .B(n10037), .Z(n10039) );
  XOR U10281 ( .A(n10038), .B(n10039), .Z(n10045) );
  NANDN U10282 ( .A(n9989), .B(n42093), .Z(n9991) );
  XOR U10283 ( .A(n42134), .B(a[240]), .Z(n10030) );
  NANDN U10284 ( .A(n10030), .B(n42095), .Z(n9990) );
  NAND U10285 ( .A(n9991), .B(n9990), .Z(n10043) );
  NANDN U10286 ( .A(n9992), .B(n42231), .Z(n9994) );
  XOR U10287 ( .A(n181), .B(a[236]), .Z(n10033) );
  NANDN U10288 ( .A(n10033), .B(n42234), .Z(n9993) );
  AND U10289 ( .A(n9994), .B(n9993), .Z(n10042) );
  XNOR U10290 ( .A(n10043), .B(n10042), .Z(n10044) );
  XNOR U10291 ( .A(n10045), .B(n10044), .Z(n10049) );
  NANDN U10292 ( .A(n9996), .B(n9995), .Z(n10000) );
  NAND U10293 ( .A(n9998), .B(n9997), .Z(n9999) );
  AND U10294 ( .A(n10000), .B(n9999), .Z(n10048) );
  XOR U10295 ( .A(n10049), .B(n10048), .Z(n10050) );
  NANDN U10296 ( .A(n10002), .B(n10001), .Z(n10006) );
  NANDN U10297 ( .A(n10004), .B(n10003), .Z(n10005) );
  NAND U10298 ( .A(n10006), .B(n10005), .Z(n10051) );
  XOR U10299 ( .A(n10050), .B(n10051), .Z(n10018) );
  OR U10300 ( .A(n10008), .B(n10007), .Z(n10012) );
  NANDN U10301 ( .A(n10010), .B(n10009), .Z(n10011) );
  NAND U10302 ( .A(n10012), .B(n10011), .Z(n10019) );
  XNOR U10303 ( .A(n10018), .B(n10019), .Z(n10020) );
  XNOR U10304 ( .A(n10021), .B(n10020), .Z(n10054) );
  XNOR U10305 ( .A(n10054), .B(sreg[1258]), .Z(n10056) );
  NAND U10306 ( .A(n10013), .B(sreg[1257]), .Z(n10017) );
  OR U10307 ( .A(n10015), .B(n10014), .Z(n10016) );
  AND U10308 ( .A(n10017), .B(n10016), .Z(n10055) );
  XOR U10309 ( .A(n10056), .B(n10055), .Z(c[1258]) );
  NANDN U10310 ( .A(n10019), .B(n10018), .Z(n10023) );
  NAND U10311 ( .A(n10021), .B(n10020), .Z(n10022) );
  NAND U10312 ( .A(n10023), .B(n10022), .Z(n10062) );
  NAND U10313 ( .A(b[0]), .B(a[243]), .Z(n10024) );
  XNOR U10314 ( .A(b[1]), .B(n10024), .Z(n10026) );
  NAND U10315 ( .A(n49), .B(a[242]), .Z(n10025) );
  AND U10316 ( .A(n10026), .B(n10025), .Z(n10079) );
  XOR U10317 ( .A(a[239]), .B(n42197), .Z(n10068) );
  NANDN U10318 ( .A(n10068), .B(n42173), .Z(n10029) );
  NANDN U10319 ( .A(n10027), .B(n42172), .Z(n10028) );
  NAND U10320 ( .A(n10029), .B(n10028), .Z(n10077) );
  NAND U10321 ( .A(b[7]), .B(a[235]), .Z(n10078) );
  XNOR U10322 ( .A(n10077), .B(n10078), .Z(n10080) );
  XOR U10323 ( .A(n10079), .B(n10080), .Z(n10086) );
  NANDN U10324 ( .A(n10030), .B(n42093), .Z(n10032) );
  XOR U10325 ( .A(n42134), .B(a[241]), .Z(n10071) );
  NANDN U10326 ( .A(n10071), .B(n42095), .Z(n10031) );
  NAND U10327 ( .A(n10032), .B(n10031), .Z(n10084) );
  NANDN U10328 ( .A(n10033), .B(n42231), .Z(n10035) );
  XOR U10329 ( .A(n181), .B(a[237]), .Z(n10074) );
  NANDN U10330 ( .A(n10074), .B(n42234), .Z(n10034) );
  AND U10331 ( .A(n10035), .B(n10034), .Z(n10083) );
  XNOR U10332 ( .A(n10084), .B(n10083), .Z(n10085) );
  XNOR U10333 ( .A(n10086), .B(n10085), .Z(n10090) );
  NANDN U10334 ( .A(n10037), .B(n10036), .Z(n10041) );
  NAND U10335 ( .A(n10039), .B(n10038), .Z(n10040) );
  AND U10336 ( .A(n10041), .B(n10040), .Z(n10089) );
  XOR U10337 ( .A(n10090), .B(n10089), .Z(n10091) );
  NANDN U10338 ( .A(n10043), .B(n10042), .Z(n10047) );
  NANDN U10339 ( .A(n10045), .B(n10044), .Z(n10046) );
  NAND U10340 ( .A(n10047), .B(n10046), .Z(n10092) );
  XOR U10341 ( .A(n10091), .B(n10092), .Z(n10059) );
  OR U10342 ( .A(n10049), .B(n10048), .Z(n10053) );
  NANDN U10343 ( .A(n10051), .B(n10050), .Z(n10052) );
  NAND U10344 ( .A(n10053), .B(n10052), .Z(n10060) );
  XNOR U10345 ( .A(n10059), .B(n10060), .Z(n10061) );
  XNOR U10346 ( .A(n10062), .B(n10061), .Z(n10095) );
  XNOR U10347 ( .A(n10095), .B(sreg[1259]), .Z(n10097) );
  NAND U10348 ( .A(n10054), .B(sreg[1258]), .Z(n10058) );
  OR U10349 ( .A(n10056), .B(n10055), .Z(n10057) );
  AND U10350 ( .A(n10058), .B(n10057), .Z(n10096) );
  XOR U10351 ( .A(n10097), .B(n10096), .Z(c[1259]) );
  NANDN U10352 ( .A(n10060), .B(n10059), .Z(n10064) );
  NAND U10353 ( .A(n10062), .B(n10061), .Z(n10063) );
  NAND U10354 ( .A(n10064), .B(n10063), .Z(n10103) );
  NAND U10355 ( .A(b[0]), .B(a[244]), .Z(n10065) );
  XNOR U10356 ( .A(b[1]), .B(n10065), .Z(n10067) );
  NAND U10357 ( .A(n49), .B(a[243]), .Z(n10066) );
  AND U10358 ( .A(n10067), .B(n10066), .Z(n10120) );
  XOR U10359 ( .A(a[240]), .B(n42197), .Z(n10109) );
  NANDN U10360 ( .A(n10109), .B(n42173), .Z(n10070) );
  NANDN U10361 ( .A(n10068), .B(n42172), .Z(n10069) );
  NAND U10362 ( .A(n10070), .B(n10069), .Z(n10118) );
  NAND U10363 ( .A(b[7]), .B(a[236]), .Z(n10119) );
  XNOR U10364 ( .A(n10118), .B(n10119), .Z(n10121) );
  XOR U10365 ( .A(n10120), .B(n10121), .Z(n10127) );
  NANDN U10366 ( .A(n10071), .B(n42093), .Z(n10073) );
  XOR U10367 ( .A(n42134), .B(a[242]), .Z(n10112) );
  NANDN U10368 ( .A(n10112), .B(n42095), .Z(n10072) );
  NAND U10369 ( .A(n10073), .B(n10072), .Z(n10125) );
  NANDN U10370 ( .A(n10074), .B(n42231), .Z(n10076) );
  XOR U10371 ( .A(n181), .B(a[238]), .Z(n10115) );
  NANDN U10372 ( .A(n10115), .B(n42234), .Z(n10075) );
  AND U10373 ( .A(n10076), .B(n10075), .Z(n10124) );
  XNOR U10374 ( .A(n10125), .B(n10124), .Z(n10126) );
  XNOR U10375 ( .A(n10127), .B(n10126), .Z(n10131) );
  NANDN U10376 ( .A(n10078), .B(n10077), .Z(n10082) );
  NAND U10377 ( .A(n10080), .B(n10079), .Z(n10081) );
  AND U10378 ( .A(n10082), .B(n10081), .Z(n10130) );
  XOR U10379 ( .A(n10131), .B(n10130), .Z(n10132) );
  NANDN U10380 ( .A(n10084), .B(n10083), .Z(n10088) );
  NANDN U10381 ( .A(n10086), .B(n10085), .Z(n10087) );
  NAND U10382 ( .A(n10088), .B(n10087), .Z(n10133) );
  XOR U10383 ( .A(n10132), .B(n10133), .Z(n10100) );
  OR U10384 ( .A(n10090), .B(n10089), .Z(n10094) );
  NANDN U10385 ( .A(n10092), .B(n10091), .Z(n10093) );
  NAND U10386 ( .A(n10094), .B(n10093), .Z(n10101) );
  XNOR U10387 ( .A(n10100), .B(n10101), .Z(n10102) );
  XNOR U10388 ( .A(n10103), .B(n10102), .Z(n10136) );
  XNOR U10389 ( .A(n10136), .B(sreg[1260]), .Z(n10138) );
  NAND U10390 ( .A(n10095), .B(sreg[1259]), .Z(n10099) );
  OR U10391 ( .A(n10097), .B(n10096), .Z(n10098) );
  AND U10392 ( .A(n10099), .B(n10098), .Z(n10137) );
  XOR U10393 ( .A(n10138), .B(n10137), .Z(c[1260]) );
  NANDN U10394 ( .A(n10101), .B(n10100), .Z(n10105) );
  NAND U10395 ( .A(n10103), .B(n10102), .Z(n10104) );
  NAND U10396 ( .A(n10105), .B(n10104), .Z(n10144) );
  NAND U10397 ( .A(b[0]), .B(a[245]), .Z(n10106) );
  XNOR U10398 ( .A(b[1]), .B(n10106), .Z(n10108) );
  NAND U10399 ( .A(n50), .B(a[244]), .Z(n10107) );
  AND U10400 ( .A(n10108), .B(n10107), .Z(n10161) );
  XOR U10401 ( .A(a[241]), .B(n42197), .Z(n10150) );
  NANDN U10402 ( .A(n10150), .B(n42173), .Z(n10111) );
  NANDN U10403 ( .A(n10109), .B(n42172), .Z(n10110) );
  NAND U10404 ( .A(n10111), .B(n10110), .Z(n10159) );
  NAND U10405 ( .A(b[7]), .B(a[237]), .Z(n10160) );
  XNOR U10406 ( .A(n10159), .B(n10160), .Z(n10162) );
  XOR U10407 ( .A(n10161), .B(n10162), .Z(n10168) );
  NANDN U10408 ( .A(n10112), .B(n42093), .Z(n10114) );
  XOR U10409 ( .A(n42134), .B(a[243]), .Z(n10153) );
  NANDN U10410 ( .A(n10153), .B(n42095), .Z(n10113) );
  NAND U10411 ( .A(n10114), .B(n10113), .Z(n10166) );
  NANDN U10412 ( .A(n10115), .B(n42231), .Z(n10117) );
  XOR U10413 ( .A(n182), .B(a[239]), .Z(n10156) );
  NANDN U10414 ( .A(n10156), .B(n42234), .Z(n10116) );
  AND U10415 ( .A(n10117), .B(n10116), .Z(n10165) );
  XNOR U10416 ( .A(n10166), .B(n10165), .Z(n10167) );
  XNOR U10417 ( .A(n10168), .B(n10167), .Z(n10172) );
  NANDN U10418 ( .A(n10119), .B(n10118), .Z(n10123) );
  NAND U10419 ( .A(n10121), .B(n10120), .Z(n10122) );
  AND U10420 ( .A(n10123), .B(n10122), .Z(n10171) );
  XOR U10421 ( .A(n10172), .B(n10171), .Z(n10173) );
  NANDN U10422 ( .A(n10125), .B(n10124), .Z(n10129) );
  NANDN U10423 ( .A(n10127), .B(n10126), .Z(n10128) );
  NAND U10424 ( .A(n10129), .B(n10128), .Z(n10174) );
  XOR U10425 ( .A(n10173), .B(n10174), .Z(n10141) );
  OR U10426 ( .A(n10131), .B(n10130), .Z(n10135) );
  NANDN U10427 ( .A(n10133), .B(n10132), .Z(n10134) );
  NAND U10428 ( .A(n10135), .B(n10134), .Z(n10142) );
  XNOR U10429 ( .A(n10141), .B(n10142), .Z(n10143) );
  XNOR U10430 ( .A(n10144), .B(n10143), .Z(n10177) );
  XNOR U10431 ( .A(n10177), .B(sreg[1261]), .Z(n10179) );
  NAND U10432 ( .A(n10136), .B(sreg[1260]), .Z(n10140) );
  OR U10433 ( .A(n10138), .B(n10137), .Z(n10139) );
  AND U10434 ( .A(n10140), .B(n10139), .Z(n10178) );
  XOR U10435 ( .A(n10179), .B(n10178), .Z(c[1261]) );
  NANDN U10436 ( .A(n10142), .B(n10141), .Z(n10146) );
  NAND U10437 ( .A(n10144), .B(n10143), .Z(n10145) );
  NAND U10438 ( .A(n10146), .B(n10145), .Z(n10185) );
  NAND U10439 ( .A(b[0]), .B(a[246]), .Z(n10147) );
  XNOR U10440 ( .A(b[1]), .B(n10147), .Z(n10149) );
  NAND U10441 ( .A(n50), .B(a[245]), .Z(n10148) );
  AND U10442 ( .A(n10149), .B(n10148), .Z(n10202) );
  XOR U10443 ( .A(a[242]), .B(n42197), .Z(n10191) );
  NANDN U10444 ( .A(n10191), .B(n42173), .Z(n10152) );
  NANDN U10445 ( .A(n10150), .B(n42172), .Z(n10151) );
  NAND U10446 ( .A(n10152), .B(n10151), .Z(n10200) );
  NAND U10447 ( .A(b[7]), .B(a[238]), .Z(n10201) );
  XNOR U10448 ( .A(n10200), .B(n10201), .Z(n10203) );
  XOR U10449 ( .A(n10202), .B(n10203), .Z(n10209) );
  NANDN U10450 ( .A(n10153), .B(n42093), .Z(n10155) );
  XOR U10451 ( .A(n42134), .B(a[244]), .Z(n10194) );
  NANDN U10452 ( .A(n10194), .B(n42095), .Z(n10154) );
  NAND U10453 ( .A(n10155), .B(n10154), .Z(n10207) );
  NANDN U10454 ( .A(n10156), .B(n42231), .Z(n10158) );
  XOR U10455 ( .A(n182), .B(a[240]), .Z(n10197) );
  NANDN U10456 ( .A(n10197), .B(n42234), .Z(n10157) );
  AND U10457 ( .A(n10158), .B(n10157), .Z(n10206) );
  XNOR U10458 ( .A(n10207), .B(n10206), .Z(n10208) );
  XNOR U10459 ( .A(n10209), .B(n10208), .Z(n10213) );
  NANDN U10460 ( .A(n10160), .B(n10159), .Z(n10164) );
  NAND U10461 ( .A(n10162), .B(n10161), .Z(n10163) );
  AND U10462 ( .A(n10164), .B(n10163), .Z(n10212) );
  XOR U10463 ( .A(n10213), .B(n10212), .Z(n10214) );
  NANDN U10464 ( .A(n10166), .B(n10165), .Z(n10170) );
  NANDN U10465 ( .A(n10168), .B(n10167), .Z(n10169) );
  NAND U10466 ( .A(n10170), .B(n10169), .Z(n10215) );
  XOR U10467 ( .A(n10214), .B(n10215), .Z(n10182) );
  OR U10468 ( .A(n10172), .B(n10171), .Z(n10176) );
  NANDN U10469 ( .A(n10174), .B(n10173), .Z(n10175) );
  NAND U10470 ( .A(n10176), .B(n10175), .Z(n10183) );
  XNOR U10471 ( .A(n10182), .B(n10183), .Z(n10184) );
  XNOR U10472 ( .A(n10185), .B(n10184), .Z(n10218) );
  XNOR U10473 ( .A(n10218), .B(sreg[1262]), .Z(n10220) );
  NAND U10474 ( .A(n10177), .B(sreg[1261]), .Z(n10181) );
  OR U10475 ( .A(n10179), .B(n10178), .Z(n10180) );
  AND U10476 ( .A(n10181), .B(n10180), .Z(n10219) );
  XOR U10477 ( .A(n10220), .B(n10219), .Z(c[1262]) );
  NANDN U10478 ( .A(n10183), .B(n10182), .Z(n10187) );
  NAND U10479 ( .A(n10185), .B(n10184), .Z(n10186) );
  NAND U10480 ( .A(n10187), .B(n10186), .Z(n10226) );
  NAND U10481 ( .A(b[0]), .B(a[247]), .Z(n10188) );
  XNOR U10482 ( .A(b[1]), .B(n10188), .Z(n10190) );
  NAND U10483 ( .A(n50), .B(a[246]), .Z(n10189) );
  AND U10484 ( .A(n10190), .B(n10189), .Z(n10243) );
  XOR U10485 ( .A(a[243]), .B(n42197), .Z(n10232) );
  NANDN U10486 ( .A(n10232), .B(n42173), .Z(n10193) );
  NANDN U10487 ( .A(n10191), .B(n42172), .Z(n10192) );
  NAND U10488 ( .A(n10193), .B(n10192), .Z(n10241) );
  NAND U10489 ( .A(b[7]), .B(a[239]), .Z(n10242) );
  XNOR U10490 ( .A(n10241), .B(n10242), .Z(n10244) );
  XOR U10491 ( .A(n10243), .B(n10244), .Z(n10250) );
  NANDN U10492 ( .A(n10194), .B(n42093), .Z(n10196) );
  XOR U10493 ( .A(n42134), .B(a[245]), .Z(n10235) );
  NANDN U10494 ( .A(n10235), .B(n42095), .Z(n10195) );
  NAND U10495 ( .A(n10196), .B(n10195), .Z(n10248) );
  NANDN U10496 ( .A(n10197), .B(n42231), .Z(n10199) );
  XOR U10497 ( .A(n182), .B(a[241]), .Z(n10238) );
  NANDN U10498 ( .A(n10238), .B(n42234), .Z(n10198) );
  AND U10499 ( .A(n10199), .B(n10198), .Z(n10247) );
  XNOR U10500 ( .A(n10248), .B(n10247), .Z(n10249) );
  XNOR U10501 ( .A(n10250), .B(n10249), .Z(n10254) );
  NANDN U10502 ( .A(n10201), .B(n10200), .Z(n10205) );
  NAND U10503 ( .A(n10203), .B(n10202), .Z(n10204) );
  AND U10504 ( .A(n10205), .B(n10204), .Z(n10253) );
  XOR U10505 ( .A(n10254), .B(n10253), .Z(n10255) );
  NANDN U10506 ( .A(n10207), .B(n10206), .Z(n10211) );
  NANDN U10507 ( .A(n10209), .B(n10208), .Z(n10210) );
  NAND U10508 ( .A(n10211), .B(n10210), .Z(n10256) );
  XOR U10509 ( .A(n10255), .B(n10256), .Z(n10223) );
  OR U10510 ( .A(n10213), .B(n10212), .Z(n10217) );
  NANDN U10511 ( .A(n10215), .B(n10214), .Z(n10216) );
  NAND U10512 ( .A(n10217), .B(n10216), .Z(n10224) );
  XNOR U10513 ( .A(n10223), .B(n10224), .Z(n10225) );
  XNOR U10514 ( .A(n10226), .B(n10225), .Z(n10259) );
  XNOR U10515 ( .A(n10259), .B(sreg[1263]), .Z(n10261) );
  NAND U10516 ( .A(n10218), .B(sreg[1262]), .Z(n10222) );
  OR U10517 ( .A(n10220), .B(n10219), .Z(n10221) );
  AND U10518 ( .A(n10222), .B(n10221), .Z(n10260) );
  XOR U10519 ( .A(n10261), .B(n10260), .Z(c[1263]) );
  NANDN U10520 ( .A(n10224), .B(n10223), .Z(n10228) );
  NAND U10521 ( .A(n10226), .B(n10225), .Z(n10227) );
  NAND U10522 ( .A(n10228), .B(n10227), .Z(n10267) );
  NAND U10523 ( .A(b[0]), .B(a[248]), .Z(n10229) );
  XNOR U10524 ( .A(b[1]), .B(n10229), .Z(n10231) );
  NAND U10525 ( .A(n50), .B(a[247]), .Z(n10230) );
  AND U10526 ( .A(n10231), .B(n10230), .Z(n10284) );
  XOR U10527 ( .A(a[244]), .B(n42197), .Z(n10273) );
  NANDN U10528 ( .A(n10273), .B(n42173), .Z(n10234) );
  NANDN U10529 ( .A(n10232), .B(n42172), .Z(n10233) );
  NAND U10530 ( .A(n10234), .B(n10233), .Z(n10282) );
  NAND U10531 ( .A(b[7]), .B(a[240]), .Z(n10283) );
  XNOR U10532 ( .A(n10282), .B(n10283), .Z(n10285) );
  XOR U10533 ( .A(n10284), .B(n10285), .Z(n10291) );
  NANDN U10534 ( .A(n10235), .B(n42093), .Z(n10237) );
  XOR U10535 ( .A(n42134), .B(a[246]), .Z(n10276) );
  NANDN U10536 ( .A(n10276), .B(n42095), .Z(n10236) );
  NAND U10537 ( .A(n10237), .B(n10236), .Z(n10289) );
  NANDN U10538 ( .A(n10238), .B(n42231), .Z(n10240) );
  XOR U10539 ( .A(n182), .B(a[242]), .Z(n10279) );
  NANDN U10540 ( .A(n10279), .B(n42234), .Z(n10239) );
  AND U10541 ( .A(n10240), .B(n10239), .Z(n10288) );
  XNOR U10542 ( .A(n10289), .B(n10288), .Z(n10290) );
  XNOR U10543 ( .A(n10291), .B(n10290), .Z(n10295) );
  NANDN U10544 ( .A(n10242), .B(n10241), .Z(n10246) );
  NAND U10545 ( .A(n10244), .B(n10243), .Z(n10245) );
  AND U10546 ( .A(n10246), .B(n10245), .Z(n10294) );
  XOR U10547 ( .A(n10295), .B(n10294), .Z(n10296) );
  NANDN U10548 ( .A(n10248), .B(n10247), .Z(n10252) );
  NANDN U10549 ( .A(n10250), .B(n10249), .Z(n10251) );
  NAND U10550 ( .A(n10252), .B(n10251), .Z(n10297) );
  XOR U10551 ( .A(n10296), .B(n10297), .Z(n10264) );
  OR U10552 ( .A(n10254), .B(n10253), .Z(n10258) );
  NANDN U10553 ( .A(n10256), .B(n10255), .Z(n10257) );
  NAND U10554 ( .A(n10258), .B(n10257), .Z(n10265) );
  XNOR U10555 ( .A(n10264), .B(n10265), .Z(n10266) );
  XNOR U10556 ( .A(n10267), .B(n10266), .Z(n10300) );
  XNOR U10557 ( .A(n10300), .B(sreg[1264]), .Z(n10302) );
  NAND U10558 ( .A(n10259), .B(sreg[1263]), .Z(n10263) );
  OR U10559 ( .A(n10261), .B(n10260), .Z(n10262) );
  AND U10560 ( .A(n10263), .B(n10262), .Z(n10301) );
  XOR U10561 ( .A(n10302), .B(n10301), .Z(c[1264]) );
  NANDN U10562 ( .A(n10265), .B(n10264), .Z(n10269) );
  NAND U10563 ( .A(n10267), .B(n10266), .Z(n10268) );
  NAND U10564 ( .A(n10269), .B(n10268), .Z(n10308) );
  NAND U10565 ( .A(b[0]), .B(a[249]), .Z(n10270) );
  XNOR U10566 ( .A(b[1]), .B(n10270), .Z(n10272) );
  NAND U10567 ( .A(n50), .B(a[248]), .Z(n10271) );
  AND U10568 ( .A(n10272), .B(n10271), .Z(n10325) );
  XOR U10569 ( .A(a[245]), .B(n42197), .Z(n10314) );
  NANDN U10570 ( .A(n10314), .B(n42173), .Z(n10275) );
  NANDN U10571 ( .A(n10273), .B(n42172), .Z(n10274) );
  NAND U10572 ( .A(n10275), .B(n10274), .Z(n10323) );
  NAND U10573 ( .A(b[7]), .B(a[241]), .Z(n10324) );
  XNOR U10574 ( .A(n10323), .B(n10324), .Z(n10326) );
  XOR U10575 ( .A(n10325), .B(n10326), .Z(n10332) );
  NANDN U10576 ( .A(n10276), .B(n42093), .Z(n10278) );
  XOR U10577 ( .A(n42134), .B(a[247]), .Z(n10317) );
  NANDN U10578 ( .A(n10317), .B(n42095), .Z(n10277) );
  NAND U10579 ( .A(n10278), .B(n10277), .Z(n10330) );
  NANDN U10580 ( .A(n10279), .B(n42231), .Z(n10281) );
  XOR U10581 ( .A(n182), .B(a[243]), .Z(n10320) );
  NANDN U10582 ( .A(n10320), .B(n42234), .Z(n10280) );
  AND U10583 ( .A(n10281), .B(n10280), .Z(n10329) );
  XNOR U10584 ( .A(n10330), .B(n10329), .Z(n10331) );
  XNOR U10585 ( .A(n10332), .B(n10331), .Z(n10336) );
  NANDN U10586 ( .A(n10283), .B(n10282), .Z(n10287) );
  NAND U10587 ( .A(n10285), .B(n10284), .Z(n10286) );
  AND U10588 ( .A(n10287), .B(n10286), .Z(n10335) );
  XOR U10589 ( .A(n10336), .B(n10335), .Z(n10337) );
  NANDN U10590 ( .A(n10289), .B(n10288), .Z(n10293) );
  NANDN U10591 ( .A(n10291), .B(n10290), .Z(n10292) );
  NAND U10592 ( .A(n10293), .B(n10292), .Z(n10338) );
  XOR U10593 ( .A(n10337), .B(n10338), .Z(n10305) );
  OR U10594 ( .A(n10295), .B(n10294), .Z(n10299) );
  NANDN U10595 ( .A(n10297), .B(n10296), .Z(n10298) );
  NAND U10596 ( .A(n10299), .B(n10298), .Z(n10306) );
  XNOR U10597 ( .A(n10305), .B(n10306), .Z(n10307) );
  XNOR U10598 ( .A(n10308), .B(n10307), .Z(n10341) );
  XNOR U10599 ( .A(n10341), .B(sreg[1265]), .Z(n10343) );
  NAND U10600 ( .A(n10300), .B(sreg[1264]), .Z(n10304) );
  OR U10601 ( .A(n10302), .B(n10301), .Z(n10303) );
  AND U10602 ( .A(n10304), .B(n10303), .Z(n10342) );
  XOR U10603 ( .A(n10343), .B(n10342), .Z(c[1265]) );
  NANDN U10604 ( .A(n10306), .B(n10305), .Z(n10310) );
  NAND U10605 ( .A(n10308), .B(n10307), .Z(n10309) );
  NAND U10606 ( .A(n10310), .B(n10309), .Z(n10349) );
  NAND U10607 ( .A(b[0]), .B(a[250]), .Z(n10311) );
  XNOR U10608 ( .A(b[1]), .B(n10311), .Z(n10313) );
  NAND U10609 ( .A(n50), .B(a[249]), .Z(n10312) );
  AND U10610 ( .A(n10313), .B(n10312), .Z(n10366) );
  XOR U10611 ( .A(a[246]), .B(n42197), .Z(n10355) );
  NANDN U10612 ( .A(n10355), .B(n42173), .Z(n10316) );
  NANDN U10613 ( .A(n10314), .B(n42172), .Z(n10315) );
  NAND U10614 ( .A(n10316), .B(n10315), .Z(n10364) );
  NAND U10615 ( .A(b[7]), .B(a[242]), .Z(n10365) );
  XNOR U10616 ( .A(n10364), .B(n10365), .Z(n10367) );
  XOR U10617 ( .A(n10366), .B(n10367), .Z(n10373) );
  NANDN U10618 ( .A(n10317), .B(n42093), .Z(n10319) );
  XOR U10619 ( .A(n42134), .B(a[248]), .Z(n10358) );
  NANDN U10620 ( .A(n10358), .B(n42095), .Z(n10318) );
  NAND U10621 ( .A(n10319), .B(n10318), .Z(n10371) );
  NANDN U10622 ( .A(n10320), .B(n42231), .Z(n10322) );
  XOR U10623 ( .A(n182), .B(a[244]), .Z(n10361) );
  NANDN U10624 ( .A(n10361), .B(n42234), .Z(n10321) );
  AND U10625 ( .A(n10322), .B(n10321), .Z(n10370) );
  XNOR U10626 ( .A(n10371), .B(n10370), .Z(n10372) );
  XNOR U10627 ( .A(n10373), .B(n10372), .Z(n10377) );
  NANDN U10628 ( .A(n10324), .B(n10323), .Z(n10328) );
  NAND U10629 ( .A(n10326), .B(n10325), .Z(n10327) );
  AND U10630 ( .A(n10328), .B(n10327), .Z(n10376) );
  XOR U10631 ( .A(n10377), .B(n10376), .Z(n10378) );
  NANDN U10632 ( .A(n10330), .B(n10329), .Z(n10334) );
  NANDN U10633 ( .A(n10332), .B(n10331), .Z(n10333) );
  NAND U10634 ( .A(n10334), .B(n10333), .Z(n10379) );
  XOR U10635 ( .A(n10378), .B(n10379), .Z(n10346) );
  OR U10636 ( .A(n10336), .B(n10335), .Z(n10340) );
  NANDN U10637 ( .A(n10338), .B(n10337), .Z(n10339) );
  NAND U10638 ( .A(n10340), .B(n10339), .Z(n10347) );
  XNOR U10639 ( .A(n10346), .B(n10347), .Z(n10348) );
  XNOR U10640 ( .A(n10349), .B(n10348), .Z(n10382) );
  XNOR U10641 ( .A(n10382), .B(sreg[1266]), .Z(n10384) );
  NAND U10642 ( .A(n10341), .B(sreg[1265]), .Z(n10345) );
  OR U10643 ( .A(n10343), .B(n10342), .Z(n10344) );
  AND U10644 ( .A(n10345), .B(n10344), .Z(n10383) );
  XOR U10645 ( .A(n10384), .B(n10383), .Z(c[1266]) );
  NANDN U10646 ( .A(n10347), .B(n10346), .Z(n10351) );
  NAND U10647 ( .A(n10349), .B(n10348), .Z(n10350) );
  NAND U10648 ( .A(n10351), .B(n10350), .Z(n10390) );
  NAND U10649 ( .A(b[0]), .B(a[251]), .Z(n10352) );
  XNOR U10650 ( .A(b[1]), .B(n10352), .Z(n10354) );
  NAND U10651 ( .A(n50), .B(a[250]), .Z(n10353) );
  AND U10652 ( .A(n10354), .B(n10353), .Z(n10407) );
  XOR U10653 ( .A(a[247]), .B(n42197), .Z(n10396) );
  NANDN U10654 ( .A(n10396), .B(n42173), .Z(n10357) );
  NANDN U10655 ( .A(n10355), .B(n42172), .Z(n10356) );
  NAND U10656 ( .A(n10357), .B(n10356), .Z(n10405) );
  NAND U10657 ( .A(b[7]), .B(a[243]), .Z(n10406) );
  XNOR U10658 ( .A(n10405), .B(n10406), .Z(n10408) );
  XOR U10659 ( .A(n10407), .B(n10408), .Z(n10414) );
  NANDN U10660 ( .A(n10358), .B(n42093), .Z(n10360) );
  XOR U10661 ( .A(n42134), .B(a[249]), .Z(n10399) );
  NANDN U10662 ( .A(n10399), .B(n42095), .Z(n10359) );
  NAND U10663 ( .A(n10360), .B(n10359), .Z(n10412) );
  NANDN U10664 ( .A(n10361), .B(n42231), .Z(n10363) );
  XOR U10665 ( .A(n182), .B(a[245]), .Z(n10402) );
  NANDN U10666 ( .A(n10402), .B(n42234), .Z(n10362) );
  AND U10667 ( .A(n10363), .B(n10362), .Z(n10411) );
  XNOR U10668 ( .A(n10412), .B(n10411), .Z(n10413) );
  XNOR U10669 ( .A(n10414), .B(n10413), .Z(n10418) );
  NANDN U10670 ( .A(n10365), .B(n10364), .Z(n10369) );
  NAND U10671 ( .A(n10367), .B(n10366), .Z(n10368) );
  AND U10672 ( .A(n10369), .B(n10368), .Z(n10417) );
  XOR U10673 ( .A(n10418), .B(n10417), .Z(n10419) );
  NANDN U10674 ( .A(n10371), .B(n10370), .Z(n10375) );
  NANDN U10675 ( .A(n10373), .B(n10372), .Z(n10374) );
  NAND U10676 ( .A(n10375), .B(n10374), .Z(n10420) );
  XOR U10677 ( .A(n10419), .B(n10420), .Z(n10387) );
  OR U10678 ( .A(n10377), .B(n10376), .Z(n10381) );
  NANDN U10679 ( .A(n10379), .B(n10378), .Z(n10380) );
  NAND U10680 ( .A(n10381), .B(n10380), .Z(n10388) );
  XNOR U10681 ( .A(n10387), .B(n10388), .Z(n10389) );
  XNOR U10682 ( .A(n10390), .B(n10389), .Z(n10423) );
  XNOR U10683 ( .A(n10423), .B(sreg[1267]), .Z(n10425) );
  NAND U10684 ( .A(n10382), .B(sreg[1266]), .Z(n10386) );
  OR U10685 ( .A(n10384), .B(n10383), .Z(n10385) );
  AND U10686 ( .A(n10386), .B(n10385), .Z(n10424) );
  XOR U10687 ( .A(n10425), .B(n10424), .Z(c[1267]) );
  NANDN U10688 ( .A(n10388), .B(n10387), .Z(n10392) );
  NAND U10689 ( .A(n10390), .B(n10389), .Z(n10391) );
  NAND U10690 ( .A(n10392), .B(n10391), .Z(n10431) );
  NAND U10691 ( .A(b[0]), .B(a[252]), .Z(n10393) );
  XNOR U10692 ( .A(b[1]), .B(n10393), .Z(n10395) );
  NAND U10693 ( .A(n51), .B(a[251]), .Z(n10394) );
  AND U10694 ( .A(n10395), .B(n10394), .Z(n10448) );
  XOR U10695 ( .A(a[248]), .B(n42197), .Z(n10437) );
  NANDN U10696 ( .A(n10437), .B(n42173), .Z(n10398) );
  NANDN U10697 ( .A(n10396), .B(n42172), .Z(n10397) );
  NAND U10698 ( .A(n10398), .B(n10397), .Z(n10446) );
  NAND U10699 ( .A(b[7]), .B(a[244]), .Z(n10447) );
  XNOR U10700 ( .A(n10446), .B(n10447), .Z(n10449) );
  XOR U10701 ( .A(n10448), .B(n10449), .Z(n10455) );
  NANDN U10702 ( .A(n10399), .B(n42093), .Z(n10401) );
  XOR U10703 ( .A(n42134), .B(a[250]), .Z(n10440) );
  NANDN U10704 ( .A(n10440), .B(n42095), .Z(n10400) );
  NAND U10705 ( .A(n10401), .B(n10400), .Z(n10453) );
  NANDN U10706 ( .A(n10402), .B(n42231), .Z(n10404) );
  XOR U10707 ( .A(n182), .B(a[246]), .Z(n10443) );
  NANDN U10708 ( .A(n10443), .B(n42234), .Z(n10403) );
  AND U10709 ( .A(n10404), .B(n10403), .Z(n10452) );
  XNOR U10710 ( .A(n10453), .B(n10452), .Z(n10454) );
  XNOR U10711 ( .A(n10455), .B(n10454), .Z(n10459) );
  NANDN U10712 ( .A(n10406), .B(n10405), .Z(n10410) );
  NAND U10713 ( .A(n10408), .B(n10407), .Z(n10409) );
  AND U10714 ( .A(n10410), .B(n10409), .Z(n10458) );
  XOR U10715 ( .A(n10459), .B(n10458), .Z(n10460) );
  NANDN U10716 ( .A(n10412), .B(n10411), .Z(n10416) );
  NANDN U10717 ( .A(n10414), .B(n10413), .Z(n10415) );
  NAND U10718 ( .A(n10416), .B(n10415), .Z(n10461) );
  XOR U10719 ( .A(n10460), .B(n10461), .Z(n10428) );
  OR U10720 ( .A(n10418), .B(n10417), .Z(n10422) );
  NANDN U10721 ( .A(n10420), .B(n10419), .Z(n10421) );
  NAND U10722 ( .A(n10422), .B(n10421), .Z(n10429) );
  XNOR U10723 ( .A(n10428), .B(n10429), .Z(n10430) );
  XNOR U10724 ( .A(n10431), .B(n10430), .Z(n10464) );
  XNOR U10725 ( .A(n10464), .B(sreg[1268]), .Z(n10466) );
  NAND U10726 ( .A(n10423), .B(sreg[1267]), .Z(n10427) );
  OR U10727 ( .A(n10425), .B(n10424), .Z(n10426) );
  AND U10728 ( .A(n10427), .B(n10426), .Z(n10465) );
  XOR U10729 ( .A(n10466), .B(n10465), .Z(c[1268]) );
  NANDN U10730 ( .A(n10429), .B(n10428), .Z(n10433) );
  NAND U10731 ( .A(n10431), .B(n10430), .Z(n10432) );
  NAND U10732 ( .A(n10433), .B(n10432), .Z(n10472) );
  NAND U10733 ( .A(b[0]), .B(a[253]), .Z(n10434) );
  XNOR U10734 ( .A(b[1]), .B(n10434), .Z(n10436) );
  NAND U10735 ( .A(n51), .B(a[252]), .Z(n10435) );
  AND U10736 ( .A(n10436), .B(n10435), .Z(n10489) );
  XOR U10737 ( .A(a[249]), .B(n42197), .Z(n10478) );
  NANDN U10738 ( .A(n10478), .B(n42173), .Z(n10439) );
  NANDN U10739 ( .A(n10437), .B(n42172), .Z(n10438) );
  NAND U10740 ( .A(n10439), .B(n10438), .Z(n10487) );
  NAND U10741 ( .A(b[7]), .B(a[245]), .Z(n10488) );
  XNOR U10742 ( .A(n10487), .B(n10488), .Z(n10490) );
  XOR U10743 ( .A(n10489), .B(n10490), .Z(n10496) );
  NANDN U10744 ( .A(n10440), .B(n42093), .Z(n10442) );
  XOR U10745 ( .A(n42134), .B(a[251]), .Z(n10481) );
  NANDN U10746 ( .A(n10481), .B(n42095), .Z(n10441) );
  NAND U10747 ( .A(n10442), .B(n10441), .Z(n10494) );
  NANDN U10748 ( .A(n10443), .B(n42231), .Z(n10445) );
  XOR U10749 ( .A(n182), .B(a[247]), .Z(n10484) );
  NANDN U10750 ( .A(n10484), .B(n42234), .Z(n10444) );
  AND U10751 ( .A(n10445), .B(n10444), .Z(n10493) );
  XNOR U10752 ( .A(n10494), .B(n10493), .Z(n10495) );
  XNOR U10753 ( .A(n10496), .B(n10495), .Z(n10500) );
  NANDN U10754 ( .A(n10447), .B(n10446), .Z(n10451) );
  NAND U10755 ( .A(n10449), .B(n10448), .Z(n10450) );
  AND U10756 ( .A(n10451), .B(n10450), .Z(n10499) );
  XOR U10757 ( .A(n10500), .B(n10499), .Z(n10501) );
  NANDN U10758 ( .A(n10453), .B(n10452), .Z(n10457) );
  NANDN U10759 ( .A(n10455), .B(n10454), .Z(n10456) );
  NAND U10760 ( .A(n10457), .B(n10456), .Z(n10502) );
  XOR U10761 ( .A(n10501), .B(n10502), .Z(n10469) );
  OR U10762 ( .A(n10459), .B(n10458), .Z(n10463) );
  NANDN U10763 ( .A(n10461), .B(n10460), .Z(n10462) );
  NAND U10764 ( .A(n10463), .B(n10462), .Z(n10470) );
  XNOR U10765 ( .A(n10469), .B(n10470), .Z(n10471) );
  XNOR U10766 ( .A(n10472), .B(n10471), .Z(n10505) );
  XNOR U10767 ( .A(n10505), .B(sreg[1269]), .Z(n10507) );
  NAND U10768 ( .A(n10464), .B(sreg[1268]), .Z(n10468) );
  OR U10769 ( .A(n10466), .B(n10465), .Z(n10467) );
  AND U10770 ( .A(n10468), .B(n10467), .Z(n10506) );
  XOR U10771 ( .A(n10507), .B(n10506), .Z(c[1269]) );
  NANDN U10772 ( .A(n10470), .B(n10469), .Z(n10474) );
  NAND U10773 ( .A(n10472), .B(n10471), .Z(n10473) );
  NAND U10774 ( .A(n10474), .B(n10473), .Z(n10513) );
  NAND U10775 ( .A(b[0]), .B(a[254]), .Z(n10475) );
  XNOR U10776 ( .A(b[1]), .B(n10475), .Z(n10477) );
  NAND U10777 ( .A(n51), .B(a[253]), .Z(n10476) );
  AND U10778 ( .A(n10477), .B(n10476), .Z(n10530) );
  XOR U10779 ( .A(a[250]), .B(n42197), .Z(n10519) );
  NANDN U10780 ( .A(n10519), .B(n42173), .Z(n10480) );
  NANDN U10781 ( .A(n10478), .B(n42172), .Z(n10479) );
  NAND U10782 ( .A(n10480), .B(n10479), .Z(n10528) );
  NAND U10783 ( .A(b[7]), .B(a[246]), .Z(n10529) );
  XNOR U10784 ( .A(n10528), .B(n10529), .Z(n10531) );
  XOR U10785 ( .A(n10530), .B(n10531), .Z(n10537) );
  NANDN U10786 ( .A(n10481), .B(n42093), .Z(n10483) );
  XOR U10787 ( .A(n42134), .B(a[252]), .Z(n10522) );
  NANDN U10788 ( .A(n10522), .B(n42095), .Z(n10482) );
  NAND U10789 ( .A(n10483), .B(n10482), .Z(n10535) );
  NANDN U10790 ( .A(n10484), .B(n42231), .Z(n10486) );
  XOR U10791 ( .A(n182), .B(a[248]), .Z(n10525) );
  NANDN U10792 ( .A(n10525), .B(n42234), .Z(n10485) );
  AND U10793 ( .A(n10486), .B(n10485), .Z(n10534) );
  XNOR U10794 ( .A(n10535), .B(n10534), .Z(n10536) );
  XNOR U10795 ( .A(n10537), .B(n10536), .Z(n10541) );
  NANDN U10796 ( .A(n10488), .B(n10487), .Z(n10492) );
  NAND U10797 ( .A(n10490), .B(n10489), .Z(n10491) );
  AND U10798 ( .A(n10492), .B(n10491), .Z(n10540) );
  XOR U10799 ( .A(n10541), .B(n10540), .Z(n10542) );
  NANDN U10800 ( .A(n10494), .B(n10493), .Z(n10498) );
  NANDN U10801 ( .A(n10496), .B(n10495), .Z(n10497) );
  NAND U10802 ( .A(n10498), .B(n10497), .Z(n10543) );
  XOR U10803 ( .A(n10542), .B(n10543), .Z(n10510) );
  OR U10804 ( .A(n10500), .B(n10499), .Z(n10504) );
  NANDN U10805 ( .A(n10502), .B(n10501), .Z(n10503) );
  NAND U10806 ( .A(n10504), .B(n10503), .Z(n10511) );
  XNOR U10807 ( .A(n10510), .B(n10511), .Z(n10512) );
  XNOR U10808 ( .A(n10513), .B(n10512), .Z(n10546) );
  XNOR U10809 ( .A(n10546), .B(sreg[1270]), .Z(n10548) );
  NAND U10810 ( .A(n10505), .B(sreg[1269]), .Z(n10509) );
  OR U10811 ( .A(n10507), .B(n10506), .Z(n10508) );
  AND U10812 ( .A(n10509), .B(n10508), .Z(n10547) );
  XOR U10813 ( .A(n10548), .B(n10547), .Z(c[1270]) );
  NANDN U10814 ( .A(n10511), .B(n10510), .Z(n10515) );
  NAND U10815 ( .A(n10513), .B(n10512), .Z(n10514) );
  NAND U10816 ( .A(n10515), .B(n10514), .Z(n10554) );
  NAND U10817 ( .A(b[0]), .B(a[255]), .Z(n10516) );
  XNOR U10818 ( .A(b[1]), .B(n10516), .Z(n10518) );
  NAND U10819 ( .A(n51), .B(a[254]), .Z(n10517) );
  AND U10820 ( .A(n10518), .B(n10517), .Z(n10571) );
  XOR U10821 ( .A(a[251]), .B(n42197), .Z(n10560) );
  NANDN U10822 ( .A(n10560), .B(n42173), .Z(n10521) );
  NANDN U10823 ( .A(n10519), .B(n42172), .Z(n10520) );
  NAND U10824 ( .A(n10521), .B(n10520), .Z(n10569) );
  NAND U10825 ( .A(b[7]), .B(a[247]), .Z(n10570) );
  XNOR U10826 ( .A(n10569), .B(n10570), .Z(n10572) );
  XOR U10827 ( .A(n10571), .B(n10572), .Z(n10578) );
  NANDN U10828 ( .A(n10522), .B(n42093), .Z(n10524) );
  XOR U10829 ( .A(n42134), .B(a[253]), .Z(n10563) );
  NANDN U10830 ( .A(n10563), .B(n42095), .Z(n10523) );
  NAND U10831 ( .A(n10524), .B(n10523), .Z(n10576) );
  NANDN U10832 ( .A(n10525), .B(n42231), .Z(n10527) );
  XOR U10833 ( .A(n182), .B(a[249]), .Z(n10566) );
  NANDN U10834 ( .A(n10566), .B(n42234), .Z(n10526) );
  AND U10835 ( .A(n10527), .B(n10526), .Z(n10575) );
  XNOR U10836 ( .A(n10576), .B(n10575), .Z(n10577) );
  XNOR U10837 ( .A(n10578), .B(n10577), .Z(n10582) );
  NANDN U10838 ( .A(n10529), .B(n10528), .Z(n10533) );
  NAND U10839 ( .A(n10531), .B(n10530), .Z(n10532) );
  AND U10840 ( .A(n10533), .B(n10532), .Z(n10581) );
  XOR U10841 ( .A(n10582), .B(n10581), .Z(n10583) );
  NANDN U10842 ( .A(n10535), .B(n10534), .Z(n10539) );
  NANDN U10843 ( .A(n10537), .B(n10536), .Z(n10538) );
  NAND U10844 ( .A(n10539), .B(n10538), .Z(n10584) );
  XOR U10845 ( .A(n10583), .B(n10584), .Z(n10551) );
  OR U10846 ( .A(n10541), .B(n10540), .Z(n10545) );
  NANDN U10847 ( .A(n10543), .B(n10542), .Z(n10544) );
  NAND U10848 ( .A(n10545), .B(n10544), .Z(n10552) );
  XNOR U10849 ( .A(n10551), .B(n10552), .Z(n10553) );
  XNOR U10850 ( .A(n10554), .B(n10553), .Z(n10587) );
  XNOR U10851 ( .A(n10587), .B(sreg[1271]), .Z(n10589) );
  NAND U10852 ( .A(n10546), .B(sreg[1270]), .Z(n10550) );
  OR U10853 ( .A(n10548), .B(n10547), .Z(n10549) );
  AND U10854 ( .A(n10550), .B(n10549), .Z(n10588) );
  XOR U10855 ( .A(n10589), .B(n10588), .Z(c[1271]) );
  NANDN U10856 ( .A(n10552), .B(n10551), .Z(n10556) );
  NAND U10857 ( .A(n10554), .B(n10553), .Z(n10555) );
  NAND U10858 ( .A(n10556), .B(n10555), .Z(n10595) );
  NAND U10859 ( .A(b[0]), .B(a[256]), .Z(n10557) );
  XNOR U10860 ( .A(b[1]), .B(n10557), .Z(n10559) );
  NAND U10861 ( .A(n51), .B(a[255]), .Z(n10558) );
  AND U10862 ( .A(n10559), .B(n10558), .Z(n10612) );
  XOR U10863 ( .A(a[252]), .B(n42197), .Z(n10601) );
  NANDN U10864 ( .A(n10601), .B(n42173), .Z(n10562) );
  NANDN U10865 ( .A(n10560), .B(n42172), .Z(n10561) );
  NAND U10866 ( .A(n10562), .B(n10561), .Z(n10610) );
  NAND U10867 ( .A(b[7]), .B(a[248]), .Z(n10611) );
  XNOR U10868 ( .A(n10610), .B(n10611), .Z(n10613) );
  XOR U10869 ( .A(n10612), .B(n10613), .Z(n10619) );
  NANDN U10870 ( .A(n10563), .B(n42093), .Z(n10565) );
  XOR U10871 ( .A(n42134), .B(a[254]), .Z(n10604) );
  NANDN U10872 ( .A(n10604), .B(n42095), .Z(n10564) );
  NAND U10873 ( .A(n10565), .B(n10564), .Z(n10617) );
  NANDN U10874 ( .A(n10566), .B(n42231), .Z(n10568) );
  XOR U10875 ( .A(n182), .B(a[250]), .Z(n10607) );
  NANDN U10876 ( .A(n10607), .B(n42234), .Z(n10567) );
  AND U10877 ( .A(n10568), .B(n10567), .Z(n10616) );
  XNOR U10878 ( .A(n10617), .B(n10616), .Z(n10618) );
  XNOR U10879 ( .A(n10619), .B(n10618), .Z(n10623) );
  NANDN U10880 ( .A(n10570), .B(n10569), .Z(n10574) );
  NAND U10881 ( .A(n10572), .B(n10571), .Z(n10573) );
  AND U10882 ( .A(n10574), .B(n10573), .Z(n10622) );
  XOR U10883 ( .A(n10623), .B(n10622), .Z(n10624) );
  NANDN U10884 ( .A(n10576), .B(n10575), .Z(n10580) );
  NANDN U10885 ( .A(n10578), .B(n10577), .Z(n10579) );
  NAND U10886 ( .A(n10580), .B(n10579), .Z(n10625) );
  XOR U10887 ( .A(n10624), .B(n10625), .Z(n10592) );
  OR U10888 ( .A(n10582), .B(n10581), .Z(n10586) );
  NANDN U10889 ( .A(n10584), .B(n10583), .Z(n10585) );
  NAND U10890 ( .A(n10586), .B(n10585), .Z(n10593) );
  XNOR U10891 ( .A(n10592), .B(n10593), .Z(n10594) );
  XNOR U10892 ( .A(n10595), .B(n10594), .Z(n10628) );
  XNOR U10893 ( .A(n10628), .B(sreg[1272]), .Z(n10630) );
  NAND U10894 ( .A(n10587), .B(sreg[1271]), .Z(n10591) );
  OR U10895 ( .A(n10589), .B(n10588), .Z(n10590) );
  AND U10896 ( .A(n10591), .B(n10590), .Z(n10629) );
  XOR U10897 ( .A(n10630), .B(n10629), .Z(c[1272]) );
  NANDN U10898 ( .A(n10593), .B(n10592), .Z(n10597) );
  NAND U10899 ( .A(n10595), .B(n10594), .Z(n10596) );
  NAND U10900 ( .A(n10597), .B(n10596), .Z(n10636) );
  NAND U10901 ( .A(b[0]), .B(a[257]), .Z(n10598) );
  XNOR U10902 ( .A(b[1]), .B(n10598), .Z(n10600) );
  NAND U10903 ( .A(n51), .B(a[256]), .Z(n10599) );
  AND U10904 ( .A(n10600), .B(n10599), .Z(n10653) );
  XOR U10905 ( .A(a[253]), .B(n42197), .Z(n10642) );
  NANDN U10906 ( .A(n10642), .B(n42173), .Z(n10603) );
  NANDN U10907 ( .A(n10601), .B(n42172), .Z(n10602) );
  NAND U10908 ( .A(n10603), .B(n10602), .Z(n10651) );
  NAND U10909 ( .A(b[7]), .B(a[249]), .Z(n10652) );
  XNOR U10910 ( .A(n10651), .B(n10652), .Z(n10654) );
  XOR U10911 ( .A(n10653), .B(n10654), .Z(n10660) );
  NANDN U10912 ( .A(n10604), .B(n42093), .Z(n10606) );
  XOR U10913 ( .A(n42134), .B(a[255]), .Z(n10645) );
  NANDN U10914 ( .A(n10645), .B(n42095), .Z(n10605) );
  NAND U10915 ( .A(n10606), .B(n10605), .Z(n10658) );
  NANDN U10916 ( .A(n10607), .B(n42231), .Z(n10609) );
  XOR U10917 ( .A(n183), .B(a[251]), .Z(n10648) );
  NANDN U10918 ( .A(n10648), .B(n42234), .Z(n10608) );
  AND U10919 ( .A(n10609), .B(n10608), .Z(n10657) );
  XNOR U10920 ( .A(n10658), .B(n10657), .Z(n10659) );
  XNOR U10921 ( .A(n10660), .B(n10659), .Z(n10664) );
  NANDN U10922 ( .A(n10611), .B(n10610), .Z(n10615) );
  NAND U10923 ( .A(n10613), .B(n10612), .Z(n10614) );
  AND U10924 ( .A(n10615), .B(n10614), .Z(n10663) );
  XOR U10925 ( .A(n10664), .B(n10663), .Z(n10665) );
  NANDN U10926 ( .A(n10617), .B(n10616), .Z(n10621) );
  NANDN U10927 ( .A(n10619), .B(n10618), .Z(n10620) );
  NAND U10928 ( .A(n10621), .B(n10620), .Z(n10666) );
  XOR U10929 ( .A(n10665), .B(n10666), .Z(n10633) );
  OR U10930 ( .A(n10623), .B(n10622), .Z(n10627) );
  NANDN U10931 ( .A(n10625), .B(n10624), .Z(n10626) );
  NAND U10932 ( .A(n10627), .B(n10626), .Z(n10634) );
  XNOR U10933 ( .A(n10633), .B(n10634), .Z(n10635) );
  XNOR U10934 ( .A(n10636), .B(n10635), .Z(n10669) );
  XNOR U10935 ( .A(n10669), .B(sreg[1273]), .Z(n10671) );
  NAND U10936 ( .A(n10628), .B(sreg[1272]), .Z(n10632) );
  OR U10937 ( .A(n10630), .B(n10629), .Z(n10631) );
  AND U10938 ( .A(n10632), .B(n10631), .Z(n10670) );
  XOR U10939 ( .A(n10671), .B(n10670), .Z(c[1273]) );
  NANDN U10940 ( .A(n10634), .B(n10633), .Z(n10638) );
  NAND U10941 ( .A(n10636), .B(n10635), .Z(n10637) );
  NAND U10942 ( .A(n10638), .B(n10637), .Z(n10677) );
  NAND U10943 ( .A(b[0]), .B(a[258]), .Z(n10639) );
  XNOR U10944 ( .A(b[1]), .B(n10639), .Z(n10641) );
  NAND U10945 ( .A(n51), .B(a[257]), .Z(n10640) );
  AND U10946 ( .A(n10641), .B(n10640), .Z(n10694) );
  XOR U10947 ( .A(a[254]), .B(n42197), .Z(n10683) );
  NANDN U10948 ( .A(n10683), .B(n42173), .Z(n10644) );
  NANDN U10949 ( .A(n10642), .B(n42172), .Z(n10643) );
  NAND U10950 ( .A(n10644), .B(n10643), .Z(n10692) );
  NAND U10951 ( .A(b[7]), .B(a[250]), .Z(n10693) );
  XNOR U10952 ( .A(n10692), .B(n10693), .Z(n10695) );
  XOR U10953 ( .A(n10694), .B(n10695), .Z(n10701) );
  NANDN U10954 ( .A(n10645), .B(n42093), .Z(n10647) );
  XOR U10955 ( .A(n42134), .B(a[256]), .Z(n10686) );
  NANDN U10956 ( .A(n10686), .B(n42095), .Z(n10646) );
  NAND U10957 ( .A(n10647), .B(n10646), .Z(n10699) );
  NANDN U10958 ( .A(n10648), .B(n42231), .Z(n10650) );
  XOR U10959 ( .A(n183), .B(a[252]), .Z(n10689) );
  NANDN U10960 ( .A(n10689), .B(n42234), .Z(n10649) );
  AND U10961 ( .A(n10650), .B(n10649), .Z(n10698) );
  XNOR U10962 ( .A(n10699), .B(n10698), .Z(n10700) );
  XNOR U10963 ( .A(n10701), .B(n10700), .Z(n10705) );
  NANDN U10964 ( .A(n10652), .B(n10651), .Z(n10656) );
  NAND U10965 ( .A(n10654), .B(n10653), .Z(n10655) );
  AND U10966 ( .A(n10656), .B(n10655), .Z(n10704) );
  XOR U10967 ( .A(n10705), .B(n10704), .Z(n10706) );
  NANDN U10968 ( .A(n10658), .B(n10657), .Z(n10662) );
  NANDN U10969 ( .A(n10660), .B(n10659), .Z(n10661) );
  NAND U10970 ( .A(n10662), .B(n10661), .Z(n10707) );
  XOR U10971 ( .A(n10706), .B(n10707), .Z(n10674) );
  OR U10972 ( .A(n10664), .B(n10663), .Z(n10668) );
  NANDN U10973 ( .A(n10666), .B(n10665), .Z(n10667) );
  NAND U10974 ( .A(n10668), .B(n10667), .Z(n10675) );
  XNOR U10975 ( .A(n10674), .B(n10675), .Z(n10676) );
  XNOR U10976 ( .A(n10677), .B(n10676), .Z(n10710) );
  XNOR U10977 ( .A(n10710), .B(sreg[1274]), .Z(n10712) );
  NAND U10978 ( .A(n10669), .B(sreg[1273]), .Z(n10673) );
  OR U10979 ( .A(n10671), .B(n10670), .Z(n10672) );
  AND U10980 ( .A(n10673), .B(n10672), .Z(n10711) );
  XOR U10981 ( .A(n10712), .B(n10711), .Z(c[1274]) );
  NANDN U10982 ( .A(n10675), .B(n10674), .Z(n10679) );
  NAND U10983 ( .A(n10677), .B(n10676), .Z(n10678) );
  NAND U10984 ( .A(n10679), .B(n10678), .Z(n10718) );
  NAND U10985 ( .A(b[0]), .B(a[259]), .Z(n10680) );
  XNOR U10986 ( .A(b[1]), .B(n10680), .Z(n10682) );
  NAND U10987 ( .A(n52), .B(a[258]), .Z(n10681) );
  AND U10988 ( .A(n10682), .B(n10681), .Z(n10735) );
  XOR U10989 ( .A(a[255]), .B(n42197), .Z(n10724) );
  NANDN U10990 ( .A(n10724), .B(n42173), .Z(n10685) );
  NANDN U10991 ( .A(n10683), .B(n42172), .Z(n10684) );
  NAND U10992 ( .A(n10685), .B(n10684), .Z(n10733) );
  NAND U10993 ( .A(b[7]), .B(a[251]), .Z(n10734) );
  XNOR U10994 ( .A(n10733), .B(n10734), .Z(n10736) );
  XOR U10995 ( .A(n10735), .B(n10736), .Z(n10742) );
  NANDN U10996 ( .A(n10686), .B(n42093), .Z(n10688) );
  XOR U10997 ( .A(n42134), .B(a[257]), .Z(n10727) );
  NANDN U10998 ( .A(n10727), .B(n42095), .Z(n10687) );
  NAND U10999 ( .A(n10688), .B(n10687), .Z(n10740) );
  NANDN U11000 ( .A(n10689), .B(n42231), .Z(n10691) );
  XOR U11001 ( .A(n183), .B(a[253]), .Z(n10730) );
  NANDN U11002 ( .A(n10730), .B(n42234), .Z(n10690) );
  AND U11003 ( .A(n10691), .B(n10690), .Z(n10739) );
  XNOR U11004 ( .A(n10740), .B(n10739), .Z(n10741) );
  XNOR U11005 ( .A(n10742), .B(n10741), .Z(n10746) );
  NANDN U11006 ( .A(n10693), .B(n10692), .Z(n10697) );
  NAND U11007 ( .A(n10695), .B(n10694), .Z(n10696) );
  AND U11008 ( .A(n10697), .B(n10696), .Z(n10745) );
  XOR U11009 ( .A(n10746), .B(n10745), .Z(n10747) );
  NANDN U11010 ( .A(n10699), .B(n10698), .Z(n10703) );
  NANDN U11011 ( .A(n10701), .B(n10700), .Z(n10702) );
  NAND U11012 ( .A(n10703), .B(n10702), .Z(n10748) );
  XOR U11013 ( .A(n10747), .B(n10748), .Z(n10715) );
  OR U11014 ( .A(n10705), .B(n10704), .Z(n10709) );
  NANDN U11015 ( .A(n10707), .B(n10706), .Z(n10708) );
  NAND U11016 ( .A(n10709), .B(n10708), .Z(n10716) );
  XNOR U11017 ( .A(n10715), .B(n10716), .Z(n10717) );
  XNOR U11018 ( .A(n10718), .B(n10717), .Z(n10751) );
  XNOR U11019 ( .A(n10751), .B(sreg[1275]), .Z(n10753) );
  NAND U11020 ( .A(n10710), .B(sreg[1274]), .Z(n10714) );
  OR U11021 ( .A(n10712), .B(n10711), .Z(n10713) );
  AND U11022 ( .A(n10714), .B(n10713), .Z(n10752) );
  XOR U11023 ( .A(n10753), .B(n10752), .Z(c[1275]) );
  NANDN U11024 ( .A(n10716), .B(n10715), .Z(n10720) );
  NAND U11025 ( .A(n10718), .B(n10717), .Z(n10719) );
  NAND U11026 ( .A(n10720), .B(n10719), .Z(n10759) );
  NAND U11027 ( .A(b[0]), .B(a[260]), .Z(n10721) );
  XNOR U11028 ( .A(b[1]), .B(n10721), .Z(n10723) );
  NAND U11029 ( .A(n52), .B(a[259]), .Z(n10722) );
  AND U11030 ( .A(n10723), .B(n10722), .Z(n10776) );
  XOR U11031 ( .A(a[256]), .B(n42197), .Z(n10765) );
  NANDN U11032 ( .A(n10765), .B(n42173), .Z(n10726) );
  NANDN U11033 ( .A(n10724), .B(n42172), .Z(n10725) );
  NAND U11034 ( .A(n10726), .B(n10725), .Z(n10774) );
  NAND U11035 ( .A(b[7]), .B(a[252]), .Z(n10775) );
  XNOR U11036 ( .A(n10774), .B(n10775), .Z(n10777) );
  XOR U11037 ( .A(n10776), .B(n10777), .Z(n10783) );
  NANDN U11038 ( .A(n10727), .B(n42093), .Z(n10729) );
  XOR U11039 ( .A(n42134), .B(a[258]), .Z(n10768) );
  NANDN U11040 ( .A(n10768), .B(n42095), .Z(n10728) );
  NAND U11041 ( .A(n10729), .B(n10728), .Z(n10781) );
  NANDN U11042 ( .A(n10730), .B(n42231), .Z(n10732) );
  XOR U11043 ( .A(n183), .B(a[254]), .Z(n10771) );
  NANDN U11044 ( .A(n10771), .B(n42234), .Z(n10731) );
  AND U11045 ( .A(n10732), .B(n10731), .Z(n10780) );
  XNOR U11046 ( .A(n10781), .B(n10780), .Z(n10782) );
  XNOR U11047 ( .A(n10783), .B(n10782), .Z(n10787) );
  NANDN U11048 ( .A(n10734), .B(n10733), .Z(n10738) );
  NAND U11049 ( .A(n10736), .B(n10735), .Z(n10737) );
  AND U11050 ( .A(n10738), .B(n10737), .Z(n10786) );
  XOR U11051 ( .A(n10787), .B(n10786), .Z(n10788) );
  NANDN U11052 ( .A(n10740), .B(n10739), .Z(n10744) );
  NANDN U11053 ( .A(n10742), .B(n10741), .Z(n10743) );
  NAND U11054 ( .A(n10744), .B(n10743), .Z(n10789) );
  XOR U11055 ( .A(n10788), .B(n10789), .Z(n10756) );
  OR U11056 ( .A(n10746), .B(n10745), .Z(n10750) );
  NANDN U11057 ( .A(n10748), .B(n10747), .Z(n10749) );
  NAND U11058 ( .A(n10750), .B(n10749), .Z(n10757) );
  XNOR U11059 ( .A(n10756), .B(n10757), .Z(n10758) );
  XNOR U11060 ( .A(n10759), .B(n10758), .Z(n10792) );
  XNOR U11061 ( .A(n10792), .B(sreg[1276]), .Z(n10794) );
  NAND U11062 ( .A(n10751), .B(sreg[1275]), .Z(n10755) );
  OR U11063 ( .A(n10753), .B(n10752), .Z(n10754) );
  AND U11064 ( .A(n10755), .B(n10754), .Z(n10793) );
  XOR U11065 ( .A(n10794), .B(n10793), .Z(c[1276]) );
  NANDN U11066 ( .A(n10757), .B(n10756), .Z(n10761) );
  NAND U11067 ( .A(n10759), .B(n10758), .Z(n10760) );
  NAND U11068 ( .A(n10761), .B(n10760), .Z(n10800) );
  NAND U11069 ( .A(b[0]), .B(a[261]), .Z(n10762) );
  XNOR U11070 ( .A(b[1]), .B(n10762), .Z(n10764) );
  NAND U11071 ( .A(n52), .B(a[260]), .Z(n10763) );
  AND U11072 ( .A(n10764), .B(n10763), .Z(n10817) );
  XOR U11073 ( .A(a[257]), .B(n42197), .Z(n10806) );
  NANDN U11074 ( .A(n10806), .B(n42173), .Z(n10767) );
  NANDN U11075 ( .A(n10765), .B(n42172), .Z(n10766) );
  NAND U11076 ( .A(n10767), .B(n10766), .Z(n10815) );
  NAND U11077 ( .A(b[7]), .B(a[253]), .Z(n10816) );
  XNOR U11078 ( .A(n10815), .B(n10816), .Z(n10818) );
  XOR U11079 ( .A(n10817), .B(n10818), .Z(n10824) );
  NANDN U11080 ( .A(n10768), .B(n42093), .Z(n10770) );
  XOR U11081 ( .A(n42134), .B(a[259]), .Z(n10809) );
  NANDN U11082 ( .A(n10809), .B(n42095), .Z(n10769) );
  NAND U11083 ( .A(n10770), .B(n10769), .Z(n10822) );
  NANDN U11084 ( .A(n10771), .B(n42231), .Z(n10773) );
  XOR U11085 ( .A(n183), .B(a[255]), .Z(n10812) );
  NANDN U11086 ( .A(n10812), .B(n42234), .Z(n10772) );
  AND U11087 ( .A(n10773), .B(n10772), .Z(n10821) );
  XNOR U11088 ( .A(n10822), .B(n10821), .Z(n10823) );
  XNOR U11089 ( .A(n10824), .B(n10823), .Z(n10828) );
  NANDN U11090 ( .A(n10775), .B(n10774), .Z(n10779) );
  NAND U11091 ( .A(n10777), .B(n10776), .Z(n10778) );
  AND U11092 ( .A(n10779), .B(n10778), .Z(n10827) );
  XOR U11093 ( .A(n10828), .B(n10827), .Z(n10829) );
  NANDN U11094 ( .A(n10781), .B(n10780), .Z(n10785) );
  NANDN U11095 ( .A(n10783), .B(n10782), .Z(n10784) );
  NAND U11096 ( .A(n10785), .B(n10784), .Z(n10830) );
  XOR U11097 ( .A(n10829), .B(n10830), .Z(n10797) );
  OR U11098 ( .A(n10787), .B(n10786), .Z(n10791) );
  NANDN U11099 ( .A(n10789), .B(n10788), .Z(n10790) );
  NAND U11100 ( .A(n10791), .B(n10790), .Z(n10798) );
  XNOR U11101 ( .A(n10797), .B(n10798), .Z(n10799) );
  XNOR U11102 ( .A(n10800), .B(n10799), .Z(n10833) );
  XNOR U11103 ( .A(n10833), .B(sreg[1277]), .Z(n10835) );
  NAND U11104 ( .A(n10792), .B(sreg[1276]), .Z(n10796) );
  OR U11105 ( .A(n10794), .B(n10793), .Z(n10795) );
  AND U11106 ( .A(n10796), .B(n10795), .Z(n10834) );
  XOR U11107 ( .A(n10835), .B(n10834), .Z(c[1277]) );
  NANDN U11108 ( .A(n10798), .B(n10797), .Z(n10802) );
  NAND U11109 ( .A(n10800), .B(n10799), .Z(n10801) );
  NAND U11110 ( .A(n10802), .B(n10801), .Z(n10841) );
  NAND U11111 ( .A(b[0]), .B(a[262]), .Z(n10803) );
  XNOR U11112 ( .A(b[1]), .B(n10803), .Z(n10805) );
  NAND U11113 ( .A(n52), .B(a[261]), .Z(n10804) );
  AND U11114 ( .A(n10805), .B(n10804), .Z(n10858) );
  XOR U11115 ( .A(a[258]), .B(n42197), .Z(n10847) );
  NANDN U11116 ( .A(n10847), .B(n42173), .Z(n10808) );
  NANDN U11117 ( .A(n10806), .B(n42172), .Z(n10807) );
  NAND U11118 ( .A(n10808), .B(n10807), .Z(n10856) );
  NAND U11119 ( .A(b[7]), .B(a[254]), .Z(n10857) );
  XNOR U11120 ( .A(n10856), .B(n10857), .Z(n10859) );
  XOR U11121 ( .A(n10858), .B(n10859), .Z(n10865) );
  NANDN U11122 ( .A(n10809), .B(n42093), .Z(n10811) );
  XOR U11123 ( .A(n42134), .B(a[260]), .Z(n10850) );
  NANDN U11124 ( .A(n10850), .B(n42095), .Z(n10810) );
  NAND U11125 ( .A(n10811), .B(n10810), .Z(n10863) );
  NANDN U11126 ( .A(n10812), .B(n42231), .Z(n10814) );
  XOR U11127 ( .A(n183), .B(a[256]), .Z(n10853) );
  NANDN U11128 ( .A(n10853), .B(n42234), .Z(n10813) );
  AND U11129 ( .A(n10814), .B(n10813), .Z(n10862) );
  XNOR U11130 ( .A(n10863), .B(n10862), .Z(n10864) );
  XNOR U11131 ( .A(n10865), .B(n10864), .Z(n10869) );
  NANDN U11132 ( .A(n10816), .B(n10815), .Z(n10820) );
  NAND U11133 ( .A(n10818), .B(n10817), .Z(n10819) );
  AND U11134 ( .A(n10820), .B(n10819), .Z(n10868) );
  XOR U11135 ( .A(n10869), .B(n10868), .Z(n10870) );
  NANDN U11136 ( .A(n10822), .B(n10821), .Z(n10826) );
  NANDN U11137 ( .A(n10824), .B(n10823), .Z(n10825) );
  NAND U11138 ( .A(n10826), .B(n10825), .Z(n10871) );
  XOR U11139 ( .A(n10870), .B(n10871), .Z(n10838) );
  OR U11140 ( .A(n10828), .B(n10827), .Z(n10832) );
  NANDN U11141 ( .A(n10830), .B(n10829), .Z(n10831) );
  NAND U11142 ( .A(n10832), .B(n10831), .Z(n10839) );
  XNOR U11143 ( .A(n10838), .B(n10839), .Z(n10840) );
  XNOR U11144 ( .A(n10841), .B(n10840), .Z(n10874) );
  XNOR U11145 ( .A(n10874), .B(sreg[1278]), .Z(n10876) );
  NAND U11146 ( .A(n10833), .B(sreg[1277]), .Z(n10837) );
  OR U11147 ( .A(n10835), .B(n10834), .Z(n10836) );
  AND U11148 ( .A(n10837), .B(n10836), .Z(n10875) );
  XOR U11149 ( .A(n10876), .B(n10875), .Z(c[1278]) );
  NANDN U11150 ( .A(n10839), .B(n10838), .Z(n10843) );
  NAND U11151 ( .A(n10841), .B(n10840), .Z(n10842) );
  NAND U11152 ( .A(n10843), .B(n10842), .Z(n10882) );
  NAND U11153 ( .A(b[0]), .B(a[263]), .Z(n10844) );
  XNOR U11154 ( .A(b[1]), .B(n10844), .Z(n10846) );
  NAND U11155 ( .A(n52), .B(a[262]), .Z(n10845) );
  AND U11156 ( .A(n10846), .B(n10845), .Z(n10899) );
  XOR U11157 ( .A(a[259]), .B(n42197), .Z(n10888) );
  NANDN U11158 ( .A(n10888), .B(n42173), .Z(n10849) );
  NANDN U11159 ( .A(n10847), .B(n42172), .Z(n10848) );
  NAND U11160 ( .A(n10849), .B(n10848), .Z(n10897) );
  NAND U11161 ( .A(b[7]), .B(a[255]), .Z(n10898) );
  XNOR U11162 ( .A(n10897), .B(n10898), .Z(n10900) );
  XOR U11163 ( .A(n10899), .B(n10900), .Z(n10906) );
  NANDN U11164 ( .A(n10850), .B(n42093), .Z(n10852) );
  XOR U11165 ( .A(n42134), .B(a[261]), .Z(n10891) );
  NANDN U11166 ( .A(n10891), .B(n42095), .Z(n10851) );
  NAND U11167 ( .A(n10852), .B(n10851), .Z(n10904) );
  NANDN U11168 ( .A(n10853), .B(n42231), .Z(n10855) );
  XOR U11169 ( .A(n183), .B(a[257]), .Z(n10894) );
  NANDN U11170 ( .A(n10894), .B(n42234), .Z(n10854) );
  AND U11171 ( .A(n10855), .B(n10854), .Z(n10903) );
  XNOR U11172 ( .A(n10904), .B(n10903), .Z(n10905) );
  XNOR U11173 ( .A(n10906), .B(n10905), .Z(n10910) );
  NANDN U11174 ( .A(n10857), .B(n10856), .Z(n10861) );
  NAND U11175 ( .A(n10859), .B(n10858), .Z(n10860) );
  AND U11176 ( .A(n10861), .B(n10860), .Z(n10909) );
  XOR U11177 ( .A(n10910), .B(n10909), .Z(n10911) );
  NANDN U11178 ( .A(n10863), .B(n10862), .Z(n10867) );
  NANDN U11179 ( .A(n10865), .B(n10864), .Z(n10866) );
  NAND U11180 ( .A(n10867), .B(n10866), .Z(n10912) );
  XOR U11181 ( .A(n10911), .B(n10912), .Z(n10879) );
  OR U11182 ( .A(n10869), .B(n10868), .Z(n10873) );
  NANDN U11183 ( .A(n10871), .B(n10870), .Z(n10872) );
  NAND U11184 ( .A(n10873), .B(n10872), .Z(n10880) );
  XNOR U11185 ( .A(n10879), .B(n10880), .Z(n10881) );
  XNOR U11186 ( .A(n10882), .B(n10881), .Z(n10915) );
  XNOR U11187 ( .A(n10915), .B(sreg[1279]), .Z(n10917) );
  NAND U11188 ( .A(n10874), .B(sreg[1278]), .Z(n10878) );
  OR U11189 ( .A(n10876), .B(n10875), .Z(n10877) );
  AND U11190 ( .A(n10878), .B(n10877), .Z(n10916) );
  XOR U11191 ( .A(n10917), .B(n10916), .Z(c[1279]) );
  NANDN U11192 ( .A(n10880), .B(n10879), .Z(n10884) );
  NAND U11193 ( .A(n10882), .B(n10881), .Z(n10883) );
  NAND U11194 ( .A(n10884), .B(n10883), .Z(n10923) );
  NAND U11195 ( .A(b[0]), .B(a[264]), .Z(n10885) );
  XNOR U11196 ( .A(b[1]), .B(n10885), .Z(n10887) );
  NAND U11197 ( .A(n52), .B(a[263]), .Z(n10886) );
  AND U11198 ( .A(n10887), .B(n10886), .Z(n10940) );
  XOR U11199 ( .A(a[260]), .B(n42197), .Z(n10929) );
  NANDN U11200 ( .A(n10929), .B(n42173), .Z(n10890) );
  NANDN U11201 ( .A(n10888), .B(n42172), .Z(n10889) );
  NAND U11202 ( .A(n10890), .B(n10889), .Z(n10938) );
  NAND U11203 ( .A(b[7]), .B(a[256]), .Z(n10939) );
  XNOR U11204 ( .A(n10938), .B(n10939), .Z(n10941) );
  XOR U11205 ( .A(n10940), .B(n10941), .Z(n10947) );
  NANDN U11206 ( .A(n10891), .B(n42093), .Z(n10893) );
  XOR U11207 ( .A(n42134), .B(a[262]), .Z(n10932) );
  NANDN U11208 ( .A(n10932), .B(n42095), .Z(n10892) );
  NAND U11209 ( .A(n10893), .B(n10892), .Z(n10945) );
  NANDN U11210 ( .A(n10894), .B(n42231), .Z(n10896) );
  XOR U11211 ( .A(n183), .B(a[258]), .Z(n10935) );
  NANDN U11212 ( .A(n10935), .B(n42234), .Z(n10895) );
  AND U11213 ( .A(n10896), .B(n10895), .Z(n10944) );
  XNOR U11214 ( .A(n10945), .B(n10944), .Z(n10946) );
  XNOR U11215 ( .A(n10947), .B(n10946), .Z(n10951) );
  NANDN U11216 ( .A(n10898), .B(n10897), .Z(n10902) );
  NAND U11217 ( .A(n10900), .B(n10899), .Z(n10901) );
  AND U11218 ( .A(n10902), .B(n10901), .Z(n10950) );
  XOR U11219 ( .A(n10951), .B(n10950), .Z(n10952) );
  NANDN U11220 ( .A(n10904), .B(n10903), .Z(n10908) );
  NANDN U11221 ( .A(n10906), .B(n10905), .Z(n10907) );
  NAND U11222 ( .A(n10908), .B(n10907), .Z(n10953) );
  XOR U11223 ( .A(n10952), .B(n10953), .Z(n10920) );
  OR U11224 ( .A(n10910), .B(n10909), .Z(n10914) );
  NANDN U11225 ( .A(n10912), .B(n10911), .Z(n10913) );
  NAND U11226 ( .A(n10914), .B(n10913), .Z(n10921) );
  XNOR U11227 ( .A(n10920), .B(n10921), .Z(n10922) );
  XNOR U11228 ( .A(n10923), .B(n10922), .Z(n10956) );
  XNOR U11229 ( .A(n10956), .B(sreg[1280]), .Z(n10958) );
  NAND U11230 ( .A(n10915), .B(sreg[1279]), .Z(n10919) );
  OR U11231 ( .A(n10917), .B(n10916), .Z(n10918) );
  AND U11232 ( .A(n10919), .B(n10918), .Z(n10957) );
  XOR U11233 ( .A(n10958), .B(n10957), .Z(c[1280]) );
  NANDN U11234 ( .A(n10921), .B(n10920), .Z(n10925) );
  NAND U11235 ( .A(n10923), .B(n10922), .Z(n10924) );
  NAND U11236 ( .A(n10925), .B(n10924), .Z(n10964) );
  NAND U11237 ( .A(b[0]), .B(a[265]), .Z(n10926) );
  XNOR U11238 ( .A(b[1]), .B(n10926), .Z(n10928) );
  NAND U11239 ( .A(n52), .B(a[264]), .Z(n10927) );
  AND U11240 ( .A(n10928), .B(n10927), .Z(n10981) );
  XOR U11241 ( .A(a[261]), .B(n42197), .Z(n10970) );
  NANDN U11242 ( .A(n10970), .B(n42173), .Z(n10931) );
  NANDN U11243 ( .A(n10929), .B(n42172), .Z(n10930) );
  NAND U11244 ( .A(n10931), .B(n10930), .Z(n10979) );
  NAND U11245 ( .A(b[7]), .B(a[257]), .Z(n10980) );
  XNOR U11246 ( .A(n10979), .B(n10980), .Z(n10982) );
  XOR U11247 ( .A(n10981), .B(n10982), .Z(n10988) );
  NANDN U11248 ( .A(n10932), .B(n42093), .Z(n10934) );
  XOR U11249 ( .A(n42134), .B(a[263]), .Z(n10973) );
  NANDN U11250 ( .A(n10973), .B(n42095), .Z(n10933) );
  NAND U11251 ( .A(n10934), .B(n10933), .Z(n10986) );
  NANDN U11252 ( .A(n10935), .B(n42231), .Z(n10937) );
  XOR U11253 ( .A(n183), .B(a[259]), .Z(n10976) );
  NANDN U11254 ( .A(n10976), .B(n42234), .Z(n10936) );
  AND U11255 ( .A(n10937), .B(n10936), .Z(n10985) );
  XNOR U11256 ( .A(n10986), .B(n10985), .Z(n10987) );
  XNOR U11257 ( .A(n10988), .B(n10987), .Z(n10992) );
  NANDN U11258 ( .A(n10939), .B(n10938), .Z(n10943) );
  NAND U11259 ( .A(n10941), .B(n10940), .Z(n10942) );
  AND U11260 ( .A(n10943), .B(n10942), .Z(n10991) );
  XOR U11261 ( .A(n10992), .B(n10991), .Z(n10993) );
  NANDN U11262 ( .A(n10945), .B(n10944), .Z(n10949) );
  NANDN U11263 ( .A(n10947), .B(n10946), .Z(n10948) );
  NAND U11264 ( .A(n10949), .B(n10948), .Z(n10994) );
  XOR U11265 ( .A(n10993), .B(n10994), .Z(n10961) );
  OR U11266 ( .A(n10951), .B(n10950), .Z(n10955) );
  NANDN U11267 ( .A(n10953), .B(n10952), .Z(n10954) );
  NAND U11268 ( .A(n10955), .B(n10954), .Z(n10962) );
  XNOR U11269 ( .A(n10961), .B(n10962), .Z(n10963) );
  XNOR U11270 ( .A(n10964), .B(n10963), .Z(n10997) );
  XNOR U11271 ( .A(n10997), .B(sreg[1281]), .Z(n10999) );
  NAND U11272 ( .A(n10956), .B(sreg[1280]), .Z(n10960) );
  OR U11273 ( .A(n10958), .B(n10957), .Z(n10959) );
  AND U11274 ( .A(n10960), .B(n10959), .Z(n10998) );
  XOR U11275 ( .A(n10999), .B(n10998), .Z(c[1281]) );
  NANDN U11276 ( .A(n10962), .B(n10961), .Z(n10966) );
  NAND U11277 ( .A(n10964), .B(n10963), .Z(n10965) );
  NAND U11278 ( .A(n10966), .B(n10965), .Z(n11005) );
  NAND U11279 ( .A(b[0]), .B(a[266]), .Z(n10967) );
  XNOR U11280 ( .A(b[1]), .B(n10967), .Z(n10969) );
  NAND U11281 ( .A(n53), .B(a[265]), .Z(n10968) );
  AND U11282 ( .A(n10969), .B(n10968), .Z(n11022) );
  XOR U11283 ( .A(a[262]), .B(n42197), .Z(n11011) );
  NANDN U11284 ( .A(n11011), .B(n42173), .Z(n10972) );
  NANDN U11285 ( .A(n10970), .B(n42172), .Z(n10971) );
  NAND U11286 ( .A(n10972), .B(n10971), .Z(n11020) );
  NAND U11287 ( .A(b[7]), .B(a[258]), .Z(n11021) );
  XNOR U11288 ( .A(n11020), .B(n11021), .Z(n11023) );
  XOR U11289 ( .A(n11022), .B(n11023), .Z(n11029) );
  NANDN U11290 ( .A(n10973), .B(n42093), .Z(n10975) );
  XOR U11291 ( .A(n42134), .B(a[264]), .Z(n11014) );
  NANDN U11292 ( .A(n11014), .B(n42095), .Z(n10974) );
  NAND U11293 ( .A(n10975), .B(n10974), .Z(n11027) );
  NANDN U11294 ( .A(n10976), .B(n42231), .Z(n10978) );
  XOR U11295 ( .A(n183), .B(a[260]), .Z(n11017) );
  NANDN U11296 ( .A(n11017), .B(n42234), .Z(n10977) );
  AND U11297 ( .A(n10978), .B(n10977), .Z(n11026) );
  XNOR U11298 ( .A(n11027), .B(n11026), .Z(n11028) );
  XNOR U11299 ( .A(n11029), .B(n11028), .Z(n11033) );
  NANDN U11300 ( .A(n10980), .B(n10979), .Z(n10984) );
  NAND U11301 ( .A(n10982), .B(n10981), .Z(n10983) );
  AND U11302 ( .A(n10984), .B(n10983), .Z(n11032) );
  XOR U11303 ( .A(n11033), .B(n11032), .Z(n11034) );
  NANDN U11304 ( .A(n10986), .B(n10985), .Z(n10990) );
  NANDN U11305 ( .A(n10988), .B(n10987), .Z(n10989) );
  NAND U11306 ( .A(n10990), .B(n10989), .Z(n11035) );
  XOR U11307 ( .A(n11034), .B(n11035), .Z(n11002) );
  OR U11308 ( .A(n10992), .B(n10991), .Z(n10996) );
  NANDN U11309 ( .A(n10994), .B(n10993), .Z(n10995) );
  NAND U11310 ( .A(n10996), .B(n10995), .Z(n11003) );
  XNOR U11311 ( .A(n11002), .B(n11003), .Z(n11004) );
  XNOR U11312 ( .A(n11005), .B(n11004), .Z(n11038) );
  XNOR U11313 ( .A(n11038), .B(sreg[1282]), .Z(n11040) );
  NAND U11314 ( .A(n10997), .B(sreg[1281]), .Z(n11001) );
  OR U11315 ( .A(n10999), .B(n10998), .Z(n11000) );
  AND U11316 ( .A(n11001), .B(n11000), .Z(n11039) );
  XOR U11317 ( .A(n11040), .B(n11039), .Z(c[1282]) );
  NANDN U11318 ( .A(n11003), .B(n11002), .Z(n11007) );
  NAND U11319 ( .A(n11005), .B(n11004), .Z(n11006) );
  NAND U11320 ( .A(n11007), .B(n11006), .Z(n11046) );
  NAND U11321 ( .A(b[0]), .B(a[267]), .Z(n11008) );
  XNOR U11322 ( .A(b[1]), .B(n11008), .Z(n11010) );
  NAND U11323 ( .A(n53), .B(a[266]), .Z(n11009) );
  AND U11324 ( .A(n11010), .B(n11009), .Z(n11063) );
  XOR U11325 ( .A(a[263]), .B(n42197), .Z(n11052) );
  NANDN U11326 ( .A(n11052), .B(n42173), .Z(n11013) );
  NANDN U11327 ( .A(n11011), .B(n42172), .Z(n11012) );
  NAND U11328 ( .A(n11013), .B(n11012), .Z(n11061) );
  NAND U11329 ( .A(b[7]), .B(a[259]), .Z(n11062) );
  XNOR U11330 ( .A(n11061), .B(n11062), .Z(n11064) );
  XOR U11331 ( .A(n11063), .B(n11064), .Z(n11070) );
  NANDN U11332 ( .A(n11014), .B(n42093), .Z(n11016) );
  XOR U11333 ( .A(n42134), .B(a[265]), .Z(n11055) );
  NANDN U11334 ( .A(n11055), .B(n42095), .Z(n11015) );
  NAND U11335 ( .A(n11016), .B(n11015), .Z(n11068) );
  NANDN U11336 ( .A(n11017), .B(n42231), .Z(n11019) );
  XOR U11337 ( .A(n183), .B(a[261]), .Z(n11058) );
  NANDN U11338 ( .A(n11058), .B(n42234), .Z(n11018) );
  AND U11339 ( .A(n11019), .B(n11018), .Z(n11067) );
  XNOR U11340 ( .A(n11068), .B(n11067), .Z(n11069) );
  XNOR U11341 ( .A(n11070), .B(n11069), .Z(n11074) );
  NANDN U11342 ( .A(n11021), .B(n11020), .Z(n11025) );
  NAND U11343 ( .A(n11023), .B(n11022), .Z(n11024) );
  AND U11344 ( .A(n11025), .B(n11024), .Z(n11073) );
  XOR U11345 ( .A(n11074), .B(n11073), .Z(n11075) );
  NANDN U11346 ( .A(n11027), .B(n11026), .Z(n11031) );
  NANDN U11347 ( .A(n11029), .B(n11028), .Z(n11030) );
  NAND U11348 ( .A(n11031), .B(n11030), .Z(n11076) );
  XOR U11349 ( .A(n11075), .B(n11076), .Z(n11043) );
  OR U11350 ( .A(n11033), .B(n11032), .Z(n11037) );
  NANDN U11351 ( .A(n11035), .B(n11034), .Z(n11036) );
  NAND U11352 ( .A(n11037), .B(n11036), .Z(n11044) );
  XNOR U11353 ( .A(n11043), .B(n11044), .Z(n11045) );
  XNOR U11354 ( .A(n11046), .B(n11045), .Z(n11079) );
  XNOR U11355 ( .A(n11079), .B(sreg[1283]), .Z(n11081) );
  NAND U11356 ( .A(n11038), .B(sreg[1282]), .Z(n11042) );
  OR U11357 ( .A(n11040), .B(n11039), .Z(n11041) );
  AND U11358 ( .A(n11042), .B(n11041), .Z(n11080) );
  XOR U11359 ( .A(n11081), .B(n11080), .Z(c[1283]) );
  NANDN U11360 ( .A(n11044), .B(n11043), .Z(n11048) );
  NAND U11361 ( .A(n11046), .B(n11045), .Z(n11047) );
  NAND U11362 ( .A(n11048), .B(n11047), .Z(n11087) );
  NAND U11363 ( .A(b[0]), .B(a[268]), .Z(n11049) );
  XNOR U11364 ( .A(b[1]), .B(n11049), .Z(n11051) );
  NAND U11365 ( .A(n53), .B(a[267]), .Z(n11050) );
  AND U11366 ( .A(n11051), .B(n11050), .Z(n11104) );
  XOR U11367 ( .A(a[264]), .B(n42197), .Z(n11093) );
  NANDN U11368 ( .A(n11093), .B(n42173), .Z(n11054) );
  NANDN U11369 ( .A(n11052), .B(n42172), .Z(n11053) );
  NAND U11370 ( .A(n11054), .B(n11053), .Z(n11102) );
  NAND U11371 ( .A(b[7]), .B(a[260]), .Z(n11103) );
  XNOR U11372 ( .A(n11102), .B(n11103), .Z(n11105) );
  XOR U11373 ( .A(n11104), .B(n11105), .Z(n11111) );
  NANDN U11374 ( .A(n11055), .B(n42093), .Z(n11057) );
  XOR U11375 ( .A(n42134), .B(a[266]), .Z(n11096) );
  NANDN U11376 ( .A(n11096), .B(n42095), .Z(n11056) );
  NAND U11377 ( .A(n11057), .B(n11056), .Z(n11109) );
  NANDN U11378 ( .A(n11058), .B(n42231), .Z(n11060) );
  XOR U11379 ( .A(n183), .B(a[262]), .Z(n11099) );
  NANDN U11380 ( .A(n11099), .B(n42234), .Z(n11059) );
  AND U11381 ( .A(n11060), .B(n11059), .Z(n11108) );
  XNOR U11382 ( .A(n11109), .B(n11108), .Z(n11110) );
  XNOR U11383 ( .A(n11111), .B(n11110), .Z(n11115) );
  NANDN U11384 ( .A(n11062), .B(n11061), .Z(n11066) );
  NAND U11385 ( .A(n11064), .B(n11063), .Z(n11065) );
  AND U11386 ( .A(n11066), .B(n11065), .Z(n11114) );
  XOR U11387 ( .A(n11115), .B(n11114), .Z(n11116) );
  NANDN U11388 ( .A(n11068), .B(n11067), .Z(n11072) );
  NANDN U11389 ( .A(n11070), .B(n11069), .Z(n11071) );
  NAND U11390 ( .A(n11072), .B(n11071), .Z(n11117) );
  XOR U11391 ( .A(n11116), .B(n11117), .Z(n11084) );
  OR U11392 ( .A(n11074), .B(n11073), .Z(n11078) );
  NANDN U11393 ( .A(n11076), .B(n11075), .Z(n11077) );
  NAND U11394 ( .A(n11078), .B(n11077), .Z(n11085) );
  XNOR U11395 ( .A(n11084), .B(n11085), .Z(n11086) );
  XNOR U11396 ( .A(n11087), .B(n11086), .Z(n11120) );
  XNOR U11397 ( .A(n11120), .B(sreg[1284]), .Z(n11122) );
  NAND U11398 ( .A(n11079), .B(sreg[1283]), .Z(n11083) );
  OR U11399 ( .A(n11081), .B(n11080), .Z(n11082) );
  AND U11400 ( .A(n11083), .B(n11082), .Z(n11121) );
  XOR U11401 ( .A(n11122), .B(n11121), .Z(c[1284]) );
  NANDN U11402 ( .A(n11085), .B(n11084), .Z(n11089) );
  NAND U11403 ( .A(n11087), .B(n11086), .Z(n11088) );
  NAND U11404 ( .A(n11089), .B(n11088), .Z(n11128) );
  NAND U11405 ( .A(b[0]), .B(a[269]), .Z(n11090) );
  XNOR U11406 ( .A(b[1]), .B(n11090), .Z(n11092) );
  NAND U11407 ( .A(n53), .B(a[268]), .Z(n11091) );
  AND U11408 ( .A(n11092), .B(n11091), .Z(n11145) );
  XOR U11409 ( .A(a[265]), .B(n42197), .Z(n11134) );
  NANDN U11410 ( .A(n11134), .B(n42173), .Z(n11095) );
  NANDN U11411 ( .A(n11093), .B(n42172), .Z(n11094) );
  NAND U11412 ( .A(n11095), .B(n11094), .Z(n11143) );
  NAND U11413 ( .A(b[7]), .B(a[261]), .Z(n11144) );
  XNOR U11414 ( .A(n11143), .B(n11144), .Z(n11146) );
  XOR U11415 ( .A(n11145), .B(n11146), .Z(n11152) );
  NANDN U11416 ( .A(n11096), .B(n42093), .Z(n11098) );
  XOR U11417 ( .A(n42134), .B(a[267]), .Z(n11137) );
  NANDN U11418 ( .A(n11137), .B(n42095), .Z(n11097) );
  NAND U11419 ( .A(n11098), .B(n11097), .Z(n11150) );
  NANDN U11420 ( .A(n11099), .B(n42231), .Z(n11101) );
  XOR U11421 ( .A(n184), .B(a[263]), .Z(n11140) );
  NANDN U11422 ( .A(n11140), .B(n42234), .Z(n11100) );
  AND U11423 ( .A(n11101), .B(n11100), .Z(n11149) );
  XNOR U11424 ( .A(n11150), .B(n11149), .Z(n11151) );
  XNOR U11425 ( .A(n11152), .B(n11151), .Z(n11156) );
  NANDN U11426 ( .A(n11103), .B(n11102), .Z(n11107) );
  NAND U11427 ( .A(n11105), .B(n11104), .Z(n11106) );
  AND U11428 ( .A(n11107), .B(n11106), .Z(n11155) );
  XOR U11429 ( .A(n11156), .B(n11155), .Z(n11157) );
  NANDN U11430 ( .A(n11109), .B(n11108), .Z(n11113) );
  NANDN U11431 ( .A(n11111), .B(n11110), .Z(n11112) );
  NAND U11432 ( .A(n11113), .B(n11112), .Z(n11158) );
  XOR U11433 ( .A(n11157), .B(n11158), .Z(n11125) );
  OR U11434 ( .A(n11115), .B(n11114), .Z(n11119) );
  NANDN U11435 ( .A(n11117), .B(n11116), .Z(n11118) );
  NAND U11436 ( .A(n11119), .B(n11118), .Z(n11126) );
  XNOR U11437 ( .A(n11125), .B(n11126), .Z(n11127) );
  XNOR U11438 ( .A(n11128), .B(n11127), .Z(n11161) );
  XNOR U11439 ( .A(n11161), .B(sreg[1285]), .Z(n11163) );
  NAND U11440 ( .A(n11120), .B(sreg[1284]), .Z(n11124) );
  OR U11441 ( .A(n11122), .B(n11121), .Z(n11123) );
  AND U11442 ( .A(n11124), .B(n11123), .Z(n11162) );
  XOR U11443 ( .A(n11163), .B(n11162), .Z(c[1285]) );
  NANDN U11444 ( .A(n11126), .B(n11125), .Z(n11130) );
  NAND U11445 ( .A(n11128), .B(n11127), .Z(n11129) );
  NAND U11446 ( .A(n11130), .B(n11129), .Z(n11169) );
  NAND U11447 ( .A(b[0]), .B(a[270]), .Z(n11131) );
  XNOR U11448 ( .A(b[1]), .B(n11131), .Z(n11133) );
  NAND U11449 ( .A(n53), .B(a[269]), .Z(n11132) );
  AND U11450 ( .A(n11133), .B(n11132), .Z(n11186) );
  XOR U11451 ( .A(a[266]), .B(n42197), .Z(n11175) );
  NANDN U11452 ( .A(n11175), .B(n42173), .Z(n11136) );
  NANDN U11453 ( .A(n11134), .B(n42172), .Z(n11135) );
  NAND U11454 ( .A(n11136), .B(n11135), .Z(n11184) );
  NAND U11455 ( .A(b[7]), .B(a[262]), .Z(n11185) );
  XNOR U11456 ( .A(n11184), .B(n11185), .Z(n11187) );
  XOR U11457 ( .A(n11186), .B(n11187), .Z(n11193) );
  NANDN U11458 ( .A(n11137), .B(n42093), .Z(n11139) );
  XOR U11459 ( .A(n42134), .B(a[268]), .Z(n11178) );
  NANDN U11460 ( .A(n11178), .B(n42095), .Z(n11138) );
  NAND U11461 ( .A(n11139), .B(n11138), .Z(n11191) );
  NANDN U11462 ( .A(n11140), .B(n42231), .Z(n11142) );
  XOR U11463 ( .A(n184), .B(a[264]), .Z(n11181) );
  NANDN U11464 ( .A(n11181), .B(n42234), .Z(n11141) );
  AND U11465 ( .A(n11142), .B(n11141), .Z(n11190) );
  XNOR U11466 ( .A(n11191), .B(n11190), .Z(n11192) );
  XNOR U11467 ( .A(n11193), .B(n11192), .Z(n11197) );
  NANDN U11468 ( .A(n11144), .B(n11143), .Z(n11148) );
  NAND U11469 ( .A(n11146), .B(n11145), .Z(n11147) );
  AND U11470 ( .A(n11148), .B(n11147), .Z(n11196) );
  XOR U11471 ( .A(n11197), .B(n11196), .Z(n11198) );
  NANDN U11472 ( .A(n11150), .B(n11149), .Z(n11154) );
  NANDN U11473 ( .A(n11152), .B(n11151), .Z(n11153) );
  NAND U11474 ( .A(n11154), .B(n11153), .Z(n11199) );
  XOR U11475 ( .A(n11198), .B(n11199), .Z(n11166) );
  OR U11476 ( .A(n11156), .B(n11155), .Z(n11160) );
  NANDN U11477 ( .A(n11158), .B(n11157), .Z(n11159) );
  NAND U11478 ( .A(n11160), .B(n11159), .Z(n11167) );
  XNOR U11479 ( .A(n11166), .B(n11167), .Z(n11168) );
  XNOR U11480 ( .A(n11169), .B(n11168), .Z(n11202) );
  XNOR U11481 ( .A(n11202), .B(sreg[1286]), .Z(n11204) );
  NAND U11482 ( .A(n11161), .B(sreg[1285]), .Z(n11165) );
  OR U11483 ( .A(n11163), .B(n11162), .Z(n11164) );
  AND U11484 ( .A(n11165), .B(n11164), .Z(n11203) );
  XOR U11485 ( .A(n11204), .B(n11203), .Z(c[1286]) );
  NANDN U11486 ( .A(n11167), .B(n11166), .Z(n11171) );
  NAND U11487 ( .A(n11169), .B(n11168), .Z(n11170) );
  NAND U11488 ( .A(n11171), .B(n11170), .Z(n11210) );
  NAND U11489 ( .A(b[0]), .B(a[271]), .Z(n11172) );
  XNOR U11490 ( .A(b[1]), .B(n11172), .Z(n11174) );
  NAND U11491 ( .A(n53), .B(a[270]), .Z(n11173) );
  AND U11492 ( .A(n11174), .B(n11173), .Z(n11227) );
  XOR U11493 ( .A(a[267]), .B(n42197), .Z(n11216) );
  NANDN U11494 ( .A(n11216), .B(n42173), .Z(n11177) );
  NANDN U11495 ( .A(n11175), .B(n42172), .Z(n11176) );
  NAND U11496 ( .A(n11177), .B(n11176), .Z(n11225) );
  NAND U11497 ( .A(b[7]), .B(a[263]), .Z(n11226) );
  XNOR U11498 ( .A(n11225), .B(n11226), .Z(n11228) );
  XOR U11499 ( .A(n11227), .B(n11228), .Z(n11234) );
  NANDN U11500 ( .A(n11178), .B(n42093), .Z(n11180) );
  XOR U11501 ( .A(n42134), .B(a[269]), .Z(n11219) );
  NANDN U11502 ( .A(n11219), .B(n42095), .Z(n11179) );
  NAND U11503 ( .A(n11180), .B(n11179), .Z(n11232) );
  NANDN U11504 ( .A(n11181), .B(n42231), .Z(n11183) );
  XOR U11505 ( .A(n184), .B(a[265]), .Z(n11222) );
  NANDN U11506 ( .A(n11222), .B(n42234), .Z(n11182) );
  AND U11507 ( .A(n11183), .B(n11182), .Z(n11231) );
  XNOR U11508 ( .A(n11232), .B(n11231), .Z(n11233) );
  XNOR U11509 ( .A(n11234), .B(n11233), .Z(n11238) );
  NANDN U11510 ( .A(n11185), .B(n11184), .Z(n11189) );
  NAND U11511 ( .A(n11187), .B(n11186), .Z(n11188) );
  AND U11512 ( .A(n11189), .B(n11188), .Z(n11237) );
  XOR U11513 ( .A(n11238), .B(n11237), .Z(n11239) );
  NANDN U11514 ( .A(n11191), .B(n11190), .Z(n11195) );
  NANDN U11515 ( .A(n11193), .B(n11192), .Z(n11194) );
  NAND U11516 ( .A(n11195), .B(n11194), .Z(n11240) );
  XOR U11517 ( .A(n11239), .B(n11240), .Z(n11207) );
  OR U11518 ( .A(n11197), .B(n11196), .Z(n11201) );
  NANDN U11519 ( .A(n11199), .B(n11198), .Z(n11200) );
  NAND U11520 ( .A(n11201), .B(n11200), .Z(n11208) );
  XNOR U11521 ( .A(n11207), .B(n11208), .Z(n11209) );
  XNOR U11522 ( .A(n11210), .B(n11209), .Z(n11243) );
  XNOR U11523 ( .A(n11243), .B(sreg[1287]), .Z(n11245) );
  NAND U11524 ( .A(n11202), .B(sreg[1286]), .Z(n11206) );
  OR U11525 ( .A(n11204), .B(n11203), .Z(n11205) );
  AND U11526 ( .A(n11206), .B(n11205), .Z(n11244) );
  XOR U11527 ( .A(n11245), .B(n11244), .Z(c[1287]) );
  NANDN U11528 ( .A(n11208), .B(n11207), .Z(n11212) );
  NAND U11529 ( .A(n11210), .B(n11209), .Z(n11211) );
  NAND U11530 ( .A(n11212), .B(n11211), .Z(n11251) );
  NAND U11531 ( .A(b[0]), .B(a[272]), .Z(n11213) );
  XNOR U11532 ( .A(b[1]), .B(n11213), .Z(n11215) );
  NAND U11533 ( .A(n53), .B(a[271]), .Z(n11214) );
  AND U11534 ( .A(n11215), .B(n11214), .Z(n11268) );
  XOR U11535 ( .A(a[268]), .B(n42197), .Z(n11257) );
  NANDN U11536 ( .A(n11257), .B(n42173), .Z(n11218) );
  NANDN U11537 ( .A(n11216), .B(n42172), .Z(n11217) );
  NAND U11538 ( .A(n11218), .B(n11217), .Z(n11266) );
  NAND U11539 ( .A(b[7]), .B(a[264]), .Z(n11267) );
  XNOR U11540 ( .A(n11266), .B(n11267), .Z(n11269) );
  XOR U11541 ( .A(n11268), .B(n11269), .Z(n11275) );
  NANDN U11542 ( .A(n11219), .B(n42093), .Z(n11221) );
  XOR U11543 ( .A(n42134), .B(a[270]), .Z(n11260) );
  NANDN U11544 ( .A(n11260), .B(n42095), .Z(n11220) );
  NAND U11545 ( .A(n11221), .B(n11220), .Z(n11273) );
  NANDN U11546 ( .A(n11222), .B(n42231), .Z(n11224) );
  XOR U11547 ( .A(n184), .B(a[266]), .Z(n11263) );
  NANDN U11548 ( .A(n11263), .B(n42234), .Z(n11223) );
  AND U11549 ( .A(n11224), .B(n11223), .Z(n11272) );
  XNOR U11550 ( .A(n11273), .B(n11272), .Z(n11274) );
  XNOR U11551 ( .A(n11275), .B(n11274), .Z(n11279) );
  NANDN U11552 ( .A(n11226), .B(n11225), .Z(n11230) );
  NAND U11553 ( .A(n11228), .B(n11227), .Z(n11229) );
  AND U11554 ( .A(n11230), .B(n11229), .Z(n11278) );
  XOR U11555 ( .A(n11279), .B(n11278), .Z(n11280) );
  NANDN U11556 ( .A(n11232), .B(n11231), .Z(n11236) );
  NANDN U11557 ( .A(n11234), .B(n11233), .Z(n11235) );
  NAND U11558 ( .A(n11236), .B(n11235), .Z(n11281) );
  XOR U11559 ( .A(n11280), .B(n11281), .Z(n11248) );
  OR U11560 ( .A(n11238), .B(n11237), .Z(n11242) );
  NANDN U11561 ( .A(n11240), .B(n11239), .Z(n11241) );
  NAND U11562 ( .A(n11242), .B(n11241), .Z(n11249) );
  XNOR U11563 ( .A(n11248), .B(n11249), .Z(n11250) );
  XNOR U11564 ( .A(n11251), .B(n11250), .Z(n11284) );
  XNOR U11565 ( .A(n11284), .B(sreg[1288]), .Z(n11286) );
  NAND U11566 ( .A(n11243), .B(sreg[1287]), .Z(n11247) );
  OR U11567 ( .A(n11245), .B(n11244), .Z(n11246) );
  AND U11568 ( .A(n11247), .B(n11246), .Z(n11285) );
  XOR U11569 ( .A(n11286), .B(n11285), .Z(c[1288]) );
  NANDN U11570 ( .A(n11249), .B(n11248), .Z(n11253) );
  NAND U11571 ( .A(n11251), .B(n11250), .Z(n11252) );
  NAND U11572 ( .A(n11253), .B(n11252), .Z(n11292) );
  NAND U11573 ( .A(b[0]), .B(a[273]), .Z(n11254) );
  XNOR U11574 ( .A(b[1]), .B(n11254), .Z(n11256) );
  NAND U11575 ( .A(n54), .B(a[272]), .Z(n11255) );
  AND U11576 ( .A(n11256), .B(n11255), .Z(n11309) );
  XOR U11577 ( .A(a[269]), .B(n42197), .Z(n11298) );
  NANDN U11578 ( .A(n11298), .B(n42173), .Z(n11259) );
  NANDN U11579 ( .A(n11257), .B(n42172), .Z(n11258) );
  NAND U11580 ( .A(n11259), .B(n11258), .Z(n11307) );
  NAND U11581 ( .A(b[7]), .B(a[265]), .Z(n11308) );
  XNOR U11582 ( .A(n11307), .B(n11308), .Z(n11310) );
  XOR U11583 ( .A(n11309), .B(n11310), .Z(n11316) );
  NANDN U11584 ( .A(n11260), .B(n42093), .Z(n11262) );
  XOR U11585 ( .A(n42134), .B(a[271]), .Z(n11301) );
  NANDN U11586 ( .A(n11301), .B(n42095), .Z(n11261) );
  NAND U11587 ( .A(n11262), .B(n11261), .Z(n11314) );
  NANDN U11588 ( .A(n11263), .B(n42231), .Z(n11265) );
  XOR U11589 ( .A(n184), .B(a[267]), .Z(n11304) );
  NANDN U11590 ( .A(n11304), .B(n42234), .Z(n11264) );
  AND U11591 ( .A(n11265), .B(n11264), .Z(n11313) );
  XNOR U11592 ( .A(n11314), .B(n11313), .Z(n11315) );
  XNOR U11593 ( .A(n11316), .B(n11315), .Z(n11320) );
  NANDN U11594 ( .A(n11267), .B(n11266), .Z(n11271) );
  NAND U11595 ( .A(n11269), .B(n11268), .Z(n11270) );
  AND U11596 ( .A(n11271), .B(n11270), .Z(n11319) );
  XOR U11597 ( .A(n11320), .B(n11319), .Z(n11321) );
  NANDN U11598 ( .A(n11273), .B(n11272), .Z(n11277) );
  NANDN U11599 ( .A(n11275), .B(n11274), .Z(n11276) );
  NAND U11600 ( .A(n11277), .B(n11276), .Z(n11322) );
  XOR U11601 ( .A(n11321), .B(n11322), .Z(n11289) );
  OR U11602 ( .A(n11279), .B(n11278), .Z(n11283) );
  NANDN U11603 ( .A(n11281), .B(n11280), .Z(n11282) );
  NAND U11604 ( .A(n11283), .B(n11282), .Z(n11290) );
  XNOR U11605 ( .A(n11289), .B(n11290), .Z(n11291) );
  XNOR U11606 ( .A(n11292), .B(n11291), .Z(n11325) );
  XNOR U11607 ( .A(n11325), .B(sreg[1289]), .Z(n11327) );
  NAND U11608 ( .A(n11284), .B(sreg[1288]), .Z(n11288) );
  OR U11609 ( .A(n11286), .B(n11285), .Z(n11287) );
  AND U11610 ( .A(n11288), .B(n11287), .Z(n11326) );
  XOR U11611 ( .A(n11327), .B(n11326), .Z(c[1289]) );
  NANDN U11612 ( .A(n11290), .B(n11289), .Z(n11294) );
  NAND U11613 ( .A(n11292), .B(n11291), .Z(n11293) );
  NAND U11614 ( .A(n11294), .B(n11293), .Z(n11333) );
  NAND U11615 ( .A(b[0]), .B(a[274]), .Z(n11295) );
  XNOR U11616 ( .A(b[1]), .B(n11295), .Z(n11297) );
  NAND U11617 ( .A(n54), .B(a[273]), .Z(n11296) );
  AND U11618 ( .A(n11297), .B(n11296), .Z(n11350) );
  XOR U11619 ( .A(a[270]), .B(n42197), .Z(n11339) );
  NANDN U11620 ( .A(n11339), .B(n42173), .Z(n11300) );
  NANDN U11621 ( .A(n11298), .B(n42172), .Z(n11299) );
  NAND U11622 ( .A(n11300), .B(n11299), .Z(n11348) );
  NAND U11623 ( .A(b[7]), .B(a[266]), .Z(n11349) );
  XNOR U11624 ( .A(n11348), .B(n11349), .Z(n11351) );
  XOR U11625 ( .A(n11350), .B(n11351), .Z(n11357) );
  NANDN U11626 ( .A(n11301), .B(n42093), .Z(n11303) );
  XOR U11627 ( .A(n42134), .B(a[272]), .Z(n11342) );
  NANDN U11628 ( .A(n11342), .B(n42095), .Z(n11302) );
  NAND U11629 ( .A(n11303), .B(n11302), .Z(n11355) );
  NANDN U11630 ( .A(n11304), .B(n42231), .Z(n11306) );
  XOR U11631 ( .A(n184), .B(a[268]), .Z(n11345) );
  NANDN U11632 ( .A(n11345), .B(n42234), .Z(n11305) );
  AND U11633 ( .A(n11306), .B(n11305), .Z(n11354) );
  XNOR U11634 ( .A(n11355), .B(n11354), .Z(n11356) );
  XNOR U11635 ( .A(n11357), .B(n11356), .Z(n11361) );
  NANDN U11636 ( .A(n11308), .B(n11307), .Z(n11312) );
  NAND U11637 ( .A(n11310), .B(n11309), .Z(n11311) );
  AND U11638 ( .A(n11312), .B(n11311), .Z(n11360) );
  XOR U11639 ( .A(n11361), .B(n11360), .Z(n11362) );
  NANDN U11640 ( .A(n11314), .B(n11313), .Z(n11318) );
  NANDN U11641 ( .A(n11316), .B(n11315), .Z(n11317) );
  NAND U11642 ( .A(n11318), .B(n11317), .Z(n11363) );
  XOR U11643 ( .A(n11362), .B(n11363), .Z(n11330) );
  OR U11644 ( .A(n11320), .B(n11319), .Z(n11324) );
  NANDN U11645 ( .A(n11322), .B(n11321), .Z(n11323) );
  NAND U11646 ( .A(n11324), .B(n11323), .Z(n11331) );
  XNOR U11647 ( .A(n11330), .B(n11331), .Z(n11332) );
  XNOR U11648 ( .A(n11333), .B(n11332), .Z(n11366) );
  XNOR U11649 ( .A(n11366), .B(sreg[1290]), .Z(n11368) );
  NAND U11650 ( .A(n11325), .B(sreg[1289]), .Z(n11329) );
  OR U11651 ( .A(n11327), .B(n11326), .Z(n11328) );
  AND U11652 ( .A(n11329), .B(n11328), .Z(n11367) );
  XOR U11653 ( .A(n11368), .B(n11367), .Z(c[1290]) );
  NANDN U11654 ( .A(n11331), .B(n11330), .Z(n11335) );
  NAND U11655 ( .A(n11333), .B(n11332), .Z(n11334) );
  NAND U11656 ( .A(n11335), .B(n11334), .Z(n11374) );
  NAND U11657 ( .A(b[0]), .B(a[275]), .Z(n11336) );
  XNOR U11658 ( .A(b[1]), .B(n11336), .Z(n11338) );
  NAND U11659 ( .A(n54), .B(a[274]), .Z(n11337) );
  AND U11660 ( .A(n11338), .B(n11337), .Z(n11391) );
  XOR U11661 ( .A(a[271]), .B(n42197), .Z(n11380) );
  NANDN U11662 ( .A(n11380), .B(n42173), .Z(n11341) );
  NANDN U11663 ( .A(n11339), .B(n42172), .Z(n11340) );
  NAND U11664 ( .A(n11341), .B(n11340), .Z(n11389) );
  NAND U11665 ( .A(b[7]), .B(a[267]), .Z(n11390) );
  XNOR U11666 ( .A(n11389), .B(n11390), .Z(n11392) );
  XOR U11667 ( .A(n11391), .B(n11392), .Z(n11398) );
  NANDN U11668 ( .A(n11342), .B(n42093), .Z(n11344) );
  XOR U11669 ( .A(n42134), .B(a[273]), .Z(n11383) );
  NANDN U11670 ( .A(n11383), .B(n42095), .Z(n11343) );
  NAND U11671 ( .A(n11344), .B(n11343), .Z(n11396) );
  NANDN U11672 ( .A(n11345), .B(n42231), .Z(n11347) );
  XOR U11673 ( .A(n184), .B(a[269]), .Z(n11386) );
  NANDN U11674 ( .A(n11386), .B(n42234), .Z(n11346) );
  AND U11675 ( .A(n11347), .B(n11346), .Z(n11395) );
  XNOR U11676 ( .A(n11396), .B(n11395), .Z(n11397) );
  XNOR U11677 ( .A(n11398), .B(n11397), .Z(n11402) );
  NANDN U11678 ( .A(n11349), .B(n11348), .Z(n11353) );
  NAND U11679 ( .A(n11351), .B(n11350), .Z(n11352) );
  AND U11680 ( .A(n11353), .B(n11352), .Z(n11401) );
  XOR U11681 ( .A(n11402), .B(n11401), .Z(n11403) );
  NANDN U11682 ( .A(n11355), .B(n11354), .Z(n11359) );
  NANDN U11683 ( .A(n11357), .B(n11356), .Z(n11358) );
  NAND U11684 ( .A(n11359), .B(n11358), .Z(n11404) );
  XOR U11685 ( .A(n11403), .B(n11404), .Z(n11371) );
  OR U11686 ( .A(n11361), .B(n11360), .Z(n11365) );
  NANDN U11687 ( .A(n11363), .B(n11362), .Z(n11364) );
  NAND U11688 ( .A(n11365), .B(n11364), .Z(n11372) );
  XNOR U11689 ( .A(n11371), .B(n11372), .Z(n11373) );
  XNOR U11690 ( .A(n11374), .B(n11373), .Z(n11407) );
  XNOR U11691 ( .A(n11407), .B(sreg[1291]), .Z(n11409) );
  NAND U11692 ( .A(n11366), .B(sreg[1290]), .Z(n11370) );
  OR U11693 ( .A(n11368), .B(n11367), .Z(n11369) );
  AND U11694 ( .A(n11370), .B(n11369), .Z(n11408) );
  XOR U11695 ( .A(n11409), .B(n11408), .Z(c[1291]) );
  NANDN U11696 ( .A(n11372), .B(n11371), .Z(n11376) );
  NAND U11697 ( .A(n11374), .B(n11373), .Z(n11375) );
  NAND U11698 ( .A(n11376), .B(n11375), .Z(n11415) );
  NAND U11699 ( .A(b[0]), .B(a[276]), .Z(n11377) );
  XNOR U11700 ( .A(b[1]), .B(n11377), .Z(n11379) );
  NAND U11701 ( .A(n54), .B(a[275]), .Z(n11378) );
  AND U11702 ( .A(n11379), .B(n11378), .Z(n11432) );
  XOR U11703 ( .A(a[272]), .B(n42197), .Z(n11421) );
  NANDN U11704 ( .A(n11421), .B(n42173), .Z(n11382) );
  NANDN U11705 ( .A(n11380), .B(n42172), .Z(n11381) );
  NAND U11706 ( .A(n11382), .B(n11381), .Z(n11430) );
  NAND U11707 ( .A(b[7]), .B(a[268]), .Z(n11431) );
  XNOR U11708 ( .A(n11430), .B(n11431), .Z(n11433) );
  XOR U11709 ( .A(n11432), .B(n11433), .Z(n11439) );
  NANDN U11710 ( .A(n11383), .B(n42093), .Z(n11385) );
  XOR U11711 ( .A(n42134), .B(a[274]), .Z(n11424) );
  NANDN U11712 ( .A(n11424), .B(n42095), .Z(n11384) );
  NAND U11713 ( .A(n11385), .B(n11384), .Z(n11437) );
  NANDN U11714 ( .A(n11386), .B(n42231), .Z(n11388) );
  XOR U11715 ( .A(n184), .B(a[270]), .Z(n11427) );
  NANDN U11716 ( .A(n11427), .B(n42234), .Z(n11387) );
  AND U11717 ( .A(n11388), .B(n11387), .Z(n11436) );
  XNOR U11718 ( .A(n11437), .B(n11436), .Z(n11438) );
  XNOR U11719 ( .A(n11439), .B(n11438), .Z(n11443) );
  NANDN U11720 ( .A(n11390), .B(n11389), .Z(n11394) );
  NAND U11721 ( .A(n11392), .B(n11391), .Z(n11393) );
  AND U11722 ( .A(n11394), .B(n11393), .Z(n11442) );
  XOR U11723 ( .A(n11443), .B(n11442), .Z(n11444) );
  NANDN U11724 ( .A(n11396), .B(n11395), .Z(n11400) );
  NANDN U11725 ( .A(n11398), .B(n11397), .Z(n11399) );
  NAND U11726 ( .A(n11400), .B(n11399), .Z(n11445) );
  XOR U11727 ( .A(n11444), .B(n11445), .Z(n11412) );
  OR U11728 ( .A(n11402), .B(n11401), .Z(n11406) );
  NANDN U11729 ( .A(n11404), .B(n11403), .Z(n11405) );
  NAND U11730 ( .A(n11406), .B(n11405), .Z(n11413) );
  XNOR U11731 ( .A(n11412), .B(n11413), .Z(n11414) );
  XNOR U11732 ( .A(n11415), .B(n11414), .Z(n11448) );
  XNOR U11733 ( .A(n11448), .B(sreg[1292]), .Z(n11450) );
  NAND U11734 ( .A(n11407), .B(sreg[1291]), .Z(n11411) );
  OR U11735 ( .A(n11409), .B(n11408), .Z(n11410) );
  AND U11736 ( .A(n11411), .B(n11410), .Z(n11449) );
  XOR U11737 ( .A(n11450), .B(n11449), .Z(c[1292]) );
  NANDN U11738 ( .A(n11413), .B(n11412), .Z(n11417) );
  NAND U11739 ( .A(n11415), .B(n11414), .Z(n11416) );
  NAND U11740 ( .A(n11417), .B(n11416), .Z(n11456) );
  NAND U11741 ( .A(b[0]), .B(a[277]), .Z(n11418) );
  XNOR U11742 ( .A(b[1]), .B(n11418), .Z(n11420) );
  NAND U11743 ( .A(n54), .B(a[276]), .Z(n11419) );
  AND U11744 ( .A(n11420), .B(n11419), .Z(n11473) );
  XOR U11745 ( .A(a[273]), .B(n42197), .Z(n11462) );
  NANDN U11746 ( .A(n11462), .B(n42173), .Z(n11423) );
  NANDN U11747 ( .A(n11421), .B(n42172), .Z(n11422) );
  NAND U11748 ( .A(n11423), .B(n11422), .Z(n11471) );
  NAND U11749 ( .A(b[7]), .B(a[269]), .Z(n11472) );
  XNOR U11750 ( .A(n11471), .B(n11472), .Z(n11474) );
  XOR U11751 ( .A(n11473), .B(n11474), .Z(n11480) );
  NANDN U11752 ( .A(n11424), .B(n42093), .Z(n11426) );
  XOR U11753 ( .A(n42134), .B(a[275]), .Z(n11465) );
  NANDN U11754 ( .A(n11465), .B(n42095), .Z(n11425) );
  NAND U11755 ( .A(n11426), .B(n11425), .Z(n11478) );
  NANDN U11756 ( .A(n11427), .B(n42231), .Z(n11429) );
  XOR U11757 ( .A(n184), .B(a[271]), .Z(n11468) );
  NANDN U11758 ( .A(n11468), .B(n42234), .Z(n11428) );
  AND U11759 ( .A(n11429), .B(n11428), .Z(n11477) );
  XNOR U11760 ( .A(n11478), .B(n11477), .Z(n11479) );
  XNOR U11761 ( .A(n11480), .B(n11479), .Z(n11484) );
  NANDN U11762 ( .A(n11431), .B(n11430), .Z(n11435) );
  NAND U11763 ( .A(n11433), .B(n11432), .Z(n11434) );
  AND U11764 ( .A(n11435), .B(n11434), .Z(n11483) );
  XOR U11765 ( .A(n11484), .B(n11483), .Z(n11485) );
  NANDN U11766 ( .A(n11437), .B(n11436), .Z(n11441) );
  NANDN U11767 ( .A(n11439), .B(n11438), .Z(n11440) );
  NAND U11768 ( .A(n11441), .B(n11440), .Z(n11486) );
  XOR U11769 ( .A(n11485), .B(n11486), .Z(n11453) );
  OR U11770 ( .A(n11443), .B(n11442), .Z(n11447) );
  NANDN U11771 ( .A(n11445), .B(n11444), .Z(n11446) );
  NAND U11772 ( .A(n11447), .B(n11446), .Z(n11454) );
  XNOR U11773 ( .A(n11453), .B(n11454), .Z(n11455) );
  XNOR U11774 ( .A(n11456), .B(n11455), .Z(n11489) );
  XNOR U11775 ( .A(n11489), .B(sreg[1293]), .Z(n11491) );
  NAND U11776 ( .A(n11448), .B(sreg[1292]), .Z(n11452) );
  OR U11777 ( .A(n11450), .B(n11449), .Z(n11451) );
  AND U11778 ( .A(n11452), .B(n11451), .Z(n11490) );
  XOR U11779 ( .A(n11491), .B(n11490), .Z(c[1293]) );
  NANDN U11780 ( .A(n11454), .B(n11453), .Z(n11458) );
  NAND U11781 ( .A(n11456), .B(n11455), .Z(n11457) );
  NAND U11782 ( .A(n11458), .B(n11457), .Z(n11497) );
  NAND U11783 ( .A(b[0]), .B(a[278]), .Z(n11459) );
  XNOR U11784 ( .A(b[1]), .B(n11459), .Z(n11461) );
  NAND U11785 ( .A(n54), .B(a[277]), .Z(n11460) );
  AND U11786 ( .A(n11461), .B(n11460), .Z(n11514) );
  XOR U11787 ( .A(a[274]), .B(n42197), .Z(n11503) );
  NANDN U11788 ( .A(n11503), .B(n42173), .Z(n11464) );
  NANDN U11789 ( .A(n11462), .B(n42172), .Z(n11463) );
  NAND U11790 ( .A(n11464), .B(n11463), .Z(n11512) );
  NAND U11791 ( .A(b[7]), .B(a[270]), .Z(n11513) );
  XNOR U11792 ( .A(n11512), .B(n11513), .Z(n11515) );
  XOR U11793 ( .A(n11514), .B(n11515), .Z(n11521) );
  NANDN U11794 ( .A(n11465), .B(n42093), .Z(n11467) );
  XOR U11795 ( .A(n42134), .B(a[276]), .Z(n11506) );
  NANDN U11796 ( .A(n11506), .B(n42095), .Z(n11466) );
  NAND U11797 ( .A(n11467), .B(n11466), .Z(n11519) );
  NANDN U11798 ( .A(n11468), .B(n42231), .Z(n11470) );
  XOR U11799 ( .A(n184), .B(a[272]), .Z(n11509) );
  NANDN U11800 ( .A(n11509), .B(n42234), .Z(n11469) );
  AND U11801 ( .A(n11470), .B(n11469), .Z(n11518) );
  XNOR U11802 ( .A(n11519), .B(n11518), .Z(n11520) );
  XNOR U11803 ( .A(n11521), .B(n11520), .Z(n11525) );
  NANDN U11804 ( .A(n11472), .B(n11471), .Z(n11476) );
  NAND U11805 ( .A(n11474), .B(n11473), .Z(n11475) );
  AND U11806 ( .A(n11476), .B(n11475), .Z(n11524) );
  XOR U11807 ( .A(n11525), .B(n11524), .Z(n11526) );
  NANDN U11808 ( .A(n11478), .B(n11477), .Z(n11482) );
  NANDN U11809 ( .A(n11480), .B(n11479), .Z(n11481) );
  NAND U11810 ( .A(n11482), .B(n11481), .Z(n11527) );
  XOR U11811 ( .A(n11526), .B(n11527), .Z(n11494) );
  OR U11812 ( .A(n11484), .B(n11483), .Z(n11488) );
  NANDN U11813 ( .A(n11486), .B(n11485), .Z(n11487) );
  NAND U11814 ( .A(n11488), .B(n11487), .Z(n11495) );
  XNOR U11815 ( .A(n11494), .B(n11495), .Z(n11496) );
  XNOR U11816 ( .A(n11497), .B(n11496), .Z(n11530) );
  XNOR U11817 ( .A(n11530), .B(sreg[1294]), .Z(n11532) );
  NAND U11818 ( .A(n11489), .B(sreg[1293]), .Z(n11493) );
  OR U11819 ( .A(n11491), .B(n11490), .Z(n11492) );
  AND U11820 ( .A(n11493), .B(n11492), .Z(n11531) );
  XOR U11821 ( .A(n11532), .B(n11531), .Z(c[1294]) );
  NANDN U11822 ( .A(n11495), .B(n11494), .Z(n11499) );
  NAND U11823 ( .A(n11497), .B(n11496), .Z(n11498) );
  NAND U11824 ( .A(n11499), .B(n11498), .Z(n11538) );
  NAND U11825 ( .A(b[0]), .B(a[279]), .Z(n11500) );
  XNOR U11826 ( .A(b[1]), .B(n11500), .Z(n11502) );
  NAND U11827 ( .A(n54), .B(a[278]), .Z(n11501) );
  AND U11828 ( .A(n11502), .B(n11501), .Z(n11555) );
  XOR U11829 ( .A(a[275]), .B(n42197), .Z(n11544) );
  NANDN U11830 ( .A(n11544), .B(n42173), .Z(n11505) );
  NANDN U11831 ( .A(n11503), .B(n42172), .Z(n11504) );
  NAND U11832 ( .A(n11505), .B(n11504), .Z(n11553) );
  NAND U11833 ( .A(b[7]), .B(a[271]), .Z(n11554) );
  XNOR U11834 ( .A(n11553), .B(n11554), .Z(n11556) );
  XOR U11835 ( .A(n11555), .B(n11556), .Z(n11562) );
  NANDN U11836 ( .A(n11506), .B(n42093), .Z(n11508) );
  XOR U11837 ( .A(n42134), .B(a[277]), .Z(n11547) );
  NANDN U11838 ( .A(n11547), .B(n42095), .Z(n11507) );
  NAND U11839 ( .A(n11508), .B(n11507), .Z(n11560) );
  NANDN U11840 ( .A(n11509), .B(n42231), .Z(n11511) );
  XOR U11841 ( .A(n184), .B(a[273]), .Z(n11550) );
  NANDN U11842 ( .A(n11550), .B(n42234), .Z(n11510) );
  AND U11843 ( .A(n11511), .B(n11510), .Z(n11559) );
  XNOR U11844 ( .A(n11560), .B(n11559), .Z(n11561) );
  XNOR U11845 ( .A(n11562), .B(n11561), .Z(n11566) );
  NANDN U11846 ( .A(n11513), .B(n11512), .Z(n11517) );
  NAND U11847 ( .A(n11515), .B(n11514), .Z(n11516) );
  AND U11848 ( .A(n11517), .B(n11516), .Z(n11565) );
  XOR U11849 ( .A(n11566), .B(n11565), .Z(n11567) );
  NANDN U11850 ( .A(n11519), .B(n11518), .Z(n11523) );
  NANDN U11851 ( .A(n11521), .B(n11520), .Z(n11522) );
  NAND U11852 ( .A(n11523), .B(n11522), .Z(n11568) );
  XOR U11853 ( .A(n11567), .B(n11568), .Z(n11535) );
  OR U11854 ( .A(n11525), .B(n11524), .Z(n11529) );
  NANDN U11855 ( .A(n11527), .B(n11526), .Z(n11528) );
  NAND U11856 ( .A(n11529), .B(n11528), .Z(n11536) );
  XNOR U11857 ( .A(n11535), .B(n11536), .Z(n11537) );
  XNOR U11858 ( .A(n11538), .B(n11537), .Z(n11571) );
  XNOR U11859 ( .A(n11571), .B(sreg[1295]), .Z(n11573) );
  NAND U11860 ( .A(n11530), .B(sreg[1294]), .Z(n11534) );
  OR U11861 ( .A(n11532), .B(n11531), .Z(n11533) );
  AND U11862 ( .A(n11534), .B(n11533), .Z(n11572) );
  XOR U11863 ( .A(n11573), .B(n11572), .Z(c[1295]) );
  NANDN U11864 ( .A(n11536), .B(n11535), .Z(n11540) );
  NAND U11865 ( .A(n11538), .B(n11537), .Z(n11539) );
  NAND U11866 ( .A(n11540), .B(n11539), .Z(n11579) );
  NAND U11867 ( .A(b[0]), .B(a[280]), .Z(n11541) );
  XNOR U11868 ( .A(b[1]), .B(n11541), .Z(n11543) );
  NAND U11869 ( .A(n55), .B(a[279]), .Z(n11542) );
  AND U11870 ( .A(n11543), .B(n11542), .Z(n11596) );
  XOR U11871 ( .A(a[276]), .B(n42197), .Z(n11585) );
  NANDN U11872 ( .A(n11585), .B(n42173), .Z(n11546) );
  NANDN U11873 ( .A(n11544), .B(n42172), .Z(n11545) );
  NAND U11874 ( .A(n11546), .B(n11545), .Z(n11594) );
  NAND U11875 ( .A(b[7]), .B(a[272]), .Z(n11595) );
  XNOR U11876 ( .A(n11594), .B(n11595), .Z(n11597) );
  XOR U11877 ( .A(n11596), .B(n11597), .Z(n11603) );
  NANDN U11878 ( .A(n11547), .B(n42093), .Z(n11549) );
  XOR U11879 ( .A(n42134), .B(a[278]), .Z(n11588) );
  NANDN U11880 ( .A(n11588), .B(n42095), .Z(n11548) );
  NAND U11881 ( .A(n11549), .B(n11548), .Z(n11601) );
  NANDN U11882 ( .A(n11550), .B(n42231), .Z(n11552) );
  XOR U11883 ( .A(n184), .B(a[274]), .Z(n11591) );
  NANDN U11884 ( .A(n11591), .B(n42234), .Z(n11551) );
  AND U11885 ( .A(n11552), .B(n11551), .Z(n11600) );
  XNOR U11886 ( .A(n11601), .B(n11600), .Z(n11602) );
  XNOR U11887 ( .A(n11603), .B(n11602), .Z(n11607) );
  NANDN U11888 ( .A(n11554), .B(n11553), .Z(n11558) );
  NAND U11889 ( .A(n11556), .B(n11555), .Z(n11557) );
  AND U11890 ( .A(n11558), .B(n11557), .Z(n11606) );
  XOR U11891 ( .A(n11607), .B(n11606), .Z(n11608) );
  NANDN U11892 ( .A(n11560), .B(n11559), .Z(n11564) );
  NANDN U11893 ( .A(n11562), .B(n11561), .Z(n11563) );
  NAND U11894 ( .A(n11564), .B(n11563), .Z(n11609) );
  XOR U11895 ( .A(n11608), .B(n11609), .Z(n11576) );
  OR U11896 ( .A(n11566), .B(n11565), .Z(n11570) );
  NANDN U11897 ( .A(n11568), .B(n11567), .Z(n11569) );
  NAND U11898 ( .A(n11570), .B(n11569), .Z(n11577) );
  XNOR U11899 ( .A(n11576), .B(n11577), .Z(n11578) );
  XNOR U11900 ( .A(n11579), .B(n11578), .Z(n11612) );
  XNOR U11901 ( .A(n11612), .B(sreg[1296]), .Z(n11614) );
  NAND U11902 ( .A(n11571), .B(sreg[1295]), .Z(n11575) );
  OR U11903 ( .A(n11573), .B(n11572), .Z(n11574) );
  AND U11904 ( .A(n11575), .B(n11574), .Z(n11613) );
  XOR U11905 ( .A(n11614), .B(n11613), .Z(c[1296]) );
  NANDN U11906 ( .A(n11577), .B(n11576), .Z(n11581) );
  NAND U11907 ( .A(n11579), .B(n11578), .Z(n11580) );
  NAND U11908 ( .A(n11581), .B(n11580), .Z(n11620) );
  NAND U11909 ( .A(b[0]), .B(a[281]), .Z(n11582) );
  XNOR U11910 ( .A(b[1]), .B(n11582), .Z(n11584) );
  NAND U11911 ( .A(n55), .B(a[280]), .Z(n11583) );
  AND U11912 ( .A(n11584), .B(n11583), .Z(n11637) );
  XOR U11913 ( .A(a[277]), .B(n42197), .Z(n11626) );
  NANDN U11914 ( .A(n11626), .B(n42173), .Z(n11587) );
  NANDN U11915 ( .A(n11585), .B(n42172), .Z(n11586) );
  NAND U11916 ( .A(n11587), .B(n11586), .Z(n11635) );
  NAND U11917 ( .A(b[7]), .B(a[273]), .Z(n11636) );
  XNOR U11918 ( .A(n11635), .B(n11636), .Z(n11638) );
  XOR U11919 ( .A(n11637), .B(n11638), .Z(n11644) );
  NANDN U11920 ( .A(n11588), .B(n42093), .Z(n11590) );
  XOR U11921 ( .A(n42134), .B(a[279]), .Z(n11629) );
  NANDN U11922 ( .A(n11629), .B(n42095), .Z(n11589) );
  NAND U11923 ( .A(n11590), .B(n11589), .Z(n11642) );
  NANDN U11924 ( .A(n11591), .B(n42231), .Z(n11593) );
  XOR U11925 ( .A(n185), .B(a[275]), .Z(n11632) );
  NANDN U11926 ( .A(n11632), .B(n42234), .Z(n11592) );
  AND U11927 ( .A(n11593), .B(n11592), .Z(n11641) );
  XNOR U11928 ( .A(n11642), .B(n11641), .Z(n11643) );
  XNOR U11929 ( .A(n11644), .B(n11643), .Z(n11648) );
  NANDN U11930 ( .A(n11595), .B(n11594), .Z(n11599) );
  NAND U11931 ( .A(n11597), .B(n11596), .Z(n11598) );
  AND U11932 ( .A(n11599), .B(n11598), .Z(n11647) );
  XOR U11933 ( .A(n11648), .B(n11647), .Z(n11649) );
  NANDN U11934 ( .A(n11601), .B(n11600), .Z(n11605) );
  NANDN U11935 ( .A(n11603), .B(n11602), .Z(n11604) );
  NAND U11936 ( .A(n11605), .B(n11604), .Z(n11650) );
  XOR U11937 ( .A(n11649), .B(n11650), .Z(n11617) );
  OR U11938 ( .A(n11607), .B(n11606), .Z(n11611) );
  NANDN U11939 ( .A(n11609), .B(n11608), .Z(n11610) );
  NAND U11940 ( .A(n11611), .B(n11610), .Z(n11618) );
  XNOR U11941 ( .A(n11617), .B(n11618), .Z(n11619) );
  XNOR U11942 ( .A(n11620), .B(n11619), .Z(n11653) );
  XNOR U11943 ( .A(n11653), .B(sreg[1297]), .Z(n11655) );
  NAND U11944 ( .A(n11612), .B(sreg[1296]), .Z(n11616) );
  OR U11945 ( .A(n11614), .B(n11613), .Z(n11615) );
  AND U11946 ( .A(n11616), .B(n11615), .Z(n11654) );
  XOR U11947 ( .A(n11655), .B(n11654), .Z(c[1297]) );
  NANDN U11948 ( .A(n11618), .B(n11617), .Z(n11622) );
  NAND U11949 ( .A(n11620), .B(n11619), .Z(n11621) );
  NAND U11950 ( .A(n11622), .B(n11621), .Z(n11661) );
  NAND U11951 ( .A(b[0]), .B(a[282]), .Z(n11623) );
  XNOR U11952 ( .A(b[1]), .B(n11623), .Z(n11625) );
  NAND U11953 ( .A(n55), .B(a[281]), .Z(n11624) );
  AND U11954 ( .A(n11625), .B(n11624), .Z(n11678) );
  XOR U11955 ( .A(a[278]), .B(n42197), .Z(n11667) );
  NANDN U11956 ( .A(n11667), .B(n42173), .Z(n11628) );
  NANDN U11957 ( .A(n11626), .B(n42172), .Z(n11627) );
  NAND U11958 ( .A(n11628), .B(n11627), .Z(n11676) );
  NAND U11959 ( .A(b[7]), .B(a[274]), .Z(n11677) );
  XNOR U11960 ( .A(n11676), .B(n11677), .Z(n11679) );
  XOR U11961 ( .A(n11678), .B(n11679), .Z(n11685) );
  NANDN U11962 ( .A(n11629), .B(n42093), .Z(n11631) );
  XOR U11963 ( .A(n42134), .B(a[280]), .Z(n11670) );
  NANDN U11964 ( .A(n11670), .B(n42095), .Z(n11630) );
  NAND U11965 ( .A(n11631), .B(n11630), .Z(n11683) );
  NANDN U11966 ( .A(n11632), .B(n42231), .Z(n11634) );
  XOR U11967 ( .A(n185), .B(a[276]), .Z(n11673) );
  NANDN U11968 ( .A(n11673), .B(n42234), .Z(n11633) );
  AND U11969 ( .A(n11634), .B(n11633), .Z(n11682) );
  XNOR U11970 ( .A(n11683), .B(n11682), .Z(n11684) );
  XNOR U11971 ( .A(n11685), .B(n11684), .Z(n11689) );
  NANDN U11972 ( .A(n11636), .B(n11635), .Z(n11640) );
  NAND U11973 ( .A(n11638), .B(n11637), .Z(n11639) );
  AND U11974 ( .A(n11640), .B(n11639), .Z(n11688) );
  XOR U11975 ( .A(n11689), .B(n11688), .Z(n11690) );
  NANDN U11976 ( .A(n11642), .B(n11641), .Z(n11646) );
  NANDN U11977 ( .A(n11644), .B(n11643), .Z(n11645) );
  NAND U11978 ( .A(n11646), .B(n11645), .Z(n11691) );
  XOR U11979 ( .A(n11690), .B(n11691), .Z(n11658) );
  OR U11980 ( .A(n11648), .B(n11647), .Z(n11652) );
  NANDN U11981 ( .A(n11650), .B(n11649), .Z(n11651) );
  NAND U11982 ( .A(n11652), .B(n11651), .Z(n11659) );
  XNOR U11983 ( .A(n11658), .B(n11659), .Z(n11660) );
  XNOR U11984 ( .A(n11661), .B(n11660), .Z(n11694) );
  XNOR U11985 ( .A(n11694), .B(sreg[1298]), .Z(n11696) );
  NAND U11986 ( .A(n11653), .B(sreg[1297]), .Z(n11657) );
  OR U11987 ( .A(n11655), .B(n11654), .Z(n11656) );
  AND U11988 ( .A(n11657), .B(n11656), .Z(n11695) );
  XOR U11989 ( .A(n11696), .B(n11695), .Z(c[1298]) );
  NANDN U11990 ( .A(n11659), .B(n11658), .Z(n11663) );
  NAND U11991 ( .A(n11661), .B(n11660), .Z(n11662) );
  NAND U11992 ( .A(n11663), .B(n11662), .Z(n11702) );
  NAND U11993 ( .A(b[0]), .B(a[283]), .Z(n11664) );
  XNOR U11994 ( .A(b[1]), .B(n11664), .Z(n11666) );
  NAND U11995 ( .A(n55), .B(a[282]), .Z(n11665) );
  AND U11996 ( .A(n11666), .B(n11665), .Z(n11719) );
  XOR U11997 ( .A(a[279]), .B(n42197), .Z(n11708) );
  NANDN U11998 ( .A(n11708), .B(n42173), .Z(n11669) );
  NANDN U11999 ( .A(n11667), .B(n42172), .Z(n11668) );
  NAND U12000 ( .A(n11669), .B(n11668), .Z(n11717) );
  NAND U12001 ( .A(b[7]), .B(a[275]), .Z(n11718) );
  XNOR U12002 ( .A(n11717), .B(n11718), .Z(n11720) );
  XOR U12003 ( .A(n11719), .B(n11720), .Z(n11726) );
  NANDN U12004 ( .A(n11670), .B(n42093), .Z(n11672) );
  XOR U12005 ( .A(n42134), .B(a[281]), .Z(n11711) );
  NANDN U12006 ( .A(n11711), .B(n42095), .Z(n11671) );
  NAND U12007 ( .A(n11672), .B(n11671), .Z(n11724) );
  NANDN U12008 ( .A(n11673), .B(n42231), .Z(n11675) );
  XOR U12009 ( .A(n185), .B(a[277]), .Z(n11714) );
  NANDN U12010 ( .A(n11714), .B(n42234), .Z(n11674) );
  AND U12011 ( .A(n11675), .B(n11674), .Z(n11723) );
  XNOR U12012 ( .A(n11724), .B(n11723), .Z(n11725) );
  XNOR U12013 ( .A(n11726), .B(n11725), .Z(n11730) );
  NANDN U12014 ( .A(n11677), .B(n11676), .Z(n11681) );
  NAND U12015 ( .A(n11679), .B(n11678), .Z(n11680) );
  AND U12016 ( .A(n11681), .B(n11680), .Z(n11729) );
  XOR U12017 ( .A(n11730), .B(n11729), .Z(n11731) );
  NANDN U12018 ( .A(n11683), .B(n11682), .Z(n11687) );
  NANDN U12019 ( .A(n11685), .B(n11684), .Z(n11686) );
  NAND U12020 ( .A(n11687), .B(n11686), .Z(n11732) );
  XOR U12021 ( .A(n11731), .B(n11732), .Z(n11699) );
  OR U12022 ( .A(n11689), .B(n11688), .Z(n11693) );
  NANDN U12023 ( .A(n11691), .B(n11690), .Z(n11692) );
  NAND U12024 ( .A(n11693), .B(n11692), .Z(n11700) );
  XNOR U12025 ( .A(n11699), .B(n11700), .Z(n11701) );
  XNOR U12026 ( .A(n11702), .B(n11701), .Z(n11735) );
  XNOR U12027 ( .A(n11735), .B(sreg[1299]), .Z(n11737) );
  NAND U12028 ( .A(n11694), .B(sreg[1298]), .Z(n11698) );
  OR U12029 ( .A(n11696), .B(n11695), .Z(n11697) );
  AND U12030 ( .A(n11698), .B(n11697), .Z(n11736) );
  XOR U12031 ( .A(n11737), .B(n11736), .Z(c[1299]) );
  NANDN U12032 ( .A(n11700), .B(n11699), .Z(n11704) );
  NAND U12033 ( .A(n11702), .B(n11701), .Z(n11703) );
  NAND U12034 ( .A(n11704), .B(n11703), .Z(n11743) );
  NAND U12035 ( .A(b[0]), .B(a[284]), .Z(n11705) );
  XNOR U12036 ( .A(b[1]), .B(n11705), .Z(n11707) );
  NAND U12037 ( .A(n55), .B(a[283]), .Z(n11706) );
  AND U12038 ( .A(n11707), .B(n11706), .Z(n11760) );
  XOR U12039 ( .A(a[280]), .B(n42197), .Z(n11749) );
  NANDN U12040 ( .A(n11749), .B(n42173), .Z(n11710) );
  NANDN U12041 ( .A(n11708), .B(n42172), .Z(n11709) );
  NAND U12042 ( .A(n11710), .B(n11709), .Z(n11758) );
  NAND U12043 ( .A(b[7]), .B(a[276]), .Z(n11759) );
  XNOR U12044 ( .A(n11758), .B(n11759), .Z(n11761) );
  XOR U12045 ( .A(n11760), .B(n11761), .Z(n11767) );
  NANDN U12046 ( .A(n11711), .B(n42093), .Z(n11713) );
  XOR U12047 ( .A(n42134), .B(a[282]), .Z(n11752) );
  NANDN U12048 ( .A(n11752), .B(n42095), .Z(n11712) );
  NAND U12049 ( .A(n11713), .B(n11712), .Z(n11765) );
  NANDN U12050 ( .A(n11714), .B(n42231), .Z(n11716) );
  XOR U12051 ( .A(n185), .B(a[278]), .Z(n11755) );
  NANDN U12052 ( .A(n11755), .B(n42234), .Z(n11715) );
  AND U12053 ( .A(n11716), .B(n11715), .Z(n11764) );
  XNOR U12054 ( .A(n11765), .B(n11764), .Z(n11766) );
  XNOR U12055 ( .A(n11767), .B(n11766), .Z(n11771) );
  NANDN U12056 ( .A(n11718), .B(n11717), .Z(n11722) );
  NAND U12057 ( .A(n11720), .B(n11719), .Z(n11721) );
  AND U12058 ( .A(n11722), .B(n11721), .Z(n11770) );
  XOR U12059 ( .A(n11771), .B(n11770), .Z(n11772) );
  NANDN U12060 ( .A(n11724), .B(n11723), .Z(n11728) );
  NANDN U12061 ( .A(n11726), .B(n11725), .Z(n11727) );
  NAND U12062 ( .A(n11728), .B(n11727), .Z(n11773) );
  XOR U12063 ( .A(n11772), .B(n11773), .Z(n11740) );
  OR U12064 ( .A(n11730), .B(n11729), .Z(n11734) );
  NANDN U12065 ( .A(n11732), .B(n11731), .Z(n11733) );
  NAND U12066 ( .A(n11734), .B(n11733), .Z(n11741) );
  XNOR U12067 ( .A(n11740), .B(n11741), .Z(n11742) );
  XNOR U12068 ( .A(n11743), .B(n11742), .Z(n11776) );
  XNOR U12069 ( .A(n11776), .B(sreg[1300]), .Z(n11778) );
  NAND U12070 ( .A(n11735), .B(sreg[1299]), .Z(n11739) );
  OR U12071 ( .A(n11737), .B(n11736), .Z(n11738) );
  AND U12072 ( .A(n11739), .B(n11738), .Z(n11777) );
  XOR U12073 ( .A(n11778), .B(n11777), .Z(c[1300]) );
  NANDN U12074 ( .A(n11741), .B(n11740), .Z(n11745) );
  NAND U12075 ( .A(n11743), .B(n11742), .Z(n11744) );
  NAND U12076 ( .A(n11745), .B(n11744), .Z(n11784) );
  NAND U12077 ( .A(b[0]), .B(a[285]), .Z(n11746) );
  XNOR U12078 ( .A(b[1]), .B(n11746), .Z(n11748) );
  NAND U12079 ( .A(n55), .B(a[284]), .Z(n11747) );
  AND U12080 ( .A(n11748), .B(n11747), .Z(n11801) );
  XOR U12081 ( .A(a[281]), .B(n42197), .Z(n11790) );
  NANDN U12082 ( .A(n11790), .B(n42173), .Z(n11751) );
  NANDN U12083 ( .A(n11749), .B(n42172), .Z(n11750) );
  NAND U12084 ( .A(n11751), .B(n11750), .Z(n11799) );
  NAND U12085 ( .A(b[7]), .B(a[277]), .Z(n11800) );
  XNOR U12086 ( .A(n11799), .B(n11800), .Z(n11802) );
  XOR U12087 ( .A(n11801), .B(n11802), .Z(n11808) );
  NANDN U12088 ( .A(n11752), .B(n42093), .Z(n11754) );
  XOR U12089 ( .A(n42134), .B(a[283]), .Z(n11793) );
  NANDN U12090 ( .A(n11793), .B(n42095), .Z(n11753) );
  NAND U12091 ( .A(n11754), .B(n11753), .Z(n11806) );
  NANDN U12092 ( .A(n11755), .B(n42231), .Z(n11757) );
  XOR U12093 ( .A(n185), .B(a[279]), .Z(n11796) );
  NANDN U12094 ( .A(n11796), .B(n42234), .Z(n11756) );
  AND U12095 ( .A(n11757), .B(n11756), .Z(n11805) );
  XNOR U12096 ( .A(n11806), .B(n11805), .Z(n11807) );
  XNOR U12097 ( .A(n11808), .B(n11807), .Z(n11812) );
  NANDN U12098 ( .A(n11759), .B(n11758), .Z(n11763) );
  NAND U12099 ( .A(n11761), .B(n11760), .Z(n11762) );
  AND U12100 ( .A(n11763), .B(n11762), .Z(n11811) );
  XOR U12101 ( .A(n11812), .B(n11811), .Z(n11813) );
  NANDN U12102 ( .A(n11765), .B(n11764), .Z(n11769) );
  NANDN U12103 ( .A(n11767), .B(n11766), .Z(n11768) );
  NAND U12104 ( .A(n11769), .B(n11768), .Z(n11814) );
  XOR U12105 ( .A(n11813), .B(n11814), .Z(n11781) );
  OR U12106 ( .A(n11771), .B(n11770), .Z(n11775) );
  NANDN U12107 ( .A(n11773), .B(n11772), .Z(n11774) );
  NAND U12108 ( .A(n11775), .B(n11774), .Z(n11782) );
  XNOR U12109 ( .A(n11781), .B(n11782), .Z(n11783) );
  XNOR U12110 ( .A(n11784), .B(n11783), .Z(n11817) );
  XNOR U12111 ( .A(n11817), .B(sreg[1301]), .Z(n11819) );
  NAND U12112 ( .A(n11776), .B(sreg[1300]), .Z(n11780) );
  OR U12113 ( .A(n11778), .B(n11777), .Z(n11779) );
  AND U12114 ( .A(n11780), .B(n11779), .Z(n11818) );
  XOR U12115 ( .A(n11819), .B(n11818), .Z(c[1301]) );
  NANDN U12116 ( .A(n11782), .B(n11781), .Z(n11786) );
  NAND U12117 ( .A(n11784), .B(n11783), .Z(n11785) );
  NAND U12118 ( .A(n11786), .B(n11785), .Z(n11825) );
  NAND U12119 ( .A(b[0]), .B(a[286]), .Z(n11787) );
  XNOR U12120 ( .A(b[1]), .B(n11787), .Z(n11789) );
  NAND U12121 ( .A(n55), .B(a[285]), .Z(n11788) );
  AND U12122 ( .A(n11789), .B(n11788), .Z(n11842) );
  XOR U12123 ( .A(a[282]), .B(n42197), .Z(n11831) );
  NANDN U12124 ( .A(n11831), .B(n42173), .Z(n11792) );
  NANDN U12125 ( .A(n11790), .B(n42172), .Z(n11791) );
  NAND U12126 ( .A(n11792), .B(n11791), .Z(n11840) );
  NAND U12127 ( .A(b[7]), .B(a[278]), .Z(n11841) );
  XNOR U12128 ( .A(n11840), .B(n11841), .Z(n11843) );
  XOR U12129 ( .A(n11842), .B(n11843), .Z(n11849) );
  NANDN U12130 ( .A(n11793), .B(n42093), .Z(n11795) );
  XOR U12131 ( .A(n42134), .B(a[284]), .Z(n11834) );
  NANDN U12132 ( .A(n11834), .B(n42095), .Z(n11794) );
  NAND U12133 ( .A(n11795), .B(n11794), .Z(n11847) );
  NANDN U12134 ( .A(n11796), .B(n42231), .Z(n11798) );
  XOR U12135 ( .A(n185), .B(a[280]), .Z(n11837) );
  NANDN U12136 ( .A(n11837), .B(n42234), .Z(n11797) );
  AND U12137 ( .A(n11798), .B(n11797), .Z(n11846) );
  XNOR U12138 ( .A(n11847), .B(n11846), .Z(n11848) );
  XNOR U12139 ( .A(n11849), .B(n11848), .Z(n11853) );
  NANDN U12140 ( .A(n11800), .B(n11799), .Z(n11804) );
  NAND U12141 ( .A(n11802), .B(n11801), .Z(n11803) );
  AND U12142 ( .A(n11804), .B(n11803), .Z(n11852) );
  XOR U12143 ( .A(n11853), .B(n11852), .Z(n11854) );
  NANDN U12144 ( .A(n11806), .B(n11805), .Z(n11810) );
  NANDN U12145 ( .A(n11808), .B(n11807), .Z(n11809) );
  NAND U12146 ( .A(n11810), .B(n11809), .Z(n11855) );
  XOR U12147 ( .A(n11854), .B(n11855), .Z(n11822) );
  OR U12148 ( .A(n11812), .B(n11811), .Z(n11816) );
  NANDN U12149 ( .A(n11814), .B(n11813), .Z(n11815) );
  NAND U12150 ( .A(n11816), .B(n11815), .Z(n11823) );
  XNOR U12151 ( .A(n11822), .B(n11823), .Z(n11824) );
  XNOR U12152 ( .A(n11825), .B(n11824), .Z(n11858) );
  XNOR U12153 ( .A(n11858), .B(sreg[1302]), .Z(n11860) );
  NAND U12154 ( .A(n11817), .B(sreg[1301]), .Z(n11821) );
  OR U12155 ( .A(n11819), .B(n11818), .Z(n11820) );
  AND U12156 ( .A(n11821), .B(n11820), .Z(n11859) );
  XOR U12157 ( .A(n11860), .B(n11859), .Z(c[1302]) );
  NANDN U12158 ( .A(n11823), .B(n11822), .Z(n11827) );
  NAND U12159 ( .A(n11825), .B(n11824), .Z(n11826) );
  NAND U12160 ( .A(n11827), .B(n11826), .Z(n11866) );
  NAND U12161 ( .A(b[0]), .B(a[287]), .Z(n11828) );
  XNOR U12162 ( .A(b[1]), .B(n11828), .Z(n11830) );
  NAND U12163 ( .A(n56), .B(a[286]), .Z(n11829) );
  AND U12164 ( .A(n11830), .B(n11829), .Z(n11883) );
  XOR U12165 ( .A(a[283]), .B(n42197), .Z(n11872) );
  NANDN U12166 ( .A(n11872), .B(n42173), .Z(n11833) );
  NANDN U12167 ( .A(n11831), .B(n42172), .Z(n11832) );
  NAND U12168 ( .A(n11833), .B(n11832), .Z(n11881) );
  NAND U12169 ( .A(b[7]), .B(a[279]), .Z(n11882) );
  XNOR U12170 ( .A(n11881), .B(n11882), .Z(n11884) );
  XOR U12171 ( .A(n11883), .B(n11884), .Z(n11890) );
  NANDN U12172 ( .A(n11834), .B(n42093), .Z(n11836) );
  XOR U12173 ( .A(n42134), .B(a[285]), .Z(n11875) );
  NANDN U12174 ( .A(n11875), .B(n42095), .Z(n11835) );
  NAND U12175 ( .A(n11836), .B(n11835), .Z(n11888) );
  NANDN U12176 ( .A(n11837), .B(n42231), .Z(n11839) );
  XOR U12177 ( .A(n185), .B(a[281]), .Z(n11878) );
  NANDN U12178 ( .A(n11878), .B(n42234), .Z(n11838) );
  AND U12179 ( .A(n11839), .B(n11838), .Z(n11887) );
  XNOR U12180 ( .A(n11888), .B(n11887), .Z(n11889) );
  XNOR U12181 ( .A(n11890), .B(n11889), .Z(n11894) );
  NANDN U12182 ( .A(n11841), .B(n11840), .Z(n11845) );
  NAND U12183 ( .A(n11843), .B(n11842), .Z(n11844) );
  AND U12184 ( .A(n11845), .B(n11844), .Z(n11893) );
  XOR U12185 ( .A(n11894), .B(n11893), .Z(n11895) );
  NANDN U12186 ( .A(n11847), .B(n11846), .Z(n11851) );
  NANDN U12187 ( .A(n11849), .B(n11848), .Z(n11850) );
  NAND U12188 ( .A(n11851), .B(n11850), .Z(n11896) );
  XOR U12189 ( .A(n11895), .B(n11896), .Z(n11863) );
  OR U12190 ( .A(n11853), .B(n11852), .Z(n11857) );
  NANDN U12191 ( .A(n11855), .B(n11854), .Z(n11856) );
  NAND U12192 ( .A(n11857), .B(n11856), .Z(n11864) );
  XNOR U12193 ( .A(n11863), .B(n11864), .Z(n11865) );
  XNOR U12194 ( .A(n11866), .B(n11865), .Z(n11899) );
  XNOR U12195 ( .A(n11899), .B(sreg[1303]), .Z(n11901) );
  NAND U12196 ( .A(n11858), .B(sreg[1302]), .Z(n11862) );
  OR U12197 ( .A(n11860), .B(n11859), .Z(n11861) );
  AND U12198 ( .A(n11862), .B(n11861), .Z(n11900) );
  XOR U12199 ( .A(n11901), .B(n11900), .Z(c[1303]) );
  NANDN U12200 ( .A(n11864), .B(n11863), .Z(n11868) );
  NAND U12201 ( .A(n11866), .B(n11865), .Z(n11867) );
  NAND U12202 ( .A(n11868), .B(n11867), .Z(n11907) );
  NAND U12203 ( .A(b[0]), .B(a[288]), .Z(n11869) );
  XNOR U12204 ( .A(b[1]), .B(n11869), .Z(n11871) );
  NAND U12205 ( .A(n56), .B(a[287]), .Z(n11870) );
  AND U12206 ( .A(n11871), .B(n11870), .Z(n11924) );
  XOR U12207 ( .A(a[284]), .B(n42197), .Z(n11913) );
  NANDN U12208 ( .A(n11913), .B(n42173), .Z(n11874) );
  NANDN U12209 ( .A(n11872), .B(n42172), .Z(n11873) );
  NAND U12210 ( .A(n11874), .B(n11873), .Z(n11922) );
  NAND U12211 ( .A(b[7]), .B(a[280]), .Z(n11923) );
  XNOR U12212 ( .A(n11922), .B(n11923), .Z(n11925) );
  XOR U12213 ( .A(n11924), .B(n11925), .Z(n11931) );
  NANDN U12214 ( .A(n11875), .B(n42093), .Z(n11877) );
  XOR U12215 ( .A(n42134), .B(a[286]), .Z(n11916) );
  NANDN U12216 ( .A(n11916), .B(n42095), .Z(n11876) );
  NAND U12217 ( .A(n11877), .B(n11876), .Z(n11929) );
  NANDN U12218 ( .A(n11878), .B(n42231), .Z(n11880) );
  XOR U12219 ( .A(n185), .B(a[282]), .Z(n11919) );
  NANDN U12220 ( .A(n11919), .B(n42234), .Z(n11879) );
  AND U12221 ( .A(n11880), .B(n11879), .Z(n11928) );
  XNOR U12222 ( .A(n11929), .B(n11928), .Z(n11930) );
  XNOR U12223 ( .A(n11931), .B(n11930), .Z(n11935) );
  NANDN U12224 ( .A(n11882), .B(n11881), .Z(n11886) );
  NAND U12225 ( .A(n11884), .B(n11883), .Z(n11885) );
  AND U12226 ( .A(n11886), .B(n11885), .Z(n11934) );
  XOR U12227 ( .A(n11935), .B(n11934), .Z(n11936) );
  NANDN U12228 ( .A(n11888), .B(n11887), .Z(n11892) );
  NANDN U12229 ( .A(n11890), .B(n11889), .Z(n11891) );
  NAND U12230 ( .A(n11892), .B(n11891), .Z(n11937) );
  XOR U12231 ( .A(n11936), .B(n11937), .Z(n11904) );
  OR U12232 ( .A(n11894), .B(n11893), .Z(n11898) );
  NANDN U12233 ( .A(n11896), .B(n11895), .Z(n11897) );
  NAND U12234 ( .A(n11898), .B(n11897), .Z(n11905) );
  XNOR U12235 ( .A(n11904), .B(n11905), .Z(n11906) );
  XNOR U12236 ( .A(n11907), .B(n11906), .Z(n11940) );
  XNOR U12237 ( .A(n11940), .B(sreg[1304]), .Z(n11942) );
  NAND U12238 ( .A(n11899), .B(sreg[1303]), .Z(n11903) );
  OR U12239 ( .A(n11901), .B(n11900), .Z(n11902) );
  AND U12240 ( .A(n11903), .B(n11902), .Z(n11941) );
  XOR U12241 ( .A(n11942), .B(n11941), .Z(c[1304]) );
  NANDN U12242 ( .A(n11905), .B(n11904), .Z(n11909) );
  NAND U12243 ( .A(n11907), .B(n11906), .Z(n11908) );
  NAND U12244 ( .A(n11909), .B(n11908), .Z(n11948) );
  NAND U12245 ( .A(b[0]), .B(a[289]), .Z(n11910) );
  XNOR U12246 ( .A(b[1]), .B(n11910), .Z(n11912) );
  NAND U12247 ( .A(n56), .B(a[288]), .Z(n11911) );
  AND U12248 ( .A(n11912), .B(n11911), .Z(n11965) );
  XOR U12249 ( .A(a[285]), .B(n42197), .Z(n11954) );
  NANDN U12250 ( .A(n11954), .B(n42173), .Z(n11915) );
  NANDN U12251 ( .A(n11913), .B(n42172), .Z(n11914) );
  NAND U12252 ( .A(n11915), .B(n11914), .Z(n11963) );
  NAND U12253 ( .A(b[7]), .B(a[281]), .Z(n11964) );
  XNOR U12254 ( .A(n11963), .B(n11964), .Z(n11966) );
  XOR U12255 ( .A(n11965), .B(n11966), .Z(n11972) );
  NANDN U12256 ( .A(n11916), .B(n42093), .Z(n11918) );
  XOR U12257 ( .A(n42134), .B(a[287]), .Z(n11957) );
  NANDN U12258 ( .A(n11957), .B(n42095), .Z(n11917) );
  NAND U12259 ( .A(n11918), .B(n11917), .Z(n11970) );
  NANDN U12260 ( .A(n11919), .B(n42231), .Z(n11921) );
  XOR U12261 ( .A(n185), .B(a[283]), .Z(n11960) );
  NANDN U12262 ( .A(n11960), .B(n42234), .Z(n11920) );
  AND U12263 ( .A(n11921), .B(n11920), .Z(n11969) );
  XNOR U12264 ( .A(n11970), .B(n11969), .Z(n11971) );
  XNOR U12265 ( .A(n11972), .B(n11971), .Z(n11976) );
  NANDN U12266 ( .A(n11923), .B(n11922), .Z(n11927) );
  NAND U12267 ( .A(n11925), .B(n11924), .Z(n11926) );
  AND U12268 ( .A(n11927), .B(n11926), .Z(n11975) );
  XOR U12269 ( .A(n11976), .B(n11975), .Z(n11977) );
  NANDN U12270 ( .A(n11929), .B(n11928), .Z(n11933) );
  NANDN U12271 ( .A(n11931), .B(n11930), .Z(n11932) );
  NAND U12272 ( .A(n11933), .B(n11932), .Z(n11978) );
  XOR U12273 ( .A(n11977), .B(n11978), .Z(n11945) );
  OR U12274 ( .A(n11935), .B(n11934), .Z(n11939) );
  NANDN U12275 ( .A(n11937), .B(n11936), .Z(n11938) );
  NAND U12276 ( .A(n11939), .B(n11938), .Z(n11946) );
  XNOR U12277 ( .A(n11945), .B(n11946), .Z(n11947) );
  XNOR U12278 ( .A(n11948), .B(n11947), .Z(n11981) );
  XNOR U12279 ( .A(n11981), .B(sreg[1305]), .Z(n11983) );
  NAND U12280 ( .A(n11940), .B(sreg[1304]), .Z(n11944) );
  OR U12281 ( .A(n11942), .B(n11941), .Z(n11943) );
  AND U12282 ( .A(n11944), .B(n11943), .Z(n11982) );
  XOR U12283 ( .A(n11983), .B(n11982), .Z(c[1305]) );
  NANDN U12284 ( .A(n11946), .B(n11945), .Z(n11950) );
  NAND U12285 ( .A(n11948), .B(n11947), .Z(n11949) );
  NAND U12286 ( .A(n11950), .B(n11949), .Z(n11989) );
  NAND U12287 ( .A(b[0]), .B(a[290]), .Z(n11951) );
  XNOR U12288 ( .A(b[1]), .B(n11951), .Z(n11953) );
  NAND U12289 ( .A(n56), .B(a[289]), .Z(n11952) );
  AND U12290 ( .A(n11953), .B(n11952), .Z(n12006) );
  XOR U12291 ( .A(a[286]), .B(n42197), .Z(n11995) );
  NANDN U12292 ( .A(n11995), .B(n42173), .Z(n11956) );
  NANDN U12293 ( .A(n11954), .B(n42172), .Z(n11955) );
  NAND U12294 ( .A(n11956), .B(n11955), .Z(n12004) );
  NAND U12295 ( .A(b[7]), .B(a[282]), .Z(n12005) );
  XNOR U12296 ( .A(n12004), .B(n12005), .Z(n12007) );
  XOR U12297 ( .A(n12006), .B(n12007), .Z(n12013) );
  NANDN U12298 ( .A(n11957), .B(n42093), .Z(n11959) );
  XOR U12299 ( .A(n42134), .B(a[288]), .Z(n11998) );
  NANDN U12300 ( .A(n11998), .B(n42095), .Z(n11958) );
  NAND U12301 ( .A(n11959), .B(n11958), .Z(n12011) );
  NANDN U12302 ( .A(n11960), .B(n42231), .Z(n11962) );
  XOR U12303 ( .A(n185), .B(a[284]), .Z(n12001) );
  NANDN U12304 ( .A(n12001), .B(n42234), .Z(n11961) );
  AND U12305 ( .A(n11962), .B(n11961), .Z(n12010) );
  XNOR U12306 ( .A(n12011), .B(n12010), .Z(n12012) );
  XNOR U12307 ( .A(n12013), .B(n12012), .Z(n12017) );
  NANDN U12308 ( .A(n11964), .B(n11963), .Z(n11968) );
  NAND U12309 ( .A(n11966), .B(n11965), .Z(n11967) );
  AND U12310 ( .A(n11968), .B(n11967), .Z(n12016) );
  XOR U12311 ( .A(n12017), .B(n12016), .Z(n12018) );
  NANDN U12312 ( .A(n11970), .B(n11969), .Z(n11974) );
  NANDN U12313 ( .A(n11972), .B(n11971), .Z(n11973) );
  NAND U12314 ( .A(n11974), .B(n11973), .Z(n12019) );
  XOR U12315 ( .A(n12018), .B(n12019), .Z(n11986) );
  OR U12316 ( .A(n11976), .B(n11975), .Z(n11980) );
  NANDN U12317 ( .A(n11978), .B(n11977), .Z(n11979) );
  NAND U12318 ( .A(n11980), .B(n11979), .Z(n11987) );
  XNOR U12319 ( .A(n11986), .B(n11987), .Z(n11988) );
  XNOR U12320 ( .A(n11989), .B(n11988), .Z(n12022) );
  XNOR U12321 ( .A(n12022), .B(sreg[1306]), .Z(n12024) );
  NAND U12322 ( .A(n11981), .B(sreg[1305]), .Z(n11985) );
  OR U12323 ( .A(n11983), .B(n11982), .Z(n11984) );
  AND U12324 ( .A(n11985), .B(n11984), .Z(n12023) );
  XOR U12325 ( .A(n12024), .B(n12023), .Z(c[1306]) );
  NANDN U12326 ( .A(n11987), .B(n11986), .Z(n11991) );
  NAND U12327 ( .A(n11989), .B(n11988), .Z(n11990) );
  NAND U12328 ( .A(n11991), .B(n11990), .Z(n12030) );
  NAND U12329 ( .A(b[0]), .B(a[291]), .Z(n11992) );
  XNOR U12330 ( .A(b[1]), .B(n11992), .Z(n11994) );
  NAND U12331 ( .A(n56), .B(a[290]), .Z(n11993) );
  AND U12332 ( .A(n11994), .B(n11993), .Z(n12047) );
  XOR U12333 ( .A(a[287]), .B(n42197), .Z(n12036) );
  NANDN U12334 ( .A(n12036), .B(n42173), .Z(n11997) );
  NANDN U12335 ( .A(n11995), .B(n42172), .Z(n11996) );
  NAND U12336 ( .A(n11997), .B(n11996), .Z(n12045) );
  NAND U12337 ( .A(b[7]), .B(a[283]), .Z(n12046) );
  XNOR U12338 ( .A(n12045), .B(n12046), .Z(n12048) );
  XOR U12339 ( .A(n12047), .B(n12048), .Z(n12054) );
  NANDN U12340 ( .A(n11998), .B(n42093), .Z(n12000) );
  XOR U12341 ( .A(n42134), .B(a[289]), .Z(n12039) );
  NANDN U12342 ( .A(n12039), .B(n42095), .Z(n11999) );
  NAND U12343 ( .A(n12000), .B(n11999), .Z(n12052) );
  NANDN U12344 ( .A(n12001), .B(n42231), .Z(n12003) );
  XOR U12345 ( .A(n185), .B(a[285]), .Z(n12042) );
  NANDN U12346 ( .A(n12042), .B(n42234), .Z(n12002) );
  AND U12347 ( .A(n12003), .B(n12002), .Z(n12051) );
  XNOR U12348 ( .A(n12052), .B(n12051), .Z(n12053) );
  XNOR U12349 ( .A(n12054), .B(n12053), .Z(n12058) );
  NANDN U12350 ( .A(n12005), .B(n12004), .Z(n12009) );
  NAND U12351 ( .A(n12007), .B(n12006), .Z(n12008) );
  AND U12352 ( .A(n12009), .B(n12008), .Z(n12057) );
  XOR U12353 ( .A(n12058), .B(n12057), .Z(n12059) );
  NANDN U12354 ( .A(n12011), .B(n12010), .Z(n12015) );
  NANDN U12355 ( .A(n12013), .B(n12012), .Z(n12014) );
  NAND U12356 ( .A(n12015), .B(n12014), .Z(n12060) );
  XOR U12357 ( .A(n12059), .B(n12060), .Z(n12027) );
  OR U12358 ( .A(n12017), .B(n12016), .Z(n12021) );
  NANDN U12359 ( .A(n12019), .B(n12018), .Z(n12020) );
  NAND U12360 ( .A(n12021), .B(n12020), .Z(n12028) );
  XNOR U12361 ( .A(n12027), .B(n12028), .Z(n12029) );
  XNOR U12362 ( .A(n12030), .B(n12029), .Z(n12063) );
  XNOR U12363 ( .A(n12063), .B(sreg[1307]), .Z(n12065) );
  NAND U12364 ( .A(n12022), .B(sreg[1306]), .Z(n12026) );
  OR U12365 ( .A(n12024), .B(n12023), .Z(n12025) );
  AND U12366 ( .A(n12026), .B(n12025), .Z(n12064) );
  XOR U12367 ( .A(n12065), .B(n12064), .Z(c[1307]) );
  NANDN U12368 ( .A(n12028), .B(n12027), .Z(n12032) );
  NAND U12369 ( .A(n12030), .B(n12029), .Z(n12031) );
  NAND U12370 ( .A(n12032), .B(n12031), .Z(n12071) );
  NAND U12371 ( .A(b[0]), .B(a[292]), .Z(n12033) );
  XNOR U12372 ( .A(b[1]), .B(n12033), .Z(n12035) );
  NAND U12373 ( .A(n56), .B(a[291]), .Z(n12034) );
  AND U12374 ( .A(n12035), .B(n12034), .Z(n12088) );
  XOR U12375 ( .A(a[288]), .B(n42197), .Z(n12077) );
  NANDN U12376 ( .A(n12077), .B(n42173), .Z(n12038) );
  NANDN U12377 ( .A(n12036), .B(n42172), .Z(n12037) );
  NAND U12378 ( .A(n12038), .B(n12037), .Z(n12086) );
  NAND U12379 ( .A(b[7]), .B(a[284]), .Z(n12087) );
  XNOR U12380 ( .A(n12086), .B(n12087), .Z(n12089) );
  XOR U12381 ( .A(n12088), .B(n12089), .Z(n12095) );
  NANDN U12382 ( .A(n12039), .B(n42093), .Z(n12041) );
  XOR U12383 ( .A(n42134), .B(a[290]), .Z(n12080) );
  NANDN U12384 ( .A(n12080), .B(n42095), .Z(n12040) );
  NAND U12385 ( .A(n12041), .B(n12040), .Z(n12093) );
  NANDN U12386 ( .A(n12042), .B(n42231), .Z(n12044) );
  XOR U12387 ( .A(n185), .B(a[286]), .Z(n12083) );
  NANDN U12388 ( .A(n12083), .B(n42234), .Z(n12043) );
  AND U12389 ( .A(n12044), .B(n12043), .Z(n12092) );
  XNOR U12390 ( .A(n12093), .B(n12092), .Z(n12094) );
  XNOR U12391 ( .A(n12095), .B(n12094), .Z(n12099) );
  NANDN U12392 ( .A(n12046), .B(n12045), .Z(n12050) );
  NAND U12393 ( .A(n12048), .B(n12047), .Z(n12049) );
  AND U12394 ( .A(n12050), .B(n12049), .Z(n12098) );
  XOR U12395 ( .A(n12099), .B(n12098), .Z(n12100) );
  NANDN U12396 ( .A(n12052), .B(n12051), .Z(n12056) );
  NANDN U12397 ( .A(n12054), .B(n12053), .Z(n12055) );
  NAND U12398 ( .A(n12056), .B(n12055), .Z(n12101) );
  XOR U12399 ( .A(n12100), .B(n12101), .Z(n12068) );
  OR U12400 ( .A(n12058), .B(n12057), .Z(n12062) );
  NANDN U12401 ( .A(n12060), .B(n12059), .Z(n12061) );
  NAND U12402 ( .A(n12062), .B(n12061), .Z(n12069) );
  XNOR U12403 ( .A(n12068), .B(n12069), .Z(n12070) );
  XNOR U12404 ( .A(n12071), .B(n12070), .Z(n12104) );
  XNOR U12405 ( .A(n12104), .B(sreg[1308]), .Z(n12106) );
  NAND U12406 ( .A(n12063), .B(sreg[1307]), .Z(n12067) );
  OR U12407 ( .A(n12065), .B(n12064), .Z(n12066) );
  AND U12408 ( .A(n12067), .B(n12066), .Z(n12105) );
  XOR U12409 ( .A(n12106), .B(n12105), .Z(c[1308]) );
  NANDN U12410 ( .A(n12069), .B(n12068), .Z(n12073) );
  NAND U12411 ( .A(n12071), .B(n12070), .Z(n12072) );
  NAND U12412 ( .A(n12073), .B(n12072), .Z(n12112) );
  NAND U12413 ( .A(b[0]), .B(a[293]), .Z(n12074) );
  XNOR U12414 ( .A(b[1]), .B(n12074), .Z(n12076) );
  NAND U12415 ( .A(n56), .B(a[292]), .Z(n12075) );
  AND U12416 ( .A(n12076), .B(n12075), .Z(n12129) );
  XOR U12417 ( .A(a[289]), .B(n42197), .Z(n12118) );
  NANDN U12418 ( .A(n12118), .B(n42173), .Z(n12079) );
  NANDN U12419 ( .A(n12077), .B(n42172), .Z(n12078) );
  NAND U12420 ( .A(n12079), .B(n12078), .Z(n12127) );
  NAND U12421 ( .A(b[7]), .B(a[285]), .Z(n12128) );
  XNOR U12422 ( .A(n12127), .B(n12128), .Z(n12130) );
  XOR U12423 ( .A(n12129), .B(n12130), .Z(n12136) );
  NANDN U12424 ( .A(n12080), .B(n42093), .Z(n12082) );
  XOR U12425 ( .A(n42134), .B(a[291]), .Z(n12121) );
  NANDN U12426 ( .A(n12121), .B(n42095), .Z(n12081) );
  NAND U12427 ( .A(n12082), .B(n12081), .Z(n12134) );
  NANDN U12428 ( .A(n12083), .B(n42231), .Z(n12085) );
  XOR U12429 ( .A(n186), .B(a[287]), .Z(n12124) );
  NANDN U12430 ( .A(n12124), .B(n42234), .Z(n12084) );
  AND U12431 ( .A(n12085), .B(n12084), .Z(n12133) );
  XNOR U12432 ( .A(n12134), .B(n12133), .Z(n12135) );
  XNOR U12433 ( .A(n12136), .B(n12135), .Z(n12140) );
  NANDN U12434 ( .A(n12087), .B(n12086), .Z(n12091) );
  NAND U12435 ( .A(n12089), .B(n12088), .Z(n12090) );
  AND U12436 ( .A(n12091), .B(n12090), .Z(n12139) );
  XOR U12437 ( .A(n12140), .B(n12139), .Z(n12141) );
  NANDN U12438 ( .A(n12093), .B(n12092), .Z(n12097) );
  NANDN U12439 ( .A(n12095), .B(n12094), .Z(n12096) );
  NAND U12440 ( .A(n12097), .B(n12096), .Z(n12142) );
  XOR U12441 ( .A(n12141), .B(n12142), .Z(n12109) );
  OR U12442 ( .A(n12099), .B(n12098), .Z(n12103) );
  NANDN U12443 ( .A(n12101), .B(n12100), .Z(n12102) );
  NAND U12444 ( .A(n12103), .B(n12102), .Z(n12110) );
  XNOR U12445 ( .A(n12109), .B(n12110), .Z(n12111) );
  XNOR U12446 ( .A(n12112), .B(n12111), .Z(n12145) );
  XNOR U12447 ( .A(n12145), .B(sreg[1309]), .Z(n12147) );
  NAND U12448 ( .A(n12104), .B(sreg[1308]), .Z(n12108) );
  OR U12449 ( .A(n12106), .B(n12105), .Z(n12107) );
  AND U12450 ( .A(n12108), .B(n12107), .Z(n12146) );
  XOR U12451 ( .A(n12147), .B(n12146), .Z(c[1309]) );
  NANDN U12452 ( .A(n12110), .B(n12109), .Z(n12114) );
  NAND U12453 ( .A(n12112), .B(n12111), .Z(n12113) );
  NAND U12454 ( .A(n12114), .B(n12113), .Z(n12153) );
  NAND U12455 ( .A(b[0]), .B(a[294]), .Z(n12115) );
  XNOR U12456 ( .A(b[1]), .B(n12115), .Z(n12117) );
  NAND U12457 ( .A(n57), .B(a[293]), .Z(n12116) );
  AND U12458 ( .A(n12117), .B(n12116), .Z(n12170) );
  XOR U12459 ( .A(a[290]), .B(n42197), .Z(n12159) );
  NANDN U12460 ( .A(n12159), .B(n42173), .Z(n12120) );
  NANDN U12461 ( .A(n12118), .B(n42172), .Z(n12119) );
  NAND U12462 ( .A(n12120), .B(n12119), .Z(n12168) );
  NAND U12463 ( .A(b[7]), .B(a[286]), .Z(n12169) );
  XNOR U12464 ( .A(n12168), .B(n12169), .Z(n12171) );
  XOR U12465 ( .A(n12170), .B(n12171), .Z(n12177) );
  NANDN U12466 ( .A(n12121), .B(n42093), .Z(n12123) );
  XOR U12467 ( .A(n42134), .B(a[292]), .Z(n12162) );
  NANDN U12468 ( .A(n12162), .B(n42095), .Z(n12122) );
  NAND U12469 ( .A(n12123), .B(n12122), .Z(n12175) );
  NANDN U12470 ( .A(n12124), .B(n42231), .Z(n12126) );
  XOR U12471 ( .A(n186), .B(a[288]), .Z(n12165) );
  NANDN U12472 ( .A(n12165), .B(n42234), .Z(n12125) );
  AND U12473 ( .A(n12126), .B(n12125), .Z(n12174) );
  XNOR U12474 ( .A(n12175), .B(n12174), .Z(n12176) );
  XNOR U12475 ( .A(n12177), .B(n12176), .Z(n12181) );
  NANDN U12476 ( .A(n12128), .B(n12127), .Z(n12132) );
  NAND U12477 ( .A(n12130), .B(n12129), .Z(n12131) );
  AND U12478 ( .A(n12132), .B(n12131), .Z(n12180) );
  XOR U12479 ( .A(n12181), .B(n12180), .Z(n12182) );
  NANDN U12480 ( .A(n12134), .B(n12133), .Z(n12138) );
  NANDN U12481 ( .A(n12136), .B(n12135), .Z(n12137) );
  NAND U12482 ( .A(n12138), .B(n12137), .Z(n12183) );
  XOR U12483 ( .A(n12182), .B(n12183), .Z(n12150) );
  OR U12484 ( .A(n12140), .B(n12139), .Z(n12144) );
  NANDN U12485 ( .A(n12142), .B(n12141), .Z(n12143) );
  NAND U12486 ( .A(n12144), .B(n12143), .Z(n12151) );
  XNOR U12487 ( .A(n12150), .B(n12151), .Z(n12152) );
  XNOR U12488 ( .A(n12153), .B(n12152), .Z(n12186) );
  XNOR U12489 ( .A(n12186), .B(sreg[1310]), .Z(n12188) );
  NAND U12490 ( .A(n12145), .B(sreg[1309]), .Z(n12149) );
  OR U12491 ( .A(n12147), .B(n12146), .Z(n12148) );
  AND U12492 ( .A(n12149), .B(n12148), .Z(n12187) );
  XOR U12493 ( .A(n12188), .B(n12187), .Z(c[1310]) );
  NANDN U12494 ( .A(n12151), .B(n12150), .Z(n12155) );
  NAND U12495 ( .A(n12153), .B(n12152), .Z(n12154) );
  NAND U12496 ( .A(n12155), .B(n12154), .Z(n12194) );
  NAND U12497 ( .A(b[0]), .B(a[295]), .Z(n12156) );
  XNOR U12498 ( .A(b[1]), .B(n12156), .Z(n12158) );
  NAND U12499 ( .A(n57), .B(a[294]), .Z(n12157) );
  AND U12500 ( .A(n12158), .B(n12157), .Z(n12211) );
  XOR U12501 ( .A(a[291]), .B(n42197), .Z(n12200) );
  NANDN U12502 ( .A(n12200), .B(n42173), .Z(n12161) );
  NANDN U12503 ( .A(n12159), .B(n42172), .Z(n12160) );
  NAND U12504 ( .A(n12161), .B(n12160), .Z(n12209) );
  NAND U12505 ( .A(b[7]), .B(a[287]), .Z(n12210) );
  XNOR U12506 ( .A(n12209), .B(n12210), .Z(n12212) );
  XOR U12507 ( .A(n12211), .B(n12212), .Z(n12218) );
  NANDN U12508 ( .A(n12162), .B(n42093), .Z(n12164) );
  XOR U12509 ( .A(n42134), .B(a[293]), .Z(n12203) );
  NANDN U12510 ( .A(n12203), .B(n42095), .Z(n12163) );
  NAND U12511 ( .A(n12164), .B(n12163), .Z(n12216) );
  NANDN U12512 ( .A(n12165), .B(n42231), .Z(n12167) );
  XOR U12513 ( .A(n186), .B(a[289]), .Z(n12206) );
  NANDN U12514 ( .A(n12206), .B(n42234), .Z(n12166) );
  AND U12515 ( .A(n12167), .B(n12166), .Z(n12215) );
  XNOR U12516 ( .A(n12216), .B(n12215), .Z(n12217) );
  XNOR U12517 ( .A(n12218), .B(n12217), .Z(n12222) );
  NANDN U12518 ( .A(n12169), .B(n12168), .Z(n12173) );
  NAND U12519 ( .A(n12171), .B(n12170), .Z(n12172) );
  AND U12520 ( .A(n12173), .B(n12172), .Z(n12221) );
  XOR U12521 ( .A(n12222), .B(n12221), .Z(n12223) );
  NANDN U12522 ( .A(n12175), .B(n12174), .Z(n12179) );
  NANDN U12523 ( .A(n12177), .B(n12176), .Z(n12178) );
  NAND U12524 ( .A(n12179), .B(n12178), .Z(n12224) );
  XOR U12525 ( .A(n12223), .B(n12224), .Z(n12191) );
  OR U12526 ( .A(n12181), .B(n12180), .Z(n12185) );
  NANDN U12527 ( .A(n12183), .B(n12182), .Z(n12184) );
  NAND U12528 ( .A(n12185), .B(n12184), .Z(n12192) );
  XNOR U12529 ( .A(n12191), .B(n12192), .Z(n12193) );
  XNOR U12530 ( .A(n12194), .B(n12193), .Z(n12227) );
  XNOR U12531 ( .A(n12227), .B(sreg[1311]), .Z(n12229) );
  NAND U12532 ( .A(n12186), .B(sreg[1310]), .Z(n12190) );
  OR U12533 ( .A(n12188), .B(n12187), .Z(n12189) );
  AND U12534 ( .A(n12190), .B(n12189), .Z(n12228) );
  XOR U12535 ( .A(n12229), .B(n12228), .Z(c[1311]) );
  NANDN U12536 ( .A(n12192), .B(n12191), .Z(n12196) );
  NAND U12537 ( .A(n12194), .B(n12193), .Z(n12195) );
  NAND U12538 ( .A(n12196), .B(n12195), .Z(n12235) );
  NAND U12539 ( .A(b[0]), .B(a[296]), .Z(n12197) );
  XNOR U12540 ( .A(b[1]), .B(n12197), .Z(n12199) );
  NAND U12541 ( .A(n57), .B(a[295]), .Z(n12198) );
  AND U12542 ( .A(n12199), .B(n12198), .Z(n12252) );
  XOR U12543 ( .A(a[292]), .B(n42197), .Z(n12241) );
  NANDN U12544 ( .A(n12241), .B(n42173), .Z(n12202) );
  NANDN U12545 ( .A(n12200), .B(n42172), .Z(n12201) );
  NAND U12546 ( .A(n12202), .B(n12201), .Z(n12250) );
  NAND U12547 ( .A(b[7]), .B(a[288]), .Z(n12251) );
  XNOR U12548 ( .A(n12250), .B(n12251), .Z(n12253) );
  XOR U12549 ( .A(n12252), .B(n12253), .Z(n12259) );
  NANDN U12550 ( .A(n12203), .B(n42093), .Z(n12205) );
  XOR U12551 ( .A(n42134), .B(a[294]), .Z(n12244) );
  NANDN U12552 ( .A(n12244), .B(n42095), .Z(n12204) );
  NAND U12553 ( .A(n12205), .B(n12204), .Z(n12257) );
  NANDN U12554 ( .A(n12206), .B(n42231), .Z(n12208) );
  XOR U12555 ( .A(n186), .B(a[290]), .Z(n12247) );
  NANDN U12556 ( .A(n12247), .B(n42234), .Z(n12207) );
  AND U12557 ( .A(n12208), .B(n12207), .Z(n12256) );
  XNOR U12558 ( .A(n12257), .B(n12256), .Z(n12258) );
  XNOR U12559 ( .A(n12259), .B(n12258), .Z(n12263) );
  NANDN U12560 ( .A(n12210), .B(n12209), .Z(n12214) );
  NAND U12561 ( .A(n12212), .B(n12211), .Z(n12213) );
  AND U12562 ( .A(n12214), .B(n12213), .Z(n12262) );
  XOR U12563 ( .A(n12263), .B(n12262), .Z(n12264) );
  NANDN U12564 ( .A(n12216), .B(n12215), .Z(n12220) );
  NANDN U12565 ( .A(n12218), .B(n12217), .Z(n12219) );
  NAND U12566 ( .A(n12220), .B(n12219), .Z(n12265) );
  XOR U12567 ( .A(n12264), .B(n12265), .Z(n12232) );
  OR U12568 ( .A(n12222), .B(n12221), .Z(n12226) );
  NANDN U12569 ( .A(n12224), .B(n12223), .Z(n12225) );
  NAND U12570 ( .A(n12226), .B(n12225), .Z(n12233) );
  XNOR U12571 ( .A(n12232), .B(n12233), .Z(n12234) );
  XNOR U12572 ( .A(n12235), .B(n12234), .Z(n12268) );
  XNOR U12573 ( .A(n12268), .B(sreg[1312]), .Z(n12270) );
  NAND U12574 ( .A(n12227), .B(sreg[1311]), .Z(n12231) );
  OR U12575 ( .A(n12229), .B(n12228), .Z(n12230) );
  AND U12576 ( .A(n12231), .B(n12230), .Z(n12269) );
  XOR U12577 ( .A(n12270), .B(n12269), .Z(c[1312]) );
  NANDN U12578 ( .A(n12233), .B(n12232), .Z(n12237) );
  NAND U12579 ( .A(n12235), .B(n12234), .Z(n12236) );
  NAND U12580 ( .A(n12237), .B(n12236), .Z(n12276) );
  NAND U12581 ( .A(b[0]), .B(a[297]), .Z(n12238) );
  XNOR U12582 ( .A(b[1]), .B(n12238), .Z(n12240) );
  NAND U12583 ( .A(n57), .B(a[296]), .Z(n12239) );
  AND U12584 ( .A(n12240), .B(n12239), .Z(n12293) );
  XOR U12585 ( .A(a[293]), .B(n42197), .Z(n12282) );
  NANDN U12586 ( .A(n12282), .B(n42173), .Z(n12243) );
  NANDN U12587 ( .A(n12241), .B(n42172), .Z(n12242) );
  NAND U12588 ( .A(n12243), .B(n12242), .Z(n12291) );
  NAND U12589 ( .A(b[7]), .B(a[289]), .Z(n12292) );
  XNOR U12590 ( .A(n12291), .B(n12292), .Z(n12294) );
  XOR U12591 ( .A(n12293), .B(n12294), .Z(n12300) );
  NANDN U12592 ( .A(n12244), .B(n42093), .Z(n12246) );
  XOR U12593 ( .A(n42134), .B(a[295]), .Z(n12285) );
  NANDN U12594 ( .A(n12285), .B(n42095), .Z(n12245) );
  NAND U12595 ( .A(n12246), .B(n12245), .Z(n12298) );
  NANDN U12596 ( .A(n12247), .B(n42231), .Z(n12249) );
  XOR U12597 ( .A(n186), .B(a[291]), .Z(n12288) );
  NANDN U12598 ( .A(n12288), .B(n42234), .Z(n12248) );
  AND U12599 ( .A(n12249), .B(n12248), .Z(n12297) );
  XNOR U12600 ( .A(n12298), .B(n12297), .Z(n12299) );
  XNOR U12601 ( .A(n12300), .B(n12299), .Z(n12304) );
  NANDN U12602 ( .A(n12251), .B(n12250), .Z(n12255) );
  NAND U12603 ( .A(n12253), .B(n12252), .Z(n12254) );
  AND U12604 ( .A(n12255), .B(n12254), .Z(n12303) );
  XOR U12605 ( .A(n12304), .B(n12303), .Z(n12305) );
  NANDN U12606 ( .A(n12257), .B(n12256), .Z(n12261) );
  NANDN U12607 ( .A(n12259), .B(n12258), .Z(n12260) );
  NAND U12608 ( .A(n12261), .B(n12260), .Z(n12306) );
  XOR U12609 ( .A(n12305), .B(n12306), .Z(n12273) );
  OR U12610 ( .A(n12263), .B(n12262), .Z(n12267) );
  NANDN U12611 ( .A(n12265), .B(n12264), .Z(n12266) );
  NAND U12612 ( .A(n12267), .B(n12266), .Z(n12274) );
  XNOR U12613 ( .A(n12273), .B(n12274), .Z(n12275) );
  XNOR U12614 ( .A(n12276), .B(n12275), .Z(n12309) );
  XNOR U12615 ( .A(n12309), .B(sreg[1313]), .Z(n12311) );
  NAND U12616 ( .A(n12268), .B(sreg[1312]), .Z(n12272) );
  OR U12617 ( .A(n12270), .B(n12269), .Z(n12271) );
  AND U12618 ( .A(n12272), .B(n12271), .Z(n12310) );
  XOR U12619 ( .A(n12311), .B(n12310), .Z(c[1313]) );
  NANDN U12620 ( .A(n12274), .B(n12273), .Z(n12278) );
  NAND U12621 ( .A(n12276), .B(n12275), .Z(n12277) );
  NAND U12622 ( .A(n12278), .B(n12277), .Z(n12317) );
  NAND U12623 ( .A(b[0]), .B(a[298]), .Z(n12279) );
  XNOR U12624 ( .A(b[1]), .B(n12279), .Z(n12281) );
  NAND U12625 ( .A(n57), .B(a[297]), .Z(n12280) );
  AND U12626 ( .A(n12281), .B(n12280), .Z(n12334) );
  XOR U12627 ( .A(a[294]), .B(n42197), .Z(n12323) );
  NANDN U12628 ( .A(n12323), .B(n42173), .Z(n12284) );
  NANDN U12629 ( .A(n12282), .B(n42172), .Z(n12283) );
  NAND U12630 ( .A(n12284), .B(n12283), .Z(n12332) );
  NAND U12631 ( .A(b[7]), .B(a[290]), .Z(n12333) );
  XNOR U12632 ( .A(n12332), .B(n12333), .Z(n12335) );
  XOR U12633 ( .A(n12334), .B(n12335), .Z(n12341) );
  NANDN U12634 ( .A(n12285), .B(n42093), .Z(n12287) );
  XOR U12635 ( .A(n42134), .B(a[296]), .Z(n12326) );
  NANDN U12636 ( .A(n12326), .B(n42095), .Z(n12286) );
  NAND U12637 ( .A(n12287), .B(n12286), .Z(n12339) );
  NANDN U12638 ( .A(n12288), .B(n42231), .Z(n12290) );
  XOR U12639 ( .A(n186), .B(a[292]), .Z(n12329) );
  NANDN U12640 ( .A(n12329), .B(n42234), .Z(n12289) );
  AND U12641 ( .A(n12290), .B(n12289), .Z(n12338) );
  XNOR U12642 ( .A(n12339), .B(n12338), .Z(n12340) );
  XNOR U12643 ( .A(n12341), .B(n12340), .Z(n12345) );
  NANDN U12644 ( .A(n12292), .B(n12291), .Z(n12296) );
  NAND U12645 ( .A(n12294), .B(n12293), .Z(n12295) );
  AND U12646 ( .A(n12296), .B(n12295), .Z(n12344) );
  XOR U12647 ( .A(n12345), .B(n12344), .Z(n12346) );
  NANDN U12648 ( .A(n12298), .B(n12297), .Z(n12302) );
  NANDN U12649 ( .A(n12300), .B(n12299), .Z(n12301) );
  NAND U12650 ( .A(n12302), .B(n12301), .Z(n12347) );
  XOR U12651 ( .A(n12346), .B(n12347), .Z(n12314) );
  OR U12652 ( .A(n12304), .B(n12303), .Z(n12308) );
  NANDN U12653 ( .A(n12306), .B(n12305), .Z(n12307) );
  NAND U12654 ( .A(n12308), .B(n12307), .Z(n12315) );
  XNOR U12655 ( .A(n12314), .B(n12315), .Z(n12316) );
  XNOR U12656 ( .A(n12317), .B(n12316), .Z(n12350) );
  XNOR U12657 ( .A(n12350), .B(sreg[1314]), .Z(n12352) );
  NAND U12658 ( .A(n12309), .B(sreg[1313]), .Z(n12313) );
  OR U12659 ( .A(n12311), .B(n12310), .Z(n12312) );
  AND U12660 ( .A(n12313), .B(n12312), .Z(n12351) );
  XOR U12661 ( .A(n12352), .B(n12351), .Z(c[1314]) );
  NANDN U12662 ( .A(n12315), .B(n12314), .Z(n12319) );
  NAND U12663 ( .A(n12317), .B(n12316), .Z(n12318) );
  NAND U12664 ( .A(n12319), .B(n12318), .Z(n12358) );
  NAND U12665 ( .A(b[0]), .B(a[299]), .Z(n12320) );
  XNOR U12666 ( .A(b[1]), .B(n12320), .Z(n12322) );
  NAND U12667 ( .A(n57), .B(a[298]), .Z(n12321) );
  AND U12668 ( .A(n12322), .B(n12321), .Z(n12375) );
  XOR U12669 ( .A(a[295]), .B(n42197), .Z(n12364) );
  NANDN U12670 ( .A(n12364), .B(n42173), .Z(n12325) );
  NANDN U12671 ( .A(n12323), .B(n42172), .Z(n12324) );
  NAND U12672 ( .A(n12325), .B(n12324), .Z(n12373) );
  NAND U12673 ( .A(b[7]), .B(a[291]), .Z(n12374) );
  XNOR U12674 ( .A(n12373), .B(n12374), .Z(n12376) );
  XOR U12675 ( .A(n12375), .B(n12376), .Z(n12382) );
  NANDN U12676 ( .A(n12326), .B(n42093), .Z(n12328) );
  XOR U12677 ( .A(n42134), .B(a[297]), .Z(n12367) );
  NANDN U12678 ( .A(n12367), .B(n42095), .Z(n12327) );
  NAND U12679 ( .A(n12328), .B(n12327), .Z(n12380) );
  NANDN U12680 ( .A(n12329), .B(n42231), .Z(n12331) );
  XOR U12681 ( .A(n186), .B(a[293]), .Z(n12370) );
  NANDN U12682 ( .A(n12370), .B(n42234), .Z(n12330) );
  AND U12683 ( .A(n12331), .B(n12330), .Z(n12379) );
  XNOR U12684 ( .A(n12380), .B(n12379), .Z(n12381) );
  XNOR U12685 ( .A(n12382), .B(n12381), .Z(n12386) );
  NANDN U12686 ( .A(n12333), .B(n12332), .Z(n12337) );
  NAND U12687 ( .A(n12335), .B(n12334), .Z(n12336) );
  AND U12688 ( .A(n12337), .B(n12336), .Z(n12385) );
  XOR U12689 ( .A(n12386), .B(n12385), .Z(n12387) );
  NANDN U12690 ( .A(n12339), .B(n12338), .Z(n12343) );
  NANDN U12691 ( .A(n12341), .B(n12340), .Z(n12342) );
  NAND U12692 ( .A(n12343), .B(n12342), .Z(n12388) );
  XOR U12693 ( .A(n12387), .B(n12388), .Z(n12355) );
  OR U12694 ( .A(n12345), .B(n12344), .Z(n12349) );
  NANDN U12695 ( .A(n12347), .B(n12346), .Z(n12348) );
  NAND U12696 ( .A(n12349), .B(n12348), .Z(n12356) );
  XNOR U12697 ( .A(n12355), .B(n12356), .Z(n12357) );
  XNOR U12698 ( .A(n12358), .B(n12357), .Z(n12391) );
  XNOR U12699 ( .A(n12391), .B(sreg[1315]), .Z(n12393) );
  NAND U12700 ( .A(n12350), .B(sreg[1314]), .Z(n12354) );
  OR U12701 ( .A(n12352), .B(n12351), .Z(n12353) );
  AND U12702 ( .A(n12354), .B(n12353), .Z(n12392) );
  XOR U12703 ( .A(n12393), .B(n12392), .Z(c[1315]) );
  NANDN U12704 ( .A(n12356), .B(n12355), .Z(n12360) );
  NAND U12705 ( .A(n12358), .B(n12357), .Z(n12359) );
  NAND U12706 ( .A(n12360), .B(n12359), .Z(n12399) );
  NAND U12707 ( .A(b[0]), .B(a[300]), .Z(n12361) );
  XNOR U12708 ( .A(b[1]), .B(n12361), .Z(n12363) );
  NAND U12709 ( .A(n57), .B(a[299]), .Z(n12362) );
  AND U12710 ( .A(n12363), .B(n12362), .Z(n12416) );
  XOR U12711 ( .A(a[296]), .B(n42197), .Z(n12405) );
  NANDN U12712 ( .A(n12405), .B(n42173), .Z(n12366) );
  NANDN U12713 ( .A(n12364), .B(n42172), .Z(n12365) );
  NAND U12714 ( .A(n12366), .B(n12365), .Z(n12414) );
  NAND U12715 ( .A(b[7]), .B(a[292]), .Z(n12415) );
  XNOR U12716 ( .A(n12414), .B(n12415), .Z(n12417) );
  XOR U12717 ( .A(n12416), .B(n12417), .Z(n12423) );
  NANDN U12718 ( .A(n12367), .B(n42093), .Z(n12369) );
  XOR U12719 ( .A(n42134), .B(a[298]), .Z(n12408) );
  NANDN U12720 ( .A(n12408), .B(n42095), .Z(n12368) );
  NAND U12721 ( .A(n12369), .B(n12368), .Z(n12421) );
  NANDN U12722 ( .A(n12370), .B(n42231), .Z(n12372) );
  XOR U12723 ( .A(n186), .B(a[294]), .Z(n12411) );
  NANDN U12724 ( .A(n12411), .B(n42234), .Z(n12371) );
  AND U12725 ( .A(n12372), .B(n12371), .Z(n12420) );
  XNOR U12726 ( .A(n12421), .B(n12420), .Z(n12422) );
  XNOR U12727 ( .A(n12423), .B(n12422), .Z(n12427) );
  NANDN U12728 ( .A(n12374), .B(n12373), .Z(n12378) );
  NAND U12729 ( .A(n12376), .B(n12375), .Z(n12377) );
  AND U12730 ( .A(n12378), .B(n12377), .Z(n12426) );
  XOR U12731 ( .A(n12427), .B(n12426), .Z(n12428) );
  NANDN U12732 ( .A(n12380), .B(n12379), .Z(n12384) );
  NANDN U12733 ( .A(n12382), .B(n12381), .Z(n12383) );
  NAND U12734 ( .A(n12384), .B(n12383), .Z(n12429) );
  XOR U12735 ( .A(n12428), .B(n12429), .Z(n12396) );
  OR U12736 ( .A(n12386), .B(n12385), .Z(n12390) );
  NANDN U12737 ( .A(n12388), .B(n12387), .Z(n12389) );
  NAND U12738 ( .A(n12390), .B(n12389), .Z(n12397) );
  XNOR U12739 ( .A(n12396), .B(n12397), .Z(n12398) );
  XNOR U12740 ( .A(n12399), .B(n12398), .Z(n12432) );
  XNOR U12741 ( .A(n12432), .B(sreg[1316]), .Z(n12434) );
  NAND U12742 ( .A(n12391), .B(sreg[1315]), .Z(n12395) );
  OR U12743 ( .A(n12393), .B(n12392), .Z(n12394) );
  AND U12744 ( .A(n12395), .B(n12394), .Z(n12433) );
  XOR U12745 ( .A(n12434), .B(n12433), .Z(c[1316]) );
  NANDN U12746 ( .A(n12397), .B(n12396), .Z(n12401) );
  NAND U12747 ( .A(n12399), .B(n12398), .Z(n12400) );
  NAND U12748 ( .A(n12401), .B(n12400), .Z(n12440) );
  NAND U12749 ( .A(b[0]), .B(a[301]), .Z(n12402) );
  XNOR U12750 ( .A(b[1]), .B(n12402), .Z(n12404) );
  NAND U12751 ( .A(n58), .B(a[300]), .Z(n12403) );
  AND U12752 ( .A(n12404), .B(n12403), .Z(n12457) );
  XOR U12753 ( .A(a[297]), .B(n42197), .Z(n12446) );
  NANDN U12754 ( .A(n12446), .B(n42173), .Z(n12407) );
  NANDN U12755 ( .A(n12405), .B(n42172), .Z(n12406) );
  NAND U12756 ( .A(n12407), .B(n12406), .Z(n12455) );
  NAND U12757 ( .A(b[7]), .B(a[293]), .Z(n12456) );
  XNOR U12758 ( .A(n12455), .B(n12456), .Z(n12458) );
  XOR U12759 ( .A(n12457), .B(n12458), .Z(n12464) );
  NANDN U12760 ( .A(n12408), .B(n42093), .Z(n12410) );
  XOR U12761 ( .A(n42134), .B(a[299]), .Z(n12449) );
  NANDN U12762 ( .A(n12449), .B(n42095), .Z(n12409) );
  NAND U12763 ( .A(n12410), .B(n12409), .Z(n12462) );
  NANDN U12764 ( .A(n12411), .B(n42231), .Z(n12413) );
  XOR U12765 ( .A(n186), .B(a[295]), .Z(n12452) );
  NANDN U12766 ( .A(n12452), .B(n42234), .Z(n12412) );
  AND U12767 ( .A(n12413), .B(n12412), .Z(n12461) );
  XNOR U12768 ( .A(n12462), .B(n12461), .Z(n12463) );
  XNOR U12769 ( .A(n12464), .B(n12463), .Z(n12468) );
  NANDN U12770 ( .A(n12415), .B(n12414), .Z(n12419) );
  NAND U12771 ( .A(n12417), .B(n12416), .Z(n12418) );
  AND U12772 ( .A(n12419), .B(n12418), .Z(n12467) );
  XOR U12773 ( .A(n12468), .B(n12467), .Z(n12469) );
  NANDN U12774 ( .A(n12421), .B(n12420), .Z(n12425) );
  NANDN U12775 ( .A(n12423), .B(n12422), .Z(n12424) );
  NAND U12776 ( .A(n12425), .B(n12424), .Z(n12470) );
  XOR U12777 ( .A(n12469), .B(n12470), .Z(n12437) );
  OR U12778 ( .A(n12427), .B(n12426), .Z(n12431) );
  NANDN U12779 ( .A(n12429), .B(n12428), .Z(n12430) );
  NAND U12780 ( .A(n12431), .B(n12430), .Z(n12438) );
  XNOR U12781 ( .A(n12437), .B(n12438), .Z(n12439) );
  XNOR U12782 ( .A(n12440), .B(n12439), .Z(n12473) );
  XNOR U12783 ( .A(n12473), .B(sreg[1317]), .Z(n12475) );
  NAND U12784 ( .A(n12432), .B(sreg[1316]), .Z(n12436) );
  OR U12785 ( .A(n12434), .B(n12433), .Z(n12435) );
  AND U12786 ( .A(n12436), .B(n12435), .Z(n12474) );
  XOR U12787 ( .A(n12475), .B(n12474), .Z(c[1317]) );
  NANDN U12788 ( .A(n12438), .B(n12437), .Z(n12442) );
  NAND U12789 ( .A(n12440), .B(n12439), .Z(n12441) );
  NAND U12790 ( .A(n12442), .B(n12441), .Z(n12481) );
  NAND U12791 ( .A(b[0]), .B(a[302]), .Z(n12443) );
  XNOR U12792 ( .A(b[1]), .B(n12443), .Z(n12445) );
  NAND U12793 ( .A(n58), .B(a[301]), .Z(n12444) );
  AND U12794 ( .A(n12445), .B(n12444), .Z(n12498) );
  XOR U12795 ( .A(a[298]), .B(n42197), .Z(n12487) );
  NANDN U12796 ( .A(n12487), .B(n42173), .Z(n12448) );
  NANDN U12797 ( .A(n12446), .B(n42172), .Z(n12447) );
  NAND U12798 ( .A(n12448), .B(n12447), .Z(n12496) );
  NAND U12799 ( .A(b[7]), .B(a[294]), .Z(n12497) );
  XNOR U12800 ( .A(n12496), .B(n12497), .Z(n12499) );
  XOR U12801 ( .A(n12498), .B(n12499), .Z(n12505) );
  NANDN U12802 ( .A(n12449), .B(n42093), .Z(n12451) );
  XOR U12803 ( .A(n42134), .B(a[300]), .Z(n12490) );
  NANDN U12804 ( .A(n12490), .B(n42095), .Z(n12450) );
  NAND U12805 ( .A(n12451), .B(n12450), .Z(n12503) );
  NANDN U12806 ( .A(n12452), .B(n42231), .Z(n12454) );
  XOR U12807 ( .A(n186), .B(a[296]), .Z(n12493) );
  NANDN U12808 ( .A(n12493), .B(n42234), .Z(n12453) );
  AND U12809 ( .A(n12454), .B(n12453), .Z(n12502) );
  XNOR U12810 ( .A(n12503), .B(n12502), .Z(n12504) );
  XNOR U12811 ( .A(n12505), .B(n12504), .Z(n12509) );
  NANDN U12812 ( .A(n12456), .B(n12455), .Z(n12460) );
  NAND U12813 ( .A(n12458), .B(n12457), .Z(n12459) );
  AND U12814 ( .A(n12460), .B(n12459), .Z(n12508) );
  XOR U12815 ( .A(n12509), .B(n12508), .Z(n12510) );
  NANDN U12816 ( .A(n12462), .B(n12461), .Z(n12466) );
  NANDN U12817 ( .A(n12464), .B(n12463), .Z(n12465) );
  NAND U12818 ( .A(n12466), .B(n12465), .Z(n12511) );
  XOR U12819 ( .A(n12510), .B(n12511), .Z(n12478) );
  OR U12820 ( .A(n12468), .B(n12467), .Z(n12472) );
  NANDN U12821 ( .A(n12470), .B(n12469), .Z(n12471) );
  NAND U12822 ( .A(n12472), .B(n12471), .Z(n12479) );
  XNOR U12823 ( .A(n12478), .B(n12479), .Z(n12480) );
  XNOR U12824 ( .A(n12481), .B(n12480), .Z(n12514) );
  XNOR U12825 ( .A(n12514), .B(sreg[1318]), .Z(n12516) );
  NAND U12826 ( .A(n12473), .B(sreg[1317]), .Z(n12477) );
  OR U12827 ( .A(n12475), .B(n12474), .Z(n12476) );
  AND U12828 ( .A(n12477), .B(n12476), .Z(n12515) );
  XOR U12829 ( .A(n12516), .B(n12515), .Z(c[1318]) );
  NANDN U12830 ( .A(n12479), .B(n12478), .Z(n12483) );
  NAND U12831 ( .A(n12481), .B(n12480), .Z(n12482) );
  NAND U12832 ( .A(n12483), .B(n12482), .Z(n12522) );
  NAND U12833 ( .A(b[0]), .B(a[303]), .Z(n12484) );
  XNOR U12834 ( .A(b[1]), .B(n12484), .Z(n12486) );
  NAND U12835 ( .A(n58), .B(a[302]), .Z(n12485) );
  AND U12836 ( .A(n12486), .B(n12485), .Z(n12539) );
  XOR U12837 ( .A(a[299]), .B(n42197), .Z(n12528) );
  NANDN U12838 ( .A(n12528), .B(n42173), .Z(n12489) );
  NANDN U12839 ( .A(n12487), .B(n42172), .Z(n12488) );
  NAND U12840 ( .A(n12489), .B(n12488), .Z(n12537) );
  NAND U12841 ( .A(b[7]), .B(a[295]), .Z(n12538) );
  XNOR U12842 ( .A(n12537), .B(n12538), .Z(n12540) );
  XOR U12843 ( .A(n12539), .B(n12540), .Z(n12546) );
  NANDN U12844 ( .A(n12490), .B(n42093), .Z(n12492) );
  XOR U12845 ( .A(n42134), .B(a[301]), .Z(n12531) );
  NANDN U12846 ( .A(n12531), .B(n42095), .Z(n12491) );
  NAND U12847 ( .A(n12492), .B(n12491), .Z(n12544) );
  NANDN U12848 ( .A(n12493), .B(n42231), .Z(n12495) );
  XOR U12849 ( .A(n186), .B(a[297]), .Z(n12534) );
  NANDN U12850 ( .A(n12534), .B(n42234), .Z(n12494) );
  AND U12851 ( .A(n12495), .B(n12494), .Z(n12543) );
  XNOR U12852 ( .A(n12544), .B(n12543), .Z(n12545) );
  XNOR U12853 ( .A(n12546), .B(n12545), .Z(n12550) );
  NANDN U12854 ( .A(n12497), .B(n12496), .Z(n12501) );
  NAND U12855 ( .A(n12499), .B(n12498), .Z(n12500) );
  AND U12856 ( .A(n12501), .B(n12500), .Z(n12549) );
  XOR U12857 ( .A(n12550), .B(n12549), .Z(n12551) );
  NANDN U12858 ( .A(n12503), .B(n12502), .Z(n12507) );
  NANDN U12859 ( .A(n12505), .B(n12504), .Z(n12506) );
  NAND U12860 ( .A(n12507), .B(n12506), .Z(n12552) );
  XOR U12861 ( .A(n12551), .B(n12552), .Z(n12519) );
  OR U12862 ( .A(n12509), .B(n12508), .Z(n12513) );
  NANDN U12863 ( .A(n12511), .B(n12510), .Z(n12512) );
  NAND U12864 ( .A(n12513), .B(n12512), .Z(n12520) );
  XNOR U12865 ( .A(n12519), .B(n12520), .Z(n12521) );
  XNOR U12866 ( .A(n12522), .B(n12521), .Z(n12555) );
  XNOR U12867 ( .A(n12555), .B(sreg[1319]), .Z(n12557) );
  NAND U12868 ( .A(n12514), .B(sreg[1318]), .Z(n12518) );
  OR U12869 ( .A(n12516), .B(n12515), .Z(n12517) );
  AND U12870 ( .A(n12518), .B(n12517), .Z(n12556) );
  XOR U12871 ( .A(n12557), .B(n12556), .Z(c[1319]) );
  NANDN U12872 ( .A(n12520), .B(n12519), .Z(n12524) );
  NAND U12873 ( .A(n12522), .B(n12521), .Z(n12523) );
  NAND U12874 ( .A(n12524), .B(n12523), .Z(n12563) );
  NAND U12875 ( .A(b[0]), .B(a[304]), .Z(n12525) );
  XNOR U12876 ( .A(b[1]), .B(n12525), .Z(n12527) );
  NAND U12877 ( .A(n58), .B(a[303]), .Z(n12526) );
  AND U12878 ( .A(n12527), .B(n12526), .Z(n12580) );
  XOR U12879 ( .A(a[300]), .B(n42197), .Z(n12569) );
  NANDN U12880 ( .A(n12569), .B(n42173), .Z(n12530) );
  NANDN U12881 ( .A(n12528), .B(n42172), .Z(n12529) );
  NAND U12882 ( .A(n12530), .B(n12529), .Z(n12578) );
  NAND U12883 ( .A(b[7]), .B(a[296]), .Z(n12579) );
  XNOR U12884 ( .A(n12578), .B(n12579), .Z(n12581) );
  XOR U12885 ( .A(n12580), .B(n12581), .Z(n12587) );
  NANDN U12886 ( .A(n12531), .B(n42093), .Z(n12533) );
  XOR U12887 ( .A(n42134), .B(a[302]), .Z(n12572) );
  NANDN U12888 ( .A(n12572), .B(n42095), .Z(n12532) );
  NAND U12889 ( .A(n12533), .B(n12532), .Z(n12585) );
  NANDN U12890 ( .A(n12534), .B(n42231), .Z(n12536) );
  XOR U12891 ( .A(n186), .B(a[298]), .Z(n12575) );
  NANDN U12892 ( .A(n12575), .B(n42234), .Z(n12535) );
  AND U12893 ( .A(n12536), .B(n12535), .Z(n12584) );
  XNOR U12894 ( .A(n12585), .B(n12584), .Z(n12586) );
  XNOR U12895 ( .A(n12587), .B(n12586), .Z(n12591) );
  NANDN U12896 ( .A(n12538), .B(n12537), .Z(n12542) );
  NAND U12897 ( .A(n12540), .B(n12539), .Z(n12541) );
  AND U12898 ( .A(n12542), .B(n12541), .Z(n12590) );
  XOR U12899 ( .A(n12591), .B(n12590), .Z(n12592) );
  NANDN U12900 ( .A(n12544), .B(n12543), .Z(n12548) );
  NANDN U12901 ( .A(n12546), .B(n12545), .Z(n12547) );
  NAND U12902 ( .A(n12548), .B(n12547), .Z(n12593) );
  XOR U12903 ( .A(n12592), .B(n12593), .Z(n12560) );
  OR U12904 ( .A(n12550), .B(n12549), .Z(n12554) );
  NANDN U12905 ( .A(n12552), .B(n12551), .Z(n12553) );
  NAND U12906 ( .A(n12554), .B(n12553), .Z(n12561) );
  XNOR U12907 ( .A(n12560), .B(n12561), .Z(n12562) );
  XNOR U12908 ( .A(n12563), .B(n12562), .Z(n12596) );
  XNOR U12909 ( .A(n12596), .B(sreg[1320]), .Z(n12598) );
  NAND U12910 ( .A(n12555), .B(sreg[1319]), .Z(n12559) );
  OR U12911 ( .A(n12557), .B(n12556), .Z(n12558) );
  AND U12912 ( .A(n12559), .B(n12558), .Z(n12597) );
  XOR U12913 ( .A(n12598), .B(n12597), .Z(c[1320]) );
  NANDN U12914 ( .A(n12561), .B(n12560), .Z(n12565) );
  NAND U12915 ( .A(n12563), .B(n12562), .Z(n12564) );
  NAND U12916 ( .A(n12565), .B(n12564), .Z(n12604) );
  NAND U12917 ( .A(b[0]), .B(a[305]), .Z(n12566) );
  XNOR U12918 ( .A(b[1]), .B(n12566), .Z(n12568) );
  NAND U12919 ( .A(n58), .B(a[304]), .Z(n12567) );
  AND U12920 ( .A(n12568), .B(n12567), .Z(n12621) );
  XOR U12921 ( .A(a[301]), .B(n42197), .Z(n12610) );
  NANDN U12922 ( .A(n12610), .B(n42173), .Z(n12571) );
  NANDN U12923 ( .A(n12569), .B(n42172), .Z(n12570) );
  NAND U12924 ( .A(n12571), .B(n12570), .Z(n12619) );
  NAND U12925 ( .A(b[7]), .B(a[297]), .Z(n12620) );
  XNOR U12926 ( .A(n12619), .B(n12620), .Z(n12622) );
  XOR U12927 ( .A(n12621), .B(n12622), .Z(n12628) );
  NANDN U12928 ( .A(n12572), .B(n42093), .Z(n12574) );
  XOR U12929 ( .A(n42134), .B(a[303]), .Z(n12613) );
  NANDN U12930 ( .A(n12613), .B(n42095), .Z(n12573) );
  NAND U12931 ( .A(n12574), .B(n12573), .Z(n12626) );
  NANDN U12932 ( .A(n12575), .B(n42231), .Z(n12577) );
  XOR U12933 ( .A(n187), .B(a[299]), .Z(n12616) );
  NANDN U12934 ( .A(n12616), .B(n42234), .Z(n12576) );
  AND U12935 ( .A(n12577), .B(n12576), .Z(n12625) );
  XNOR U12936 ( .A(n12626), .B(n12625), .Z(n12627) );
  XNOR U12937 ( .A(n12628), .B(n12627), .Z(n12632) );
  NANDN U12938 ( .A(n12579), .B(n12578), .Z(n12583) );
  NAND U12939 ( .A(n12581), .B(n12580), .Z(n12582) );
  AND U12940 ( .A(n12583), .B(n12582), .Z(n12631) );
  XOR U12941 ( .A(n12632), .B(n12631), .Z(n12633) );
  NANDN U12942 ( .A(n12585), .B(n12584), .Z(n12589) );
  NANDN U12943 ( .A(n12587), .B(n12586), .Z(n12588) );
  NAND U12944 ( .A(n12589), .B(n12588), .Z(n12634) );
  XOR U12945 ( .A(n12633), .B(n12634), .Z(n12601) );
  OR U12946 ( .A(n12591), .B(n12590), .Z(n12595) );
  NANDN U12947 ( .A(n12593), .B(n12592), .Z(n12594) );
  NAND U12948 ( .A(n12595), .B(n12594), .Z(n12602) );
  XNOR U12949 ( .A(n12601), .B(n12602), .Z(n12603) );
  XNOR U12950 ( .A(n12604), .B(n12603), .Z(n12637) );
  XNOR U12951 ( .A(n12637), .B(sreg[1321]), .Z(n12639) );
  NAND U12952 ( .A(n12596), .B(sreg[1320]), .Z(n12600) );
  OR U12953 ( .A(n12598), .B(n12597), .Z(n12599) );
  AND U12954 ( .A(n12600), .B(n12599), .Z(n12638) );
  XOR U12955 ( .A(n12639), .B(n12638), .Z(c[1321]) );
  NANDN U12956 ( .A(n12602), .B(n12601), .Z(n12606) );
  NAND U12957 ( .A(n12604), .B(n12603), .Z(n12605) );
  NAND U12958 ( .A(n12606), .B(n12605), .Z(n12645) );
  NAND U12959 ( .A(b[0]), .B(a[306]), .Z(n12607) );
  XNOR U12960 ( .A(b[1]), .B(n12607), .Z(n12609) );
  NAND U12961 ( .A(n58), .B(a[305]), .Z(n12608) );
  AND U12962 ( .A(n12609), .B(n12608), .Z(n12662) );
  XOR U12963 ( .A(a[302]), .B(n42197), .Z(n12651) );
  NANDN U12964 ( .A(n12651), .B(n42173), .Z(n12612) );
  NANDN U12965 ( .A(n12610), .B(n42172), .Z(n12611) );
  NAND U12966 ( .A(n12612), .B(n12611), .Z(n12660) );
  NAND U12967 ( .A(b[7]), .B(a[298]), .Z(n12661) );
  XNOR U12968 ( .A(n12660), .B(n12661), .Z(n12663) );
  XOR U12969 ( .A(n12662), .B(n12663), .Z(n12669) );
  NANDN U12970 ( .A(n12613), .B(n42093), .Z(n12615) );
  XOR U12971 ( .A(n42134), .B(a[304]), .Z(n12654) );
  NANDN U12972 ( .A(n12654), .B(n42095), .Z(n12614) );
  NAND U12973 ( .A(n12615), .B(n12614), .Z(n12667) );
  NANDN U12974 ( .A(n12616), .B(n42231), .Z(n12618) );
  XOR U12975 ( .A(n187), .B(a[300]), .Z(n12657) );
  NANDN U12976 ( .A(n12657), .B(n42234), .Z(n12617) );
  AND U12977 ( .A(n12618), .B(n12617), .Z(n12666) );
  XNOR U12978 ( .A(n12667), .B(n12666), .Z(n12668) );
  XNOR U12979 ( .A(n12669), .B(n12668), .Z(n12673) );
  NANDN U12980 ( .A(n12620), .B(n12619), .Z(n12624) );
  NAND U12981 ( .A(n12622), .B(n12621), .Z(n12623) );
  AND U12982 ( .A(n12624), .B(n12623), .Z(n12672) );
  XOR U12983 ( .A(n12673), .B(n12672), .Z(n12674) );
  NANDN U12984 ( .A(n12626), .B(n12625), .Z(n12630) );
  NANDN U12985 ( .A(n12628), .B(n12627), .Z(n12629) );
  NAND U12986 ( .A(n12630), .B(n12629), .Z(n12675) );
  XOR U12987 ( .A(n12674), .B(n12675), .Z(n12642) );
  OR U12988 ( .A(n12632), .B(n12631), .Z(n12636) );
  NANDN U12989 ( .A(n12634), .B(n12633), .Z(n12635) );
  NAND U12990 ( .A(n12636), .B(n12635), .Z(n12643) );
  XNOR U12991 ( .A(n12642), .B(n12643), .Z(n12644) );
  XNOR U12992 ( .A(n12645), .B(n12644), .Z(n12678) );
  XNOR U12993 ( .A(n12678), .B(sreg[1322]), .Z(n12680) );
  NAND U12994 ( .A(n12637), .B(sreg[1321]), .Z(n12641) );
  OR U12995 ( .A(n12639), .B(n12638), .Z(n12640) );
  AND U12996 ( .A(n12641), .B(n12640), .Z(n12679) );
  XOR U12997 ( .A(n12680), .B(n12679), .Z(c[1322]) );
  NANDN U12998 ( .A(n12643), .B(n12642), .Z(n12647) );
  NAND U12999 ( .A(n12645), .B(n12644), .Z(n12646) );
  NAND U13000 ( .A(n12647), .B(n12646), .Z(n12686) );
  NAND U13001 ( .A(b[0]), .B(a[307]), .Z(n12648) );
  XNOR U13002 ( .A(b[1]), .B(n12648), .Z(n12650) );
  NAND U13003 ( .A(n58), .B(a[306]), .Z(n12649) );
  AND U13004 ( .A(n12650), .B(n12649), .Z(n12703) );
  XOR U13005 ( .A(a[303]), .B(n42197), .Z(n12692) );
  NANDN U13006 ( .A(n12692), .B(n42173), .Z(n12653) );
  NANDN U13007 ( .A(n12651), .B(n42172), .Z(n12652) );
  NAND U13008 ( .A(n12653), .B(n12652), .Z(n12701) );
  NAND U13009 ( .A(b[7]), .B(a[299]), .Z(n12702) );
  XNOR U13010 ( .A(n12701), .B(n12702), .Z(n12704) );
  XOR U13011 ( .A(n12703), .B(n12704), .Z(n12710) );
  NANDN U13012 ( .A(n12654), .B(n42093), .Z(n12656) );
  XOR U13013 ( .A(n42134), .B(a[305]), .Z(n12695) );
  NANDN U13014 ( .A(n12695), .B(n42095), .Z(n12655) );
  NAND U13015 ( .A(n12656), .B(n12655), .Z(n12708) );
  NANDN U13016 ( .A(n12657), .B(n42231), .Z(n12659) );
  XOR U13017 ( .A(n187), .B(a[301]), .Z(n12698) );
  NANDN U13018 ( .A(n12698), .B(n42234), .Z(n12658) );
  AND U13019 ( .A(n12659), .B(n12658), .Z(n12707) );
  XNOR U13020 ( .A(n12708), .B(n12707), .Z(n12709) );
  XNOR U13021 ( .A(n12710), .B(n12709), .Z(n12714) );
  NANDN U13022 ( .A(n12661), .B(n12660), .Z(n12665) );
  NAND U13023 ( .A(n12663), .B(n12662), .Z(n12664) );
  AND U13024 ( .A(n12665), .B(n12664), .Z(n12713) );
  XOR U13025 ( .A(n12714), .B(n12713), .Z(n12715) );
  NANDN U13026 ( .A(n12667), .B(n12666), .Z(n12671) );
  NANDN U13027 ( .A(n12669), .B(n12668), .Z(n12670) );
  NAND U13028 ( .A(n12671), .B(n12670), .Z(n12716) );
  XOR U13029 ( .A(n12715), .B(n12716), .Z(n12683) );
  OR U13030 ( .A(n12673), .B(n12672), .Z(n12677) );
  NANDN U13031 ( .A(n12675), .B(n12674), .Z(n12676) );
  NAND U13032 ( .A(n12677), .B(n12676), .Z(n12684) );
  XNOR U13033 ( .A(n12683), .B(n12684), .Z(n12685) );
  XNOR U13034 ( .A(n12686), .B(n12685), .Z(n12719) );
  XNOR U13035 ( .A(n12719), .B(sreg[1323]), .Z(n12721) );
  NAND U13036 ( .A(n12678), .B(sreg[1322]), .Z(n12682) );
  OR U13037 ( .A(n12680), .B(n12679), .Z(n12681) );
  AND U13038 ( .A(n12682), .B(n12681), .Z(n12720) );
  XOR U13039 ( .A(n12721), .B(n12720), .Z(c[1323]) );
  NANDN U13040 ( .A(n12684), .B(n12683), .Z(n12688) );
  NAND U13041 ( .A(n12686), .B(n12685), .Z(n12687) );
  NAND U13042 ( .A(n12688), .B(n12687), .Z(n12727) );
  NAND U13043 ( .A(b[0]), .B(a[308]), .Z(n12689) );
  XNOR U13044 ( .A(b[1]), .B(n12689), .Z(n12691) );
  NAND U13045 ( .A(n59), .B(a[307]), .Z(n12690) );
  AND U13046 ( .A(n12691), .B(n12690), .Z(n12744) );
  XOR U13047 ( .A(a[304]), .B(n42197), .Z(n12733) );
  NANDN U13048 ( .A(n12733), .B(n42173), .Z(n12694) );
  NANDN U13049 ( .A(n12692), .B(n42172), .Z(n12693) );
  NAND U13050 ( .A(n12694), .B(n12693), .Z(n12742) );
  NAND U13051 ( .A(b[7]), .B(a[300]), .Z(n12743) );
  XNOR U13052 ( .A(n12742), .B(n12743), .Z(n12745) );
  XOR U13053 ( .A(n12744), .B(n12745), .Z(n12751) );
  NANDN U13054 ( .A(n12695), .B(n42093), .Z(n12697) );
  XOR U13055 ( .A(n42134), .B(a[306]), .Z(n12736) );
  NANDN U13056 ( .A(n12736), .B(n42095), .Z(n12696) );
  NAND U13057 ( .A(n12697), .B(n12696), .Z(n12749) );
  NANDN U13058 ( .A(n12698), .B(n42231), .Z(n12700) );
  XOR U13059 ( .A(n187), .B(a[302]), .Z(n12739) );
  NANDN U13060 ( .A(n12739), .B(n42234), .Z(n12699) );
  AND U13061 ( .A(n12700), .B(n12699), .Z(n12748) );
  XNOR U13062 ( .A(n12749), .B(n12748), .Z(n12750) );
  XNOR U13063 ( .A(n12751), .B(n12750), .Z(n12755) );
  NANDN U13064 ( .A(n12702), .B(n12701), .Z(n12706) );
  NAND U13065 ( .A(n12704), .B(n12703), .Z(n12705) );
  AND U13066 ( .A(n12706), .B(n12705), .Z(n12754) );
  XOR U13067 ( .A(n12755), .B(n12754), .Z(n12756) );
  NANDN U13068 ( .A(n12708), .B(n12707), .Z(n12712) );
  NANDN U13069 ( .A(n12710), .B(n12709), .Z(n12711) );
  NAND U13070 ( .A(n12712), .B(n12711), .Z(n12757) );
  XOR U13071 ( .A(n12756), .B(n12757), .Z(n12724) );
  OR U13072 ( .A(n12714), .B(n12713), .Z(n12718) );
  NANDN U13073 ( .A(n12716), .B(n12715), .Z(n12717) );
  NAND U13074 ( .A(n12718), .B(n12717), .Z(n12725) );
  XNOR U13075 ( .A(n12724), .B(n12725), .Z(n12726) );
  XNOR U13076 ( .A(n12727), .B(n12726), .Z(n12760) );
  XNOR U13077 ( .A(n12760), .B(sreg[1324]), .Z(n12762) );
  NAND U13078 ( .A(n12719), .B(sreg[1323]), .Z(n12723) );
  OR U13079 ( .A(n12721), .B(n12720), .Z(n12722) );
  AND U13080 ( .A(n12723), .B(n12722), .Z(n12761) );
  XOR U13081 ( .A(n12762), .B(n12761), .Z(c[1324]) );
  NANDN U13082 ( .A(n12725), .B(n12724), .Z(n12729) );
  NAND U13083 ( .A(n12727), .B(n12726), .Z(n12728) );
  NAND U13084 ( .A(n12729), .B(n12728), .Z(n12768) );
  NAND U13085 ( .A(b[0]), .B(a[309]), .Z(n12730) );
  XNOR U13086 ( .A(b[1]), .B(n12730), .Z(n12732) );
  NAND U13087 ( .A(n59), .B(a[308]), .Z(n12731) );
  AND U13088 ( .A(n12732), .B(n12731), .Z(n12785) );
  XOR U13089 ( .A(a[305]), .B(n42197), .Z(n12774) );
  NANDN U13090 ( .A(n12774), .B(n42173), .Z(n12735) );
  NANDN U13091 ( .A(n12733), .B(n42172), .Z(n12734) );
  NAND U13092 ( .A(n12735), .B(n12734), .Z(n12783) );
  NAND U13093 ( .A(b[7]), .B(a[301]), .Z(n12784) );
  XNOR U13094 ( .A(n12783), .B(n12784), .Z(n12786) );
  XOR U13095 ( .A(n12785), .B(n12786), .Z(n12792) );
  NANDN U13096 ( .A(n12736), .B(n42093), .Z(n12738) );
  XOR U13097 ( .A(n42134), .B(a[307]), .Z(n12777) );
  NANDN U13098 ( .A(n12777), .B(n42095), .Z(n12737) );
  NAND U13099 ( .A(n12738), .B(n12737), .Z(n12790) );
  NANDN U13100 ( .A(n12739), .B(n42231), .Z(n12741) );
  XOR U13101 ( .A(n187), .B(a[303]), .Z(n12780) );
  NANDN U13102 ( .A(n12780), .B(n42234), .Z(n12740) );
  AND U13103 ( .A(n12741), .B(n12740), .Z(n12789) );
  XNOR U13104 ( .A(n12790), .B(n12789), .Z(n12791) );
  XNOR U13105 ( .A(n12792), .B(n12791), .Z(n12796) );
  NANDN U13106 ( .A(n12743), .B(n12742), .Z(n12747) );
  NAND U13107 ( .A(n12745), .B(n12744), .Z(n12746) );
  AND U13108 ( .A(n12747), .B(n12746), .Z(n12795) );
  XOR U13109 ( .A(n12796), .B(n12795), .Z(n12797) );
  NANDN U13110 ( .A(n12749), .B(n12748), .Z(n12753) );
  NANDN U13111 ( .A(n12751), .B(n12750), .Z(n12752) );
  NAND U13112 ( .A(n12753), .B(n12752), .Z(n12798) );
  XOR U13113 ( .A(n12797), .B(n12798), .Z(n12765) );
  OR U13114 ( .A(n12755), .B(n12754), .Z(n12759) );
  NANDN U13115 ( .A(n12757), .B(n12756), .Z(n12758) );
  NAND U13116 ( .A(n12759), .B(n12758), .Z(n12766) );
  XNOR U13117 ( .A(n12765), .B(n12766), .Z(n12767) );
  XNOR U13118 ( .A(n12768), .B(n12767), .Z(n12801) );
  XNOR U13119 ( .A(n12801), .B(sreg[1325]), .Z(n12803) );
  NAND U13120 ( .A(n12760), .B(sreg[1324]), .Z(n12764) );
  OR U13121 ( .A(n12762), .B(n12761), .Z(n12763) );
  AND U13122 ( .A(n12764), .B(n12763), .Z(n12802) );
  XOR U13123 ( .A(n12803), .B(n12802), .Z(c[1325]) );
  NANDN U13124 ( .A(n12766), .B(n12765), .Z(n12770) );
  NAND U13125 ( .A(n12768), .B(n12767), .Z(n12769) );
  NAND U13126 ( .A(n12770), .B(n12769), .Z(n12809) );
  NAND U13127 ( .A(b[0]), .B(a[310]), .Z(n12771) );
  XNOR U13128 ( .A(b[1]), .B(n12771), .Z(n12773) );
  NAND U13129 ( .A(n59), .B(a[309]), .Z(n12772) );
  AND U13130 ( .A(n12773), .B(n12772), .Z(n12826) );
  XOR U13131 ( .A(a[306]), .B(n42197), .Z(n12815) );
  NANDN U13132 ( .A(n12815), .B(n42173), .Z(n12776) );
  NANDN U13133 ( .A(n12774), .B(n42172), .Z(n12775) );
  NAND U13134 ( .A(n12776), .B(n12775), .Z(n12824) );
  NAND U13135 ( .A(b[7]), .B(a[302]), .Z(n12825) );
  XNOR U13136 ( .A(n12824), .B(n12825), .Z(n12827) );
  XOR U13137 ( .A(n12826), .B(n12827), .Z(n12833) );
  NANDN U13138 ( .A(n12777), .B(n42093), .Z(n12779) );
  XOR U13139 ( .A(n42134), .B(a[308]), .Z(n12818) );
  NANDN U13140 ( .A(n12818), .B(n42095), .Z(n12778) );
  NAND U13141 ( .A(n12779), .B(n12778), .Z(n12831) );
  NANDN U13142 ( .A(n12780), .B(n42231), .Z(n12782) );
  XOR U13143 ( .A(n187), .B(a[304]), .Z(n12821) );
  NANDN U13144 ( .A(n12821), .B(n42234), .Z(n12781) );
  AND U13145 ( .A(n12782), .B(n12781), .Z(n12830) );
  XNOR U13146 ( .A(n12831), .B(n12830), .Z(n12832) );
  XNOR U13147 ( .A(n12833), .B(n12832), .Z(n12837) );
  NANDN U13148 ( .A(n12784), .B(n12783), .Z(n12788) );
  NAND U13149 ( .A(n12786), .B(n12785), .Z(n12787) );
  AND U13150 ( .A(n12788), .B(n12787), .Z(n12836) );
  XOR U13151 ( .A(n12837), .B(n12836), .Z(n12838) );
  NANDN U13152 ( .A(n12790), .B(n12789), .Z(n12794) );
  NANDN U13153 ( .A(n12792), .B(n12791), .Z(n12793) );
  NAND U13154 ( .A(n12794), .B(n12793), .Z(n12839) );
  XOR U13155 ( .A(n12838), .B(n12839), .Z(n12806) );
  OR U13156 ( .A(n12796), .B(n12795), .Z(n12800) );
  NANDN U13157 ( .A(n12798), .B(n12797), .Z(n12799) );
  NAND U13158 ( .A(n12800), .B(n12799), .Z(n12807) );
  XNOR U13159 ( .A(n12806), .B(n12807), .Z(n12808) );
  XNOR U13160 ( .A(n12809), .B(n12808), .Z(n12842) );
  XNOR U13161 ( .A(n12842), .B(sreg[1326]), .Z(n12844) );
  NAND U13162 ( .A(n12801), .B(sreg[1325]), .Z(n12805) );
  OR U13163 ( .A(n12803), .B(n12802), .Z(n12804) );
  AND U13164 ( .A(n12805), .B(n12804), .Z(n12843) );
  XOR U13165 ( .A(n12844), .B(n12843), .Z(c[1326]) );
  NANDN U13166 ( .A(n12807), .B(n12806), .Z(n12811) );
  NAND U13167 ( .A(n12809), .B(n12808), .Z(n12810) );
  NAND U13168 ( .A(n12811), .B(n12810), .Z(n12850) );
  NAND U13169 ( .A(b[0]), .B(a[311]), .Z(n12812) );
  XNOR U13170 ( .A(b[1]), .B(n12812), .Z(n12814) );
  NAND U13171 ( .A(n59), .B(a[310]), .Z(n12813) );
  AND U13172 ( .A(n12814), .B(n12813), .Z(n12867) );
  XOR U13173 ( .A(a[307]), .B(n42197), .Z(n12856) );
  NANDN U13174 ( .A(n12856), .B(n42173), .Z(n12817) );
  NANDN U13175 ( .A(n12815), .B(n42172), .Z(n12816) );
  NAND U13176 ( .A(n12817), .B(n12816), .Z(n12865) );
  NAND U13177 ( .A(b[7]), .B(a[303]), .Z(n12866) );
  XNOR U13178 ( .A(n12865), .B(n12866), .Z(n12868) );
  XOR U13179 ( .A(n12867), .B(n12868), .Z(n12874) );
  NANDN U13180 ( .A(n12818), .B(n42093), .Z(n12820) );
  XOR U13181 ( .A(n42134), .B(a[309]), .Z(n12859) );
  NANDN U13182 ( .A(n12859), .B(n42095), .Z(n12819) );
  NAND U13183 ( .A(n12820), .B(n12819), .Z(n12872) );
  NANDN U13184 ( .A(n12821), .B(n42231), .Z(n12823) );
  XOR U13185 ( .A(n187), .B(a[305]), .Z(n12862) );
  NANDN U13186 ( .A(n12862), .B(n42234), .Z(n12822) );
  AND U13187 ( .A(n12823), .B(n12822), .Z(n12871) );
  XNOR U13188 ( .A(n12872), .B(n12871), .Z(n12873) );
  XNOR U13189 ( .A(n12874), .B(n12873), .Z(n12878) );
  NANDN U13190 ( .A(n12825), .B(n12824), .Z(n12829) );
  NAND U13191 ( .A(n12827), .B(n12826), .Z(n12828) );
  AND U13192 ( .A(n12829), .B(n12828), .Z(n12877) );
  XOR U13193 ( .A(n12878), .B(n12877), .Z(n12879) );
  NANDN U13194 ( .A(n12831), .B(n12830), .Z(n12835) );
  NANDN U13195 ( .A(n12833), .B(n12832), .Z(n12834) );
  NAND U13196 ( .A(n12835), .B(n12834), .Z(n12880) );
  XOR U13197 ( .A(n12879), .B(n12880), .Z(n12847) );
  OR U13198 ( .A(n12837), .B(n12836), .Z(n12841) );
  NANDN U13199 ( .A(n12839), .B(n12838), .Z(n12840) );
  NAND U13200 ( .A(n12841), .B(n12840), .Z(n12848) );
  XNOR U13201 ( .A(n12847), .B(n12848), .Z(n12849) );
  XNOR U13202 ( .A(n12850), .B(n12849), .Z(n12883) );
  XNOR U13203 ( .A(n12883), .B(sreg[1327]), .Z(n12885) );
  NAND U13204 ( .A(n12842), .B(sreg[1326]), .Z(n12846) );
  OR U13205 ( .A(n12844), .B(n12843), .Z(n12845) );
  AND U13206 ( .A(n12846), .B(n12845), .Z(n12884) );
  XOR U13207 ( .A(n12885), .B(n12884), .Z(c[1327]) );
  NANDN U13208 ( .A(n12848), .B(n12847), .Z(n12852) );
  NAND U13209 ( .A(n12850), .B(n12849), .Z(n12851) );
  NAND U13210 ( .A(n12852), .B(n12851), .Z(n12891) );
  NAND U13211 ( .A(b[0]), .B(a[312]), .Z(n12853) );
  XNOR U13212 ( .A(b[1]), .B(n12853), .Z(n12855) );
  NAND U13213 ( .A(n59), .B(a[311]), .Z(n12854) );
  AND U13214 ( .A(n12855), .B(n12854), .Z(n12908) );
  XOR U13215 ( .A(a[308]), .B(n42197), .Z(n12897) );
  NANDN U13216 ( .A(n12897), .B(n42173), .Z(n12858) );
  NANDN U13217 ( .A(n12856), .B(n42172), .Z(n12857) );
  NAND U13218 ( .A(n12858), .B(n12857), .Z(n12906) );
  NAND U13219 ( .A(b[7]), .B(a[304]), .Z(n12907) );
  XNOR U13220 ( .A(n12906), .B(n12907), .Z(n12909) );
  XOR U13221 ( .A(n12908), .B(n12909), .Z(n12915) );
  NANDN U13222 ( .A(n12859), .B(n42093), .Z(n12861) );
  XOR U13223 ( .A(n42134), .B(a[310]), .Z(n12900) );
  NANDN U13224 ( .A(n12900), .B(n42095), .Z(n12860) );
  NAND U13225 ( .A(n12861), .B(n12860), .Z(n12913) );
  NANDN U13226 ( .A(n12862), .B(n42231), .Z(n12864) );
  XOR U13227 ( .A(n187), .B(a[306]), .Z(n12903) );
  NANDN U13228 ( .A(n12903), .B(n42234), .Z(n12863) );
  AND U13229 ( .A(n12864), .B(n12863), .Z(n12912) );
  XNOR U13230 ( .A(n12913), .B(n12912), .Z(n12914) );
  XNOR U13231 ( .A(n12915), .B(n12914), .Z(n12919) );
  NANDN U13232 ( .A(n12866), .B(n12865), .Z(n12870) );
  NAND U13233 ( .A(n12868), .B(n12867), .Z(n12869) );
  AND U13234 ( .A(n12870), .B(n12869), .Z(n12918) );
  XOR U13235 ( .A(n12919), .B(n12918), .Z(n12920) );
  NANDN U13236 ( .A(n12872), .B(n12871), .Z(n12876) );
  NANDN U13237 ( .A(n12874), .B(n12873), .Z(n12875) );
  NAND U13238 ( .A(n12876), .B(n12875), .Z(n12921) );
  XOR U13239 ( .A(n12920), .B(n12921), .Z(n12888) );
  OR U13240 ( .A(n12878), .B(n12877), .Z(n12882) );
  NANDN U13241 ( .A(n12880), .B(n12879), .Z(n12881) );
  NAND U13242 ( .A(n12882), .B(n12881), .Z(n12889) );
  XNOR U13243 ( .A(n12888), .B(n12889), .Z(n12890) );
  XNOR U13244 ( .A(n12891), .B(n12890), .Z(n12924) );
  XNOR U13245 ( .A(n12924), .B(sreg[1328]), .Z(n12926) );
  NAND U13246 ( .A(n12883), .B(sreg[1327]), .Z(n12887) );
  OR U13247 ( .A(n12885), .B(n12884), .Z(n12886) );
  AND U13248 ( .A(n12887), .B(n12886), .Z(n12925) );
  XOR U13249 ( .A(n12926), .B(n12925), .Z(c[1328]) );
  NANDN U13250 ( .A(n12889), .B(n12888), .Z(n12893) );
  NAND U13251 ( .A(n12891), .B(n12890), .Z(n12892) );
  NAND U13252 ( .A(n12893), .B(n12892), .Z(n12932) );
  NAND U13253 ( .A(b[0]), .B(a[313]), .Z(n12894) );
  XNOR U13254 ( .A(b[1]), .B(n12894), .Z(n12896) );
  NAND U13255 ( .A(n59), .B(a[312]), .Z(n12895) );
  AND U13256 ( .A(n12896), .B(n12895), .Z(n12949) );
  XOR U13257 ( .A(a[309]), .B(n42197), .Z(n12938) );
  NANDN U13258 ( .A(n12938), .B(n42173), .Z(n12899) );
  NANDN U13259 ( .A(n12897), .B(n42172), .Z(n12898) );
  NAND U13260 ( .A(n12899), .B(n12898), .Z(n12947) );
  NAND U13261 ( .A(b[7]), .B(a[305]), .Z(n12948) );
  XNOR U13262 ( .A(n12947), .B(n12948), .Z(n12950) );
  XOR U13263 ( .A(n12949), .B(n12950), .Z(n12956) );
  NANDN U13264 ( .A(n12900), .B(n42093), .Z(n12902) );
  XOR U13265 ( .A(n42134), .B(a[311]), .Z(n12941) );
  NANDN U13266 ( .A(n12941), .B(n42095), .Z(n12901) );
  NAND U13267 ( .A(n12902), .B(n12901), .Z(n12954) );
  NANDN U13268 ( .A(n12903), .B(n42231), .Z(n12905) );
  XOR U13269 ( .A(n187), .B(a[307]), .Z(n12944) );
  NANDN U13270 ( .A(n12944), .B(n42234), .Z(n12904) );
  AND U13271 ( .A(n12905), .B(n12904), .Z(n12953) );
  XNOR U13272 ( .A(n12954), .B(n12953), .Z(n12955) );
  XNOR U13273 ( .A(n12956), .B(n12955), .Z(n12960) );
  NANDN U13274 ( .A(n12907), .B(n12906), .Z(n12911) );
  NAND U13275 ( .A(n12909), .B(n12908), .Z(n12910) );
  AND U13276 ( .A(n12911), .B(n12910), .Z(n12959) );
  XOR U13277 ( .A(n12960), .B(n12959), .Z(n12961) );
  NANDN U13278 ( .A(n12913), .B(n12912), .Z(n12917) );
  NANDN U13279 ( .A(n12915), .B(n12914), .Z(n12916) );
  NAND U13280 ( .A(n12917), .B(n12916), .Z(n12962) );
  XOR U13281 ( .A(n12961), .B(n12962), .Z(n12929) );
  OR U13282 ( .A(n12919), .B(n12918), .Z(n12923) );
  NANDN U13283 ( .A(n12921), .B(n12920), .Z(n12922) );
  NAND U13284 ( .A(n12923), .B(n12922), .Z(n12930) );
  XNOR U13285 ( .A(n12929), .B(n12930), .Z(n12931) );
  XNOR U13286 ( .A(n12932), .B(n12931), .Z(n12965) );
  XNOR U13287 ( .A(n12965), .B(sreg[1329]), .Z(n12967) );
  NAND U13288 ( .A(n12924), .B(sreg[1328]), .Z(n12928) );
  OR U13289 ( .A(n12926), .B(n12925), .Z(n12927) );
  AND U13290 ( .A(n12928), .B(n12927), .Z(n12966) );
  XOR U13291 ( .A(n12967), .B(n12966), .Z(c[1329]) );
  NANDN U13292 ( .A(n12930), .B(n12929), .Z(n12934) );
  NAND U13293 ( .A(n12932), .B(n12931), .Z(n12933) );
  NAND U13294 ( .A(n12934), .B(n12933), .Z(n12973) );
  NAND U13295 ( .A(b[0]), .B(a[314]), .Z(n12935) );
  XNOR U13296 ( .A(b[1]), .B(n12935), .Z(n12937) );
  NAND U13297 ( .A(n59), .B(a[313]), .Z(n12936) );
  AND U13298 ( .A(n12937), .B(n12936), .Z(n12990) );
  XOR U13299 ( .A(a[310]), .B(n42197), .Z(n12979) );
  NANDN U13300 ( .A(n12979), .B(n42173), .Z(n12940) );
  NANDN U13301 ( .A(n12938), .B(n42172), .Z(n12939) );
  NAND U13302 ( .A(n12940), .B(n12939), .Z(n12988) );
  NAND U13303 ( .A(b[7]), .B(a[306]), .Z(n12989) );
  XNOR U13304 ( .A(n12988), .B(n12989), .Z(n12991) );
  XOR U13305 ( .A(n12990), .B(n12991), .Z(n12997) );
  NANDN U13306 ( .A(n12941), .B(n42093), .Z(n12943) );
  XOR U13307 ( .A(n42134), .B(a[312]), .Z(n12982) );
  NANDN U13308 ( .A(n12982), .B(n42095), .Z(n12942) );
  NAND U13309 ( .A(n12943), .B(n12942), .Z(n12995) );
  NANDN U13310 ( .A(n12944), .B(n42231), .Z(n12946) );
  XOR U13311 ( .A(n187), .B(a[308]), .Z(n12985) );
  NANDN U13312 ( .A(n12985), .B(n42234), .Z(n12945) );
  AND U13313 ( .A(n12946), .B(n12945), .Z(n12994) );
  XNOR U13314 ( .A(n12995), .B(n12994), .Z(n12996) );
  XNOR U13315 ( .A(n12997), .B(n12996), .Z(n13001) );
  NANDN U13316 ( .A(n12948), .B(n12947), .Z(n12952) );
  NAND U13317 ( .A(n12950), .B(n12949), .Z(n12951) );
  AND U13318 ( .A(n12952), .B(n12951), .Z(n13000) );
  XOR U13319 ( .A(n13001), .B(n13000), .Z(n13002) );
  NANDN U13320 ( .A(n12954), .B(n12953), .Z(n12958) );
  NANDN U13321 ( .A(n12956), .B(n12955), .Z(n12957) );
  NAND U13322 ( .A(n12958), .B(n12957), .Z(n13003) );
  XOR U13323 ( .A(n13002), .B(n13003), .Z(n12970) );
  OR U13324 ( .A(n12960), .B(n12959), .Z(n12964) );
  NANDN U13325 ( .A(n12962), .B(n12961), .Z(n12963) );
  NAND U13326 ( .A(n12964), .B(n12963), .Z(n12971) );
  XNOR U13327 ( .A(n12970), .B(n12971), .Z(n12972) );
  XNOR U13328 ( .A(n12973), .B(n12972), .Z(n13006) );
  XNOR U13329 ( .A(n13006), .B(sreg[1330]), .Z(n13008) );
  NAND U13330 ( .A(n12965), .B(sreg[1329]), .Z(n12969) );
  OR U13331 ( .A(n12967), .B(n12966), .Z(n12968) );
  AND U13332 ( .A(n12969), .B(n12968), .Z(n13007) );
  XOR U13333 ( .A(n13008), .B(n13007), .Z(c[1330]) );
  NANDN U13334 ( .A(n12971), .B(n12970), .Z(n12975) );
  NAND U13335 ( .A(n12973), .B(n12972), .Z(n12974) );
  NAND U13336 ( .A(n12975), .B(n12974), .Z(n13014) );
  NAND U13337 ( .A(b[0]), .B(a[315]), .Z(n12976) );
  XNOR U13338 ( .A(b[1]), .B(n12976), .Z(n12978) );
  NAND U13339 ( .A(n60), .B(a[314]), .Z(n12977) );
  AND U13340 ( .A(n12978), .B(n12977), .Z(n13031) );
  XOR U13341 ( .A(a[311]), .B(n42197), .Z(n13020) );
  NANDN U13342 ( .A(n13020), .B(n42173), .Z(n12981) );
  NANDN U13343 ( .A(n12979), .B(n42172), .Z(n12980) );
  NAND U13344 ( .A(n12981), .B(n12980), .Z(n13029) );
  NAND U13345 ( .A(b[7]), .B(a[307]), .Z(n13030) );
  XNOR U13346 ( .A(n13029), .B(n13030), .Z(n13032) );
  XOR U13347 ( .A(n13031), .B(n13032), .Z(n13038) );
  NANDN U13348 ( .A(n12982), .B(n42093), .Z(n12984) );
  XOR U13349 ( .A(n42134), .B(a[313]), .Z(n13023) );
  NANDN U13350 ( .A(n13023), .B(n42095), .Z(n12983) );
  NAND U13351 ( .A(n12984), .B(n12983), .Z(n13036) );
  NANDN U13352 ( .A(n12985), .B(n42231), .Z(n12987) );
  XOR U13353 ( .A(n187), .B(a[309]), .Z(n13026) );
  NANDN U13354 ( .A(n13026), .B(n42234), .Z(n12986) );
  AND U13355 ( .A(n12987), .B(n12986), .Z(n13035) );
  XNOR U13356 ( .A(n13036), .B(n13035), .Z(n13037) );
  XNOR U13357 ( .A(n13038), .B(n13037), .Z(n13042) );
  NANDN U13358 ( .A(n12989), .B(n12988), .Z(n12993) );
  NAND U13359 ( .A(n12991), .B(n12990), .Z(n12992) );
  AND U13360 ( .A(n12993), .B(n12992), .Z(n13041) );
  XOR U13361 ( .A(n13042), .B(n13041), .Z(n13043) );
  NANDN U13362 ( .A(n12995), .B(n12994), .Z(n12999) );
  NANDN U13363 ( .A(n12997), .B(n12996), .Z(n12998) );
  NAND U13364 ( .A(n12999), .B(n12998), .Z(n13044) );
  XOR U13365 ( .A(n13043), .B(n13044), .Z(n13011) );
  OR U13366 ( .A(n13001), .B(n13000), .Z(n13005) );
  NANDN U13367 ( .A(n13003), .B(n13002), .Z(n13004) );
  NAND U13368 ( .A(n13005), .B(n13004), .Z(n13012) );
  XNOR U13369 ( .A(n13011), .B(n13012), .Z(n13013) );
  XNOR U13370 ( .A(n13014), .B(n13013), .Z(n13047) );
  XNOR U13371 ( .A(n13047), .B(sreg[1331]), .Z(n13049) );
  NAND U13372 ( .A(n13006), .B(sreg[1330]), .Z(n13010) );
  OR U13373 ( .A(n13008), .B(n13007), .Z(n13009) );
  AND U13374 ( .A(n13010), .B(n13009), .Z(n13048) );
  XOR U13375 ( .A(n13049), .B(n13048), .Z(c[1331]) );
  NANDN U13376 ( .A(n13012), .B(n13011), .Z(n13016) );
  NAND U13377 ( .A(n13014), .B(n13013), .Z(n13015) );
  NAND U13378 ( .A(n13016), .B(n13015), .Z(n13055) );
  NAND U13379 ( .A(b[0]), .B(a[316]), .Z(n13017) );
  XNOR U13380 ( .A(b[1]), .B(n13017), .Z(n13019) );
  NAND U13381 ( .A(n60), .B(a[315]), .Z(n13018) );
  AND U13382 ( .A(n13019), .B(n13018), .Z(n13072) );
  XOR U13383 ( .A(a[312]), .B(n42197), .Z(n13061) );
  NANDN U13384 ( .A(n13061), .B(n42173), .Z(n13022) );
  NANDN U13385 ( .A(n13020), .B(n42172), .Z(n13021) );
  NAND U13386 ( .A(n13022), .B(n13021), .Z(n13070) );
  NAND U13387 ( .A(b[7]), .B(a[308]), .Z(n13071) );
  XNOR U13388 ( .A(n13070), .B(n13071), .Z(n13073) );
  XOR U13389 ( .A(n13072), .B(n13073), .Z(n13079) );
  NANDN U13390 ( .A(n13023), .B(n42093), .Z(n13025) );
  XOR U13391 ( .A(n42134), .B(a[314]), .Z(n13064) );
  NANDN U13392 ( .A(n13064), .B(n42095), .Z(n13024) );
  NAND U13393 ( .A(n13025), .B(n13024), .Z(n13077) );
  NANDN U13394 ( .A(n13026), .B(n42231), .Z(n13028) );
  XOR U13395 ( .A(n187), .B(a[310]), .Z(n13067) );
  NANDN U13396 ( .A(n13067), .B(n42234), .Z(n13027) );
  AND U13397 ( .A(n13028), .B(n13027), .Z(n13076) );
  XNOR U13398 ( .A(n13077), .B(n13076), .Z(n13078) );
  XNOR U13399 ( .A(n13079), .B(n13078), .Z(n13083) );
  NANDN U13400 ( .A(n13030), .B(n13029), .Z(n13034) );
  NAND U13401 ( .A(n13032), .B(n13031), .Z(n13033) );
  AND U13402 ( .A(n13034), .B(n13033), .Z(n13082) );
  XOR U13403 ( .A(n13083), .B(n13082), .Z(n13084) );
  NANDN U13404 ( .A(n13036), .B(n13035), .Z(n13040) );
  NANDN U13405 ( .A(n13038), .B(n13037), .Z(n13039) );
  NAND U13406 ( .A(n13040), .B(n13039), .Z(n13085) );
  XOR U13407 ( .A(n13084), .B(n13085), .Z(n13052) );
  OR U13408 ( .A(n13042), .B(n13041), .Z(n13046) );
  NANDN U13409 ( .A(n13044), .B(n13043), .Z(n13045) );
  NAND U13410 ( .A(n13046), .B(n13045), .Z(n13053) );
  XNOR U13411 ( .A(n13052), .B(n13053), .Z(n13054) );
  XNOR U13412 ( .A(n13055), .B(n13054), .Z(n13088) );
  XNOR U13413 ( .A(n13088), .B(sreg[1332]), .Z(n13090) );
  NAND U13414 ( .A(n13047), .B(sreg[1331]), .Z(n13051) );
  OR U13415 ( .A(n13049), .B(n13048), .Z(n13050) );
  AND U13416 ( .A(n13051), .B(n13050), .Z(n13089) );
  XOR U13417 ( .A(n13090), .B(n13089), .Z(c[1332]) );
  NANDN U13418 ( .A(n13053), .B(n13052), .Z(n13057) );
  NAND U13419 ( .A(n13055), .B(n13054), .Z(n13056) );
  NAND U13420 ( .A(n13057), .B(n13056), .Z(n13096) );
  NAND U13421 ( .A(b[0]), .B(a[317]), .Z(n13058) );
  XNOR U13422 ( .A(b[1]), .B(n13058), .Z(n13060) );
  NAND U13423 ( .A(n60), .B(a[316]), .Z(n13059) );
  AND U13424 ( .A(n13060), .B(n13059), .Z(n13113) );
  XOR U13425 ( .A(a[313]), .B(n42197), .Z(n13102) );
  NANDN U13426 ( .A(n13102), .B(n42173), .Z(n13063) );
  NANDN U13427 ( .A(n13061), .B(n42172), .Z(n13062) );
  NAND U13428 ( .A(n13063), .B(n13062), .Z(n13111) );
  NAND U13429 ( .A(b[7]), .B(a[309]), .Z(n13112) );
  XNOR U13430 ( .A(n13111), .B(n13112), .Z(n13114) );
  XOR U13431 ( .A(n13113), .B(n13114), .Z(n13120) );
  NANDN U13432 ( .A(n13064), .B(n42093), .Z(n13066) );
  XOR U13433 ( .A(n42134), .B(a[315]), .Z(n13105) );
  NANDN U13434 ( .A(n13105), .B(n42095), .Z(n13065) );
  NAND U13435 ( .A(n13066), .B(n13065), .Z(n13118) );
  NANDN U13436 ( .A(n13067), .B(n42231), .Z(n13069) );
  XOR U13437 ( .A(n188), .B(a[311]), .Z(n13108) );
  NANDN U13438 ( .A(n13108), .B(n42234), .Z(n13068) );
  AND U13439 ( .A(n13069), .B(n13068), .Z(n13117) );
  XNOR U13440 ( .A(n13118), .B(n13117), .Z(n13119) );
  XNOR U13441 ( .A(n13120), .B(n13119), .Z(n13124) );
  NANDN U13442 ( .A(n13071), .B(n13070), .Z(n13075) );
  NAND U13443 ( .A(n13073), .B(n13072), .Z(n13074) );
  AND U13444 ( .A(n13075), .B(n13074), .Z(n13123) );
  XOR U13445 ( .A(n13124), .B(n13123), .Z(n13125) );
  NANDN U13446 ( .A(n13077), .B(n13076), .Z(n13081) );
  NANDN U13447 ( .A(n13079), .B(n13078), .Z(n13080) );
  NAND U13448 ( .A(n13081), .B(n13080), .Z(n13126) );
  XOR U13449 ( .A(n13125), .B(n13126), .Z(n13093) );
  OR U13450 ( .A(n13083), .B(n13082), .Z(n13087) );
  NANDN U13451 ( .A(n13085), .B(n13084), .Z(n13086) );
  NAND U13452 ( .A(n13087), .B(n13086), .Z(n13094) );
  XNOR U13453 ( .A(n13093), .B(n13094), .Z(n13095) );
  XNOR U13454 ( .A(n13096), .B(n13095), .Z(n13129) );
  XNOR U13455 ( .A(n13129), .B(sreg[1333]), .Z(n13131) );
  NAND U13456 ( .A(n13088), .B(sreg[1332]), .Z(n13092) );
  OR U13457 ( .A(n13090), .B(n13089), .Z(n13091) );
  AND U13458 ( .A(n13092), .B(n13091), .Z(n13130) );
  XOR U13459 ( .A(n13131), .B(n13130), .Z(c[1333]) );
  NANDN U13460 ( .A(n13094), .B(n13093), .Z(n13098) );
  NAND U13461 ( .A(n13096), .B(n13095), .Z(n13097) );
  NAND U13462 ( .A(n13098), .B(n13097), .Z(n13137) );
  NAND U13463 ( .A(b[0]), .B(a[318]), .Z(n13099) );
  XNOR U13464 ( .A(b[1]), .B(n13099), .Z(n13101) );
  NAND U13465 ( .A(n60), .B(a[317]), .Z(n13100) );
  AND U13466 ( .A(n13101), .B(n13100), .Z(n13154) );
  XOR U13467 ( .A(a[314]), .B(n42197), .Z(n13143) );
  NANDN U13468 ( .A(n13143), .B(n42173), .Z(n13104) );
  NANDN U13469 ( .A(n13102), .B(n42172), .Z(n13103) );
  NAND U13470 ( .A(n13104), .B(n13103), .Z(n13152) );
  NAND U13471 ( .A(b[7]), .B(a[310]), .Z(n13153) );
  XNOR U13472 ( .A(n13152), .B(n13153), .Z(n13155) );
  XOR U13473 ( .A(n13154), .B(n13155), .Z(n13161) );
  NANDN U13474 ( .A(n13105), .B(n42093), .Z(n13107) );
  XOR U13475 ( .A(n42134), .B(a[316]), .Z(n13146) );
  NANDN U13476 ( .A(n13146), .B(n42095), .Z(n13106) );
  NAND U13477 ( .A(n13107), .B(n13106), .Z(n13159) );
  NANDN U13478 ( .A(n13108), .B(n42231), .Z(n13110) );
  XOR U13479 ( .A(n188), .B(a[312]), .Z(n13149) );
  NANDN U13480 ( .A(n13149), .B(n42234), .Z(n13109) );
  AND U13481 ( .A(n13110), .B(n13109), .Z(n13158) );
  XNOR U13482 ( .A(n13159), .B(n13158), .Z(n13160) );
  XNOR U13483 ( .A(n13161), .B(n13160), .Z(n13165) );
  NANDN U13484 ( .A(n13112), .B(n13111), .Z(n13116) );
  NAND U13485 ( .A(n13114), .B(n13113), .Z(n13115) );
  AND U13486 ( .A(n13116), .B(n13115), .Z(n13164) );
  XOR U13487 ( .A(n13165), .B(n13164), .Z(n13166) );
  NANDN U13488 ( .A(n13118), .B(n13117), .Z(n13122) );
  NANDN U13489 ( .A(n13120), .B(n13119), .Z(n13121) );
  NAND U13490 ( .A(n13122), .B(n13121), .Z(n13167) );
  XOR U13491 ( .A(n13166), .B(n13167), .Z(n13134) );
  OR U13492 ( .A(n13124), .B(n13123), .Z(n13128) );
  NANDN U13493 ( .A(n13126), .B(n13125), .Z(n13127) );
  NAND U13494 ( .A(n13128), .B(n13127), .Z(n13135) );
  XNOR U13495 ( .A(n13134), .B(n13135), .Z(n13136) );
  XNOR U13496 ( .A(n13137), .B(n13136), .Z(n13170) );
  XNOR U13497 ( .A(n13170), .B(sreg[1334]), .Z(n13172) );
  NAND U13498 ( .A(n13129), .B(sreg[1333]), .Z(n13133) );
  OR U13499 ( .A(n13131), .B(n13130), .Z(n13132) );
  AND U13500 ( .A(n13133), .B(n13132), .Z(n13171) );
  XOR U13501 ( .A(n13172), .B(n13171), .Z(c[1334]) );
  NANDN U13502 ( .A(n13135), .B(n13134), .Z(n13139) );
  NAND U13503 ( .A(n13137), .B(n13136), .Z(n13138) );
  NAND U13504 ( .A(n13139), .B(n13138), .Z(n13178) );
  NAND U13505 ( .A(b[0]), .B(a[319]), .Z(n13140) );
  XNOR U13506 ( .A(b[1]), .B(n13140), .Z(n13142) );
  NAND U13507 ( .A(n60), .B(a[318]), .Z(n13141) );
  AND U13508 ( .A(n13142), .B(n13141), .Z(n13195) );
  XOR U13509 ( .A(a[315]), .B(n42197), .Z(n13184) );
  NANDN U13510 ( .A(n13184), .B(n42173), .Z(n13145) );
  NANDN U13511 ( .A(n13143), .B(n42172), .Z(n13144) );
  NAND U13512 ( .A(n13145), .B(n13144), .Z(n13193) );
  NAND U13513 ( .A(b[7]), .B(a[311]), .Z(n13194) );
  XNOR U13514 ( .A(n13193), .B(n13194), .Z(n13196) );
  XOR U13515 ( .A(n13195), .B(n13196), .Z(n13202) );
  NANDN U13516 ( .A(n13146), .B(n42093), .Z(n13148) );
  XOR U13517 ( .A(n42134), .B(a[317]), .Z(n13187) );
  NANDN U13518 ( .A(n13187), .B(n42095), .Z(n13147) );
  NAND U13519 ( .A(n13148), .B(n13147), .Z(n13200) );
  NANDN U13520 ( .A(n13149), .B(n42231), .Z(n13151) );
  XOR U13521 ( .A(n188), .B(a[313]), .Z(n13190) );
  NANDN U13522 ( .A(n13190), .B(n42234), .Z(n13150) );
  AND U13523 ( .A(n13151), .B(n13150), .Z(n13199) );
  XNOR U13524 ( .A(n13200), .B(n13199), .Z(n13201) );
  XNOR U13525 ( .A(n13202), .B(n13201), .Z(n13206) );
  NANDN U13526 ( .A(n13153), .B(n13152), .Z(n13157) );
  NAND U13527 ( .A(n13155), .B(n13154), .Z(n13156) );
  AND U13528 ( .A(n13157), .B(n13156), .Z(n13205) );
  XOR U13529 ( .A(n13206), .B(n13205), .Z(n13207) );
  NANDN U13530 ( .A(n13159), .B(n13158), .Z(n13163) );
  NANDN U13531 ( .A(n13161), .B(n13160), .Z(n13162) );
  NAND U13532 ( .A(n13163), .B(n13162), .Z(n13208) );
  XOR U13533 ( .A(n13207), .B(n13208), .Z(n13175) );
  OR U13534 ( .A(n13165), .B(n13164), .Z(n13169) );
  NANDN U13535 ( .A(n13167), .B(n13166), .Z(n13168) );
  NAND U13536 ( .A(n13169), .B(n13168), .Z(n13176) );
  XNOR U13537 ( .A(n13175), .B(n13176), .Z(n13177) );
  XNOR U13538 ( .A(n13178), .B(n13177), .Z(n13211) );
  XNOR U13539 ( .A(n13211), .B(sreg[1335]), .Z(n13213) );
  NAND U13540 ( .A(n13170), .B(sreg[1334]), .Z(n13174) );
  OR U13541 ( .A(n13172), .B(n13171), .Z(n13173) );
  AND U13542 ( .A(n13174), .B(n13173), .Z(n13212) );
  XOR U13543 ( .A(n13213), .B(n13212), .Z(c[1335]) );
  NANDN U13544 ( .A(n13176), .B(n13175), .Z(n13180) );
  NAND U13545 ( .A(n13178), .B(n13177), .Z(n13179) );
  NAND U13546 ( .A(n13180), .B(n13179), .Z(n13219) );
  NAND U13547 ( .A(b[0]), .B(a[320]), .Z(n13181) );
  XNOR U13548 ( .A(b[1]), .B(n13181), .Z(n13183) );
  NAND U13549 ( .A(n60), .B(a[319]), .Z(n13182) );
  AND U13550 ( .A(n13183), .B(n13182), .Z(n13236) );
  XOR U13551 ( .A(a[316]), .B(n42197), .Z(n13225) );
  NANDN U13552 ( .A(n13225), .B(n42173), .Z(n13186) );
  NANDN U13553 ( .A(n13184), .B(n42172), .Z(n13185) );
  NAND U13554 ( .A(n13186), .B(n13185), .Z(n13234) );
  NAND U13555 ( .A(b[7]), .B(a[312]), .Z(n13235) );
  XNOR U13556 ( .A(n13234), .B(n13235), .Z(n13237) );
  XOR U13557 ( .A(n13236), .B(n13237), .Z(n13243) );
  NANDN U13558 ( .A(n13187), .B(n42093), .Z(n13189) );
  XOR U13559 ( .A(n42134), .B(a[318]), .Z(n13228) );
  NANDN U13560 ( .A(n13228), .B(n42095), .Z(n13188) );
  NAND U13561 ( .A(n13189), .B(n13188), .Z(n13241) );
  NANDN U13562 ( .A(n13190), .B(n42231), .Z(n13192) );
  XOR U13563 ( .A(n188), .B(a[314]), .Z(n13231) );
  NANDN U13564 ( .A(n13231), .B(n42234), .Z(n13191) );
  AND U13565 ( .A(n13192), .B(n13191), .Z(n13240) );
  XNOR U13566 ( .A(n13241), .B(n13240), .Z(n13242) );
  XNOR U13567 ( .A(n13243), .B(n13242), .Z(n13247) );
  NANDN U13568 ( .A(n13194), .B(n13193), .Z(n13198) );
  NAND U13569 ( .A(n13196), .B(n13195), .Z(n13197) );
  AND U13570 ( .A(n13198), .B(n13197), .Z(n13246) );
  XOR U13571 ( .A(n13247), .B(n13246), .Z(n13248) );
  NANDN U13572 ( .A(n13200), .B(n13199), .Z(n13204) );
  NANDN U13573 ( .A(n13202), .B(n13201), .Z(n13203) );
  NAND U13574 ( .A(n13204), .B(n13203), .Z(n13249) );
  XOR U13575 ( .A(n13248), .B(n13249), .Z(n13216) );
  OR U13576 ( .A(n13206), .B(n13205), .Z(n13210) );
  NANDN U13577 ( .A(n13208), .B(n13207), .Z(n13209) );
  NAND U13578 ( .A(n13210), .B(n13209), .Z(n13217) );
  XNOR U13579 ( .A(n13216), .B(n13217), .Z(n13218) );
  XNOR U13580 ( .A(n13219), .B(n13218), .Z(n13252) );
  XNOR U13581 ( .A(n13252), .B(sreg[1336]), .Z(n13254) );
  NAND U13582 ( .A(n13211), .B(sreg[1335]), .Z(n13215) );
  OR U13583 ( .A(n13213), .B(n13212), .Z(n13214) );
  AND U13584 ( .A(n13215), .B(n13214), .Z(n13253) );
  XOR U13585 ( .A(n13254), .B(n13253), .Z(c[1336]) );
  NANDN U13586 ( .A(n13217), .B(n13216), .Z(n13221) );
  NAND U13587 ( .A(n13219), .B(n13218), .Z(n13220) );
  NAND U13588 ( .A(n13221), .B(n13220), .Z(n13260) );
  NAND U13589 ( .A(b[0]), .B(a[321]), .Z(n13222) );
  XNOR U13590 ( .A(b[1]), .B(n13222), .Z(n13224) );
  NAND U13591 ( .A(n60), .B(a[320]), .Z(n13223) );
  AND U13592 ( .A(n13224), .B(n13223), .Z(n13277) );
  XOR U13593 ( .A(a[317]), .B(n42197), .Z(n13266) );
  NANDN U13594 ( .A(n13266), .B(n42173), .Z(n13227) );
  NANDN U13595 ( .A(n13225), .B(n42172), .Z(n13226) );
  NAND U13596 ( .A(n13227), .B(n13226), .Z(n13275) );
  NAND U13597 ( .A(b[7]), .B(a[313]), .Z(n13276) );
  XNOR U13598 ( .A(n13275), .B(n13276), .Z(n13278) );
  XOR U13599 ( .A(n13277), .B(n13278), .Z(n13284) );
  NANDN U13600 ( .A(n13228), .B(n42093), .Z(n13230) );
  XOR U13601 ( .A(n42134), .B(a[319]), .Z(n13269) );
  NANDN U13602 ( .A(n13269), .B(n42095), .Z(n13229) );
  NAND U13603 ( .A(n13230), .B(n13229), .Z(n13282) );
  NANDN U13604 ( .A(n13231), .B(n42231), .Z(n13233) );
  XOR U13605 ( .A(n188), .B(a[315]), .Z(n13272) );
  NANDN U13606 ( .A(n13272), .B(n42234), .Z(n13232) );
  AND U13607 ( .A(n13233), .B(n13232), .Z(n13281) );
  XNOR U13608 ( .A(n13282), .B(n13281), .Z(n13283) );
  XNOR U13609 ( .A(n13284), .B(n13283), .Z(n13288) );
  NANDN U13610 ( .A(n13235), .B(n13234), .Z(n13239) );
  NAND U13611 ( .A(n13237), .B(n13236), .Z(n13238) );
  AND U13612 ( .A(n13239), .B(n13238), .Z(n13287) );
  XOR U13613 ( .A(n13288), .B(n13287), .Z(n13289) );
  NANDN U13614 ( .A(n13241), .B(n13240), .Z(n13245) );
  NANDN U13615 ( .A(n13243), .B(n13242), .Z(n13244) );
  NAND U13616 ( .A(n13245), .B(n13244), .Z(n13290) );
  XOR U13617 ( .A(n13289), .B(n13290), .Z(n13257) );
  OR U13618 ( .A(n13247), .B(n13246), .Z(n13251) );
  NANDN U13619 ( .A(n13249), .B(n13248), .Z(n13250) );
  NAND U13620 ( .A(n13251), .B(n13250), .Z(n13258) );
  XNOR U13621 ( .A(n13257), .B(n13258), .Z(n13259) );
  XNOR U13622 ( .A(n13260), .B(n13259), .Z(n13293) );
  XNOR U13623 ( .A(n13293), .B(sreg[1337]), .Z(n13295) );
  NAND U13624 ( .A(n13252), .B(sreg[1336]), .Z(n13256) );
  OR U13625 ( .A(n13254), .B(n13253), .Z(n13255) );
  AND U13626 ( .A(n13256), .B(n13255), .Z(n13294) );
  XOR U13627 ( .A(n13295), .B(n13294), .Z(c[1337]) );
  NANDN U13628 ( .A(n13258), .B(n13257), .Z(n13262) );
  NAND U13629 ( .A(n13260), .B(n13259), .Z(n13261) );
  NAND U13630 ( .A(n13262), .B(n13261), .Z(n13301) );
  NAND U13631 ( .A(b[0]), .B(a[322]), .Z(n13263) );
  XNOR U13632 ( .A(b[1]), .B(n13263), .Z(n13265) );
  NAND U13633 ( .A(n61), .B(a[321]), .Z(n13264) );
  AND U13634 ( .A(n13265), .B(n13264), .Z(n13318) );
  XOR U13635 ( .A(a[318]), .B(n42197), .Z(n13307) );
  NANDN U13636 ( .A(n13307), .B(n42173), .Z(n13268) );
  NANDN U13637 ( .A(n13266), .B(n42172), .Z(n13267) );
  NAND U13638 ( .A(n13268), .B(n13267), .Z(n13316) );
  NAND U13639 ( .A(b[7]), .B(a[314]), .Z(n13317) );
  XNOR U13640 ( .A(n13316), .B(n13317), .Z(n13319) );
  XOR U13641 ( .A(n13318), .B(n13319), .Z(n13325) );
  NANDN U13642 ( .A(n13269), .B(n42093), .Z(n13271) );
  XOR U13643 ( .A(n42134), .B(a[320]), .Z(n13310) );
  NANDN U13644 ( .A(n13310), .B(n42095), .Z(n13270) );
  NAND U13645 ( .A(n13271), .B(n13270), .Z(n13323) );
  NANDN U13646 ( .A(n13272), .B(n42231), .Z(n13274) );
  XOR U13647 ( .A(n188), .B(a[316]), .Z(n13313) );
  NANDN U13648 ( .A(n13313), .B(n42234), .Z(n13273) );
  AND U13649 ( .A(n13274), .B(n13273), .Z(n13322) );
  XNOR U13650 ( .A(n13323), .B(n13322), .Z(n13324) );
  XNOR U13651 ( .A(n13325), .B(n13324), .Z(n13329) );
  NANDN U13652 ( .A(n13276), .B(n13275), .Z(n13280) );
  NAND U13653 ( .A(n13278), .B(n13277), .Z(n13279) );
  AND U13654 ( .A(n13280), .B(n13279), .Z(n13328) );
  XOR U13655 ( .A(n13329), .B(n13328), .Z(n13330) );
  NANDN U13656 ( .A(n13282), .B(n13281), .Z(n13286) );
  NANDN U13657 ( .A(n13284), .B(n13283), .Z(n13285) );
  NAND U13658 ( .A(n13286), .B(n13285), .Z(n13331) );
  XOR U13659 ( .A(n13330), .B(n13331), .Z(n13298) );
  OR U13660 ( .A(n13288), .B(n13287), .Z(n13292) );
  NANDN U13661 ( .A(n13290), .B(n13289), .Z(n13291) );
  NAND U13662 ( .A(n13292), .B(n13291), .Z(n13299) );
  XNOR U13663 ( .A(n13298), .B(n13299), .Z(n13300) );
  XNOR U13664 ( .A(n13301), .B(n13300), .Z(n13334) );
  XNOR U13665 ( .A(n13334), .B(sreg[1338]), .Z(n13336) );
  NAND U13666 ( .A(n13293), .B(sreg[1337]), .Z(n13297) );
  OR U13667 ( .A(n13295), .B(n13294), .Z(n13296) );
  AND U13668 ( .A(n13297), .B(n13296), .Z(n13335) );
  XOR U13669 ( .A(n13336), .B(n13335), .Z(c[1338]) );
  NANDN U13670 ( .A(n13299), .B(n13298), .Z(n13303) );
  NAND U13671 ( .A(n13301), .B(n13300), .Z(n13302) );
  NAND U13672 ( .A(n13303), .B(n13302), .Z(n13342) );
  NAND U13673 ( .A(b[0]), .B(a[323]), .Z(n13304) );
  XNOR U13674 ( .A(b[1]), .B(n13304), .Z(n13306) );
  NAND U13675 ( .A(n61), .B(a[322]), .Z(n13305) );
  AND U13676 ( .A(n13306), .B(n13305), .Z(n13359) );
  XOR U13677 ( .A(a[319]), .B(n42197), .Z(n13348) );
  NANDN U13678 ( .A(n13348), .B(n42173), .Z(n13309) );
  NANDN U13679 ( .A(n13307), .B(n42172), .Z(n13308) );
  NAND U13680 ( .A(n13309), .B(n13308), .Z(n13357) );
  NAND U13681 ( .A(b[7]), .B(a[315]), .Z(n13358) );
  XNOR U13682 ( .A(n13357), .B(n13358), .Z(n13360) );
  XOR U13683 ( .A(n13359), .B(n13360), .Z(n13366) );
  NANDN U13684 ( .A(n13310), .B(n42093), .Z(n13312) );
  XOR U13685 ( .A(n42134), .B(a[321]), .Z(n13351) );
  NANDN U13686 ( .A(n13351), .B(n42095), .Z(n13311) );
  NAND U13687 ( .A(n13312), .B(n13311), .Z(n13364) );
  NANDN U13688 ( .A(n13313), .B(n42231), .Z(n13315) );
  XOR U13689 ( .A(n188), .B(a[317]), .Z(n13354) );
  NANDN U13690 ( .A(n13354), .B(n42234), .Z(n13314) );
  AND U13691 ( .A(n13315), .B(n13314), .Z(n13363) );
  XNOR U13692 ( .A(n13364), .B(n13363), .Z(n13365) );
  XNOR U13693 ( .A(n13366), .B(n13365), .Z(n13370) );
  NANDN U13694 ( .A(n13317), .B(n13316), .Z(n13321) );
  NAND U13695 ( .A(n13319), .B(n13318), .Z(n13320) );
  AND U13696 ( .A(n13321), .B(n13320), .Z(n13369) );
  XOR U13697 ( .A(n13370), .B(n13369), .Z(n13371) );
  NANDN U13698 ( .A(n13323), .B(n13322), .Z(n13327) );
  NANDN U13699 ( .A(n13325), .B(n13324), .Z(n13326) );
  NAND U13700 ( .A(n13327), .B(n13326), .Z(n13372) );
  XOR U13701 ( .A(n13371), .B(n13372), .Z(n13339) );
  OR U13702 ( .A(n13329), .B(n13328), .Z(n13333) );
  NANDN U13703 ( .A(n13331), .B(n13330), .Z(n13332) );
  NAND U13704 ( .A(n13333), .B(n13332), .Z(n13340) );
  XNOR U13705 ( .A(n13339), .B(n13340), .Z(n13341) );
  XNOR U13706 ( .A(n13342), .B(n13341), .Z(n13375) );
  XNOR U13707 ( .A(n13375), .B(sreg[1339]), .Z(n13377) );
  NAND U13708 ( .A(n13334), .B(sreg[1338]), .Z(n13338) );
  OR U13709 ( .A(n13336), .B(n13335), .Z(n13337) );
  AND U13710 ( .A(n13338), .B(n13337), .Z(n13376) );
  XOR U13711 ( .A(n13377), .B(n13376), .Z(c[1339]) );
  NANDN U13712 ( .A(n13340), .B(n13339), .Z(n13344) );
  NAND U13713 ( .A(n13342), .B(n13341), .Z(n13343) );
  NAND U13714 ( .A(n13344), .B(n13343), .Z(n13383) );
  NAND U13715 ( .A(b[0]), .B(a[324]), .Z(n13345) );
  XNOR U13716 ( .A(b[1]), .B(n13345), .Z(n13347) );
  NAND U13717 ( .A(n61), .B(a[323]), .Z(n13346) );
  AND U13718 ( .A(n13347), .B(n13346), .Z(n13400) );
  XOR U13719 ( .A(a[320]), .B(n42197), .Z(n13389) );
  NANDN U13720 ( .A(n13389), .B(n42173), .Z(n13350) );
  NANDN U13721 ( .A(n13348), .B(n42172), .Z(n13349) );
  NAND U13722 ( .A(n13350), .B(n13349), .Z(n13398) );
  NAND U13723 ( .A(b[7]), .B(a[316]), .Z(n13399) );
  XNOR U13724 ( .A(n13398), .B(n13399), .Z(n13401) );
  XOR U13725 ( .A(n13400), .B(n13401), .Z(n13407) );
  NANDN U13726 ( .A(n13351), .B(n42093), .Z(n13353) );
  XOR U13727 ( .A(n42134), .B(a[322]), .Z(n13392) );
  NANDN U13728 ( .A(n13392), .B(n42095), .Z(n13352) );
  NAND U13729 ( .A(n13353), .B(n13352), .Z(n13405) );
  NANDN U13730 ( .A(n13354), .B(n42231), .Z(n13356) );
  XOR U13731 ( .A(n188), .B(a[318]), .Z(n13395) );
  NANDN U13732 ( .A(n13395), .B(n42234), .Z(n13355) );
  AND U13733 ( .A(n13356), .B(n13355), .Z(n13404) );
  XNOR U13734 ( .A(n13405), .B(n13404), .Z(n13406) );
  XNOR U13735 ( .A(n13407), .B(n13406), .Z(n13411) );
  NANDN U13736 ( .A(n13358), .B(n13357), .Z(n13362) );
  NAND U13737 ( .A(n13360), .B(n13359), .Z(n13361) );
  AND U13738 ( .A(n13362), .B(n13361), .Z(n13410) );
  XOR U13739 ( .A(n13411), .B(n13410), .Z(n13412) );
  NANDN U13740 ( .A(n13364), .B(n13363), .Z(n13368) );
  NANDN U13741 ( .A(n13366), .B(n13365), .Z(n13367) );
  NAND U13742 ( .A(n13368), .B(n13367), .Z(n13413) );
  XOR U13743 ( .A(n13412), .B(n13413), .Z(n13380) );
  OR U13744 ( .A(n13370), .B(n13369), .Z(n13374) );
  NANDN U13745 ( .A(n13372), .B(n13371), .Z(n13373) );
  NAND U13746 ( .A(n13374), .B(n13373), .Z(n13381) );
  XNOR U13747 ( .A(n13380), .B(n13381), .Z(n13382) );
  XNOR U13748 ( .A(n13383), .B(n13382), .Z(n13416) );
  XNOR U13749 ( .A(n13416), .B(sreg[1340]), .Z(n13418) );
  NAND U13750 ( .A(n13375), .B(sreg[1339]), .Z(n13379) );
  OR U13751 ( .A(n13377), .B(n13376), .Z(n13378) );
  AND U13752 ( .A(n13379), .B(n13378), .Z(n13417) );
  XOR U13753 ( .A(n13418), .B(n13417), .Z(c[1340]) );
  NANDN U13754 ( .A(n13381), .B(n13380), .Z(n13385) );
  NAND U13755 ( .A(n13383), .B(n13382), .Z(n13384) );
  NAND U13756 ( .A(n13385), .B(n13384), .Z(n13424) );
  NAND U13757 ( .A(b[0]), .B(a[325]), .Z(n13386) );
  XNOR U13758 ( .A(b[1]), .B(n13386), .Z(n13388) );
  NAND U13759 ( .A(n61), .B(a[324]), .Z(n13387) );
  AND U13760 ( .A(n13388), .B(n13387), .Z(n13441) );
  XOR U13761 ( .A(a[321]), .B(n42197), .Z(n13430) );
  NANDN U13762 ( .A(n13430), .B(n42173), .Z(n13391) );
  NANDN U13763 ( .A(n13389), .B(n42172), .Z(n13390) );
  NAND U13764 ( .A(n13391), .B(n13390), .Z(n13439) );
  NAND U13765 ( .A(b[7]), .B(a[317]), .Z(n13440) );
  XNOR U13766 ( .A(n13439), .B(n13440), .Z(n13442) );
  XOR U13767 ( .A(n13441), .B(n13442), .Z(n13448) );
  NANDN U13768 ( .A(n13392), .B(n42093), .Z(n13394) );
  XOR U13769 ( .A(n42134), .B(a[323]), .Z(n13433) );
  NANDN U13770 ( .A(n13433), .B(n42095), .Z(n13393) );
  NAND U13771 ( .A(n13394), .B(n13393), .Z(n13446) );
  NANDN U13772 ( .A(n13395), .B(n42231), .Z(n13397) );
  XOR U13773 ( .A(n188), .B(a[319]), .Z(n13436) );
  NANDN U13774 ( .A(n13436), .B(n42234), .Z(n13396) );
  AND U13775 ( .A(n13397), .B(n13396), .Z(n13445) );
  XNOR U13776 ( .A(n13446), .B(n13445), .Z(n13447) );
  XNOR U13777 ( .A(n13448), .B(n13447), .Z(n13452) );
  NANDN U13778 ( .A(n13399), .B(n13398), .Z(n13403) );
  NAND U13779 ( .A(n13401), .B(n13400), .Z(n13402) );
  AND U13780 ( .A(n13403), .B(n13402), .Z(n13451) );
  XOR U13781 ( .A(n13452), .B(n13451), .Z(n13453) );
  NANDN U13782 ( .A(n13405), .B(n13404), .Z(n13409) );
  NANDN U13783 ( .A(n13407), .B(n13406), .Z(n13408) );
  NAND U13784 ( .A(n13409), .B(n13408), .Z(n13454) );
  XOR U13785 ( .A(n13453), .B(n13454), .Z(n13421) );
  OR U13786 ( .A(n13411), .B(n13410), .Z(n13415) );
  NANDN U13787 ( .A(n13413), .B(n13412), .Z(n13414) );
  NAND U13788 ( .A(n13415), .B(n13414), .Z(n13422) );
  XNOR U13789 ( .A(n13421), .B(n13422), .Z(n13423) );
  XNOR U13790 ( .A(n13424), .B(n13423), .Z(n13457) );
  XNOR U13791 ( .A(n13457), .B(sreg[1341]), .Z(n13459) );
  NAND U13792 ( .A(n13416), .B(sreg[1340]), .Z(n13420) );
  OR U13793 ( .A(n13418), .B(n13417), .Z(n13419) );
  AND U13794 ( .A(n13420), .B(n13419), .Z(n13458) );
  XOR U13795 ( .A(n13459), .B(n13458), .Z(c[1341]) );
  NANDN U13796 ( .A(n13422), .B(n13421), .Z(n13426) );
  NAND U13797 ( .A(n13424), .B(n13423), .Z(n13425) );
  NAND U13798 ( .A(n13426), .B(n13425), .Z(n13465) );
  NAND U13799 ( .A(b[0]), .B(a[326]), .Z(n13427) );
  XNOR U13800 ( .A(b[1]), .B(n13427), .Z(n13429) );
  NAND U13801 ( .A(n61), .B(a[325]), .Z(n13428) );
  AND U13802 ( .A(n13429), .B(n13428), .Z(n13482) );
  XOR U13803 ( .A(a[322]), .B(n42197), .Z(n13471) );
  NANDN U13804 ( .A(n13471), .B(n42173), .Z(n13432) );
  NANDN U13805 ( .A(n13430), .B(n42172), .Z(n13431) );
  NAND U13806 ( .A(n13432), .B(n13431), .Z(n13480) );
  NAND U13807 ( .A(b[7]), .B(a[318]), .Z(n13481) );
  XNOR U13808 ( .A(n13480), .B(n13481), .Z(n13483) );
  XOR U13809 ( .A(n13482), .B(n13483), .Z(n13489) );
  NANDN U13810 ( .A(n13433), .B(n42093), .Z(n13435) );
  XOR U13811 ( .A(n42134), .B(a[324]), .Z(n13474) );
  NANDN U13812 ( .A(n13474), .B(n42095), .Z(n13434) );
  NAND U13813 ( .A(n13435), .B(n13434), .Z(n13487) );
  NANDN U13814 ( .A(n13436), .B(n42231), .Z(n13438) );
  XOR U13815 ( .A(n188), .B(a[320]), .Z(n13477) );
  NANDN U13816 ( .A(n13477), .B(n42234), .Z(n13437) );
  AND U13817 ( .A(n13438), .B(n13437), .Z(n13486) );
  XNOR U13818 ( .A(n13487), .B(n13486), .Z(n13488) );
  XNOR U13819 ( .A(n13489), .B(n13488), .Z(n13493) );
  NANDN U13820 ( .A(n13440), .B(n13439), .Z(n13444) );
  NAND U13821 ( .A(n13442), .B(n13441), .Z(n13443) );
  AND U13822 ( .A(n13444), .B(n13443), .Z(n13492) );
  XOR U13823 ( .A(n13493), .B(n13492), .Z(n13494) );
  NANDN U13824 ( .A(n13446), .B(n13445), .Z(n13450) );
  NANDN U13825 ( .A(n13448), .B(n13447), .Z(n13449) );
  NAND U13826 ( .A(n13450), .B(n13449), .Z(n13495) );
  XOR U13827 ( .A(n13494), .B(n13495), .Z(n13462) );
  OR U13828 ( .A(n13452), .B(n13451), .Z(n13456) );
  NANDN U13829 ( .A(n13454), .B(n13453), .Z(n13455) );
  NAND U13830 ( .A(n13456), .B(n13455), .Z(n13463) );
  XNOR U13831 ( .A(n13462), .B(n13463), .Z(n13464) );
  XNOR U13832 ( .A(n13465), .B(n13464), .Z(n13498) );
  XNOR U13833 ( .A(n13498), .B(sreg[1342]), .Z(n13500) );
  NAND U13834 ( .A(n13457), .B(sreg[1341]), .Z(n13461) );
  OR U13835 ( .A(n13459), .B(n13458), .Z(n13460) );
  AND U13836 ( .A(n13461), .B(n13460), .Z(n13499) );
  XOR U13837 ( .A(n13500), .B(n13499), .Z(c[1342]) );
  NANDN U13838 ( .A(n13463), .B(n13462), .Z(n13467) );
  NAND U13839 ( .A(n13465), .B(n13464), .Z(n13466) );
  NAND U13840 ( .A(n13467), .B(n13466), .Z(n13506) );
  NAND U13841 ( .A(b[0]), .B(a[327]), .Z(n13468) );
  XNOR U13842 ( .A(b[1]), .B(n13468), .Z(n13470) );
  NAND U13843 ( .A(n61), .B(a[326]), .Z(n13469) );
  AND U13844 ( .A(n13470), .B(n13469), .Z(n13523) );
  XOR U13845 ( .A(a[323]), .B(n42197), .Z(n13512) );
  NANDN U13846 ( .A(n13512), .B(n42173), .Z(n13473) );
  NANDN U13847 ( .A(n13471), .B(n42172), .Z(n13472) );
  NAND U13848 ( .A(n13473), .B(n13472), .Z(n13521) );
  NAND U13849 ( .A(b[7]), .B(a[319]), .Z(n13522) );
  XNOR U13850 ( .A(n13521), .B(n13522), .Z(n13524) );
  XOR U13851 ( .A(n13523), .B(n13524), .Z(n13530) );
  NANDN U13852 ( .A(n13474), .B(n42093), .Z(n13476) );
  XOR U13853 ( .A(n42134), .B(a[325]), .Z(n13515) );
  NANDN U13854 ( .A(n13515), .B(n42095), .Z(n13475) );
  NAND U13855 ( .A(n13476), .B(n13475), .Z(n13528) );
  NANDN U13856 ( .A(n13477), .B(n42231), .Z(n13479) );
  XOR U13857 ( .A(n188), .B(a[321]), .Z(n13518) );
  NANDN U13858 ( .A(n13518), .B(n42234), .Z(n13478) );
  AND U13859 ( .A(n13479), .B(n13478), .Z(n13527) );
  XNOR U13860 ( .A(n13528), .B(n13527), .Z(n13529) );
  XNOR U13861 ( .A(n13530), .B(n13529), .Z(n13534) );
  NANDN U13862 ( .A(n13481), .B(n13480), .Z(n13485) );
  NAND U13863 ( .A(n13483), .B(n13482), .Z(n13484) );
  AND U13864 ( .A(n13485), .B(n13484), .Z(n13533) );
  XOR U13865 ( .A(n13534), .B(n13533), .Z(n13535) );
  NANDN U13866 ( .A(n13487), .B(n13486), .Z(n13491) );
  NANDN U13867 ( .A(n13489), .B(n13488), .Z(n13490) );
  NAND U13868 ( .A(n13491), .B(n13490), .Z(n13536) );
  XOR U13869 ( .A(n13535), .B(n13536), .Z(n13503) );
  OR U13870 ( .A(n13493), .B(n13492), .Z(n13497) );
  NANDN U13871 ( .A(n13495), .B(n13494), .Z(n13496) );
  NAND U13872 ( .A(n13497), .B(n13496), .Z(n13504) );
  XNOR U13873 ( .A(n13503), .B(n13504), .Z(n13505) );
  XNOR U13874 ( .A(n13506), .B(n13505), .Z(n13539) );
  XNOR U13875 ( .A(n13539), .B(sreg[1343]), .Z(n13541) );
  NAND U13876 ( .A(n13498), .B(sreg[1342]), .Z(n13502) );
  OR U13877 ( .A(n13500), .B(n13499), .Z(n13501) );
  AND U13878 ( .A(n13502), .B(n13501), .Z(n13540) );
  XOR U13879 ( .A(n13541), .B(n13540), .Z(c[1343]) );
  NANDN U13880 ( .A(n13504), .B(n13503), .Z(n13508) );
  NAND U13881 ( .A(n13506), .B(n13505), .Z(n13507) );
  NAND U13882 ( .A(n13508), .B(n13507), .Z(n13547) );
  NAND U13883 ( .A(b[0]), .B(a[328]), .Z(n13509) );
  XNOR U13884 ( .A(b[1]), .B(n13509), .Z(n13511) );
  NAND U13885 ( .A(n61), .B(a[327]), .Z(n13510) );
  AND U13886 ( .A(n13511), .B(n13510), .Z(n13564) );
  XOR U13887 ( .A(a[324]), .B(n42197), .Z(n13553) );
  NANDN U13888 ( .A(n13553), .B(n42173), .Z(n13514) );
  NANDN U13889 ( .A(n13512), .B(n42172), .Z(n13513) );
  NAND U13890 ( .A(n13514), .B(n13513), .Z(n13562) );
  NAND U13891 ( .A(b[7]), .B(a[320]), .Z(n13563) );
  XNOR U13892 ( .A(n13562), .B(n13563), .Z(n13565) );
  XOR U13893 ( .A(n13564), .B(n13565), .Z(n13571) );
  NANDN U13894 ( .A(n13515), .B(n42093), .Z(n13517) );
  XOR U13895 ( .A(n42134), .B(a[326]), .Z(n13556) );
  NANDN U13896 ( .A(n13556), .B(n42095), .Z(n13516) );
  NAND U13897 ( .A(n13517), .B(n13516), .Z(n13569) );
  NANDN U13898 ( .A(n13518), .B(n42231), .Z(n13520) );
  XOR U13899 ( .A(n188), .B(a[322]), .Z(n13559) );
  NANDN U13900 ( .A(n13559), .B(n42234), .Z(n13519) );
  AND U13901 ( .A(n13520), .B(n13519), .Z(n13568) );
  XNOR U13902 ( .A(n13569), .B(n13568), .Z(n13570) );
  XNOR U13903 ( .A(n13571), .B(n13570), .Z(n13575) );
  NANDN U13904 ( .A(n13522), .B(n13521), .Z(n13526) );
  NAND U13905 ( .A(n13524), .B(n13523), .Z(n13525) );
  AND U13906 ( .A(n13526), .B(n13525), .Z(n13574) );
  XOR U13907 ( .A(n13575), .B(n13574), .Z(n13576) );
  NANDN U13908 ( .A(n13528), .B(n13527), .Z(n13532) );
  NANDN U13909 ( .A(n13530), .B(n13529), .Z(n13531) );
  NAND U13910 ( .A(n13532), .B(n13531), .Z(n13577) );
  XOR U13911 ( .A(n13576), .B(n13577), .Z(n13544) );
  OR U13912 ( .A(n13534), .B(n13533), .Z(n13538) );
  NANDN U13913 ( .A(n13536), .B(n13535), .Z(n13537) );
  NAND U13914 ( .A(n13538), .B(n13537), .Z(n13545) );
  XNOR U13915 ( .A(n13544), .B(n13545), .Z(n13546) );
  XNOR U13916 ( .A(n13547), .B(n13546), .Z(n13580) );
  XNOR U13917 ( .A(n13580), .B(sreg[1344]), .Z(n13582) );
  NAND U13918 ( .A(n13539), .B(sreg[1343]), .Z(n13543) );
  OR U13919 ( .A(n13541), .B(n13540), .Z(n13542) );
  AND U13920 ( .A(n13543), .B(n13542), .Z(n13581) );
  XOR U13921 ( .A(n13582), .B(n13581), .Z(c[1344]) );
  NANDN U13922 ( .A(n13545), .B(n13544), .Z(n13549) );
  NAND U13923 ( .A(n13547), .B(n13546), .Z(n13548) );
  NAND U13924 ( .A(n13549), .B(n13548), .Z(n13588) );
  NAND U13925 ( .A(b[0]), .B(a[329]), .Z(n13550) );
  XNOR U13926 ( .A(b[1]), .B(n13550), .Z(n13552) );
  NAND U13927 ( .A(n62), .B(a[328]), .Z(n13551) );
  AND U13928 ( .A(n13552), .B(n13551), .Z(n13605) );
  XOR U13929 ( .A(a[325]), .B(n42197), .Z(n13594) );
  NANDN U13930 ( .A(n13594), .B(n42173), .Z(n13555) );
  NANDN U13931 ( .A(n13553), .B(n42172), .Z(n13554) );
  NAND U13932 ( .A(n13555), .B(n13554), .Z(n13603) );
  NAND U13933 ( .A(b[7]), .B(a[321]), .Z(n13604) );
  XNOR U13934 ( .A(n13603), .B(n13604), .Z(n13606) );
  XOR U13935 ( .A(n13605), .B(n13606), .Z(n13612) );
  NANDN U13936 ( .A(n13556), .B(n42093), .Z(n13558) );
  XOR U13937 ( .A(n42134), .B(a[327]), .Z(n13597) );
  NANDN U13938 ( .A(n13597), .B(n42095), .Z(n13557) );
  NAND U13939 ( .A(n13558), .B(n13557), .Z(n13610) );
  NANDN U13940 ( .A(n13559), .B(n42231), .Z(n13561) );
  XOR U13941 ( .A(n189), .B(a[323]), .Z(n13600) );
  NANDN U13942 ( .A(n13600), .B(n42234), .Z(n13560) );
  AND U13943 ( .A(n13561), .B(n13560), .Z(n13609) );
  XNOR U13944 ( .A(n13610), .B(n13609), .Z(n13611) );
  XNOR U13945 ( .A(n13612), .B(n13611), .Z(n13616) );
  NANDN U13946 ( .A(n13563), .B(n13562), .Z(n13567) );
  NAND U13947 ( .A(n13565), .B(n13564), .Z(n13566) );
  AND U13948 ( .A(n13567), .B(n13566), .Z(n13615) );
  XOR U13949 ( .A(n13616), .B(n13615), .Z(n13617) );
  NANDN U13950 ( .A(n13569), .B(n13568), .Z(n13573) );
  NANDN U13951 ( .A(n13571), .B(n13570), .Z(n13572) );
  NAND U13952 ( .A(n13573), .B(n13572), .Z(n13618) );
  XOR U13953 ( .A(n13617), .B(n13618), .Z(n13585) );
  OR U13954 ( .A(n13575), .B(n13574), .Z(n13579) );
  NANDN U13955 ( .A(n13577), .B(n13576), .Z(n13578) );
  NAND U13956 ( .A(n13579), .B(n13578), .Z(n13586) );
  XNOR U13957 ( .A(n13585), .B(n13586), .Z(n13587) );
  XNOR U13958 ( .A(n13588), .B(n13587), .Z(n13621) );
  XNOR U13959 ( .A(n13621), .B(sreg[1345]), .Z(n13623) );
  NAND U13960 ( .A(n13580), .B(sreg[1344]), .Z(n13584) );
  OR U13961 ( .A(n13582), .B(n13581), .Z(n13583) );
  AND U13962 ( .A(n13584), .B(n13583), .Z(n13622) );
  XOR U13963 ( .A(n13623), .B(n13622), .Z(c[1345]) );
  NANDN U13964 ( .A(n13586), .B(n13585), .Z(n13590) );
  NAND U13965 ( .A(n13588), .B(n13587), .Z(n13589) );
  NAND U13966 ( .A(n13590), .B(n13589), .Z(n13629) );
  NAND U13967 ( .A(b[0]), .B(a[330]), .Z(n13591) );
  XNOR U13968 ( .A(b[1]), .B(n13591), .Z(n13593) );
  NAND U13969 ( .A(n62), .B(a[329]), .Z(n13592) );
  AND U13970 ( .A(n13593), .B(n13592), .Z(n13646) );
  XOR U13971 ( .A(a[326]), .B(n42197), .Z(n13635) );
  NANDN U13972 ( .A(n13635), .B(n42173), .Z(n13596) );
  NANDN U13973 ( .A(n13594), .B(n42172), .Z(n13595) );
  NAND U13974 ( .A(n13596), .B(n13595), .Z(n13644) );
  NAND U13975 ( .A(b[7]), .B(a[322]), .Z(n13645) );
  XNOR U13976 ( .A(n13644), .B(n13645), .Z(n13647) );
  XOR U13977 ( .A(n13646), .B(n13647), .Z(n13653) );
  NANDN U13978 ( .A(n13597), .B(n42093), .Z(n13599) );
  XOR U13979 ( .A(n42134), .B(a[328]), .Z(n13638) );
  NANDN U13980 ( .A(n13638), .B(n42095), .Z(n13598) );
  NAND U13981 ( .A(n13599), .B(n13598), .Z(n13651) );
  NANDN U13982 ( .A(n13600), .B(n42231), .Z(n13602) );
  XOR U13983 ( .A(n189), .B(a[324]), .Z(n13641) );
  NANDN U13984 ( .A(n13641), .B(n42234), .Z(n13601) );
  AND U13985 ( .A(n13602), .B(n13601), .Z(n13650) );
  XNOR U13986 ( .A(n13651), .B(n13650), .Z(n13652) );
  XNOR U13987 ( .A(n13653), .B(n13652), .Z(n13657) );
  NANDN U13988 ( .A(n13604), .B(n13603), .Z(n13608) );
  NAND U13989 ( .A(n13606), .B(n13605), .Z(n13607) );
  AND U13990 ( .A(n13608), .B(n13607), .Z(n13656) );
  XOR U13991 ( .A(n13657), .B(n13656), .Z(n13658) );
  NANDN U13992 ( .A(n13610), .B(n13609), .Z(n13614) );
  NANDN U13993 ( .A(n13612), .B(n13611), .Z(n13613) );
  NAND U13994 ( .A(n13614), .B(n13613), .Z(n13659) );
  XOR U13995 ( .A(n13658), .B(n13659), .Z(n13626) );
  OR U13996 ( .A(n13616), .B(n13615), .Z(n13620) );
  NANDN U13997 ( .A(n13618), .B(n13617), .Z(n13619) );
  NAND U13998 ( .A(n13620), .B(n13619), .Z(n13627) );
  XNOR U13999 ( .A(n13626), .B(n13627), .Z(n13628) );
  XNOR U14000 ( .A(n13629), .B(n13628), .Z(n13662) );
  XNOR U14001 ( .A(n13662), .B(sreg[1346]), .Z(n13664) );
  NAND U14002 ( .A(n13621), .B(sreg[1345]), .Z(n13625) );
  OR U14003 ( .A(n13623), .B(n13622), .Z(n13624) );
  AND U14004 ( .A(n13625), .B(n13624), .Z(n13663) );
  XOR U14005 ( .A(n13664), .B(n13663), .Z(c[1346]) );
  NANDN U14006 ( .A(n13627), .B(n13626), .Z(n13631) );
  NAND U14007 ( .A(n13629), .B(n13628), .Z(n13630) );
  NAND U14008 ( .A(n13631), .B(n13630), .Z(n13670) );
  NAND U14009 ( .A(b[0]), .B(a[331]), .Z(n13632) );
  XNOR U14010 ( .A(b[1]), .B(n13632), .Z(n13634) );
  NAND U14011 ( .A(n62), .B(a[330]), .Z(n13633) );
  AND U14012 ( .A(n13634), .B(n13633), .Z(n13687) );
  XOR U14013 ( .A(a[327]), .B(n42197), .Z(n13676) );
  NANDN U14014 ( .A(n13676), .B(n42173), .Z(n13637) );
  NANDN U14015 ( .A(n13635), .B(n42172), .Z(n13636) );
  NAND U14016 ( .A(n13637), .B(n13636), .Z(n13685) );
  NAND U14017 ( .A(b[7]), .B(a[323]), .Z(n13686) );
  XNOR U14018 ( .A(n13685), .B(n13686), .Z(n13688) );
  XOR U14019 ( .A(n13687), .B(n13688), .Z(n13694) );
  NANDN U14020 ( .A(n13638), .B(n42093), .Z(n13640) );
  XOR U14021 ( .A(n42134), .B(a[329]), .Z(n13679) );
  NANDN U14022 ( .A(n13679), .B(n42095), .Z(n13639) );
  NAND U14023 ( .A(n13640), .B(n13639), .Z(n13692) );
  NANDN U14024 ( .A(n13641), .B(n42231), .Z(n13643) );
  XOR U14025 ( .A(n189), .B(a[325]), .Z(n13682) );
  NANDN U14026 ( .A(n13682), .B(n42234), .Z(n13642) );
  AND U14027 ( .A(n13643), .B(n13642), .Z(n13691) );
  XNOR U14028 ( .A(n13692), .B(n13691), .Z(n13693) );
  XNOR U14029 ( .A(n13694), .B(n13693), .Z(n13698) );
  NANDN U14030 ( .A(n13645), .B(n13644), .Z(n13649) );
  NAND U14031 ( .A(n13647), .B(n13646), .Z(n13648) );
  AND U14032 ( .A(n13649), .B(n13648), .Z(n13697) );
  XOR U14033 ( .A(n13698), .B(n13697), .Z(n13699) );
  NANDN U14034 ( .A(n13651), .B(n13650), .Z(n13655) );
  NANDN U14035 ( .A(n13653), .B(n13652), .Z(n13654) );
  NAND U14036 ( .A(n13655), .B(n13654), .Z(n13700) );
  XOR U14037 ( .A(n13699), .B(n13700), .Z(n13667) );
  OR U14038 ( .A(n13657), .B(n13656), .Z(n13661) );
  NANDN U14039 ( .A(n13659), .B(n13658), .Z(n13660) );
  NAND U14040 ( .A(n13661), .B(n13660), .Z(n13668) );
  XNOR U14041 ( .A(n13667), .B(n13668), .Z(n13669) );
  XNOR U14042 ( .A(n13670), .B(n13669), .Z(n13703) );
  XNOR U14043 ( .A(n13703), .B(sreg[1347]), .Z(n13705) );
  NAND U14044 ( .A(n13662), .B(sreg[1346]), .Z(n13666) );
  OR U14045 ( .A(n13664), .B(n13663), .Z(n13665) );
  AND U14046 ( .A(n13666), .B(n13665), .Z(n13704) );
  XOR U14047 ( .A(n13705), .B(n13704), .Z(c[1347]) );
  NANDN U14048 ( .A(n13668), .B(n13667), .Z(n13672) );
  NAND U14049 ( .A(n13670), .B(n13669), .Z(n13671) );
  NAND U14050 ( .A(n13672), .B(n13671), .Z(n13711) );
  NAND U14051 ( .A(b[0]), .B(a[332]), .Z(n13673) );
  XNOR U14052 ( .A(b[1]), .B(n13673), .Z(n13675) );
  NAND U14053 ( .A(n62), .B(a[331]), .Z(n13674) );
  AND U14054 ( .A(n13675), .B(n13674), .Z(n13728) );
  XOR U14055 ( .A(a[328]), .B(n42197), .Z(n13717) );
  NANDN U14056 ( .A(n13717), .B(n42173), .Z(n13678) );
  NANDN U14057 ( .A(n13676), .B(n42172), .Z(n13677) );
  NAND U14058 ( .A(n13678), .B(n13677), .Z(n13726) );
  NAND U14059 ( .A(b[7]), .B(a[324]), .Z(n13727) );
  XNOR U14060 ( .A(n13726), .B(n13727), .Z(n13729) );
  XOR U14061 ( .A(n13728), .B(n13729), .Z(n13735) );
  NANDN U14062 ( .A(n13679), .B(n42093), .Z(n13681) );
  XOR U14063 ( .A(n42134), .B(a[330]), .Z(n13720) );
  NANDN U14064 ( .A(n13720), .B(n42095), .Z(n13680) );
  NAND U14065 ( .A(n13681), .B(n13680), .Z(n13733) );
  NANDN U14066 ( .A(n13682), .B(n42231), .Z(n13684) );
  XOR U14067 ( .A(n189), .B(a[326]), .Z(n13723) );
  NANDN U14068 ( .A(n13723), .B(n42234), .Z(n13683) );
  AND U14069 ( .A(n13684), .B(n13683), .Z(n13732) );
  XNOR U14070 ( .A(n13733), .B(n13732), .Z(n13734) );
  XNOR U14071 ( .A(n13735), .B(n13734), .Z(n13739) );
  NANDN U14072 ( .A(n13686), .B(n13685), .Z(n13690) );
  NAND U14073 ( .A(n13688), .B(n13687), .Z(n13689) );
  AND U14074 ( .A(n13690), .B(n13689), .Z(n13738) );
  XOR U14075 ( .A(n13739), .B(n13738), .Z(n13740) );
  NANDN U14076 ( .A(n13692), .B(n13691), .Z(n13696) );
  NANDN U14077 ( .A(n13694), .B(n13693), .Z(n13695) );
  NAND U14078 ( .A(n13696), .B(n13695), .Z(n13741) );
  XOR U14079 ( .A(n13740), .B(n13741), .Z(n13708) );
  OR U14080 ( .A(n13698), .B(n13697), .Z(n13702) );
  NANDN U14081 ( .A(n13700), .B(n13699), .Z(n13701) );
  NAND U14082 ( .A(n13702), .B(n13701), .Z(n13709) );
  XNOR U14083 ( .A(n13708), .B(n13709), .Z(n13710) );
  XNOR U14084 ( .A(n13711), .B(n13710), .Z(n13744) );
  XNOR U14085 ( .A(n13744), .B(sreg[1348]), .Z(n13746) );
  NAND U14086 ( .A(n13703), .B(sreg[1347]), .Z(n13707) );
  OR U14087 ( .A(n13705), .B(n13704), .Z(n13706) );
  AND U14088 ( .A(n13707), .B(n13706), .Z(n13745) );
  XOR U14089 ( .A(n13746), .B(n13745), .Z(c[1348]) );
  NANDN U14090 ( .A(n13709), .B(n13708), .Z(n13713) );
  NAND U14091 ( .A(n13711), .B(n13710), .Z(n13712) );
  NAND U14092 ( .A(n13713), .B(n13712), .Z(n13752) );
  NAND U14093 ( .A(b[0]), .B(a[333]), .Z(n13714) );
  XNOR U14094 ( .A(b[1]), .B(n13714), .Z(n13716) );
  NAND U14095 ( .A(n62), .B(a[332]), .Z(n13715) );
  AND U14096 ( .A(n13716), .B(n13715), .Z(n13769) );
  XOR U14097 ( .A(a[329]), .B(n42197), .Z(n13758) );
  NANDN U14098 ( .A(n13758), .B(n42173), .Z(n13719) );
  NANDN U14099 ( .A(n13717), .B(n42172), .Z(n13718) );
  NAND U14100 ( .A(n13719), .B(n13718), .Z(n13767) );
  NAND U14101 ( .A(b[7]), .B(a[325]), .Z(n13768) );
  XNOR U14102 ( .A(n13767), .B(n13768), .Z(n13770) );
  XOR U14103 ( .A(n13769), .B(n13770), .Z(n13776) );
  NANDN U14104 ( .A(n13720), .B(n42093), .Z(n13722) );
  XOR U14105 ( .A(n42134), .B(a[331]), .Z(n13761) );
  NANDN U14106 ( .A(n13761), .B(n42095), .Z(n13721) );
  NAND U14107 ( .A(n13722), .B(n13721), .Z(n13774) );
  NANDN U14108 ( .A(n13723), .B(n42231), .Z(n13725) );
  XOR U14109 ( .A(n189), .B(a[327]), .Z(n13764) );
  NANDN U14110 ( .A(n13764), .B(n42234), .Z(n13724) );
  AND U14111 ( .A(n13725), .B(n13724), .Z(n13773) );
  XNOR U14112 ( .A(n13774), .B(n13773), .Z(n13775) );
  XNOR U14113 ( .A(n13776), .B(n13775), .Z(n13780) );
  NANDN U14114 ( .A(n13727), .B(n13726), .Z(n13731) );
  NAND U14115 ( .A(n13729), .B(n13728), .Z(n13730) );
  AND U14116 ( .A(n13731), .B(n13730), .Z(n13779) );
  XOR U14117 ( .A(n13780), .B(n13779), .Z(n13781) );
  NANDN U14118 ( .A(n13733), .B(n13732), .Z(n13737) );
  NANDN U14119 ( .A(n13735), .B(n13734), .Z(n13736) );
  NAND U14120 ( .A(n13737), .B(n13736), .Z(n13782) );
  XOR U14121 ( .A(n13781), .B(n13782), .Z(n13749) );
  OR U14122 ( .A(n13739), .B(n13738), .Z(n13743) );
  NANDN U14123 ( .A(n13741), .B(n13740), .Z(n13742) );
  NAND U14124 ( .A(n13743), .B(n13742), .Z(n13750) );
  XNOR U14125 ( .A(n13749), .B(n13750), .Z(n13751) );
  XNOR U14126 ( .A(n13752), .B(n13751), .Z(n13785) );
  XNOR U14127 ( .A(n13785), .B(sreg[1349]), .Z(n13787) );
  NAND U14128 ( .A(n13744), .B(sreg[1348]), .Z(n13748) );
  OR U14129 ( .A(n13746), .B(n13745), .Z(n13747) );
  AND U14130 ( .A(n13748), .B(n13747), .Z(n13786) );
  XOR U14131 ( .A(n13787), .B(n13786), .Z(c[1349]) );
  NANDN U14132 ( .A(n13750), .B(n13749), .Z(n13754) );
  NAND U14133 ( .A(n13752), .B(n13751), .Z(n13753) );
  NAND U14134 ( .A(n13754), .B(n13753), .Z(n13793) );
  NAND U14135 ( .A(b[0]), .B(a[334]), .Z(n13755) );
  XNOR U14136 ( .A(b[1]), .B(n13755), .Z(n13757) );
  NAND U14137 ( .A(n62), .B(a[333]), .Z(n13756) );
  AND U14138 ( .A(n13757), .B(n13756), .Z(n13810) );
  XOR U14139 ( .A(a[330]), .B(n42197), .Z(n13799) );
  NANDN U14140 ( .A(n13799), .B(n42173), .Z(n13760) );
  NANDN U14141 ( .A(n13758), .B(n42172), .Z(n13759) );
  NAND U14142 ( .A(n13760), .B(n13759), .Z(n13808) );
  NAND U14143 ( .A(b[7]), .B(a[326]), .Z(n13809) );
  XNOR U14144 ( .A(n13808), .B(n13809), .Z(n13811) );
  XOR U14145 ( .A(n13810), .B(n13811), .Z(n13817) );
  NANDN U14146 ( .A(n13761), .B(n42093), .Z(n13763) );
  XOR U14147 ( .A(n42134), .B(a[332]), .Z(n13802) );
  NANDN U14148 ( .A(n13802), .B(n42095), .Z(n13762) );
  NAND U14149 ( .A(n13763), .B(n13762), .Z(n13815) );
  NANDN U14150 ( .A(n13764), .B(n42231), .Z(n13766) );
  XOR U14151 ( .A(n189), .B(a[328]), .Z(n13805) );
  NANDN U14152 ( .A(n13805), .B(n42234), .Z(n13765) );
  AND U14153 ( .A(n13766), .B(n13765), .Z(n13814) );
  XNOR U14154 ( .A(n13815), .B(n13814), .Z(n13816) );
  XNOR U14155 ( .A(n13817), .B(n13816), .Z(n13821) );
  NANDN U14156 ( .A(n13768), .B(n13767), .Z(n13772) );
  NAND U14157 ( .A(n13770), .B(n13769), .Z(n13771) );
  AND U14158 ( .A(n13772), .B(n13771), .Z(n13820) );
  XOR U14159 ( .A(n13821), .B(n13820), .Z(n13822) );
  NANDN U14160 ( .A(n13774), .B(n13773), .Z(n13778) );
  NANDN U14161 ( .A(n13776), .B(n13775), .Z(n13777) );
  NAND U14162 ( .A(n13778), .B(n13777), .Z(n13823) );
  XOR U14163 ( .A(n13822), .B(n13823), .Z(n13790) );
  OR U14164 ( .A(n13780), .B(n13779), .Z(n13784) );
  NANDN U14165 ( .A(n13782), .B(n13781), .Z(n13783) );
  NAND U14166 ( .A(n13784), .B(n13783), .Z(n13791) );
  XNOR U14167 ( .A(n13790), .B(n13791), .Z(n13792) );
  XNOR U14168 ( .A(n13793), .B(n13792), .Z(n13826) );
  XNOR U14169 ( .A(n13826), .B(sreg[1350]), .Z(n13828) );
  NAND U14170 ( .A(n13785), .B(sreg[1349]), .Z(n13789) );
  OR U14171 ( .A(n13787), .B(n13786), .Z(n13788) );
  AND U14172 ( .A(n13789), .B(n13788), .Z(n13827) );
  XOR U14173 ( .A(n13828), .B(n13827), .Z(c[1350]) );
  NANDN U14174 ( .A(n13791), .B(n13790), .Z(n13795) );
  NAND U14175 ( .A(n13793), .B(n13792), .Z(n13794) );
  NAND U14176 ( .A(n13795), .B(n13794), .Z(n13834) );
  NAND U14177 ( .A(b[0]), .B(a[335]), .Z(n13796) );
  XNOR U14178 ( .A(b[1]), .B(n13796), .Z(n13798) );
  NAND U14179 ( .A(n62), .B(a[334]), .Z(n13797) );
  AND U14180 ( .A(n13798), .B(n13797), .Z(n13851) );
  XOR U14181 ( .A(a[331]), .B(n42197), .Z(n13840) );
  NANDN U14182 ( .A(n13840), .B(n42173), .Z(n13801) );
  NANDN U14183 ( .A(n13799), .B(n42172), .Z(n13800) );
  NAND U14184 ( .A(n13801), .B(n13800), .Z(n13849) );
  NAND U14185 ( .A(b[7]), .B(a[327]), .Z(n13850) );
  XNOR U14186 ( .A(n13849), .B(n13850), .Z(n13852) );
  XOR U14187 ( .A(n13851), .B(n13852), .Z(n13858) );
  NANDN U14188 ( .A(n13802), .B(n42093), .Z(n13804) );
  XOR U14189 ( .A(n42134), .B(a[333]), .Z(n13843) );
  NANDN U14190 ( .A(n13843), .B(n42095), .Z(n13803) );
  NAND U14191 ( .A(n13804), .B(n13803), .Z(n13856) );
  NANDN U14192 ( .A(n13805), .B(n42231), .Z(n13807) );
  XOR U14193 ( .A(n189), .B(a[329]), .Z(n13846) );
  NANDN U14194 ( .A(n13846), .B(n42234), .Z(n13806) );
  AND U14195 ( .A(n13807), .B(n13806), .Z(n13855) );
  XNOR U14196 ( .A(n13856), .B(n13855), .Z(n13857) );
  XNOR U14197 ( .A(n13858), .B(n13857), .Z(n13862) );
  NANDN U14198 ( .A(n13809), .B(n13808), .Z(n13813) );
  NAND U14199 ( .A(n13811), .B(n13810), .Z(n13812) );
  AND U14200 ( .A(n13813), .B(n13812), .Z(n13861) );
  XOR U14201 ( .A(n13862), .B(n13861), .Z(n13863) );
  NANDN U14202 ( .A(n13815), .B(n13814), .Z(n13819) );
  NANDN U14203 ( .A(n13817), .B(n13816), .Z(n13818) );
  NAND U14204 ( .A(n13819), .B(n13818), .Z(n13864) );
  XOR U14205 ( .A(n13863), .B(n13864), .Z(n13831) );
  OR U14206 ( .A(n13821), .B(n13820), .Z(n13825) );
  NANDN U14207 ( .A(n13823), .B(n13822), .Z(n13824) );
  NAND U14208 ( .A(n13825), .B(n13824), .Z(n13832) );
  XNOR U14209 ( .A(n13831), .B(n13832), .Z(n13833) );
  XNOR U14210 ( .A(n13834), .B(n13833), .Z(n13867) );
  XNOR U14211 ( .A(n13867), .B(sreg[1351]), .Z(n13869) );
  NAND U14212 ( .A(n13826), .B(sreg[1350]), .Z(n13830) );
  OR U14213 ( .A(n13828), .B(n13827), .Z(n13829) );
  AND U14214 ( .A(n13830), .B(n13829), .Z(n13868) );
  XOR U14215 ( .A(n13869), .B(n13868), .Z(c[1351]) );
  NANDN U14216 ( .A(n13832), .B(n13831), .Z(n13836) );
  NAND U14217 ( .A(n13834), .B(n13833), .Z(n13835) );
  NAND U14218 ( .A(n13836), .B(n13835), .Z(n13875) );
  NAND U14219 ( .A(b[0]), .B(a[336]), .Z(n13837) );
  XNOR U14220 ( .A(b[1]), .B(n13837), .Z(n13839) );
  NAND U14221 ( .A(n63), .B(a[335]), .Z(n13838) );
  AND U14222 ( .A(n13839), .B(n13838), .Z(n13892) );
  XOR U14223 ( .A(a[332]), .B(n42197), .Z(n13881) );
  NANDN U14224 ( .A(n13881), .B(n42173), .Z(n13842) );
  NANDN U14225 ( .A(n13840), .B(n42172), .Z(n13841) );
  NAND U14226 ( .A(n13842), .B(n13841), .Z(n13890) );
  NAND U14227 ( .A(b[7]), .B(a[328]), .Z(n13891) );
  XNOR U14228 ( .A(n13890), .B(n13891), .Z(n13893) );
  XOR U14229 ( .A(n13892), .B(n13893), .Z(n13899) );
  NANDN U14230 ( .A(n13843), .B(n42093), .Z(n13845) );
  XOR U14231 ( .A(n42134), .B(a[334]), .Z(n13884) );
  NANDN U14232 ( .A(n13884), .B(n42095), .Z(n13844) );
  NAND U14233 ( .A(n13845), .B(n13844), .Z(n13897) );
  NANDN U14234 ( .A(n13846), .B(n42231), .Z(n13848) );
  XOR U14235 ( .A(n189), .B(a[330]), .Z(n13887) );
  NANDN U14236 ( .A(n13887), .B(n42234), .Z(n13847) );
  AND U14237 ( .A(n13848), .B(n13847), .Z(n13896) );
  XNOR U14238 ( .A(n13897), .B(n13896), .Z(n13898) );
  XNOR U14239 ( .A(n13899), .B(n13898), .Z(n13903) );
  NANDN U14240 ( .A(n13850), .B(n13849), .Z(n13854) );
  NAND U14241 ( .A(n13852), .B(n13851), .Z(n13853) );
  AND U14242 ( .A(n13854), .B(n13853), .Z(n13902) );
  XOR U14243 ( .A(n13903), .B(n13902), .Z(n13904) );
  NANDN U14244 ( .A(n13856), .B(n13855), .Z(n13860) );
  NANDN U14245 ( .A(n13858), .B(n13857), .Z(n13859) );
  NAND U14246 ( .A(n13860), .B(n13859), .Z(n13905) );
  XOR U14247 ( .A(n13904), .B(n13905), .Z(n13872) );
  OR U14248 ( .A(n13862), .B(n13861), .Z(n13866) );
  NANDN U14249 ( .A(n13864), .B(n13863), .Z(n13865) );
  NAND U14250 ( .A(n13866), .B(n13865), .Z(n13873) );
  XNOR U14251 ( .A(n13872), .B(n13873), .Z(n13874) );
  XNOR U14252 ( .A(n13875), .B(n13874), .Z(n13908) );
  XNOR U14253 ( .A(n13908), .B(sreg[1352]), .Z(n13910) );
  NAND U14254 ( .A(n13867), .B(sreg[1351]), .Z(n13871) );
  OR U14255 ( .A(n13869), .B(n13868), .Z(n13870) );
  AND U14256 ( .A(n13871), .B(n13870), .Z(n13909) );
  XOR U14257 ( .A(n13910), .B(n13909), .Z(c[1352]) );
  NANDN U14258 ( .A(n13873), .B(n13872), .Z(n13877) );
  NAND U14259 ( .A(n13875), .B(n13874), .Z(n13876) );
  NAND U14260 ( .A(n13877), .B(n13876), .Z(n13916) );
  NAND U14261 ( .A(b[0]), .B(a[337]), .Z(n13878) );
  XNOR U14262 ( .A(b[1]), .B(n13878), .Z(n13880) );
  NAND U14263 ( .A(n63), .B(a[336]), .Z(n13879) );
  AND U14264 ( .A(n13880), .B(n13879), .Z(n13933) );
  XOR U14265 ( .A(a[333]), .B(n42197), .Z(n13922) );
  NANDN U14266 ( .A(n13922), .B(n42173), .Z(n13883) );
  NANDN U14267 ( .A(n13881), .B(n42172), .Z(n13882) );
  NAND U14268 ( .A(n13883), .B(n13882), .Z(n13931) );
  NAND U14269 ( .A(b[7]), .B(a[329]), .Z(n13932) );
  XNOR U14270 ( .A(n13931), .B(n13932), .Z(n13934) );
  XOR U14271 ( .A(n13933), .B(n13934), .Z(n13940) );
  NANDN U14272 ( .A(n13884), .B(n42093), .Z(n13886) );
  XOR U14273 ( .A(n42134), .B(a[335]), .Z(n13925) );
  NANDN U14274 ( .A(n13925), .B(n42095), .Z(n13885) );
  NAND U14275 ( .A(n13886), .B(n13885), .Z(n13938) );
  NANDN U14276 ( .A(n13887), .B(n42231), .Z(n13889) );
  XOR U14277 ( .A(n189), .B(a[331]), .Z(n13928) );
  NANDN U14278 ( .A(n13928), .B(n42234), .Z(n13888) );
  AND U14279 ( .A(n13889), .B(n13888), .Z(n13937) );
  XNOR U14280 ( .A(n13938), .B(n13937), .Z(n13939) );
  XNOR U14281 ( .A(n13940), .B(n13939), .Z(n13944) );
  NANDN U14282 ( .A(n13891), .B(n13890), .Z(n13895) );
  NAND U14283 ( .A(n13893), .B(n13892), .Z(n13894) );
  AND U14284 ( .A(n13895), .B(n13894), .Z(n13943) );
  XOR U14285 ( .A(n13944), .B(n13943), .Z(n13945) );
  NANDN U14286 ( .A(n13897), .B(n13896), .Z(n13901) );
  NANDN U14287 ( .A(n13899), .B(n13898), .Z(n13900) );
  NAND U14288 ( .A(n13901), .B(n13900), .Z(n13946) );
  XOR U14289 ( .A(n13945), .B(n13946), .Z(n13913) );
  OR U14290 ( .A(n13903), .B(n13902), .Z(n13907) );
  NANDN U14291 ( .A(n13905), .B(n13904), .Z(n13906) );
  NAND U14292 ( .A(n13907), .B(n13906), .Z(n13914) );
  XNOR U14293 ( .A(n13913), .B(n13914), .Z(n13915) );
  XNOR U14294 ( .A(n13916), .B(n13915), .Z(n13949) );
  XNOR U14295 ( .A(n13949), .B(sreg[1353]), .Z(n13951) );
  NAND U14296 ( .A(n13908), .B(sreg[1352]), .Z(n13912) );
  OR U14297 ( .A(n13910), .B(n13909), .Z(n13911) );
  AND U14298 ( .A(n13912), .B(n13911), .Z(n13950) );
  XOR U14299 ( .A(n13951), .B(n13950), .Z(c[1353]) );
  NANDN U14300 ( .A(n13914), .B(n13913), .Z(n13918) );
  NAND U14301 ( .A(n13916), .B(n13915), .Z(n13917) );
  NAND U14302 ( .A(n13918), .B(n13917), .Z(n13957) );
  NAND U14303 ( .A(b[0]), .B(a[338]), .Z(n13919) );
  XNOR U14304 ( .A(b[1]), .B(n13919), .Z(n13921) );
  NAND U14305 ( .A(n63), .B(a[337]), .Z(n13920) );
  AND U14306 ( .A(n13921), .B(n13920), .Z(n13974) );
  XOR U14307 ( .A(a[334]), .B(n42197), .Z(n13963) );
  NANDN U14308 ( .A(n13963), .B(n42173), .Z(n13924) );
  NANDN U14309 ( .A(n13922), .B(n42172), .Z(n13923) );
  NAND U14310 ( .A(n13924), .B(n13923), .Z(n13972) );
  NAND U14311 ( .A(b[7]), .B(a[330]), .Z(n13973) );
  XNOR U14312 ( .A(n13972), .B(n13973), .Z(n13975) );
  XOR U14313 ( .A(n13974), .B(n13975), .Z(n13981) );
  NANDN U14314 ( .A(n13925), .B(n42093), .Z(n13927) );
  XOR U14315 ( .A(n42134), .B(a[336]), .Z(n13966) );
  NANDN U14316 ( .A(n13966), .B(n42095), .Z(n13926) );
  NAND U14317 ( .A(n13927), .B(n13926), .Z(n13979) );
  NANDN U14318 ( .A(n13928), .B(n42231), .Z(n13930) );
  XOR U14319 ( .A(n189), .B(a[332]), .Z(n13969) );
  NANDN U14320 ( .A(n13969), .B(n42234), .Z(n13929) );
  AND U14321 ( .A(n13930), .B(n13929), .Z(n13978) );
  XNOR U14322 ( .A(n13979), .B(n13978), .Z(n13980) );
  XNOR U14323 ( .A(n13981), .B(n13980), .Z(n13985) );
  NANDN U14324 ( .A(n13932), .B(n13931), .Z(n13936) );
  NAND U14325 ( .A(n13934), .B(n13933), .Z(n13935) );
  AND U14326 ( .A(n13936), .B(n13935), .Z(n13984) );
  XOR U14327 ( .A(n13985), .B(n13984), .Z(n13986) );
  NANDN U14328 ( .A(n13938), .B(n13937), .Z(n13942) );
  NANDN U14329 ( .A(n13940), .B(n13939), .Z(n13941) );
  NAND U14330 ( .A(n13942), .B(n13941), .Z(n13987) );
  XOR U14331 ( .A(n13986), .B(n13987), .Z(n13954) );
  OR U14332 ( .A(n13944), .B(n13943), .Z(n13948) );
  NANDN U14333 ( .A(n13946), .B(n13945), .Z(n13947) );
  NAND U14334 ( .A(n13948), .B(n13947), .Z(n13955) );
  XNOR U14335 ( .A(n13954), .B(n13955), .Z(n13956) );
  XNOR U14336 ( .A(n13957), .B(n13956), .Z(n13990) );
  XNOR U14337 ( .A(n13990), .B(sreg[1354]), .Z(n13992) );
  NAND U14338 ( .A(n13949), .B(sreg[1353]), .Z(n13953) );
  OR U14339 ( .A(n13951), .B(n13950), .Z(n13952) );
  AND U14340 ( .A(n13953), .B(n13952), .Z(n13991) );
  XOR U14341 ( .A(n13992), .B(n13991), .Z(c[1354]) );
  NANDN U14342 ( .A(n13955), .B(n13954), .Z(n13959) );
  NAND U14343 ( .A(n13957), .B(n13956), .Z(n13958) );
  NAND U14344 ( .A(n13959), .B(n13958), .Z(n13998) );
  NAND U14345 ( .A(b[0]), .B(a[339]), .Z(n13960) );
  XNOR U14346 ( .A(b[1]), .B(n13960), .Z(n13962) );
  NAND U14347 ( .A(n63), .B(a[338]), .Z(n13961) );
  AND U14348 ( .A(n13962), .B(n13961), .Z(n14015) );
  XOR U14349 ( .A(a[335]), .B(n42197), .Z(n14004) );
  NANDN U14350 ( .A(n14004), .B(n42173), .Z(n13965) );
  NANDN U14351 ( .A(n13963), .B(n42172), .Z(n13964) );
  NAND U14352 ( .A(n13965), .B(n13964), .Z(n14013) );
  NAND U14353 ( .A(b[7]), .B(a[331]), .Z(n14014) );
  XNOR U14354 ( .A(n14013), .B(n14014), .Z(n14016) );
  XOR U14355 ( .A(n14015), .B(n14016), .Z(n14022) );
  NANDN U14356 ( .A(n13966), .B(n42093), .Z(n13968) );
  XOR U14357 ( .A(n42134), .B(a[337]), .Z(n14007) );
  NANDN U14358 ( .A(n14007), .B(n42095), .Z(n13967) );
  NAND U14359 ( .A(n13968), .B(n13967), .Z(n14020) );
  NANDN U14360 ( .A(n13969), .B(n42231), .Z(n13971) );
  XOR U14361 ( .A(n189), .B(a[333]), .Z(n14010) );
  NANDN U14362 ( .A(n14010), .B(n42234), .Z(n13970) );
  AND U14363 ( .A(n13971), .B(n13970), .Z(n14019) );
  XNOR U14364 ( .A(n14020), .B(n14019), .Z(n14021) );
  XNOR U14365 ( .A(n14022), .B(n14021), .Z(n14026) );
  NANDN U14366 ( .A(n13973), .B(n13972), .Z(n13977) );
  NAND U14367 ( .A(n13975), .B(n13974), .Z(n13976) );
  AND U14368 ( .A(n13977), .B(n13976), .Z(n14025) );
  XOR U14369 ( .A(n14026), .B(n14025), .Z(n14027) );
  NANDN U14370 ( .A(n13979), .B(n13978), .Z(n13983) );
  NANDN U14371 ( .A(n13981), .B(n13980), .Z(n13982) );
  NAND U14372 ( .A(n13983), .B(n13982), .Z(n14028) );
  XOR U14373 ( .A(n14027), .B(n14028), .Z(n13995) );
  OR U14374 ( .A(n13985), .B(n13984), .Z(n13989) );
  NANDN U14375 ( .A(n13987), .B(n13986), .Z(n13988) );
  NAND U14376 ( .A(n13989), .B(n13988), .Z(n13996) );
  XNOR U14377 ( .A(n13995), .B(n13996), .Z(n13997) );
  XNOR U14378 ( .A(n13998), .B(n13997), .Z(n14031) );
  XNOR U14379 ( .A(n14031), .B(sreg[1355]), .Z(n14033) );
  NAND U14380 ( .A(n13990), .B(sreg[1354]), .Z(n13994) );
  OR U14381 ( .A(n13992), .B(n13991), .Z(n13993) );
  AND U14382 ( .A(n13994), .B(n13993), .Z(n14032) );
  XOR U14383 ( .A(n14033), .B(n14032), .Z(c[1355]) );
  NANDN U14384 ( .A(n13996), .B(n13995), .Z(n14000) );
  NAND U14385 ( .A(n13998), .B(n13997), .Z(n13999) );
  NAND U14386 ( .A(n14000), .B(n13999), .Z(n14039) );
  NAND U14387 ( .A(b[0]), .B(a[340]), .Z(n14001) );
  XNOR U14388 ( .A(b[1]), .B(n14001), .Z(n14003) );
  NAND U14389 ( .A(n63), .B(a[339]), .Z(n14002) );
  AND U14390 ( .A(n14003), .B(n14002), .Z(n14056) );
  XOR U14391 ( .A(a[336]), .B(n42197), .Z(n14045) );
  NANDN U14392 ( .A(n14045), .B(n42173), .Z(n14006) );
  NANDN U14393 ( .A(n14004), .B(n42172), .Z(n14005) );
  NAND U14394 ( .A(n14006), .B(n14005), .Z(n14054) );
  NAND U14395 ( .A(b[7]), .B(a[332]), .Z(n14055) );
  XNOR U14396 ( .A(n14054), .B(n14055), .Z(n14057) );
  XOR U14397 ( .A(n14056), .B(n14057), .Z(n14063) );
  NANDN U14398 ( .A(n14007), .B(n42093), .Z(n14009) );
  XOR U14399 ( .A(n42134), .B(a[338]), .Z(n14048) );
  NANDN U14400 ( .A(n14048), .B(n42095), .Z(n14008) );
  NAND U14401 ( .A(n14009), .B(n14008), .Z(n14061) );
  NANDN U14402 ( .A(n14010), .B(n42231), .Z(n14012) );
  XOR U14403 ( .A(n189), .B(a[334]), .Z(n14051) );
  NANDN U14404 ( .A(n14051), .B(n42234), .Z(n14011) );
  AND U14405 ( .A(n14012), .B(n14011), .Z(n14060) );
  XNOR U14406 ( .A(n14061), .B(n14060), .Z(n14062) );
  XNOR U14407 ( .A(n14063), .B(n14062), .Z(n14067) );
  NANDN U14408 ( .A(n14014), .B(n14013), .Z(n14018) );
  NAND U14409 ( .A(n14016), .B(n14015), .Z(n14017) );
  AND U14410 ( .A(n14018), .B(n14017), .Z(n14066) );
  XOR U14411 ( .A(n14067), .B(n14066), .Z(n14068) );
  NANDN U14412 ( .A(n14020), .B(n14019), .Z(n14024) );
  NANDN U14413 ( .A(n14022), .B(n14021), .Z(n14023) );
  NAND U14414 ( .A(n14024), .B(n14023), .Z(n14069) );
  XOR U14415 ( .A(n14068), .B(n14069), .Z(n14036) );
  OR U14416 ( .A(n14026), .B(n14025), .Z(n14030) );
  NANDN U14417 ( .A(n14028), .B(n14027), .Z(n14029) );
  NAND U14418 ( .A(n14030), .B(n14029), .Z(n14037) );
  XNOR U14419 ( .A(n14036), .B(n14037), .Z(n14038) );
  XNOR U14420 ( .A(n14039), .B(n14038), .Z(n14072) );
  XNOR U14421 ( .A(n14072), .B(sreg[1356]), .Z(n14074) );
  NAND U14422 ( .A(n14031), .B(sreg[1355]), .Z(n14035) );
  OR U14423 ( .A(n14033), .B(n14032), .Z(n14034) );
  AND U14424 ( .A(n14035), .B(n14034), .Z(n14073) );
  XOR U14425 ( .A(n14074), .B(n14073), .Z(c[1356]) );
  NANDN U14426 ( .A(n14037), .B(n14036), .Z(n14041) );
  NAND U14427 ( .A(n14039), .B(n14038), .Z(n14040) );
  NAND U14428 ( .A(n14041), .B(n14040), .Z(n14080) );
  NAND U14429 ( .A(b[0]), .B(a[341]), .Z(n14042) );
  XNOR U14430 ( .A(b[1]), .B(n14042), .Z(n14044) );
  NAND U14431 ( .A(n63), .B(a[340]), .Z(n14043) );
  AND U14432 ( .A(n14044), .B(n14043), .Z(n14097) );
  XOR U14433 ( .A(a[337]), .B(n42197), .Z(n14086) );
  NANDN U14434 ( .A(n14086), .B(n42173), .Z(n14047) );
  NANDN U14435 ( .A(n14045), .B(n42172), .Z(n14046) );
  NAND U14436 ( .A(n14047), .B(n14046), .Z(n14095) );
  NAND U14437 ( .A(b[7]), .B(a[333]), .Z(n14096) );
  XNOR U14438 ( .A(n14095), .B(n14096), .Z(n14098) );
  XOR U14439 ( .A(n14097), .B(n14098), .Z(n14104) );
  NANDN U14440 ( .A(n14048), .B(n42093), .Z(n14050) );
  XOR U14441 ( .A(n42134), .B(a[339]), .Z(n14089) );
  NANDN U14442 ( .A(n14089), .B(n42095), .Z(n14049) );
  NAND U14443 ( .A(n14050), .B(n14049), .Z(n14102) );
  NANDN U14444 ( .A(n14051), .B(n42231), .Z(n14053) );
  XOR U14445 ( .A(n190), .B(a[335]), .Z(n14092) );
  NANDN U14446 ( .A(n14092), .B(n42234), .Z(n14052) );
  AND U14447 ( .A(n14053), .B(n14052), .Z(n14101) );
  XNOR U14448 ( .A(n14102), .B(n14101), .Z(n14103) );
  XNOR U14449 ( .A(n14104), .B(n14103), .Z(n14108) );
  NANDN U14450 ( .A(n14055), .B(n14054), .Z(n14059) );
  NAND U14451 ( .A(n14057), .B(n14056), .Z(n14058) );
  AND U14452 ( .A(n14059), .B(n14058), .Z(n14107) );
  XOR U14453 ( .A(n14108), .B(n14107), .Z(n14109) );
  NANDN U14454 ( .A(n14061), .B(n14060), .Z(n14065) );
  NANDN U14455 ( .A(n14063), .B(n14062), .Z(n14064) );
  NAND U14456 ( .A(n14065), .B(n14064), .Z(n14110) );
  XOR U14457 ( .A(n14109), .B(n14110), .Z(n14077) );
  OR U14458 ( .A(n14067), .B(n14066), .Z(n14071) );
  NANDN U14459 ( .A(n14069), .B(n14068), .Z(n14070) );
  NAND U14460 ( .A(n14071), .B(n14070), .Z(n14078) );
  XNOR U14461 ( .A(n14077), .B(n14078), .Z(n14079) );
  XNOR U14462 ( .A(n14080), .B(n14079), .Z(n14113) );
  XNOR U14463 ( .A(n14113), .B(sreg[1357]), .Z(n14115) );
  NAND U14464 ( .A(n14072), .B(sreg[1356]), .Z(n14076) );
  OR U14465 ( .A(n14074), .B(n14073), .Z(n14075) );
  AND U14466 ( .A(n14076), .B(n14075), .Z(n14114) );
  XOR U14467 ( .A(n14115), .B(n14114), .Z(c[1357]) );
  NANDN U14468 ( .A(n14078), .B(n14077), .Z(n14082) );
  NAND U14469 ( .A(n14080), .B(n14079), .Z(n14081) );
  NAND U14470 ( .A(n14082), .B(n14081), .Z(n14121) );
  NAND U14471 ( .A(b[0]), .B(a[342]), .Z(n14083) );
  XNOR U14472 ( .A(b[1]), .B(n14083), .Z(n14085) );
  NAND U14473 ( .A(n63), .B(a[341]), .Z(n14084) );
  AND U14474 ( .A(n14085), .B(n14084), .Z(n14138) );
  XOR U14475 ( .A(a[338]), .B(n42197), .Z(n14127) );
  NANDN U14476 ( .A(n14127), .B(n42173), .Z(n14088) );
  NANDN U14477 ( .A(n14086), .B(n42172), .Z(n14087) );
  NAND U14478 ( .A(n14088), .B(n14087), .Z(n14136) );
  NAND U14479 ( .A(b[7]), .B(a[334]), .Z(n14137) );
  XNOR U14480 ( .A(n14136), .B(n14137), .Z(n14139) );
  XOR U14481 ( .A(n14138), .B(n14139), .Z(n14145) );
  NANDN U14482 ( .A(n14089), .B(n42093), .Z(n14091) );
  XOR U14483 ( .A(n42134), .B(a[340]), .Z(n14130) );
  NANDN U14484 ( .A(n14130), .B(n42095), .Z(n14090) );
  NAND U14485 ( .A(n14091), .B(n14090), .Z(n14143) );
  NANDN U14486 ( .A(n14092), .B(n42231), .Z(n14094) );
  XOR U14487 ( .A(n190), .B(a[336]), .Z(n14133) );
  NANDN U14488 ( .A(n14133), .B(n42234), .Z(n14093) );
  AND U14489 ( .A(n14094), .B(n14093), .Z(n14142) );
  XNOR U14490 ( .A(n14143), .B(n14142), .Z(n14144) );
  XNOR U14491 ( .A(n14145), .B(n14144), .Z(n14149) );
  NANDN U14492 ( .A(n14096), .B(n14095), .Z(n14100) );
  NAND U14493 ( .A(n14098), .B(n14097), .Z(n14099) );
  AND U14494 ( .A(n14100), .B(n14099), .Z(n14148) );
  XOR U14495 ( .A(n14149), .B(n14148), .Z(n14150) );
  NANDN U14496 ( .A(n14102), .B(n14101), .Z(n14106) );
  NANDN U14497 ( .A(n14104), .B(n14103), .Z(n14105) );
  NAND U14498 ( .A(n14106), .B(n14105), .Z(n14151) );
  XOR U14499 ( .A(n14150), .B(n14151), .Z(n14118) );
  OR U14500 ( .A(n14108), .B(n14107), .Z(n14112) );
  NANDN U14501 ( .A(n14110), .B(n14109), .Z(n14111) );
  NAND U14502 ( .A(n14112), .B(n14111), .Z(n14119) );
  XNOR U14503 ( .A(n14118), .B(n14119), .Z(n14120) );
  XNOR U14504 ( .A(n14121), .B(n14120), .Z(n14154) );
  XNOR U14505 ( .A(n14154), .B(sreg[1358]), .Z(n14156) );
  NAND U14506 ( .A(n14113), .B(sreg[1357]), .Z(n14117) );
  OR U14507 ( .A(n14115), .B(n14114), .Z(n14116) );
  AND U14508 ( .A(n14117), .B(n14116), .Z(n14155) );
  XOR U14509 ( .A(n14156), .B(n14155), .Z(c[1358]) );
  NANDN U14510 ( .A(n14119), .B(n14118), .Z(n14123) );
  NAND U14511 ( .A(n14121), .B(n14120), .Z(n14122) );
  NAND U14512 ( .A(n14123), .B(n14122), .Z(n14162) );
  NAND U14513 ( .A(b[0]), .B(a[343]), .Z(n14124) );
  XNOR U14514 ( .A(b[1]), .B(n14124), .Z(n14126) );
  NAND U14515 ( .A(n64), .B(a[342]), .Z(n14125) );
  AND U14516 ( .A(n14126), .B(n14125), .Z(n14179) );
  XOR U14517 ( .A(a[339]), .B(n42197), .Z(n14168) );
  NANDN U14518 ( .A(n14168), .B(n42173), .Z(n14129) );
  NANDN U14519 ( .A(n14127), .B(n42172), .Z(n14128) );
  NAND U14520 ( .A(n14129), .B(n14128), .Z(n14177) );
  NAND U14521 ( .A(b[7]), .B(a[335]), .Z(n14178) );
  XNOR U14522 ( .A(n14177), .B(n14178), .Z(n14180) );
  XOR U14523 ( .A(n14179), .B(n14180), .Z(n14186) );
  NANDN U14524 ( .A(n14130), .B(n42093), .Z(n14132) );
  XOR U14525 ( .A(n42134), .B(a[341]), .Z(n14171) );
  NANDN U14526 ( .A(n14171), .B(n42095), .Z(n14131) );
  NAND U14527 ( .A(n14132), .B(n14131), .Z(n14184) );
  NANDN U14528 ( .A(n14133), .B(n42231), .Z(n14135) );
  XOR U14529 ( .A(n190), .B(a[337]), .Z(n14174) );
  NANDN U14530 ( .A(n14174), .B(n42234), .Z(n14134) );
  AND U14531 ( .A(n14135), .B(n14134), .Z(n14183) );
  XNOR U14532 ( .A(n14184), .B(n14183), .Z(n14185) );
  XNOR U14533 ( .A(n14186), .B(n14185), .Z(n14190) );
  NANDN U14534 ( .A(n14137), .B(n14136), .Z(n14141) );
  NAND U14535 ( .A(n14139), .B(n14138), .Z(n14140) );
  AND U14536 ( .A(n14141), .B(n14140), .Z(n14189) );
  XOR U14537 ( .A(n14190), .B(n14189), .Z(n14191) );
  NANDN U14538 ( .A(n14143), .B(n14142), .Z(n14147) );
  NANDN U14539 ( .A(n14145), .B(n14144), .Z(n14146) );
  NAND U14540 ( .A(n14147), .B(n14146), .Z(n14192) );
  XOR U14541 ( .A(n14191), .B(n14192), .Z(n14159) );
  OR U14542 ( .A(n14149), .B(n14148), .Z(n14153) );
  NANDN U14543 ( .A(n14151), .B(n14150), .Z(n14152) );
  NAND U14544 ( .A(n14153), .B(n14152), .Z(n14160) );
  XNOR U14545 ( .A(n14159), .B(n14160), .Z(n14161) );
  XNOR U14546 ( .A(n14162), .B(n14161), .Z(n14195) );
  XNOR U14547 ( .A(n14195), .B(sreg[1359]), .Z(n14197) );
  NAND U14548 ( .A(n14154), .B(sreg[1358]), .Z(n14158) );
  OR U14549 ( .A(n14156), .B(n14155), .Z(n14157) );
  AND U14550 ( .A(n14158), .B(n14157), .Z(n14196) );
  XOR U14551 ( .A(n14197), .B(n14196), .Z(c[1359]) );
  NANDN U14552 ( .A(n14160), .B(n14159), .Z(n14164) );
  NAND U14553 ( .A(n14162), .B(n14161), .Z(n14163) );
  NAND U14554 ( .A(n14164), .B(n14163), .Z(n14203) );
  NAND U14555 ( .A(b[0]), .B(a[344]), .Z(n14165) );
  XNOR U14556 ( .A(b[1]), .B(n14165), .Z(n14167) );
  NAND U14557 ( .A(n64), .B(a[343]), .Z(n14166) );
  AND U14558 ( .A(n14167), .B(n14166), .Z(n14220) );
  XOR U14559 ( .A(a[340]), .B(n42197), .Z(n14209) );
  NANDN U14560 ( .A(n14209), .B(n42173), .Z(n14170) );
  NANDN U14561 ( .A(n14168), .B(n42172), .Z(n14169) );
  NAND U14562 ( .A(n14170), .B(n14169), .Z(n14218) );
  NAND U14563 ( .A(b[7]), .B(a[336]), .Z(n14219) );
  XNOR U14564 ( .A(n14218), .B(n14219), .Z(n14221) );
  XOR U14565 ( .A(n14220), .B(n14221), .Z(n14227) );
  NANDN U14566 ( .A(n14171), .B(n42093), .Z(n14173) );
  XOR U14567 ( .A(n42134), .B(a[342]), .Z(n14212) );
  NANDN U14568 ( .A(n14212), .B(n42095), .Z(n14172) );
  NAND U14569 ( .A(n14173), .B(n14172), .Z(n14225) );
  NANDN U14570 ( .A(n14174), .B(n42231), .Z(n14176) );
  XOR U14571 ( .A(n190), .B(a[338]), .Z(n14215) );
  NANDN U14572 ( .A(n14215), .B(n42234), .Z(n14175) );
  AND U14573 ( .A(n14176), .B(n14175), .Z(n14224) );
  XNOR U14574 ( .A(n14225), .B(n14224), .Z(n14226) );
  XNOR U14575 ( .A(n14227), .B(n14226), .Z(n14231) );
  NANDN U14576 ( .A(n14178), .B(n14177), .Z(n14182) );
  NAND U14577 ( .A(n14180), .B(n14179), .Z(n14181) );
  AND U14578 ( .A(n14182), .B(n14181), .Z(n14230) );
  XOR U14579 ( .A(n14231), .B(n14230), .Z(n14232) );
  NANDN U14580 ( .A(n14184), .B(n14183), .Z(n14188) );
  NANDN U14581 ( .A(n14186), .B(n14185), .Z(n14187) );
  NAND U14582 ( .A(n14188), .B(n14187), .Z(n14233) );
  XOR U14583 ( .A(n14232), .B(n14233), .Z(n14200) );
  OR U14584 ( .A(n14190), .B(n14189), .Z(n14194) );
  NANDN U14585 ( .A(n14192), .B(n14191), .Z(n14193) );
  NAND U14586 ( .A(n14194), .B(n14193), .Z(n14201) );
  XNOR U14587 ( .A(n14200), .B(n14201), .Z(n14202) );
  XNOR U14588 ( .A(n14203), .B(n14202), .Z(n14236) );
  XNOR U14589 ( .A(n14236), .B(sreg[1360]), .Z(n14238) );
  NAND U14590 ( .A(n14195), .B(sreg[1359]), .Z(n14199) );
  OR U14591 ( .A(n14197), .B(n14196), .Z(n14198) );
  AND U14592 ( .A(n14199), .B(n14198), .Z(n14237) );
  XOR U14593 ( .A(n14238), .B(n14237), .Z(c[1360]) );
  NANDN U14594 ( .A(n14201), .B(n14200), .Z(n14205) );
  NAND U14595 ( .A(n14203), .B(n14202), .Z(n14204) );
  NAND U14596 ( .A(n14205), .B(n14204), .Z(n14244) );
  NAND U14597 ( .A(b[0]), .B(a[345]), .Z(n14206) );
  XNOR U14598 ( .A(b[1]), .B(n14206), .Z(n14208) );
  NAND U14599 ( .A(n64), .B(a[344]), .Z(n14207) );
  AND U14600 ( .A(n14208), .B(n14207), .Z(n14261) );
  XOR U14601 ( .A(a[341]), .B(n42197), .Z(n14250) );
  NANDN U14602 ( .A(n14250), .B(n42173), .Z(n14211) );
  NANDN U14603 ( .A(n14209), .B(n42172), .Z(n14210) );
  NAND U14604 ( .A(n14211), .B(n14210), .Z(n14259) );
  NAND U14605 ( .A(b[7]), .B(a[337]), .Z(n14260) );
  XNOR U14606 ( .A(n14259), .B(n14260), .Z(n14262) );
  XOR U14607 ( .A(n14261), .B(n14262), .Z(n14268) );
  NANDN U14608 ( .A(n14212), .B(n42093), .Z(n14214) );
  XOR U14609 ( .A(n42134), .B(a[343]), .Z(n14253) );
  NANDN U14610 ( .A(n14253), .B(n42095), .Z(n14213) );
  NAND U14611 ( .A(n14214), .B(n14213), .Z(n14266) );
  NANDN U14612 ( .A(n14215), .B(n42231), .Z(n14217) );
  XOR U14613 ( .A(n190), .B(a[339]), .Z(n14256) );
  NANDN U14614 ( .A(n14256), .B(n42234), .Z(n14216) );
  AND U14615 ( .A(n14217), .B(n14216), .Z(n14265) );
  XNOR U14616 ( .A(n14266), .B(n14265), .Z(n14267) );
  XNOR U14617 ( .A(n14268), .B(n14267), .Z(n14272) );
  NANDN U14618 ( .A(n14219), .B(n14218), .Z(n14223) );
  NAND U14619 ( .A(n14221), .B(n14220), .Z(n14222) );
  AND U14620 ( .A(n14223), .B(n14222), .Z(n14271) );
  XOR U14621 ( .A(n14272), .B(n14271), .Z(n14273) );
  NANDN U14622 ( .A(n14225), .B(n14224), .Z(n14229) );
  NANDN U14623 ( .A(n14227), .B(n14226), .Z(n14228) );
  NAND U14624 ( .A(n14229), .B(n14228), .Z(n14274) );
  XOR U14625 ( .A(n14273), .B(n14274), .Z(n14241) );
  OR U14626 ( .A(n14231), .B(n14230), .Z(n14235) );
  NANDN U14627 ( .A(n14233), .B(n14232), .Z(n14234) );
  NAND U14628 ( .A(n14235), .B(n14234), .Z(n14242) );
  XNOR U14629 ( .A(n14241), .B(n14242), .Z(n14243) );
  XNOR U14630 ( .A(n14244), .B(n14243), .Z(n14277) );
  XNOR U14631 ( .A(n14277), .B(sreg[1361]), .Z(n14279) );
  NAND U14632 ( .A(n14236), .B(sreg[1360]), .Z(n14240) );
  OR U14633 ( .A(n14238), .B(n14237), .Z(n14239) );
  AND U14634 ( .A(n14240), .B(n14239), .Z(n14278) );
  XOR U14635 ( .A(n14279), .B(n14278), .Z(c[1361]) );
  NANDN U14636 ( .A(n14242), .B(n14241), .Z(n14246) );
  NAND U14637 ( .A(n14244), .B(n14243), .Z(n14245) );
  NAND U14638 ( .A(n14246), .B(n14245), .Z(n14285) );
  NAND U14639 ( .A(b[0]), .B(a[346]), .Z(n14247) );
  XNOR U14640 ( .A(b[1]), .B(n14247), .Z(n14249) );
  NAND U14641 ( .A(n64), .B(a[345]), .Z(n14248) );
  AND U14642 ( .A(n14249), .B(n14248), .Z(n14302) );
  XOR U14643 ( .A(a[342]), .B(n42197), .Z(n14291) );
  NANDN U14644 ( .A(n14291), .B(n42173), .Z(n14252) );
  NANDN U14645 ( .A(n14250), .B(n42172), .Z(n14251) );
  NAND U14646 ( .A(n14252), .B(n14251), .Z(n14300) );
  NAND U14647 ( .A(b[7]), .B(a[338]), .Z(n14301) );
  XNOR U14648 ( .A(n14300), .B(n14301), .Z(n14303) );
  XOR U14649 ( .A(n14302), .B(n14303), .Z(n14309) );
  NANDN U14650 ( .A(n14253), .B(n42093), .Z(n14255) );
  XOR U14651 ( .A(n42134), .B(a[344]), .Z(n14294) );
  NANDN U14652 ( .A(n14294), .B(n42095), .Z(n14254) );
  NAND U14653 ( .A(n14255), .B(n14254), .Z(n14307) );
  NANDN U14654 ( .A(n14256), .B(n42231), .Z(n14258) );
  XOR U14655 ( .A(n190), .B(a[340]), .Z(n14297) );
  NANDN U14656 ( .A(n14297), .B(n42234), .Z(n14257) );
  AND U14657 ( .A(n14258), .B(n14257), .Z(n14306) );
  XNOR U14658 ( .A(n14307), .B(n14306), .Z(n14308) );
  XNOR U14659 ( .A(n14309), .B(n14308), .Z(n14313) );
  NANDN U14660 ( .A(n14260), .B(n14259), .Z(n14264) );
  NAND U14661 ( .A(n14262), .B(n14261), .Z(n14263) );
  AND U14662 ( .A(n14264), .B(n14263), .Z(n14312) );
  XOR U14663 ( .A(n14313), .B(n14312), .Z(n14314) );
  NANDN U14664 ( .A(n14266), .B(n14265), .Z(n14270) );
  NANDN U14665 ( .A(n14268), .B(n14267), .Z(n14269) );
  NAND U14666 ( .A(n14270), .B(n14269), .Z(n14315) );
  XOR U14667 ( .A(n14314), .B(n14315), .Z(n14282) );
  OR U14668 ( .A(n14272), .B(n14271), .Z(n14276) );
  NANDN U14669 ( .A(n14274), .B(n14273), .Z(n14275) );
  NAND U14670 ( .A(n14276), .B(n14275), .Z(n14283) );
  XNOR U14671 ( .A(n14282), .B(n14283), .Z(n14284) );
  XNOR U14672 ( .A(n14285), .B(n14284), .Z(n14318) );
  XNOR U14673 ( .A(n14318), .B(sreg[1362]), .Z(n14320) );
  NAND U14674 ( .A(n14277), .B(sreg[1361]), .Z(n14281) );
  OR U14675 ( .A(n14279), .B(n14278), .Z(n14280) );
  AND U14676 ( .A(n14281), .B(n14280), .Z(n14319) );
  XOR U14677 ( .A(n14320), .B(n14319), .Z(c[1362]) );
  NANDN U14678 ( .A(n14283), .B(n14282), .Z(n14287) );
  NAND U14679 ( .A(n14285), .B(n14284), .Z(n14286) );
  NAND U14680 ( .A(n14287), .B(n14286), .Z(n14326) );
  NAND U14681 ( .A(b[0]), .B(a[347]), .Z(n14288) );
  XNOR U14682 ( .A(b[1]), .B(n14288), .Z(n14290) );
  NAND U14683 ( .A(n64), .B(a[346]), .Z(n14289) );
  AND U14684 ( .A(n14290), .B(n14289), .Z(n14343) );
  XOR U14685 ( .A(a[343]), .B(n42197), .Z(n14332) );
  NANDN U14686 ( .A(n14332), .B(n42173), .Z(n14293) );
  NANDN U14687 ( .A(n14291), .B(n42172), .Z(n14292) );
  NAND U14688 ( .A(n14293), .B(n14292), .Z(n14341) );
  NAND U14689 ( .A(b[7]), .B(a[339]), .Z(n14342) );
  XNOR U14690 ( .A(n14341), .B(n14342), .Z(n14344) );
  XOR U14691 ( .A(n14343), .B(n14344), .Z(n14350) );
  NANDN U14692 ( .A(n14294), .B(n42093), .Z(n14296) );
  XOR U14693 ( .A(n42134), .B(a[345]), .Z(n14335) );
  NANDN U14694 ( .A(n14335), .B(n42095), .Z(n14295) );
  NAND U14695 ( .A(n14296), .B(n14295), .Z(n14348) );
  NANDN U14696 ( .A(n14297), .B(n42231), .Z(n14299) );
  XOR U14697 ( .A(n190), .B(a[341]), .Z(n14338) );
  NANDN U14698 ( .A(n14338), .B(n42234), .Z(n14298) );
  AND U14699 ( .A(n14299), .B(n14298), .Z(n14347) );
  XNOR U14700 ( .A(n14348), .B(n14347), .Z(n14349) );
  XNOR U14701 ( .A(n14350), .B(n14349), .Z(n14354) );
  NANDN U14702 ( .A(n14301), .B(n14300), .Z(n14305) );
  NAND U14703 ( .A(n14303), .B(n14302), .Z(n14304) );
  AND U14704 ( .A(n14305), .B(n14304), .Z(n14353) );
  XOR U14705 ( .A(n14354), .B(n14353), .Z(n14355) );
  NANDN U14706 ( .A(n14307), .B(n14306), .Z(n14311) );
  NANDN U14707 ( .A(n14309), .B(n14308), .Z(n14310) );
  NAND U14708 ( .A(n14311), .B(n14310), .Z(n14356) );
  XOR U14709 ( .A(n14355), .B(n14356), .Z(n14323) );
  OR U14710 ( .A(n14313), .B(n14312), .Z(n14317) );
  NANDN U14711 ( .A(n14315), .B(n14314), .Z(n14316) );
  NAND U14712 ( .A(n14317), .B(n14316), .Z(n14324) );
  XNOR U14713 ( .A(n14323), .B(n14324), .Z(n14325) );
  XNOR U14714 ( .A(n14326), .B(n14325), .Z(n14359) );
  XNOR U14715 ( .A(n14359), .B(sreg[1363]), .Z(n14361) );
  NAND U14716 ( .A(n14318), .B(sreg[1362]), .Z(n14322) );
  OR U14717 ( .A(n14320), .B(n14319), .Z(n14321) );
  AND U14718 ( .A(n14322), .B(n14321), .Z(n14360) );
  XOR U14719 ( .A(n14361), .B(n14360), .Z(c[1363]) );
  NANDN U14720 ( .A(n14324), .B(n14323), .Z(n14328) );
  NAND U14721 ( .A(n14326), .B(n14325), .Z(n14327) );
  NAND U14722 ( .A(n14328), .B(n14327), .Z(n14367) );
  NAND U14723 ( .A(b[0]), .B(a[348]), .Z(n14329) );
  XNOR U14724 ( .A(b[1]), .B(n14329), .Z(n14331) );
  NAND U14725 ( .A(n64), .B(a[347]), .Z(n14330) );
  AND U14726 ( .A(n14331), .B(n14330), .Z(n14384) );
  XOR U14727 ( .A(a[344]), .B(n42197), .Z(n14373) );
  NANDN U14728 ( .A(n14373), .B(n42173), .Z(n14334) );
  NANDN U14729 ( .A(n14332), .B(n42172), .Z(n14333) );
  NAND U14730 ( .A(n14334), .B(n14333), .Z(n14382) );
  NAND U14731 ( .A(b[7]), .B(a[340]), .Z(n14383) );
  XNOR U14732 ( .A(n14382), .B(n14383), .Z(n14385) );
  XOR U14733 ( .A(n14384), .B(n14385), .Z(n14391) );
  NANDN U14734 ( .A(n14335), .B(n42093), .Z(n14337) );
  XOR U14735 ( .A(n42134), .B(a[346]), .Z(n14376) );
  NANDN U14736 ( .A(n14376), .B(n42095), .Z(n14336) );
  NAND U14737 ( .A(n14337), .B(n14336), .Z(n14389) );
  NANDN U14738 ( .A(n14338), .B(n42231), .Z(n14340) );
  XOR U14739 ( .A(n190), .B(a[342]), .Z(n14379) );
  NANDN U14740 ( .A(n14379), .B(n42234), .Z(n14339) );
  AND U14741 ( .A(n14340), .B(n14339), .Z(n14388) );
  XNOR U14742 ( .A(n14389), .B(n14388), .Z(n14390) );
  XNOR U14743 ( .A(n14391), .B(n14390), .Z(n14395) );
  NANDN U14744 ( .A(n14342), .B(n14341), .Z(n14346) );
  NAND U14745 ( .A(n14344), .B(n14343), .Z(n14345) );
  AND U14746 ( .A(n14346), .B(n14345), .Z(n14394) );
  XOR U14747 ( .A(n14395), .B(n14394), .Z(n14396) );
  NANDN U14748 ( .A(n14348), .B(n14347), .Z(n14352) );
  NANDN U14749 ( .A(n14350), .B(n14349), .Z(n14351) );
  NAND U14750 ( .A(n14352), .B(n14351), .Z(n14397) );
  XOR U14751 ( .A(n14396), .B(n14397), .Z(n14364) );
  OR U14752 ( .A(n14354), .B(n14353), .Z(n14358) );
  NANDN U14753 ( .A(n14356), .B(n14355), .Z(n14357) );
  NAND U14754 ( .A(n14358), .B(n14357), .Z(n14365) );
  XNOR U14755 ( .A(n14364), .B(n14365), .Z(n14366) );
  XNOR U14756 ( .A(n14367), .B(n14366), .Z(n14400) );
  XNOR U14757 ( .A(n14400), .B(sreg[1364]), .Z(n14402) );
  NAND U14758 ( .A(n14359), .B(sreg[1363]), .Z(n14363) );
  OR U14759 ( .A(n14361), .B(n14360), .Z(n14362) );
  AND U14760 ( .A(n14363), .B(n14362), .Z(n14401) );
  XOR U14761 ( .A(n14402), .B(n14401), .Z(c[1364]) );
  NANDN U14762 ( .A(n14365), .B(n14364), .Z(n14369) );
  NAND U14763 ( .A(n14367), .B(n14366), .Z(n14368) );
  NAND U14764 ( .A(n14369), .B(n14368), .Z(n14408) );
  NAND U14765 ( .A(b[0]), .B(a[349]), .Z(n14370) );
  XNOR U14766 ( .A(b[1]), .B(n14370), .Z(n14372) );
  NAND U14767 ( .A(n64), .B(a[348]), .Z(n14371) );
  AND U14768 ( .A(n14372), .B(n14371), .Z(n14425) );
  XOR U14769 ( .A(a[345]), .B(n42197), .Z(n14414) );
  NANDN U14770 ( .A(n14414), .B(n42173), .Z(n14375) );
  NANDN U14771 ( .A(n14373), .B(n42172), .Z(n14374) );
  NAND U14772 ( .A(n14375), .B(n14374), .Z(n14423) );
  NAND U14773 ( .A(b[7]), .B(a[341]), .Z(n14424) );
  XNOR U14774 ( .A(n14423), .B(n14424), .Z(n14426) );
  XOR U14775 ( .A(n14425), .B(n14426), .Z(n14432) );
  NANDN U14776 ( .A(n14376), .B(n42093), .Z(n14378) );
  XOR U14777 ( .A(n42134), .B(a[347]), .Z(n14417) );
  NANDN U14778 ( .A(n14417), .B(n42095), .Z(n14377) );
  NAND U14779 ( .A(n14378), .B(n14377), .Z(n14430) );
  NANDN U14780 ( .A(n14379), .B(n42231), .Z(n14381) );
  XOR U14781 ( .A(n190), .B(a[343]), .Z(n14420) );
  NANDN U14782 ( .A(n14420), .B(n42234), .Z(n14380) );
  AND U14783 ( .A(n14381), .B(n14380), .Z(n14429) );
  XNOR U14784 ( .A(n14430), .B(n14429), .Z(n14431) );
  XNOR U14785 ( .A(n14432), .B(n14431), .Z(n14436) );
  NANDN U14786 ( .A(n14383), .B(n14382), .Z(n14387) );
  NAND U14787 ( .A(n14385), .B(n14384), .Z(n14386) );
  AND U14788 ( .A(n14387), .B(n14386), .Z(n14435) );
  XOR U14789 ( .A(n14436), .B(n14435), .Z(n14437) );
  NANDN U14790 ( .A(n14389), .B(n14388), .Z(n14393) );
  NANDN U14791 ( .A(n14391), .B(n14390), .Z(n14392) );
  NAND U14792 ( .A(n14393), .B(n14392), .Z(n14438) );
  XOR U14793 ( .A(n14437), .B(n14438), .Z(n14405) );
  OR U14794 ( .A(n14395), .B(n14394), .Z(n14399) );
  NANDN U14795 ( .A(n14397), .B(n14396), .Z(n14398) );
  NAND U14796 ( .A(n14399), .B(n14398), .Z(n14406) );
  XNOR U14797 ( .A(n14405), .B(n14406), .Z(n14407) );
  XNOR U14798 ( .A(n14408), .B(n14407), .Z(n14441) );
  XNOR U14799 ( .A(n14441), .B(sreg[1365]), .Z(n14443) );
  NAND U14800 ( .A(n14400), .B(sreg[1364]), .Z(n14404) );
  OR U14801 ( .A(n14402), .B(n14401), .Z(n14403) );
  AND U14802 ( .A(n14404), .B(n14403), .Z(n14442) );
  XOR U14803 ( .A(n14443), .B(n14442), .Z(c[1365]) );
  NANDN U14804 ( .A(n14406), .B(n14405), .Z(n14410) );
  NAND U14805 ( .A(n14408), .B(n14407), .Z(n14409) );
  NAND U14806 ( .A(n14410), .B(n14409), .Z(n14449) );
  NAND U14807 ( .A(b[0]), .B(a[350]), .Z(n14411) );
  XNOR U14808 ( .A(b[1]), .B(n14411), .Z(n14413) );
  NAND U14809 ( .A(n65), .B(a[349]), .Z(n14412) );
  AND U14810 ( .A(n14413), .B(n14412), .Z(n14466) );
  XOR U14811 ( .A(a[346]), .B(n42197), .Z(n14455) );
  NANDN U14812 ( .A(n14455), .B(n42173), .Z(n14416) );
  NANDN U14813 ( .A(n14414), .B(n42172), .Z(n14415) );
  NAND U14814 ( .A(n14416), .B(n14415), .Z(n14464) );
  NAND U14815 ( .A(b[7]), .B(a[342]), .Z(n14465) );
  XNOR U14816 ( .A(n14464), .B(n14465), .Z(n14467) );
  XOR U14817 ( .A(n14466), .B(n14467), .Z(n14473) );
  NANDN U14818 ( .A(n14417), .B(n42093), .Z(n14419) );
  XOR U14819 ( .A(n42134), .B(a[348]), .Z(n14458) );
  NANDN U14820 ( .A(n14458), .B(n42095), .Z(n14418) );
  NAND U14821 ( .A(n14419), .B(n14418), .Z(n14471) );
  NANDN U14822 ( .A(n14420), .B(n42231), .Z(n14422) );
  XOR U14823 ( .A(n190), .B(a[344]), .Z(n14461) );
  NANDN U14824 ( .A(n14461), .B(n42234), .Z(n14421) );
  AND U14825 ( .A(n14422), .B(n14421), .Z(n14470) );
  XNOR U14826 ( .A(n14471), .B(n14470), .Z(n14472) );
  XNOR U14827 ( .A(n14473), .B(n14472), .Z(n14477) );
  NANDN U14828 ( .A(n14424), .B(n14423), .Z(n14428) );
  NAND U14829 ( .A(n14426), .B(n14425), .Z(n14427) );
  AND U14830 ( .A(n14428), .B(n14427), .Z(n14476) );
  XOR U14831 ( .A(n14477), .B(n14476), .Z(n14478) );
  NANDN U14832 ( .A(n14430), .B(n14429), .Z(n14434) );
  NANDN U14833 ( .A(n14432), .B(n14431), .Z(n14433) );
  NAND U14834 ( .A(n14434), .B(n14433), .Z(n14479) );
  XOR U14835 ( .A(n14478), .B(n14479), .Z(n14446) );
  OR U14836 ( .A(n14436), .B(n14435), .Z(n14440) );
  NANDN U14837 ( .A(n14438), .B(n14437), .Z(n14439) );
  NAND U14838 ( .A(n14440), .B(n14439), .Z(n14447) );
  XNOR U14839 ( .A(n14446), .B(n14447), .Z(n14448) );
  XNOR U14840 ( .A(n14449), .B(n14448), .Z(n14482) );
  XNOR U14841 ( .A(n14482), .B(sreg[1366]), .Z(n14484) );
  NAND U14842 ( .A(n14441), .B(sreg[1365]), .Z(n14445) );
  OR U14843 ( .A(n14443), .B(n14442), .Z(n14444) );
  AND U14844 ( .A(n14445), .B(n14444), .Z(n14483) );
  XOR U14845 ( .A(n14484), .B(n14483), .Z(c[1366]) );
  NANDN U14846 ( .A(n14447), .B(n14446), .Z(n14451) );
  NAND U14847 ( .A(n14449), .B(n14448), .Z(n14450) );
  NAND U14848 ( .A(n14451), .B(n14450), .Z(n14490) );
  NAND U14849 ( .A(b[0]), .B(a[351]), .Z(n14452) );
  XNOR U14850 ( .A(b[1]), .B(n14452), .Z(n14454) );
  NAND U14851 ( .A(n65), .B(a[350]), .Z(n14453) );
  AND U14852 ( .A(n14454), .B(n14453), .Z(n14507) );
  XOR U14853 ( .A(a[347]), .B(n42197), .Z(n14496) );
  NANDN U14854 ( .A(n14496), .B(n42173), .Z(n14457) );
  NANDN U14855 ( .A(n14455), .B(n42172), .Z(n14456) );
  NAND U14856 ( .A(n14457), .B(n14456), .Z(n14505) );
  NAND U14857 ( .A(b[7]), .B(a[343]), .Z(n14506) );
  XNOR U14858 ( .A(n14505), .B(n14506), .Z(n14508) );
  XOR U14859 ( .A(n14507), .B(n14508), .Z(n14514) );
  NANDN U14860 ( .A(n14458), .B(n42093), .Z(n14460) );
  XOR U14861 ( .A(n42134), .B(a[349]), .Z(n14499) );
  NANDN U14862 ( .A(n14499), .B(n42095), .Z(n14459) );
  NAND U14863 ( .A(n14460), .B(n14459), .Z(n14512) );
  NANDN U14864 ( .A(n14461), .B(n42231), .Z(n14463) );
  XOR U14865 ( .A(n190), .B(a[345]), .Z(n14502) );
  NANDN U14866 ( .A(n14502), .B(n42234), .Z(n14462) );
  AND U14867 ( .A(n14463), .B(n14462), .Z(n14511) );
  XNOR U14868 ( .A(n14512), .B(n14511), .Z(n14513) );
  XNOR U14869 ( .A(n14514), .B(n14513), .Z(n14518) );
  NANDN U14870 ( .A(n14465), .B(n14464), .Z(n14469) );
  NAND U14871 ( .A(n14467), .B(n14466), .Z(n14468) );
  AND U14872 ( .A(n14469), .B(n14468), .Z(n14517) );
  XOR U14873 ( .A(n14518), .B(n14517), .Z(n14519) );
  NANDN U14874 ( .A(n14471), .B(n14470), .Z(n14475) );
  NANDN U14875 ( .A(n14473), .B(n14472), .Z(n14474) );
  NAND U14876 ( .A(n14475), .B(n14474), .Z(n14520) );
  XOR U14877 ( .A(n14519), .B(n14520), .Z(n14487) );
  OR U14878 ( .A(n14477), .B(n14476), .Z(n14481) );
  NANDN U14879 ( .A(n14479), .B(n14478), .Z(n14480) );
  NAND U14880 ( .A(n14481), .B(n14480), .Z(n14488) );
  XNOR U14881 ( .A(n14487), .B(n14488), .Z(n14489) );
  XNOR U14882 ( .A(n14490), .B(n14489), .Z(n14523) );
  XNOR U14883 ( .A(n14523), .B(sreg[1367]), .Z(n14525) );
  NAND U14884 ( .A(n14482), .B(sreg[1366]), .Z(n14486) );
  OR U14885 ( .A(n14484), .B(n14483), .Z(n14485) );
  AND U14886 ( .A(n14486), .B(n14485), .Z(n14524) );
  XOR U14887 ( .A(n14525), .B(n14524), .Z(c[1367]) );
  NANDN U14888 ( .A(n14488), .B(n14487), .Z(n14492) );
  NAND U14889 ( .A(n14490), .B(n14489), .Z(n14491) );
  NAND U14890 ( .A(n14492), .B(n14491), .Z(n14531) );
  NAND U14891 ( .A(b[0]), .B(a[352]), .Z(n14493) );
  XNOR U14892 ( .A(b[1]), .B(n14493), .Z(n14495) );
  NAND U14893 ( .A(n65), .B(a[351]), .Z(n14494) );
  AND U14894 ( .A(n14495), .B(n14494), .Z(n14548) );
  XOR U14895 ( .A(a[348]), .B(n42197), .Z(n14537) );
  NANDN U14896 ( .A(n14537), .B(n42173), .Z(n14498) );
  NANDN U14897 ( .A(n14496), .B(n42172), .Z(n14497) );
  NAND U14898 ( .A(n14498), .B(n14497), .Z(n14546) );
  NAND U14899 ( .A(b[7]), .B(a[344]), .Z(n14547) );
  XNOR U14900 ( .A(n14546), .B(n14547), .Z(n14549) );
  XOR U14901 ( .A(n14548), .B(n14549), .Z(n14555) );
  NANDN U14902 ( .A(n14499), .B(n42093), .Z(n14501) );
  XOR U14903 ( .A(n42134), .B(a[350]), .Z(n14540) );
  NANDN U14904 ( .A(n14540), .B(n42095), .Z(n14500) );
  NAND U14905 ( .A(n14501), .B(n14500), .Z(n14553) );
  NANDN U14906 ( .A(n14502), .B(n42231), .Z(n14504) );
  XOR U14907 ( .A(n190), .B(a[346]), .Z(n14543) );
  NANDN U14908 ( .A(n14543), .B(n42234), .Z(n14503) );
  AND U14909 ( .A(n14504), .B(n14503), .Z(n14552) );
  XNOR U14910 ( .A(n14553), .B(n14552), .Z(n14554) );
  XNOR U14911 ( .A(n14555), .B(n14554), .Z(n14559) );
  NANDN U14912 ( .A(n14506), .B(n14505), .Z(n14510) );
  NAND U14913 ( .A(n14508), .B(n14507), .Z(n14509) );
  AND U14914 ( .A(n14510), .B(n14509), .Z(n14558) );
  XOR U14915 ( .A(n14559), .B(n14558), .Z(n14560) );
  NANDN U14916 ( .A(n14512), .B(n14511), .Z(n14516) );
  NANDN U14917 ( .A(n14514), .B(n14513), .Z(n14515) );
  NAND U14918 ( .A(n14516), .B(n14515), .Z(n14561) );
  XOR U14919 ( .A(n14560), .B(n14561), .Z(n14528) );
  OR U14920 ( .A(n14518), .B(n14517), .Z(n14522) );
  NANDN U14921 ( .A(n14520), .B(n14519), .Z(n14521) );
  NAND U14922 ( .A(n14522), .B(n14521), .Z(n14529) );
  XNOR U14923 ( .A(n14528), .B(n14529), .Z(n14530) );
  XNOR U14924 ( .A(n14531), .B(n14530), .Z(n14564) );
  XNOR U14925 ( .A(n14564), .B(sreg[1368]), .Z(n14566) );
  NAND U14926 ( .A(n14523), .B(sreg[1367]), .Z(n14527) );
  OR U14927 ( .A(n14525), .B(n14524), .Z(n14526) );
  AND U14928 ( .A(n14527), .B(n14526), .Z(n14565) );
  XOR U14929 ( .A(n14566), .B(n14565), .Z(c[1368]) );
  NANDN U14930 ( .A(n14529), .B(n14528), .Z(n14533) );
  NAND U14931 ( .A(n14531), .B(n14530), .Z(n14532) );
  NAND U14932 ( .A(n14533), .B(n14532), .Z(n14572) );
  NAND U14933 ( .A(b[0]), .B(a[353]), .Z(n14534) );
  XNOR U14934 ( .A(b[1]), .B(n14534), .Z(n14536) );
  NAND U14935 ( .A(n65), .B(a[352]), .Z(n14535) );
  AND U14936 ( .A(n14536), .B(n14535), .Z(n14589) );
  XOR U14937 ( .A(a[349]), .B(n42197), .Z(n14578) );
  NANDN U14938 ( .A(n14578), .B(n42173), .Z(n14539) );
  NANDN U14939 ( .A(n14537), .B(n42172), .Z(n14538) );
  NAND U14940 ( .A(n14539), .B(n14538), .Z(n14587) );
  NAND U14941 ( .A(b[7]), .B(a[345]), .Z(n14588) );
  XNOR U14942 ( .A(n14587), .B(n14588), .Z(n14590) );
  XOR U14943 ( .A(n14589), .B(n14590), .Z(n14596) );
  NANDN U14944 ( .A(n14540), .B(n42093), .Z(n14542) );
  XOR U14945 ( .A(n42134), .B(a[351]), .Z(n14581) );
  NANDN U14946 ( .A(n14581), .B(n42095), .Z(n14541) );
  NAND U14947 ( .A(n14542), .B(n14541), .Z(n14594) );
  NANDN U14948 ( .A(n14543), .B(n42231), .Z(n14545) );
  XOR U14949 ( .A(n191), .B(a[347]), .Z(n14584) );
  NANDN U14950 ( .A(n14584), .B(n42234), .Z(n14544) );
  AND U14951 ( .A(n14545), .B(n14544), .Z(n14593) );
  XNOR U14952 ( .A(n14594), .B(n14593), .Z(n14595) );
  XNOR U14953 ( .A(n14596), .B(n14595), .Z(n14600) );
  NANDN U14954 ( .A(n14547), .B(n14546), .Z(n14551) );
  NAND U14955 ( .A(n14549), .B(n14548), .Z(n14550) );
  AND U14956 ( .A(n14551), .B(n14550), .Z(n14599) );
  XOR U14957 ( .A(n14600), .B(n14599), .Z(n14601) );
  NANDN U14958 ( .A(n14553), .B(n14552), .Z(n14557) );
  NANDN U14959 ( .A(n14555), .B(n14554), .Z(n14556) );
  NAND U14960 ( .A(n14557), .B(n14556), .Z(n14602) );
  XOR U14961 ( .A(n14601), .B(n14602), .Z(n14569) );
  OR U14962 ( .A(n14559), .B(n14558), .Z(n14563) );
  NANDN U14963 ( .A(n14561), .B(n14560), .Z(n14562) );
  NAND U14964 ( .A(n14563), .B(n14562), .Z(n14570) );
  XNOR U14965 ( .A(n14569), .B(n14570), .Z(n14571) );
  XNOR U14966 ( .A(n14572), .B(n14571), .Z(n14605) );
  XNOR U14967 ( .A(n14605), .B(sreg[1369]), .Z(n14607) );
  NAND U14968 ( .A(n14564), .B(sreg[1368]), .Z(n14568) );
  OR U14969 ( .A(n14566), .B(n14565), .Z(n14567) );
  AND U14970 ( .A(n14568), .B(n14567), .Z(n14606) );
  XOR U14971 ( .A(n14607), .B(n14606), .Z(c[1369]) );
  NANDN U14972 ( .A(n14570), .B(n14569), .Z(n14574) );
  NAND U14973 ( .A(n14572), .B(n14571), .Z(n14573) );
  NAND U14974 ( .A(n14574), .B(n14573), .Z(n14613) );
  NAND U14975 ( .A(b[0]), .B(a[354]), .Z(n14575) );
  XNOR U14976 ( .A(b[1]), .B(n14575), .Z(n14577) );
  NAND U14977 ( .A(n65), .B(a[353]), .Z(n14576) );
  AND U14978 ( .A(n14577), .B(n14576), .Z(n14630) );
  XOR U14979 ( .A(a[350]), .B(n42197), .Z(n14619) );
  NANDN U14980 ( .A(n14619), .B(n42173), .Z(n14580) );
  NANDN U14981 ( .A(n14578), .B(n42172), .Z(n14579) );
  NAND U14982 ( .A(n14580), .B(n14579), .Z(n14628) );
  NAND U14983 ( .A(b[7]), .B(a[346]), .Z(n14629) );
  XNOR U14984 ( .A(n14628), .B(n14629), .Z(n14631) );
  XOR U14985 ( .A(n14630), .B(n14631), .Z(n14637) );
  NANDN U14986 ( .A(n14581), .B(n42093), .Z(n14583) );
  XOR U14987 ( .A(n42134), .B(a[352]), .Z(n14622) );
  NANDN U14988 ( .A(n14622), .B(n42095), .Z(n14582) );
  NAND U14989 ( .A(n14583), .B(n14582), .Z(n14635) );
  NANDN U14990 ( .A(n14584), .B(n42231), .Z(n14586) );
  XOR U14991 ( .A(n191), .B(a[348]), .Z(n14625) );
  NANDN U14992 ( .A(n14625), .B(n42234), .Z(n14585) );
  AND U14993 ( .A(n14586), .B(n14585), .Z(n14634) );
  XNOR U14994 ( .A(n14635), .B(n14634), .Z(n14636) );
  XNOR U14995 ( .A(n14637), .B(n14636), .Z(n14641) );
  NANDN U14996 ( .A(n14588), .B(n14587), .Z(n14592) );
  NAND U14997 ( .A(n14590), .B(n14589), .Z(n14591) );
  AND U14998 ( .A(n14592), .B(n14591), .Z(n14640) );
  XOR U14999 ( .A(n14641), .B(n14640), .Z(n14642) );
  NANDN U15000 ( .A(n14594), .B(n14593), .Z(n14598) );
  NANDN U15001 ( .A(n14596), .B(n14595), .Z(n14597) );
  NAND U15002 ( .A(n14598), .B(n14597), .Z(n14643) );
  XOR U15003 ( .A(n14642), .B(n14643), .Z(n14610) );
  OR U15004 ( .A(n14600), .B(n14599), .Z(n14604) );
  NANDN U15005 ( .A(n14602), .B(n14601), .Z(n14603) );
  NAND U15006 ( .A(n14604), .B(n14603), .Z(n14611) );
  XNOR U15007 ( .A(n14610), .B(n14611), .Z(n14612) );
  XNOR U15008 ( .A(n14613), .B(n14612), .Z(n14646) );
  XNOR U15009 ( .A(n14646), .B(sreg[1370]), .Z(n14648) );
  NAND U15010 ( .A(n14605), .B(sreg[1369]), .Z(n14609) );
  OR U15011 ( .A(n14607), .B(n14606), .Z(n14608) );
  AND U15012 ( .A(n14609), .B(n14608), .Z(n14647) );
  XOR U15013 ( .A(n14648), .B(n14647), .Z(c[1370]) );
  NANDN U15014 ( .A(n14611), .B(n14610), .Z(n14615) );
  NAND U15015 ( .A(n14613), .B(n14612), .Z(n14614) );
  NAND U15016 ( .A(n14615), .B(n14614), .Z(n14654) );
  NAND U15017 ( .A(b[0]), .B(a[355]), .Z(n14616) );
  XNOR U15018 ( .A(b[1]), .B(n14616), .Z(n14618) );
  NAND U15019 ( .A(n65), .B(a[354]), .Z(n14617) );
  AND U15020 ( .A(n14618), .B(n14617), .Z(n14671) );
  XOR U15021 ( .A(a[351]), .B(n42197), .Z(n14660) );
  NANDN U15022 ( .A(n14660), .B(n42173), .Z(n14621) );
  NANDN U15023 ( .A(n14619), .B(n42172), .Z(n14620) );
  NAND U15024 ( .A(n14621), .B(n14620), .Z(n14669) );
  NAND U15025 ( .A(b[7]), .B(a[347]), .Z(n14670) );
  XNOR U15026 ( .A(n14669), .B(n14670), .Z(n14672) );
  XOR U15027 ( .A(n14671), .B(n14672), .Z(n14678) );
  NANDN U15028 ( .A(n14622), .B(n42093), .Z(n14624) );
  XOR U15029 ( .A(n42134), .B(a[353]), .Z(n14663) );
  NANDN U15030 ( .A(n14663), .B(n42095), .Z(n14623) );
  NAND U15031 ( .A(n14624), .B(n14623), .Z(n14676) );
  NANDN U15032 ( .A(n14625), .B(n42231), .Z(n14627) );
  XOR U15033 ( .A(n191), .B(a[349]), .Z(n14666) );
  NANDN U15034 ( .A(n14666), .B(n42234), .Z(n14626) );
  AND U15035 ( .A(n14627), .B(n14626), .Z(n14675) );
  XNOR U15036 ( .A(n14676), .B(n14675), .Z(n14677) );
  XNOR U15037 ( .A(n14678), .B(n14677), .Z(n14682) );
  NANDN U15038 ( .A(n14629), .B(n14628), .Z(n14633) );
  NAND U15039 ( .A(n14631), .B(n14630), .Z(n14632) );
  AND U15040 ( .A(n14633), .B(n14632), .Z(n14681) );
  XOR U15041 ( .A(n14682), .B(n14681), .Z(n14683) );
  NANDN U15042 ( .A(n14635), .B(n14634), .Z(n14639) );
  NANDN U15043 ( .A(n14637), .B(n14636), .Z(n14638) );
  NAND U15044 ( .A(n14639), .B(n14638), .Z(n14684) );
  XOR U15045 ( .A(n14683), .B(n14684), .Z(n14651) );
  OR U15046 ( .A(n14641), .B(n14640), .Z(n14645) );
  NANDN U15047 ( .A(n14643), .B(n14642), .Z(n14644) );
  NAND U15048 ( .A(n14645), .B(n14644), .Z(n14652) );
  XNOR U15049 ( .A(n14651), .B(n14652), .Z(n14653) );
  XNOR U15050 ( .A(n14654), .B(n14653), .Z(n14687) );
  XNOR U15051 ( .A(n14687), .B(sreg[1371]), .Z(n14689) );
  NAND U15052 ( .A(n14646), .B(sreg[1370]), .Z(n14650) );
  OR U15053 ( .A(n14648), .B(n14647), .Z(n14649) );
  AND U15054 ( .A(n14650), .B(n14649), .Z(n14688) );
  XOR U15055 ( .A(n14689), .B(n14688), .Z(c[1371]) );
  NANDN U15056 ( .A(n14652), .B(n14651), .Z(n14656) );
  NAND U15057 ( .A(n14654), .B(n14653), .Z(n14655) );
  NAND U15058 ( .A(n14656), .B(n14655), .Z(n14695) );
  NAND U15059 ( .A(b[0]), .B(a[356]), .Z(n14657) );
  XNOR U15060 ( .A(b[1]), .B(n14657), .Z(n14659) );
  NAND U15061 ( .A(n65), .B(a[355]), .Z(n14658) );
  AND U15062 ( .A(n14659), .B(n14658), .Z(n14712) );
  XOR U15063 ( .A(a[352]), .B(n42197), .Z(n14701) );
  NANDN U15064 ( .A(n14701), .B(n42173), .Z(n14662) );
  NANDN U15065 ( .A(n14660), .B(n42172), .Z(n14661) );
  NAND U15066 ( .A(n14662), .B(n14661), .Z(n14710) );
  NAND U15067 ( .A(b[7]), .B(a[348]), .Z(n14711) );
  XNOR U15068 ( .A(n14710), .B(n14711), .Z(n14713) );
  XOR U15069 ( .A(n14712), .B(n14713), .Z(n14719) );
  NANDN U15070 ( .A(n14663), .B(n42093), .Z(n14665) );
  XOR U15071 ( .A(n42134), .B(a[354]), .Z(n14704) );
  NANDN U15072 ( .A(n14704), .B(n42095), .Z(n14664) );
  NAND U15073 ( .A(n14665), .B(n14664), .Z(n14717) );
  NANDN U15074 ( .A(n14666), .B(n42231), .Z(n14668) );
  XOR U15075 ( .A(n191), .B(a[350]), .Z(n14707) );
  NANDN U15076 ( .A(n14707), .B(n42234), .Z(n14667) );
  AND U15077 ( .A(n14668), .B(n14667), .Z(n14716) );
  XNOR U15078 ( .A(n14717), .B(n14716), .Z(n14718) );
  XNOR U15079 ( .A(n14719), .B(n14718), .Z(n14723) );
  NANDN U15080 ( .A(n14670), .B(n14669), .Z(n14674) );
  NAND U15081 ( .A(n14672), .B(n14671), .Z(n14673) );
  AND U15082 ( .A(n14674), .B(n14673), .Z(n14722) );
  XOR U15083 ( .A(n14723), .B(n14722), .Z(n14724) );
  NANDN U15084 ( .A(n14676), .B(n14675), .Z(n14680) );
  NANDN U15085 ( .A(n14678), .B(n14677), .Z(n14679) );
  NAND U15086 ( .A(n14680), .B(n14679), .Z(n14725) );
  XOR U15087 ( .A(n14724), .B(n14725), .Z(n14692) );
  OR U15088 ( .A(n14682), .B(n14681), .Z(n14686) );
  NANDN U15089 ( .A(n14684), .B(n14683), .Z(n14685) );
  NAND U15090 ( .A(n14686), .B(n14685), .Z(n14693) );
  XNOR U15091 ( .A(n14692), .B(n14693), .Z(n14694) );
  XNOR U15092 ( .A(n14695), .B(n14694), .Z(n14728) );
  XNOR U15093 ( .A(n14728), .B(sreg[1372]), .Z(n14730) );
  NAND U15094 ( .A(n14687), .B(sreg[1371]), .Z(n14691) );
  OR U15095 ( .A(n14689), .B(n14688), .Z(n14690) );
  AND U15096 ( .A(n14691), .B(n14690), .Z(n14729) );
  XOR U15097 ( .A(n14730), .B(n14729), .Z(c[1372]) );
  NANDN U15098 ( .A(n14693), .B(n14692), .Z(n14697) );
  NAND U15099 ( .A(n14695), .B(n14694), .Z(n14696) );
  NAND U15100 ( .A(n14697), .B(n14696), .Z(n14736) );
  NAND U15101 ( .A(b[0]), .B(a[357]), .Z(n14698) );
  XNOR U15102 ( .A(b[1]), .B(n14698), .Z(n14700) );
  NAND U15103 ( .A(n66), .B(a[356]), .Z(n14699) );
  AND U15104 ( .A(n14700), .B(n14699), .Z(n14753) );
  XOR U15105 ( .A(a[353]), .B(n42197), .Z(n14742) );
  NANDN U15106 ( .A(n14742), .B(n42173), .Z(n14703) );
  NANDN U15107 ( .A(n14701), .B(n42172), .Z(n14702) );
  NAND U15108 ( .A(n14703), .B(n14702), .Z(n14751) );
  NAND U15109 ( .A(b[7]), .B(a[349]), .Z(n14752) );
  XNOR U15110 ( .A(n14751), .B(n14752), .Z(n14754) );
  XOR U15111 ( .A(n14753), .B(n14754), .Z(n14760) );
  NANDN U15112 ( .A(n14704), .B(n42093), .Z(n14706) );
  XOR U15113 ( .A(n42134), .B(a[355]), .Z(n14745) );
  NANDN U15114 ( .A(n14745), .B(n42095), .Z(n14705) );
  NAND U15115 ( .A(n14706), .B(n14705), .Z(n14758) );
  NANDN U15116 ( .A(n14707), .B(n42231), .Z(n14709) );
  XOR U15117 ( .A(n191), .B(a[351]), .Z(n14748) );
  NANDN U15118 ( .A(n14748), .B(n42234), .Z(n14708) );
  AND U15119 ( .A(n14709), .B(n14708), .Z(n14757) );
  XNOR U15120 ( .A(n14758), .B(n14757), .Z(n14759) );
  XNOR U15121 ( .A(n14760), .B(n14759), .Z(n14764) );
  NANDN U15122 ( .A(n14711), .B(n14710), .Z(n14715) );
  NAND U15123 ( .A(n14713), .B(n14712), .Z(n14714) );
  AND U15124 ( .A(n14715), .B(n14714), .Z(n14763) );
  XOR U15125 ( .A(n14764), .B(n14763), .Z(n14765) );
  NANDN U15126 ( .A(n14717), .B(n14716), .Z(n14721) );
  NANDN U15127 ( .A(n14719), .B(n14718), .Z(n14720) );
  NAND U15128 ( .A(n14721), .B(n14720), .Z(n14766) );
  XOR U15129 ( .A(n14765), .B(n14766), .Z(n14733) );
  OR U15130 ( .A(n14723), .B(n14722), .Z(n14727) );
  NANDN U15131 ( .A(n14725), .B(n14724), .Z(n14726) );
  NAND U15132 ( .A(n14727), .B(n14726), .Z(n14734) );
  XNOR U15133 ( .A(n14733), .B(n14734), .Z(n14735) );
  XNOR U15134 ( .A(n14736), .B(n14735), .Z(n14769) );
  XNOR U15135 ( .A(n14769), .B(sreg[1373]), .Z(n14771) );
  NAND U15136 ( .A(n14728), .B(sreg[1372]), .Z(n14732) );
  OR U15137 ( .A(n14730), .B(n14729), .Z(n14731) );
  AND U15138 ( .A(n14732), .B(n14731), .Z(n14770) );
  XOR U15139 ( .A(n14771), .B(n14770), .Z(c[1373]) );
  NANDN U15140 ( .A(n14734), .B(n14733), .Z(n14738) );
  NAND U15141 ( .A(n14736), .B(n14735), .Z(n14737) );
  NAND U15142 ( .A(n14738), .B(n14737), .Z(n14777) );
  NAND U15143 ( .A(b[0]), .B(a[358]), .Z(n14739) );
  XNOR U15144 ( .A(b[1]), .B(n14739), .Z(n14741) );
  NAND U15145 ( .A(n66), .B(a[357]), .Z(n14740) );
  AND U15146 ( .A(n14741), .B(n14740), .Z(n14794) );
  XOR U15147 ( .A(a[354]), .B(n42197), .Z(n14783) );
  NANDN U15148 ( .A(n14783), .B(n42173), .Z(n14744) );
  NANDN U15149 ( .A(n14742), .B(n42172), .Z(n14743) );
  NAND U15150 ( .A(n14744), .B(n14743), .Z(n14792) );
  NAND U15151 ( .A(b[7]), .B(a[350]), .Z(n14793) );
  XNOR U15152 ( .A(n14792), .B(n14793), .Z(n14795) );
  XOR U15153 ( .A(n14794), .B(n14795), .Z(n14801) );
  NANDN U15154 ( .A(n14745), .B(n42093), .Z(n14747) );
  XOR U15155 ( .A(n42134), .B(a[356]), .Z(n14786) );
  NANDN U15156 ( .A(n14786), .B(n42095), .Z(n14746) );
  NAND U15157 ( .A(n14747), .B(n14746), .Z(n14799) );
  NANDN U15158 ( .A(n14748), .B(n42231), .Z(n14750) );
  XOR U15159 ( .A(n191), .B(a[352]), .Z(n14789) );
  NANDN U15160 ( .A(n14789), .B(n42234), .Z(n14749) );
  AND U15161 ( .A(n14750), .B(n14749), .Z(n14798) );
  XNOR U15162 ( .A(n14799), .B(n14798), .Z(n14800) );
  XNOR U15163 ( .A(n14801), .B(n14800), .Z(n14805) );
  NANDN U15164 ( .A(n14752), .B(n14751), .Z(n14756) );
  NAND U15165 ( .A(n14754), .B(n14753), .Z(n14755) );
  AND U15166 ( .A(n14756), .B(n14755), .Z(n14804) );
  XOR U15167 ( .A(n14805), .B(n14804), .Z(n14806) );
  NANDN U15168 ( .A(n14758), .B(n14757), .Z(n14762) );
  NANDN U15169 ( .A(n14760), .B(n14759), .Z(n14761) );
  NAND U15170 ( .A(n14762), .B(n14761), .Z(n14807) );
  XOR U15171 ( .A(n14806), .B(n14807), .Z(n14774) );
  OR U15172 ( .A(n14764), .B(n14763), .Z(n14768) );
  NANDN U15173 ( .A(n14766), .B(n14765), .Z(n14767) );
  NAND U15174 ( .A(n14768), .B(n14767), .Z(n14775) );
  XNOR U15175 ( .A(n14774), .B(n14775), .Z(n14776) );
  XNOR U15176 ( .A(n14777), .B(n14776), .Z(n14810) );
  XNOR U15177 ( .A(n14810), .B(sreg[1374]), .Z(n14812) );
  NAND U15178 ( .A(n14769), .B(sreg[1373]), .Z(n14773) );
  OR U15179 ( .A(n14771), .B(n14770), .Z(n14772) );
  AND U15180 ( .A(n14773), .B(n14772), .Z(n14811) );
  XOR U15181 ( .A(n14812), .B(n14811), .Z(c[1374]) );
  NANDN U15182 ( .A(n14775), .B(n14774), .Z(n14779) );
  NAND U15183 ( .A(n14777), .B(n14776), .Z(n14778) );
  NAND U15184 ( .A(n14779), .B(n14778), .Z(n14818) );
  NAND U15185 ( .A(b[0]), .B(a[359]), .Z(n14780) );
  XNOR U15186 ( .A(b[1]), .B(n14780), .Z(n14782) );
  NAND U15187 ( .A(n66), .B(a[358]), .Z(n14781) );
  AND U15188 ( .A(n14782), .B(n14781), .Z(n14835) );
  XOR U15189 ( .A(a[355]), .B(n42197), .Z(n14824) );
  NANDN U15190 ( .A(n14824), .B(n42173), .Z(n14785) );
  NANDN U15191 ( .A(n14783), .B(n42172), .Z(n14784) );
  NAND U15192 ( .A(n14785), .B(n14784), .Z(n14833) );
  NAND U15193 ( .A(b[7]), .B(a[351]), .Z(n14834) );
  XNOR U15194 ( .A(n14833), .B(n14834), .Z(n14836) );
  XOR U15195 ( .A(n14835), .B(n14836), .Z(n14842) );
  NANDN U15196 ( .A(n14786), .B(n42093), .Z(n14788) );
  XOR U15197 ( .A(n42134), .B(a[357]), .Z(n14827) );
  NANDN U15198 ( .A(n14827), .B(n42095), .Z(n14787) );
  NAND U15199 ( .A(n14788), .B(n14787), .Z(n14840) );
  NANDN U15200 ( .A(n14789), .B(n42231), .Z(n14791) );
  XOR U15201 ( .A(n191), .B(a[353]), .Z(n14830) );
  NANDN U15202 ( .A(n14830), .B(n42234), .Z(n14790) );
  AND U15203 ( .A(n14791), .B(n14790), .Z(n14839) );
  XNOR U15204 ( .A(n14840), .B(n14839), .Z(n14841) );
  XNOR U15205 ( .A(n14842), .B(n14841), .Z(n14846) );
  NANDN U15206 ( .A(n14793), .B(n14792), .Z(n14797) );
  NAND U15207 ( .A(n14795), .B(n14794), .Z(n14796) );
  AND U15208 ( .A(n14797), .B(n14796), .Z(n14845) );
  XOR U15209 ( .A(n14846), .B(n14845), .Z(n14847) );
  NANDN U15210 ( .A(n14799), .B(n14798), .Z(n14803) );
  NANDN U15211 ( .A(n14801), .B(n14800), .Z(n14802) );
  NAND U15212 ( .A(n14803), .B(n14802), .Z(n14848) );
  XOR U15213 ( .A(n14847), .B(n14848), .Z(n14815) );
  OR U15214 ( .A(n14805), .B(n14804), .Z(n14809) );
  NANDN U15215 ( .A(n14807), .B(n14806), .Z(n14808) );
  NAND U15216 ( .A(n14809), .B(n14808), .Z(n14816) );
  XNOR U15217 ( .A(n14815), .B(n14816), .Z(n14817) );
  XNOR U15218 ( .A(n14818), .B(n14817), .Z(n14851) );
  XNOR U15219 ( .A(n14851), .B(sreg[1375]), .Z(n14853) );
  NAND U15220 ( .A(n14810), .B(sreg[1374]), .Z(n14814) );
  OR U15221 ( .A(n14812), .B(n14811), .Z(n14813) );
  AND U15222 ( .A(n14814), .B(n14813), .Z(n14852) );
  XOR U15223 ( .A(n14853), .B(n14852), .Z(c[1375]) );
  NANDN U15224 ( .A(n14816), .B(n14815), .Z(n14820) );
  NAND U15225 ( .A(n14818), .B(n14817), .Z(n14819) );
  NAND U15226 ( .A(n14820), .B(n14819), .Z(n14859) );
  NAND U15227 ( .A(b[0]), .B(a[360]), .Z(n14821) );
  XNOR U15228 ( .A(b[1]), .B(n14821), .Z(n14823) );
  NAND U15229 ( .A(n66), .B(a[359]), .Z(n14822) );
  AND U15230 ( .A(n14823), .B(n14822), .Z(n14876) );
  XOR U15231 ( .A(a[356]), .B(n42197), .Z(n14865) );
  NANDN U15232 ( .A(n14865), .B(n42173), .Z(n14826) );
  NANDN U15233 ( .A(n14824), .B(n42172), .Z(n14825) );
  NAND U15234 ( .A(n14826), .B(n14825), .Z(n14874) );
  NAND U15235 ( .A(b[7]), .B(a[352]), .Z(n14875) );
  XNOR U15236 ( .A(n14874), .B(n14875), .Z(n14877) );
  XOR U15237 ( .A(n14876), .B(n14877), .Z(n14883) );
  NANDN U15238 ( .A(n14827), .B(n42093), .Z(n14829) );
  XOR U15239 ( .A(n42134), .B(a[358]), .Z(n14868) );
  NANDN U15240 ( .A(n14868), .B(n42095), .Z(n14828) );
  NAND U15241 ( .A(n14829), .B(n14828), .Z(n14881) );
  NANDN U15242 ( .A(n14830), .B(n42231), .Z(n14832) );
  XOR U15243 ( .A(n191), .B(a[354]), .Z(n14871) );
  NANDN U15244 ( .A(n14871), .B(n42234), .Z(n14831) );
  AND U15245 ( .A(n14832), .B(n14831), .Z(n14880) );
  XNOR U15246 ( .A(n14881), .B(n14880), .Z(n14882) );
  XNOR U15247 ( .A(n14883), .B(n14882), .Z(n14887) );
  NANDN U15248 ( .A(n14834), .B(n14833), .Z(n14838) );
  NAND U15249 ( .A(n14836), .B(n14835), .Z(n14837) );
  AND U15250 ( .A(n14838), .B(n14837), .Z(n14886) );
  XOR U15251 ( .A(n14887), .B(n14886), .Z(n14888) );
  NANDN U15252 ( .A(n14840), .B(n14839), .Z(n14844) );
  NANDN U15253 ( .A(n14842), .B(n14841), .Z(n14843) );
  NAND U15254 ( .A(n14844), .B(n14843), .Z(n14889) );
  XOR U15255 ( .A(n14888), .B(n14889), .Z(n14856) );
  OR U15256 ( .A(n14846), .B(n14845), .Z(n14850) );
  NANDN U15257 ( .A(n14848), .B(n14847), .Z(n14849) );
  NAND U15258 ( .A(n14850), .B(n14849), .Z(n14857) );
  XNOR U15259 ( .A(n14856), .B(n14857), .Z(n14858) );
  XNOR U15260 ( .A(n14859), .B(n14858), .Z(n14892) );
  XNOR U15261 ( .A(n14892), .B(sreg[1376]), .Z(n14894) );
  NAND U15262 ( .A(n14851), .B(sreg[1375]), .Z(n14855) );
  OR U15263 ( .A(n14853), .B(n14852), .Z(n14854) );
  AND U15264 ( .A(n14855), .B(n14854), .Z(n14893) );
  XOR U15265 ( .A(n14894), .B(n14893), .Z(c[1376]) );
  NANDN U15266 ( .A(n14857), .B(n14856), .Z(n14861) );
  NAND U15267 ( .A(n14859), .B(n14858), .Z(n14860) );
  NAND U15268 ( .A(n14861), .B(n14860), .Z(n14900) );
  NAND U15269 ( .A(b[0]), .B(a[361]), .Z(n14862) );
  XNOR U15270 ( .A(b[1]), .B(n14862), .Z(n14864) );
  NAND U15271 ( .A(n66), .B(a[360]), .Z(n14863) );
  AND U15272 ( .A(n14864), .B(n14863), .Z(n14917) );
  XOR U15273 ( .A(a[357]), .B(n42197), .Z(n14906) );
  NANDN U15274 ( .A(n14906), .B(n42173), .Z(n14867) );
  NANDN U15275 ( .A(n14865), .B(n42172), .Z(n14866) );
  NAND U15276 ( .A(n14867), .B(n14866), .Z(n14915) );
  NAND U15277 ( .A(b[7]), .B(a[353]), .Z(n14916) );
  XNOR U15278 ( .A(n14915), .B(n14916), .Z(n14918) );
  XOR U15279 ( .A(n14917), .B(n14918), .Z(n14924) );
  NANDN U15280 ( .A(n14868), .B(n42093), .Z(n14870) );
  XOR U15281 ( .A(n42134), .B(a[359]), .Z(n14909) );
  NANDN U15282 ( .A(n14909), .B(n42095), .Z(n14869) );
  NAND U15283 ( .A(n14870), .B(n14869), .Z(n14922) );
  NANDN U15284 ( .A(n14871), .B(n42231), .Z(n14873) );
  XOR U15285 ( .A(n191), .B(a[355]), .Z(n14912) );
  NANDN U15286 ( .A(n14912), .B(n42234), .Z(n14872) );
  AND U15287 ( .A(n14873), .B(n14872), .Z(n14921) );
  XNOR U15288 ( .A(n14922), .B(n14921), .Z(n14923) );
  XNOR U15289 ( .A(n14924), .B(n14923), .Z(n14928) );
  NANDN U15290 ( .A(n14875), .B(n14874), .Z(n14879) );
  NAND U15291 ( .A(n14877), .B(n14876), .Z(n14878) );
  AND U15292 ( .A(n14879), .B(n14878), .Z(n14927) );
  XOR U15293 ( .A(n14928), .B(n14927), .Z(n14929) );
  NANDN U15294 ( .A(n14881), .B(n14880), .Z(n14885) );
  NANDN U15295 ( .A(n14883), .B(n14882), .Z(n14884) );
  NAND U15296 ( .A(n14885), .B(n14884), .Z(n14930) );
  XOR U15297 ( .A(n14929), .B(n14930), .Z(n14897) );
  OR U15298 ( .A(n14887), .B(n14886), .Z(n14891) );
  NANDN U15299 ( .A(n14889), .B(n14888), .Z(n14890) );
  NAND U15300 ( .A(n14891), .B(n14890), .Z(n14898) );
  XNOR U15301 ( .A(n14897), .B(n14898), .Z(n14899) );
  XNOR U15302 ( .A(n14900), .B(n14899), .Z(n14933) );
  XNOR U15303 ( .A(n14933), .B(sreg[1377]), .Z(n14935) );
  NAND U15304 ( .A(n14892), .B(sreg[1376]), .Z(n14896) );
  OR U15305 ( .A(n14894), .B(n14893), .Z(n14895) );
  AND U15306 ( .A(n14896), .B(n14895), .Z(n14934) );
  XOR U15307 ( .A(n14935), .B(n14934), .Z(c[1377]) );
  NANDN U15308 ( .A(n14898), .B(n14897), .Z(n14902) );
  NAND U15309 ( .A(n14900), .B(n14899), .Z(n14901) );
  NAND U15310 ( .A(n14902), .B(n14901), .Z(n14941) );
  NAND U15311 ( .A(b[0]), .B(a[362]), .Z(n14903) );
  XNOR U15312 ( .A(b[1]), .B(n14903), .Z(n14905) );
  NAND U15313 ( .A(n66), .B(a[361]), .Z(n14904) );
  AND U15314 ( .A(n14905), .B(n14904), .Z(n14958) );
  XOR U15315 ( .A(a[358]), .B(n42197), .Z(n14947) );
  NANDN U15316 ( .A(n14947), .B(n42173), .Z(n14908) );
  NANDN U15317 ( .A(n14906), .B(n42172), .Z(n14907) );
  NAND U15318 ( .A(n14908), .B(n14907), .Z(n14956) );
  NAND U15319 ( .A(b[7]), .B(a[354]), .Z(n14957) );
  XNOR U15320 ( .A(n14956), .B(n14957), .Z(n14959) );
  XOR U15321 ( .A(n14958), .B(n14959), .Z(n14965) );
  NANDN U15322 ( .A(n14909), .B(n42093), .Z(n14911) );
  XOR U15323 ( .A(n42134), .B(a[360]), .Z(n14950) );
  NANDN U15324 ( .A(n14950), .B(n42095), .Z(n14910) );
  NAND U15325 ( .A(n14911), .B(n14910), .Z(n14963) );
  NANDN U15326 ( .A(n14912), .B(n42231), .Z(n14914) );
  XOR U15327 ( .A(n191), .B(a[356]), .Z(n14953) );
  NANDN U15328 ( .A(n14953), .B(n42234), .Z(n14913) );
  AND U15329 ( .A(n14914), .B(n14913), .Z(n14962) );
  XNOR U15330 ( .A(n14963), .B(n14962), .Z(n14964) );
  XNOR U15331 ( .A(n14965), .B(n14964), .Z(n14969) );
  NANDN U15332 ( .A(n14916), .B(n14915), .Z(n14920) );
  NAND U15333 ( .A(n14918), .B(n14917), .Z(n14919) );
  AND U15334 ( .A(n14920), .B(n14919), .Z(n14968) );
  XOR U15335 ( .A(n14969), .B(n14968), .Z(n14970) );
  NANDN U15336 ( .A(n14922), .B(n14921), .Z(n14926) );
  NANDN U15337 ( .A(n14924), .B(n14923), .Z(n14925) );
  NAND U15338 ( .A(n14926), .B(n14925), .Z(n14971) );
  XOR U15339 ( .A(n14970), .B(n14971), .Z(n14938) );
  OR U15340 ( .A(n14928), .B(n14927), .Z(n14932) );
  NANDN U15341 ( .A(n14930), .B(n14929), .Z(n14931) );
  NAND U15342 ( .A(n14932), .B(n14931), .Z(n14939) );
  XNOR U15343 ( .A(n14938), .B(n14939), .Z(n14940) );
  XNOR U15344 ( .A(n14941), .B(n14940), .Z(n14974) );
  XNOR U15345 ( .A(n14974), .B(sreg[1378]), .Z(n14976) );
  NAND U15346 ( .A(n14933), .B(sreg[1377]), .Z(n14937) );
  OR U15347 ( .A(n14935), .B(n14934), .Z(n14936) );
  AND U15348 ( .A(n14937), .B(n14936), .Z(n14975) );
  XOR U15349 ( .A(n14976), .B(n14975), .Z(c[1378]) );
  NANDN U15350 ( .A(n14939), .B(n14938), .Z(n14943) );
  NAND U15351 ( .A(n14941), .B(n14940), .Z(n14942) );
  NAND U15352 ( .A(n14943), .B(n14942), .Z(n14982) );
  NAND U15353 ( .A(b[0]), .B(a[363]), .Z(n14944) );
  XNOR U15354 ( .A(b[1]), .B(n14944), .Z(n14946) );
  NAND U15355 ( .A(n66), .B(a[362]), .Z(n14945) );
  AND U15356 ( .A(n14946), .B(n14945), .Z(n14999) );
  XOR U15357 ( .A(a[359]), .B(n42197), .Z(n14988) );
  NANDN U15358 ( .A(n14988), .B(n42173), .Z(n14949) );
  NANDN U15359 ( .A(n14947), .B(n42172), .Z(n14948) );
  NAND U15360 ( .A(n14949), .B(n14948), .Z(n14997) );
  NAND U15361 ( .A(b[7]), .B(a[355]), .Z(n14998) );
  XNOR U15362 ( .A(n14997), .B(n14998), .Z(n15000) );
  XOR U15363 ( .A(n14999), .B(n15000), .Z(n15006) );
  NANDN U15364 ( .A(n14950), .B(n42093), .Z(n14952) );
  XOR U15365 ( .A(n42134), .B(a[361]), .Z(n14991) );
  NANDN U15366 ( .A(n14991), .B(n42095), .Z(n14951) );
  NAND U15367 ( .A(n14952), .B(n14951), .Z(n15004) );
  NANDN U15368 ( .A(n14953), .B(n42231), .Z(n14955) );
  XOR U15369 ( .A(n191), .B(a[357]), .Z(n14994) );
  NANDN U15370 ( .A(n14994), .B(n42234), .Z(n14954) );
  AND U15371 ( .A(n14955), .B(n14954), .Z(n15003) );
  XNOR U15372 ( .A(n15004), .B(n15003), .Z(n15005) );
  XNOR U15373 ( .A(n15006), .B(n15005), .Z(n15010) );
  NANDN U15374 ( .A(n14957), .B(n14956), .Z(n14961) );
  NAND U15375 ( .A(n14959), .B(n14958), .Z(n14960) );
  AND U15376 ( .A(n14961), .B(n14960), .Z(n15009) );
  XOR U15377 ( .A(n15010), .B(n15009), .Z(n15011) );
  NANDN U15378 ( .A(n14963), .B(n14962), .Z(n14967) );
  NANDN U15379 ( .A(n14965), .B(n14964), .Z(n14966) );
  NAND U15380 ( .A(n14967), .B(n14966), .Z(n15012) );
  XOR U15381 ( .A(n15011), .B(n15012), .Z(n14979) );
  OR U15382 ( .A(n14969), .B(n14968), .Z(n14973) );
  NANDN U15383 ( .A(n14971), .B(n14970), .Z(n14972) );
  NAND U15384 ( .A(n14973), .B(n14972), .Z(n14980) );
  XNOR U15385 ( .A(n14979), .B(n14980), .Z(n14981) );
  XNOR U15386 ( .A(n14982), .B(n14981), .Z(n15015) );
  XNOR U15387 ( .A(n15015), .B(sreg[1379]), .Z(n15017) );
  NAND U15388 ( .A(n14974), .B(sreg[1378]), .Z(n14978) );
  OR U15389 ( .A(n14976), .B(n14975), .Z(n14977) );
  AND U15390 ( .A(n14978), .B(n14977), .Z(n15016) );
  XOR U15391 ( .A(n15017), .B(n15016), .Z(c[1379]) );
  NANDN U15392 ( .A(n14980), .B(n14979), .Z(n14984) );
  NAND U15393 ( .A(n14982), .B(n14981), .Z(n14983) );
  NAND U15394 ( .A(n14984), .B(n14983), .Z(n15023) );
  NAND U15395 ( .A(b[0]), .B(a[364]), .Z(n14985) );
  XNOR U15396 ( .A(b[1]), .B(n14985), .Z(n14987) );
  NAND U15397 ( .A(n67), .B(a[363]), .Z(n14986) );
  AND U15398 ( .A(n14987), .B(n14986), .Z(n15040) );
  XOR U15399 ( .A(a[360]), .B(n42197), .Z(n15029) );
  NANDN U15400 ( .A(n15029), .B(n42173), .Z(n14990) );
  NANDN U15401 ( .A(n14988), .B(n42172), .Z(n14989) );
  NAND U15402 ( .A(n14990), .B(n14989), .Z(n15038) );
  NAND U15403 ( .A(b[7]), .B(a[356]), .Z(n15039) );
  XNOR U15404 ( .A(n15038), .B(n15039), .Z(n15041) );
  XOR U15405 ( .A(n15040), .B(n15041), .Z(n15047) );
  NANDN U15406 ( .A(n14991), .B(n42093), .Z(n14993) );
  XOR U15407 ( .A(n42134), .B(a[362]), .Z(n15032) );
  NANDN U15408 ( .A(n15032), .B(n42095), .Z(n14992) );
  NAND U15409 ( .A(n14993), .B(n14992), .Z(n15045) );
  NANDN U15410 ( .A(n14994), .B(n42231), .Z(n14996) );
  XOR U15411 ( .A(n191), .B(a[358]), .Z(n15035) );
  NANDN U15412 ( .A(n15035), .B(n42234), .Z(n14995) );
  AND U15413 ( .A(n14996), .B(n14995), .Z(n15044) );
  XNOR U15414 ( .A(n15045), .B(n15044), .Z(n15046) );
  XNOR U15415 ( .A(n15047), .B(n15046), .Z(n15051) );
  NANDN U15416 ( .A(n14998), .B(n14997), .Z(n15002) );
  NAND U15417 ( .A(n15000), .B(n14999), .Z(n15001) );
  AND U15418 ( .A(n15002), .B(n15001), .Z(n15050) );
  XOR U15419 ( .A(n15051), .B(n15050), .Z(n15052) );
  NANDN U15420 ( .A(n15004), .B(n15003), .Z(n15008) );
  NANDN U15421 ( .A(n15006), .B(n15005), .Z(n15007) );
  NAND U15422 ( .A(n15008), .B(n15007), .Z(n15053) );
  XOR U15423 ( .A(n15052), .B(n15053), .Z(n15020) );
  OR U15424 ( .A(n15010), .B(n15009), .Z(n15014) );
  NANDN U15425 ( .A(n15012), .B(n15011), .Z(n15013) );
  NAND U15426 ( .A(n15014), .B(n15013), .Z(n15021) );
  XNOR U15427 ( .A(n15020), .B(n15021), .Z(n15022) );
  XNOR U15428 ( .A(n15023), .B(n15022), .Z(n15056) );
  XNOR U15429 ( .A(n15056), .B(sreg[1380]), .Z(n15058) );
  NAND U15430 ( .A(n15015), .B(sreg[1379]), .Z(n15019) );
  OR U15431 ( .A(n15017), .B(n15016), .Z(n15018) );
  AND U15432 ( .A(n15019), .B(n15018), .Z(n15057) );
  XOR U15433 ( .A(n15058), .B(n15057), .Z(c[1380]) );
  NANDN U15434 ( .A(n15021), .B(n15020), .Z(n15025) );
  NAND U15435 ( .A(n15023), .B(n15022), .Z(n15024) );
  NAND U15436 ( .A(n15025), .B(n15024), .Z(n15064) );
  NAND U15437 ( .A(b[0]), .B(a[365]), .Z(n15026) );
  XNOR U15438 ( .A(b[1]), .B(n15026), .Z(n15028) );
  NAND U15439 ( .A(n67), .B(a[364]), .Z(n15027) );
  AND U15440 ( .A(n15028), .B(n15027), .Z(n15081) );
  XOR U15441 ( .A(a[361]), .B(n42197), .Z(n15070) );
  NANDN U15442 ( .A(n15070), .B(n42173), .Z(n15031) );
  NANDN U15443 ( .A(n15029), .B(n42172), .Z(n15030) );
  NAND U15444 ( .A(n15031), .B(n15030), .Z(n15079) );
  NAND U15445 ( .A(b[7]), .B(a[357]), .Z(n15080) );
  XNOR U15446 ( .A(n15079), .B(n15080), .Z(n15082) );
  XOR U15447 ( .A(n15081), .B(n15082), .Z(n15088) );
  NANDN U15448 ( .A(n15032), .B(n42093), .Z(n15034) );
  XOR U15449 ( .A(n42134), .B(a[363]), .Z(n15073) );
  NANDN U15450 ( .A(n15073), .B(n42095), .Z(n15033) );
  NAND U15451 ( .A(n15034), .B(n15033), .Z(n15086) );
  NANDN U15452 ( .A(n15035), .B(n42231), .Z(n15037) );
  XOR U15453 ( .A(n192), .B(a[359]), .Z(n15076) );
  NANDN U15454 ( .A(n15076), .B(n42234), .Z(n15036) );
  AND U15455 ( .A(n15037), .B(n15036), .Z(n15085) );
  XNOR U15456 ( .A(n15086), .B(n15085), .Z(n15087) );
  XNOR U15457 ( .A(n15088), .B(n15087), .Z(n15092) );
  NANDN U15458 ( .A(n15039), .B(n15038), .Z(n15043) );
  NAND U15459 ( .A(n15041), .B(n15040), .Z(n15042) );
  AND U15460 ( .A(n15043), .B(n15042), .Z(n15091) );
  XOR U15461 ( .A(n15092), .B(n15091), .Z(n15093) );
  NANDN U15462 ( .A(n15045), .B(n15044), .Z(n15049) );
  NANDN U15463 ( .A(n15047), .B(n15046), .Z(n15048) );
  NAND U15464 ( .A(n15049), .B(n15048), .Z(n15094) );
  XOR U15465 ( .A(n15093), .B(n15094), .Z(n15061) );
  OR U15466 ( .A(n15051), .B(n15050), .Z(n15055) );
  NANDN U15467 ( .A(n15053), .B(n15052), .Z(n15054) );
  NAND U15468 ( .A(n15055), .B(n15054), .Z(n15062) );
  XNOR U15469 ( .A(n15061), .B(n15062), .Z(n15063) );
  XNOR U15470 ( .A(n15064), .B(n15063), .Z(n15097) );
  XNOR U15471 ( .A(n15097), .B(sreg[1381]), .Z(n15099) );
  NAND U15472 ( .A(n15056), .B(sreg[1380]), .Z(n15060) );
  OR U15473 ( .A(n15058), .B(n15057), .Z(n15059) );
  AND U15474 ( .A(n15060), .B(n15059), .Z(n15098) );
  XOR U15475 ( .A(n15099), .B(n15098), .Z(c[1381]) );
  NANDN U15476 ( .A(n15062), .B(n15061), .Z(n15066) );
  NAND U15477 ( .A(n15064), .B(n15063), .Z(n15065) );
  NAND U15478 ( .A(n15066), .B(n15065), .Z(n15105) );
  NAND U15479 ( .A(b[0]), .B(a[366]), .Z(n15067) );
  XNOR U15480 ( .A(b[1]), .B(n15067), .Z(n15069) );
  NAND U15481 ( .A(n67), .B(a[365]), .Z(n15068) );
  AND U15482 ( .A(n15069), .B(n15068), .Z(n15122) );
  XOR U15483 ( .A(a[362]), .B(n42197), .Z(n15111) );
  NANDN U15484 ( .A(n15111), .B(n42173), .Z(n15072) );
  NANDN U15485 ( .A(n15070), .B(n42172), .Z(n15071) );
  NAND U15486 ( .A(n15072), .B(n15071), .Z(n15120) );
  NAND U15487 ( .A(b[7]), .B(a[358]), .Z(n15121) );
  XNOR U15488 ( .A(n15120), .B(n15121), .Z(n15123) );
  XOR U15489 ( .A(n15122), .B(n15123), .Z(n15129) );
  NANDN U15490 ( .A(n15073), .B(n42093), .Z(n15075) );
  XOR U15491 ( .A(n42134), .B(a[364]), .Z(n15114) );
  NANDN U15492 ( .A(n15114), .B(n42095), .Z(n15074) );
  NAND U15493 ( .A(n15075), .B(n15074), .Z(n15127) );
  NANDN U15494 ( .A(n15076), .B(n42231), .Z(n15078) );
  XOR U15495 ( .A(n192), .B(a[360]), .Z(n15117) );
  NANDN U15496 ( .A(n15117), .B(n42234), .Z(n15077) );
  AND U15497 ( .A(n15078), .B(n15077), .Z(n15126) );
  XNOR U15498 ( .A(n15127), .B(n15126), .Z(n15128) );
  XNOR U15499 ( .A(n15129), .B(n15128), .Z(n15133) );
  NANDN U15500 ( .A(n15080), .B(n15079), .Z(n15084) );
  NAND U15501 ( .A(n15082), .B(n15081), .Z(n15083) );
  AND U15502 ( .A(n15084), .B(n15083), .Z(n15132) );
  XOR U15503 ( .A(n15133), .B(n15132), .Z(n15134) );
  NANDN U15504 ( .A(n15086), .B(n15085), .Z(n15090) );
  NANDN U15505 ( .A(n15088), .B(n15087), .Z(n15089) );
  NAND U15506 ( .A(n15090), .B(n15089), .Z(n15135) );
  XOR U15507 ( .A(n15134), .B(n15135), .Z(n15102) );
  OR U15508 ( .A(n15092), .B(n15091), .Z(n15096) );
  NANDN U15509 ( .A(n15094), .B(n15093), .Z(n15095) );
  NAND U15510 ( .A(n15096), .B(n15095), .Z(n15103) );
  XNOR U15511 ( .A(n15102), .B(n15103), .Z(n15104) );
  XNOR U15512 ( .A(n15105), .B(n15104), .Z(n15138) );
  XNOR U15513 ( .A(n15138), .B(sreg[1382]), .Z(n15140) );
  NAND U15514 ( .A(n15097), .B(sreg[1381]), .Z(n15101) );
  OR U15515 ( .A(n15099), .B(n15098), .Z(n15100) );
  AND U15516 ( .A(n15101), .B(n15100), .Z(n15139) );
  XOR U15517 ( .A(n15140), .B(n15139), .Z(c[1382]) );
  NANDN U15518 ( .A(n15103), .B(n15102), .Z(n15107) );
  NAND U15519 ( .A(n15105), .B(n15104), .Z(n15106) );
  NAND U15520 ( .A(n15107), .B(n15106), .Z(n15146) );
  NAND U15521 ( .A(b[0]), .B(a[367]), .Z(n15108) );
  XNOR U15522 ( .A(b[1]), .B(n15108), .Z(n15110) );
  NAND U15523 ( .A(n67), .B(a[366]), .Z(n15109) );
  AND U15524 ( .A(n15110), .B(n15109), .Z(n15163) );
  XOR U15525 ( .A(a[363]), .B(n42197), .Z(n15152) );
  NANDN U15526 ( .A(n15152), .B(n42173), .Z(n15113) );
  NANDN U15527 ( .A(n15111), .B(n42172), .Z(n15112) );
  NAND U15528 ( .A(n15113), .B(n15112), .Z(n15161) );
  NAND U15529 ( .A(b[7]), .B(a[359]), .Z(n15162) );
  XNOR U15530 ( .A(n15161), .B(n15162), .Z(n15164) );
  XOR U15531 ( .A(n15163), .B(n15164), .Z(n15170) );
  NANDN U15532 ( .A(n15114), .B(n42093), .Z(n15116) );
  XOR U15533 ( .A(n42134), .B(a[365]), .Z(n15155) );
  NANDN U15534 ( .A(n15155), .B(n42095), .Z(n15115) );
  NAND U15535 ( .A(n15116), .B(n15115), .Z(n15168) );
  NANDN U15536 ( .A(n15117), .B(n42231), .Z(n15119) );
  XOR U15537 ( .A(n192), .B(a[361]), .Z(n15158) );
  NANDN U15538 ( .A(n15158), .B(n42234), .Z(n15118) );
  AND U15539 ( .A(n15119), .B(n15118), .Z(n15167) );
  XNOR U15540 ( .A(n15168), .B(n15167), .Z(n15169) );
  XNOR U15541 ( .A(n15170), .B(n15169), .Z(n15174) );
  NANDN U15542 ( .A(n15121), .B(n15120), .Z(n15125) );
  NAND U15543 ( .A(n15123), .B(n15122), .Z(n15124) );
  AND U15544 ( .A(n15125), .B(n15124), .Z(n15173) );
  XOR U15545 ( .A(n15174), .B(n15173), .Z(n15175) );
  NANDN U15546 ( .A(n15127), .B(n15126), .Z(n15131) );
  NANDN U15547 ( .A(n15129), .B(n15128), .Z(n15130) );
  NAND U15548 ( .A(n15131), .B(n15130), .Z(n15176) );
  XOR U15549 ( .A(n15175), .B(n15176), .Z(n15143) );
  OR U15550 ( .A(n15133), .B(n15132), .Z(n15137) );
  NANDN U15551 ( .A(n15135), .B(n15134), .Z(n15136) );
  NAND U15552 ( .A(n15137), .B(n15136), .Z(n15144) );
  XNOR U15553 ( .A(n15143), .B(n15144), .Z(n15145) );
  XNOR U15554 ( .A(n15146), .B(n15145), .Z(n15179) );
  XNOR U15555 ( .A(n15179), .B(sreg[1383]), .Z(n15181) );
  NAND U15556 ( .A(n15138), .B(sreg[1382]), .Z(n15142) );
  OR U15557 ( .A(n15140), .B(n15139), .Z(n15141) );
  AND U15558 ( .A(n15142), .B(n15141), .Z(n15180) );
  XOR U15559 ( .A(n15181), .B(n15180), .Z(c[1383]) );
  NANDN U15560 ( .A(n15144), .B(n15143), .Z(n15148) );
  NAND U15561 ( .A(n15146), .B(n15145), .Z(n15147) );
  NAND U15562 ( .A(n15148), .B(n15147), .Z(n15187) );
  NAND U15563 ( .A(b[0]), .B(a[368]), .Z(n15149) );
  XNOR U15564 ( .A(b[1]), .B(n15149), .Z(n15151) );
  NAND U15565 ( .A(n67), .B(a[367]), .Z(n15150) );
  AND U15566 ( .A(n15151), .B(n15150), .Z(n15204) );
  XOR U15567 ( .A(a[364]), .B(n42197), .Z(n15193) );
  NANDN U15568 ( .A(n15193), .B(n42173), .Z(n15154) );
  NANDN U15569 ( .A(n15152), .B(n42172), .Z(n15153) );
  NAND U15570 ( .A(n15154), .B(n15153), .Z(n15202) );
  NAND U15571 ( .A(b[7]), .B(a[360]), .Z(n15203) );
  XNOR U15572 ( .A(n15202), .B(n15203), .Z(n15205) );
  XOR U15573 ( .A(n15204), .B(n15205), .Z(n15211) );
  NANDN U15574 ( .A(n15155), .B(n42093), .Z(n15157) );
  XOR U15575 ( .A(n42134), .B(a[366]), .Z(n15196) );
  NANDN U15576 ( .A(n15196), .B(n42095), .Z(n15156) );
  NAND U15577 ( .A(n15157), .B(n15156), .Z(n15209) );
  NANDN U15578 ( .A(n15158), .B(n42231), .Z(n15160) );
  XOR U15579 ( .A(n192), .B(a[362]), .Z(n15199) );
  NANDN U15580 ( .A(n15199), .B(n42234), .Z(n15159) );
  AND U15581 ( .A(n15160), .B(n15159), .Z(n15208) );
  XNOR U15582 ( .A(n15209), .B(n15208), .Z(n15210) );
  XNOR U15583 ( .A(n15211), .B(n15210), .Z(n15215) );
  NANDN U15584 ( .A(n15162), .B(n15161), .Z(n15166) );
  NAND U15585 ( .A(n15164), .B(n15163), .Z(n15165) );
  AND U15586 ( .A(n15166), .B(n15165), .Z(n15214) );
  XOR U15587 ( .A(n15215), .B(n15214), .Z(n15216) );
  NANDN U15588 ( .A(n15168), .B(n15167), .Z(n15172) );
  NANDN U15589 ( .A(n15170), .B(n15169), .Z(n15171) );
  NAND U15590 ( .A(n15172), .B(n15171), .Z(n15217) );
  XOR U15591 ( .A(n15216), .B(n15217), .Z(n15184) );
  OR U15592 ( .A(n15174), .B(n15173), .Z(n15178) );
  NANDN U15593 ( .A(n15176), .B(n15175), .Z(n15177) );
  NAND U15594 ( .A(n15178), .B(n15177), .Z(n15185) );
  XNOR U15595 ( .A(n15184), .B(n15185), .Z(n15186) );
  XNOR U15596 ( .A(n15187), .B(n15186), .Z(n15220) );
  XNOR U15597 ( .A(n15220), .B(sreg[1384]), .Z(n15222) );
  NAND U15598 ( .A(n15179), .B(sreg[1383]), .Z(n15183) );
  OR U15599 ( .A(n15181), .B(n15180), .Z(n15182) );
  AND U15600 ( .A(n15183), .B(n15182), .Z(n15221) );
  XOR U15601 ( .A(n15222), .B(n15221), .Z(c[1384]) );
  NANDN U15602 ( .A(n15185), .B(n15184), .Z(n15189) );
  NAND U15603 ( .A(n15187), .B(n15186), .Z(n15188) );
  NAND U15604 ( .A(n15189), .B(n15188), .Z(n15228) );
  NAND U15605 ( .A(b[0]), .B(a[369]), .Z(n15190) );
  XNOR U15606 ( .A(b[1]), .B(n15190), .Z(n15192) );
  NAND U15607 ( .A(n67), .B(a[368]), .Z(n15191) );
  AND U15608 ( .A(n15192), .B(n15191), .Z(n15245) );
  XOR U15609 ( .A(a[365]), .B(n42197), .Z(n15234) );
  NANDN U15610 ( .A(n15234), .B(n42173), .Z(n15195) );
  NANDN U15611 ( .A(n15193), .B(n42172), .Z(n15194) );
  NAND U15612 ( .A(n15195), .B(n15194), .Z(n15243) );
  NAND U15613 ( .A(b[7]), .B(a[361]), .Z(n15244) );
  XNOR U15614 ( .A(n15243), .B(n15244), .Z(n15246) );
  XOR U15615 ( .A(n15245), .B(n15246), .Z(n15252) );
  NANDN U15616 ( .A(n15196), .B(n42093), .Z(n15198) );
  XOR U15617 ( .A(n42134), .B(a[367]), .Z(n15237) );
  NANDN U15618 ( .A(n15237), .B(n42095), .Z(n15197) );
  NAND U15619 ( .A(n15198), .B(n15197), .Z(n15250) );
  NANDN U15620 ( .A(n15199), .B(n42231), .Z(n15201) );
  XOR U15621 ( .A(n192), .B(a[363]), .Z(n15240) );
  NANDN U15622 ( .A(n15240), .B(n42234), .Z(n15200) );
  AND U15623 ( .A(n15201), .B(n15200), .Z(n15249) );
  XNOR U15624 ( .A(n15250), .B(n15249), .Z(n15251) );
  XNOR U15625 ( .A(n15252), .B(n15251), .Z(n15256) );
  NANDN U15626 ( .A(n15203), .B(n15202), .Z(n15207) );
  NAND U15627 ( .A(n15205), .B(n15204), .Z(n15206) );
  AND U15628 ( .A(n15207), .B(n15206), .Z(n15255) );
  XOR U15629 ( .A(n15256), .B(n15255), .Z(n15257) );
  NANDN U15630 ( .A(n15209), .B(n15208), .Z(n15213) );
  NANDN U15631 ( .A(n15211), .B(n15210), .Z(n15212) );
  NAND U15632 ( .A(n15213), .B(n15212), .Z(n15258) );
  XOR U15633 ( .A(n15257), .B(n15258), .Z(n15225) );
  OR U15634 ( .A(n15215), .B(n15214), .Z(n15219) );
  NANDN U15635 ( .A(n15217), .B(n15216), .Z(n15218) );
  NAND U15636 ( .A(n15219), .B(n15218), .Z(n15226) );
  XNOR U15637 ( .A(n15225), .B(n15226), .Z(n15227) );
  XNOR U15638 ( .A(n15228), .B(n15227), .Z(n15261) );
  XNOR U15639 ( .A(n15261), .B(sreg[1385]), .Z(n15263) );
  NAND U15640 ( .A(n15220), .B(sreg[1384]), .Z(n15224) );
  OR U15641 ( .A(n15222), .B(n15221), .Z(n15223) );
  AND U15642 ( .A(n15224), .B(n15223), .Z(n15262) );
  XOR U15643 ( .A(n15263), .B(n15262), .Z(c[1385]) );
  NANDN U15644 ( .A(n15226), .B(n15225), .Z(n15230) );
  NAND U15645 ( .A(n15228), .B(n15227), .Z(n15229) );
  NAND U15646 ( .A(n15230), .B(n15229), .Z(n15269) );
  NAND U15647 ( .A(b[0]), .B(a[370]), .Z(n15231) );
  XNOR U15648 ( .A(b[1]), .B(n15231), .Z(n15233) );
  NAND U15649 ( .A(n67), .B(a[369]), .Z(n15232) );
  AND U15650 ( .A(n15233), .B(n15232), .Z(n15286) );
  XOR U15651 ( .A(a[366]), .B(n42197), .Z(n15275) );
  NANDN U15652 ( .A(n15275), .B(n42173), .Z(n15236) );
  NANDN U15653 ( .A(n15234), .B(n42172), .Z(n15235) );
  NAND U15654 ( .A(n15236), .B(n15235), .Z(n15284) );
  NAND U15655 ( .A(b[7]), .B(a[362]), .Z(n15285) );
  XNOR U15656 ( .A(n15284), .B(n15285), .Z(n15287) );
  XOR U15657 ( .A(n15286), .B(n15287), .Z(n15293) );
  NANDN U15658 ( .A(n15237), .B(n42093), .Z(n15239) );
  XOR U15659 ( .A(n42134), .B(a[368]), .Z(n15278) );
  NANDN U15660 ( .A(n15278), .B(n42095), .Z(n15238) );
  NAND U15661 ( .A(n15239), .B(n15238), .Z(n15291) );
  NANDN U15662 ( .A(n15240), .B(n42231), .Z(n15242) );
  XOR U15663 ( .A(n192), .B(a[364]), .Z(n15281) );
  NANDN U15664 ( .A(n15281), .B(n42234), .Z(n15241) );
  AND U15665 ( .A(n15242), .B(n15241), .Z(n15290) );
  XNOR U15666 ( .A(n15291), .B(n15290), .Z(n15292) );
  XNOR U15667 ( .A(n15293), .B(n15292), .Z(n15297) );
  NANDN U15668 ( .A(n15244), .B(n15243), .Z(n15248) );
  NAND U15669 ( .A(n15246), .B(n15245), .Z(n15247) );
  AND U15670 ( .A(n15248), .B(n15247), .Z(n15296) );
  XOR U15671 ( .A(n15297), .B(n15296), .Z(n15298) );
  NANDN U15672 ( .A(n15250), .B(n15249), .Z(n15254) );
  NANDN U15673 ( .A(n15252), .B(n15251), .Z(n15253) );
  NAND U15674 ( .A(n15254), .B(n15253), .Z(n15299) );
  XOR U15675 ( .A(n15298), .B(n15299), .Z(n15266) );
  OR U15676 ( .A(n15256), .B(n15255), .Z(n15260) );
  NANDN U15677 ( .A(n15258), .B(n15257), .Z(n15259) );
  NAND U15678 ( .A(n15260), .B(n15259), .Z(n15267) );
  XNOR U15679 ( .A(n15266), .B(n15267), .Z(n15268) );
  XNOR U15680 ( .A(n15269), .B(n15268), .Z(n15302) );
  XNOR U15681 ( .A(n15302), .B(sreg[1386]), .Z(n15304) );
  NAND U15682 ( .A(n15261), .B(sreg[1385]), .Z(n15265) );
  OR U15683 ( .A(n15263), .B(n15262), .Z(n15264) );
  AND U15684 ( .A(n15265), .B(n15264), .Z(n15303) );
  XOR U15685 ( .A(n15304), .B(n15303), .Z(c[1386]) );
  NANDN U15686 ( .A(n15267), .B(n15266), .Z(n15271) );
  NAND U15687 ( .A(n15269), .B(n15268), .Z(n15270) );
  NAND U15688 ( .A(n15271), .B(n15270), .Z(n15310) );
  NAND U15689 ( .A(b[0]), .B(a[371]), .Z(n15272) );
  XNOR U15690 ( .A(b[1]), .B(n15272), .Z(n15274) );
  NAND U15691 ( .A(n68), .B(a[370]), .Z(n15273) );
  AND U15692 ( .A(n15274), .B(n15273), .Z(n15327) );
  XOR U15693 ( .A(a[367]), .B(n42197), .Z(n15316) );
  NANDN U15694 ( .A(n15316), .B(n42173), .Z(n15277) );
  NANDN U15695 ( .A(n15275), .B(n42172), .Z(n15276) );
  NAND U15696 ( .A(n15277), .B(n15276), .Z(n15325) );
  NAND U15697 ( .A(b[7]), .B(a[363]), .Z(n15326) );
  XNOR U15698 ( .A(n15325), .B(n15326), .Z(n15328) );
  XOR U15699 ( .A(n15327), .B(n15328), .Z(n15334) );
  NANDN U15700 ( .A(n15278), .B(n42093), .Z(n15280) );
  XOR U15701 ( .A(n42134), .B(a[369]), .Z(n15319) );
  NANDN U15702 ( .A(n15319), .B(n42095), .Z(n15279) );
  NAND U15703 ( .A(n15280), .B(n15279), .Z(n15332) );
  NANDN U15704 ( .A(n15281), .B(n42231), .Z(n15283) );
  XOR U15705 ( .A(n192), .B(a[365]), .Z(n15322) );
  NANDN U15706 ( .A(n15322), .B(n42234), .Z(n15282) );
  AND U15707 ( .A(n15283), .B(n15282), .Z(n15331) );
  XNOR U15708 ( .A(n15332), .B(n15331), .Z(n15333) );
  XNOR U15709 ( .A(n15334), .B(n15333), .Z(n15338) );
  NANDN U15710 ( .A(n15285), .B(n15284), .Z(n15289) );
  NAND U15711 ( .A(n15287), .B(n15286), .Z(n15288) );
  AND U15712 ( .A(n15289), .B(n15288), .Z(n15337) );
  XOR U15713 ( .A(n15338), .B(n15337), .Z(n15339) );
  NANDN U15714 ( .A(n15291), .B(n15290), .Z(n15295) );
  NANDN U15715 ( .A(n15293), .B(n15292), .Z(n15294) );
  NAND U15716 ( .A(n15295), .B(n15294), .Z(n15340) );
  XOR U15717 ( .A(n15339), .B(n15340), .Z(n15307) );
  OR U15718 ( .A(n15297), .B(n15296), .Z(n15301) );
  NANDN U15719 ( .A(n15299), .B(n15298), .Z(n15300) );
  NAND U15720 ( .A(n15301), .B(n15300), .Z(n15308) );
  XNOR U15721 ( .A(n15307), .B(n15308), .Z(n15309) );
  XNOR U15722 ( .A(n15310), .B(n15309), .Z(n15343) );
  XNOR U15723 ( .A(n15343), .B(sreg[1387]), .Z(n15345) );
  NAND U15724 ( .A(n15302), .B(sreg[1386]), .Z(n15306) );
  OR U15725 ( .A(n15304), .B(n15303), .Z(n15305) );
  AND U15726 ( .A(n15306), .B(n15305), .Z(n15344) );
  XOR U15727 ( .A(n15345), .B(n15344), .Z(c[1387]) );
  NANDN U15728 ( .A(n15308), .B(n15307), .Z(n15312) );
  NAND U15729 ( .A(n15310), .B(n15309), .Z(n15311) );
  NAND U15730 ( .A(n15312), .B(n15311), .Z(n15351) );
  NAND U15731 ( .A(b[0]), .B(a[372]), .Z(n15313) );
  XNOR U15732 ( .A(b[1]), .B(n15313), .Z(n15315) );
  NAND U15733 ( .A(n68), .B(a[371]), .Z(n15314) );
  AND U15734 ( .A(n15315), .B(n15314), .Z(n15368) );
  XOR U15735 ( .A(a[368]), .B(n42197), .Z(n15357) );
  NANDN U15736 ( .A(n15357), .B(n42173), .Z(n15318) );
  NANDN U15737 ( .A(n15316), .B(n42172), .Z(n15317) );
  NAND U15738 ( .A(n15318), .B(n15317), .Z(n15366) );
  NAND U15739 ( .A(b[7]), .B(a[364]), .Z(n15367) );
  XNOR U15740 ( .A(n15366), .B(n15367), .Z(n15369) );
  XOR U15741 ( .A(n15368), .B(n15369), .Z(n15375) );
  NANDN U15742 ( .A(n15319), .B(n42093), .Z(n15321) );
  XOR U15743 ( .A(n42134), .B(a[370]), .Z(n15360) );
  NANDN U15744 ( .A(n15360), .B(n42095), .Z(n15320) );
  NAND U15745 ( .A(n15321), .B(n15320), .Z(n15373) );
  NANDN U15746 ( .A(n15322), .B(n42231), .Z(n15324) );
  XOR U15747 ( .A(n192), .B(a[366]), .Z(n15363) );
  NANDN U15748 ( .A(n15363), .B(n42234), .Z(n15323) );
  AND U15749 ( .A(n15324), .B(n15323), .Z(n15372) );
  XNOR U15750 ( .A(n15373), .B(n15372), .Z(n15374) );
  XNOR U15751 ( .A(n15375), .B(n15374), .Z(n15379) );
  NANDN U15752 ( .A(n15326), .B(n15325), .Z(n15330) );
  NAND U15753 ( .A(n15328), .B(n15327), .Z(n15329) );
  AND U15754 ( .A(n15330), .B(n15329), .Z(n15378) );
  XOR U15755 ( .A(n15379), .B(n15378), .Z(n15380) );
  NANDN U15756 ( .A(n15332), .B(n15331), .Z(n15336) );
  NANDN U15757 ( .A(n15334), .B(n15333), .Z(n15335) );
  NAND U15758 ( .A(n15336), .B(n15335), .Z(n15381) );
  XOR U15759 ( .A(n15380), .B(n15381), .Z(n15348) );
  OR U15760 ( .A(n15338), .B(n15337), .Z(n15342) );
  NANDN U15761 ( .A(n15340), .B(n15339), .Z(n15341) );
  NAND U15762 ( .A(n15342), .B(n15341), .Z(n15349) );
  XNOR U15763 ( .A(n15348), .B(n15349), .Z(n15350) );
  XNOR U15764 ( .A(n15351), .B(n15350), .Z(n15384) );
  XNOR U15765 ( .A(n15384), .B(sreg[1388]), .Z(n15386) );
  NAND U15766 ( .A(n15343), .B(sreg[1387]), .Z(n15347) );
  OR U15767 ( .A(n15345), .B(n15344), .Z(n15346) );
  AND U15768 ( .A(n15347), .B(n15346), .Z(n15385) );
  XOR U15769 ( .A(n15386), .B(n15385), .Z(c[1388]) );
  NANDN U15770 ( .A(n15349), .B(n15348), .Z(n15353) );
  NAND U15771 ( .A(n15351), .B(n15350), .Z(n15352) );
  NAND U15772 ( .A(n15353), .B(n15352), .Z(n15392) );
  NAND U15773 ( .A(b[0]), .B(a[373]), .Z(n15354) );
  XNOR U15774 ( .A(b[1]), .B(n15354), .Z(n15356) );
  NAND U15775 ( .A(n68), .B(a[372]), .Z(n15355) );
  AND U15776 ( .A(n15356), .B(n15355), .Z(n15409) );
  XOR U15777 ( .A(a[369]), .B(n42197), .Z(n15398) );
  NANDN U15778 ( .A(n15398), .B(n42173), .Z(n15359) );
  NANDN U15779 ( .A(n15357), .B(n42172), .Z(n15358) );
  NAND U15780 ( .A(n15359), .B(n15358), .Z(n15407) );
  NAND U15781 ( .A(b[7]), .B(a[365]), .Z(n15408) );
  XNOR U15782 ( .A(n15407), .B(n15408), .Z(n15410) );
  XOR U15783 ( .A(n15409), .B(n15410), .Z(n15416) );
  NANDN U15784 ( .A(n15360), .B(n42093), .Z(n15362) );
  XOR U15785 ( .A(n42134), .B(a[371]), .Z(n15401) );
  NANDN U15786 ( .A(n15401), .B(n42095), .Z(n15361) );
  NAND U15787 ( .A(n15362), .B(n15361), .Z(n15414) );
  NANDN U15788 ( .A(n15363), .B(n42231), .Z(n15365) );
  XOR U15789 ( .A(n192), .B(a[367]), .Z(n15404) );
  NANDN U15790 ( .A(n15404), .B(n42234), .Z(n15364) );
  AND U15791 ( .A(n15365), .B(n15364), .Z(n15413) );
  XNOR U15792 ( .A(n15414), .B(n15413), .Z(n15415) );
  XNOR U15793 ( .A(n15416), .B(n15415), .Z(n15420) );
  NANDN U15794 ( .A(n15367), .B(n15366), .Z(n15371) );
  NAND U15795 ( .A(n15369), .B(n15368), .Z(n15370) );
  AND U15796 ( .A(n15371), .B(n15370), .Z(n15419) );
  XOR U15797 ( .A(n15420), .B(n15419), .Z(n15421) );
  NANDN U15798 ( .A(n15373), .B(n15372), .Z(n15377) );
  NANDN U15799 ( .A(n15375), .B(n15374), .Z(n15376) );
  NAND U15800 ( .A(n15377), .B(n15376), .Z(n15422) );
  XOR U15801 ( .A(n15421), .B(n15422), .Z(n15389) );
  OR U15802 ( .A(n15379), .B(n15378), .Z(n15383) );
  NANDN U15803 ( .A(n15381), .B(n15380), .Z(n15382) );
  NAND U15804 ( .A(n15383), .B(n15382), .Z(n15390) );
  XNOR U15805 ( .A(n15389), .B(n15390), .Z(n15391) );
  XNOR U15806 ( .A(n15392), .B(n15391), .Z(n15425) );
  XNOR U15807 ( .A(n15425), .B(sreg[1389]), .Z(n15427) );
  NAND U15808 ( .A(n15384), .B(sreg[1388]), .Z(n15388) );
  OR U15809 ( .A(n15386), .B(n15385), .Z(n15387) );
  AND U15810 ( .A(n15388), .B(n15387), .Z(n15426) );
  XOR U15811 ( .A(n15427), .B(n15426), .Z(c[1389]) );
  NANDN U15812 ( .A(n15390), .B(n15389), .Z(n15394) );
  NAND U15813 ( .A(n15392), .B(n15391), .Z(n15393) );
  NAND U15814 ( .A(n15394), .B(n15393), .Z(n15433) );
  NAND U15815 ( .A(b[0]), .B(a[374]), .Z(n15395) );
  XNOR U15816 ( .A(b[1]), .B(n15395), .Z(n15397) );
  NAND U15817 ( .A(n68), .B(a[373]), .Z(n15396) );
  AND U15818 ( .A(n15397), .B(n15396), .Z(n15450) );
  XOR U15819 ( .A(a[370]), .B(n42197), .Z(n15439) );
  NANDN U15820 ( .A(n15439), .B(n42173), .Z(n15400) );
  NANDN U15821 ( .A(n15398), .B(n42172), .Z(n15399) );
  NAND U15822 ( .A(n15400), .B(n15399), .Z(n15448) );
  NAND U15823 ( .A(b[7]), .B(a[366]), .Z(n15449) );
  XNOR U15824 ( .A(n15448), .B(n15449), .Z(n15451) );
  XOR U15825 ( .A(n15450), .B(n15451), .Z(n15457) );
  NANDN U15826 ( .A(n15401), .B(n42093), .Z(n15403) );
  XOR U15827 ( .A(n42134), .B(a[372]), .Z(n15442) );
  NANDN U15828 ( .A(n15442), .B(n42095), .Z(n15402) );
  NAND U15829 ( .A(n15403), .B(n15402), .Z(n15455) );
  NANDN U15830 ( .A(n15404), .B(n42231), .Z(n15406) );
  XOR U15831 ( .A(n192), .B(a[368]), .Z(n15445) );
  NANDN U15832 ( .A(n15445), .B(n42234), .Z(n15405) );
  AND U15833 ( .A(n15406), .B(n15405), .Z(n15454) );
  XNOR U15834 ( .A(n15455), .B(n15454), .Z(n15456) );
  XNOR U15835 ( .A(n15457), .B(n15456), .Z(n15461) );
  NANDN U15836 ( .A(n15408), .B(n15407), .Z(n15412) );
  NAND U15837 ( .A(n15410), .B(n15409), .Z(n15411) );
  AND U15838 ( .A(n15412), .B(n15411), .Z(n15460) );
  XOR U15839 ( .A(n15461), .B(n15460), .Z(n15462) );
  NANDN U15840 ( .A(n15414), .B(n15413), .Z(n15418) );
  NANDN U15841 ( .A(n15416), .B(n15415), .Z(n15417) );
  NAND U15842 ( .A(n15418), .B(n15417), .Z(n15463) );
  XOR U15843 ( .A(n15462), .B(n15463), .Z(n15430) );
  OR U15844 ( .A(n15420), .B(n15419), .Z(n15424) );
  NANDN U15845 ( .A(n15422), .B(n15421), .Z(n15423) );
  NAND U15846 ( .A(n15424), .B(n15423), .Z(n15431) );
  XNOR U15847 ( .A(n15430), .B(n15431), .Z(n15432) );
  XNOR U15848 ( .A(n15433), .B(n15432), .Z(n15466) );
  XNOR U15849 ( .A(n15466), .B(sreg[1390]), .Z(n15468) );
  NAND U15850 ( .A(n15425), .B(sreg[1389]), .Z(n15429) );
  OR U15851 ( .A(n15427), .B(n15426), .Z(n15428) );
  AND U15852 ( .A(n15429), .B(n15428), .Z(n15467) );
  XOR U15853 ( .A(n15468), .B(n15467), .Z(c[1390]) );
  NANDN U15854 ( .A(n15431), .B(n15430), .Z(n15435) );
  NAND U15855 ( .A(n15433), .B(n15432), .Z(n15434) );
  NAND U15856 ( .A(n15435), .B(n15434), .Z(n15474) );
  NAND U15857 ( .A(b[0]), .B(a[375]), .Z(n15436) );
  XNOR U15858 ( .A(b[1]), .B(n15436), .Z(n15438) );
  NAND U15859 ( .A(n68), .B(a[374]), .Z(n15437) );
  AND U15860 ( .A(n15438), .B(n15437), .Z(n15491) );
  XOR U15861 ( .A(a[371]), .B(n42197), .Z(n15480) );
  NANDN U15862 ( .A(n15480), .B(n42173), .Z(n15441) );
  NANDN U15863 ( .A(n15439), .B(n42172), .Z(n15440) );
  NAND U15864 ( .A(n15441), .B(n15440), .Z(n15489) );
  NAND U15865 ( .A(b[7]), .B(a[367]), .Z(n15490) );
  XNOR U15866 ( .A(n15489), .B(n15490), .Z(n15492) );
  XOR U15867 ( .A(n15491), .B(n15492), .Z(n15498) );
  NANDN U15868 ( .A(n15442), .B(n42093), .Z(n15444) );
  XOR U15869 ( .A(n42134), .B(a[373]), .Z(n15483) );
  NANDN U15870 ( .A(n15483), .B(n42095), .Z(n15443) );
  NAND U15871 ( .A(n15444), .B(n15443), .Z(n15496) );
  NANDN U15872 ( .A(n15445), .B(n42231), .Z(n15447) );
  XOR U15873 ( .A(n192), .B(a[369]), .Z(n15486) );
  NANDN U15874 ( .A(n15486), .B(n42234), .Z(n15446) );
  AND U15875 ( .A(n15447), .B(n15446), .Z(n15495) );
  XNOR U15876 ( .A(n15496), .B(n15495), .Z(n15497) );
  XNOR U15877 ( .A(n15498), .B(n15497), .Z(n15502) );
  NANDN U15878 ( .A(n15449), .B(n15448), .Z(n15453) );
  NAND U15879 ( .A(n15451), .B(n15450), .Z(n15452) );
  AND U15880 ( .A(n15453), .B(n15452), .Z(n15501) );
  XOR U15881 ( .A(n15502), .B(n15501), .Z(n15503) );
  NANDN U15882 ( .A(n15455), .B(n15454), .Z(n15459) );
  NANDN U15883 ( .A(n15457), .B(n15456), .Z(n15458) );
  NAND U15884 ( .A(n15459), .B(n15458), .Z(n15504) );
  XOR U15885 ( .A(n15503), .B(n15504), .Z(n15471) );
  OR U15886 ( .A(n15461), .B(n15460), .Z(n15465) );
  NANDN U15887 ( .A(n15463), .B(n15462), .Z(n15464) );
  NAND U15888 ( .A(n15465), .B(n15464), .Z(n15472) );
  XNOR U15889 ( .A(n15471), .B(n15472), .Z(n15473) );
  XNOR U15890 ( .A(n15474), .B(n15473), .Z(n15507) );
  XNOR U15891 ( .A(n15507), .B(sreg[1391]), .Z(n15509) );
  NAND U15892 ( .A(n15466), .B(sreg[1390]), .Z(n15470) );
  OR U15893 ( .A(n15468), .B(n15467), .Z(n15469) );
  AND U15894 ( .A(n15470), .B(n15469), .Z(n15508) );
  XOR U15895 ( .A(n15509), .B(n15508), .Z(c[1391]) );
  NANDN U15896 ( .A(n15472), .B(n15471), .Z(n15476) );
  NAND U15897 ( .A(n15474), .B(n15473), .Z(n15475) );
  NAND U15898 ( .A(n15476), .B(n15475), .Z(n15515) );
  NAND U15899 ( .A(b[0]), .B(a[376]), .Z(n15477) );
  XNOR U15900 ( .A(b[1]), .B(n15477), .Z(n15479) );
  NAND U15901 ( .A(n68), .B(a[375]), .Z(n15478) );
  AND U15902 ( .A(n15479), .B(n15478), .Z(n15532) );
  XOR U15903 ( .A(a[372]), .B(n42197), .Z(n15521) );
  NANDN U15904 ( .A(n15521), .B(n42173), .Z(n15482) );
  NANDN U15905 ( .A(n15480), .B(n42172), .Z(n15481) );
  NAND U15906 ( .A(n15482), .B(n15481), .Z(n15530) );
  NAND U15907 ( .A(b[7]), .B(a[368]), .Z(n15531) );
  XNOR U15908 ( .A(n15530), .B(n15531), .Z(n15533) );
  XOR U15909 ( .A(n15532), .B(n15533), .Z(n15539) );
  NANDN U15910 ( .A(n15483), .B(n42093), .Z(n15485) );
  XOR U15911 ( .A(n42134), .B(a[374]), .Z(n15524) );
  NANDN U15912 ( .A(n15524), .B(n42095), .Z(n15484) );
  NAND U15913 ( .A(n15485), .B(n15484), .Z(n15537) );
  NANDN U15914 ( .A(n15486), .B(n42231), .Z(n15488) );
  XOR U15915 ( .A(n192), .B(a[370]), .Z(n15527) );
  NANDN U15916 ( .A(n15527), .B(n42234), .Z(n15487) );
  AND U15917 ( .A(n15488), .B(n15487), .Z(n15536) );
  XNOR U15918 ( .A(n15537), .B(n15536), .Z(n15538) );
  XNOR U15919 ( .A(n15539), .B(n15538), .Z(n15543) );
  NANDN U15920 ( .A(n15490), .B(n15489), .Z(n15494) );
  NAND U15921 ( .A(n15492), .B(n15491), .Z(n15493) );
  AND U15922 ( .A(n15494), .B(n15493), .Z(n15542) );
  XOR U15923 ( .A(n15543), .B(n15542), .Z(n15544) );
  NANDN U15924 ( .A(n15496), .B(n15495), .Z(n15500) );
  NANDN U15925 ( .A(n15498), .B(n15497), .Z(n15499) );
  NAND U15926 ( .A(n15500), .B(n15499), .Z(n15545) );
  XOR U15927 ( .A(n15544), .B(n15545), .Z(n15512) );
  OR U15928 ( .A(n15502), .B(n15501), .Z(n15506) );
  NANDN U15929 ( .A(n15504), .B(n15503), .Z(n15505) );
  NAND U15930 ( .A(n15506), .B(n15505), .Z(n15513) );
  XNOR U15931 ( .A(n15512), .B(n15513), .Z(n15514) );
  XNOR U15932 ( .A(n15515), .B(n15514), .Z(n15548) );
  XNOR U15933 ( .A(n15548), .B(sreg[1392]), .Z(n15550) );
  NAND U15934 ( .A(n15507), .B(sreg[1391]), .Z(n15511) );
  OR U15935 ( .A(n15509), .B(n15508), .Z(n15510) );
  AND U15936 ( .A(n15511), .B(n15510), .Z(n15549) );
  XOR U15937 ( .A(n15550), .B(n15549), .Z(c[1392]) );
  NANDN U15938 ( .A(n15513), .B(n15512), .Z(n15517) );
  NAND U15939 ( .A(n15515), .B(n15514), .Z(n15516) );
  NAND U15940 ( .A(n15517), .B(n15516), .Z(n15556) );
  NAND U15941 ( .A(b[0]), .B(a[377]), .Z(n15518) );
  XNOR U15942 ( .A(b[1]), .B(n15518), .Z(n15520) );
  NAND U15943 ( .A(n68), .B(a[376]), .Z(n15519) );
  AND U15944 ( .A(n15520), .B(n15519), .Z(n15573) );
  XOR U15945 ( .A(a[373]), .B(n42197), .Z(n15562) );
  NANDN U15946 ( .A(n15562), .B(n42173), .Z(n15523) );
  NANDN U15947 ( .A(n15521), .B(n42172), .Z(n15522) );
  NAND U15948 ( .A(n15523), .B(n15522), .Z(n15571) );
  NAND U15949 ( .A(b[7]), .B(a[369]), .Z(n15572) );
  XNOR U15950 ( .A(n15571), .B(n15572), .Z(n15574) );
  XOR U15951 ( .A(n15573), .B(n15574), .Z(n15580) );
  NANDN U15952 ( .A(n15524), .B(n42093), .Z(n15526) );
  XOR U15953 ( .A(n42134), .B(a[375]), .Z(n15565) );
  NANDN U15954 ( .A(n15565), .B(n42095), .Z(n15525) );
  NAND U15955 ( .A(n15526), .B(n15525), .Z(n15578) );
  NANDN U15956 ( .A(n15527), .B(n42231), .Z(n15529) );
  XOR U15957 ( .A(n193), .B(a[371]), .Z(n15568) );
  NANDN U15958 ( .A(n15568), .B(n42234), .Z(n15528) );
  AND U15959 ( .A(n15529), .B(n15528), .Z(n15577) );
  XNOR U15960 ( .A(n15578), .B(n15577), .Z(n15579) );
  XNOR U15961 ( .A(n15580), .B(n15579), .Z(n15584) );
  NANDN U15962 ( .A(n15531), .B(n15530), .Z(n15535) );
  NAND U15963 ( .A(n15533), .B(n15532), .Z(n15534) );
  AND U15964 ( .A(n15535), .B(n15534), .Z(n15583) );
  XOR U15965 ( .A(n15584), .B(n15583), .Z(n15585) );
  NANDN U15966 ( .A(n15537), .B(n15536), .Z(n15541) );
  NANDN U15967 ( .A(n15539), .B(n15538), .Z(n15540) );
  NAND U15968 ( .A(n15541), .B(n15540), .Z(n15586) );
  XOR U15969 ( .A(n15585), .B(n15586), .Z(n15553) );
  OR U15970 ( .A(n15543), .B(n15542), .Z(n15547) );
  NANDN U15971 ( .A(n15545), .B(n15544), .Z(n15546) );
  NAND U15972 ( .A(n15547), .B(n15546), .Z(n15554) );
  XNOR U15973 ( .A(n15553), .B(n15554), .Z(n15555) );
  XNOR U15974 ( .A(n15556), .B(n15555), .Z(n15589) );
  XNOR U15975 ( .A(n15589), .B(sreg[1393]), .Z(n15591) );
  NAND U15976 ( .A(n15548), .B(sreg[1392]), .Z(n15552) );
  OR U15977 ( .A(n15550), .B(n15549), .Z(n15551) );
  AND U15978 ( .A(n15552), .B(n15551), .Z(n15590) );
  XOR U15979 ( .A(n15591), .B(n15590), .Z(c[1393]) );
  NANDN U15980 ( .A(n15554), .B(n15553), .Z(n15558) );
  NAND U15981 ( .A(n15556), .B(n15555), .Z(n15557) );
  NAND U15982 ( .A(n15558), .B(n15557), .Z(n15597) );
  NAND U15983 ( .A(b[0]), .B(a[378]), .Z(n15559) );
  XNOR U15984 ( .A(b[1]), .B(n15559), .Z(n15561) );
  NAND U15985 ( .A(n69), .B(a[377]), .Z(n15560) );
  AND U15986 ( .A(n15561), .B(n15560), .Z(n15614) );
  XOR U15987 ( .A(a[374]), .B(n42197), .Z(n15603) );
  NANDN U15988 ( .A(n15603), .B(n42173), .Z(n15564) );
  NANDN U15989 ( .A(n15562), .B(n42172), .Z(n15563) );
  NAND U15990 ( .A(n15564), .B(n15563), .Z(n15612) );
  NAND U15991 ( .A(b[7]), .B(a[370]), .Z(n15613) );
  XNOR U15992 ( .A(n15612), .B(n15613), .Z(n15615) );
  XOR U15993 ( .A(n15614), .B(n15615), .Z(n15621) );
  NANDN U15994 ( .A(n15565), .B(n42093), .Z(n15567) );
  XOR U15995 ( .A(n42134), .B(a[376]), .Z(n15606) );
  NANDN U15996 ( .A(n15606), .B(n42095), .Z(n15566) );
  NAND U15997 ( .A(n15567), .B(n15566), .Z(n15619) );
  NANDN U15998 ( .A(n15568), .B(n42231), .Z(n15570) );
  XOR U15999 ( .A(n193), .B(a[372]), .Z(n15609) );
  NANDN U16000 ( .A(n15609), .B(n42234), .Z(n15569) );
  AND U16001 ( .A(n15570), .B(n15569), .Z(n15618) );
  XNOR U16002 ( .A(n15619), .B(n15618), .Z(n15620) );
  XNOR U16003 ( .A(n15621), .B(n15620), .Z(n15625) );
  NANDN U16004 ( .A(n15572), .B(n15571), .Z(n15576) );
  NAND U16005 ( .A(n15574), .B(n15573), .Z(n15575) );
  AND U16006 ( .A(n15576), .B(n15575), .Z(n15624) );
  XOR U16007 ( .A(n15625), .B(n15624), .Z(n15626) );
  NANDN U16008 ( .A(n15578), .B(n15577), .Z(n15582) );
  NANDN U16009 ( .A(n15580), .B(n15579), .Z(n15581) );
  NAND U16010 ( .A(n15582), .B(n15581), .Z(n15627) );
  XOR U16011 ( .A(n15626), .B(n15627), .Z(n15594) );
  OR U16012 ( .A(n15584), .B(n15583), .Z(n15588) );
  NANDN U16013 ( .A(n15586), .B(n15585), .Z(n15587) );
  NAND U16014 ( .A(n15588), .B(n15587), .Z(n15595) );
  XNOR U16015 ( .A(n15594), .B(n15595), .Z(n15596) );
  XNOR U16016 ( .A(n15597), .B(n15596), .Z(n15630) );
  XNOR U16017 ( .A(n15630), .B(sreg[1394]), .Z(n15632) );
  NAND U16018 ( .A(n15589), .B(sreg[1393]), .Z(n15593) );
  OR U16019 ( .A(n15591), .B(n15590), .Z(n15592) );
  AND U16020 ( .A(n15593), .B(n15592), .Z(n15631) );
  XOR U16021 ( .A(n15632), .B(n15631), .Z(c[1394]) );
  NANDN U16022 ( .A(n15595), .B(n15594), .Z(n15599) );
  NAND U16023 ( .A(n15597), .B(n15596), .Z(n15598) );
  NAND U16024 ( .A(n15599), .B(n15598), .Z(n15638) );
  NAND U16025 ( .A(b[0]), .B(a[379]), .Z(n15600) );
  XNOR U16026 ( .A(b[1]), .B(n15600), .Z(n15602) );
  NAND U16027 ( .A(n69), .B(a[378]), .Z(n15601) );
  AND U16028 ( .A(n15602), .B(n15601), .Z(n15655) );
  XOR U16029 ( .A(a[375]), .B(n42197), .Z(n15644) );
  NANDN U16030 ( .A(n15644), .B(n42173), .Z(n15605) );
  NANDN U16031 ( .A(n15603), .B(n42172), .Z(n15604) );
  NAND U16032 ( .A(n15605), .B(n15604), .Z(n15653) );
  NAND U16033 ( .A(b[7]), .B(a[371]), .Z(n15654) );
  XNOR U16034 ( .A(n15653), .B(n15654), .Z(n15656) );
  XOR U16035 ( .A(n15655), .B(n15656), .Z(n15662) );
  NANDN U16036 ( .A(n15606), .B(n42093), .Z(n15608) );
  XOR U16037 ( .A(n42134), .B(a[377]), .Z(n15647) );
  NANDN U16038 ( .A(n15647), .B(n42095), .Z(n15607) );
  NAND U16039 ( .A(n15608), .B(n15607), .Z(n15660) );
  NANDN U16040 ( .A(n15609), .B(n42231), .Z(n15611) );
  XOR U16041 ( .A(n193), .B(a[373]), .Z(n15650) );
  NANDN U16042 ( .A(n15650), .B(n42234), .Z(n15610) );
  AND U16043 ( .A(n15611), .B(n15610), .Z(n15659) );
  XNOR U16044 ( .A(n15660), .B(n15659), .Z(n15661) );
  XNOR U16045 ( .A(n15662), .B(n15661), .Z(n15666) );
  NANDN U16046 ( .A(n15613), .B(n15612), .Z(n15617) );
  NAND U16047 ( .A(n15615), .B(n15614), .Z(n15616) );
  AND U16048 ( .A(n15617), .B(n15616), .Z(n15665) );
  XOR U16049 ( .A(n15666), .B(n15665), .Z(n15667) );
  NANDN U16050 ( .A(n15619), .B(n15618), .Z(n15623) );
  NANDN U16051 ( .A(n15621), .B(n15620), .Z(n15622) );
  NAND U16052 ( .A(n15623), .B(n15622), .Z(n15668) );
  XOR U16053 ( .A(n15667), .B(n15668), .Z(n15635) );
  OR U16054 ( .A(n15625), .B(n15624), .Z(n15629) );
  NANDN U16055 ( .A(n15627), .B(n15626), .Z(n15628) );
  NAND U16056 ( .A(n15629), .B(n15628), .Z(n15636) );
  XNOR U16057 ( .A(n15635), .B(n15636), .Z(n15637) );
  XNOR U16058 ( .A(n15638), .B(n15637), .Z(n15671) );
  XNOR U16059 ( .A(n15671), .B(sreg[1395]), .Z(n15673) );
  NAND U16060 ( .A(n15630), .B(sreg[1394]), .Z(n15634) );
  OR U16061 ( .A(n15632), .B(n15631), .Z(n15633) );
  AND U16062 ( .A(n15634), .B(n15633), .Z(n15672) );
  XOR U16063 ( .A(n15673), .B(n15672), .Z(c[1395]) );
  NANDN U16064 ( .A(n15636), .B(n15635), .Z(n15640) );
  NAND U16065 ( .A(n15638), .B(n15637), .Z(n15639) );
  NAND U16066 ( .A(n15640), .B(n15639), .Z(n15679) );
  NAND U16067 ( .A(b[0]), .B(a[380]), .Z(n15641) );
  XNOR U16068 ( .A(b[1]), .B(n15641), .Z(n15643) );
  NAND U16069 ( .A(n69), .B(a[379]), .Z(n15642) );
  AND U16070 ( .A(n15643), .B(n15642), .Z(n15696) );
  XOR U16071 ( .A(a[376]), .B(n42197), .Z(n15685) );
  NANDN U16072 ( .A(n15685), .B(n42173), .Z(n15646) );
  NANDN U16073 ( .A(n15644), .B(n42172), .Z(n15645) );
  NAND U16074 ( .A(n15646), .B(n15645), .Z(n15694) );
  NAND U16075 ( .A(b[7]), .B(a[372]), .Z(n15695) );
  XNOR U16076 ( .A(n15694), .B(n15695), .Z(n15697) );
  XOR U16077 ( .A(n15696), .B(n15697), .Z(n15703) );
  NANDN U16078 ( .A(n15647), .B(n42093), .Z(n15649) );
  XOR U16079 ( .A(n42134), .B(a[378]), .Z(n15688) );
  NANDN U16080 ( .A(n15688), .B(n42095), .Z(n15648) );
  NAND U16081 ( .A(n15649), .B(n15648), .Z(n15701) );
  NANDN U16082 ( .A(n15650), .B(n42231), .Z(n15652) );
  XOR U16083 ( .A(n193), .B(a[374]), .Z(n15691) );
  NANDN U16084 ( .A(n15691), .B(n42234), .Z(n15651) );
  AND U16085 ( .A(n15652), .B(n15651), .Z(n15700) );
  XNOR U16086 ( .A(n15701), .B(n15700), .Z(n15702) );
  XNOR U16087 ( .A(n15703), .B(n15702), .Z(n15707) );
  NANDN U16088 ( .A(n15654), .B(n15653), .Z(n15658) );
  NAND U16089 ( .A(n15656), .B(n15655), .Z(n15657) );
  AND U16090 ( .A(n15658), .B(n15657), .Z(n15706) );
  XOR U16091 ( .A(n15707), .B(n15706), .Z(n15708) );
  NANDN U16092 ( .A(n15660), .B(n15659), .Z(n15664) );
  NANDN U16093 ( .A(n15662), .B(n15661), .Z(n15663) );
  NAND U16094 ( .A(n15664), .B(n15663), .Z(n15709) );
  XOR U16095 ( .A(n15708), .B(n15709), .Z(n15676) );
  OR U16096 ( .A(n15666), .B(n15665), .Z(n15670) );
  NANDN U16097 ( .A(n15668), .B(n15667), .Z(n15669) );
  NAND U16098 ( .A(n15670), .B(n15669), .Z(n15677) );
  XNOR U16099 ( .A(n15676), .B(n15677), .Z(n15678) );
  XNOR U16100 ( .A(n15679), .B(n15678), .Z(n15712) );
  XNOR U16101 ( .A(n15712), .B(sreg[1396]), .Z(n15714) );
  NAND U16102 ( .A(n15671), .B(sreg[1395]), .Z(n15675) );
  OR U16103 ( .A(n15673), .B(n15672), .Z(n15674) );
  AND U16104 ( .A(n15675), .B(n15674), .Z(n15713) );
  XOR U16105 ( .A(n15714), .B(n15713), .Z(c[1396]) );
  NANDN U16106 ( .A(n15677), .B(n15676), .Z(n15681) );
  NAND U16107 ( .A(n15679), .B(n15678), .Z(n15680) );
  NAND U16108 ( .A(n15681), .B(n15680), .Z(n15720) );
  NAND U16109 ( .A(b[0]), .B(a[381]), .Z(n15682) );
  XNOR U16110 ( .A(b[1]), .B(n15682), .Z(n15684) );
  NAND U16111 ( .A(n69), .B(a[380]), .Z(n15683) );
  AND U16112 ( .A(n15684), .B(n15683), .Z(n15737) );
  XOR U16113 ( .A(a[377]), .B(n42197), .Z(n15726) );
  NANDN U16114 ( .A(n15726), .B(n42173), .Z(n15687) );
  NANDN U16115 ( .A(n15685), .B(n42172), .Z(n15686) );
  NAND U16116 ( .A(n15687), .B(n15686), .Z(n15735) );
  NAND U16117 ( .A(b[7]), .B(a[373]), .Z(n15736) );
  XNOR U16118 ( .A(n15735), .B(n15736), .Z(n15738) );
  XOR U16119 ( .A(n15737), .B(n15738), .Z(n15744) );
  NANDN U16120 ( .A(n15688), .B(n42093), .Z(n15690) );
  XOR U16121 ( .A(n42134), .B(a[379]), .Z(n15729) );
  NANDN U16122 ( .A(n15729), .B(n42095), .Z(n15689) );
  NAND U16123 ( .A(n15690), .B(n15689), .Z(n15742) );
  NANDN U16124 ( .A(n15691), .B(n42231), .Z(n15693) );
  XOR U16125 ( .A(n193), .B(a[375]), .Z(n15732) );
  NANDN U16126 ( .A(n15732), .B(n42234), .Z(n15692) );
  AND U16127 ( .A(n15693), .B(n15692), .Z(n15741) );
  XNOR U16128 ( .A(n15742), .B(n15741), .Z(n15743) );
  XNOR U16129 ( .A(n15744), .B(n15743), .Z(n15748) );
  NANDN U16130 ( .A(n15695), .B(n15694), .Z(n15699) );
  NAND U16131 ( .A(n15697), .B(n15696), .Z(n15698) );
  AND U16132 ( .A(n15699), .B(n15698), .Z(n15747) );
  XOR U16133 ( .A(n15748), .B(n15747), .Z(n15749) );
  NANDN U16134 ( .A(n15701), .B(n15700), .Z(n15705) );
  NANDN U16135 ( .A(n15703), .B(n15702), .Z(n15704) );
  NAND U16136 ( .A(n15705), .B(n15704), .Z(n15750) );
  XOR U16137 ( .A(n15749), .B(n15750), .Z(n15717) );
  OR U16138 ( .A(n15707), .B(n15706), .Z(n15711) );
  NANDN U16139 ( .A(n15709), .B(n15708), .Z(n15710) );
  NAND U16140 ( .A(n15711), .B(n15710), .Z(n15718) );
  XNOR U16141 ( .A(n15717), .B(n15718), .Z(n15719) );
  XNOR U16142 ( .A(n15720), .B(n15719), .Z(n15753) );
  XNOR U16143 ( .A(n15753), .B(sreg[1397]), .Z(n15755) );
  NAND U16144 ( .A(n15712), .B(sreg[1396]), .Z(n15716) );
  OR U16145 ( .A(n15714), .B(n15713), .Z(n15715) );
  AND U16146 ( .A(n15716), .B(n15715), .Z(n15754) );
  XOR U16147 ( .A(n15755), .B(n15754), .Z(c[1397]) );
  NANDN U16148 ( .A(n15718), .B(n15717), .Z(n15722) );
  NAND U16149 ( .A(n15720), .B(n15719), .Z(n15721) );
  NAND U16150 ( .A(n15722), .B(n15721), .Z(n15761) );
  NAND U16151 ( .A(b[0]), .B(a[382]), .Z(n15723) );
  XNOR U16152 ( .A(b[1]), .B(n15723), .Z(n15725) );
  NAND U16153 ( .A(n69), .B(a[381]), .Z(n15724) );
  AND U16154 ( .A(n15725), .B(n15724), .Z(n15778) );
  XOR U16155 ( .A(a[378]), .B(n42197), .Z(n15767) );
  NANDN U16156 ( .A(n15767), .B(n42173), .Z(n15728) );
  NANDN U16157 ( .A(n15726), .B(n42172), .Z(n15727) );
  NAND U16158 ( .A(n15728), .B(n15727), .Z(n15776) );
  NAND U16159 ( .A(b[7]), .B(a[374]), .Z(n15777) );
  XNOR U16160 ( .A(n15776), .B(n15777), .Z(n15779) );
  XOR U16161 ( .A(n15778), .B(n15779), .Z(n15785) );
  NANDN U16162 ( .A(n15729), .B(n42093), .Z(n15731) );
  XOR U16163 ( .A(n42134), .B(a[380]), .Z(n15770) );
  NANDN U16164 ( .A(n15770), .B(n42095), .Z(n15730) );
  NAND U16165 ( .A(n15731), .B(n15730), .Z(n15783) );
  NANDN U16166 ( .A(n15732), .B(n42231), .Z(n15734) );
  XOR U16167 ( .A(n193), .B(a[376]), .Z(n15773) );
  NANDN U16168 ( .A(n15773), .B(n42234), .Z(n15733) );
  AND U16169 ( .A(n15734), .B(n15733), .Z(n15782) );
  XNOR U16170 ( .A(n15783), .B(n15782), .Z(n15784) );
  XNOR U16171 ( .A(n15785), .B(n15784), .Z(n15789) );
  NANDN U16172 ( .A(n15736), .B(n15735), .Z(n15740) );
  NAND U16173 ( .A(n15738), .B(n15737), .Z(n15739) );
  AND U16174 ( .A(n15740), .B(n15739), .Z(n15788) );
  XOR U16175 ( .A(n15789), .B(n15788), .Z(n15790) );
  NANDN U16176 ( .A(n15742), .B(n15741), .Z(n15746) );
  NANDN U16177 ( .A(n15744), .B(n15743), .Z(n15745) );
  NAND U16178 ( .A(n15746), .B(n15745), .Z(n15791) );
  XOR U16179 ( .A(n15790), .B(n15791), .Z(n15758) );
  OR U16180 ( .A(n15748), .B(n15747), .Z(n15752) );
  NANDN U16181 ( .A(n15750), .B(n15749), .Z(n15751) );
  NAND U16182 ( .A(n15752), .B(n15751), .Z(n15759) );
  XNOR U16183 ( .A(n15758), .B(n15759), .Z(n15760) );
  XNOR U16184 ( .A(n15761), .B(n15760), .Z(n15794) );
  XNOR U16185 ( .A(n15794), .B(sreg[1398]), .Z(n15796) );
  NAND U16186 ( .A(n15753), .B(sreg[1397]), .Z(n15757) );
  OR U16187 ( .A(n15755), .B(n15754), .Z(n15756) );
  AND U16188 ( .A(n15757), .B(n15756), .Z(n15795) );
  XOR U16189 ( .A(n15796), .B(n15795), .Z(c[1398]) );
  NANDN U16190 ( .A(n15759), .B(n15758), .Z(n15763) );
  NAND U16191 ( .A(n15761), .B(n15760), .Z(n15762) );
  NAND U16192 ( .A(n15763), .B(n15762), .Z(n15802) );
  NAND U16193 ( .A(b[0]), .B(a[383]), .Z(n15764) );
  XNOR U16194 ( .A(b[1]), .B(n15764), .Z(n15766) );
  NAND U16195 ( .A(n69), .B(a[382]), .Z(n15765) );
  AND U16196 ( .A(n15766), .B(n15765), .Z(n15819) );
  XOR U16197 ( .A(a[379]), .B(n42197), .Z(n15808) );
  NANDN U16198 ( .A(n15808), .B(n42173), .Z(n15769) );
  NANDN U16199 ( .A(n15767), .B(n42172), .Z(n15768) );
  NAND U16200 ( .A(n15769), .B(n15768), .Z(n15817) );
  NAND U16201 ( .A(b[7]), .B(a[375]), .Z(n15818) );
  XNOR U16202 ( .A(n15817), .B(n15818), .Z(n15820) );
  XOR U16203 ( .A(n15819), .B(n15820), .Z(n15826) );
  NANDN U16204 ( .A(n15770), .B(n42093), .Z(n15772) );
  XOR U16205 ( .A(n42134), .B(a[381]), .Z(n15811) );
  NANDN U16206 ( .A(n15811), .B(n42095), .Z(n15771) );
  NAND U16207 ( .A(n15772), .B(n15771), .Z(n15824) );
  NANDN U16208 ( .A(n15773), .B(n42231), .Z(n15775) );
  XOR U16209 ( .A(n193), .B(a[377]), .Z(n15814) );
  NANDN U16210 ( .A(n15814), .B(n42234), .Z(n15774) );
  AND U16211 ( .A(n15775), .B(n15774), .Z(n15823) );
  XNOR U16212 ( .A(n15824), .B(n15823), .Z(n15825) );
  XNOR U16213 ( .A(n15826), .B(n15825), .Z(n15830) );
  NANDN U16214 ( .A(n15777), .B(n15776), .Z(n15781) );
  NAND U16215 ( .A(n15779), .B(n15778), .Z(n15780) );
  AND U16216 ( .A(n15781), .B(n15780), .Z(n15829) );
  XOR U16217 ( .A(n15830), .B(n15829), .Z(n15831) );
  NANDN U16218 ( .A(n15783), .B(n15782), .Z(n15787) );
  NANDN U16219 ( .A(n15785), .B(n15784), .Z(n15786) );
  NAND U16220 ( .A(n15787), .B(n15786), .Z(n15832) );
  XOR U16221 ( .A(n15831), .B(n15832), .Z(n15799) );
  OR U16222 ( .A(n15789), .B(n15788), .Z(n15793) );
  NANDN U16223 ( .A(n15791), .B(n15790), .Z(n15792) );
  NAND U16224 ( .A(n15793), .B(n15792), .Z(n15800) );
  XNOR U16225 ( .A(n15799), .B(n15800), .Z(n15801) );
  XNOR U16226 ( .A(n15802), .B(n15801), .Z(n15835) );
  XNOR U16227 ( .A(n15835), .B(sreg[1399]), .Z(n15837) );
  NAND U16228 ( .A(n15794), .B(sreg[1398]), .Z(n15798) );
  OR U16229 ( .A(n15796), .B(n15795), .Z(n15797) );
  AND U16230 ( .A(n15798), .B(n15797), .Z(n15836) );
  XOR U16231 ( .A(n15837), .B(n15836), .Z(c[1399]) );
  NANDN U16232 ( .A(n15800), .B(n15799), .Z(n15804) );
  NAND U16233 ( .A(n15802), .B(n15801), .Z(n15803) );
  NAND U16234 ( .A(n15804), .B(n15803), .Z(n15843) );
  NAND U16235 ( .A(b[0]), .B(a[384]), .Z(n15805) );
  XNOR U16236 ( .A(b[1]), .B(n15805), .Z(n15807) );
  NAND U16237 ( .A(n69), .B(a[383]), .Z(n15806) );
  AND U16238 ( .A(n15807), .B(n15806), .Z(n15860) );
  XOR U16239 ( .A(a[380]), .B(n42197), .Z(n15849) );
  NANDN U16240 ( .A(n15849), .B(n42173), .Z(n15810) );
  NANDN U16241 ( .A(n15808), .B(n42172), .Z(n15809) );
  NAND U16242 ( .A(n15810), .B(n15809), .Z(n15858) );
  NAND U16243 ( .A(b[7]), .B(a[376]), .Z(n15859) );
  XNOR U16244 ( .A(n15858), .B(n15859), .Z(n15861) );
  XOR U16245 ( .A(n15860), .B(n15861), .Z(n15867) );
  NANDN U16246 ( .A(n15811), .B(n42093), .Z(n15813) );
  XOR U16247 ( .A(n42134), .B(a[382]), .Z(n15852) );
  NANDN U16248 ( .A(n15852), .B(n42095), .Z(n15812) );
  NAND U16249 ( .A(n15813), .B(n15812), .Z(n15865) );
  NANDN U16250 ( .A(n15814), .B(n42231), .Z(n15816) );
  XOR U16251 ( .A(n193), .B(a[378]), .Z(n15855) );
  NANDN U16252 ( .A(n15855), .B(n42234), .Z(n15815) );
  AND U16253 ( .A(n15816), .B(n15815), .Z(n15864) );
  XNOR U16254 ( .A(n15865), .B(n15864), .Z(n15866) );
  XNOR U16255 ( .A(n15867), .B(n15866), .Z(n15871) );
  NANDN U16256 ( .A(n15818), .B(n15817), .Z(n15822) );
  NAND U16257 ( .A(n15820), .B(n15819), .Z(n15821) );
  AND U16258 ( .A(n15822), .B(n15821), .Z(n15870) );
  XOR U16259 ( .A(n15871), .B(n15870), .Z(n15872) );
  NANDN U16260 ( .A(n15824), .B(n15823), .Z(n15828) );
  NANDN U16261 ( .A(n15826), .B(n15825), .Z(n15827) );
  NAND U16262 ( .A(n15828), .B(n15827), .Z(n15873) );
  XOR U16263 ( .A(n15872), .B(n15873), .Z(n15840) );
  OR U16264 ( .A(n15830), .B(n15829), .Z(n15834) );
  NANDN U16265 ( .A(n15832), .B(n15831), .Z(n15833) );
  NAND U16266 ( .A(n15834), .B(n15833), .Z(n15841) );
  XNOR U16267 ( .A(n15840), .B(n15841), .Z(n15842) );
  XNOR U16268 ( .A(n15843), .B(n15842), .Z(n15876) );
  XNOR U16269 ( .A(n15876), .B(sreg[1400]), .Z(n15878) );
  NAND U16270 ( .A(n15835), .B(sreg[1399]), .Z(n15839) );
  OR U16271 ( .A(n15837), .B(n15836), .Z(n15838) );
  AND U16272 ( .A(n15839), .B(n15838), .Z(n15877) );
  XOR U16273 ( .A(n15878), .B(n15877), .Z(c[1400]) );
  NANDN U16274 ( .A(n15841), .B(n15840), .Z(n15845) );
  NAND U16275 ( .A(n15843), .B(n15842), .Z(n15844) );
  NAND U16276 ( .A(n15845), .B(n15844), .Z(n15884) );
  NAND U16277 ( .A(b[0]), .B(a[385]), .Z(n15846) );
  XNOR U16278 ( .A(b[1]), .B(n15846), .Z(n15848) );
  NAND U16279 ( .A(n70), .B(a[384]), .Z(n15847) );
  AND U16280 ( .A(n15848), .B(n15847), .Z(n15901) );
  XOR U16281 ( .A(a[381]), .B(n42197), .Z(n15890) );
  NANDN U16282 ( .A(n15890), .B(n42173), .Z(n15851) );
  NANDN U16283 ( .A(n15849), .B(n42172), .Z(n15850) );
  NAND U16284 ( .A(n15851), .B(n15850), .Z(n15899) );
  NAND U16285 ( .A(b[7]), .B(a[377]), .Z(n15900) );
  XNOR U16286 ( .A(n15899), .B(n15900), .Z(n15902) );
  XOR U16287 ( .A(n15901), .B(n15902), .Z(n15908) );
  NANDN U16288 ( .A(n15852), .B(n42093), .Z(n15854) );
  XOR U16289 ( .A(n42134), .B(a[383]), .Z(n15893) );
  NANDN U16290 ( .A(n15893), .B(n42095), .Z(n15853) );
  NAND U16291 ( .A(n15854), .B(n15853), .Z(n15906) );
  NANDN U16292 ( .A(n15855), .B(n42231), .Z(n15857) );
  XOR U16293 ( .A(n193), .B(a[379]), .Z(n15896) );
  NANDN U16294 ( .A(n15896), .B(n42234), .Z(n15856) );
  AND U16295 ( .A(n15857), .B(n15856), .Z(n15905) );
  XNOR U16296 ( .A(n15906), .B(n15905), .Z(n15907) );
  XNOR U16297 ( .A(n15908), .B(n15907), .Z(n15912) );
  NANDN U16298 ( .A(n15859), .B(n15858), .Z(n15863) );
  NAND U16299 ( .A(n15861), .B(n15860), .Z(n15862) );
  AND U16300 ( .A(n15863), .B(n15862), .Z(n15911) );
  XOR U16301 ( .A(n15912), .B(n15911), .Z(n15913) );
  NANDN U16302 ( .A(n15865), .B(n15864), .Z(n15869) );
  NANDN U16303 ( .A(n15867), .B(n15866), .Z(n15868) );
  NAND U16304 ( .A(n15869), .B(n15868), .Z(n15914) );
  XOR U16305 ( .A(n15913), .B(n15914), .Z(n15881) );
  OR U16306 ( .A(n15871), .B(n15870), .Z(n15875) );
  NANDN U16307 ( .A(n15873), .B(n15872), .Z(n15874) );
  NAND U16308 ( .A(n15875), .B(n15874), .Z(n15882) );
  XNOR U16309 ( .A(n15881), .B(n15882), .Z(n15883) );
  XNOR U16310 ( .A(n15884), .B(n15883), .Z(n15917) );
  XNOR U16311 ( .A(n15917), .B(sreg[1401]), .Z(n15919) );
  NAND U16312 ( .A(n15876), .B(sreg[1400]), .Z(n15880) );
  OR U16313 ( .A(n15878), .B(n15877), .Z(n15879) );
  AND U16314 ( .A(n15880), .B(n15879), .Z(n15918) );
  XOR U16315 ( .A(n15919), .B(n15918), .Z(c[1401]) );
  NANDN U16316 ( .A(n15882), .B(n15881), .Z(n15886) );
  NAND U16317 ( .A(n15884), .B(n15883), .Z(n15885) );
  NAND U16318 ( .A(n15886), .B(n15885), .Z(n15925) );
  NAND U16319 ( .A(b[0]), .B(a[386]), .Z(n15887) );
  XNOR U16320 ( .A(b[1]), .B(n15887), .Z(n15889) );
  NAND U16321 ( .A(n70), .B(a[385]), .Z(n15888) );
  AND U16322 ( .A(n15889), .B(n15888), .Z(n15942) );
  XOR U16323 ( .A(a[382]), .B(n42197), .Z(n15931) );
  NANDN U16324 ( .A(n15931), .B(n42173), .Z(n15892) );
  NANDN U16325 ( .A(n15890), .B(n42172), .Z(n15891) );
  NAND U16326 ( .A(n15892), .B(n15891), .Z(n15940) );
  NAND U16327 ( .A(b[7]), .B(a[378]), .Z(n15941) );
  XNOR U16328 ( .A(n15940), .B(n15941), .Z(n15943) );
  XOR U16329 ( .A(n15942), .B(n15943), .Z(n15949) );
  NANDN U16330 ( .A(n15893), .B(n42093), .Z(n15895) );
  XOR U16331 ( .A(n42134), .B(a[384]), .Z(n15934) );
  NANDN U16332 ( .A(n15934), .B(n42095), .Z(n15894) );
  NAND U16333 ( .A(n15895), .B(n15894), .Z(n15947) );
  NANDN U16334 ( .A(n15896), .B(n42231), .Z(n15898) );
  XOR U16335 ( .A(n193), .B(a[380]), .Z(n15937) );
  NANDN U16336 ( .A(n15937), .B(n42234), .Z(n15897) );
  AND U16337 ( .A(n15898), .B(n15897), .Z(n15946) );
  XNOR U16338 ( .A(n15947), .B(n15946), .Z(n15948) );
  XNOR U16339 ( .A(n15949), .B(n15948), .Z(n15953) );
  NANDN U16340 ( .A(n15900), .B(n15899), .Z(n15904) );
  NAND U16341 ( .A(n15902), .B(n15901), .Z(n15903) );
  AND U16342 ( .A(n15904), .B(n15903), .Z(n15952) );
  XOR U16343 ( .A(n15953), .B(n15952), .Z(n15954) );
  NANDN U16344 ( .A(n15906), .B(n15905), .Z(n15910) );
  NANDN U16345 ( .A(n15908), .B(n15907), .Z(n15909) );
  NAND U16346 ( .A(n15910), .B(n15909), .Z(n15955) );
  XOR U16347 ( .A(n15954), .B(n15955), .Z(n15922) );
  OR U16348 ( .A(n15912), .B(n15911), .Z(n15916) );
  NANDN U16349 ( .A(n15914), .B(n15913), .Z(n15915) );
  NAND U16350 ( .A(n15916), .B(n15915), .Z(n15923) );
  XNOR U16351 ( .A(n15922), .B(n15923), .Z(n15924) );
  XNOR U16352 ( .A(n15925), .B(n15924), .Z(n15958) );
  XNOR U16353 ( .A(n15958), .B(sreg[1402]), .Z(n15960) );
  NAND U16354 ( .A(n15917), .B(sreg[1401]), .Z(n15921) );
  OR U16355 ( .A(n15919), .B(n15918), .Z(n15920) );
  AND U16356 ( .A(n15921), .B(n15920), .Z(n15959) );
  XOR U16357 ( .A(n15960), .B(n15959), .Z(c[1402]) );
  NANDN U16358 ( .A(n15923), .B(n15922), .Z(n15927) );
  NAND U16359 ( .A(n15925), .B(n15924), .Z(n15926) );
  NAND U16360 ( .A(n15927), .B(n15926), .Z(n15966) );
  NAND U16361 ( .A(b[0]), .B(a[387]), .Z(n15928) );
  XNOR U16362 ( .A(b[1]), .B(n15928), .Z(n15930) );
  NAND U16363 ( .A(n70), .B(a[386]), .Z(n15929) );
  AND U16364 ( .A(n15930), .B(n15929), .Z(n15983) );
  XOR U16365 ( .A(a[383]), .B(n42197), .Z(n15972) );
  NANDN U16366 ( .A(n15972), .B(n42173), .Z(n15933) );
  NANDN U16367 ( .A(n15931), .B(n42172), .Z(n15932) );
  NAND U16368 ( .A(n15933), .B(n15932), .Z(n15981) );
  NAND U16369 ( .A(b[7]), .B(a[379]), .Z(n15982) );
  XNOR U16370 ( .A(n15981), .B(n15982), .Z(n15984) );
  XOR U16371 ( .A(n15983), .B(n15984), .Z(n15990) );
  NANDN U16372 ( .A(n15934), .B(n42093), .Z(n15936) );
  XOR U16373 ( .A(n42134), .B(a[385]), .Z(n15975) );
  NANDN U16374 ( .A(n15975), .B(n42095), .Z(n15935) );
  NAND U16375 ( .A(n15936), .B(n15935), .Z(n15988) );
  NANDN U16376 ( .A(n15937), .B(n42231), .Z(n15939) );
  XOR U16377 ( .A(n193), .B(a[381]), .Z(n15978) );
  NANDN U16378 ( .A(n15978), .B(n42234), .Z(n15938) );
  AND U16379 ( .A(n15939), .B(n15938), .Z(n15987) );
  XNOR U16380 ( .A(n15988), .B(n15987), .Z(n15989) );
  XNOR U16381 ( .A(n15990), .B(n15989), .Z(n15994) );
  NANDN U16382 ( .A(n15941), .B(n15940), .Z(n15945) );
  NAND U16383 ( .A(n15943), .B(n15942), .Z(n15944) );
  AND U16384 ( .A(n15945), .B(n15944), .Z(n15993) );
  XOR U16385 ( .A(n15994), .B(n15993), .Z(n15995) );
  NANDN U16386 ( .A(n15947), .B(n15946), .Z(n15951) );
  NANDN U16387 ( .A(n15949), .B(n15948), .Z(n15950) );
  NAND U16388 ( .A(n15951), .B(n15950), .Z(n15996) );
  XOR U16389 ( .A(n15995), .B(n15996), .Z(n15963) );
  OR U16390 ( .A(n15953), .B(n15952), .Z(n15957) );
  NANDN U16391 ( .A(n15955), .B(n15954), .Z(n15956) );
  NAND U16392 ( .A(n15957), .B(n15956), .Z(n15964) );
  XNOR U16393 ( .A(n15963), .B(n15964), .Z(n15965) );
  XNOR U16394 ( .A(n15966), .B(n15965), .Z(n15999) );
  XNOR U16395 ( .A(n15999), .B(sreg[1403]), .Z(n16001) );
  NAND U16396 ( .A(n15958), .B(sreg[1402]), .Z(n15962) );
  OR U16397 ( .A(n15960), .B(n15959), .Z(n15961) );
  AND U16398 ( .A(n15962), .B(n15961), .Z(n16000) );
  XOR U16399 ( .A(n16001), .B(n16000), .Z(c[1403]) );
  NANDN U16400 ( .A(n15964), .B(n15963), .Z(n15968) );
  NAND U16401 ( .A(n15966), .B(n15965), .Z(n15967) );
  NAND U16402 ( .A(n15968), .B(n15967), .Z(n16007) );
  NAND U16403 ( .A(b[0]), .B(a[388]), .Z(n15969) );
  XNOR U16404 ( .A(b[1]), .B(n15969), .Z(n15971) );
  NAND U16405 ( .A(n70), .B(a[387]), .Z(n15970) );
  AND U16406 ( .A(n15971), .B(n15970), .Z(n16024) );
  XOR U16407 ( .A(a[384]), .B(n42197), .Z(n16013) );
  NANDN U16408 ( .A(n16013), .B(n42173), .Z(n15974) );
  NANDN U16409 ( .A(n15972), .B(n42172), .Z(n15973) );
  NAND U16410 ( .A(n15974), .B(n15973), .Z(n16022) );
  NAND U16411 ( .A(b[7]), .B(a[380]), .Z(n16023) );
  XNOR U16412 ( .A(n16022), .B(n16023), .Z(n16025) );
  XOR U16413 ( .A(n16024), .B(n16025), .Z(n16031) );
  NANDN U16414 ( .A(n15975), .B(n42093), .Z(n15977) );
  XOR U16415 ( .A(n42134), .B(a[386]), .Z(n16016) );
  NANDN U16416 ( .A(n16016), .B(n42095), .Z(n15976) );
  NAND U16417 ( .A(n15977), .B(n15976), .Z(n16029) );
  NANDN U16418 ( .A(n15978), .B(n42231), .Z(n15980) );
  XOR U16419 ( .A(n193), .B(a[382]), .Z(n16019) );
  NANDN U16420 ( .A(n16019), .B(n42234), .Z(n15979) );
  AND U16421 ( .A(n15980), .B(n15979), .Z(n16028) );
  XNOR U16422 ( .A(n16029), .B(n16028), .Z(n16030) );
  XNOR U16423 ( .A(n16031), .B(n16030), .Z(n16035) );
  NANDN U16424 ( .A(n15982), .B(n15981), .Z(n15986) );
  NAND U16425 ( .A(n15984), .B(n15983), .Z(n15985) );
  AND U16426 ( .A(n15986), .B(n15985), .Z(n16034) );
  XOR U16427 ( .A(n16035), .B(n16034), .Z(n16036) );
  NANDN U16428 ( .A(n15988), .B(n15987), .Z(n15992) );
  NANDN U16429 ( .A(n15990), .B(n15989), .Z(n15991) );
  NAND U16430 ( .A(n15992), .B(n15991), .Z(n16037) );
  XOR U16431 ( .A(n16036), .B(n16037), .Z(n16004) );
  OR U16432 ( .A(n15994), .B(n15993), .Z(n15998) );
  NANDN U16433 ( .A(n15996), .B(n15995), .Z(n15997) );
  NAND U16434 ( .A(n15998), .B(n15997), .Z(n16005) );
  XNOR U16435 ( .A(n16004), .B(n16005), .Z(n16006) );
  XNOR U16436 ( .A(n16007), .B(n16006), .Z(n16040) );
  XNOR U16437 ( .A(n16040), .B(sreg[1404]), .Z(n16042) );
  NAND U16438 ( .A(n15999), .B(sreg[1403]), .Z(n16003) );
  OR U16439 ( .A(n16001), .B(n16000), .Z(n16002) );
  AND U16440 ( .A(n16003), .B(n16002), .Z(n16041) );
  XOR U16441 ( .A(n16042), .B(n16041), .Z(c[1404]) );
  NANDN U16442 ( .A(n16005), .B(n16004), .Z(n16009) );
  NAND U16443 ( .A(n16007), .B(n16006), .Z(n16008) );
  NAND U16444 ( .A(n16009), .B(n16008), .Z(n16048) );
  NAND U16445 ( .A(b[0]), .B(a[389]), .Z(n16010) );
  XNOR U16446 ( .A(b[1]), .B(n16010), .Z(n16012) );
  NAND U16447 ( .A(n70), .B(a[388]), .Z(n16011) );
  AND U16448 ( .A(n16012), .B(n16011), .Z(n16065) );
  XOR U16449 ( .A(a[385]), .B(n42197), .Z(n16054) );
  NANDN U16450 ( .A(n16054), .B(n42173), .Z(n16015) );
  NANDN U16451 ( .A(n16013), .B(n42172), .Z(n16014) );
  NAND U16452 ( .A(n16015), .B(n16014), .Z(n16063) );
  NAND U16453 ( .A(b[7]), .B(a[381]), .Z(n16064) );
  XNOR U16454 ( .A(n16063), .B(n16064), .Z(n16066) );
  XOR U16455 ( .A(n16065), .B(n16066), .Z(n16072) );
  NANDN U16456 ( .A(n16016), .B(n42093), .Z(n16018) );
  XOR U16457 ( .A(n42134), .B(a[387]), .Z(n16057) );
  NANDN U16458 ( .A(n16057), .B(n42095), .Z(n16017) );
  NAND U16459 ( .A(n16018), .B(n16017), .Z(n16070) );
  NANDN U16460 ( .A(n16019), .B(n42231), .Z(n16021) );
  XOR U16461 ( .A(n194), .B(a[383]), .Z(n16060) );
  NANDN U16462 ( .A(n16060), .B(n42234), .Z(n16020) );
  AND U16463 ( .A(n16021), .B(n16020), .Z(n16069) );
  XNOR U16464 ( .A(n16070), .B(n16069), .Z(n16071) );
  XNOR U16465 ( .A(n16072), .B(n16071), .Z(n16076) );
  NANDN U16466 ( .A(n16023), .B(n16022), .Z(n16027) );
  NAND U16467 ( .A(n16025), .B(n16024), .Z(n16026) );
  AND U16468 ( .A(n16027), .B(n16026), .Z(n16075) );
  XOR U16469 ( .A(n16076), .B(n16075), .Z(n16077) );
  NANDN U16470 ( .A(n16029), .B(n16028), .Z(n16033) );
  NANDN U16471 ( .A(n16031), .B(n16030), .Z(n16032) );
  NAND U16472 ( .A(n16033), .B(n16032), .Z(n16078) );
  XOR U16473 ( .A(n16077), .B(n16078), .Z(n16045) );
  OR U16474 ( .A(n16035), .B(n16034), .Z(n16039) );
  NANDN U16475 ( .A(n16037), .B(n16036), .Z(n16038) );
  NAND U16476 ( .A(n16039), .B(n16038), .Z(n16046) );
  XNOR U16477 ( .A(n16045), .B(n16046), .Z(n16047) );
  XNOR U16478 ( .A(n16048), .B(n16047), .Z(n16081) );
  XNOR U16479 ( .A(n16081), .B(sreg[1405]), .Z(n16083) );
  NAND U16480 ( .A(n16040), .B(sreg[1404]), .Z(n16044) );
  OR U16481 ( .A(n16042), .B(n16041), .Z(n16043) );
  AND U16482 ( .A(n16044), .B(n16043), .Z(n16082) );
  XOR U16483 ( .A(n16083), .B(n16082), .Z(c[1405]) );
  NANDN U16484 ( .A(n16046), .B(n16045), .Z(n16050) );
  NAND U16485 ( .A(n16048), .B(n16047), .Z(n16049) );
  NAND U16486 ( .A(n16050), .B(n16049), .Z(n16089) );
  NAND U16487 ( .A(b[0]), .B(a[390]), .Z(n16051) );
  XNOR U16488 ( .A(b[1]), .B(n16051), .Z(n16053) );
  NAND U16489 ( .A(n70), .B(a[389]), .Z(n16052) );
  AND U16490 ( .A(n16053), .B(n16052), .Z(n16106) );
  XOR U16491 ( .A(a[386]), .B(n42197), .Z(n16095) );
  NANDN U16492 ( .A(n16095), .B(n42173), .Z(n16056) );
  NANDN U16493 ( .A(n16054), .B(n42172), .Z(n16055) );
  NAND U16494 ( .A(n16056), .B(n16055), .Z(n16104) );
  NAND U16495 ( .A(b[7]), .B(a[382]), .Z(n16105) );
  XNOR U16496 ( .A(n16104), .B(n16105), .Z(n16107) );
  XOR U16497 ( .A(n16106), .B(n16107), .Z(n16113) );
  NANDN U16498 ( .A(n16057), .B(n42093), .Z(n16059) );
  XOR U16499 ( .A(n42134), .B(a[388]), .Z(n16098) );
  NANDN U16500 ( .A(n16098), .B(n42095), .Z(n16058) );
  NAND U16501 ( .A(n16059), .B(n16058), .Z(n16111) );
  NANDN U16502 ( .A(n16060), .B(n42231), .Z(n16062) );
  XOR U16503 ( .A(n194), .B(a[384]), .Z(n16101) );
  NANDN U16504 ( .A(n16101), .B(n42234), .Z(n16061) );
  AND U16505 ( .A(n16062), .B(n16061), .Z(n16110) );
  XNOR U16506 ( .A(n16111), .B(n16110), .Z(n16112) );
  XNOR U16507 ( .A(n16113), .B(n16112), .Z(n16117) );
  NANDN U16508 ( .A(n16064), .B(n16063), .Z(n16068) );
  NAND U16509 ( .A(n16066), .B(n16065), .Z(n16067) );
  AND U16510 ( .A(n16068), .B(n16067), .Z(n16116) );
  XOR U16511 ( .A(n16117), .B(n16116), .Z(n16118) );
  NANDN U16512 ( .A(n16070), .B(n16069), .Z(n16074) );
  NANDN U16513 ( .A(n16072), .B(n16071), .Z(n16073) );
  NAND U16514 ( .A(n16074), .B(n16073), .Z(n16119) );
  XOR U16515 ( .A(n16118), .B(n16119), .Z(n16086) );
  OR U16516 ( .A(n16076), .B(n16075), .Z(n16080) );
  NANDN U16517 ( .A(n16078), .B(n16077), .Z(n16079) );
  NAND U16518 ( .A(n16080), .B(n16079), .Z(n16087) );
  XNOR U16519 ( .A(n16086), .B(n16087), .Z(n16088) );
  XNOR U16520 ( .A(n16089), .B(n16088), .Z(n16122) );
  XNOR U16521 ( .A(n16122), .B(sreg[1406]), .Z(n16124) );
  NAND U16522 ( .A(n16081), .B(sreg[1405]), .Z(n16085) );
  OR U16523 ( .A(n16083), .B(n16082), .Z(n16084) );
  AND U16524 ( .A(n16085), .B(n16084), .Z(n16123) );
  XOR U16525 ( .A(n16124), .B(n16123), .Z(c[1406]) );
  NANDN U16526 ( .A(n16087), .B(n16086), .Z(n16091) );
  NAND U16527 ( .A(n16089), .B(n16088), .Z(n16090) );
  NAND U16528 ( .A(n16091), .B(n16090), .Z(n16130) );
  NAND U16529 ( .A(b[0]), .B(a[391]), .Z(n16092) );
  XNOR U16530 ( .A(b[1]), .B(n16092), .Z(n16094) );
  NAND U16531 ( .A(n70), .B(a[390]), .Z(n16093) );
  AND U16532 ( .A(n16094), .B(n16093), .Z(n16147) );
  XOR U16533 ( .A(a[387]), .B(n42197), .Z(n16136) );
  NANDN U16534 ( .A(n16136), .B(n42173), .Z(n16097) );
  NANDN U16535 ( .A(n16095), .B(n42172), .Z(n16096) );
  NAND U16536 ( .A(n16097), .B(n16096), .Z(n16145) );
  NAND U16537 ( .A(b[7]), .B(a[383]), .Z(n16146) );
  XNOR U16538 ( .A(n16145), .B(n16146), .Z(n16148) );
  XOR U16539 ( .A(n16147), .B(n16148), .Z(n16154) );
  NANDN U16540 ( .A(n16098), .B(n42093), .Z(n16100) );
  XOR U16541 ( .A(n42134), .B(a[389]), .Z(n16139) );
  NANDN U16542 ( .A(n16139), .B(n42095), .Z(n16099) );
  NAND U16543 ( .A(n16100), .B(n16099), .Z(n16152) );
  NANDN U16544 ( .A(n16101), .B(n42231), .Z(n16103) );
  XOR U16545 ( .A(n194), .B(a[385]), .Z(n16142) );
  NANDN U16546 ( .A(n16142), .B(n42234), .Z(n16102) );
  AND U16547 ( .A(n16103), .B(n16102), .Z(n16151) );
  XNOR U16548 ( .A(n16152), .B(n16151), .Z(n16153) );
  XNOR U16549 ( .A(n16154), .B(n16153), .Z(n16158) );
  NANDN U16550 ( .A(n16105), .B(n16104), .Z(n16109) );
  NAND U16551 ( .A(n16107), .B(n16106), .Z(n16108) );
  AND U16552 ( .A(n16109), .B(n16108), .Z(n16157) );
  XOR U16553 ( .A(n16158), .B(n16157), .Z(n16159) );
  NANDN U16554 ( .A(n16111), .B(n16110), .Z(n16115) );
  NANDN U16555 ( .A(n16113), .B(n16112), .Z(n16114) );
  NAND U16556 ( .A(n16115), .B(n16114), .Z(n16160) );
  XOR U16557 ( .A(n16159), .B(n16160), .Z(n16127) );
  OR U16558 ( .A(n16117), .B(n16116), .Z(n16121) );
  NANDN U16559 ( .A(n16119), .B(n16118), .Z(n16120) );
  NAND U16560 ( .A(n16121), .B(n16120), .Z(n16128) );
  XNOR U16561 ( .A(n16127), .B(n16128), .Z(n16129) );
  XNOR U16562 ( .A(n16130), .B(n16129), .Z(n16163) );
  XNOR U16563 ( .A(n16163), .B(sreg[1407]), .Z(n16165) );
  NAND U16564 ( .A(n16122), .B(sreg[1406]), .Z(n16126) );
  OR U16565 ( .A(n16124), .B(n16123), .Z(n16125) );
  AND U16566 ( .A(n16126), .B(n16125), .Z(n16164) );
  XOR U16567 ( .A(n16165), .B(n16164), .Z(c[1407]) );
  NANDN U16568 ( .A(n16128), .B(n16127), .Z(n16132) );
  NAND U16569 ( .A(n16130), .B(n16129), .Z(n16131) );
  NAND U16570 ( .A(n16132), .B(n16131), .Z(n16171) );
  NAND U16571 ( .A(b[0]), .B(a[392]), .Z(n16133) );
  XNOR U16572 ( .A(b[1]), .B(n16133), .Z(n16135) );
  NAND U16573 ( .A(n71), .B(a[391]), .Z(n16134) );
  AND U16574 ( .A(n16135), .B(n16134), .Z(n16188) );
  XOR U16575 ( .A(a[388]), .B(n42197), .Z(n16177) );
  NANDN U16576 ( .A(n16177), .B(n42173), .Z(n16138) );
  NANDN U16577 ( .A(n16136), .B(n42172), .Z(n16137) );
  NAND U16578 ( .A(n16138), .B(n16137), .Z(n16186) );
  NAND U16579 ( .A(b[7]), .B(a[384]), .Z(n16187) );
  XNOR U16580 ( .A(n16186), .B(n16187), .Z(n16189) );
  XOR U16581 ( .A(n16188), .B(n16189), .Z(n16195) );
  NANDN U16582 ( .A(n16139), .B(n42093), .Z(n16141) );
  XOR U16583 ( .A(n42134), .B(a[390]), .Z(n16180) );
  NANDN U16584 ( .A(n16180), .B(n42095), .Z(n16140) );
  NAND U16585 ( .A(n16141), .B(n16140), .Z(n16193) );
  NANDN U16586 ( .A(n16142), .B(n42231), .Z(n16144) );
  XOR U16587 ( .A(n194), .B(a[386]), .Z(n16183) );
  NANDN U16588 ( .A(n16183), .B(n42234), .Z(n16143) );
  AND U16589 ( .A(n16144), .B(n16143), .Z(n16192) );
  XNOR U16590 ( .A(n16193), .B(n16192), .Z(n16194) );
  XNOR U16591 ( .A(n16195), .B(n16194), .Z(n16199) );
  NANDN U16592 ( .A(n16146), .B(n16145), .Z(n16150) );
  NAND U16593 ( .A(n16148), .B(n16147), .Z(n16149) );
  AND U16594 ( .A(n16150), .B(n16149), .Z(n16198) );
  XOR U16595 ( .A(n16199), .B(n16198), .Z(n16200) );
  NANDN U16596 ( .A(n16152), .B(n16151), .Z(n16156) );
  NANDN U16597 ( .A(n16154), .B(n16153), .Z(n16155) );
  NAND U16598 ( .A(n16156), .B(n16155), .Z(n16201) );
  XOR U16599 ( .A(n16200), .B(n16201), .Z(n16168) );
  OR U16600 ( .A(n16158), .B(n16157), .Z(n16162) );
  NANDN U16601 ( .A(n16160), .B(n16159), .Z(n16161) );
  NAND U16602 ( .A(n16162), .B(n16161), .Z(n16169) );
  XNOR U16603 ( .A(n16168), .B(n16169), .Z(n16170) );
  XNOR U16604 ( .A(n16171), .B(n16170), .Z(n16204) );
  XNOR U16605 ( .A(n16204), .B(sreg[1408]), .Z(n16206) );
  NAND U16606 ( .A(n16163), .B(sreg[1407]), .Z(n16167) );
  OR U16607 ( .A(n16165), .B(n16164), .Z(n16166) );
  AND U16608 ( .A(n16167), .B(n16166), .Z(n16205) );
  XOR U16609 ( .A(n16206), .B(n16205), .Z(c[1408]) );
  NANDN U16610 ( .A(n16169), .B(n16168), .Z(n16173) );
  NAND U16611 ( .A(n16171), .B(n16170), .Z(n16172) );
  NAND U16612 ( .A(n16173), .B(n16172), .Z(n16212) );
  NAND U16613 ( .A(b[0]), .B(a[393]), .Z(n16174) );
  XNOR U16614 ( .A(b[1]), .B(n16174), .Z(n16176) );
  NAND U16615 ( .A(n71), .B(a[392]), .Z(n16175) );
  AND U16616 ( .A(n16176), .B(n16175), .Z(n16229) );
  XOR U16617 ( .A(a[389]), .B(n42197), .Z(n16218) );
  NANDN U16618 ( .A(n16218), .B(n42173), .Z(n16179) );
  NANDN U16619 ( .A(n16177), .B(n42172), .Z(n16178) );
  NAND U16620 ( .A(n16179), .B(n16178), .Z(n16227) );
  NAND U16621 ( .A(b[7]), .B(a[385]), .Z(n16228) );
  XNOR U16622 ( .A(n16227), .B(n16228), .Z(n16230) );
  XOR U16623 ( .A(n16229), .B(n16230), .Z(n16236) );
  NANDN U16624 ( .A(n16180), .B(n42093), .Z(n16182) );
  XOR U16625 ( .A(n42134), .B(a[391]), .Z(n16221) );
  NANDN U16626 ( .A(n16221), .B(n42095), .Z(n16181) );
  NAND U16627 ( .A(n16182), .B(n16181), .Z(n16234) );
  NANDN U16628 ( .A(n16183), .B(n42231), .Z(n16185) );
  XOR U16629 ( .A(n194), .B(a[387]), .Z(n16224) );
  NANDN U16630 ( .A(n16224), .B(n42234), .Z(n16184) );
  AND U16631 ( .A(n16185), .B(n16184), .Z(n16233) );
  XNOR U16632 ( .A(n16234), .B(n16233), .Z(n16235) );
  XNOR U16633 ( .A(n16236), .B(n16235), .Z(n16240) );
  NANDN U16634 ( .A(n16187), .B(n16186), .Z(n16191) );
  NAND U16635 ( .A(n16189), .B(n16188), .Z(n16190) );
  AND U16636 ( .A(n16191), .B(n16190), .Z(n16239) );
  XOR U16637 ( .A(n16240), .B(n16239), .Z(n16241) );
  NANDN U16638 ( .A(n16193), .B(n16192), .Z(n16197) );
  NANDN U16639 ( .A(n16195), .B(n16194), .Z(n16196) );
  NAND U16640 ( .A(n16197), .B(n16196), .Z(n16242) );
  XOR U16641 ( .A(n16241), .B(n16242), .Z(n16209) );
  OR U16642 ( .A(n16199), .B(n16198), .Z(n16203) );
  NANDN U16643 ( .A(n16201), .B(n16200), .Z(n16202) );
  NAND U16644 ( .A(n16203), .B(n16202), .Z(n16210) );
  XNOR U16645 ( .A(n16209), .B(n16210), .Z(n16211) );
  XNOR U16646 ( .A(n16212), .B(n16211), .Z(n16245) );
  XNOR U16647 ( .A(n16245), .B(sreg[1409]), .Z(n16247) );
  NAND U16648 ( .A(n16204), .B(sreg[1408]), .Z(n16208) );
  OR U16649 ( .A(n16206), .B(n16205), .Z(n16207) );
  AND U16650 ( .A(n16208), .B(n16207), .Z(n16246) );
  XOR U16651 ( .A(n16247), .B(n16246), .Z(c[1409]) );
  NANDN U16652 ( .A(n16210), .B(n16209), .Z(n16214) );
  NAND U16653 ( .A(n16212), .B(n16211), .Z(n16213) );
  NAND U16654 ( .A(n16214), .B(n16213), .Z(n16253) );
  NAND U16655 ( .A(b[0]), .B(a[394]), .Z(n16215) );
  XNOR U16656 ( .A(b[1]), .B(n16215), .Z(n16217) );
  NAND U16657 ( .A(n71), .B(a[393]), .Z(n16216) );
  AND U16658 ( .A(n16217), .B(n16216), .Z(n16270) );
  XOR U16659 ( .A(a[390]), .B(n42197), .Z(n16259) );
  NANDN U16660 ( .A(n16259), .B(n42173), .Z(n16220) );
  NANDN U16661 ( .A(n16218), .B(n42172), .Z(n16219) );
  NAND U16662 ( .A(n16220), .B(n16219), .Z(n16268) );
  NAND U16663 ( .A(b[7]), .B(a[386]), .Z(n16269) );
  XNOR U16664 ( .A(n16268), .B(n16269), .Z(n16271) );
  XOR U16665 ( .A(n16270), .B(n16271), .Z(n16277) );
  NANDN U16666 ( .A(n16221), .B(n42093), .Z(n16223) );
  XOR U16667 ( .A(n42134), .B(a[392]), .Z(n16262) );
  NANDN U16668 ( .A(n16262), .B(n42095), .Z(n16222) );
  NAND U16669 ( .A(n16223), .B(n16222), .Z(n16275) );
  NANDN U16670 ( .A(n16224), .B(n42231), .Z(n16226) );
  XOR U16671 ( .A(n194), .B(a[388]), .Z(n16265) );
  NANDN U16672 ( .A(n16265), .B(n42234), .Z(n16225) );
  AND U16673 ( .A(n16226), .B(n16225), .Z(n16274) );
  XNOR U16674 ( .A(n16275), .B(n16274), .Z(n16276) );
  XNOR U16675 ( .A(n16277), .B(n16276), .Z(n16281) );
  NANDN U16676 ( .A(n16228), .B(n16227), .Z(n16232) );
  NAND U16677 ( .A(n16230), .B(n16229), .Z(n16231) );
  AND U16678 ( .A(n16232), .B(n16231), .Z(n16280) );
  XOR U16679 ( .A(n16281), .B(n16280), .Z(n16282) );
  NANDN U16680 ( .A(n16234), .B(n16233), .Z(n16238) );
  NANDN U16681 ( .A(n16236), .B(n16235), .Z(n16237) );
  NAND U16682 ( .A(n16238), .B(n16237), .Z(n16283) );
  XOR U16683 ( .A(n16282), .B(n16283), .Z(n16250) );
  OR U16684 ( .A(n16240), .B(n16239), .Z(n16244) );
  NANDN U16685 ( .A(n16242), .B(n16241), .Z(n16243) );
  NAND U16686 ( .A(n16244), .B(n16243), .Z(n16251) );
  XNOR U16687 ( .A(n16250), .B(n16251), .Z(n16252) );
  XNOR U16688 ( .A(n16253), .B(n16252), .Z(n16286) );
  XNOR U16689 ( .A(n16286), .B(sreg[1410]), .Z(n16288) );
  NAND U16690 ( .A(n16245), .B(sreg[1409]), .Z(n16249) );
  OR U16691 ( .A(n16247), .B(n16246), .Z(n16248) );
  AND U16692 ( .A(n16249), .B(n16248), .Z(n16287) );
  XOR U16693 ( .A(n16288), .B(n16287), .Z(c[1410]) );
  NANDN U16694 ( .A(n16251), .B(n16250), .Z(n16255) );
  NAND U16695 ( .A(n16253), .B(n16252), .Z(n16254) );
  NAND U16696 ( .A(n16255), .B(n16254), .Z(n16294) );
  NAND U16697 ( .A(b[0]), .B(a[395]), .Z(n16256) );
  XNOR U16698 ( .A(b[1]), .B(n16256), .Z(n16258) );
  NAND U16699 ( .A(n71), .B(a[394]), .Z(n16257) );
  AND U16700 ( .A(n16258), .B(n16257), .Z(n16311) );
  XOR U16701 ( .A(a[391]), .B(n42197), .Z(n16300) );
  NANDN U16702 ( .A(n16300), .B(n42173), .Z(n16261) );
  NANDN U16703 ( .A(n16259), .B(n42172), .Z(n16260) );
  NAND U16704 ( .A(n16261), .B(n16260), .Z(n16309) );
  NAND U16705 ( .A(b[7]), .B(a[387]), .Z(n16310) );
  XNOR U16706 ( .A(n16309), .B(n16310), .Z(n16312) );
  XOR U16707 ( .A(n16311), .B(n16312), .Z(n16318) );
  NANDN U16708 ( .A(n16262), .B(n42093), .Z(n16264) );
  XOR U16709 ( .A(n42134), .B(a[393]), .Z(n16303) );
  NANDN U16710 ( .A(n16303), .B(n42095), .Z(n16263) );
  NAND U16711 ( .A(n16264), .B(n16263), .Z(n16316) );
  NANDN U16712 ( .A(n16265), .B(n42231), .Z(n16267) );
  XOR U16713 ( .A(n194), .B(a[389]), .Z(n16306) );
  NANDN U16714 ( .A(n16306), .B(n42234), .Z(n16266) );
  AND U16715 ( .A(n16267), .B(n16266), .Z(n16315) );
  XNOR U16716 ( .A(n16316), .B(n16315), .Z(n16317) );
  XNOR U16717 ( .A(n16318), .B(n16317), .Z(n16322) );
  NANDN U16718 ( .A(n16269), .B(n16268), .Z(n16273) );
  NAND U16719 ( .A(n16271), .B(n16270), .Z(n16272) );
  AND U16720 ( .A(n16273), .B(n16272), .Z(n16321) );
  XOR U16721 ( .A(n16322), .B(n16321), .Z(n16323) );
  NANDN U16722 ( .A(n16275), .B(n16274), .Z(n16279) );
  NANDN U16723 ( .A(n16277), .B(n16276), .Z(n16278) );
  NAND U16724 ( .A(n16279), .B(n16278), .Z(n16324) );
  XOR U16725 ( .A(n16323), .B(n16324), .Z(n16291) );
  OR U16726 ( .A(n16281), .B(n16280), .Z(n16285) );
  NANDN U16727 ( .A(n16283), .B(n16282), .Z(n16284) );
  NAND U16728 ( .A(n16285), .B(n16284), .Z(n16292) );
  XNOR U16729 ( .A(n16291), .B(n16292), .Z(n16293) );
  XNOR U16730 ( .A(n16294), .B(n16293), .Z(n16327) );
  XNOR U16731 ( .A(n16327), .B(sreg[1411]), .Z(n16329) );
  NAND U16732 ( .A(n16286), .B(sreg[1410]), .Z(n16290) );
  OR U16733 ( .A(n16288), .B(n16287), .Z(n16289) );
  AND U16734 ( .A(n16290), .B(n16289), .Z(n16328) );
  XOR U16735 ( .A(n16329), .B(n16328), .Z(c[1411]) );
  NANDN U16736 ( .A(n16292), .B(n16291), .Z(n16296) );
  NAND U16737 ( .A(n16294), .B(n16293), .Z(n16295) );
  NAND U16738 ( .A(n16296), .B(n16295), .Z(n16335) );
  NAND U16739 ( .A(b[0]), .B(a[396]), .Z(n16297) );
  XNOR U16740 ( .A(b[1]), .B(n16297), .Z(n16299) );
  NAND U16741 ( .A(n71), .B(a[395]), .Z(n16298) );
  AND U16742 ( .A(n16299), .B(n16298), .Z(n16352) );
  XOR U16743 ( .A(a[392]), .B(n42197), .Z(n16341) );
  NANDN U16744 ( .A(n16341), .B(n42173), .Z(n16302) );
  NANDN U16745 ( .A(n16300), .B(n42172), .Z(n16301) );
  NAND U16746 ( .A(n16302), .B(n16301), .Z(n16350) );
  NAND U16747 ( .A(b[7]), .B(a[388]), .Z(n16351) );
  XNOR U16748 ( .A(n16350), .B(n16351), .Z(n16353) );
  XOR U16749 ( .A(n16352), .B(n16353), .Z(n16359) );
  NANDN U16750 ( .A(n16303), .B(n42093), .Z(n16305) );
  XOR U16751 ( .A(n42134), .B(a[394]), .Z(n16344) );
  NANDN U16752 ( .A(n16344), .B(n42095), .Z(n16304) );
  NAND U16753 ( .A(n16305), .B(n16304), .Z(n16357) );
  NANDN U16754 ( .A(n16306), .B(n42231), .Z(n16308) );
  XOR U16755 ( .A(n194), .B(a[390]), .Z(n16347) );
  NANDN U16756 ( .A(n16347), .B(n42234), .Z(n16307) );
  AND U16757 ( .A(n16308), .B(n16307), .Z(n16356) );
  XNOR U16758 ( .A(n16357), .B(n16356), .Z(n16358) );
  XNOR U16759 ( .A(n16359), .B(n16358), .Z(n16363) );
  NANDN U16760 ( .A(n16310), .B(n16309), .Z(n16314) );
  NAND U16761 ( .A(n16312), .B(n16311), .Z(n16313) );
  AND U16762 ( .A(n16314), .B(n16313), .Z(n16362) );
  XOR U16763 ( .A(n16363), .B(n16362), .Z(n16364) );
  NANDN U16764 ( .A(n16316), .B(n16315), .Z(n16320) );
  NANDN U16765 ( .A(n16318), .B(n16317), .Z(n16319) );
  NAND U16766 ( .A(n16320), .B(n16319), .Z(n16365) );
  XOR U16767 ( .A(n16364), .B(n16365), .Z(n16332) );
  OR U16768 ( .A(n16322), .B(n16321), .Z(n16326) );
  NANDN U16769 ( .A(n16324), .B(n16323), .Z(n16325) );
  NAND U16770 ( .A(n16326), .B(n16325), .Z(n16333) );
  XNOR U16771 ( .A(n16332), .B(n16333), .Z(n16334) );
  XNOR U16772 ( .A(n16335), .B(n16334), .Z(n16368) );
  XNOR U16773 ( .A(n16368), .B(sreg[1412]), .Z(n16370) );
  NAND U16774 ( .A(n16327), .B(sreg[1411]), .Z(n16331) );
  OR U16775 ( .A(n16329), .B(n16328), .Z(n16330) );
  AND U16776 ( .A(n16331), .B(n16330), .Z(n16369) );
  XOR U16777 ( .A(n16370), .B(n16369), .Z(c[1412]) );
  NANDN U16778 ( .A(n16333), .B(n16332), .Z(n16337) );
  NAND U16779 ( .A(n16335), .B(n16334), .Z(n16336) );
  NAND U16780 ( .A(n16337), .B(n16336), .Z(n16376) );
  NAND U16781 ( .A(b[0]), .B(a[397]), .Z(n16338) );
  XNOR U16782 ( .A(b[1]), .B(n16338), .Z(n16340) );
  NAND U16783 ( .A(n71), .B(a[396]), .Z(n16339) );
  AND U16784 ( .A(n16340), .B(n16339), .Z(n16393) );
  XOR U16785 ( .A(a[393]), .B(n42197), .Z(n16382) );
  NANDN U16786 ( .A(n16382), .B(n42173), .Z(n16343) );
  NANDN U16787 ( .A(n16341), .B(n42172), .Z(n16342) );
  NAND U16788 ( .A(n16343), .B(n16342), .Z(n16391) );
  NAND U16789 ( .A(b[7]), .B(a[389]), .Z(n16392) );
  XNOR U16790 ( .A(n16391), .B(n16392), .Z(n16394) );
  XOR U16791 ( .A(n16393), .B(n16394), .Z(n16400) );
  NANDN U16792 ( .A(n16344), .B(n42093), .Z(n16346) );
  XOR U16793 ( .A(n42134), .B(a[395]), .Z(n16385) );
  NANDN U16794 ( .A(n16385), .B(n42095), .Z(n16345) );
  NAND U16795 ( .A(n16346), .B(n16345), .Z(n16398) );
  NANDN U16796 ( .A(n16347), .B(n42231), .Z(n16349) );
  XOR U16797 ( .A(n194), .B(a[391]), .Z(n16388) );
  NANDN U16798 ( .A(n16388), .B(n42234), .Z(n16348) );
  AND U16799 ( .A(n16349), .B(n16348), .Z(n16397) );
  XNOR U16800 ( .A(n16398), .B(n16397), .Z(n16399) );
  XNOR U16801 ( .A(n16400), .B(n16399), .Z(n16404) );
  NANDN U16802 ( .A(n16351), .B(n16350), .Z(n16355) );
  NAND U16803 ( .A(n16353), .B(n16352), .Z(n16354) );
  AND U16804 ( .A(n16355), .B(n16354), .Z(n16403) );
  XOR U16805 ( .A(n16404), .B(n16403), .Z(n16405) );
  NANDN U16806 ( .A(n16357), .B(n16356), .Z(n16361) );
  NANDN U16807 ( .A(n16359), .B(n16358), .Z(n16360) );
  NAND U16808 ( .A(n16361), .B(n16360), .Z(n16406) );
  XOR U16809 ( .A(n16405), .B(n16406), .Z(n16373) );
  OR U16810 ( .A(n16363), .B(n16362), .Z(n16367) );
  NANDN U16811 ( .A(n16365), .B(n16364), .Z(n16366) );
  NAND U16812 ( .A(n16367), .B(n16366), .Z(n16374) );
  XNOR U16813 ( .A(n16373), .B(n16374), .Z(n16375) );
  XNOR U16814 ( .A(n16376), .B(n16375), .Z(n16409) );
  XNOR U16815 ( .A(n16409), .B(sreg[1413]), .Z(n16411) );
  NAND U16816 ( .A(n16368), .B(sreg[1412]), .Z(n16372) );
  OR U16817 ( .A(n16370), .B(n16369), .Z(n16371) );
  AND U16818 ( .A(n16372), .B(n16371), .Z(n16410) );
  XOR U16819 ( .A(n16411), .B(n16410), .Z(c[1413]) );
  NANDN U16820 ( .A(n16374), .B(n16373), .Z(n16378) );
  NAND U16821 ( .A(n16376), .B(n16375), .Z(n16377) );
  NAND U16822 ( .A(n16378), .B(n16377), .Z(n16417) );
  NAND U16823 ( .A(b[0]), .B(a[398]), .Z(n16379) );
  XNOR U16824 ( .A(b[1]), .B(n16379), .Z(n16381) );
  NAND U16825 ( .A(n71), .B(a[397]), .Z(n16380) );
  AND U16826 ( .A(n16381), .B(n16380), .Z(n16434) );
  XOR U16827 ( .A(a[394]), .B(n42197), .Z(n16423) );
  NANDN U16828 ( .A(n16423), .B(n42173), .Z(n16384) );
  NANDN U16829 ( .A(n16382), .B(n42172), .Z(n16383) );
  NAND U16830 ( .A(n16384), .B(n16383), .Z(n16432) );
  NAND U16831 ( .A(b[7]), .B(a[390]), .Z(n16433) );
  XNOR U16832 ( .A(n16432), .B(n16433), .Z(n16435) );
  XOR U16833 ( .A(n16434), .B(n16435), .Z(n16441) );
  NANDN U16834 ( .A(n16385), .B(n42093), .Z(n16387) );
  XOR U16835 ( .A(n42134), .B(a[396]), .Z(n16426) );
  NANDN U16836 ( .A(n16426), .B(n42095), .Z(n16386) );
  NAND U16837 ( .A(n16387), .B(n16386), .Z(n16439) );
  NANDN U16838 ( .A(n16388), .B(n42231), .Z(n16390) );
  XOR U16839 ( .A(n194), .B(a[392]), .Z(n16429) );
  NANDN U16840 ( .A(n16429), .B(n42234), .Z(n16389) );
  AND U16841 ( .A(n16390), .B(n16389), .Z(n16438) );
  XNOR U16842 ( .A(n16439), .B(n16438), .Z(n16440) );
  XNOR U16843 ( .A(n16441), .B(n16440), .Z(n16445) );
  NANDN U16844 ( .A(n16392), .B(n16391), .Z(n16396) );
  NAND U16845 ( .A(n16394), .B(n16393), .Z(n16395) );
  AND U16846 ( .A(n16396), .B(n16395), .Z(n16444) );
  XOR U16847 ( .A(n16445), .B(n16444), .Z(n16446) );
  NANDN U16848 ( .A(n16398), .B(n16397), .Z(n16402) );
  NANDN U16849 ( .A(n16400), .B(n16399), .Z(n16401) );
  NAND U16850 ( .A(n16402), .B(n16401), .Z(n16447) );
  XOR U16851 ( .A(n16446), .B(n16447), .Z(n16414) );
  OR U16852 ( .A(n16404), .B(n16403), .Z(n16408) );
  NANDN U16853 ( .A(n16406), .B(n16405), .Z(n16407) );
  NAND U16854 ( .A(n16408), .B(n16407), .Z(n16415) );
  XNOR U16855 ( .A(n16414), .B(n16415), .Z(n16416) );
  XNOR U16856 ( .A(n16417), .B(n16416), .Z(n16450) );
  XNOR U16857 ( .A(n16450), .B(sreg[1414]), .Z(n16452) );
  NAND U16858 ( .A(n16409), .B(sreg[1413]), .Z(n16413) );
  OR U16859 ( .A(n16411), .B(n16410), .Z(n16412) );
  AND U16860 ( .A(n16413), .B(n16412), .Z(n16451) );
  XOR U16861 ( .A(n16452), .B(n16451), .Z(c[1414]) );
  NANDN U16862 ( .A(n16415), .B(n16414), .Z(n16419) );
  NAND U16863 ( .A(n16417), .B(n16416), .Z(n16418) );
  NAND U16864 ( .A(n16419), .B(n16418), .Z(n16458) );
  NAND U16865 ( .A(b[0]), .B(a[399]), .Z(n16420) );
  XNOR U16866 ( .A(b[1]), .B(n16420), .Z(n16422) );
  NAND U16867 ( .A(n72), .B(a[398]), .Z(n16421) );
  AND U16868 ( .A(n16422), .B(n16421), .Z(n16475) );
  XOR U16869 ( .A(a[395]), .B(n42197), .Z(n16464) );
  NANDN U16870 ( .A(n16464), .B(n42173), .Z(n16425) );
  NANDN U16871 ( .A(n16423), .B(n42172), .Z(n16424) );
  NAND U16872 ( .A(n16425), .B(n16424), .Z(n16473) );
  NAND U16873 ( .A(b[7]), .B(a[391]), .Z(n16474) );
  XNOR U16874 ( .A(n16473), .B(n16474), .Z(n16476) );
  XOR U16875 ( .A(n16475), .B(n16476), .Z(n16482) );
  NANDN U16876 ( .A(n16426), .B(n42093), .Z(n16428) );
  XOR U16877 ( .A(n42134), .B(a[397]), .Z(n16467) );
  NANDN U16878 ( .A(n16467), .B(n42095), .Z(n16427) );
  NAND U16879 ( .A(n16428), .B(n16427), .Z(n16480) );
  NANDN U16880 ( .A(n16429), .B(n42231), .Z(n16431) );
  XOR U16881 ( .A(n194), .B(a[393]), .Z(n16470) );
  NANDN U16882 ( .A(n16470), .B(n42234), .Z(n16430) );
  AND U16883 ( .A(n16431), .B(n16430), .Z(n16479) );
  XNOR U16884 ( .A(n16480), .B(n16479), .Z(n16481) );
  XNOR U16885 ( .A(n16482), .B(n16481), .Z(n16486) );
  NANDN U16886 ( .A(n16433), .B(n16432), .Z(n16437) );
  NAND U16887 ( .A(n16435), .B(n16434), .Z(n16436) );
  AND U16888 ( .A(n16437), .B(n16436), .Z(n16485) );
  XOR U16889 ( .A(n16486), .B(n16485), .Z(n16487) );
  NANDN U16890 ( .A(n16439), .B(n16438), .Z(n16443) );
  NANDN U16891 ( .A(n16441), .B(n16440), .Z(n16442) );
  NAND U16892 ( .A(n16443), .B(n16442), .Z(n16488) );
  XOR U16893 ( .A(n16487), .B(n16488), .Z(n16455) );
  OR U16894 ( .A(n16445), .B(n16444), .Z(n16449) );
  NANDN U16895 ( .A(n16447), .B(n16446), .Z(n16448) );
  NAND U16896 ( .A(n16449), .B(n16448), .Z(n16456) );
  XNOR U16897 ( .A(n16455), .B(n16456), .Z(n16457) );
  XNOR U16898 ( .A(n16458), .B(n16457), .Z(n16491) );
  XNOR U16899 ( .A(n16491), .B(sreg[1415]), .Z(n16493) );
  NAND U16900 ( .A(n16450), .B(sreg[1414]), .Z(n16454) );
  OR U16901 ( .A(n16452), .B(n16451), .Z(n16453) );
  AND U16902 ( .A(n16454), .B(n16453), .Z(n16492) );
  XOR U16903 ( .A(n16493), .B(n16492), .Z(c[1415]) );
  NANDN U16904 ( .A(n16456), .B(n16455), .Z(n16460) );
  NAND U16905 ( .A(n16458), .B(n16457), .Z(n16459) );
  NAND U16906 ( .A(n16460), .B(n16459), .Z(n16499) );
  NAND U16907 ( .A(b[0]), .B(a[400]), .Z(n16461) );
  XNOR U16908 ( .A(b[1]), .B(n16461), .Z(n16463) );
  NAND U16909 ( .A(n72), .B(a[399]), .Z(n16462) );
  AND U16910 ( .A(n16463), .B(n16462), .Z(n16516) );
  XOR U16911 ( .A(a[396]), .B(n42197), .Z(n16505) );
  NANDN U16912 ( .A(n16505), .B(n42173), .Z(n16466) );
  NANDN U16913 ( .A(n16464), .B(n42172), .Z(n16465) );
  NAND U16914 ( .A(n16466), .B(n16465), .Z(n16514) );
  NAND U16915 ( .A(b[7]), .B(a[392]), .Z(n16515) );
  XNOR U16916 ( .A(n16514), .B(n16515), .Z(n16517) );
  XOR U16917 ( .A(n16516), .B(n16517), .Z(n16523) );
  NANDN U16918 ( .A(n16467), .B(n42093), .Z(n16469) );
  XOR U16919 ( .A(n42134), .B(a[398]), .Z(n16508) );
  NANDN U16920 ( .A(n16508), .B(n42095), .Z(n16468) );
  NAND U16921 ( .A(n16469), .B(n16468), .Z(n16521) );
  NANDN U16922 ( .A(n16470), .B(n42231), .Z(n16472) );
  XOR U16923 ( .A(n194), .B(a[394]), .Z(n16511) );
  NANDN U16924 ( .A(n16511), .B(n42234), .Z(n16471) );
  AND U16925 ( .A(n16472), .B(n16471), .Z(n16520) );
  XNOR U16926 ( .A(n16521), .B(n16520), .Z(n16522) );
  XNOR U16927 ( .A(n16523), .B(n16522), .Z(n16527) );
  NANDN U16928 ( .A(n16474), .B(n16473), .Z(n16478) );
  NAND U16929 ( .A(n16476), .B(n16475), .Z(n16477) );
  AND U16930 ( .A(n16478), .B(n16477), .Z(n16526) );
  XOR U16931 ( .A(n16527), .B(n16526), .Z(n16528) );
  NANDN U16932 ( .A(n16480), .B(n16479), .Z(n16484) );
  NANDN U16933 ( .A(n16482), .B(n16481), .Z(n16483) );
  NAND U16934 ( .A(n16484), .B(n16483), .Z(n16529) );
  XOR U16935 ( .A(n16528), .B(n16529), .Z(n16496) );
  OR U16936 ( .A(n16486), .B(n16485), .Z(n16490) );
  NANDN U16937 ( .A(n16488), .B(n16487), .Z(n16489) );
  NAND U16938 ( .A(n16490), .B(n16489), .Z(n16497) );
  XNOR U16939 ( .A(n16496), .B(n16497), .Z(n16498) );
  XNOR U16940 ( .A(n16499), .B(n16498), .Z(n16532) );
  XNOR U16941 ( .A(n16532), .B(sreg[1416]), .Z(n16534) );
  NAND U16942 ( .A(n16491), .B(sreg[1415]), .Z(n16495) );
  OR U16943 ( .A(n16493), .B(n16492), .Z(n16494) );
  AND U16944 ( .A(n16495), .B(n16494), .Z(n16533) );
  XOR U16945 ( .A(n16534), .B(n16533), .Z(c[1416]) );
  NANDN U16946 ( .A(n16497), .B(n16496), .Z(n16501) );
  NAND U16947 ( .A(n16499), .B(n16498), .Z(n16500) );
  NAND U16948 ( .A(n16501), .B(n16500), .Z(n16540) );
  NAND U16949 ( .A(b[0]), .B(a[401]), .Z(n16502) );
  XNOR U16950 ( .A(b[1]), .B(n16502), .Z(n16504) );
  NAND U16951 ( .A(n72), .B(a[400]), .Z(n16503) );
  AND U16952 ( .A(n16504), .B(n16503), .Z(n16557) );
  XOR U16953 ( .A(a[397]), .B(n42197), .Z(n16546) );
  NANDN U16954 ( .A(n16546), .B(n42173), .Z(n16507) );
  NANDN U16955 ( .A(n16505), .B(n42172), .Z(n16506) );
  NAND U16956 ( .A(n16507), .B(n16506), .Z(n16555) );
  NAND U16957 ( .A(b[7]), .B(a[393]), .Z(n16556) );
  XNOR U16958 ( .A(n16555), .B(n16556), .Z(n16558) );
  XOR U16959 ( .A(n16557), .B(n16558), .Z(n16564) );
  NANDN U16960 ( .A(n16508), .B(n42093), .Z(n16510) );
  XOR U16961 ( .A(n42134), .B(a[399]), .Z(n16549) );
  NANDN U16962 ( .A(n16549), .B(n42095), .Z(n16509) );
  NAND U16963 ( .A(n16510), .B(n16509), .Z(n16562) );
  NANDN U16964 ( .A(n16511), .B(n42231), .Z(n16513) );
  XOR U16965 ( .A(n195), .B(a[395]), .Z(n16552) );
  NANDN U16966 ( .A(n16552), .B(n42234), .Z(n16512) );
  AND U16967 ( .A(n16513), .B(n16512), .Z(n16561) );
  XNOR U16968 ( .A(n16562), .B(n16561), .Z(n16563) );
  XNOR U16969 ( .A(n16564), .B(n16563), .Z(n16568) );
  NANDN U16970 ( .A(n16515), .B(n16514), .Z(n16519) );
  NAND U16971 ( .A(n16517), .B(n16516), .Z(n16518) );
  AND U16972 ( .A(n16519), .B(n16518), .Z(n16567) );
  XOR U16973 ( .A(n16568), .B(n16567), .Z(n16569) );
  NANDN U16974 ( .A(n16521), .B(n16520), .Z(n16525) );
  NANDN U16975 ( .A(n16523), .B(n16522), .Z(n16524) );
  NAND U16976 ( .A(n16525), .B(n16524), .Z(n16570) );
  XOR U16977 ( .A(n16569), .B(n16570), .Z(n16537) );
  OR U16978 ( .A(n16527), .B(n16526), .Z(n16531) );
  NANDN U16979 ( .A(n16529), .B(n16528), .Z(n16530) );
  NAND U16980 ( .A(n16531), .B(n16530), .Z(n16538) );
  XNOR U16981 ( .A(n16537), .B(n16538), .Z(n16539) );
  XNOR U16982 ( .A(n16540), .B(n16539), .Z(n16573) );
  XNOR U16983 ( .A(n16573), .B(sreg[1417]), .Z(n16575) );
  NAND U16984 ( .A(n16532), .B(sreg[1416]), .Z(n16536) );
  OR U16985 ( .A(n16534), .B(n16533), .Z(n16535) );
  AND U16986 ( .A(n16536), .B(n16535), .Z(n16574) );
  XOR U16987 ( .A(n16575), .B(n16574), .Z(c[1417]) );
  NANDN U16988 ( .A(n16538), .B(n16537), .Z(n16542) );
  NAND U16989 ( .A(n16540), .B(n16539), .Z(n16541) );
  NAND U16990 ( .A(n16542), .B(n16541), .Z(n16581) );
  NAND U16991 ( .A(b[0]), .B(a[402]), .Z(n16543) );
  XNOR U16992 ( .A(b[1]), .B(n16543), .Z(n16545) );
  NAND U16993 ( .A(n72), .B(a[401]), .Z(n16544) );
  AND U16994 ( .A(n16545), .B(n16544), .Z(n16598) );
  XOR U16995 ( .A(a[398]), .B(n42197), .Z(n16587) );
  NANDN U16996 ( .A(n16587), .B(n42173), .Z(n16548) );
  NANDN U16997 ( .A(n16546), .B(n42172), .Z(n16547) );
  NAND U16998 ( .A(n16548), .B(n16547), .Z(n16596) );
  NAND U16999 ( .A(b[7]), .B(a[394]), .Z(n16597) );
  XNOR U17000 ( .A(n16596), .B(n16597), .Z(n16599) );
  XOR U17001 ( .A(n16598), .B(n16599), .Z(n16605) );
  NANDN U17002 ( .A(n16549), .B(n42093), .Z(n16551) );
  XOR U17003 ( .A(n42134), .B(a[400]), .Z(n16590) );
  NANDN U17004 ( .A(n16590), .B(n42095), .Z(n16550) );
  NAND U17005 ( .A(n16551), .B(n16550), .Z(n16603) );
  NANDN U17006 ( .A(n16552), .B(n42231), .Z(n16554) );
  XOR U17007 ( .A(n195), .B(a[396]), .Z(n16593) );
  NANDN U17008 ( .A(n16593), .B(n42234), .Z(n16553) );
  AND U17009 ( .A(n16554), .B(n16553), .Z(n16602) );
  XNOR U17010 ( .A(n16603), .B(n16602), .Z(n16604) );
  XNOR U17011 ( .A(n16605), .B(n16604), .Z(n16609) );
  NANDN U17012 ( .A(n16556), .B(n16555), .Z(n16560) );
  NAND U17013 ( .A(n16558), .B(n16557), .Z(n16559) );
  AND U17014 ( .A(n16560), .B(n16559), .Z(n16608) );
  XOR U17015 ( .A(n16609), .B(n16608), .Z(n16610) );
  NANDN U17016 ( .A(n16562), .B(n16561), .Z(n16566) );
  NANDN U17017 ( .A(n16564), .B(n16563), .Z(n16565) );
  NAND U17018 ( .A(n16566), .B(n16565), .Z(n16611) );
  XOR U17019 ( .A(n16610), .B(n16611), .Z(n16578) );
  OR U17020 ( .A(n16568), .B(n16567), .Z(n16572) );
  NANDN U17021 ( .A(n16570), .B(n16569), .Z(n16571) );
  NAND U17022 ( .A(n16572), .B(n16571), .Z(n16579) );
  XNOR U17023 ( .A(n16578), .B(n16579), .Z(n16580) );
  XNOR U17024 ( .A(n16581), .B(n16580), .Z(n16614) );
  XNOR U17025 ( .A(n16614), .B(sreg[1418]), .Z(n16616) );
  NAND U17026 ( .A(n16573), .B(sreg[1417]), .Z(n16577) );
  OR U17027 ( .A(n16575), .B(n16574), .Z(n16576) );
  AND U17028 ( .A(n16577), .B(n16576), .Z(n16615) );
  XOR U17029 ( .A(n16616), .B(n16615), .Z(c[1418]) );
  NANDN U17030 ( .A(n16579), .B(n16578), .Z(n16583) );
  NAND U17031 ( .A(n16581), .B(n16580), .Z(n16582) );
  NAND U17032 ( .A(n16583), .B(n16582), .Z(n16622) );
  NAND U17033 ( .A(b[0]), .B(a[403]), .Z(n16584) );
  XNOR U17034 ( .A(b[1]), .B(n16584), .Z(n16586) );
  NAND U17035 ( .A(n72), .B(a[402]), .Z(n16585) );
  AND U17036 ( .A(n16586), .B(n16585), .Z(n16639) );
  XOR U17037 ( .A(a[399]), .B(n42197), .Z(n16628) );
  NANDN U17038 ( .A(n16628), .B(n42173), .Z(n16589) );
  NANDN U17039 ( .A(n16587), .B(n42172), .Z(n16588) );
  NAND U17040 ( .A(n16589), .B(n16588), .Z(n16637) );
  NAND U17041 ( .A(b[7]), .B(a[395]), .Z(n16638) );
  XNOR U17042 ( .A(n16637), .B(n16638), .Z(n16640) );
  XOR U17043 ( .A(n16639), .B(n16640), .Z(n16646) );
  NANDN U17044 ( .A(n16590), .B(n42093), .Z(n16592) );
  XOR U17045 ( .A(n42134), .B(a[401]), .Z(n16631) );
  NANDN U17046 ( .A(n16631), .B(n42095), .Z(n16591) );
  NAND U17047 ( .A(n16592), .B(n16591), .Z(n16644) );
  NANDN U17048 ( .A(n16593), .B(n42231), .Z(n16595) );
  XOR U17049 ( .A(n195), .B(a[397]), .Z(n16634) );
  NANDN U17050 ( .A(n16634), .B(n42234), .Z(n16594) );
  AND U17051 ( .A(n16595), .B(n16594), .Z(n16643) );
  XNOR U17052 ( .A(n16644), .B(n16643), .Z(n16645) );
  XNOR U17053 ( .A(n16646), .B(n16645), .Z(n16650) );
  NANDN U17054 ( .A(n16597), .B(n16596), .Z(n16601) );
  NAND U17055 ( .A(n16599), .B(n16598), .Z(n16600) );
  AND U17056 ( .A(n16601), .B(n16600), .Z(n16649) );
  XOR U17057 ( .A(n16650), .B(n16649), .Z(n16651) );
  NANDN U17058 ( .A(n16603), .B(n16602), .Z(n16607) );
  NANDN U17059 ( .A(n16605), .B(n16604), .Z(n16606) );
  NAND U17060 ( .A(n16607), .B(n16606), .Z(n16652) );
  XOR U17061 ( .A(n16651), .B(n16652), .Z(n16619) );
  OR U17062 ( .A(n16609), .B(n16608), .Z(n16613) );
  NANDN U17063 ( .A(n16611), .B(n16610), .Z(n16612) );
  NAND U17064 ( .A(n16613), .B(n16612), .Z(n16620) );
  XNOR U17065 ( .A(n16619), .B(n16620), .Z(n16621) );
  XNOR U17066 ( .A(n16622), .B(n16621), .Z(n16655) );
  XNOR U17067 ( .A(n16655), .B(sreg[1419]), .Z(n16657) );
  NAND U17068 ( .A(n16614), .B(sreg[1418]), .Z(n16618) );
  OR U17069 ( .A(n16616), .B(n16615), .Z(n16617) );
  AND U17070 ( .A(n16618), .B(n16617), .Z(n16656) );
  XOR U17071 ( .A(n16657), .B(n16656), .Z(c[1419]) );
  NANDN U17072 ( .A(n16620), .B(n16619), .Z(n16624) );
  NAND U17073 ( .A(n16622), .B(n16621), .Z(n16623) );
  NAND U17074 ( .A(n16624), .B(n16623), .Z(n16663) );
  NAND U17075 ( .A(b[0]), .B(a[404]), .Z(n16625) );
  XNOR U17076 ( .A(b[1]), .B(n16625), .Z(n16627) );
  NAND U17077 ( .A(n72), .B(a[403]), .Z(n16626) );
  AND U17078 ( .A(n16627), .B(n16626), .Z(n16680) );
  XOR U17079 ( .A(a[400]), .B(n42197), .Z(n16669) );
  NANDN U17080 ( .A(n16669), .B(n42173), .Z(n16630) );
  NANDN U17081 ( .A(n16628), .B(n42172), .Z(n16629) );
  NAND U17082 ( .A(n16630), .B(n16629), .Z(n16678) );
  NAND U17083 ( .A(b[7]), .B(a[396]), .Z(n16679) );
  XNOR U17084 ( .A(n16678), .B(n16679), .Z(n16681) );
  XOR U17085 ( .A(n16680), .B(n16681), .Z(n16687) );
  NANDN U17086 ( .A(n16631), .B(n42093), .Z(n16633) );
  XOR U17087 ( .A(n42134), .B(a[402]), .Z(n16672) );
  NANDN U17088 ( .A(n16672), .B(n42095), .Z(n16632) );
  NAND U17089 ( .A(n16633), .B(n16632), .Z(n16685) );
  NANDN U17090 ( .A(n16634), .B(n42231), .Z(n16636) );
  XOR U17091 ( .A(n195), .B(a[398]), .Z(n16675) );
  NANDN U17092 ( .A(n16675), .B(n42234), .Z(n16635) );
  AND U17093 ( .A(n16636), .B(n16635), .Z(n16684) );
  XNOR U17094 ( .A(n16685), .B(n16684), .Z(n16686) );
  XNOR U17095 ( .A(n16687), .B(n16686), .Z(n16691) );
  NANDN U17096 ( .A(n16638), .B(n16637), .Z(n16642) );
  NAND U17097 ( .A(n16640), .B(n16639), .Z(n16641) );
  AND U17098 ( .A(n16642), .B(n16641), .Z(n16690) );
  XOR U17099 ( .A(n16691), .B(n16690), .Z(n16692) );
  NANDN U17100 ( .A(n16644), .B(n16643), .Z(n16648) );
  NANDN U17101 ( .A(n16646), .B(n16645), .Z(n16647) );
  NAND U17102 ( .A(n16648), .B(n16647), .Z(n16693) );
  XOR U17103 ( .A(n16692), .B(n16693), .Z(n16660) );
  OR U17104 ( .A(n16650), .B(n16649), .Z(n16654) );
  NANDN U17105 ( .A(n16652), .B(n16651), .Z(n16653) );
  NAND U17106 ( .A(n16654), .B(n16653), .Z(n16661) );
  XNOR U17107 ( .A(n16660), .B(n16661), .Z(n16662) );
  XNOR U17108 ( .A(n16663), .B(n16662), .Z(n16696) );
  XNOR U17109 ( .A(n16696), .B(sreg[1420]), .Z(n16698) );
  NAND U17110 ( .A(n16655), .B(sreg[1419]), .Z(n16659) );
  OR U17111 ( .A(n16657), .B(n16656), .Z(n16658) );
  AND U17112 ( .A(n16659), .B(n16658), .Z(n16697) );
  XOR U17113 ( .A(n16698), .B(n16697), .Z(c[1420]) );
  NANDN U17114 ( .A(n16661), .B(n16660), .Z(n16665) );
  NAND U17115 ( .A(n16663), .B(n16662), .Z(n16664) );
  NAND U17116 ( .A(n16665), .B(n16664), .Z(n16704) );
  NAND U17117 ( .A(b[0]), .B(a[405]), .Z(n16666) );
  XNOR U17118 ( .A(b[1]), .B(n16666), .Z(n16668) );
  NAND U17119 ( .A(n72), .B(a[404]), .Z(n16667) );
  AND U17120 ( .A(n16668), .B(n16667), .Z(n16721) );
  XOR U17121 ( .A(a[401]), .B(n42197), .Z(n16710) );
  NANDN U17122 ( .A(n16710), .B(n42173), .Z(n16671) );
  NANDN U17123 ( .A(n16669), .B(n42172), .Z(n16670) );
  NAND U17124 ( .A(n16671), .B(n16670), .Z(n16719) );
  NAND U17125 ( .A(b[7]), .B(a[397]), .Z(n16720) );
  XNOR U17126 ( .A(n16719), .B(n16720), .Z(n16722) );
  XOR U17127 ( .A(n16721), .B(n16722), .Z(n16728) );
  NANDN U17128 ( .A(n16672), .B(n42093), .Z(n16674) );
  XOR U17129 ( .A(n42134), .B(a[403]), .Z(n16713) );
  NANDN U17130 ( .A(n16713), .B(n42095), .Z(n16673) );
  NAND U17131 ( .A(n16674), .B(n16673), .Z(n16726) );
  NANDN U17132 ( .A(n16675), .B(n42231), .Z(n16677) );
  XOR U17133 ( .A(n195), .B(a[399]), .Z(n16716) );
  NANDN U17134 ( .A(n16716), .B(n42234), .Z(n16676) );
  AND U17135 ( .A(n16677), .B(n16676), .Z(n16725) );
  XNOR U17136 ( .A(n16726), .B(n16725), .Z(n16727) );
  XNOR U17137 ( .A(n16728), .B(n16727), .Z(n16732) );
  NANDN U17138 ( .A(n16679), .B(n16678), .Z(n16683) );
  NAND U17139 ( .A(n16681), .B(n16680), .Z(n16682) );
  AND U17140 ( .A(n16683), .B(n16682), .Z(n16731) );
  XOR U17141 ( .A(n16732), .B(n16731), .Z(n16733) );
  NANDN U17142 ( .A(n16685), .B(n16684), .Z(n16689) );
  NANDN U17143 ( .A(n16687), .B(n16686), .Z(n16688) );
  NAND U17144 ( .A(n16689), .B(n16688), .Z(n16734) );
  XOR U17145 ( .A(n16733), .B(n16734), .Z(n16701) );
  OR U17146 ( .A(n16691), .B(n16690), .Z(n16695) );
  NANDN U17147 ( .A(n16693), .B(n16692), .Z(n16694) );
  NAND U17148 ( .A(n16695), .B(n16694), .Z(n16702) );
  XNOR U17149 ( .A(n16701), .B(n16702), .Z(n16703) );
  XNOR U17150 ( .A(n16704), .B(n16703), .Z(n16737) );
  XNOR U17151 ( .A(n16737), .B(sreg[1421]), .Z(n16739) );
  NAND U17152 ( .A(n16696), .B(sreg[1420]), .Z(n16700) );
  OR U17153 ( .A(n16698), .B(n16697), .Z(n16699) );
  AND U17154 ( .A(n16700), .B(n16699), .Z(n16738) );
  XOR U17155 ( .A(n16739), .B(n16738), .Z(c[1421]) );
  NANDN U17156 ( .A(n16702), .B(n16701), .Z(n16706) );
  NAND U17157 ( .A(n16704), .B(n16703), .Z(n16705) );
  NAND U17158 ( .A(n16706), .B(n16705), .Z(n16745) );
  NAND U17159 ( .A(b[0]), .B(a[406]), .Z(n16707) );
  XNOR U17160 ( .A(b[1]), .B(n16707), .Z(n16709) );
  NAND U17161 ( .A(n73), .B(a[405]), .Z(n16708) );
  AND U17162 ( .A(n16709), .B(n16708), .Z(n16762) );
  XOR U17163 ( .A(a[402]), .B(n42197), .Z(n16751) );
  NANDN U17164 ( .A(n16751), .B(n42173), .Z(n16712) );
  NANDN U17165 ( .A(n16710), .B(n42172), .Z(n16711) );
  NAND U17166 ( .A(n16712), .B(n16711), .Z(n16760) );
  NAND U17167 ( .A(b[7]), .B(a[398]), .Z(n16761) );
  XNOR U17168 ( .A(n16760), .B(n16761), .Z(n16763) );
  XOR U17169 ( .A(n16762), .B(n16763), .Z(n16769) );
  NANDN U17170 ( .A(n16713), .B(n42093), .Z(n16715) );
  XOR U17171 ( .A(n42134), .B(a[404]), .Z(n16754) );
  NANDN U17172 ( .A(n16754), .B(n42095), .Z(n16714) );
  NAND U17173 ( .A(n16715), .B(n16714), .Z(n16767) );
  NANDN U17174 ( .A(n16716), .B(n42231), .Z(n16718) );
  XOR U17175 ( .A(n195), .B(a[400]), .Z(n16757) );
  NANDN U17176 ( .A(n16757), .B(n42234), .Z(n16717) );
  AND U17177 ( .A(n16718), .B(n16717), .Z(n16766) );
  XNOR U17178 ( .A(n16767), .B(n16766), .Z(n16768) );
  XNOR U17179 ( .A(n16769), .B(n16768), .Z(n16773) );
  NANDN U17180 ( .A(n16720), .B(n16719), .Z(n16724) );
  NAND U17181 ( .A(n16722), .B(n16721), .Z(n16723) );
  AND U17182 ( .A(n16724), .B(n16723), .Z(n16772) );
  XOR U17183 ( .A(n16773), .B(n16772), .Z(n16774) );
  NANDN U17184 ( .A(n16726), .B(n16725), .Z(n16730) );
  NANDN U17185 ( .A(n16728), .B(n16727), .Z(n16729) );
  NAND U17186 ( .A(n16730), .B(n16729), .Z(n16775) );
  XOR U17187 ( .A(n16774), .B(n16775), .Z(n16742) );
  OR U17188 ( .A(n16732), .B(n16731), .Z(n16736) );
  NANDN U17189 ( .A(n16734), .B(n16733), .Z(n16735) );
  NAND U17190 ( .A(n16736), .B(n16735), .Z(n16743) );
  XNOR U17191 ( .A(n16742), .B(n16743), .Z(n16744) );
  XNOR U17192 ( .A(n16745), .B(n16744), .Z(n16778) );
  XNOR U17193 ( .A(n16778), .B(sreg[1422]), .Z(n16780) );
  NAND U17194 ( .A(n16737), .B(sreg[1421]), .Z(n16741) );
  OR U17195 ( .A(n16739), .B(n16738), .Z(n16740) );
  AND U17196 ( .A(n16741), .B(n16740), .Z(n16779) );
  XOR U17197 ( .A(n16780), .B(n16779), .Z(c[1422]) );
  NANDN U17198 ( .A(n16743), .B(n16742), .Z(n16747) );
  NAND U17199 ( .A(n16745), .B(n16744), .Z(n16746) );
  NAND U17200 ( .A(n16747), .B(n16746), .Z(n16786) );
  NAND U17201 ( .A(b[0]), .B(a[407]), .Z(n16748) );
  XNOR U17202 ( .A(b[1]), .B(n16748), .Z(n16750) );
  NAND U17203 ( .A(n73), .B(a[406]), .Z(n16749) );
  AND U17204 ( .A(n16750), .B(n16749), .Z(n16803) );
  XOR U17205 ( .A(a[403]), .B(n42197), .Z(n16792) );
  NANDN U17206 ( .A(n16792), .B(n42173), .Z(n16753) );
  NANDN U17207 ( .A(n16751), .B(n42172), .Z(n16752) );
  NAND U17208 ( .A(n16753), .B(n16752), .Z(n16801) );
  NAND U17209 ( .A(b[7]), .B(a[399]), .Z(n16802) );
  XNOR U17210 ( .A(n16801), .B(n16802), .Z(n16804) );
  XOR U17211 ( .A(n16803), .B(n16804), .Z(n16810) );
  NANDN U17212 ( .A(n16754), .B(n42093), .Z(n16756) );
  XOR U17213 ( .A(n42134), .B(a[405]), .Z(n16795) );
  NANDN U17214 ( .A(n16795), .B(n42095), .Z(n16755) );
  NAND U17215 ( .A(n16756), .B(n16755), .Z(n16808) );
  NANDN U17216 ( .A(n16757), .B(n42231), .Z(n16759) );
  XOR U17217 ( .A(n195), .B(a[401]), .Z(n16798) );
  NANDN U17218 ( .A(n16798), .B(n42234), .Z(n16758) );
  AND U17219 ( .A(n16759), .B(n16758), .Z(n16807) );
  XNOR U17220 ( .A(n16808), .B(n16807), .Z(n16809) );
  XNOR U17221 ( .A(n16810), .B(n16809), .Z(n16814) );
  NANDN U17222 ( .A(n16761), .B(n16760), .Z(n16765) );
  NAND U17223 ( .A(n16763), .B(n16762), .Z(n16764) );
  AND U17224 ( .A(n16765), .B(n16764), .Z(n16813) );
  XOR U17225 ( .A(n16814), .B(n16813), .Z(n16815) );
  NANDN U17226 ( .A(n16767), .B(n16766), .Z(n16771) );
  NANDN U17227 ( .A(n16769), .B(n16768), .Z(n16770) );
  NAND U17228 ( .A(n16771), .B(n16770), .Z(n16816) );
  XOR U17229 ( .A(n16815), .B(n16816), .Z(n16783) );
  OR U17230 ( .A(n16773), .B(n16772), .Z(n16777) );
  NANDN U17231 ( .A(n16775), .B(n16774), .Z(n16776) );
  NAND U17232 ( .A(n16777), .B(n16776), .Z(n16784) );
  XNOR U17233 ( .A(n16783), .B(n16784), .Z(n16785) );
  XNOR U17234 ( .A(n16786), .B(n16785), .Z(n16819) );
  XNOR U17235 ( .A(n16819), .B(sreg[1423]), .Z(n16821) );
  NAND U17236 ( .A(n16778), .B(sreg[1422]), .Z(n16782) );
  OR U17237 ( .A(n16780), .B(n16779), .Z(n16781) );
  AND U17238 ( .A(n16782), .B(n16781), .Z(n16820) );
  XOR U17239 ( .A(n16821), .B(n16820), .Z(c[1423]) );
  NANDN U17240 ( .A(n16784), .B(n16783), .Z(n16788) );
  NAND U17241 ( .A(n16786), .B(n16785), .Z(n16787) );
  NAND U17242 ( .A(n16788), .B(n16787), .Z(n16827) );
  NAND U17243 ( .A(b[0]), .B(a[408]), .Z(n16789) );
  XNOR U17244 ( .A(b[1]), .B(n16789), .Z(n16791) );
  NAND U17245 ( .A(n73), .B(a[407]), .Z(n16790) );
  AND U17246 ( .A(n16791), .B(n16790), .Z(n16844) );
  XOR U17247 ( .A(a[404]), .B(n42197), .Z(n16833) );
  NANDN U17248 ( .A(n16833), .B(n42173), .Z(n16794) );
  NANDN U17249 ( .A(n16792), .B(n42172), .Z(n16793) );
  NAND U17250 ( .A(n16794), .B(n16793), .Z(n16842) );
  NAND U17251 ( .A(b[7]), .B(a[400]), .Z(n16843) );
  XNOR U17252 ( .A(n16842), .B(n16843), .Z(n16845) );
  XOR U17253 ( .A(n16844), .B(n16845), .Z(n16851) );
  NANDN U17254 ( .A(n16795), .B(n42093), .Z(n16797) );
  XOR U17255 ( .A(n42134), .B(a[406]), .Z(n16836) );
  NANDN U17256 ( .A(n16836), .B(n42095), .Z(n16796) );
  NAND U17257 ( .A(n16797), .B(n16796), .Z(n16849) );
  NANDN U17258 ( .A(n16798), .B(n42231), .Z(n16800) );
  XOR U17259 ( .A(n195), .B(a[402]), .Z(n16839) );
  NANDN U17260 ( .A(n16839), .B(n42234), .Z(n16799) );
  AND U17261 ( .A(n16800), .B(n16799), .Z(n16848) );
  XNOR U17262 ( .A(n16849), .B(n16848), .Z(n16850) );
  XNOR U17263 ( .A(n16851), .B(n16850), .Z(n16855) );
  NANDN U17264 ( .A(n16802), .B(n16801), .Z(n16806) );
  NAND U17265 ( .A(n16804), .B(n16803), .Z(n16805) );
  AND U17266 ( .A(n16806), .B(n16805), .Z(n16854) );
  XOR U17267 ( .A(n16855), .B(n16854), .Z(n16856) );
  NANDN U17268 ( .A(n16808), .B(n16807), .Z(n16812) );
  NANDN U17269 ( .A(n16810), .B(n16809), .Z(n16811) );
  NAND U17270 ( .A(n16812), .B(n16811), .Z(n16857) );
  XOR U17271 ( .A(n16856), .B(n16857), .Z(n16824) );
  OR U17272 ( .A(n16814), .B(n16813), .Z(n16818) );
  NANDN U17273 ( .A(n16816), .B(n16815), .Z(n16817) );
  NAND U17274 ( .A(n16818), .B(n16817), .Z(n16825) );
  XNOR U17275 ( .A(n16824), .B(n16825), .Z(n16826) );
  XNOR U17276 ( .A(n16827), .B(n16826), .Z(n16860) );
  XNOR U17277 ( .A(n16860), .B(sreg[1424]), .Z(n16862) );
  NAND U17278 ( .A(n16819), .B(sreg[1423]), .Z(n16823) );
  OR U17279 ( .A(n16821), .B(n16820), .Z(n16822) );
  AND U17280 ( .A(n16823), .B(n16822), .Z(n16861) );
  XOR U17281 ( .A(n16862), .B(n16861), .Z(c[1424]) );
  NANDN U17282 ( .A(n16825), .B(n16824), .Z(n16829) );
  NAND U17283 ( .A(n16827), .B(n16826), .Z(n16828) );
  NAND U17284 ( .A(n16829), .B(n16828), .Z(n16868) );
  NAND U17285 ( .A(b[0]), .B(a[409]), .Z(n16830) );
  XNOR U17286 ( .A(b[1]), .B(n16830), .Z(n16832) );
  NAND U17287 ( .A(n73), .B(a[408]), .Z(n16831) );
  AND U17288 ( .A(n16832), .B(n16831), .Z(n16885) );
  XOR U17289 ( .A(a[405]), .B(n42197), .Z(n16874) );
  NANDN U17290 ( .A(n16874), .B(n42173), .Z(n16835) );
  NANDN U17291 ( .A(n16833), .B(n42172), .Z(n16834) );
  NAND U17292 ( .A(n16835), .B(n16834), .Z(n16883) );
  NAND U17293 ( .A(b[7]), .B(a[401]), .Z(n16884) );
  XNOR U17294 ( .A(n16883), .B(n16884), .Z(n16886) );
  XOR U17295 ( .A(n16885), .B(n16886), .Z(n16892) );
  NANDN U17296 ( .A(n16836), .B(n42093), .Z(n16838) );
  XOR U17297 ( .A(n42134), .B(a[407]), .Z(n16877) );
  NANDN U17298 ( .A(n16877), .B(n42095), .Z(n16837) );
  NAND U17299 ( .A(n16838), .B(n16837), .Z(n16890) );
  NANDN U17300 ( .A(n16839), .B(n42231), .Z(n16841) );
  XOR U17301 ( .A(n195), .B(a[403]), .Z(n16880) );
  NANDN U17302 ( .A(n16880), .B(n42234), .Z(n16840) );
  AND U17303 ( .A(n16841), .B(n16840), .Z(n16889) );
  XNOR U17304 ( .A(n16890), .B(n16889), .Z(n16891) );
  XNOR U17305 ( .A(n16892), .B(n16891), .Z(n16896) );
  NANDN U17306 ( .A(n16843), .B(n16842), .Z(n16847) );
  NAND U17307 ( .A(n16845), .B(n16844), .Z(n16846) );
  AND U17308 ( .A(n16847), .B(n16846), .Z(n16895) );
  XOR U17309 ( .A(n16896), .B(n16895), .Z(n16897) );
  NANDN U17310 ( .A(n16849), .B(n16848), .Z(n16853) );
  NANDN U17311 ( .A(n16851), .B(n16850), .Z(n16852) );
  NAND U17312 ( .A(n16853), .B(n16852), .Z(n16898) );
  XOR U17313 ( .A(n16897), .B(n16898), .Z(n16865) );
  OR U17314 ( .A(n16855), .B(n16854), .Z(n16859) );
  NANDN U17315 ( .A(n16857), .B(n16856), .Z(n16858) );
  NAND U17316 ( .A(n16859), .B(n16858), .Z(n16866) );
  XNOR U17317 ( .A(n16865), .B(n16866), .Z(n16867) );
  XNOR U17318 ( .A(n16868), .B(n16867), .Z(n16901) );
  XNOR U17319 ( .A(n16901), .B(sreg[1425]), .Z(n16903) );
  NAND U17320 ( .A(n16860), .B(sreg[1424]), .Z(n16864) );
  OR U17321 ( .A(n16862), .B(n16861), .Z(n16863) );
  AND U17322 ( .A(n16864), .B(n16863), .Z(n16902) );
  XOR U17323 ( .A(n16903), .B(n16902), .Z(c[1425]) );
  NANDN U17324 ( .A(n16866), .B(n16865), .Z(n16870) );
  NAND U17325 ( .A(n16868), .B(n16867), .Z(n16869) );
  NAND U17326 ( .A(n16870), .B(n16869), .Z(n16909) );
  NAND U17327 ( .A(b[0]), .B(a[410]), .Z(n16871) );
  XNOR U17328 ( .A(b[1]), .B(n16871), .Z(n16873) );
  NAND U17329 ( .A(n73), .B(a[409]), .Z(n16872) );
  AND U17330 ( .A(n16873), .B(n16872), .Z(n16926) );
  XOR U17331 ( .A(a[406]), .B(n42197), .Z(n16915) );
  NANDN U17332 ( .A(n16915), .B(n42173), .Z(n16876) );
  NANDN U17333 ( .A(n16874), .B(n42172), .Z(n16875) );
  NAND U17334 ( .A(n16876), .B(n16875), .Z(n16924) );
  NAND U17335 ( .A(b[7]), .B(a[402]), .Z(n16925) );
  XNOR U17336 ( .A(n16924), .B(n16925), .Z(n16927) );
  XOR U17337 ( .A(n16926), .B(n16927), .Z(n16933) );
  NANDN U17338 ( .A(n16877), .B(n42093), .Z(n16879) );
  XOR U17339 ( .A(n42134), .B(a[408]), .Z(n16918) );
  NANDN U17340 ( .A(n16918), .B(n42095), .Z(n16878) );
  NAND U17341 ( .A(n16879), .B(n16878), .Z(n16931) );
  NANDN U17342 ( .A(n16880), .B(n42231), .Z(n16882) );
  XOR U17343 ( .A(n195), .B(a[404]), .Z(n16921) );
  NANDN U17344 ( .A(n16921), .B(n42234), .Z(n16881) );
  AND U17345 ( .A(n16882), .B(n16881), .Z(n16930) );
  XNOR U17346 ( .A(n16931), .B(n16930), .Z(n16932) );
  XNOR U17347 ( .A(n16933), .B(n16932), .Z(n16937) );
  NANDN U17348 ( .A(n16884), .B(n16883), .Z(n16888) );
  NAND U17349 ( .A(n16886), .B(n16885), .Z(n16887) );
  AND U17350 ( .A(n16888), .B(n16887), .Z(n16936) );
  XOR U17351 ( .A(n16937), .B(n16936), .Z(n16938) );
  NANDN U17352 ( .A(n16890), .B(n16889), .Z(n16894) );
  NANDN U17353 ( .A(n16892), .B(n16891), .Z(n16893) );
  NAND U17354 ( .A(n16894), .B(n16893), .Z(n16939) );
  XOR U17355 ( .A(n16938), .B(n16939), .Z(n16906) );
  OR U17356 ( .A(n16896), .B(n16895), .Z(n16900) );
  NANDN U17357 ( .A(n16898), .B(n16897), .Z(n16899) );
  NAND U17358 ( .A(n16900), .B(n16899), .Z(n16907) );
  XNOR U17359 ( .A(n16906), .B(n16907), .Z(n16908) );
  XNOR U17360 ( .A(n16909), .B(n16908), .Z(n16942) );
  XNOR U17361 ( .A(n16942), .B(sreg[1426]), .Z(n16944) );
  NAND U17362 ( .A(n16901), .B(sreg[1425]), .Z(n16905) );
  OR U17363 ( .A(n16903), .B(n16902), .Z(n16904) );
  AND U17364 ( .A(n16905), .B(n16904), .Z(n16943) );
  XOR U17365 ( .A(n16944), .B(n16943), .Z(c[1426]) );
  NANDN U17366 ( .A(n16907), .B(n16906), .Z(n16911) );
  NAND U17367 ( .A(n16909), .B(n16908), .Z(n16910) );
  NAND U17368 ( .A(n16911), .B(n16910), .Z(n16950) );
  NAND U17369 ( .A(b[0]), .B(a[411]), .Z(n16912) );
  XNOR U17370 ( .A(b[1]), .B(n16912), .Z(n16914) );
  NAND U17371 ( .A(n73), .B(a[410]), .Z(n16913) );
  AND U17372 ( .A(n16914), .B(n16913), .Z(n16967) );
  XOR U17373 ( .A(a[407]), .B(n42197), .Z(n16956) );
  NANDN U17374 ( .A(n16956), .B(n42173), .Z(n16917) );
  NANDN U17375 ( .A(n16915), .B(n42172), .Z(n16916) );
  NAND U17376 ( .A(n16917), .B(n16916), .Z(n16965) );
  NAND U17377 ( .A(b[7]), .B(a[403]), .Z(n16966) );
  XNOR U17378 ( .A(n16965), .B(n16966), .Z(n16968) );
  XOR U17379 ( .A(n16967), .B(n16968), .Z(n16974) );
  NANDN U17380 ( .A(n16918), .B(n42093), .Z(n16920) );
  XOR U17381 ( .A(n42134), .B(a[409]), .Z(n16959) );
  NANDN U17382 ( .A(n16959), .B(n42095), .Z(n16919) );
  NAND U17383 ( .A(n16920), .B(n16919), .Z(n16972) );
  NANDN U17384 ( .A(n16921), .B(n42231), .Z(n16923) );
  XOR U17385 ( .A(n195), .B(a[405]), .Z(n16962) );
  NANDN U17386 ( .A(n16962), .B(n42234), .Z(n16922) );
  AND U17387 ( .A(n16923), .B(n16922), .Z(n16971) );
  XNOR U17388 ( .A(n16972), .B(n16971), .Z(n16973) );
  XNOR U17389 ( .A(n16974), .B(n16973), .Z(n16978) );
  NANDN U17390 ( .A(n16925), .B(n16924), .Z(n16929) );
  NAND U17391 ( .A(n16927), .B(n16926), .Z(n16928) );
  AND U17392 ( .A(n16929), .B(n16928), .Z(n16977) );
  XOR U17393 ( .A(n16978), .B(n16977), .Z(n16979) );
  NANDN U17394 ( .A(n16931), .B(n16930), .Z(n16935) );
  NANDN U17395 ( .A(n16933), .B(n16932), .Z(n16934) );
  NAND U17396 ( .A(n16935), .B(n16934), .Z(n16980) );
  XOR U17397 ( .A(n16979), .B(n16980), .Z(n16947) );
  OR U17398 ( .A(n16937), .B(n16936), .Z(n16941) );
  NANDN U17399 ( .A(n16939), .B(n16938), .Z(n16940) );
  NAND U17400 ( .A(n16941), .B(n16940), .Z(n16948) );
  XNOR U17401 ( .A(n16947), .B(n16948), .Z(n16949) );
  XNOR U17402 ( .A(n16950), .B(n16949), .Z(n16983) );
  XNOR U17403 ( .A(n16983), .B(sreg[1427]), .Z(n16985) );
  NAND U17404 ( .A(n16942), .B(sreg[1426]), .Z(n16946) );
  OR U17405 ( .A(n16944), .B(n16943), .Z(n16945) );
  AND U17406 ( .A(n16946), .B(n16945), .Z(n16984) );
  XOR U17407 ( .A(n16985), .B(n16984), .Z(c[1427]) );
  NANDN U17408 ( .A(n16948), .B(n16947), .Z(n16952) );
  NAND U17409 ( .A(n16950), .B(n16949), .Z(n16951) );
  NAND U17410 ( .A(n16952), .B(n16951), .Z(n16991) );
  NAND U17411 ( .A(b[0]), .B(a[412]), .Z(n16953) );
  XNOR U17412 ( .A(b[1]), .B(n16953), .Z(n16955) );
  NAND U17413 ( .A(n73), .B(a[411]), .Z(n16954) );
  AND U17414 ( .A(n16955), .B(n16954), .Z(n17008) );
  XOR U17415 ( .A(a[408]), .B(n42197), .Z(n16997) );
  NANDN U17416 ( .A(n16997), .B(n42173), .Z(n16958) );
  NANDN U17417 ( .A(n16956), .B(n42172), .Z(n16957) );
  NAND U17418 ( .A(n16958), .B(n16957), .Z(n17006) );
  NAND U17419 ( .A(b[7]), .B(a[404]), .Z(n17007) );
  XNOR U17420 ( .A(n17006), .B(n17007), .Z(n17009) );
  XOR U17421 ( .A(n17008), .B(n17009), .Z(n17015) );
  NANDN U17422 ( .A(n16959), .B(n42093), .Z(n16961) );
  XOR U17423 ( .A(n42134), .B(a[410]), .Z(n17000) );
  NANDN U17424 ( .A(n17000), .B(n42095), .Z(n16960) );
  NAND U17425 ( .A(n16961), .B(n16960), .Z(n17013) );
  NANDN U17426 ( .A(n16962), .B(n42231), .Z(n16964) );
  XOR U17427 ( .A(n195), .B(a[406]), .Z(n17003) );
  NANDN U17428 ( .A(n17003), .B(n42234), .Z(n16963) );
  AND U17429 ( .A(n16964), .B(n16963), .Z(n17012) );
  XNOR U17430 ( .A(n17013), .B(n17012), .Z(n17014) );
  XNOR U17431 ( .A(n17015), .B(n17014), .Z(n17019) );
  NANDN U17432 ( .A(n16966), .B(n16965), .Z(n16970) );
  NAND U17433 ( .A(n16968), .B(n16967), .Z(n16969) );
  AND U17434 ( .A(n16970), .B(n16969), .Z(n17018) );
  XOR U17435 ( .A(n17019), .B(n17018), .Z(n17020) );
  NANDN U17436 ( .A(n16972), .B(n16971), .Z(n16976) );
  NANDN U17437 ( .A(n16974), .B(n16973), .Z(n16975) );
  NAND U17438 ( .A(n16976), .B(n16975), .Z(n17021) );
  XOR U17439 ( .A(n17020), .B(n17021), .Z(n16988) );
  OR U17440 ( .A(n16978), .B(n16977), .Z(n16982) );
  NANDN U17441 ( .A(n16980), .B(n16979), .Z(n16981) );
  NAND U17442 ( .A(n16982), .B(n16981), .Z(n16989) );
  XNOR U17443 ( .A(n16988), .B(n16989), .Z(n16990) );
  XNOR U17444 ( .A(n16991), .B(n16990), .Z(n17024) );
  XNOR U17445 ( .A(n17024), .B(sreg[1428]), .Z(n17026) );
  NAND U17446 ( .A(n16983), .B(sreg[1427]), .Z(n16987) );
  OR U17447 ( .A(n16985), .B(n16984), .Z(n16986) );
  AND U17448 ( .A(n16987), .B(n16986), .Z(n17025) );
  XOR U17449 ( .A(n17026), .B(n17025), .Z(c[1428]) );
  NANDN U17450 ( .A(n16989), .B(n16988), .Z(n16993) );
  NAND U17451 ( .A(n16991), .B(n16990), .Z(n16992) );
  NAND U17452 ( .A(n16993), .B(n16992), .Z(n17032) );
  NAND U17453 ( .A(b[0]), .B(a[413]), .Z(n16994) );
  XNOR U17454 ( .A(b[1]), .B(n16994), .Z(n16996) );
  NAND U17455 ( .A(n74), .B(a[412]), .Z(n16995) );
  AND U17456 ( .A(n16996), .B(n16995), .Z(n17049) );
  XOR U17457 ( .A(a[409]), .B(n42197), .Z(n17038) );
  NANDN U17458 ( .A(n17038), .B(n42173), .Z(n16999) );
  NANDN U17459 ( .A(n16997), .B(n42172), .Z(n16998) );
  NAND U17460 ( .A(n16999), .B(n16998), .Z(n17047) );
  NAND U17461 ( .A(b[7]), .B(a[405]), .Z(n17048) );
  XNOR U17462 ( .A(n17047), .B(n17048), .Z(n17050) );
  XOR U17463 ( .A(n17049), .B(n17050), .Z(n17056) );
  NANDN U17464 ( .A(n17000), .B(n42093), .Z(n17002) );
  XOR U17465 ( .A(n42134), .B(a[411]), .Z(n17041) );
  NANDN U17466 ( .A(n17041), .B(n42095), .Z(n17001) );
  NAND U17467 ( .A(n17002), .B(n17001), .Z(n17054) );
  NANDN U17468 ( .A(n17003), .B(n42231), .Z(n17005) );
  XOR U17469 ( .A(n196), .B(a[407]), .Z(n17044) );
  NANDN U17470 ( .A(n17044), .B(n42234), .Z(n17004) );
  AND U17471 ( .A(n17005), .B(n17004), .Z(n17053) );
  XNOR U17472 ( .A(n17054), .B(n17053), .Z(n17055) );
  XNOR U17473 ( .A(n17056), .B(n17055), .Z(n17060) );
  NANDN U17474 ( .A(n17007), .B(n17006), .Z(n17011) );
  NAND U17475 ( .A(n17009), .B(n17008), .Z(n17010) );
  AND U17476 ( .A(n17011), .B(n17010), .Z(n17059) );
  XOR U17477 ( .A(n17060), .B(n17059), .Z(n17061) );
  NANDN U17478 ( .A(n17013), .B(n17012), .Z(n17017) );
  NANDN U17479 ( .A(n17015), .B(n17014), .Z(n17016) );
  NAND U17480 ( .A(n17017), .B(n17016), .Z(n17062) );
  XOR U17481 ( .A(n17061), .B(n17062), .Z(n17029) );
  OR U17482 ( .A(n17019), .B(n17018), .Z(n17023) );
  NANDN U17483 ( .A(n17021), .B(n17020), .Z(n17022) );
  NAND U17484 ( .A(n17023), .B(n17022), .Z(n17030) );
  XNOR U17485 ( .A(n17029), .B(n17030), .Z(n17031) );
  XNOR U17486 ( .A(n17032), .B(n17031), .Z(n17065) );
  XNOR U17487 ( .A(n17065), .B(sreg[1429]), .Z(n17067) );
  NAND U17488 ( .A(n17024), .B(sreg[1428]), .Z(n17028) );
  OR U17489 ( .A(n17026), .B(n17025), .Z(n17027) );
  AND U17490 ( .A(n17028), .B(n17027), .Z(n17066) );
  XOR U17491 ( .A(n17067), .B(n17066), .Z(c[1429]) );
  NANDN U17492 ( .A(n17030), .B(n17029), .Z(n17034) );
  NAND U17493 ( .A(n17032), .B(n17031), .Z(n17033) );
  NAND U17494 ( .A(n17034), .B(n17033), .Z(n17073) );
  NAND U17495 ( .A(b[0]), .B(a[414]), .Z(n17035) );
  XNOR U17496 ( .A(b[1]), .B(n17035), .Z(n17037) );
  NAND U17497 ( .A(n74), .B(a[413]), .Z(n17036) );
  AND U17498 ( .A(n17037), .B(n17036), .Z(n17090) );
  XOR U17499 ( .A(a[410]), .B(n42197), .Z(n17079) );
  NANDN U17500 ( .A(n17079), .B(n42173), .Z(n17040) );
  NANDN U17501 ( .A(n17038), .B(n42172), .Z(n17039) );
  NAND U17502 ( .A(n17040), .B(n17039), .Z(n17088) );
  NAND U17503 ( .A(b[7]), .B(a[406]), .Z(n17089) );
  XNOR U17504 ( .A(n17088), .B(n17089), .Z(n17091) );
  XOR U17505 ( .A(n17090), .B(n17091), .Z(n17097) );
  NANDN U17506 ( .A(n17041), .B(n42093), .Z(n17043) );
  XOR U17507 ( .A(n42134), .B(a[412]), .Z(n17082) );
  NANDN U17508 ( .A(n17082), .B(n42095), .Z(n17042) );
  NAND U17509 ( .A(n17043), .B(n17042), .Z(n17095) );
  NANDN U17510 ( .A(n17044), .B(n42231), .Z(n17046) );
  XOR U17511 ( .A(n196), .B(a[408]), .Z(n17085) );
  NANDN U17512 ( .A(n17085), .B(n42234), .Z(n17045) );
  AND U17513 ( .A(n17046), .B(n17045), .Z(n17094) );
  XNOR U17514 ( .A(n17095), .B(n17094), .Z(n17096) );
  XNOR U17515 ( .A(n17097), .B(n17096), .Z(n17101) );
  NANDN U17516 ( .A(n17048), .B(n17047), .Z(n17052) );
  NAND U17517 ( .A(n17050), .B(n17049), .Z(n17051) );
  AND U17518 ( .A(n17052), .B(n17051), .Z(n17100) );
  XOR U17519 ( .A(n17101), .B(n17100), .Z(n17102) );
  NANDN U17520 ( .A(n17054), .B(n17053), .Z(n17058) );
  NANDN U17521 ( .A(n17056), .B(n17055), .Z(n17057) );
  NAND U17522 ( .A(n17058), .B(n17057), .Z(n17103) );
  XOR U17523 ( .A(n17102), .B(n17103), .Z(n17070) );
  OR U17524 ( .A(n17060), .B(n17059), .Z(n17064) );
  NANDN U17525 ( .A(n17062), .B(n17061), .Z(n17063) );
  NAND U17526 ( .A(n17064), .B(n17063), .Z(n17071) );
  XNOR U17527 ( .A(n17070), .B(n17071), .Z(n17072) );
  XNOR U17528 ( .A(n17073), .B(n17072), .Z(n17106) );
  XNOR U17529 ( .A(n17106), .B(sreg[1430]), .Z(n17108) );
  NAND U17530 ( .A(n17065), .B(sreg[1429]), .Z(n17069) );
  OR U17531 ( .A(n17067), .B(n17066), .Z(n17068) );
  AND U17532 ( .A(n17069), .B(n17068), .Z(n17107) );
  XOR U17533 ( .A(n17108), .B(n17107), .Z(c[1430]) );
  NANDN U17534 ( .A(n17071), .B(n17070), .Z(n17075) );
  NAND U17535 ( .A(n17073), .B(n17072), .Z(n17074) );
  NAND U17536 ( .A(n17075), .B(n17074), .Z(n17114) );
  NAND U17537 ( .A(b[0]), .B(a[415]), .Z(n17076) );
  XNOR U17538 ( .A(b[1]), .B(n17076), .Z(n17078) );
  NAND U17539 ( .A(n74), .B(a[414]), .Z(n17077) );
  AND U17540 ( .A(n17078), .B(n17077), .Z(n17131) );
  XOR U17541 ( .A(a[411]), .B(n42197), .Z(n17120) );
  NANDN U17542 ( .A(n17120), .B(n42173), .Z(n17081) );
  NANDN U17543 ( .A(n17079), .B(n42172), .Z(n17080) );
  NAND U17544 ( .A(n17081), .B(n17080), .Z(n17129) );
  NAND U17545 ( .A(b[7]), .B(a[407]), .Z(n17130) );
  XNOR U17546 ( .A(n17129), .B(n17130), .Z(n17132) );
  XOR U17547 ( .A(n17131), .B(n17132), .Z(n17138) );
  NANDN U17548 ( .A(n17082), .B(n42093), .Z(n17084) );
  XOR U17549 ( .A(n42134), .B(a[413]), .Z(n17123) );
  NANDN U17550 ( .A(n17123), .B(n42095), .Z(n17083) );
  NAND U17551 ( .A(n17084), .B(n17083), .Z(n17136) );
  NANDN U17552 ( .A(n17085), .B(n42231), .Z(n17087) );
  XOR U17553 ( .A(n196), .B(a[409]), .Z(n17126) );
  NANDN U17554 ( .A(n17126), .B(n42234), .Z(n17086) );
  AND U17555 ( .A(n17087), .B(n17086), .Z(n17135) );
  XNOR U17556 ( .A(n17136), .B(n17135), .Z(n17137) );
  XNOR U17557 ( .A(n17138), .B(n17137), .Z(n17142) );
  NANDN U17558 ( .A(n17089), .B(n17088), .Z(n17093) );
  NAND U17559 ( .A(n17091), .B(n17090), .Z(n17092) );
  AND U17560 ( .A(n17093), .B(n17092), .Z(n17141) );
  XOR U17561 ( .A(n17142), .B(n17141), .Z(n17143) );
  NANDN U17562 ( .A(n17095), .B(n17094), .Z(n17099) );
  NANDN U17563 ( .A(n17097), .B(n17096), .Z(n17098) );
  NAND U17564 ( .A(n17099), .B(n17098), .Z(n17144) );
  XOR U17565 ( .A(n17143), .B(n17144), .Z(n17111) );
  OR U17566 ( .A(n17101), .B(n17100), .Z(n17105) );
  NANDN U17567 ( .A(n17103), .B(n17102), .Z(n17104) );
  NAND U17568 ( .A(n17105), .B(n17104), .Z(n17112) );
  XNOR U17569 ( .A(n17111), .B(n17112), .Z(n17113) );
  XNOR U17570 ( .A(n17114), .B(n17113), .Z(n17147) );
  XNOR U17571 ( .A(n17147), .B(sreg[1431]), .Z(n17149) );
  NAND U17572 ( .A(n17106), .B(sreg[1430]), .Z(n17110) );
  OR U17573 ( .A(n17108), .B(n17107), .Z(n17109) );
  AND U17574 ( .A(n17110), .B(n17109), .Z(n17148) );
  XOR U17575 ( .A(n17149), .B(n17148), .Z(c[1431]) );
  NANDN U17576 ( .A(n17112), .B(n17111), .Z(n17116) );
  NAND U17577 ( .A(n17114), .B(n17113), .Z(n17115) );
  NAND U17578 ( .A(n17116), .B(n17115), .Z(n17155) );
  NAND U17579 ( .A(b[0]), .B(a[416]), .Z(n17117) );
  XNOR U17580 ( .A(b[1]), .B(n17117), .Z(n17119) );
  NAND U17581 ( .A(n74), .B(a[415]), .Z(n17118) );
  AND U17582 ( .A(n17119), .B(n17118), .Z(n17172) );
  XOR U17583 ( .A(a[412]), .B(n42197), .Z(n17161) );
  NANDN U17584 ( .A(n17161), .B(n42173), .Z(n17122) );
  NANDN U17585 ( .A(n17120), .B(n42172), .Z(n17121) );
  NAND U17586 ( .A(n17122), .B(n17121), .Z(n17170) );
  NAND U17587 ( .A(b[7]), .B(a[408]), .Z(n17171) );
  XNOR U17588 ( .A(n17170), .B(n17171), .Z(n17173) );
  XOR U17589 ( .A(n17172), .B(n17173), .Z(n17179) );
  NANDN U17590 ( .A(n17123), .B(n42093), .Z(n17125) );
  XOR U17591 ( .A(n42134), .B(a[414]), .Z(n17164) );
  NANDN U17592 ( .A(n17164), .B(n42095), .Z(n17124) );
  NAND U17593 ( .A(n17125), .B(n17124), .Z(n17177) );
  NANDN U17594 ( .A(n17126), .B(n42231), .Z(n17128) );
  XOR U17595 ( .A(n196), .B(a[410]), .Z(n17167) );
  NANDN U17596 ( .A(n17167), .B(n42234), .Z(n17127) );
  AND U17597 ( .A(n17128), .B(n17127), .Z(n17176) );
  XNOR U17598 ( .A(n17177), .B(n17176), .Z(n17178) );
  XNOR U17599 ( .A(n17179), .B(n17178), .Z(n17183) );
  NANDN U17600 ( .A(n17130), .B(n17129), .Z(n17134) );
  NAND U17601 ( .A(n17132), .B(n17131), .Z(n17133) );
  AND U17602 ( .A(n17134), .B(n17133), .Z(n17182) );
  XOR U17603 ( .A(n17183), .B(n17182), .Z(n17184) );
  NANDN U17604 ( .A(n17136), .B(n17135), .Z(n17140) );
  NANDN U17605 ( .A(n17138), .B(n17137), .Z(n17139) );
  NAND U17606 ( .A(n17140), .B(n17139), .Z(n17185) );
  XOR U17607 ( .A(n17184), .B(n17185), .Z(n17152) );
  OR U17608 ( .A(n17142), .B(n17141), .Z(n17146) );
  NANDN U17609 ( .A(n17144), .B(n17143), .Z(n17145) );
  NAND U17610 ( .A(n17146), .B(n17145), .Z(n17153) );
  XNOR U17611 ( .A(n17152), .B(n17153), .Z(n17154) );
  XNOR U17612 ( .A(n17155), .B(n17154), .Z(n17188) );
  XNOR U17613 ( .A(n17188), .B(sreg[1432]), .Z(n17190) );
  NAND U17614 ( .A(n17147), .B(sreg[1431]), .Z(n17151) );
  OR U17615 ( .A(n17149), .B(n17148), .Z(n17150) );
  AND U17616 ( .A(n17151), .B(n17150), .Z(n17189) );
  XOR U17617 ( .A(n17190), .B(n17189), .Z(c[1432]) );
  NANDN U17618 ( .A(n17153), .B(n17152), .Z(n17157) );
  NAND U17619 ( .A(n17155), .B(n17154), .Z(n17156) );
  NAND U17620 ( .A(n17157), .B(n17156), .Z(n17196) );
  NAND U17621 ( .A(b[0]), .B(a[417]), .Z(n17158) );
  XNOR U17622 ( .A(b[1]), .B(n17158), .Z(n17160) );
  NAND U17623 ( .A(n74), .B(a[416]), .Z(n17159) );
  AND U17624 ( .A(n17160), .B(n17159), .Z(n17213) );
  XOR U17625 ( .A(a[413]), .B(n42197), .Z(n17202) );
  NANDN U17626 ( .A(n17202), .B(n42173), .Z(n17163) );
  NANDN U17627 ( .A(n17161), .B(n42172), .Z(n17162) );
  NAND U17628 ( .A(n17163), .B(n17162), .Z(n17211) );
  NAND U17629 ( .A(b[7]), .B(a[409]), .Z(n17212) );
  XNOR U17630 ( .A(n17211), .B(n17212), .Z(n17214) );
  XOR U17631 ( .A(n17213), .B(n17214), .Z(n17220) );
  NANDN U17632 ( .A(n17164), .B(n42093), .Z(n17166) );
  XOR U17633 ( .A(n42134), .B(a[415]), .Z(n17205) );
  NANDN U17634 ( .A(n17205), .B(n42095), .Z(n17165) );
  NAND U17635 ( .A(n17166), .B(n17165), .Z(n17218) );
  NANDN U17636 ( .A(n17167), .B(n42231), .Z(n17169) );
  XOR U17637 ( .A(n196), .B(a[411]), .Z(n17208) );
  NANDN U17638 ( .A(n17208), .B(n42234), .Z(n17168) );
  AND U17639 ( .A(n17169), .B(n17168), .Z(n17217) );
  XNOR U17640 ( .A(n17218), .B(n17217), .Z(n17219) );
  XNOR U17641 ( .A(n17220), .B(n17219), .Z(n17224) );
  NANDN U17642 ( .A(n17171), .B(n17170), .Z(n17175) );
  NAND U17643 ( .A(n17173), .B(n17172), .Z(n17174) );
  AND U17644 ( .A(n17175), .B(n17174), .Z(n17223) );
  XOR U17645 ( .A(n17224), .B(n17223), .Z(n17225) );
  NANDN U17646 ( .A(n17177), .B(n17176), .Z(n17181) );
  NANDN U17647 ( .A(n17179), .B(n17178), .Z(n17180) );
  NAND U17648 ( .A(n17181), .B(n17180), .Z(n17226) );
  XOR U17649 ( .A(n17225), .B(n17226), .Z(n17193) );
  OR U17650 ( .A(n17183), .B(n17182), .Z(n17187) );
  NANDN U17651 ( .A(n17185), .B(n17184), .Z(n17186) );
  NAND U17652 ( .A(n17187), .B(n17186), .Z(n17194) );
  XNOR U17653 ( .A(n17193), .B(n17194), .Z(n17195) );
  XNOR U17654 ( .A(n17196), .B(n17195), .Z(n17229) );
  XNOR U17655 ( .A(n17229), .B(sreg[1433]), .Z(n17231) );
  NAND U17656 ( .A(n17188), .B(sreg[1432]), .Z(n17192) );
  OR U17657 ( .A(n17190), .B(n17189), .Z(n17191) );
  AND U17658 ( .A(n17192), .B(n17191), .Z(n17230) );
  XOR U17659 ( .A(n17231), .B(n17230), .Z(c[1433]) );
  NANDN U17660 ( .A(n17194), .B(n17193), .Z(n17198) );
  NAND U17661 ( .A(n17196), .B(n17195), .Z(n17197) );
  NAND U17662 ( .A(n17198), .B(n17197), .Z(n17237) );
  NAND U17663 ( .A(b[0]), .B(a[418]), .Z(n17199) );
  XNOR U17664 ( .A(b[1]), .B(n17199), .Z(n17201) );
  NAND U17665 ( .A(n74), .B(a[417]), .Z(n17200) );
  AND U17666 ( .A(n17201), .B(n17200), .Z(n17254) );
  XOR U17667 ( .A(a[414]), .B(n42197), .Z(n17243) );
  NANDN U17668 ( .A(n17243), .B(n42173), .Z(n17204) );
  NANDN U17669 ( .A(n17202), .B(n42172), .Z(n17203) );
  NAND U17670 ( .A(n17204), .B(n17203), .Z(n17252) );
  NAND U17671 ( .A(b[7]), .B(a[410]), .Z(n17253) );
  XNOR U17672 ( .A(n17252), .B(n17253), .Z(n17255) );
  XOR U17673 ( .A(n17254), .B(n17255), .Z(n17261) );
  NANDN U17674 ( .A(n17205), .B(n42093), .Z(n17207) );
  XOR U17675 ( .A(n42134), .B(a[416]), .Z(n17246) );
  NANDN U17676 ( .A(n17246), .B(n42095), .Z(n17206) );
  NAND U17677 ( .A(n17207), .B(n17206), .Z(n17259) );
  NANDN U17678 ( .A(n17208), .B(n42231), .Z(n17210) );
  XOR U17679 ( .A(n196), .B(a[412]), .Z(n17249) );
  NANDN U17680 ( .A(n17249), .B(n42234), .Z(n17209) );
  AND U17681 ( .A(n17210), .B(n17209), .Z(n17258) );
  XNOR U17682 ( .A(n17259), .B(n17258), .Z(n17260) );
  XNOR U17683 ( .A(n17261), .B(n17260), .Z(n17265) );
  NANDN U17684 ( .A(n17212), .B(n17211), .Z(n17216) );
  NAND U17685 ( .A(n17214), .B(n17213), .Z(n17215) );
  AND U17686 ( .A(n17216), .B(n17215), .Z(n17264) );
  XOR U17687 ( .A(n17265), .B(n17264), .Z(n17266) );
  NANDN U17688 ( .A(n17218), .B(n17217), .Z(n17222) );
  NANDN U17689 ( .A(n17220), .B(n17219), .Z(n17221) );
  NAND U17690 ( .A(n17222), .B(n17221), .Z(n17267) );
  XOR U17691 ( .A(n17266), .B(n17267), .Z(n17234) );
  OR U17692 ( .A(n17224), .B(n17223), .Z(n17228) );
  NANDN U17693 ( .A(n17226), .B(n17225), .Z(n17227) );
  NAND U17694 ( .A(n17228), .B(n17227), .Z(n17235) );
  XNOR U17695 ( .A(n17234), .B(n17235), .Z(n17236) );
  XNOR U17696 ( .A(n17237), .B(n17236), .Z(n17270) );
  XNOR U17697 ( .A(n17270), .B(sreg[1434]), .Z(n17272) );
  NAND U17698 ( .A(n17229), .B(sreg[1433]), .Z(n17233) );
  OR U17699 ( .A(n17231), .B(n17230), .Z(n17232) );
  AND U17700 ( .A(n17233), .B(n17232), .Z(n17271) );
  XOR U17701 ( .A(n17272), .B(n17271), .Z(c[1434]) );
  NANDN U17702 ( .A(n17235), .B(n17234), .Z(n17239) );
  NAND U17703 ( .A(n17237), .B(n17236), .Z(n17238) );
  NAND U17704 ( .A(n17239), .B(n17238), .Z(n17278) );
  NAND U17705 ( .A(b[0]), .B(a[419]), .Z(n17240) );
  XNOR U17706 ( .A(b[1]), .B(n17240), .Z(n17242) );
  NAND U17707 ( .A(n74), .B(a[418]), .Z(n17241) );
  AND U17708 ( .A(n17242), .B(n17241), .Z(n17295) );
  XOR U17709 ( .A(a[415]), .B(n42197), .Z(n17284) );
  NANDN U17710 ( .A(n17284), .B(n42173), .Z(n17245) );
  NANDN U17711 ( .A(n17243), .B(n42172), .Z(n17244) );
  NAND U17712 ( .A(n17245), .B(n17244), .Z(n17293) );
  NAND U17713 ( .A(b[7]), .B(a[411]), .Z(n17294) );
  XNOR U17714 ( .A(n17293), .B(n17294), .Z(n17296) );
  XOR U17715 ( .A(n17295), .B(n17296), .Z(n17302) );
  NANDN U17716 ( .A(n17246), .B(n42093), .Z(n17248) );
  XOR U17717 ( .A(n42134), .B(a[417]), .Z(n17287) );
  NANDN U17718 ( .A(n17287), .B(n42095), .Z(n17247) );
  NAND U17719 ( .A(n17248), .B(n17247), .Z(n17300) );
  NANDN U17720 ( .A(n17249), .B(n42231), .Z(n17251) );
  XOR U17721 ( .A(n196), .B(a[413]), .Z(n17290) );
  NANDN U17722 ( .A(n17290), .B(n42234), .Z(n17250) );
  AND U17723 ( .A(n17251), .B(n17250), .Z(n17299) );
  XNOR U17724 ( .A(n17300), .B(n17299), .Z(n17301) );
  XNOR U17725 ( .A(n17302), .B(n17301), .Z(n17306) );
  NANDN U17726 ( .A(n17253), .B(n17252), .Z(n17257) );
  NAND U17727 ( .A(n17255), .B(n17254), .Z(n17256) );
  AND U17728 ( .A(n17257), .B(n17256), .Z(n17305) );
  XOR U17729 ( .A(n17306), .B(n17305), .Z(n17307) );
  NANDN U17730 ( .A(n17259), .B(n17258), .Z(n17263) );
  NANDN U17731 ( .A(n17261), .B(n17260), .Z(n17262) );
  NAND U17732 ( .A(n17263), .B(n17262), .Z(n17308) );
  XOR U17733 ( .A(n17307), .B(n17308), .Z(n17275) );
  OR U17734 ( .A(n17265), .B(n17264), .Z(n17269) );
  NANDN U17735 ( .A(n17267), .B(n17266), .Z(n17268) );
  NAND U17736 ( .A(n17269), .B(n17268), .Z(n17276) );
  XNOR U17737 ( .A(n17275), .B(n17276), .Z(n17277) );
  XNOR U17738 ( .A(n17278), .B(n17277), .Z(n17311) );
  XNOR U17739 ( .A(n17311), .B(sreg[1435]), .Z(n17313) );
  NAND U17740 ( .A(n17270), .B(sreg[1434]), .Z(n17274) );
  OR U17741 ( .A(n17272), .B(n17271), .Z(n17273) );
  AND U17742 ( .A(n17274), .B(n17273), .Z(n17312) );
  XOR U17743 ( .A(n17313), .B(n17312), .Z(c[1435]) );
  NANDN U17744 ( .A(n17276), .B(n17275), .Z(n17280) );
  NAND U17745 ( .A(n17278), .B(n17277), .Z(n17279) );
  NAND U17746 ( .A(n17280), .B(n17279), .Z(n17319) );
  NAND U17747 ( .A(b[0]), .B(a[420]), .Z(n17281) );
  XNOR U17748 ( .A(b[1]), .B(n17281), .Z(n17283) );
  NAND U17749 ( .A(n75), .B(a[419]), .Z(n17282) );
  AND U17750 ( .A(n17283), .B(n17282), .Z(n17336) );
  XOR U17751 ( .A(a[416]), .B(n42197), .Z(n17325) );
  NANDN U17752 ( .A(n17325), .B(n42173), .Z(n17286) );
  NANDN U17753 ( .A(n17284), .B(n42172), .Z(n17285) );
  NAND U17754 ( .A(n17286), .B(n17285), .Z(n17334) );
  NAND U17755 ( .A(b[7]), .B(a[412]), .Z(n17335) );
  XNOR U17756 ( .A(n17334), .B(n17335), .Z(n17337) );
  XOR U17757 ( .A(n17336), .B(n17337), .Z(n17343) );
  NANDN U17758 ( .A(n17287), .B(n42093), .Z(n17289) );
  XOR U17759 ( .A(n42134), .B(a[418]), .Z(n17328) );
  NANDN U17760 ( .A(n17328), .B(n42095), .Z(n17288) );
  NAND U17761 ( .A(n17289), .B(n17288), .Z(n17341) );
  NANDN U17762 ( .A(n17290), .B(n42231), .Z(n17292) );
  XOR U17763 ( .A(n196), .B(a[414]), .Z(n17331) );
  NANDN U17764 ( .A(n17331), .B(n42234), .Z(n17291) );
  AND U17765 ( .A(n17292), .B(n17291), .Z(n17340) );
  XNOR U17766 ( .A(n17341), .B(n17340), .Z(n17342) );
  XNOR U17767 ( .A(n17343), .B(n17342), .Z(n17347) );
  NANDN U17768 ( .A(n17294), .B(n17293), .Z(n17298) );
  NAND U17769 ( .A(n17296), .B(n17295), .Z(n17297) );
  AND U17770 ( .A(n17298), .B(n17297), .Z(n17346) );
  XOR U17771 ( .A(n17347), .B(n17346), .Z(n17348) );
  NANDN U17772 ( .A(n17300), .B(n17299), .Z(n17304) );
  NANDN U17773 ( .A(n17302), .B(n17301), .Z(n17303) );
  NAND U17774 ( .A(n17304), .B(n17303), .Z(n17349) );
  XOR U17775 ( .A(n17348), .B(n17349), .Z(n17316) );
  OR U17776 ( .A(n17306), .B(n17305), .Z(n17310) );
  NANDN U17777 ( .A(n17308), .B(n17307), .Z(n17309) );
  NAND U17778 ( .A(n17310), .B(n17309), .Z(n17317) );
  XNOR U17779 ( .A(n17316), .B(n17317), .Z(n17318) );
  XNOR U17780 ( .A(n17319), .B(n17318), .Z(n17352) );
  XNOR U17781 ( .A(n17352), .B(sreg[1436]), .Z(n17354) );
  NAND U17782 ( .A(n17311), .B(sreg[1435]), .Z(n17315) );
  OR U17783 ( .A(n17313), .B(n17312), .Z(n17314) );
  AND U17784 ( .A(n17315), .B(n17314), .Z(n17353) );
  XOR U17785 ( .A(n17354), .B(n17353), .Z(c[1436]) );
  NANDN U17786 ( .A(n17317), .B(n17316), .Z(n17321) );
  NAND U17787 ( .A(n17319), .B(n17318), .Z(n17320) );
  NAND U17788 ( .A(n17321), .B(n17320), .Z(n17360) );
  NAND U17789 ( .A(b[0]), .B(a[421]), .Z(n17322) );
  XNOR U17790 ( .A(b[1]), .B(n17322), .Z(n17324) );
  NAND U17791 ( .A(n75), .B(a[420]), .Z(n17323) );
  AND U17792 ( .A(n17324), .B(n17323), .Z(n17377) );
  XOR U17793 ( .A(a[417]), .B(n42197), .Z(n17366) );
  NANDN U17794 ( .A(n17366), .B(n42173), .Z(n17327) );
  NANDN U17795 ( .A(n17325), .B(n42172), .Z(n17326) );
  NAND U17796 ( .A(n17327), .B(n17326), .Z(n17375) );
  NAND U17797 ( .A(b[7]), .B(a[413]), .Z(n17376) );
  XNOR U17798 ( .A(n17375), .B(n17376), .Z(n17378) );
  XOR U17799 ( .A(n17377), .B(n17378), .Z(n17384) );
  NANDN U17800 ( .A(n17328), .B(n42093), .Z(n17330) );
  XOR U17801 ( .A(n42134), .B(a[419]), .Z(n17369) );
  NANDN U17802 ( .A(n17369), .B(n42095), .Z(n17329) );
  NAND U17803 ( .A(n17330), .B(n17329), .Z(n17382) );
  NANDN U17804 ( .A(n17331), .B(n42231), .Z(n17333) );
  XOR U17805 ( .A(n196), .B(a[415]), .Z(n17372) );
  NANDN U17806 ( .A(n17372), .B(n42234), .Z(n17332) );
  AND U17807 ( .A(n17333), .B(n17332), .Z(n17381) );
  XNOR U17808 ( .A(n17382), .B(n17381), .Z(n17383) );
  XNOR U17809 ( .A(n17384), .B(n17383), .Z(n17388) );
  NANDN U17810 ( .A(n17335), .B(n17334), .Z(n17339) );
  NAND U17811 ( .A(n17337), .B(n17336), .Z(n17338) );
  AND U17812 ( .A(n17339), .B(n17338), .Z(n17387) );
  XOR U17813 ( .A(n17388), .B(n17387), .Z(n17389) );
  NANDN U17814 ( .A(n17341), .B(n17340), .Z(n17345) );
  NANDN U17815 ( .A(n17343), .B(n17342), .Z(n17344) );
  NAND U17816 ( .A(n17345), .B(n17344), .Z(n17390) );
  XOR U17817 ( .A(n17389), .B(n17390), .Z(n17357) );
  OR U17818 ( .A(n17347), .B(n17346), .Z(n17351) );
  NANDN U17819 ( .A(n17349), .B(n17348), .Z(n17350) );
  NAND U17820 ( .A(n17351), .B(n17350), .Z(n17358) );
  XNOR U17821 ( .A(n17357), .B(n17358), .Z(n17359) );
  XNOR U17822 ( .A(n17360), .B(n17359), .Z(n17393) );
  XNOR U17823 ( .A(n17393), .B(sreg[1437]), .Z(n17395) );
  NAND U17824 ( .A(n17352), .B(sreg[1436]), .Z(n17356) );
  OR U17825 ( .A(n17354), .B(n17353), .Z(n17355) );
  AND U17826 ( .A(n17356), .B(n17355), .Z(n17394) );
  XOR U17827 ( .A(n17395), .B(n17394), .Z(c[1437]) );
  NANDN U17828 ( .A(n17358), .B(n17357), .Z(n17362) );
  NAND U17829 ( .A(n17360), .B(n17359), .Z(n17361) );
  NAND U17830 ( .A(n17362), .B(n17361), .Z(n17401) );
  NAND U17831 ( .A(b[0]), .B(a[422]), .Z(n17363) );
  XNOR U17832 ( .A(b[1]), .B(n17363), .Z(n17365) );
  NAND U17833 ( .A(n75), .B(a[421]), .Z(n17364) );
  AND U17834 ( .A(n17365), .B(n17364), .Z(n17418) );
  XOR U17835 ( .A(a[418]), .B(n42197), .Z(n17407) );
  NANDN U17836 ( .A(n17407), .B(n42173), .Z(n17368) );
  NANDN U17837 ( .A(n17366), .B(n42172), .Z(n17367) );
  NAND U17838 ( .A(n17368), .B(n17367), .Z(n17416) );
  NAND U17839 ( .A(b[7]), .B(a[414]), .Z(n17417) );
  XNOR U17840 ( .A(n17416), .B(n17417), .Z(n17419) );
  XOR U17841 ( .A(n17418), .B(n17419), .Z(n17425) );
  NANDN U17842 ( .A(n17369), .B(n42093), .Z(n17371) );
  XOR U17843 ( .A(n42134), .B(a[420]), .Z(n17410) );
  NANDN U17844 ( .A(n17410), .B(n42095), .Z(n17370) );
  NAND U17845 ( .A(n17371), .B(n17370), .Z(n17423) );
  NANDN U17846 ( .A(n17372), .B(n42231), .Z(n17374) );
  XOR U17847 ( .A(n196), .B(a[416]), .Z(n17413) );
  NANDN U17848 ( .A(n17413), .B(n42234), .Z(n17373) );
  AND U17849 ( .A(n17374), .B(n17373), .Z(n17422) );
  XNOR U17850 ( .A(n17423), .B(n17422), .Z(n17424) );
  XNOR U17851 ( .A(n17425), .B(n17424), .Z(n17429) );
  NANDN U17852 ( .A(n17376), .B(n17375), .Z(n17380) );
  NAND U17853 ( .A(n17378), .B(n17377), .Z(n17379) );
  AND U17854 ( .A(n17380), .B(n17379), .Z(n17428) );
  XOR U17855 ( .A(n17429), .B(n17428), .Z(n17430) );
  NANDN U17856 ( .A(n17382), .B(n17381), .Z(n17386) );
  NANDN U17857 ( .A(n17384), .B(n17383), .Z(n17385) );
  NAND U17858 ( .A(n17386), .B(n17385), .Z(n17431) );
  XOR U17859 ( .A(n17430), .B(n17431), .Z(n17398) );
  OR U17860 ( .A(n17388), .B(n17387), .Z(n17392) );
  NANDN U17861 ( .A(n17390), .B(n17389), .Z(n17391) );
  NAND U17862 ( .A(n17392), .B(n17391), .Z(n17399) );
  XNOR U17863 ( .A(n17398), .B(n17399), .Z(n17400) );
  XNOR U17864 ( .A(n17401), .B(n17400), .Z(n17434) );
  XNOR U17865 ( .A(n17434), .B(sreg[1438]), .Z(n17436) );
  NAND U17866 ( .A(n17393), .B(sreg[1437]), .Z(n17397) );
  OR U17867 ( .A(n17395), .B(n17394), .Z(n17396) );
  AND U17868 ( .A(n17397), .B(n17396), .Z(n17435) );
  XOR U17869 ( .A(n17436), .B(n17435), .Z(c[1438]) );
  NANDN U17870 ( .A(n17399), .B(n17398), .Z(n17403) );
  NAND U17871 ( .A(n17401), .B(n17400), .Z(n17402) );
  NAND U17872 ( .A(n17403), .B(n17402), .Z(n17442) );
  NAND U17873 ( .A(b[0]), .B(a[423]), .Z(n17404) );
  XNOR U17874 ( .A(b[1]), .B(n17404), .Z(n17406) );
  NAND U17875 ( .A(n75), .B(a[422]), .Z(n17405) );
  AND U17876 ( .A(n17406), .B(n17405), .Z(n17459) );
  XOR U17877 ( .A(a[419]), .B(n42197), .Z(n17448) );
  NANDN U17878 ( .A(n17448), .B(n42173), .Z(n17409) );
  NANDN U17879 ( .A(n17407), .B(n42172), .Z(n17408) );
  NAND U17880 ( .A(n17409), .B(n17408), .Z(n17457) );
  NAND U17881 ( .A(b[7]), .B(a[415]), .Z(n17458) );
  XNOR U17882 ( .A(n17457), .B(n17458), .Z(n17460) );
  XOR U17883 ( .A(n17459), .B(n17460), .Z(n17466) );
  NANDN U17884 ( .A(n17410), .B(n42093), .Z(n17412) );
  XOR U17885 ( .A(n42134), .B(a[421]), .Z(n17451) );
  NANDN U17886 ( .A(n17451), .B(n42095), .Z(n17411) );
  NAND U17887 ( .A(n17412), .B(n17411), .Z(n17464) );
  NANDN U17888 ( .A(n17413), .B(n42231), .Z(n17415) );
  XOR U17889 ( .A(n196), .B(a[417]), .Z(n17454) );
  NANDN U17890 ( .A(n17454), .B(n42234), .Z(n17414) );
  AND U17891 ( .A(n17415), .B(n17414), .Z(n17463) );
  XNOR U17892 ( .A(n17464), .B(n17463), .Z(n17465) );
  XNOR U17893 ( .A(n17466), .B(n17465), .Z(n17470) );
  NANDN U17894 ( .A(n17417), .B(n17416), .Z(n17421) );
  NAND U17895 ( .A(n17419), .B(n17418), .Z(n17420) );
  AND U17896 ( .A(n17421), .B(n17420), .Z(n17469) );
  XOR U17897 ( .A(n17470), .B(n17469), .Z(n17471) );
  NANDN U17898 ( .A(n17423), .B(n17422), .Z(n17427) );
  NANDN U17899 ( .A(n17425), .B(n17424), .Z(n17426) );
  NAND U17900 ( .A(n17427), .B(n17426), .Z(n17472) );
  XOR U17901 ( .A(n17471), .B(n17472), .Z(n17439) );
  OR U17902 ( .A(n17429), .B(n17428), .Z(n17433) );
  NANDN U17903 ( .A(n17431), .B(n17430), .Z(n17432) );
  NAND U17904 ( .A(n17433), .B(n17432), .Z(n17440) );
  XNOR U17905 ( .A(n17439), .B(n17440), .Z(n17441) );
  XNOR U17906 ( .A(n17442), .B(n17441), .Z(n17475) );
  XNOR U17907 ( .A(n17475), .B(sreg[1439]), .Z(n17477) );
  NAND U17908 ( .A(n17434), .B(sreg[1438]), .Z(n17438) );
  OR U17909 ( .A(n17436), .B(n17435), .Z(n17437) );
  AND U17910 ( .A(n17438), .B(n17437), .Z(n17476) );
  XOR U17911 ( .A(n17477), .B(n17476), .Z(c[1439]) );
  NANDN U17912 ( .A(n17440), .B(n17439), .Z(n17444) );
  NAND U17913 ( .A(n17442), .B(n17441), .Z(n17443) );
  NAND U17914 ( .A(n17444), .B(n17443), .Z(n17483) );
  NAND U17915 ( .A(b[0]), .B(a[424]), .Z(n17445) );
  XNOR U17916 ( .A(b[1]), .B(n17445), .Z(n17447) );
  NAND U17917 ( .A(n75), .B(a[423]), .Z(n17446) );
  AND U17918 ( .A(n17447), .B(n17446), .Z(n17500) );
  XOR U17919 ( .A(a[420]), .B(n42197), .Z(n17489) );
  NANDN U17920 ( .A(n17489), .B(n42173), .Z(n17450) );
  NANDN U17921 ( .A(n17448), .B(n42172), .Z(n17449) );
  NAND U17922 ( .A(n17450), .B(n17449), .Z(n17498) );
  NAND U17923 ( .A(b[7]), .B(a[416]), .Z(n17499) );
  XNOR U17924 ( .A(n17498), .B(n17499), .Z(n17501) );
  XOR U17925 ( .A(n17500), .B(n17501), .Z(n17507) );
  NANDN U17926 ( .A(n17451), .B(n42093), .Z(n17453) );
  XOR U17927 ( .A(n42134), .B(a[422]), .Z(n17492) );
  NANDN U17928 ( .A(n17492), .B(n42095), .Z(n17452) );
  NAND U17929 ( .A(n17453), .B(n17452), .Z(n17505) );
  NANDN U17930 ( .A(n17454), .B(n42231), .Z(n17456) );
  XOR U17931 ( .A(n196), .B(a[418]), .Z(n17495) );
  NANDN U17932 ( .A(n17495), .B(n42234), .Z(n17455) );
  AND U17933 ( .A(n17456), .B(n17455), .Z(n17504) );
  XNOR U17934 ( .A(n17505), .B(n17504), .Z(n17506) );
  XNOR U17935 ( .A(n17507), .B(n17506), .Z(n17511) );
  NANDN U17936 ( .A(n17458), .B(n17457), .Z(n17462) );
  NAND U17937 ( .A(n17460), .B(n17459), .Z(n17461) );
  AND U17938 ( .A(n17462), .B(n17461), .Z(n17510) );
  XOR U17939 ( .A(n17511), .B(n17510), .Z(n17512) );
  NANDN U17940 ( .A(n17464), .B(n17463), .Z(n17468) );
  NANDN U17941 ( .A(n17466), .B(n17465), .Z(n17467) );
  NAND U17942 ( .A(n17468), .B(n17467), .Z(n17513) );
  XOR U17943 ( .A(n17512), .B(n17513), .Z(n17480) );
  OR U17944 ( .A(n17470), .B(n17469), .Z(n17474) );
  NANDN U17945 ( .A(n17472), .B(n17471), .Z(n17473) );
  NAND U17946 ( .A(n17474), .B(n17473), .Z(n17481) );
  XNOR U17947 ( .A(n17480), .B(n17481), .Z(n17482) );
  XNOR U17948 ( .A(n17483), .B(n17482), .Z(n17516) );
  XNOR U17949 ( .A(n17516), .B(sreg[1440]), .Z(n17518) );
  NAND U17950 ( .A(n17475), .B(sreg[1439]), .Z(n17479) );
  OR U17951 ( .A(n17477), .B(n17476), .Z(n17478) );
  AND U17952 ( .A(n17479), .B(n17478), .Z(n17517) );
  XOR U17953 ( .A(n17518), .B(n17517), .Z(c[1440]) );
  NANDN U17954 ( .A(n17481), .B(n17480), .Z(n17485) );
  NAND U17955 ( .A(n17483), .B(n17482), .Z(n17484) );
  NAND U17956 ( .A(n17485), .B(n17484), .Z(n17524) );
  NAND U17957 ( .A(b[0]), .B(a[425]), .Z(n17486) );
  XNOR U17958 ( .A(b[1]), .B(n17486), .Z(n17488) );
  NAND U17959 ( .A(n75), .B(a[424]), .Z(n17487) );
  AND U17960 ( .A(n17488), .B(n17487), .Z(n17541) );
  XOR U17961 ( .A(a[421]), .B(n42197), .Z(n17530) );
  NANDN U17962 ( .A(n17530), .B(n42173), .Z(n17491) );
  NANDN U17963 ( .A(n17489), .B(n42172), .Z(n17490) );
  NAND U17964 ( .A(n17491), .B(n17490), .Z(n17539) );
  NAND U17965 ( .A(b[7]), .B(a[417]), .Z(n17540) );
  XNOR U17966 ( .A(n17539), .B(n17540), .Z(n17542) );
  XOR U17967 ( .A(n17541), .B(n17542), .Z(n17548) );
  NANDN U17968 ( .A(n17492), .B(n42093), .Z(n17494) );
  XOR U17969 ( .A(n42134), .B(a[423]), .Z(n17533) );
  NANDN U17970 ( .A(n17533), .B(n42095), .Z(n17493) );
  NAND U17971 ( .A(n17494), .B(n17493), .Z(n17546) );
  NANDN U17972 ( .A(n17495), .B(n42231), .Z(n17497) );
  XOR U17973 ( .A(n197), .B(a[419]), .Z(n17536) );
  NANDN U17974 ( .A(n17536), .B(n42234), .Z(n17496) );
  AND U17975 ( .A(n17497), .B(n17496), .Z(n17545) );
  XNOR U17976 ( .A(n17546), .B(n17545), .Z(n17547) );
  XNOR U17977 ( .A(n17548), .B(n17547), .Z(n17552) );
  NANDN U17978 ( .A(n17499), .B(n17498), .Z(n17503) );
  NAND U17979 ( .A(n17501), .B(n17500), .Z(n17502) );
  AND U17980 ( .A(n17503), .B(n17502), .Z(n17551) );
  XOR U17981 ( .A(n17552), .B(n17551), .Z(n17553) );
  NANDN U17982 ( .A(n17505), .B(n17504), .Z(n17509) );
  NANDN U17983 ( .A(n17507), .B(n17506), .Z(n17508) );
  NAND U17984 ( .A(n17509), .B(n17508), .Z(n17554) );
  XOR U17985 ( .A(n17553), .B(n17554), .Z(n17521) );
  OR U17986 ( .A(n17511), .B(n17510), .Z(n17515) );
  NANDN U17987 ( .A(n17513), .B(n17512), .Z(n17514) );
  NAND U17988 ( .A(n17515), .B(n17514), .Z(n17522) );
  XNOR U17989 ( .A(n17521), .B(n17522), .Z(n17523) );
  XNOR U17990 ( .A(n17524), .B(n17523), .Z(n17557) );
  XNOR U17991 ( .A(n17557), .B(sreg[1441]), .Z(n17559) );
  NAND U17992 ( .A(n17516), .B(sreg[1440]), .Z(n17520) );
  OR U17993 ( .A(n17518), .B(n17517), .Z(n17519) );
  AND U17994 ( .A(n17520), .B(n17519), .Z(n17558) );
  XOR U17995 ( .A(n17559), .B(n17558), .Z(c[1441]) );
  NANDN U17996 ( .A(n17522), .B(n17521), .Z(n17526) );
  NAND U17997 ( .A(n17524), .B(n17523), .Z(n17525) );
  NAND U17998 ( .A(n17526), .B(n17525), .Z(n17565) );
  NAND U17999 ( .A(b[0]), .B(a[426]), .Z(n17527) );
  XNOR U18000 ( .A(b[1]), .B(n17527), .Z(n17529) );
  NAND U18001 ( .A(n75), .B(a[425]), .Z(n17528) );
  AND U18002 ( .A(n17529), .B(n17528), .Z(n17582) );
  XOR U18003 ( .A(a[422]), .B(n42197), .Z(n17571) );
  NANDN U18004 ( .A(n17571), .B(n42173), .Z(n17532) );
  NANDN U18005 ( .A(n17530), .B(n42172), .Z(n17531) );
  NAND U18006 ( .A(n17532), .B(n17531), .Z(n17580) );
  NAND U18007 ( .A(b[7]), .B(a[418]), .Z(n17581) );
  XNOR U18008 ( .A(n17580), .B(n17581), .Z(n17583) );
  XOR U18009 ( .A(n17582), .B(n17583), .Z(n17589) );
  NANDN U18010 ( .A(n17533), .B(n42093), .Z(n17535) );
  XOR U18011 ( .A(n42134), .B(a[424]), .Z(n17574) );
  NANDN U18012 ( .A(n17574), .B(n42095), .Z(n17534) );
  NAND U18013 ( .A(n17535), .B(n17534), .Z(n17587) );
  NANDN U18014 ( .A(n17536), .B(n42231), .Z(n17538) );
  XOR U18015 ( .A(n197), .B(a[420]), .Z(n17577) );
  NANDN U18016 ( .A(n17577), .B(n42234), .Z(n17537) );
  AND U18017 ( .A(n17538), .B(n17537), .Z(n17586) );
  XNOR U18018 ( .A(n17587), .B(n17586), .Z(n17588) );
  XNOR U18019 ( .A(n17589), .B(n17588), .Z(n17593) );
  NANDN U18020 ( .A(n17540), .B(n17539), .Z(n17544) );
  NAND U18021 ( .A(n17542), .B(n17541), .Z(n17543) );
  AND U18022 ( .A(n17544), .B(n17543), .Z(n17592) );
  XOR U18023 ( .A(n17593), .B(n17592), .Z(n17594) );
  NANDN U18024 ( .A(n17546), .B(n17545), .Z(n17550) );
  NANDN U18025 ( .A(n17548), .B(n17547), .Z(n17549) );
  NAND U18026 ( .A(n17550), .B(n17549), .Z(n17595) );
  XOR U18027 ( .A(n17594), .B(n17595), .Z(n17562) );
  OR U18028 ( .A(n17552), .B(n17551), .Z(n17556) );
  NANDN U18029 ( .A(n17554), .B(n17553), .Z(n17555) );
  NAND U18030 ( .A(n17556), .B(n17555), .Z(n17563) );
  XNOR U18031 ( .A(n17562), .B(n17563), .Z(n17564) );
  XNOR U18032 ( .A(n17565), .B(n17564), .Z(n17598) );
  XNOR U18033 ( .A(n17598), .B(sreg[1442]), .Z(n17600) );
  NAND U18034 ( .A(n17557), .B(sreg[1441]), .Z(n17561) );
  OR U18035 ( .A(n17559), .B(n17558), .Z(n17560) );
  AND U18036 ( .A(n17561), .B(n17560), .Z(n17599) );
  XOR U18037 ( .A(n17600), .B(n17599), .Z(c[1442]) );
  NANDN U18038 ( .A(n17563), .B(n17562), .Z(n17567) );
  NAND U18039 ( .A(n17565), .B(n17564), .Z(n17566) );
  NAND U18040 ( .A(n17567), .B(n17566), .Z(n17606) );
  NAND U18041 ( .A(b[0]), .B(a[427]), .Z(n17568) );
  XNOR U18042 ( .A(b[1]), .B(n17568), .Z(n17570) );
  NAND U18043 ( .A(n76), .B(a[426]), .Z(n17569) );
  AND U18044 ( .A(n17570), .B(n17569), .Z(n17623) );
  XOR U18045 ( .A(a[423]), .B(n42197), .Z(n17612) );
  NANDN U18046 ( .A(n17612), .B(n42173), .Z(n17573) );
  NANDN U18047 ( .A(n17571), .B(n42172), .Z(n17572) );
  NAND U18048 ( .A(n17573), .B(n17572), .Z(n17621) );
  NAND U18049 ( .A(b[7]), .B(a[419]), .Z(n17622) );
  XNOR U18050 ( .A(n17621), .B(n17622), .Z(n17624) );
  XOR U18051 ( .A(n17623), .B(n17624), .Z(n17630) );
  NANDN U18052 ( .A(n17574), .B(n42093), .Z(n17576) );
  XOR U18053 ( .A(n42134), .B(a[425]), .Z(n17615) );
  NANDN U18054 ( .A(n17615), .B(n42095), .Z(n17575) );
  NAND U18055 ( .A(n17576), .B(n17575), .Z(n17628) );
  NANDN U18056 ( .A(n17577), .B(n42231), .Z(n17579) );
  XOR U18057 ( .A(n197), .B(a[421]), .Z(n17618) );
  NANDN U18058 ( .A(n17618), .B(n42234), .Z(n17578) );
  AND U18059 ( .A(n17579), .B(n17578), .Z(n17627) );
  XNOR U18060 ( .A(n17628), .B(n17627), .Z(n17629) );
  XNOR U18061 ( .A(n17630), .B(n17629), .Z(n17634) );
  NANDN U18062 ( .A(n17581), .B(n17580), .Z(n17585) );
  NAND U18063 ( .A(n17583), .B(n17582), .Z(n17584) );
  AND U18064 ( .A(n17585), .B(n17584), .Z(n17633) );
  XOR U18065 ( .A(n17634), .B(n17633), .Z(n17635) );
  NANDN U18066 ( .A(n17587), .B(n17586), .Z(n17591) );
  NANDN U18067 ( .A(n17589), .B(n17588), .Z(n17590) );
  NAND U18068 ( .A(n17591), .B(n17590), .Z(n17636) );
  XOR U18069 ( .A(n17635), .B(n17636), .Z(n17603) );
  OR U18070 ( .A(n17593), .B(n17592), .Z(n17597) );
  NANDN U18071 ( .A(n17595), .B(n17594), .Z(n17596) );
  NAND U18072 ( .A(n17597), .B(n17596), .Z(n17604) );
  XNOR U18073 ( .A(n17603), .B(n17604), .Z(n17605) );
  XNOR U18074 ( .A(n17606), .B(n17605), .Z(n17639) );
  XNOR U18075 ( .A(n17639), .B(sreg[1443]), .Z(n17641) );
  NAND U18076 ( .A(n17598), .B(sreg[1442]), .Z(n17602) );
  OR U18077 ( .A(n17600), .B(n17599), .Z(n17601) );
  AND U18078 ( .A(n17602), .B(n17601), .Z(n17640) );
  XOR U18079 ( .A(n17641), .B(n17640), .Z(c[1443]) );
  NANDN U18080 ( .A(n17604), .B(n17603), .Z(n17608) );
  NAND U18081 ( .A(n17606), .B(n17605), .Z(n17607) );
  NAND U18082 ( .A(n17608), .B(n17607), .Z(n17647) );
  NAND U18083 ( .A(b[0]), .B(a[428]), .Z(n17609) );
  XNOR U18084 ( .A(b[1]), .B(n17609), .Z(n17611) );
  NAND U18085 ( .A(n76), .B(a[427]), .Z(n17610) );
  AND U18086 ( .A(n17611), .B(n17610), .Z(n17664) );
  XOR U18087 ( .A(a[424]), .B(n42197), .Z(n17653) );
  NANDN U18088 ( .A(n17653), .B(n42173), .Z(n17614) );
  NANDN U18089 ( .A(n17612), .B(n42172), .Z(n17613) );
  NAND U18090 ( .A(n17614), .B(n17613), .Z(n17662) );
  NAND U18091 ( .A(b[7]), .B(a[420]), .Z(n17663) );
  XNOR U18092 ( .A(n17662), .B(n17663), .Z(n17665) );
  XOR U18093 ( .A(n17664), .B(n17665), .Z(n17671) );
  NANDN U18094 ( .A(n17615), .B(n42093), .Z(n17617) );
  XOR U18095 ( .A(n42134), .B(a[426]), .Z(n17656) );
  NANDN U18096 ( .A(n17656), .B(n42095), .Z(n17616) );
  NAND U18097 ( .A(n17617), .B(n17616), .Z(n17669) );
  NANDN U18098 ( .A(n17618), .B(n42231), .Z(n17620) );
  XOR U18099 ( .A(n197), .B(a[422]), .Z(n17659) );
  NANDN U18100 ( .A(n17659), .B(n42234), .Z(n17619) );
  AND U18101 ( .A(n17620), .B(n17619), .Z(n17668) );
  XNOR U18102 ( .A(n17669), .B(n17668), .Z(n17670) );
  XNOR U18103 ( .A(n17671), .B(n17670), .Z(n17675) );
  NANDN U18104 ( .A(n17622), .B(n17621), .Z(n17626) );
  NAND U18105 ( .A(n17624), .B(n17623), .Z(n17625) );
  AND U18106 ( .A(n17626), .B(n17625), .Z(n17674) );
  XOR U18107 ( .A(n17675), .B(n17674), .Z(n17676) );
  NANDN U18108 ( .A(n17628), .B(n17627), .Z(n17632) );
  NANDN U18109 ( .A(n17630), .B(n17629), .Z(n17631) );
  NAND U18110 ( .A(n17632), .B(n17631), .Z(n17677) );
  XOR U18111 ( .A(n17676), .B(n17677), .Z(n17644) );
  OR U18112 ( .A(n17634), .B(n17633), .Z(n17638) );
  NANDN U18113 ( .A(n17636), .B(n17635), .Z(n17637) );
  NAND U18114 ( .A(n17638), .B(n17637), .Z(n17645) );
  XNOR U18115 ( .A(n17644), .B(n17645), .Z(n17646) );
  XNOR U18116 ( .A(n17647), .B(n17646), .Z(n17680) );
  XNOR U18117 ( .A(n17680), .B(sreg[1444]), .Z(n17682) );
  NAND U18118 ( .A(n17639), .B(sreg[1443]), .Z(n17643) );
  OR U18119 ( .A(n17641), .B(n17640), .Z(n17642) );
  AND U18120 ( .A(n17643), .B(n17642), .Z(n17681) );
  XOR U18121 ( .A(n17682), .B(n17681), .Z(c[1444]) );
  NANDN U18122 ( .A(n17645), .B(n17644), .Z(n17649) );
  NAND U18123 ( .A(n17647), .B(n17646), .Z(n17648) );
  NAND U18124 ( .A(n17649), .B(n17648), .Z(n17688) );
  NAND U18125 ( .A(b[0]), .B(a[429]), .Z(n17650) );
  XNOR U18126 ( .A(b[1]), .B(n17650), .Z(n17652) );
  NAND U18127 ( .A(n76), .B(a[428]), .Z(n17651) );
  AND U18128 ( .A(n17652), .B(n17651), .Z(n17705) );
  XOR U18129 ( .A(a[425]), .B(n42197), .Z(n17694) );
  NANDN U18130 ( .A(n17694), .B(n42173), .Z(n17655) );
  NANDN U18131 ( .A(n17653), .B(n42172), .Z(n17654) );
  NAND U18132 ( .A(n17655), .B(n17654), .Z(n17703) );
  NAND U18133 ( .A(b[7]), .B(a[421]), .Z(n17704) );
  XNOR U18134 ( .A(n17703), .B(n17704), .Z(n17706) );
  XOR U18135 ( .A(n17705), .B(n17706), .Z(n17712) );
  NANDN U18136 ( .A(n17656), .B(n42093), .Z(n17658) );
  XOR U18137 ( .A(n42134), .B(a[427]), .Z(n17697) );
  NANDN U18138 ( .A(n17697), .B(n42095), .Z(n17657) );
  NAND U18139 ( .A(n17658), .B(n17657), .Z(n17710) );
  NANDN U18140 ( .A(n17659), .B(n42231), .Z(n17661) );
  XOR U18141 ( .A(n197), .B(a[423]), .Z(n17700) );
  NANDN U18142 ( .A(n17700), .B(n42234), .Z(n17660) );
  AND U18143 ( .A(n17661), .B(n17660), .Z(n17709) );
  XNOR U18144 ( .A(n17710), .B(n17709), .Z(n17711) );
  XNOR U18145 ( .A(n17712), .B(n17711), .Z(n17716) );
  NANDN U18146 ( .A(n17663), .B(n17662), .Z(n17667) );
  NAND U18147 ( .A(n17665), .B(n17664), .Z(n17666) );
  AND U18148 ( .A(n17667), .B(n17666), .Z(n17715) );
  XOR U18149 ( .A(n17716), .B(n17715), .Z(n17717) );
  NANDN U18150 ( .A(n17669), .B(n17668), .Z(n17673) );
  NANDN U18151 ( .A(n17671), .B(n17670), .Z(n17672) );
  NAND U18152 ( .A(n17673), .B(n17672), .Z(n17718) );
  XOR U18153 ( .A(n17717), .B(n17718), .Z(n17685) );
  OR U18154 ( .A(n17675), .B(n17674), .Z(n17679) );
  NANDN U18155 ( .A(n17677), .B(n17676), .Z(n17678) );
  NAND U18156 ( .A(n17679), .B(n17678), .Z(n17686) );
  XNOR U18157 ( .A(n17685), .B(n17686), .Z(n17687) );
  XNOR U18158 ( .A(n17688), .B(n17687), .Z(n17721) );
  XNOR U18159 ( .A(n17721), .B(sreg[1445]), .Z(n17723) );
  NAND U18160 ( .A(n17680), .B(sreg[1444]), .Z(n17684) );
  OR U18161 ( .A(n17682), .B(n17681), .Z(n17683) );
  AND U18162 ( .A(n17684), .B(n17683), .Z(n17722) );
  XOR U18163 ( .A(n17723), .B(n17722), .Z(c[1445]) );
  NANDN U18164 ( .A(n17686), .B(n17685), .Z(n17690) );
  NAND U18165 ( .A(n17688), .B(n17687), .Z(n17689) );
  NAND U18166 ( .A(n17690), .B(n17689), .Z(n17729) );
  NAND U18167 ( .A(b[0]), .B(a[430]), .Z(n17691) );
  XNOR U18168 ( .A(b[1]), .B(n17691), .Z(n17693) );
  NAND U18169 ( .A(n76), .B(a[429]), .Z(n17692) );
  AND U18170 ( .A(n17693), .B(n17692), .Z(n17746) );
  XOR U18171 ( .A(a[426]), .B(n42197), .Z(n17735) );
  NANDN U18172 ( .A(n17735), .B(n42173), .Z(n17696) );
  NANDN U18173 ( .A(n17694), .B(n42172), .Z(n17695) );
  NAND U18174 ( .A(n17696), .B(n17695), .Z(n17744) );
  NAND U18175 ( .A(b[7]), .B(a[422]), .Z(n17745) );
  XNOR U18176 ( .A(n17744), .B(n17745), .Z(n17747) );
  XOR U18177 ( .A(n17746), .B(n17747), .Z(n17753) );
  NANDN U18178 ( .A(n17697), .B(n42093), .Z(n17699) );
  XOR U18179 ( .A(n42134), .B(a[428]), .Z(n17738) );
  NANDN U18180 ( .A(n17738), .B(n42095), .Z(n17698) );
  NAND U18181 ( .A(n17699), .B(n17698), .Z(n17751) );
  NANDN U18182 ( .A(n17700), .B(n42231), .Z(n17702) );
  XOR U18183 ( .A(n197), .B(a[424]), .Z(n17741) );
  NANDN U18184 ( .A(n17741), .B(n42234), .Z(n17701) );
  AND U18185 ( .A(n17702), .B(n17701), .Z(n17750) );
  XNOR U18186 ( .A(n17751), .B(n17750), .Z(n17752) );
  XNOR U18187 ( .A(n17753), .B(n17752), .Z(n17757) );
  NANDN U18188 ( .A(n17704), .B(n17703), .Z(n17708) );
  NAND U18189 ( .A(n17706), .B(n17705), .Z(n17707) );
  AND U18190 ( .A(n17708), .B(n17707), .Z(n17756) );
  XOR U18191 ( .A(n17757), .B(n17756), .Z(n17758) );
  NANDN U18192 ( .A(n17710), .B(n17709), .Z(n17714) );
  NANDN U18193 ( .A(n17712), .B(n17711), .Z(n17713) );
  NAND U18194 ( .A(n17714), .B(n17713), .Z(n17759) );
  XOR U18195 ( .A(n17758), .B(n17759), .Z(n17726) );
  OR U18196 ( .A(n17716), .B(n17715), .Z(n17720) );
  NANDN U18197 ( .A(n17718), .B(n17717), .Z(n17719) );
  NAND U18198 ( .A(n17720), .B(n17719), .Z(n17727) );
  XNOR U18199 ( .A(n17726), .B(n17727), .Z(n17728) );
  XNOR U18200 ( .A(n17729), .B(n17728), .Z(n17762) );
  XNOR U18201 ( .A(n17762), .B(sreg[1446]), .Z(n17764) );
  NAND U18202 ( .A(n17721), .B(sreg[1445]), .Z(n17725) );
  OR U18203 ( .A(n17723), .B(n17722), .Z(n17724) );
  AND U18204 ( .A(n17725), .B(n17724), .Z(n17763) );
  XOR U18205 ( .A(n17764), .B(n17763), .Z(c[1446]) );
  NANDN U18206 ( .A(n17727), .B(n17726), .Z(n17731) );
  NAND U18207 ( .A(n17729), .B(n17728), .Z(n17730) );
  NAND U18208 ( .A(n17731), .B(n17730), .Z(n17770) );
  NAND U18209 ( .A(b[0]), .B(a[431]), .Z(n17732) );
  XNOR U18210 ( .A(b[1]), .B(n17732), .Z(n17734) );
  NAND U18211 ( .A(n76), .B(a[430]), .Z(n17733) );
  AND U18212 ( .A(n17734), .B(n17733), .Z(n17787) );
  XOR U18213 ( .A(a[427]), .B(n42197), .Z(n17776) );
  NANDN U18214 ( .A(n17776), .B(n42173), .Z(n17737) );
  NANDN U18215 ( .A(n17735), .B(n42172), .Z(n17736) );
  NAND U18216 ( .A(n17737), .B(n17736), .Z(n17785) );
  NAND U18217 ( .A(b[7]), .B(a[423]), .Z(n17786) );
  XNOR U18218 ( .A(n17785), .B(n17786), .Z(n17788) );
  XOR U18219 ( .A(n17787), .B(n17788), .Z(n17794) );
  NANDN U18220 ( .A(n17738), .B(n42093), .Z(n17740) );
  XOR U18221 ( .A(n42134), .B(a[429]), .Z(n17779) );
  NANDN U18222 ( .A(n17779), .B(n42095), .Z(n17739) );
  NAND U18223 ( .A(n17740), .B(n17739), .Z(n17792) );
  NANDN U18224 ( .A(n17741), .B(n42231), .Z(n17743) );
  XOR U18225 ( .A(n197), .B(a[425]), .Z(n17782) );
  NANDN U18226 ( .A(n17782), .B(n42234), .Z(n17742) );
  AND U18227 ( .A(n17743), .B(n17742), .Z(n17791) );
  XNOR U18228 ( .A(n17792), .B(n17791), .Z(n17793) );
  XNOR U18229 ( .A(n17794), .B(n17793), .Z(n17798) );
  NANDN U18230 ( .A(n17745), .B(n17744), .Z(n17749) );
  NAND U18231 ( .A(n17747), .B(n17746), .Z(n17748) );
  AND U18232 ( .A(n17749), .B(n17748), .Z(n17797) );
  XOR U18233 ( .A(n17798), .B(n17797), .Z(n17799) );
  NANDN U18234 ( .A(n17751), .B(n17750), .Z(n17755) );
  NANDN U18235 ( .A(n17753), .B(n17752), .Z(n17754) );
  NAND U18236 ( .A(n17755), .B(n17754), .Z(n17800) );
  XOR U18237 ( .A(n17799), .B(n17800), .Z(n17767) );
  OR U18238 ( .A(n17757), .B(n17756), .Z(n17761) );
  NANDN U18239 ( .A(n17759), .B(n17758), .Z(n17760) );
  NAND U18240 ( .A(n17761), .B(n17760), .Z(n17768) );
  XNOR U18241 ( .A(n17767), .B(n17768), .Z(n17769) );
  XNOR U18242 ( .A(n17770), .B(n17769), .Z(n17803) );
  XNOR U18243 ( .A(n17803), .B(sreg[1447]), .Z(n17805) );
  NAND U18244 ( .A(n17762), .B(sreg[1446]), .Z(n17766) );
  OR U18245 ( .A(n17764), .B(n17763), .Z(n17765) );
  AND U18246 ( .A(n17766), .B(n17765), .Z(n17804) );
  XOR U18247 ( .A(n17805), .B(n17804), .Z(c[1447]) );
  NANDN U18248 ( .A(n17768), .B(n17767), .Z(n17772) );
  NAND U18249 ( .A(n17770), .B(n17769), .Z(n17771) );
  NAND U18250 ( .A(n17772), .B(n17771), .Z(n17811) );
  NAND U18251 ( .A(b[0]), .B(a[432]), .Z(n17773) );
  XNOR U18252 ( .A(b[1]), .B(n17773), .Z(n17775) );
  NAND U18253 ( .A(n76), .B(a[431]), .Z(n17774) );
  AND U18254 ( .A(n17775), .B(n17774), .Z(n17828) );
  XOR U18255 ( .A(a[428]), .B(n42197), .Z(n17817) );
  NANDN U18256 ( .A(n17817), .B(n42173), .Z(n17778) );
  NANDN U18257 ( .A(n17776), .B(n42172), .Z(n17777) );
  NAND U18258 ( .A(n17778), .B(n17777), .Z(n17826) );
  NAND U18259 ( .A(b[7]), .B(a[424]), .Z(n17827) );
  XNOR U18260 ( .A(n17826), .B(n17827), .Z(n17829) );
  XOR U18261 ( .A(n17828), .B(n17829), .Z(n17835) );
  NANDN U18262 ( .A(n17779), .B(n42093), .Z(n17781) );
  XOR U18263 ( .A(n42134), .B(a[430]), .Z(n17820) );
  NANDN U18264 ( .A(n17820), .B(n42095), .Z(n17780) );
  NAND U18265 ( .A(n17781), .B(n17780), .Z(n17833) );
  NANDN U18266 ( .A(n17782), .B(n42231), .Z(n17784) );
  XOR U18267 ( .A(n197), .B(a[426]), .Z(n17823) );
  NANDN U18268 ( .A(n17823), .B(n42234), .Z(n17783) );
  AND U18269 ( .A(n17784), .B(n17783), .Z(n17832) );
  XNOR U18270 ( .A(n17833), .B(n17832), .Z(n17834) );
  XNOR U18271 ( .A(n17835), .B(n17834), .Z(n17839) );
  NANDN U18272 ( .A(n17786), .B(n17785), .Z(n17790) );
  NAND U18273 ( .A(n17788), .B(n17787), .Z(n17789) );
  AND U18274 ( .A(n17790), .B(n17789), .Z(n17838) );
  XOR U18275 ( .A(n17839), .B(n17838), .Z(n17840) );
  NANDN U18276 ( .A(n17792), .B(n17791), .Z(n17796) );
  NANDN U18277 ( .A(n17794), .B(n17793), .Z(n17795) );
  NAND U18278 ( .A(n17796), .B(n17795), .Z(n17841) );
  XOR U18279 ( .A(n17840), .B(n17841), .Z(n17808) );
  OR U18280 ( .A(n17798), .B(n17797), .Z(n17802) );
  NANDN U18281 ( .A(n17800), .B(n17799), .Z(n17801) );
  NAND U18282 ( .A(n17802), .B(n17801), .Z(n17809) );
  XNOR U18283 ( .A(n17808), .B(n17809), .Z(n17810) );
  XNOR U18284 ( .A(n17811), .B(n17810), .Z(n17844) );
  XNOR U18285 ( .A(n17844), .B(sreg[1448]), .Z(n17846) );
  NAND U18286 ( .A(n17803), .B(sreg[1447]), .Z(n17807) );
  OR U18287 ( .A(n17805), .B(n17804), .Z(n17806) );
  AND U18288 ( .A(n17807), .B(n17806), .Z(n17845) );
  XOR U18289 ( .A(n17846), .B(n17845), .Z(c[1448]) );
  NANDN U18290 ( .A(n17809), .B(n17808), .Z(n17813) );
  NAND U18291 ( .A(n17811), .B(n17810), .Z(n17812) );
  NAND U18292 ( .A(n17813), .B(n17812), .Z(n17852) );
  NAND U18293 ( .A(b[0]), .B(a[433]), .Z(n17814) );
  XNOR U18294 ( .A(b[1]), .B(n17814), .Z(n17816) );
  NAND U18295 ( .A(n76), .B(a[432]), .Z(n17815) );
  AND U18296 ( .A(n17816), .B(n17815), .Z(n17869) );
  XOR U18297 ( .A(a[429]), .B(n42197), .Z(n17858) );
  NANDN U18298 ( .A(n17858), .B(n42173), .Z(n17819) );
  NANDN U18299 ( .A(n17817), .B(n42172), .Z(n17818) );
  NAND U18300 ( .A(n17819), .B(n17818), .Z(n17867) );
  NAND U18301 ( .A(b[7]), .B(a[425]), .Z(n17868) );
  XNOR U18302 ( .A(n17867), .B(n17868), .Z(n17870) );
  XOR U18303 ( .A(n17869), .B(n17870), .Z(n17876) );
  NANDN U18304 ( .A(n17820), .B(n42093), .Z(n17822) );
  XOR U18305 ( .A(n42134), .B(a[431]), .Z(n17861) );
  NANDN U18306 ( .A(n17861), .B(n42095), .Z(n17821) );
  NAND U18307 ( .A(n17822), .B(n17821), .Z(n17874) );
  NANDN U18308 ( .A(n17823), .B(n42231), .Z(n17825) );
  XOR U18309 ( .A(n197), .B(a[427]), .Z(n17864) );
  NANDN U18310 ( .A(n17864), .B(n42234), .Z(n17824) );
  AND U18311 ( .A(n17825), .B(n17824), .Z(n17873) );
  XNOR U18312 ( .A(n17874), .B(n17873), .Z(n17875) );
  XNOR U18313 ( .A(n17876), .B(n17875), .Z(n17880) );
  NANDN U18314 ( .A(n17827), .B(n17826), .Z(n17831) );
  NAND U18315 ( .A(n17829), .B(n17828), .Z(n17830) );
  AND U18316 ( .A(n17831), .B(n17830), .Z(n17879) );
  XOR U18317 ( .A(n17880), .B(n17879), .Z(n17881) );
  NANDN U18318 ( .A(n17833), .B(n17832), .Z(n17837) );
  NANDN U18319 ( .A(n17835), .B(n17834), .Z(n17836) );
  NAND U18320 ( .A(n17837), .B(n17836), .Z(n17882) );
  XOR U18321 ( .A(n17881), .B(n17882), .Z(n17849) );
  OR U18322 ( .A(n17839), .B(n17838), .Z(n17843) );
  NANDN U18323 ( .A(n17841), .B(n17840), .Z(n17842) );
  NAND U18324 ( .A(n17843), .B(n17842), .Z(n17850) );
  XNOR U18325 ( .A(n17849), .B(n17850), .Z(n17851) );
  XNOR U18326 ( .A(n17852), .B(n17851), .Z(n17885) );
  XNOR U18327 ( .A(n17885), .B(sreg[1449]), .Z(n17887) );
  NAND U18328 ( .A(n17844), .B(sreg[1448]), .Z(n17848) );
  OR U18329 ( .A(n17846), .B(n17845), .Z(n17847) );
  AND U18330 ( .A(n17848), .B(n17847), .Z(n17886) );
  XOR U18331 ( .A(n17887), .B(n17886), .Z(c[1449]) );
  NANDN U18332 ( .A(n17850), .B(n17849), .Z(n17854) );
  NAND U18333 ( .A(n17852), .B(n17851), .Z(n17853) );
  NAND U18334 ( .A(n17854), .B(n17853), .Z(n17893) );
  NAND U18335 ( .A(b[0]), .B(a[434]), .Z(n17855) );
  XNOR U18336 ( .A(b[1]), .B(n17855), .Z(n17857) );
  NAND U18337 ( .A(n77), .B(a[433]), .Z(n17856) );
  AND U18338 ( .A(n17857), .B(n17856), .Z(n17910) );
  XOR U18339 ( .A(a[430]), .B(n42197), .Z(n17899) );
  NANDN U18340 ( .A(n17899), .B(n42173), .Z(n17860) );
  NANDN U18341 ( .A(n17858), .B(n42172), .Z(n17859) );
  NAND U18342 ( .A(n17860), .B(n17859), .Z(n17908) );
  NAND U18343 ( .A(b[7]), .B(a[426]), .Z(n17909) );
  XNOR U18344 ( .A(n17908), .B(n17909), .Z(n17911) );
  XOR U18345 ( .A(n17910), .B(n17911), .Z(n17917) );
  NANDN U18346 ( .A(n17861), .B(n42093), .Z(n17863) );
  XOR U18347 ( .A(n42134), .B(a[432]), .Z(n17902) );
  NANDN U18348 ( .A(n17902), .B(n42095), .Z(n17862) );
  NAND U18349 ( .A(n17863), .B(n17862), .Z(n17915) );
  NANDN U18350 ( .A(n17864), .B(n42231), .Z(n17866) );
  XOR U18351 ( .A(n197), .B(a[428]), .Z(n17905) );
  NANDN U18352 ( .A(n17905), .B(n42234), .Z(n17865) );
  AND U18353 ( .A(n17866), .B(n17865), .Z(n17914) );
  XNOR U18354 ( .A(n17915), .B(n17914), .Z(n17916) );
  XNOR U18355 ( .A(n17917), .B(n17916), .Z(n17921) );
  NANDN U18356 ( .A(n17868), .B(n17867), .Z(n17872) );
  NAND U18357 ( .A(n17870), .B(n17869), .Z(n17871) );
  AND U18358 ( .A(n17872), .B(n17871), .Z(n17920) );
  XOR U18359 ( .A(n17921), .B(n17920), .Z(n17922) );
  NANDN U18360 ( .A(n17874), .B(n17873), .Z(n17878) );
  NANDN U18361 ( .A(n17876), .B(n17875), .Z(n17877) );
  NAND U18362 ( .A(n17878), .B(n17877), .Z(n17923) );
  XOR U18363 ( .A(n17922), .B(n17923), .Z(n17890) );
  OR U18364 ( .A(n17880), .B(n17879), .Z(n17884) );
  NANDN U18365 ( .A(n17882), .B(n17881), .Z(n17883) );
  NAND U18366 ( .A(n17884), .B(n17883), .Z(n17891) );
  XNOR U18367 ( .A(n17890), .B(n17891), .Z(n17892) );
  XNOR U18368 ( .A(n17893), .B(n17892), .Z(n17926) );
  XNOR U18369 ( .A(n17926), .B(sreg[1450]), .Z(n17928) );
  NAND U18370 ( .A(n17885), .B(sreg[1449]), .Z(n17889) );
  OR U18371 ( .A(n17887), .B(n17886), .Z(n17888) );
  AND U18372 ( .A(n17889), .B(n17888), .Z(n17927) );
  XOR U18373 ( .A(n17928), .B(n17927), .Z(c[1450]) );
  NANDN U18374 ( .A(n17891), .B(n17890), .Z(n17895) );
  NAND U18375 ( .A(n17893), .B(n17892), .Z(n17894) );
  NAND U18376 ( .A(n17895), .B(n17894), .Z(n17934) );
  NAND U18377 ( .A(b[0]), .B(a[435]), .Z(n17896) );
  XNOR U18378 ( .A(b[1]), .B(n17896), .Z(n17898) );
  NAND U18379 ( .A(n77), .B(a[434]), .Z(n17897) );
  AND U18380 ( .A(n17898), .B(n17897), .Z(n17951) );
  XOR U18381 ( .A(a[431]), .B(n42197), .Z(n17940) );
  NANDN U18382 ( .A(n17940), .B(n42173), .Z(n17901) );
  NANDN U18383 ( .A(n17899), .B(n42172), .Z(n17900) );
  NAND U18384 ( .A(n17901), .B(n17900), .Z(n17949) );
  NAND U18385 ( .A(b[7]), .B(a[427]), .Z(n17950) );
  XNOR U18386 ( .A(n17949), .B(n17950), .Z(n17952) );
  XOR U18387 ( .A(n17951), .B(n17952), .Z(n17958) );
  NANDN U18388 ( .A(n17902), .B(n42093), .Z(n17904) );
  XOR U18389 ( .A(n42134), .B(a[433]), .Z(n17943) );
  NANDN U18390 ( .A(n17943), .B(n42095), .Z(n17903) );
  NAND U18391 ( .A(n17904), .B(n17903), .Z(n17956) );
  NANDN U18392 ( .A(n17905), .B(n42231), .Z(n17907) );
  XOR U18393 ( .A(n197), .B(a[429]), .Z(n17946) );
  NANDN U18394 ( .A(n17946), .B(n42234), .Z(n17906) );
  AND U18395 ( .A(n17907), .B(n17906), .Z(n17955) );
  XNOR U18396 ( .A(n17956), .B(n17955), .Z(n17957) );
  XNOR U18397 ( .A(n17958), .B(n17957), .Z(n17962) );
  NANDN U18398 ( .A(n17909), .B(n17908), .Z(n17913) );
  NAND U18399 ( .A(n17911), .B(n17910), .Z(n17912) );
  AND U18400 ( .A(n17913), .B(n17912), .Z(n17961) );
  XOR U18401 ( .A(n17962), .B(n17961), .Z(n17963) );
  NANDN U18402 ( .A(n17915), .B(n17914), .Z(n17919) );
  NANDN U18403 ( .A(n17917), .B(n17916), .Z(n17918) );
  NAND U18404 ( .A(n17919), .B(n17918), .Z(n17964) );
  XOR U18405 ( .A(n17963), .B(n17964), .Z(n17931) );
  OR U18406 ( .A(n17921), .B(n17920), .Z(n17925) );
  NANDN U18407 ( .A(n17923), .B(n17922), .Z(n17924) );
  NAND U18408 ( .A(n17925), .B(n17924), .Z(n17932) );
  XNOR U18409 ( .A(n17931), .B(n17932), .Z(n17933) );
  XNOR U18410 ( .A(n17934), .B(n17933), .Z(n17967) );
  XNOR U18411 ( .A(n17967), .B(sreg[1451]), .Z(n17969) );
  NAND U18412 ( .A(n17926), .B(sreg[1450]), .Z(n17930) );
  OR U18413 ( .A(n17928), .B(n17927), .Z(n17929) );
  AND U18414 ( .A(n17930), .B(n17929), .Z(n17968) );
  XOR U18415 ( .A(n17969), .B(n17968), .Z(c[1451]) );
  NANDN U18416 ( .A(n17932), .B(n17931), .Z(n17936) );
  NAND U18417 ( .A(n17934), .B(n17933), .Z(n17935) );
  NAND U18418 ( .A(n17936), .B(n17935), .Z(n17975) );
  NAND U18419 ( .A(b[0]), .B(a[436]), .Z(n17937) );
  XNOR U18420 ( .A(b[1]), .B(n17937), .Z(n17939) );
  NAND U18421 ( .A(n77), .B(a[435]), .Z(n17938) );
  AND U18422 ( .A(n17939), .B(n17938), .Z(n17992) );
  XOR U18423 ( .A(a[432]), .B(n42197), .Z(n17981) );
  NANDN U18424 ( .A(n17981), .B(n42173), .Z(n17942) );
  NANDN U18425 ( .A(n17940), .B(n42172), .Z(n17941) );
  NAND U18426 ( .A(n17942), .B(n17941), .Z(n17990) );
  NAND U18427 ( .A(b[7]), .B(a[428]), .Z(n17991) );
  XNOR U18428 ( .A(n17990), .B(n17991), .Z(n17993) );
  XOR U18429 ( .A(n17992), .B(n17993), .Z(n17999) );
  NANDN U18430 ( .A(n17943), .B(n42093), .Z(n17945) );
  XOR U18431 ( .A(n42134), .B(a[434]), .Z(n17984) );
  NANDN U18432 ( .A(n17984), .B(n42095), .Z(n17944) );
  NAND U18433 ( .A(n17945), .B(n17944), .Z(n17997) );
  NANDN U18434 ( .A(n17946), .B(n42231), .Z(n17948) );
  XOR U18435 ( .A(n197), .B(a[430]), .Z(n17987) );
  NANDN U18436 ( .A(n17987), .B(n42234), .Z(n17947) );
  AND U18437 ( .A(n17948), .B(n17947), .Z(n17996) );
  XNOR U18438 ( .A(n17997), .B(n17996), .Z(n17998) );
  XNOR U18439 ( .A(n17999), .B(n17998), .Z(n18003) );
  NANDN U18440 ( .A(n17950), .B(n17949), .Z(n17954) );
  NAND U18441 ( .A(n17952), .B(n17951), .Z(n17953) );
  AND U18442 ( .A(n17954), .B(n17953), .Z(n18002) );
  XOR U18443 ( .A(n18003), .B(n18002), .Z(n18004) );
  NANDN U18444 ( .A(n17956), .B(n17955), .Z(n17960) );
  NANDN U18445 ( .A(n17958), .B(n17957), .Z(n17959) );
  NAND U18446 ( .A(n17960), .B(n17959), .Z(n18005) );
  XOR U18447 ( .A(n18004), .B(n18005), .Z(n17972) );
  OR U18448 ( .A(n17962), .B(n17961), .Z(n17966) );
  NANDN U18449 ( .A(n17964), .B(n17963), .Z(n17965) );
  NAND U18450 ( .A(n17966), .B(n17965), .Z(n17973) );
  XNOR U18451 ( .A(n17972), .B(n17973), .Z(n17974) );
  XNOR U18452 ( .A(n17975), .B(n17974), .Z(n18008) );
  XNOR U18453 ( .A(n18008), .B(sreg[1452]), .Z(n18010) );
  NAND U18454 ( .A(n17967), .B(sreg[1451]), .Z(n17971) );
  OR U18455 ( .A(n17969), .B(n17968), .Z(n17970) );
  AND U18456 ( .A(n17971), .B(n17970), .Z(n18009) );
  XOR U18457 ( .A(n18010), .B(n18009), .Z(c[1452]) );
  NANDN U18458 ( .A(n17973), .B(n17972), .Z(n17977) );
  NAND U18459 ( .A(n17975), .B(n17974), .Z(n17976) );
  NAND U18460 ( .A(n17977), .B(n17976), .Z(n18016) );
  NAND U18461 ( .A(b[0]), .B(a[437]), .Z(n17978) );
  XNOR U18462 ( .A(b[1]), .B(n17978), .Z(n17980) );
  NAND U18463 ( .A(n77), .B(a[436]), .Z(n17979) );
  AND U18464 ( .A(n17980), .B(n17979), .Z(n18033) );
  XOR U18465 ( .A(a[433]), .B(n42197), .Z(n18022) );
  NANDN U18466 ( .A(n18022), .B(n42173), .Z(n17983) );
  NANDN U18467 ( .A(n17981), .B(n42172), .Z(n17982) );
  NAND U18468 ( .A(n17983), .B(n17982), .Z(n18031) );
  NAND U18469 ( .A(b[7]), .B(a[429]), .Z(n18032) );
  XNOR U18470 ( .A(n18031), .B(n18032), .Z(n18034) );
  XOR U18471 ( .A(n18033), .B(n18034), .Z(n18040) );
  NANDN U18472 ( .A(n17984), .B(n42093), .Z(n17986) );
  XOR U18473 ( .A(n42134), .B(a[435]), .Z(n18025) );
  NANDN U18474 ( .A(n18025), .B(n42095), .Z(n17985) );
  NAND U18475 ( .A(n17986), .B(n17985), .Z(n18038) );
  NANDN U18476 ( .A(n17987), .B(n42231), .Z(n17989) );
  XOR U18477 ( .A(n198), .B(a[431]), .Z(n18028) );
  NANDN U18478 ( .A(n18028), .B(n42234), .Z(n17988) );
  AND U18479 ( .A(n17989), .B(n17988), .Z(n18037) );
  XNOR U18480 ( .A(n18038), .B(n18037), .Z(n18039) );
  XNOR U18481 ( .A(n18040), .B(n18039), .Z(n18044) );
  NANDN U18482 ( .A(n17991), .B(n17990), .Z(n17995) );
  NAND U18483 ( .A(n17993), .B(n17992), .Z(n17994) );
  AND U18484 ( .A(n17995), .B(n17994), .Z(n18043) );
  XOR U18485 ( .A(n18044), .B(n18043), .Z(n18045) );
  NANDN U18486 ( .A(n17997), .B(n17996), .Z(n18001) );
  NANDN U18487 ( .A(n17999), .B(n17998), .Z(n18000) );
  NAND U18488 ( .A(n18001), .B(n18000), .Z(n18046) );
  XOR U18489 ( .A(n18045), .B(n18046), .Z(n18013) );
  OR U18490 ( .A(n18003), .B(n18002), .Z(n18007) );
  NANDN U18491 ( .A(n18005), .B(n18004), .Z(n18006) );
  NAND U18492 ( .A(n18007), .B(n18006), .Z(n18014) );
  XNOR U18493 ( .A(n18013), .B(n18014), .Z(n18015) );
  XNOR U18494 ( .A(n18016), .B(n18015), .Z(n18049) );
  XNOR U18495 ( .A(n18049), .B(sreg[1453]), .Z(n18051) );
  NAND U18496 ( .A(n18008), .B(sreg[1452]), .Z(n18012) );
  OR U18497 ( .A(n18010), .B(n18009), .Z(n18011) );
  AND U18498 ( .A(n18012), .B(n18011), .Z(n18050) );
  XOR U18499 ( .A(n18051), .B(n18050), .Z(c[1453]) );
  NANDN U18500 ( .A(n18014), .B(n18013), .Z(n18018) );
  NAND U18501 ( .A(n18016), .B(n18015), .Z(n18017) );
  NAND U18502 ( .A(n18018), .B(n18017), .Z(n18057) );
  NAND U18503 ( .A(b[0]), .B(a[438]), .Z(n18019) );
  XNOR U18504 ( .A(b[1]), .B(n18019), .Z(n18021) );
  NAND U18505 ( .A(n77), .B(a[437]), .Z(n18020) );
  AND U18506 ( .A(n18021), .B(n18020), .Z(n18074) );
  XOR U18507 ( .A(a[434]), .B(n42197), .Z(n18063) );
  NANDN U18508 ( .A(n18063), .B(n42173), .Z(n18024) );
  NANDN U18509 ( .A(n18022), .B(n42172), .Z(n18023) );
  NAND U18510 ( .A(n18024), .B(n18023), .Z(n18072) );
  NAND U18511 ( .A(b[7]), .B(a[430]), .Z(n18073) );
  XNOR U18512 ( .A(n18072), .B(n18073), .Z(n18075) );
  XOR U18513 ( .A(n18074), .B(n18075), .Z(n18081) );
  NANDN U18514 ( .A(n18025), .B(n42093), .Z(n18027) );
  XOR U18515 ( .A(n42134), .B(a[436]), .Z(n18066) );
  NANDN U18516 ( .A(n18066), .B(n42095), .Z(n18026) );
  NAND U18517 ( .A(n18027), .B(n18026), .Z(n18079) );
  NANDN U18518 ( .A(n18028), .B(n42231), .Z(n18030) );
  XOR U18519 ( .A(n198), .B(a[432]), .Z(n18069) );
  NANDN U18520 ( .A(n18069), .B(n42234), .Z(n18029) );
  AND U18521 ( .A(n18030), .B(n18029), .Z(n18078) );
  XNOR U18522 ( .A(n18079), .B(n18078), .Z(n18080) );
  XNOR U18523 ( .A(n18081), .B(n18080), .Z(n18085) );
  NANDN U18524 ( .A(n18032), .B(n18031), .Z(n18036) );
  NAND U18525 ( .A(n18034), .B(n18033), .Z(n18035) );
  AND U18526 ( .A(n18036), .B(n18035), .Z(n18084) );
  XOR U18527 ( .A(n18085), .B(n18084), .Z(n18086) );
  NANDN U18528 ( .A(n18038), .B(n18037), .Z(n18042) );
  NANDN U18529 ( .A(n18040), .B(n18039), .Z(n18041) );
  NAND U18530 ( .A(n18042), .B(n18041), .Z(n18087) );
  XOR U18531 ( .A(n18086), .B(n18087), .Z(n18054) );
  OR U18532 ( .A(n18044), .B(n18043), .Z(n18048) );
  NANDN U18533 ( .A(n18046), .B(n18045), .Z(n18047) );
  NAND U18534 ( .A(n18048), .B(n18047), .Z(n18055) );
  XNOR U18535 ( .A(n18054), .B(n18055), .Z(n18056) );
  XNOR U18536 ( .A(n18057), .B(n18056), .Z(n18090) );
  XNOR U18537 ( .A(n18090), .B(sreg[1454]), .Z(n18092) );
  NAND U18538 ( .A(n18049), .B(sreg[1453]), .Z(n18053) );
  OR U18539 ( .A(n18051), .B(n18050), .Z(n18052) );
  AND U18540 ( .A(n18053), .B(n18052), .Z(n18091) );
  XOR U18541 ( .A(n18092), .B(n18091), .Z(c[1454]) );
  NANDN U18542 ( .A(n18055), .B(n18054), .Z(n18059) );
  NAND U18543 ( .A(n18057), .B(n18056), .Z(n18058) );
  NAND U18544 ( .A(n18059), .B(n18058), .Z(n18098) );
  NAND U18545 ( .A(b[0]), .B(a[439]), .Z(n18060) );
  XNOR U18546 ( .A(b[1]), .B(n18060), .Z(n18062) );
  NAND U18547 ( .A(n77), .B(a[438]), .Z(n18061) );
  AND U18548 ( .A(n18062), .B(n18061), .Z(n18115) );
  XOR U18549 ( .A(a[435]), .B(n42197), .Z(n18104) );
  NANDN U18550 ( .A(n18104), .B(n42173), .Z(n18065) );
  NANDN U18551 ( .A(n18063), .B(n42172), .Z(n18064) );
  NAND U18552 ( .A(n18065), .B(n18064), .Z(n18113) );
  NAND U18553 ( .A(b[7]), .B(a[431]), .Z(n18114) );
  XNOR U18554 ( .A(n18113), .B(n18114), .Z(n18116) );
  XOR U18555 ( .A(n18115), .B(n18116), .Z(n18122) );
  NANDN U18556 ( .A(n18066), .B(n42093), .Z(n18068) );
  XOR U18557 ( .A(n42134), .B(a[437]), .Z(n18107) );
  NANDN U18558 ( .A(n18107), .B(n42095), .Z(n18067) );
  NAND U18559 ( .A(n18068), .B(n18067), .Z(n18120) );
  NANDN U18560 ( .A(n18069), .B(n42231), .Z(n18071) );
  XOR U18561 ( .A(n198), .B(a[433]), .Z(n18110) );
  NANDN U18562 ( .A(n18110), .B(n42234), .Z(n18070) );
  AND U18563 ( .A(n18071), .B(n18070), .Z(n18119) );
  XNOR U18564 ( .A(n18120), .B(n18119), .Z(n18121) );
  XNOR U18565 ( .A(n18122), .B(n18121), .Z(n18126) );
  NANDN U18566 ( .A(n18073), .B(n18072), .Z(n18077) );
  NAND U18567 ( .A(n18075), .B(n18074), .Z(n18076) );
  AND U18568 ( .A(n18077), .B(n18076), .Z(n18125) );
  XOR U18569 ( .A(n18126), .B(n18125), .Z(n18127) );
  NANDN U18570 ( .A(n18079), .B(n18078), .Z(n18083) );
  NANDN U18571 ( .A(n18081), .B(n18080), .Z(n18082) );
  NAND U18572 ( .A(n18083), .B(n18082), .Z(n18128) );
  XOR U18573 ( .A(n18127), .B(n18128), .Z(n18095) );
  OR U18574 ( .A(n18085), .B(n18084), .Z(n18089) );
  NANDN U18575 ( .A(n18087), .B(n18086), .Z(n18088) );
  NAND U18576 ( .A(n18089), .B(n18088), .Z(n18096) );
  XNOR U18577 ( .A(n18095), .B(n18096), .Z(n18097) );
  XNOR U18578 ( .A(n18098), .B(n18097), .Z(n18131) );
  XNOR U18579 ( .A(n18131), .B(sreg[1455]), .Z(n18133) );
  NAND U18580 ( .A(n18090), .B(sreg[1454]), .Z(n18094) );
  OR U18581 ( .A(n18092), .B(n18091), .Z(n18093) );
  AND U18582 ( .A(n18094), .B(n18093), .Z(n18132) );
  XOR U18583 ( .A(n18133), .B(n18132), .Z(c[1455]) );
  NANDN U18584 ( .A(n18096), .B(n18095), .Z(n18100) );
  NAND U18585 ( .A(n18098), .B(n18097), .Z(n18099) );
  NAND U18586 ( .A(n18100), .B(n18099), .Z(n18139) );
  NAND U18587 ( .A(b[0]), .B(a[440]), .Z(n18101) );
  XNOR U18588 ( .A(b[1]), .B(n18101), .Z(n18103) );
  NAND U18589 ( .A(n77), .B(a[439]), .Z(n18102) );
  AND U18590 ( .A(n18103), .B(n18102), .Z(n18156) );
  XOR U18591 ( .A(a[436]), .B(n42197), .Z(n18145) );
  NANDN U18592 ( .A(n18145), .B(n42173), .Z(n18106) );
  NANDN U18593 ( .A(n18104), .B(n42172), .Z(n18105) );
  NAND U18594 ( .A(n18106), .B(n18105), .Z(n18154) );
  NAND U18595 ( .A(b[7]), .B(a[432]), .Z(n18155) );
  XNOR U18596 ( .A(n18154), .B(n18155), .Z(n18157) );
  XOR U18597 ( .A(n18156), .B(n18157), .Z(n18163) );
  NANDN U18598 ( .A(n18107), .B(n42093), .Z(n18109) );
  XOR U18599 ( .A(n42134), .B(a[438]), .Z(n18148) );
  NANDN U18600 ( .A(n18148), .B(n42095), .Z(n18108) );
  NAND U18601 ( .A(n18109), .B(n18108), .Z(n18161) );
  NANDN U18602 ( .A(n18110), .B(n42231), .Z(n18112) );
  XOR U18603 ( .A(n198), .B(a[434]), .Z(n18151) );
  NANDN U18604 ( .A(n18151), .B(n42234), .Z(n18111) );
  AND U18605 ( .A(n18112), .B(n18111), .Z(n18160) );
  XNOR U18606 ( .A(n18161), .B(n18160), .Z(n18162) );
  XNOR U18607 ( .A(n18163), .B(n18162), .Z(n18167) );
  NANDN U18608 ( .A(n18114), .B(n18113), .Z(n18118) );
  NAND U18609 ( .A(n18116), .B(n18115), .Z(n18117) );
  AND U18610 ( .A(n18118), .B(n18117), .Z(n18166) );
  XOR U18611 ( .A(n18167), .B(n18166), .Z(n18168) );
  NANDN U18612 ( .A(n18120), .B(n18119), .Z(n18124) );
  NANDN U18613 ( .A(n18122), .B(n18121), .Z(n18123) );
  NAND U18614 ( .A(n18124), .B(n18123), .Z(n18169) );
  XOR U18615 ( .A(n18168), .B(n18169), .Z(n18136) );
  OR U18616 ( .A(n18126), .B(n18125), .Z(n18130) );
  NANDN U18617 ( .A(n18128), .B(n18127), .Z(n18129) );
  NAND U18618 ( .A(n18130), .B(n18129), .Z(n18137) );
  XNOR U18619 ( .A(n18136), .B(n18137), .Z(n18138) );
  XNOR U18620 ( .A(n18139), .B(n18138), .Z(n18172) );
  XNOR U18621 ( .A(n18172), .B(sreg[1456]), .Z(n18174) );
  NAND U18622 ( .A(n18131), .B(sreg[1455]), .Z(n18135) );
  OR U18623 ( .A(n18133), .B(n18132), .Z(n18134) );
  AND U18624 ( .A(n18135), .B(n18134), .Z(n18173) );
  XOR U18625 ( .A(n18174), .B(n18173), .Z(c[1456]) );
  NANDN U18626 ( .A(n18137), .B(n18136), .Z(n18141) );
  NAND U18627 ( .A(n18139), .B(n18138), .Z(n18140) );
  NAND U18628 ( .A(n18141), .B(n18140), .Z(n18180) );
  NAND U18629 ( .A(b[0]), .B(a[441]), .Z(n18142) );
  XNOR U18630 ( .A(b[1]), .B(n18142), .Z(n18144) );
  NAND U18631 ( .A(n78), .B(a[440]), .Z(n18143) );
  AND U18632 ( .A(n18144), .B(n18143), .Z(n18197) );
  XOR U18633 ( .A(a[437]), .B(n42197), .Z(n18186) );
  NANDN U18634 ( .A(n18186), .B(n42173), .Z(n18147) );
  NANDN U18635 ( .A(n18145), .B(n42172), .Z(n18146) );
  NAND U18636 ( .A(n18147), .B(n18146), .Z(n18195) );
  NAND U18637 ( .A(b[7]), .B(a[433]), .Z(n18196) );
  XNOR U18638 ( .A(n18195), .B(n18196), .Z(n18198) );
  XOR U18639 ( .A(n18197), .B(n18198), .Z(n18204) );
  NANDN U18640 ( .A(n18148), .B(n42093), .Z(n18150) );
  XOR U18641 ( .A(n42134), .B(a[439]), .Z(n18189) );
  NANDN U18642 ( .A(n18189), .B(n42095), .Z(n18149) );
  NAND U18643 ( .A(n18150), .B(n18149), .Z(n18202) );
  NANDN U18644 ( .A(n18151), .B(n42231), .Z(n18153) );
  XOR U18645 ( .A(n198), .B(a[435]), .Z(n18192) );
  NANDN U18646 ( .A(n18192), .B(n42234), .Z(n18152) );
  AND U18647 ( .A(n18153), .B(n18152), .Z(n18201) );
  XNOR U18648 ( .A(n18202), .B(n18201), .Z(n18203) );
  XNOR U18649 ( .A(n18204), .B(n18203), .Z(n18208) );
  NANDN U18650 ( .A(n18155), .B(n18154), .Z(n18159) );
  NAND U18651 ( .A(n18157), .B(n18156), .Z(n18158) );
  AND U18652 ( .A(n18159), .B(n18158), .Z(n18207) );
  XOR U18653 ( .A(n18208), .B(n18207), .Z(n18209) );
  NANDN U18654 ( .A(n18161), .B(n18160), .Z(n18165) );
  NANDN U18655 ( .A(n18163), .B(n18162), .Z(n18164) );
  NAND U18656 ( .A(n18165), .B(n18164), .Z(n18210) );
  XOR U18657 ( .A(n18209), .B(n18210), .Z(n18177) );
  OR U18658 ( .A(n18167), .B(n18166), .Z(n18171) );
  NANDN U18659 ( .A(n18169), .B(n18168), .Z(n18170) );
  NAND U18660 ( .A(n18171), .B(n18170), .Z(n18178) );
  XNOR U18661 ( .A(n18177), .B(n18178), .Z(n18179) );
  XNOR U18662 ( .A(n18180), .B(n18179), .Z(n18213) );
  XNOR U18663 ( .A(n18213), .B(sreg[1457]), .Z(n18215) );
  NAND U18664 ( .A(n18172), .B(sreg[1456]), .Z(n18176) );
  OR U18665 ( .A(n18174), .B(n18173), .Z(n18175) );
  AND U18666 ( .A(n18176), .B(n18175), .Z(n18214) );
  XOR U18667 ( .A(n18215), .B(n18214), .Z(c[1457]) );
  NANDN U18668 ( .A(n18178), .B(n18177), .Z(n18182) );
  NAND U18669 ( .A(n18180), .B(n18179), .Z(n18181) );
  NAND U18670 ( .A(n18182), .B(n18181), .Z(n18221) );
  NAND U18671 ( .A(b[0]), .B(a[442]), .Z(n18183) );
  XNOR U18672 ( .A(b[1]), .B(n18183), .Z(n18185) );
  NAND U18673 ( .A(n78), .B(a[441]), .Z(n18184) );
  AND U18674 ( .A(n18185), .B(n18184), .Z(n18238) );
  XOR U18675 ( .A(a[438]), .B(n42197), .Z(n18227) );
  NANDN U18676 ( .A(n18227), .B(n42173), .Z(n18188) );
  NANDN U18677 ( .A(n18186), .B(n42172), .Z(n18187) );
  NAND U18678 ( .A(n18188), .B(n18187), .Z(n18236) );
  NAND U18679 ( .A(b[7]), .B(a[434]), .Z(n18237) );
  XNOR U18680 ( .A(n18236), .B(n18237), .Z(n18239) );
  XOR U18681 ( .A(n18238), .B(n18239), .Z(n18245) );
  NANDN U18682 ( .A(n18189), .B(n42093), .Z(n18191) );
  XOR U18683 ( .A(n42134), .B(a[440]), .Z(n18230) );
  NANDN U18684 ( .A(n18230), .B(n42095), .Z(n18190) );
  NAND U18685 ( .A(n18191), .B(n18190), .Z(n18243) );
  NANDN U18686 ( .A(n18192), .B(n42231), .Z(n18194) );
  XOR U18687 ( .A(n198), .B(a[436]), .Z(n18233) );
  NANDN U18688 ( .A(n18233), .B(n42234), .Z(n18193) );
  AND U18689 ( .A(n18194), .B(n18193), .Z(n18242) );
  XNOR U18690 ( .A(n18243), .B(n18242), .Z(n18244) );
  XNOR U18691 ( .A(n18245), .B(n18244), .Z(n18249) );
  NANDN U18692 ( .A(n18196), .B(n18195), .Z(n18200) );
  NAND U18693 ( .A(n18198), .B(n18197), .Z(n18199) );
  AND U18694 ( .A(n18200), .B(n18199), .Z(n18248) );
  XOR U18695 ( .A(n18249), .B(n18248), .Z(n18250) );
  NANDN U18696 ( .A(n18202), .B(n18201), .Z(n18206) );
  NANDN U18697 ( .A(n18204), .B(n18203), .Z(n18205) );
  NAND U18698 ( .A(n18206), .B(n18205), .Z(n18251) );
  XOR U18699 ( .A(n18250), .B(n18251), .Z(n18218) );
  OR U18700 ( .A(n18208), .B(n18207), .Z(n18212) );
  NANDN U18701 ( .A(n18210), .B(n18209), .Z(n18211) );
  NAND U18702 ( .A(n18212), .B(n18211), .Z(n18219) );
  XNOR U18703 ( .A(n18218), .B(n18219), .Z(n18220) );
  XNOR U18704 ( .A(n18221), .B(n18220), .Z(n18254) );
  XNOR U18705 ( .A(n18254), .B(sreg[1458]), .Z(n18256) );
  NAND U18706 ( .A(n18213), .B(sreg[1457]), .Z(n18217) );
  OR U18707 ( .A(n18215), .B(n18214), .Z(n18216) );
  AND U18708 ( .A(n18217), .B(n18216), .Z(n18255) );
  XOR U18709 ( .A(n18256), .B(n18255), .Z(c[1458]) );
  NANDN U18710 ( .A(n18219), .B(n18218), .Z(n18223) );
  NAND U18711 ( .A(n18221), .B(n18220), .Z(n18222) );
  NAND U18712 ( .A(n18223), .B(n18222), .Z(n18262) );
  NAND U18713 ( .A(b[0]), .B(a[443]), .Z(n18224) );
  XNOR U18714 ( .A(b[1]), .B(n18224), .Z(n18226) );
  NAND U18715 ( .A(n78), .B(a[442]), .Z(n18225) );
  AND U18716 ( .A(n18226), .B(n18225), .Z(n18279) );
  XOR U18717 ( .A(a[439]), .B(n42197), .Z(n18268) );
  NANDN U18718 ( .A(n18268), .B(n42173), .Z(n18229) );
  NANDN U18719 ( .A(n18227), .B(n42172), .Z(n18228) );
  NAND U18720 ( .A(n18229), .B(n18228), .Z(n18277) );
  NAND U18721 ( .A(b[7]), .B(a[435]), .Z(n18278) );
  XNOR U18722 ( .A(n18277), .B(n18278), .Z(n18280) );
  XOR U18723 ( .A(n18279), .B(n18280), .Z(n18286) );
  NANDN U18724 ( .A(n18230), .B(n42093), .Z(n18232) );
  XOR U18725 ( .A(n42134), .B(a[441]), .Z(n18271) );
  NANDN U18726 ( .A(n18271), .B(n42095), .Z(n18231) );
  NAND U18727 ( .A(n18232), .B(n18231), .Z(n18284) );
  NANDN U18728 ( .A(n18233), .B(n42231), .Z(n18235) );
  XOR U18729 ( .A(n198), .B(a[437]), .Z(n18274) );
  NANDN U18730 ( .A(n18274), .B(n42234), .Z(n18234) );
  AND U18731 ( .A(n18235), .B(n18234), .Z(n18283) );
  XNOR U18732 ( .A(n18284), .B(n18283), .Z(n18285) );
  XNOR U18733 ( .A(n18286), .B(n18285), .Z(n18290) );
  NANDN U18734 ( .A(n18237), .B(n18236), .Z(n18241) );
  NAND U18735 ( .A(n18239), .B(n18238), .Z(n18240) );
  AND U18736 ( .A(n18241), .B(n18240), .Z(n18289) );
  XOR U18737 ( .A(n18290), .B(n18289), .Z(n18291) );
  NANDN U18738 ( .A(n18243), .B(n18242), .Z(n18247) );
  NANDN U18739 ( .A(n18245), .B(n18244), .Z(n18246) );
  NAND U18740 ( .A(n18247), .B(n18246), .Z(n18292) );
  XOR U18741 ( .A(n18291), .B(n18292), .Z(n18259) );
  OR U18742 ( .A(n18249), .B(n18248), .Z(n18253) );
  NANDN U18743 ( .A(n18251), .B(n18250), .Z(n18252) );
  NAND U18744 ( .A(n18253), .B(n18252), .Z(n18260) );
  XNOR U18745 ( .A(n18259), .B(n18260), .Z(n18261) );
  XNOR U18746 ( .A(n18262), .B(n18261), .Z(n18295) );
  XNOR U18747 ( .A(n18295), .B(sreg[1459]), .Z(n18297) );
  NAND U18748 ( .A(n18254), .B(sreg[1458]), .Z(n18258) );
  OR U18749 ( .A(n18256), .B(n18255), .Z(n18257) );
  AND U18750 ( .A(n18258), .B(n18257), .Z(n18296) );
  XOR U18751 ( .A(n18297), .B(n18296), .Z(c[1459]) );
  NANDN U18752 ( .A(n18260), .B(n18259), .Z(n18264) );
  NAND U18753 ( .A(n18262), .B(n18261), .Z(n18263) );
  NAND U18754 ( .A(n18264), .B(n18263), .Z(n18303) );
  NAND U18755 ( .A(b[0]), .B(a[444]), .Z(n18265) );
  XNOR U18756 ( .A(b[1]), .B(n18265), .Z(n18267) );
  NAND U18757 ( .A(n78), .B(a[443]), .Z(n18266) );
  AND U18758 ( .A(n18267), .B(n18266), .Z(n18320) );
  XOR U18759 ( .A(a[440]), .B(n42197), .Z(n18309) );
  NANDN U18760 ( .A(n18309), .B(n42173), .Z(n18270) );
  NANDN U18761 ( .A(n18268), .B(n42172), .Z(n18269) );
  NAND U18762 ( .A(n18270), .B(n18269), .Z(n18318) );
  NAND U18763 ( .A(b[7]), .B(a[436]), .Z(n18319) );
  XNOR U18764 ( .A(n18318), .B(n18319), .Z(n18321) );
  XOR U18765 ( .A(n18320), .B(n18321), .Z(n18327) );
  NANDN U18766 ( .A(n18271), .B(n42093), .Z(n18273) );
  XOR U18767 ( .A(n42134), .B(a[442]), .Z(n18312) );
  NANDN U18768 ( .A(n18312), .B(n42095), .Z(n18272) );
  NAND U18769 ( .A(n18273), .B(n18272), .Z(n18325) );
  NANDN U18770 ( .A(n18274), .B(n42231), .Z(n18276) );
  XOR U18771 ( .A(n198), .B(a[438]), .Z(n18315) );
  NANDN U18772 ( .A(n18315), .B(n42234), .Z(n18275) );
  AND U18773 ( .A(n18276), .B(n18275), .Z(n18324) );
  XNOR U18774 ( .A(n18325), .B(n18324), .Z(n18326) );
  XNOR U18775 ( .A(n18327), .B(n18326), .Z(n18331) );
  NANDN U18776 ( .A(n18278), .B(n18277), .Z(n18282) );
  NAND U18777 ( .A(n18280), .B(n18279), .Z(n18281) );
  AND U18778 ( .A(n18282), .B(n18281), .Z(n18330) );
  XOR U18779 ( .A(n18331), .B(n18330), .Z(n18332) );
  NANDN U18780 ( .A(n18284), .B(n18283), .Z(n18288) );
  NANDN U18781 ( .A(n18286), .B(n18285), .Z(n18287) );
  NAND U18782 ( .A(n18288), .B(n18287), .Z(n18333) );
  XOR U18783 ( .A(n18332), .B(n18333), .Z(n18300) );
  OR U18784 ( .A(n18290), .B(n18289), .Z(n18294) );
  NANDN U18785 ( .A(n18292), .B(n18291), .Z(n18293) );
  NAND U18786 ( .A(n18294), .B(n18293), .Z(n18301) );
  XNOR U18787 ( .A(n18300), .B(n18301), .Z(n18302) );
  XNOR U18788 ( .A(n18303), .B(n18302), .Z(n18336) );
  XNOR U18789 ( .A(n18336), .B(sreg[1460]), .Z(n18338) );
  NAND U18790 ( .A(n18295), .B(sreg[1459]), .Z(n18299) );
  OR U18791 ( .A(n18297), .B(n18296), .Z(n18298) );
  AND U18792 ( .A(n18299), .B(n18298), .Z(n18337) );
  XOR U18793 ( .A(n18338), .B(n18337), .Z(c[1460]) );
  NANDN U18794 ( .A(n18301), .B(n18300), .Z(n18305) );
  NAND U18795 ( .A(n18303), .B(n18302), .Z(n18304) );
  NAND U18796 ( .A(n18305), .B(n18304), .Z(n18344) );
  NAND U18797 ( .A(b[0]), .B(a[445]), .Z(n18306) );
  XNOR U18798 ( .A(b[1]), .B(n18306), .Z(n18308) );
  NAND U18799 ( .A(n78), .B(a[444]), .Z(n18307) );
  AND U18800 ( .A(n18308), .B(n18307), .Z(n18361) );
  XOR U18801 ( .A(a[441]), .B(n42197), .Z(n18350) );
  NANDN U18802 ( .A(n18350), .B(n42173), .Z(n18311) );
  NANDN U18803 ( .A(n18309), .B(n42172), .Z(n18310) );
  NAND U18804 ( .A(n18311), .B(n18310), .Z(n18359) );
  NAND U18805 ( .A(b[7]), .B(a[437]), .Z(n18360) );
  XNOR U18806 ( .A(n18359), .B(n18360), .Z(n18362) );
  XOR U18807 ( .A(n18361), .B(n18362), .Z(n18368) );
  NANDN U18808 ( .A(n18312), .B(n42093), .Z(n18314) );
  XOR U18809 ( .A(n42134), .B(a[443]), .Z(n18353) );
  NANDN U18810 ( .A(n18353), .B(n42095), .Z(n18313) );
  NAND U18811 ( .A(n18314), .B(n18313), .Z(n18366) );
  NANDN U18812 ( .A(n18315), .B(n42231), .Z(n18317) );
  XOR U18813 ( .A(n198), .B(a[439]), .Z(n18356) );
  NANDN U18814 ( .A(n18356), .B(n42234), .Z(n18316) );
  AND U18815 ( .A(n18317), .B(n18316), .Z(n18365) );
  XNOR U18816 ( .A(n18366), .B(n18365), .Z(n18367) );
  XNOR U18817 ( .A(n18368), .B(n18367), .Z(n18372) );
  NANDN U18818 ( .A(n18319), .B(n18318), .Z(n18323) );
  NAND U18819 ( .A(n18321), .B(n18320), .Z(n18322) );
  AND U18820 ( .A(n18323), .B(n18322), .Z(n18371) );
  XOR U18821 ( .A(n18372), .B(n18371), .Z(n18373) );
  NANDN U18822 ( .A(n18325), .B(n18324), .Z(n18329) );
  NANDN U18823 ( .A(n18327), .B(n18326), .Z(n18328) );
  NAND U18824 ( .A(n18329), .B(n18328), .Z(n18374) );
  XOR U18825 ( .A(n18373), .B(n18374), .Z(n18341) );
  OR U18826 ( .A(n18331), .B(n18330), .Z(n18335) );
  NANDN U18827 ( .A(n18333), .B(n18332), .Z(n18334) );
  NAND U18828 ( .A(n18335), .B(n18334), .Z(n18342) );
  XNOR U18829 ( .A(n18341), .B(n18342), .Z(n18343) );
  XNOR U18830 ( .A(n18344), .B(n18343), .Z(n18377) );
  XNOR U18831 ( .A(n18377), .B(sreg[1461]), .Z(n18379) );
  NAND U18832 ( .A(n18336), .B(sreg[1460]), .Z(n18340) );
  OR U18833 ( .A(n18338), .B(n18337), .Z(n18339) );
  AND U18834 ( .A(n18340), .B(n18339), .Z(n18378) );
  XOR U18835 ( .A(n18379), .B(n18378), .Z(c[1461]) );
  NANDN U18836 ( .A(n18342), .B(n18341), .Z(n18346) );
  NAND U18837 ( .A(n18344), .B(n18343), .Z(n18345) );
  NAND U18838 ( .A(n18346), .B(n18345), .Z(n18385) );
  NAND U18839 ( .A(b[0]), .B(a[446]), .Z(n18347) );
  XNOR U18840 ( .A(b[1]), .B(n18347), .Z(n18349) );
  NAND U18841 ( .A(n78), .B(a[445]), .Z(n18348) );
  AND U18842 ( .A(n18349), .B(n18348), .Z(n18402) );
  XOR U18843 ( .A(a[442]), .B(n42197), .Z(n18391) );
  NANDN U18844 ( .A(n18391), .B(n42173), .Z(n18352) );
  NANDN U18845 ( .A(n18350), .B(n42172), .Z(n18351) );
  NAND U18846 ( .A(n18352), .B(n18351), .Z(n18400) );
  NAND U18847 ( .A(b[7]), .B(a[438]), .Z(n18401) );
  XNOR U18848 ( .A(n18400), .B(n18401), .Z(n18403) );
  XOR U18849 ( .A(n18402), .B(n18403), .Z(n18409) );
  NANDN U18850 ( .A(n18353), .B(n42093), .Z(n18355) );
  XOR U18851 ( .A(n42134), .B(a[444]), .Z(n18394) );
  NANDN U18852 ( .A(n18394), .B(n42095), .Z(n18354) );
  NAND U18853 ( .A(n18355), .B(n18354), .Z(n18407) );
  NANDN U18854 ( .A(n18356), .B(n42231), .Z(n18358) );
  XOR U18855 ( .A(n198), .B(a[440]), .Z(n18397) );
  NANDN U18856 ( .A(n18397), .B(n42234), .Z(n18357) );
  AND U18857 ( .A(n18358), .B(n18357), .Z(n18406) );
  XNOR U18858 ( .A(n18407), .B(n18406), .Z(n18408) );
  XNOR U18859 ( .A(n18409), .B(n18408), .Z(n18413) );
  NANDN U18860 ( .A(n18360), .B(n18359), .Z(n18364) );
  NAND U18861 ( .A(n18362), .B(n18361), .Z(n18363) );
  AND U18862 ( .A(n18364), .B(n18363), .Z(n18412) );
  XOR U18863 ( .A(n18413), .B(n18412), .Z(n18414) );
  NANDN U18864 ( .A(n18366), .B(n18365), .Z(n18370) );
  NANDN U18865 ( .A(n18368), .B(n18367), .Z(n18369) );
  NAND U18866 ( .A(n18370), .B(n18369), .Z(n18415) );
  XOR U18867 ( .A(n18414), .B(n18415), .Z(n18382) );
  OR U18868 ( .A(n18372), .B(n18371), .Z(n18376) );
  NANDN U18869 ( .A(n18374), .B(n18373), .Z(n18375) );
  NAND U18870 ( .A(n18376), .B(n18375), .Z(n18383) );
  XNOR U18871 ( .A(n18382), .B(n18383), .Z(n18384) );
  XNOR U18872 ( .A(n18385), .B(n18384), .Z(n18418) );
  XNOR U18873 ( .A(n18418), .B(sreg[1462]), .Z(n18420) );
  NAND U18874 ( .A(n18377), .B(sreg[1461]), .Z(n18381) );
  OR U18875 ( .A(n18379), .B(n18378), .Z(n18380) );
  AND U18876 ( .A(n18381), .B(n18380), .Z(n18419) );
  XOR U18877 ( .A(n18420), .B(n18419), .Z(c[1462]) );
  NANDN U18878 ( .A(n18383), .B(n18382), .Z(n18387) );
  NAND U18879 ( .A(n18385), .B(n18384), .Z(n18386) );
  NAND U18880 ( .A(n18387), .B(n18386), .Z(n18426) );
  NAND U18881 ( .A(b[0]), .B(a[447]), .Z(n18388) );
  XNOR U18882 ( .A(b[1]), .B(n18388), .Z(n18390) );
  NAND U18883 ( .A(n78), .B(a[446]), .Z(n18389) );
  AND U18884 ( .A(n18390), .B(n18389), .Z(n18443) );
  XOR U18885 ( .A(a[443]), .B(n42197), .Z(n18432) );
  NANDN U18886 ( .A(n18432), .B(n42173), .Z(n18393) );
  NANDN U18887 ( .A(n18391), .B(n42172), .Z(n18392) );
  NAND U18888 ( .A(n18393), .B(n18392), .Z(n18441) );
  NAND U18889 ( .A(b[7]), .B(a[439]), .Z(n18442) );
  XNOR U18890 ( .A(n18441), .B(n18442), .Z(n18444) );
  XOR U18891 ( .A(n18443), .B(n18444), .Z(n18450) );
  NANDN U18892 ( .A(n18394), .B(n42093), .Z(n18396) );
  XOR U18893 ( .A(n42134), .B(a[445]), .Z(n18435) );
  NANDN U18894 ( .A(n18435), .B(n42095), .Z(n18395) );
  NAND U18895 ( .A(n18396), .B(n18395), .Z(n18448) );
  NANDN U18896 ( .A(n18397), .B(n42231), .Z(n18399) );
  XOR U18897 ( .A(n198), .B(a[441]), .Z(n18438) );
  NANDN U18898 ( .A(n18438), .B(n42234), .Z(n18398) );
  AND U18899 ( .A(n18399), .B(n18398), .Z(n18447) );
  XNOR U18900 ( .A(n18448), .B(n18447), .Z(n18449) );
  XNOR U18901 ( .A(n18450), .B(n18449), .Z(n18454) );
  NANDN U18902 ( .A(n18401), .B(n18400), .Z(n18405) );
  NAND U18903 ( .A(n18403), .B(n18402), .Z(n18404) );
  AND U18904 ( .A(n18405), .B(n18404), .Z(n18453) );
  XOR U18905 ( .A(n18454), .B(n18453), .Z(n18455) );
  NANDN U18906 ( .A(n18407), .B(n18406), .Z(n18411) );
  NANDN U18907 ( .A(n18409), .B(n18408), .Z(n18410) );
  NAND U18908 ( .A(n18411), .B(n18410), .Z(n18456) );
  XOR U18909 ( .A(n18455), .B(n18456), .Z(n18423) );
  OR U18910 ( .A(n18413), .B(n18412), .Z(n18417) );
  NANDN U18911 ( .A(n18415), .B(n18414), .Z(n18416) );
  NAND U18912 ( .A(n18417), .B(n18416), .Z(n18424) );
  XNOR U18913 ( .A(n18423), .B(n18424), .Z(n18425) );
  XNOR U18914 ( .A(n18426), .B(n18425), .Z(n18459) );
  XNOR U18915 ( .A(n18459), .B(sreg[1463]), .Z(n18461) );
  NAND U18916 ( .A(n18418), .B(sreg[1462]), .Z(n18422) );
  OR U18917 ( .A(n18420), .B(n18419), .Z(n18421) );
  AND U18918 ( .A(n18422), .B(n18421), .Z(n18460) );
  XOR U18919 ( .A(n18461), .B(n18460), .Z(c[1463]) );
  NANDN U18920 ( .A(n18424), .B(n18423), .Z(n18428) );
  NAND U18921 ( .A(n18426), .B(n18425), .Z(n18427) );
  NAND U18922 ( .A(n18428), .B(n18427), .Z(n18467) );
  NAND U18923 ( .A(b[0]), .B(a[448]), .Z(n18429) );
  XNOR U18924 ( .A(b[1]), .B(n18429), .Z(n18431) );
  NAND U18925 ( .A(n79), .B(a[447]), .Z(n18430) );
  AND U18926 ( .A(n18431), .B(n18430), .Z(n18484) );
  XOR U18927 ( .A(a[444]), .B(n42197), .Z(n18473) );
  NANDN U18928 ( .A(n18473), .B(n42173), .Z(n18434) );
  NANDN U18929 ( .A(n18432), .B(n42172), .Z(n18433) );
  NAND U18930 ( .A(n18434), .B(n18433), .Z(n18482) );
  NAND U18931 ( .A(b[7]), .B(a[440]), .Z(n18483) );
  XNOR U18932 ( .A(n18482), .B(n18483), .Z(n18485) );
  XOR U18933 ( .A(n18484), .B(n18485), .Z(n18491) );
  NANDN U18934 ( .A(n18435), .B(n42093), .Z(n18437) );
  XOR U18935 ( .A(n42134), .B(a[446]), .Z(n18476) );
  NANDN U18936 ( .A(n18476), .B(n42095), .Z(n18436) );
  NAND U18937 ( .A(n18437), .B(n18436), .Z(n18489) );
  NANDN U18938 ( .A(n18438), .B(n42231), .Z(n18440) );
  XOR U18939 ( .A(n198), .B(a[442]), .Z(n18479) );
  NANDN U18940 ( .A(n18479), .B(n42234), .Z(n18439) );
  AND U18941 ( .A(n18440), .B(n18439), .Z(n18488) );
  XNOR U18942 ( .A(n18489), .B(n18488), .Z(n18490) );
  XNOR U18943 ( .A(n18491), .B(n18490), .Z(n18495) );
  NANDN U18944 ( .A(n18442), .B(n18441), .Z(n18446) );
  NAND U18945 ( .A(n18444), .B(n18443), .Z(n18445) );
  AND U18946 ( .A(n18446), .B(n18445), .Z(n18494) );
  XOR U18947 ( .A(n18495), .B(n18494), .Z(n18496) );
  NANDN U18948 ( .A(n18448), .B(n18447), .Z(n18452) );
  NANDN U18949 ( .A(n18450), .B(n18449), .Z(n18451) );
  NAND U18950 ( .A(n18452), .B(n18451), .Z(n18497) );
  XOR U18951 ( .A(n18496), .B(n18497), .Z(n18464) );
  OR U18952 ( .A(n18454), .B(n18453), .Z(n18458) );
  NANDN U18953 ( .A(n18456), .B(n18455), .Z(n18457) );
  NAND U18954 ( .A(n18458), .B(n18457), .Z(n18465) );
  XNOR U18955 ( .A(n18464), .B(n18465), .Z(n18466) );
  XNOR U18956 ( .A(n18467), .B(n18466), .Z(n18500) );
  XNOR U18957 ( .A(n18500), .B(sreg[1464]), .Z(n18502) );
  NAND U18958 ( .A(n18459), .B(sreg[1463]), .Z(n18463) );
  OR U18959 ( .A(n18461), .B(n18460), .Z(n18462) );
  AND U18960 ( .A(n18463), .B(n18462), .Z(n18501) );
  XOR U18961 ( .A(n18502), .B(n18501), .Z(c[1464]) );
  NANDN U18962 ( .A(n18465), .B(n18464), .Z(n18469) );
  NAND U18963 ( .A(n18467), .B(n18466), .Z(n18468) );
  NAND U18964 ( .A(n18469), .B(n18468), .Z(n18508) );
  NAND U18965 ( .A(b[0]), .B(a[449]), .Z(n18470) );
  XNOR U18966 ( .A(b[1]), .B(n18470), .Z(n18472) );
  NAND U18967 ( .A(n79), .B(a[448]), .Z(n18471) );
  AND U18968 ( .A(n18472), .B(n18471), .Z(n18525) );
  XOR U18969 ( .A(a[445]), .B(n42197), .Z(n18514) );
  NANDN U18970 ( .A(n18514), .B(n42173), .Z(n18475) );
  NANDN U18971 ( .A(n18473), .B(n42172), .Z(n18474) );
  NAND U18972 ( .A(n18475), .B(n18474), .Z(n18523) );
  NAND U18973 ( .A(b[7]), .B(a[441]), .Z(n18524) );
  XNOR U18974 ( .A(n18523), .B(n18524), .Z(n18526) );
  XOR U18975 ( .A(n18525), .B(n18526), .Z(n18532) );
  NANDN U18976 ( .A(n18476), .B(n42093), .Z(n18478) );
  XOR U18977 ( .A(n42134), .B(a[447]), .Z(n18517) );
  NANDN U18978 ( .A(n18517), .B(n42095), .Z(n18477) );
  NAND U18979 ( .A(n18478), .B(n18477), .Z(n18530) );
  NANDN U18980 ( .A(n18479), .B(n42231), .Z(n18481) );
  XOR U18981 ( .A(n199), .B(a[443]), .Z(n18520) );
  NANDN U18982 ( .A(n18520), .B(n42234), .Z(n18480) );
  AND U18983 ( .A(n18481), .B(n18480), .Z(n18529) );
  XNOR U18984 ( .A(n18530), .B(n18529), .Z(n18531) );
  XNOR U18985 ( .A(n18532), .B(n18531), .Z(n18536) );
  NANDN U18986 ( .A(n18483), .B(n18482), .Z(n18487) );
  NAND U18987 ( .A(n18485), .B(n18484), .Z(n18486) );
  AND U18988 ( .A(n18487), .B(n18486), .Z(n18535) );
  XOR U18989 ( .A(n18536), .B(n18535), .Z(n18537) );
  NANDN U18990 ( .A(n18489), .B(n18488), .Z(n18493) );
  NANDN U18991 ( .A(n18491), .B(n18490), .Z(n18492) );
  NAND U18992 ( .A(n18493), .B(n18492), .Z(n18538) );
  XOR U18993 ( .A(n18537), .B(n18538), .Z(n18505) );
  OR U18994 ( .A(n18495), .B(n18494), .Z(n18499) );
  NANDN U18995 ( .A(n18497), .B(n18496), .Z(n18498) );
  NAND U18996 ( .A(n18499), .B(n18498), .Z(n18506) );
  XNOR U18997 ( .A(n18505), .B(n18506), .Z(n18507) );
  XNOR U18998 ( .A(n18508), .B(n18507), .Z(n18541) );
  XNOR U18999 ( .A(n18541), .B(sreg[1465]), .Z(n18543) );
  NAND U19000 ( .A(n18500), .B(sreg[1464]), .Z(n18504) );
  OR U19001 ( .A(n18502), .B(n18501), .Z(n18503) );
  AND U19002 ( .A(n18504), .B(n18503), .Z(n18542) );
  XOR U19003 ( .A(n18543), .B(n18542), .Z(c[1465]) );
  NANDN U19004 ( .A(n18506), .B(n18505), .Z(n18510) );
  NAND U19005 ( .A(n18508), .B(n18507), .Z(n18509) );
  NAND U19006 ( .A(n18510), .B(n18509), .Z(n18549) );
  NAND U19007 ( .A(b[0]), .B(a[450]), .Z(n18511) );
  XNOR U19008 ( .A(b[1]), .B(n18511), .Z(n18513) );
  NAND U19009 ( .A(n79), .B(a[449]), .Z(n18512) );
  AND U19010 ( .A(n18513), .B(n18512), .Z(n18566) );
  XOR U19011 ( .A(a[446]), .B(n42197), .Z(n18555) );
  NANDN U19012 ( .A(n18555), .B(n42173), .Z(n18516) );
  NANDN U19013 ( .A(n18514), .B(n42172), .Z(n18515) );
  NAND U19014 ( .A(n18516), .B(n18515), .Z(n18564) );
  NAND U19015 ( .A(b[7]), .B(a[442]), .Z(n18565) );
  XNOR U19016 ( .A(n18564), .B(n18565), .Z(n18567) );
  XOR U19017 ( .A(n18566), .B(n18567), .Z(n18573) );
  NANDN U19018 ( .A(n18517), .B(n42093), .Z(n18519) );
  XOR U19019 ( .A(n42134), .B(a[448]), .Z(n18558) );
  NANDN U19020 ( .A(n18558), .B(n42095), .Z(n18518) );
  NAND U19021 ( .A(n18519), .B(n18518), .Z(n18571) );
  NANDN U19022 ( .A(n18520), .B(n42231), .Z(n18522) );
  XOR U19023 ( .A(n199), .B(a[444]), .Z(n18561) );
  NANDN U19024 ( .A(n18561), .B(n42234), .Z(n18521) );
  AND U19025 ( .A(n18522), .B(n18521), .Z(n18570) );
  XNOR U19026 ( .A(n18571), .B(n18570), .Z(n18572) );
  XNOR U19027 ( .A(n18573), .B(n18572), .Z(n18577) );
  NANDN U19028 ( .A(n18524), .B(n18523), .Z(n18528) );
  NAND U19029 ( .A(n18526), .B(n18525), .Z(n18527) );
  AND U19030 ( .A(n18528), .B(n18527), .Z(n18576) );
  XOR U19031 ( .A(n18577), .B(n18576), .Z(n18578) );
  NANDN U19032 ( .A(n18530), .B(n18529), .Z(n18534) );
  NANDN U19033 ( .A(n18532), .B(n18531), .Z(n18533) );
  NAND U19034 ( .A(n18534), .B(n18533), .Z(n18579) );
  XOR U19035 ( .A(n18578), .B(n18579), .Z(n18546) );
  OR U19036 ( .A(n18536), .B(n18535), .Z(n18540) );
  NANDN U19037 ( .A(n18538), .B(n18537), .Z(n18539) );
  NAND U19038 ( .A(n18540), .B(n18539), .Z(n18547) );
  XNOR U19039 ( .A(n18546), .B(n18547), .Z(n18548) );
  XNOR U19040 ( .A(n18549), .B(n18548), .Z(n18582) );
  XNOR U19041 ( .A(n18582), .B(sreg[1466]), .Z(n18584) );
  NAND U19042 ( .A(n18541), .B(sreg[1465]), .Z(n18545) );
  OR U19043 ( .A(n18543), .B(n18542), .Z(n18544) );
  AND U19044 ( .A(n18545), .B(n18544), .Z(n18583) );
  XOR U19045 ( .A(n18584), .B(n18583), .Z(c[1466]) );
  NANDN U19046 ( .A(n18547), .B(n18546), .Z(n18551) );
  NAND U19047 ( .A(n18549), .B(n18548), .Z(n18550) );
  NAND U19048 ( .A(n18551), .B(n18550), .Z(n18590) );
  NAND U19049 ( .A(b[0]), .B(a[451]), .Z(n18552) );
  XNOR U19050 ( .A(b[1]), .B(n18552), .Z(n18554) );
  NAND U19051 ( .A(n79), .B(a[450]), .Z(n18553) );
  AND U19052 ( .A(n18554), .B(n18553), .Z(n18607) );
  XOR U19053 ( .A(a[447]), .B(n42197), .Z(n18596) );
  NANDN U19054 ( .A(n18596), .B(n42173), .Z(n18557) );
  NANDN U19055 ( .A(n18555), .B(n42172), .Z(n18556) );
  NAND U19056 ( .A(n18557), .B(n18556), .Z(n18605) );
  NAND U19057 ( .A(b[7]), .B(a[443]), .Z(n18606) );
  XNOR U19058 ( .A(n18605), .B(n18606), .Z(n18608) );
  XOR U19059 ( .A(n18607), .B(n18608), .Z(n18614) );
  NANDN U19060 ( .A(n18558), .B(n42093), .Z(n18560) );
  XOR U19061 ( .A(n42134), .B(a[449]), .Z(n18599) );
  NANDN U19062 ( .A(n18599), .B(n42095), .Z(n18559) );
  NAND U19063 ( .A(n18560), .B(n18559), .Z(n18612) );
  NANDN U19064 ( .A(n18561), .B(n42231), .Z(n18563) );
  XOR U19065 ( .A(n199), .B(a[445]), .Z(n18602) );
  NANDN U19066 ( .A(n18602), .B(n42234), .Z(n18562) );
  AND U19067 ( .A(n18563), .B(n18562), .Z(n18611) );
  XNOR U19068 ( .A(n18612), .B(n18611), .Z(n18613) );
  XNOR U19069 ( .A(n18614), .B(n18613), .Z(n18618) );
  NANDN U19070 ( .A(n18565), .B(n18564), .Z(n18569) );
  NAND U19071 ( .A(n18567), .B(n18566), .Z(n18568) );
  AND U19072 ( .A(n18569), .B(n18568), .Z(n18617) );
  XOR U19073 ( .A(n18618), .B(n18617), .Z(n18619) );
  NANDN U19074 ( .A(n18571), .B(n18570), .Z(n18575) );
  NANDN U19075 ( .A(n18573), .B(n18572), .Z(n18574) );
  NAND U19076 ( .A(n18575), .B(n18574), .Z(n18620) );
  XOR U19077 ( .A(n18619), .B(n18620), .Z(n18587) );
  OR U19078 ( .A(n18577), .B(n18576), .Z(n18581) );
  NANDN U19079 ( .A(n18579), .B(n18578), .Z(n18580) );
  NAND U19080 ( .A(n18581), .B(n18580), .Z(n18588) );
  XNOR U19081 ( .A(n18587), .B(n18588), .Z(n18589) );
  XNOR U19082 ( .A(n18590), .B(n18589), .Z(n18623) );
  XNOR U19083 ( .A(n18623), .B(sreg[1467]), .Z(n18625) );
  NAND U19084 ( .A(n18582), .B(sreg[1466]), .Z(n18586) );
  OR U19085 ( .A(n18584), .B(n18583), .Z(n18585) );
  AND U19086 ( .A(n18586), .B(n18585), .Z(n18624) );
  XOR U19087 ( .A(n18625), .B(n18624), .Z(c[1467]) );
  NANDN U19088 ( .A(n18588), .B(n18587), .Z(n18592) );
  NAND U19089 ( .A(n18590), .B(n18589), .Z(n18591) );
  NAND U19090 ( .A(n18592), .B(n18591), .Z(n18631) );
  NAND U19091 ( .A(b[0]), .B(a[452]), .Z(n18593) );
  XNOR U19092 ( .A(b[1]), .B(n18593), .Z(n18595) );
  NAND U19093 ( .A(n79), .B(a[451]), .Z(n18594) );
  AND U19094 ( .A(n18595), .B(n18594), .Z(n18648) );
  XOR U19095 ( .A(a[448]), .B(n42197), .Z(n18637) );
  NANDN U19096 ( .A(n18637), .B(n42173), .Z(n18598) );
  NANDN U19097 ( .A(n18596), .B(n42172), .Z(n18597) );
  NAND U19098 ( .A(n18598), .B(n18597), .Z(n18646) );
  NAND U19099 ( .A(b[7]), .B(a[444]), .Z(n18647) );
  XNOR U19100 ( .A(n18646), .B(n18647), .Z(n18649) );
  XOR U19101 ( .A(n18648), .B(n18649), .Z(n18655) );
  NANDN U19102 ( .A(n18599), .B(n42093), .Z(n18601) );
  XOR U19103 ( .A(n42134), .B(a[450]), .Z(n18640) );
  NANDN U19104 ( .A(n18640), .B(n42095), .Z(n18600) );
  NAND U19105 ( .A(n18601), .B(n18600), .Z(n18653) );
  NANDN U19106 ( .A(n18602), .B(n42231), .Z(n18604) );
  XOR U19107 ( .A(n199), .B(a[446]), .Z(n18643) );
  NANDN U19108 ( .A(n18643), .B(n42234), .Z(n18603) );
  AND U19109 ( .A(n18604), .B(n18603), .Z(n18652) );
  XNOR U19110 ( .A(n18653), .B(n18652), .Z(n18654) );
  XNOR U19111 ( .A(n18655), .B(n18654), .Z(n18659) );
  NANDN U19112 ( .A(n18606), .B(n18605), .Z(n18610) );
  NAND U19113 ( .A(n18608), .B(n18607), .Z(n18609) );
  AND U19114 ( .A(n18610), .B(n18609), .Z(n18658) );
  XOR U19115 ( .A(n18659), .B(n18658), .Z(n18660) );
  NANDN U19116 ( .A(n18612), .B(n18611), .Z(n18616) );
  NANDN U19117 ( .A(n18614), .B(n18613), .Z(n18615) );
  NAND U19118 ( .A(n18616), .B(n18615), .Z(n18661) );
  XOR U19119 ( .A(n18660), .B(n18661), .Z(n18628) );
  OR U19120 ( .A(n18618), .B(n18617), .Z(n18622) );
  NANDN U19121 ( .A(n18620), .B(n18619), .Z(n18621) );
  NAND U19122 ( .A(n18622), .B(n18621), .Z(n18629) );
  XNOR U19123 ( .A(n18628), .B(n18629), .Z(n18630) );
  XNOR U19124 ( .A(n18631), .B(n18630), .Z(n18664) );
  XNOR U19125 ( .A(n18664), .B(sreg[1468]), .Z(n18666) );
  NAND U19126 ( .A(n18623), .B(sreg[1467]), .Z(n18627) );
  OR U19127 ( .A(n18625), .B(n18624), .Z(n18626) );
  AND U19128 ( .A(n18627), .B(n18626), .Z(n18665) );
  XOR U19129 ( .A(n18666), .B(n18665), .Z(c[1468]) );
  NANDN U19130 ( .A(n18629), .B(n18628), .Z(n18633) );
  NAND U19131 ( .A(n18631), .B(n18630), .Z(n18632) );
  NAND U19132 ( .A(n18633), .B(n18632), .Z(n18672) );
  NAND U19133 ( .A(b[0]), .B(a[453]), .Z(n18634) );
  XNOR U19134 ( .A(b[1]), .B(n18634), .Z(n18636) );
  NAND U19135 ( .A(n79), .B(a[452]), .Z(n18635) );
  AND U19136 ( .A(n18636), .B(n18635), .Z(n18689) );
  XOR U19137 ( .A(a[449]), .B(n42197), .Z(n18678) );
  NANDN U19138 ( .A(n18678), .B(n42173), .Z(n18639) );
  NANDN U19139 ( .A(n18637), .B(n42172), .Z(n18638) );
  NAND U19140 ( .A(n18639), .B(n18638), .Z(n18687) );
  NAND U19141 ( .A(b[7]), .B(a[445]), .Z(n18688) );
  XNOR U19142 ( .A(n18687), .B(n18688), .Z(n18690) );
  XOR U19143 ( .A(n18689), .B(n18690), .Z(n18696) );
  NANDN U19144 ( .A(n18640), .B(n42093), .Z(n18642) );
  XOR U19145 ( .A(n42134), .B(a[451]), .Z(n18681) );
  NANDN U19146 ( .A(n18681), .B(n42095), .Z(n18641) );
  NAND U19147 ( .A(n18642), .B(n18641), .Z(n18694) );
  NANDN U19148 ( .A(n18643), .B(n42231), .Z(n18645) );
  XOR U19149 ( .A(n199), .B(a[447]), .Z(n18684) );
  NANDN U19150 ( .A(n18684), .B(n42234), .Z(n18644) );
  AND U19151 ( .A(n18645), .B(n18644), .Z(n18693) );
  XNOR U19152 ( .A(n18694), .B(n18693), .Z(n18695) );
  XNOR U19153 ( .A(n18696), .B(n18695), .Z(n18700) );
  NANDN U19154 ( .A(n18647), .B(n18646), .Z(n18651) );
  NAND U19155 ( .A(n18649), .B(n18648), .Z(n18650) );
  AND U19156 ( .A(n18651), .B(n18650), .Z(n18699) );
  XOR U19157 ( .A(n18700), .B(n18699), .Z(n18701) );
  NANDN U19158 ( .A(n18653), .B(n18652), .Z(n18657) );
  NANDN U19159 ( .A(n18655), .B(n18654), .Z(n18656) );
  NAND U19160 ( .A(n18657), .B(n18656), .Z(n18702) );
  XOR U19161 ( .A(n18701), .B(n18702), .Z(n18669) );
  OR U19162 ( .A(n18659), .B(n18658), .Z(n18663) );
  NANDN U19163 ( .A(n18661), .B(n18660), .Z(n18662) );
  NAND U19164 ( .A(n18663), .B(n18662), .Z(n18670) );
  XNOR U19165 ( .A(n18669), .B(n18670), .Z(n18671) );
  XNOR U19166 ( .A(n18672), .B(n18671), .Z(n18705) );
  XNOR U19167 ( .A(n18705), .B(sreg[1469]), .Z(n18707) );
  NAND U19168 ( .A(n18664), .B(sreg[1468]), .Z(n18668) );
  OR U19169 ( .A(n18666), .B(n18665), .Z(n18667) );
  AND U19170 ( .A(n18668), .B(n18667), .Z(n18706) );
  XOR U19171 ( .A(n18707), .B(n18706), .Z(c[1469]) );
  NANDN U19172 ( .A(n18670), .B(n18669), .Z(n18674) );
  NAND U19173 ( .A(n18672), .B(n18671), .Z(n18673) );
  NAND U19174 ( .A(n18674), .B(n18673), .Z(n18713) );
  NAND U19175 ( .A(b[0]), .B(a[454]), .Z(n18675) );
  XNOR U19176 ( .A(b[1]), .B(n18675), .Z(n18677) );
  NAND U19177 ( .A(n79), .B(a[453]), .Z(n18676) );
  AND U19178 ( .A(n18677), .B(n18676), .Z(n18730) );
  XOR U19179 ( .A(a[450]), .B(n42197), .Z(n18719) );
  NANDN U19180 ( .A(n18719), .B(n42173), .Z(n18680) );
  NANDN U19181 ( .A(n18678), .B(n42172), .Z(n18679) );
  NAND U19182 ( .A(n18680), .B(n18679), .Z(n18728) );
  NAND U19183 ( .A(b[7]), .B(a[446]), .Z(n18729) );
  XNOR U19184 ( .A(n18728), .B(n18729), .Z(n18731) );
  XOR U19185 ( .A(n18730), .B(n18731), .Z(n18737) );
  NANDN U19186 ( .A(n18681), .B(n42093), .Z(n18683) );
  XOR U19187 ( .A(n42134), .B(a[452]), .Z(n18722) );
  NANDN U19188 ( .A(n18722), .B(n42095), .Z(n18682) );
  NAND U19189 ( .A(n18683), .B(n18682), .Z(n18735) );
  NANDN U19190 ( .A(n18684), .B(n42231), .Z(n18686) );
  XOR U19191 ( .A(n199), .B(a[448]), .Z(n18725) );
  NANDN U19192 ( .A(n18725), .B(n42234), .Z(n18685) );
  AND U19193 ( .A(n18686), .B(n18685), .Z(n18734) );
  XNOR U19194 ( .A(n18735), .B(n18734), .Z(n18736) );
  XNOR U19195 ( .A(n18737), .B(n18736), .Z(n18741) );
  NANDN U19196 ( .A(n18688), .B(n18687), .Z(n18692) );
  NAND U19197 ( .A(n18690), .B(n18689), .Z(n18691) );
  AND U19198 ( .A(n18692), .B(n18691), .Z(n18740) );
  XOR U19199 ( .A(n18741), .B(n18740), .Z(n18742) );
  NANDN U19200 ( .A(n18694), .B(n18693), .Z(n18698) );
  NANDN U19201 ( .A(n18696), .B(n18695), .Z(n18697) );
  NAND U19202 ( .A(n18698), .B(n18697), .Z(n18743) );
  XOR U19203 ( .A(n18742), .B(n18743), .Z(n18710) );
  OR U19204 ( .A(n18700), .B(n18699), .Z(n18704) );
  NANDN U19205 ( .A(n18702), .B(n18701), .Z(n18703) );
  NAND U19206 ( .A(n18704), .B(n18703), .Z(n18711) );
  XNOR U19207 ( .A(n18710), .B(n18711), .Z(n18712) );
  XNOR U19208 ( .A(n18713), .B(n18712), .Z(n18746) );
  XNOR U19209 ( .A(n18746), .B(sreg[1470]), .Z(n18748) );
  NAND U19210 ( .A(n18705), .B(sreg[1469]), .Z(n18709) );
  OR U19211 ( .A(n18707), .B(n18706), .Z(n18708) );
  AND U19212 ( .A(n18709), .B(n18708), .Z(n18747) );
  XOR U19213 ( .A(n18748), .B(n18747), .Z(c[1470]) );
  NANDN U19214 ( .A(n18711), .B(n18710), .Z(n18715) );
  NAND U19215 ( .A(n18713), .B(n18712), .Z(n18714) );
  NAND U19216 ( .A(n18715), .B(n18714), .Z(n18754) );
  NAND U19217 ( .A(b[0]), .B(a[455]), .Z(n18716) );
  XNOR U19218 ( .A(b[1]), .B(n18716), .Z(n18718) );
  NAND U19219 ( .A(n80), .B(a[454]), .Z(n18717) );
  AND U19220 ( .A(n18718), .B(n18717), .Z(n18771) );
  XOR U19221 ( .A(a[451]), .B(n42197), .Z(n18760) );
  NANDN U19222 ( .A(n18760), .B(n42173), .Z(n18721) );
  NANDN U19223 ( .A(n18719), .B(n42172), .Z(n18720) );
  NAND U19224 ( .A(n18721), .B(n18720), .Z(n18769) );
  NAND U19225 ( .A(b[7]), .B(a[447]), .Z(n18770) );
  XNOR U19226 ( .A(n18769), .B(n18770), .Z(n18772) );
  XOR U19227 ( .A(n18771), .B(n18772), .Z(n18778) );
  NANDN U19228 ( .A(n18722), .B(n42093), .Z(n18724) );
  XOR U19229 ( .A(n42134), .B(a[453]), .Z(n18763) );
  NANDN U19230 ( .A(n18763), .B(n42095), .Z(n18723) );
  NAND U19231 ( .A(n18724), .B(n18723), .Z(n18776) );
  NANDN U19232 ( .A(n18725), .B(n42231), .Z(n18727) );
  XOR U19233 ( .A(n199), .B(a[449]), .Z(n18766) );
  NANDN U19234 ( .A(n18766), .B(n42234), .Z(n18726) );
  AND U19235 ( .A(n18727), .B(n18726), .Z(n18775) );
  XNOR U19236 ( .A(n18776), .B(n18775), .Z(n18777) );
  XNOR U19237 ( .A(n18778), .B(n18777), .Z(n18782) );
  NANDN U19238 ( .A(n18729), .B(n18728), .Z(n18733) );
  NAND U19239 ( .A(n18731), .B(n18730), .Z(n18732) );
  AND U19240 ( .A(n18733), .B(n18732), .Z(n18781) );
  XOR U19241 ( .A(n18782), .B(n18781), .Z(n18783) );
  NANDN U19242 ( .A(n18735), .B(n18734), .Z(n18739) );
  NANDN U19243 ( .A(n18737), .B(n18736), .Z(n18738) );
  NAND U19244 ( .A(n18739), .B(n18738), .Z(n18784) );
  XOR U19245 ( .A(n18783), .B(n18784), .Z(n18751) );
  OR U19246 ( .A(n18741), .B(n18740), .Z(n18745) );
  NANDN U19247 ( .A(n18743), .B(n18742), .Z(n18744) );
  NAND U19248 ( .A(n18745), .B(n18744), .Z(n18752) );
  XNOR U19249 ( .A(n18751), .B(n18752), .Z(n18753) );
  XNOR U19250 ( .A(n18754), .B(n18753), .Z(n18787) );
  XNOR U19251 ( .A(n18787), .B(sreg[1471]), .Z(n18789) );
  NAND U19252 ( .A(n18746), .B(sreg[1470]), .Z(n18750) );
  OR U19253 ( .A(n18748), .B(n18747), .Z(n18749) );
  AND U19254 ( .A(n18750), .B(n18749), .Z(n18788) );
  XOR U19255 ( .A(n18789), .B(n18788), .Z(c[1471]) );
  NANDN U19256 ( .A(n18752), .B(n18751), .Z(n18756) );
  NAND U19257 ( .A(n18754), .B(n18753), .Z(n18755) );
  NAND U19258 ( .A(n18756), .B(n18755), .Z(n18795) );
  NAND U19259 ( .A(b[0]), .B(a[456]), .Z(n18757) );
  XNOR U19260 ( .A(b[1]), .B(n18757), .Z(n18759) );
  NAND U19261 ( .A(n80), .B(a[455]), .Z(n18758) );
  AND U19262 ( .A(n18759), .B(n18758), .Z(n18812) );
  XOR U19263 ( .A(a[452]), .B(n42197), .Z(n18801) );
  NANDN U19264 ( .A(n18801), .B(n42173), .Z(n18762) );
  NANDN U19265 ( .A(n18760), .B(n42172), .Z(n18761) );
  NAND U19266 ( .A(n18762), .B(n18761), .Z(n18810) );
  NAND U19267 ( .A(b[7]), .B(a[448]), .Z(n18811) );
  XNOR U19268 ( .A(n18810), .B(n18811), .Z(n18813) );
  XOR U19269 ( .A(n18812), .B(n18813), .Z(n18819) );
  NANDN U19270 ( .A(n18763), .B(n42093), .Z(n18765) );
  XOR U19271 ( .A(n42134), .B(a[454]), .Z(n18804) );
  NANDN U19272 ( .A(n18804), .B(n42095), .Z(n18764) );
  NAND U19273 ( .A(n18765), .B(n18764), .Z(n18817) );
  NANDN U19274 ( .A(n18766), .B(n42231), .Z(n18768) );
  XOR U19275 ( .A(n199), .B(a[450]), .Z(n18807) );
  NANDN U19276 ( .A(n18807), .B(n42234), .Z(n18767) );
  AND U19277 ( .A(n18768), .B(n18767), .Z(n18816) );
  XNOR U19278 ( .A(n18817), .B(n18816), .Z(n18818) );
  XNOR U19279 ( .A(n18819), .B(n18818), .Z(n18823) );
  NANDN U19280 ( .A(n18770), .B(n18769), .Z(n18774) );
  NAND U19281 ( .A(n18772), .B(n18771), .Z(n18773) );
  AND U19282 ( .A(n18774), .B(n18773), .Z(n18822) );
  XOR U19283 ( .A(n18823), .B(n18822), .Z(n18824) );
  NANDN U19284 ( .A(n18776), .B(n18775), .Z(n18780) );
  NANDN U19285 ( .A(n18778), .B(n18777), .Z(n18779) );
  NAND U19286 ( .A(n18780), .B(n18779), .Z(n18825) );
  XOR U19287 ( .A(n18824), .B(n18825), .Z(n18792) );
  OR U19288 ( .A(n18782), .B(n18781), .Z(n18786) );
  NANDN U19289 ( .A(n18784), .B(n18783), .Z(n18785) );
  NAND U19290 ( .A(n18786), .B(n18785), .Z(n18793) );
  XNOR U19291 ( .A(n18792), .B(n18793), .Z(n18794) );
  XNOR U19292 ( .A(n18795), .B(n18794), .Z(n18828) );
  XNOR U19293 ( .A(n18828), .B(sreg[1472]), .Z(n18830) );
  NAND U19294 ( .A(n18787), .B(sreg[1471]), .Z(n18791) );
  OR U19295 ( .A(n18789), .B(n18788), .Z(n18790) );
  AND U19296 ( .A(n18791), .B(n18790), .Z(n18829) );
  XOR U19297 ( .A(n18830), .B(n18829), .Z(c[1472]) );
  NANDN U19298 ( .A(n18793), .B(n18792), .Z(n18797) );
  NAND U19299 ( .A(n18795), .B(n18794), .Z(n18796) );
  NAND U19300 ( .A(n18797), .B(n18796), .Z(n18836) );
  NAND U19301 ( .A(b[0]), .B(a[457]), .Z(n18798) );
  XNOR U19302 ( .A(b[1]), .B(n18798), .Z(n18800) );
  NAND U19303 ( .A(n80), .B(a[456]), .Z(n18799) );
  AND U19304 ( .A(n18800), .B(n18799), .Z(n18853) );
  XOR U19305 ( .A(a[453]), .B(n42197), .Z(n18842) );
  NANDN U19306 ( .A(n18842), .B(n42173), .Z(n18803) );
  NANDN U19307 ( .A(n18801), .B(n42172), .Z(n18802) );
  NAND U19308 ( .A(n18803), .B(n18802), .Z(n18851) );
  NAND U19309 ( .A(b[7]), .B(a[449]), .Z(n18852) );
  XNOR U19310 ( .A(n18851), .B(n18852), .Z(n18854) );
  XOR U19311 ( .A(n18853), .B(n18854), .Z(n18860) );
  NANDN U19312 ( .A(n18804), .B(n42093), .Z(n18806) );
  XOR U19313 ( .A(n42134), .B(a[455]), .Z(n18845) );
  NANDN U19314 ( .A(n18845), .B(n42095), .Z(n18805) );
  NAND U19315 ( .A(n18806), .B(n18805), .Z(n18858) );
  NANDN U19316 ( .A(n18807), .B(n42231), .Z(n18809) );
  XOR U19317 ( .A(n199), .B(a[451]), .Z(n18848) );
  NANDN U19318 ( .A(n18848), .B(n42234), .Z(n18808) );
  AND U19319 ( .A(n18809), .B(n18808), .Z(n18857) );
  XNOR U19320 ( .A(n18858), .B(n18857), .Z(n18859) );
  XNOR U19321 ( .A(n18860), .B(n18859), .Z(n18864) );
  NANDN U19322 ( .A(n18811), .B(n18810), .Z(n18815) );
  NAND U19323 ( .A(n18813), .B(n18812), .Z(n18814) );
  AND U19324 ( .A(n18815), .B(n18814), .Z(n18863) );
  XOR U19325 ( .A(n18864), .B(n18863), .Z(n18865) );
  NANDN U19326 ( .A(n18817), .B(n18816), .Z(n18821) );
  NANDN U19327 ( .A(n18819), .B(n18818), .Z(n18820) );
  NAND U19328 ( .A(n18821), .B(n18820), .Z(n18866) );
  XOR U19329 ( .A(n18865), .B(n18866), .Z(n18833) );
  OR U19330 ( .A(n18823), .B(n18822), .Z(n18827) );
  NANDN U19331 ( .A(n18825), .B(n18824), .Z(n18826) );
  NAND U19332 ( .A(n18827), .B(n18826), .Z(n18834) );
  XNOR U19333 ( .A(n18833), .B(n18834), .Z(n18835) );
  XNOR U19334 ( .A(n18836), .B(n18835), .Z(n18869) );
  XNOR U19335 ( .A(n18869), .B(sreg[1473]), .Z(n18871) );
  NAND U19336 ( .A(n18828), .B(sreg[1472]), .Z(n18832) );
  OR U19337 ( .A(n18830), .B(n18829), .Z(n18831) );
  AND U19338 ( .A(n18832), .B(n18831), .Z(n18870) );
  XOR U19339 ( .A(n18871), .B(n18870), .Z(c[1473]) );
  NANDN U19340 ( .A(n18834), .B(n18833), .Z(n18838) );
  NAND U19341 ( .A(n18836), .B(n18835), .Z(n18837) );
  NAND U19342 ( .A(n18838), .B(n18837), .Z(n18877) );
  NAND U19343 ( .A(b[0]), .B(a[458]), .Z(n18839) );
  XNOR U19344 ( .A(b[1]), .B(n18839), .Z(n18841) );
  NAND U19345 ( .A(n80), .B(a[457]), .Z(n18840) );
  AND U19346 ( .A(n18841), .B(n18840), .Z(n18894) );
  XOR U19347 ( .A(a[454]), .B(n42197), .Z(n18883) );
  NANDN U19348 ( .A(n18883), .B(n42173), .Z(n18844) );
  NANDN U19349 ( .A(n18842), .B(n42172), .Z(n18843) );
  NAND U19350 ( .A(n18844), .B(n18843), .Z(n18892) );
  NAND U19351 ( .A(b[7]), .B(a[450]), .Z(n18893) );
  XNOR U19352 ( .A(n18892), .B(n18893), .Z(n18895) );
  XOR U19353 ( .A(n18894), .B(n18895), .Z(n18901) );
  NANDN U19354 ( .A(n18845), .B(n42093), .Z(n18847) );
  XOR U19355 ( .A(n42134), .B(a[456]), .Z(n18886) );
  NANDN U19356 ( .A(n18886), .B(n42095), .Z(n18846) );
  NAND U19357 ( .A(n18847), .B(n18846), .Z(n18899) );
  NANDN U19358 ( .A(n18848), .B(n42231), .Z(n18850) );
  XOR U19359 ( .A(n199), .B(a[452]), .Z(n18889) );
  NANDN U19360 ( .A(n18889), .B(n42234), .Z(n18849) );
  AND U19361 ( .A(n18850), .B(n18849), .Z(n18898) );
  XNOR U19362 ( .A(n18899), .B(n18898), .Z(n18900) );
  XNOR U19363 ( .A(n18901), .B(n18900), .Z(n18905) );
  NANDN U19364 ( .A(n18852), .B(n18851), .Z(n18856) );
  NAND U19365 ( .A(n18854), .B(n18853), .Z(n18855) );
  AND U19366 ( .A(n18856), .B(n18855), .Z(n18904) );
  XOR U19367 ( .A(n18905), .B(n18904), .Z(n18906) );
  NANDN U19368 ( .A(n18858), .B(n18857), .Z(n18862) );
  NANDN U19369 ( .A(n18860), .B(n18859), .Z(n18861) );
  NAND U19370 ( .A(n18862), .B(n18861), .Z(n18907) );
  XOR U19371 ( .A(n18906), .B(n18907), .Z(n18874) );
  OR U19372 ( .A(n18864), .B(n18863), .Z(n18868) );
  NANDN U19373 ( .A(n18866), .B(n18865), .Z(n18867) );
  NAND U19374 ( .A(n18868), .B(n18867), .Z(n18875) );
  XNOR U19375 ( .A(n18874), .B(n18875), .Z(n18876) );
  XNOR U19376 ( .A(n18877), .B(n18876), .Z(n18910) );
  XNOR U19377 ( .A(n18910), .B(sreg[1474]), .Z(n18912) );
  NAND U19378 ( .A(n18869), .B(sreg[1473]), .Z(n18873) );
  OR U19379 ( .A(n18871), .B(n18870), .Z(n18872) );
  AND U19380 ( .A(n18873), .B(n18872), .Z(n18911) );
  XOR U19381 ( .A(n18912), .B(n18911), .Z(c[1474]) );
  NANDN U19382 ( .A(n18875), .B(n18874), .Z(n18879) );
  NAND U19383 ( .A(n18877), .B(n18876), .Z(n18878) );
  NAND U19384 ( .A(n18879), .B(n18878), .Z(n18918) );
  NAND U19385 ( .A(b[0]), .B(a[459]), .Z(n18880) );
  XNOR U19386 ( .A(b[1]), .B(n18880), .Z(n18882) );
  NAND U19387 ( .A(n80), .B(a[458]), .Z(n18881) );
  AND U19388 ( .A(n18882), .B(n18881), .Z(n18935) );
  XOR U19389 ( .A(a[455]), .B(n42197), .Z(n18924) );
  NANDN U19390 ( .A(n18924), .B(n42173), .Z(n18885) );
  NANDN U19391 ( .A(n18883), .B(n42172), .Z(n18884) );
  NAND U19392 ( .A(n18885), .B(n18884), .Z(n18933) );
  NAND U19393 ( .A(b[7]), .B(a[451]), .Z(n18934) );
  XNOR U19394 ( .A(n18933), .B(n18934), .Z(n18936) );
  XOR U19395 ( .A(n18935), .B(n18936), .Z(n18942) );
  NANDN U19396 ( .A(n18886), .B(n42093), .Z(n18888) );
  XOR U19397 ( .A(n42134), .B(a[457]), .Z(n18927) );
  NANDN U19398 ( .A(n18927), .B(n42095), .Z(n18887) );
  NAND U19399 ( .A(n18888), .B(n18887), .Z(n18940) );
  NANDN U19400 ( .A(n18889), .B(n42231), .Z(n18891) );
  XOR U19401 ( .A(n199), .B(a[453]), .Z(n18930) );
  NANDN U19402 ( .A(n18930), .B(n42234), .Z(n18890) );
  AND U19403 ( .A(n18891), .B(n18890), .Z(n18939) );
  XNOR U19404 ( .A(n18940), .B(n18939), .Z(n18941) );
  XNOR U19405 ( .A(n18942), .B(n18941), .Z(n18946) );
  NANDN U19406 ( .A(n18893), .B(n18892), .Z(n18897) );
  NAND U19407 ( .A(n18895), .B(n18894), .Z(n18896) );
  AND U19408 ( .A(n18897), .B(n18896), .Z(n18945) );
  XOR U19409 ( .A(n18946), .B(n18945), .Z(n18947) );
  NANDN U19410 ( .A(n18899), .B(n18898), .Z(n18903) );
  NANDN U19411 ( .A(n18901), .B(n18900), .Z(n18902) );
  NAND U19412 ( .A(n18903), .B(n18902), .Z(n18948) );
  XOR U19413 ( .A(n18947), .B(n18948), .Z(n18915) );
  OR U19414 ( .A(n18905), .B(n18904), .Z(n18909) );
  NANDN U19415 ( .A(n18907), .B(n18906), .Z(n18908) );
  NAND U19416 ( .A(n18909), .B(n18908), .Z(n18916) );
  XNOR U19417 ( .A(n18915), .B(n18916), .Z(n18917) );
  XNOR U19418 ( .A(n18918), .B(n18917), .Z(n18951) );
  XNOR U19419 ( .A(n18951), .B(sreg[1475]), .Z(n18953) );
  NAND U19420 ( .A(n18910), .B(sreg[1474]), .Z(n18914) );
  OR U19421 ( .A(n18912), .B(n18911), .Z(n18913) );
  AND U19422 ( .A(n18914), .B(n18913), .Z(n18952) );
  XOR U19423 ( .A(n18953), .B(n18952), .Z(c[1475]) );
  NANDN U19424 ( .A(n18916), .B(n18915), .Z(n18920) );
  NAND U19425 ( .A(n18918), .B(n18917), .Z(n18919) );
  NAND U19426 ( .A(n18920), .B(n18919), .Z(n18959) );
  NAND U19427 ( .A(b[0]), .B(a[460]), .Z(n18921) );
  XNOR U19428 ( .A(b[1]), .B(n18921), .Z(n18923) );
  NAND U19429 ( .A(n80), .B(a[459]), .Z(n18922) );
  AND U19430 ( .A(n18923), .B(n18922), .Z(n18976) );
  XOR U19431 ( .A(a[456]), .B(n42197), .Z(n18965) );
  NANDN U19432 ( .A(n18965), .B(n42173), .Z(n18926) );
  NANDN U19433 ( .A(n18924), .B(n42172), .Z(n18925) );
  NAND U19434 ( .A(n18926), .B(n18925), .Z(n18974) );
  NAND U19435 ( .A(b[7]), .B(a[452]), .Z(n18975) );
  XNOR U19436 ( .A(n18974), .B(n18975), .Z(n18977) );
  XOR U19437 ( .A(n18976), .B(n18977), .Z(n18983) );
  NANDN U19438 ( .A(n18927), .B(n42093), .Z(n18929) );
  XOR U19439 ( .A(n42134), .B(a[458]), .Z(n18968) );
  NANDN U19440 ( .A(n18968), .B(n42095), .Z(n18928) );
  NAND U19441 ( .A(n18929), .B(n18928), .Z(n18981) );
  NANDN U19442 ( .A(n18930), .B(n42231), .Z(n18932) );
  XOR U19443 ( .A(n199), .B(a[454]), .Z(n18971) );
  NANDN U19444 ( .A(n18971), .B(n42234), .Z(n18931) );
  AND U19445 ( .A(n18932), .B(n18931), .Z(n18980) );
  XNOR U19446 ( .A(n18981), .B(n18980), .Z(n18982) );
  XNOR U19447 ( .A(n18983), .B(n18982), .Z(n18987) );
  NANDN U19448 ( .A(n18934), .B(n18933), .Z(n18938) );
  NAND U19449 ( .A(n18936), .B(n18935), .Z(n18937) );
  AND U19450 ( .A(n18938), .B(n18937), .Z(n18986) );
  XOR U19451 ( .A(n18987), .B(n18986), .Z(n18988) );
  NANDN U19452 ( .A(n18940), .B(n18939), .Z(n18944) );
  NANDN U19453 ( .A(n18942), .B(n18941), .Z(n18943) );
  NAND U19454 ( .A(n18944), .B(n18943), .Z(n18989) );
  XOR U19455 ( .A(n18988), .B(n18989), .Z(n18956) );
  OR U19456 ( .A(n18946), .B(n18945), .Z(n18950) );
  NANDN U19457 ( .A(n18948), .B(n18947), .Z(n18949) );
  NAND U19458 ( .A(n18950), .B(n18949), .Z(n18957) );
  XNOR U19459 ( .A(n18956), .B(n18957), .Z(n18958) );
  XNOR U19460 ( .A(n18959), .B(n18958), .Z(n18992) );
  XNOR U19461 ( .A(n18992), .B(sreg[1476]), .Z(n18994) );
  NAND U19462 ( .A(n18951), .B(sreg[1475]), .Z(n18955) );
  OR U19463 ( .A(n18953), .B(n18952), .Z(n18954) );
  AND U19464 ( .A(n18955), .B(n18954), .Z(n18993) );
  XOR U19465 ( .A(n18994), .B(n18993), .Z(c[1476]) );
  NANDN U19466 ( .A(n18957), .B(n18956), .Z(n18961) );
  NAND U19467 ( .A(n18959), .B(n18958), .Z(n18960) );
  NAND U19468 ( .A(n18961), .B(n18960), .Z(n19000) );
  NAND U19469 ( .A(b[0]), .B(a[461]), .Z(n18962) );
  XNOR U19470 ( .A(b[1]), .B(n18962), .Z(n18964) );
  NAND U19471 ( .A(n80), .B(a[460]), .Z(n18963) );
  AND U19472 ( .A(n18964), .B(n18963), .Z(n19017) );
  XOR U19473 ( .A(a[457]), .B(n42197), .Z(n19006) );
  NANDN U19474 ( .A(n19006), .B(n42173), .Z(n18967) );
  NANDN U19475 ( .A(n18965), .B(n42172), .Z(n18966) );
  NAND U19476 ( .A(n18967), .B(n18966), .Z(n19015) );
  NAND U19477 ( .A(b[7]), .B(a[453]), .Z(n19016) );
  XNOR U19478 ( .A(n19015), .B(n19016), .Z(n19018) );
  XOR U19479 ( .A(n19017), .B(n19018), .Z(n19024) );
  NANDN U19480 ( .A(n18968), .B(n42093), .Z(n18970) );
  XOR U19481 ( .A(n42134), .B(a[459]), .Z(n19009) );
  NANDN U19482 ( .A(n19009), .B(n42095), .Z(n18969) );
  NAND U19483 ( .A(n18970), .B(n18969), .Z(n19022) );
  NANDN U19484 ( .A(n18971), .B(n42231), .Z(n18973) );
  XOR U19485 ( .A(n200), .B(a[455]), .Z(n19012) );
  NANDN U19486 ( .A(n19012), .B(n42234), .Z(n18972) );
  AND U19487 ( .A(n18973), .B(n18972), .Z(n19021) );
  XNOR U19488 ( .A(n19022), .B(n19021), .Z(n19023) );
  XNOR U19489 ( .A(n19024), .B(n19023), .Z(n19028) );
  NANDN U19490 ( .A(n18975), .B(n18974), .Z(n18979) );
  NAND U19491 ( .A(n18977), .B(n18976), .Z(n18978) );
  AND U19492 ( .A(n18979), .B(n18978), .Z(n19027) );
  XOR U19493 ( .A(n19028), .B(n19027), .Z(n19029) );
  NANDN U19494 ( .A(n18981), .B(n18980), .Z(n18985) );
  NANDN U19495 ( .A(n18983), .B(n18982), .Z(n18984) );
  NAND U19496 ( .A(n18985), .B(n18984), .Z(n19030) );
  XOR U19497 ( .A(n19029), .B(n19030), .Z(n18997) );
  OR U19498 ( .A(n18987), .B(n18986), .Z(n18991) );
  NANDN U19499 ( .A(n18989), .B(n18988), .Z(n18990) );
  NAND U19500 ( .A(n18991), .B(n18990), .Z(n18998) );
  XNOR U19501 ( .A(n18997), .B(n18998), .Z(n18999) );
  XNOR U19502 ( .A(n19000), .B(n18999), .Z(n19033) );
  XNOR U19503 ( .A(n19033), .B(sreg[1477]), .Z(n19035) );
  NAND U19504 ( .A(n18992), .B(sreg[1476]), .Z(n18996) );
  OR U19505 ( .A(n18994), .B(n18993), .Z(n18995) );
  AND U19506 ( .A(n18996), .B(n18995), .Z(n19034) );
  XOR U19507 ( .A(n19035), .B(n19034), .Z(c[1477]) );
  NANDN U19508 ( .A(n18998), .B(n18997), .Z(n19002) );
  NAND U19509 ( .A(n19000), .B(n18999), .Z(n19001) );
  NAND U19510 ( .A(n19002), .B(n19001), .Z(n19041) );
  NAND U19511 ( .A(b[0]), .B(a[462]), .Z(n19003) );
  XNOR U19512 ( .A(b[1]), .B(n19003), .Z(n19005) );
  NAND U19513 ( .A(n81), .B(a[461]), .Z(n19004) );
  AND U19514 ( .A(n19005), .B(n19004), .Z(n19058) );
  XOR U19515 ( .A(a[458]), .B(n42197), .Z(n19047) );
  NANDN U19516 ( .A(n19047), .B(n42173), .Z(n19008) );
  NANDN U19517 ( .A(n19006), .B(n42172), .Z(n19007) );
  NAND U19518 ( .A(n19008), .B(n19007), .Z(n19056) );
  NAND U19519 ( .A(b[7]), .B(a[454]), .Z(n19057) );
  XNOR U19520 ( .A(n19056), .B(n19057), .Z(n19059) );
  XOR U19521 ( .A(n19058), .B(n19059), .Z(n19065) );
  NANDN U19522 ( .A(n19009), .B(n42093), .Z(n19011) );
  XOR U19523 ( .A(n42134), .B(a[460]), .Z(n19050) );
  NANDN U19524 ( .A(n19050), .B(n42095), .Z(n19010) );
  NAND U19525 ( .A(n19011), .B(n19010), .Z(n19063) );
  NANDN U19526 ( .A(n19012), .B(n42231), .Z(n19014) );
  XOR U19527 ( .A(n200), .B(a[456]), .Z(n19053) );
  NANDN U19528 ( .A(n19053), .B(n42234), .Z(n19013) );
  AND U19529 ( .A(n19014), .B(n19013), .Z(n19062) );
  XNOR U19530 ( .A(n19063), .B(n19062), .Z(n19064) );
  XNOR U19531 ( .A(n19065), .B(n19064), .Z(n19069) );
  NANDN U19532 ( .A(n19016), .B(n19015), .Z(n19020) );
  NAND U19533 ( .A(n19018), .B(n19017), .Z(n19019) );
  AND U19534 ( .A(n19020), .B(n19019), .Z(n19068) );
  XOR U19535 ( .A(n19069), .B(n19068), .Z(n19070) );
  NANDN U19536 ( .A(n19022), .B(n19021), .Z(n19026) );
  NANDN U19537 ( .A(n19024), .B(n19023), .Z(n19025) );
  NAND U19538 ( .A(n19026), .B(n19025), .Z(n19071) );
  XOR U19539 ( .A(n19070), .B(n19071), .Z(n19038) );
  OR U19540 ( .A(n19028), .B(n19027), .Z(n19032) );
  NANDN U19541 ( .A(n19030), .B(n19029), .Z(n19031) );
  NAND U19542 ( .A(n19032), .B(n19031), .Z(n19039) );
  XNOR U19543 ( .A(n19038), .B(n19039), .Z(n19040) );
  XNOR U19544 ( .A(n19041), .B(n19040), .Z(n19074) );
  XNOR U19545 ( .A(n19074), .B(sreg[1478]), .Z(n19076) );
  NAND U19546 ( .A(n19033), .B(sreg[1477]), .Z(n19037) );
  OR U19547 ( .A(n19035), .B(n19034), .Z(n19036) );
  AND U19548 ( .A(n19037), .B(n19036), .Z(n19075) );
  XOR U19549 ( .A(n19076), .B(n19075), .Z(c[1478]) );
  NANDN U19550 ( .A(n19039), .B(n19038), .Z(n19043) );
  NAND U19551 ( .A(n19041), .B(n19040), .Z(n19042) );
  NAND U19552 ( .A(n19043), .B(n19042), .Z(n19082) );
  NAND U19553 ( .A(b[0]), .B(a[463]), .Z(n19044) );
  XNOR U19554 ( .A(b[1]), .B(n19044), .Z(n19046) );
  NAND U19555 ( .A(n81), .B(a[462]), .Z(n19045) );
  AND U19556 ( .A(n19046), .B(n19045), .Z(n19099) );
  XOR U19557 ( .A(a[459]), .B(n42197), .Z(n19088) );
  NANDN U19558 ( .A(n19088), .B(n42173), .Z(n19049) );
  NANDN U19559 ( .A(n19047), .B(n42172), .Z(n19048) );
  NAND U19560 ( .A(n19049), .B(n19048), .Z(n19097) );
  NAND U19561 ( .A(b[7]), .B(a[455]), .Z(n19098) );
  XNOR U19562 ( .A(n19097), .B(n19098), .Z(n19100) );
  XOR U19563 ( .A(n19099), .B(n19100), .Z(n19106) );
  NANDN U19564 ( .A(n19050), .B(n42093), .Z(n19052) );
  XOR U19565 ( .A(n42134), .B(a[461]), .Z(n19091) );
  NANDN U19566 ( .A(n19091), .B(n42095), .Z(n19051) );
  NAND U19567 ( .A(n19052), .B(n19051), .Z(n19104) );
  NANDN U19568 ( .A(n19053), .B(n42231), .Z(n19055) );
  XOR U19569 ( .A(n200), .B(a[457]), .Z(n19094) );
  NANDN U19570 ( .A(n19094), .B(n42234), .Z(n19054) );
  AND U19571 ( .A(n19055), .B(n19054), .Z(n19103) );
  XNOR U19572 ( .A(n19104), .B(n19103), .Z(n19105) );
  XNOR U19573 ( .A(n19106), .B(n19105), .Z(n19110) );
  NANDN U19574 ( .A(n19057), .B(n19056), .Z(n19061) );
  NAND U19575 ( .A(n19059), .B(n19058), .Z(n19060) );
  AND U19576 ( .A(n19061), .B(n19060), .Z(n19109) );
  XOR U19577 ( .A(n19110), .B(n19109), .Z(n19111) );
  NANDN U19578 ( .A(n19063), .B(n19062), .Z(n19067) );
  NANDN U19579 ( .A(n19065), .B(n19064), .Z(n19066) );
  NAND U19580 ( .A(n19067), .B(n19066), .Z(n19112) );
  XOR U19581 ( .A(n19111), .B(n19112), .Z(n19079) );
  OR U19582 ( .A(n19069), .B(n19068), .Z(n19073) );
  NANDN U19583 ( .A(n19071), .B(n19070), .Z(n19072) );
  NAND U19584 ( .A(n19073), .B(n19072), .Z(n19080) );
  XNOR U19585 ( .A(n19079), .B(n19080), .Z(n19081) );
  XNOR U19586 ( .A(n19082), .B(n19081), .Z(n19115) );
  XNOR U19587 ( .A(n19115), .B(sreg[1479]), .Z(n19117) );
  NAND U19588 ( .A(n19074), .B(sreg[1478]), .Z(n19078) );
  OR U19589 ( .A(n19076), .B(n19075), .Z(n19077) );
  AND U19590 ( .A(n19078), .B(n19077), .Z(n19116) );
  XOR U19591 ( .A(n19117), .B(n19116), .Z(c[1479]) );
  NANDN U19592 ( .A(n19080), .B(n19079), .Z(n19084) );
  NAND U19593 ( .A(n19082), .B(n19081), .Z(n19083) );
  NAND U19594 ( .A(n19084), .B(n19083), .Z(n19123) );
  NAND U19595 ( .A(b[0]), .B(a[464]), .Z(n19085) );
  XNOR U19596 ( .A(b[1]), .B(n19085), .Z(n19087) );
  NAND U19597 ( .A(n81), .B(a[463]), .Z(n19086) );
  AND U19598 ( .A(n19087), .B(n19086), .Z(n19140) );
  XOR U19599 ( .A(a[460]), .B(n42197), .Z(n19129) );
  NANDN U19600 ( .A(n19129), .B(n42173), .Z(n19090) );
  NANDN U19601 ( .A(n19088), .B(n42172), .Z(n19089) );
  NAND U19602 ( .A(n19090), .B(n19089), .Z(n19138) );
  NAND U19603 ( .A(b[7]), .B(a[456]), .Z(n19139) );
  XNOR U19604 ( .A(n19138), .B(n19139), .Z(n19141) );
  XOR U19605 ( .A(n19140), .B(n19141), .Z(n19147) );
  NANDN U19606 ( .A(n19091), .B(n42093), .Z(n19093) );
  XOR U19607 ( .A(n42134), .B(a[462]), .Z(n19132) );
  NANDN U19608 ( .A(n19132), .B(n42095), .Z(n19092) );
  NAND U19609 ( .A(n19093), .B(n19092), .Z(n19145) );
  NANDN U19610 ( .A(n19094), .B(n42231), .Z(n19096) );
  XOR U19611 ( .A(n200), .B(a[458]), .Z(n19135) );
  NANDN U19612 ( .A(n19135), .B(n42234), .Z(n19095) );
  AND U19613 ( .A(n19096), .B(n19095), .Z(n19144) );
  XNOR U19614 ( .A(n19145), .B(n19144), .Z(n19146) );
  XNOR U19615 ( .A(n19147), .B(n19146), .Z(n19151) );
  NANDN U19616 ( .A(n19098), .B(n19097), .Z(n19102) );
  NAND U19617 ( .A(n19100), .B(n19099), .Z(n19101) );
  AND U19618 ( .A(n19102), .B(n19101), .Z(n19150) );
  XOR U19619 ( .A(n19151), .B(n19150), .Z(n19152) );
  NANDN U19620 ( .A(n19104), .B(n19103), .Z(n19108) );
  NANDN U19621 ( .A(n19106), .B(n19105), .Z(n19107) );
  NAND U19622 ( .A(n19108), .B(n19107), .Z(n19153) );
  XOR U19623 ( .A(n19152), .B(n19153), .Z(n19120) );
  OR U19624 ( .A(n19110), .B(n19109), .Z(n19114) );
  NANDN U19625 ( .A(n19112), .B(n19111), .Z(n19113) );
  NAND U19626 ( .A(n19114), .B(n19113), .Z(n19121) );
  XNOR U19627 ( .A(n19120), .B(n19121), .Z(n19122) );
  XNOR U19628 ( .A(n19123), .B(n19122), .Z(n19156) );
  XNOR U19629 ( .A(n19156), .B(sreg[1480]), .Z(n19158) );
  NAND U19630 ( .A(n19115), .B(sreg[1479]), .Z(n19119) );
  OR U19631 ( .A(n19117), .B(n19116), .Z(n19118) );
  AND U19632 ( .A(n19119), .B(n19118), .Z(n19157) );
  XOR U19633 ( .A(n19158), .B(n19157), .Z(c[1480]) );
  NANDN U19634 ( .A(n19121), .B(n19120), .Z(n19125) );
  NAND U19635 ( .A(n19123), .B(n19122), .Z(n19124) );
  NAND U19636 ( .A(n19125), .B(n19124), .Z(n19164) );
  NAND U19637 ( .A(b[0]), .B(a[465]), .Z(n19126) );
  XNOR U19638 ( .A(b[1]), .B(n19126), .Z(n19128) );
  NAND U19639 ( .A(n81), .B(a[464]), .Z(n19127) );
  AND U19640 ( .A(n19128), .B(n19127), .Z(n19181) );
  XOR U19641 ( .A(a[461]), .B(n42197), .Z(n19170) );
  NANDN U19642 ( .A(n19170), .B(n42173), .Z(n19131) );
  NANDN U19643 ( .A(n19129), .B(n42172), .Z(n19130) );
  NAND U19644 ( .A(n19131), .B(n19130), .Z(n19179) );
  NAND U19645 ( .A(b[7]), .B(a[457]), .Z(n19180) );
  XNOR U19646 ( .A(n19179), .B(n19180), .Z(n19182) );
  XOR U19647 ( .A(n19181), .B(n19182), .Z(n19188) );
  NANDN U19648 ( .A(n19132), .B(n42093), .Z(n19134) );
  XOR U19649 ( .A(n42134), .B(a[463]), .Z(n19173) );
  NANDN U19650 ( .A(n19173), .B(n42095), .Z(n19133) );
  NAND U19651 ( .A(n19134), .B(n19133), .Z(n19186) );
  NANDN U19652 ( .A(n19135), .B(n42231), .Z(n19137) );
  XOR U19653 ( .A(n200), .B(a[459]), .Z(n19176) );
  NANDN U19654 ( .A(n19176), .B(n42234), .Z(n19136) );
  AND U19655 ( .A(n19137), .B(n19136), .Z(n19185) );
  XNOR U19656 ( .A(n19186), .B(n19185), .Z(n19187) );
  XNOR U19657 ( .A(n19188), .B(n19187), .Z(n19192) );
  NANDN U19658 ( .A(n19139), .B(n19138), .Z(n19143) );
  NAND U19659 ( .A(n19141), .B(n19140), .Z(n19142) );
  AND U19660 ( .A(n19143), .B(n19142), .Z(n19191) );
  XOR U19661 ( .A(n19192), .B(n19191), .Z(n19193) );
  NANDN U19662 ( .A(n19145), .B(n19144), .Z(n19149) );
  NANDN U19663 ( .A(n19147), .B(n19146), .Z(n19148) );
  NAND U19664 ( .A(n19149), .B(n19148), .Z(n19194) );
  XOR U19665 ( .A(n19193), .B(n19194), .Z(n19161) );
  OR U19666 ( .A(n19151), .B(n19150), .Z(n19155) );
  NANDN U19667 ( .A(n19153), .B(n19152), .Z(n19154) );
  NAND U19668 ( .A(n19155), .B(n19154), .Z(n19162) );
  XNOR U19669 ( .A(n19161), .B(n19162), .Z(n19163) );
  XNOR U19670 ( .A(n19164), .B(n19163), .Z(n19197) );
  XNOR U19671 ( .A(n19197), .B(sreg[1481]), .Z(n19199) );
  NAND U19672 ( .A(n19156), .B(sreg[1480]), .Z(n19160) );
  OR U19673 ( .A(n19158), .B(n19157), .Z(n19159) );
  AND U19674 ( .A(n19160), .B(n19159), .Z(n19198) );
  XOR U19675 ( .A(n19199), .B(n19198), .Z(c[1481]) );
  NANDN U19676 ( .A(n19162), .B(n19161), .Z(n19166) );
  NAND U19677 ( .A(n19164), .B(n19163), .Z(n19165) );
  NAND U19678 ( .A(n19166), .B(n19165), .Z(n19205) );
  NAND U19679 ( .A(b[0]), .B(a[466]), .Z(n19167) );
  XNOR U19680 ( .A(b[1]), .B(n19167), .Z(n19169) );
  NAND U19681 ( .A(n81), .B(a[465]), .Z(n19168) );
  AND U19682 ( .A(n19169), .B(n19168), .Z(n19222) );
  XOR U19683 ( .A(a[462]), .B(n42197), .Z(n19211) );
  NANDN U19684 ( .A(n19211), .B(n42173), .Z(n19172) );
  NANDN U19685 ( .A(n19170), .B(n42172), .Z(n19171) );
  NAND U19686 ( .A(n19172), .B(n19171), .Z(n19220) );
  NAND U19687 ( .A(b[7]), .B(a[458]), .Z(n19221) );
  XNOR U19688 ( .A(n19220), .B(n19221), .Z(n19223) );
  XOR U19689 ( .A(n19222), .B(n19223), .Z(n19229) );
  NANDN U19690 ( .A(n19173), .B(n42093), .Z(n19175) );
  XOR U19691 ( .A(n42134), .B(a[464]), .Z(n19214) );
  NANDN U19692 ( .A(n19214), .B(n42095), .Z(n19174) );
  NAND U19693 ( .A(n19175), .B(n19174), .Z(n19227) );
  NANDN U19694 ( .A(n19176), .B(n42231), .Z(n19178) );
  XOR U19695 ( .A(n200), .B(a[460]), .Z(n19217) );
  NANDN U19696 ( .A(n19217), .B(n42234), .Z(n19177) );
  AND U19697 ( .A(n19178), .B(n19177), .Z(n19226) );
  XNOR U19698 ( .A(n19227), .B(n19226), .Z(n19228) );
  XNOR U19699 ( .A(n19229), .B(n19228), .Z(n19233) );
  NANDN U19700 ( .A(n19180), .B(n19179), .Z(n19184) );
  NAND U19701 ( .A(n19182), .B(n19181), .Z(n19183) );
  AND U19702 ( .A(n19184), .B(n19183), .Z(n19232) );
  XOR U19703 ( .A(n19233), .B(n19232), .Z(n19234) );
  NANDN U19704 ( .A(n19186), .B(n19185), .Z(n19190) );
  NANDN U19705 ( .A(n19188), .B(n19187), .Z(n19189) );
  NAND U19706 ( .A(n19190), .B(n19189), .Z(n19235) );
  XOR U19707 ( .A(n19234), .B(n19235), .Z(n19202) );
  OR U19708 ( .A(n19192), .B(n19191), .Z(n19196) );
  NANDN U19709 ( .A(n19194), .B(n19193), .Z(n19195) );
  NAND U19710 ( .A(n19196), .B(n19195), .Z(n19203) );
  XNOR U19711 ( .A(n19202), .B(n19203), .Z(n19204) );
  XNOR U19712 ( .A(n19205), .B(n19204), .Z(n19238) );
  XNOR U19713 ( .A(n19238), .B(sreg[1482]), .Z(n19240) );
  NAND U19714 ( .A(n19197), .B(sreg[1481]), .Z(n19201) );
  OR U19715 ( .A(n19199), .B(n19198), .Z(n19200) );
  AND U19716 ( .A(n19201), .B(n19200), .Z(n19239) );
  XOR U19717 ( .A(n19240), .B(n19239), .Z(c[1482]) );
  NANDN U19718 ( .A(n19203), .B(n19202), .Z(n19207) );
  NAND U19719 ( .A(n19205), .B(n19204), .Z(n19206) );
  NAND U19720 ( .A(n19207), .B(n19206), .Z(n19246) );
  NAND U19721 ( .A(b[0]), .B(a[467]), .Z(n19208) );
  XNOR U19722 ( .A(b[1]), .B(n19208), .Z(n19210) );
  NAND U19723 ( .A(n81), .B(a[466]), .Z(n19209) );
  AND U19724 ( .A(n19210), .B(n19209), .Z(n19263) );
  XOR U19725 ( .A(a[463]), .B(n42197), .Z(n19252) );
  NANDN U19726 ( .A(n19252), .B(n42173), .Z(n19213) );
  NANDN U19727 ( .A(n19211), .B(n42172), .Z(n19212) );
  NAND U19728 ( .A(n19213), .B(n19212), .Z(n19261) );
  NAND U19729 ( .A(b[7]), .B(a[459]), .Z(n19262) );
  XNOR U19730 ( .A(n19261), .B(n19262), .Z(n19264) );
  XOR U19731 ( .A(n19263), .B(n19264), .Z(n19270) );
  NANDN U19732 ( .A(n19214), .B(n42093), .Z(n19216) );
  XOR U19733 ( .A(n42134), .B(a[465]), .Z(n19255) );
  NANDN U19734 ( .A(n19255), .B(n42095), .Z(n19215) );
  NAND U19735 ( .A(n19216), .B(n19215), .Z(n19268) );
  NANDN U19736 ( .A(n19217), .B(n42231), .Z(n19219) );
  XOR U19737 ( .A(n200), .B(a[461]), .Z(n19258) );
  NANDN U19738 ( .A(n19258), .B(n42234), .Z(n19218) );
  AND U19739 ( .A(n19219), .B(n19218), .Z(n19267) );
  XNOR U19740 ( .A(n19268), .B(n19267), .Z(n19269) );
  XNOR U19741 ( .A(n19270), .B(n19269), .Z(n19274) );
  NANDN U19742 ( .A(n19221), .B(n19220), .Z(n19225) );
  NAND U19743 ( .A(n19223), .B(n19222), .Z(n19224) );
  AND U19744 ( .A(n19225), .B(n19224), .Z(n19273) );
  XOR U19745 ( .A(n19274), .B(n19273), .Z(n19275) );
  NANDN U19746 ( .A(n19227), .B(n19226), .Z(n19231) );
  NANDN U19747 ( .A(n19229), .B(n19228), .Z(n19230) );
  NAND U19748 ( .A(n19231), .B(n19230), .Z(n19276) );
  XOR U19749 ( .A(n19275), .B(n19276), .Z(n19243) );
  OR U19750 ( .A(n19233), .B(n19232), .Z(n19237) );
  NANDN U19751 ( .A(n19235), .B(n19234), .Z(n19236) );
  NAND U19752 ( .A(n19237), .B(n19236), .Z(n19244) );
  XNOR U19753 ( .A(n19243), .B(n19244), .Z(n19245) );
  XNOR U19754 ( .A(n19246), .B(n19245), .Z(n19279) );
  XNOR U19755 ( .A(n19279), .B(sreg[1483]), .Z(n19281) );
  NAND U19756 ( .A(n19238), .B(sreg[1482]), .Z(n19242) );
  OR U19757 ( .A(n19240), .B(n19239), .Z(n19241) );
  AND U19758 ( .A(n19242), .B(n19241), .Z(n19280) );
  XOR U19759 ( .A(n19281), .B(n19280), .Z(c[1483]) );
  NANDN U19760 ( .A(n19244), .B(n19243), .Z(n19248) );
  NAND U19761 ( .A(n19246), .B(n19245), .Z(n19247) );
  NAND U19762 ( .A(n19248), .B(n19247), .Z(n19287) );
  NAND U19763 ( .A(b[0]), .B(a[468]), .Z(n19249) );
  XNOR U19764 ( .A(b[1]), .B(n19249), .Z(n19251) );
  NAND U19765 ( .A(n81), .B(a[467]), .Z(n19250) );
  AND U19766 ( .A(n19251), .B(n19250), .Z(n19304) );
  XOR U19767 ( .A(a[464]), .B(n42197), .Z(n19293) );
  NANDN U19768 ( .A(n19293), .B(n42173), .Z(n19254) );
  NANDN U19769 ( .A(n19252), .B(n42172), .Z(n19253) );
  NAND U19770 ( .A(n19254), .B(n19253), .Z(n19302) );
  NAND U19771 ( .A(b[7]), .B(a[460]), .Z(n19303) );
  XNOR U19772 ( .A(n19302), .B(n19303), .Z(n19305) );
  XOR U19773 ( .A(n19304), .B(n19305), .Z(n19311) );
  NANDN U19774 ( .A(n19255), .B(n42093), .Z(n19257) );
  XOR U19775 ( .A(n42134), .B(a[466]), .Z(n19296) );
  NANDN U19776 ( .A(n19296), .B(n42095), .Z(n19256) );
  NAND U19777 ( .A(n19257), .B(n19256), .Z(n19309) );
  NANDN U19778 ( .A(n19258), .B(n42231), .Z(n19260) );
  XOR U19779 ( .A(n200), .B(a[462]), .Z(n19299) );
  NANDN U19780 ( .A(n19299), .B(n42234), .Z(n19259) );
  AND U19781 ( .A(n19260), .B(n19259), .Z(n19308) );
  XNOR U19782 ( .A(n19309), .B(n19308), .Z(n19310) );
  XNOR U19783 ( .A(n19311), .B(n19310), .Z(n19315) );
  NANDN U19784 ( .A(n19262), .B(n19261), .Z(n19266) );
  NAND U19785 ( .A(n19264), .B(n19263), .Z(n19265) );
  AND U19786 ( .A(n19266), .B(n19265), .Z(n19314) );
  XOR U19787 ( .A(n19315), .B(n19314), .Z(n19316) );
  NANDN U19788 ( .A(n19268), .B(n19267), .Z(n19272) );
  NANDN U19789 ( .A(n19270), .B(n19269), .Z(n19271) );
  NAND U19790 ( .A(n19272), .B(n19271), .Z(n19317) );
  XOR U19791 ( .A(n19316), .B(n19317), .Z(n19284) );
  OR U19792 ( .A(n19274), .B(n19273), .Z(n19278) );
  NANDN U19793 ( .A(n19276), .B(n19275), .Z(n19277) );
  NAND U19794 ( .A(n19278), .B(n19277), .Z(n19285) );
  XNOR U19795 ( .A(n19284), .B(n19285), .Z(n19286) );
  XNOR U19796 ( .A(n19287), .B(n19286), .Z(n19320) );
  XNOR U19797 ( .A(n19320), .B(sreg[1484]), .Z(n19322) );
  NAND U19798 ( .A(n19279), .B(sreg[1483]), .Z(n19283) );
  OR U19799 ( .A(n19281), .B(n19280), .Z(n19282) );
  AND U19800 ( .A(n19283), .B(n19282), .Z(n19321) );
  XOR U19801 ( .A(n19322), .B(n19321), .Z(c[1484]) );
  NANDN U19802 ( .A(n19285), .B(n19284), .Z(n19289) );
  NAND U19803 ( .A(n19287), .B(n19286), .Z(n19288) );
  NAND U19804 ( .A(n19289), .B(n19288), .Z(n19328) );
  NAND U19805 ( .A(b[0]), .B(a[469]), .Z(n19290) );
  XNOR U19806 ( .A(b[1]), .B(n19290), .Z(n19292) );
  NAND U19807 ( .A(n82), .B(a[468]), .Z(n19291) );
  AND U19808 ( .A(n19292), .B(n19291), .Z(n19345) );
  XOR U19809 ( .A(a[465]), .B(n42197), .Z(n19334) );
  NANDN U19810 ( .A(n19334), .B(n42173), .Z(n19295) );
  NANDN U19811 ( .A(n19293), .B(n42172), .Z(n19294) );
  NAND U19812 ( .A(n19295), .B(n19294), .Z(n19343) );
  NAND U19813 ( .A(b[7]), .B(a[461]), .Z(n19344) );
  XNOR U19814 ( .A(n19343), .B(n19344), .Z(n19346) );
  XOR U19815 ( .A(n19345), .B(n19346), .Z(n19352) );
  NANDN U19816 ( .A(n19296), .B(n42093), .Z(n19298) );
  XOR U19817 ( .A(n42134), .B(a[467]), .Z(n19337) );
  NANDN U19818 ( .A(n19337), .B(n42095), .Z(n19297) );
  NAND U19819 ( .A(n19298), .B(n19297), .Z(n19350) );
  NANDN U19820 ( .A(n19299), .B(n42231), .Z(n19301) );
  XOR U19821 ( .A(n200), .B(a[463]), .Z(n19340) );
  NANDN U19822 ( .A(n19340), .B(n42234), .Z(n19300) );
  AND U19823 ( .A(n19301), .B(n19300), .Z(n19349) );
  XNOR U19824 ( .A(n19350), .B(n19349), .Z(n19351) );
  XNOR U19825 ( .A(n19352), .B(n19351), .Z(n19356) );
  NANDN U19826 ( .A(n19303), .B(n19302), .Z(n19307) );
  NAND U19827 ( .A(n19305), .B(n19304), .Z(n19306) );
  AND U19828 ( .A(n19307), .B(n19306), .Z(n19355) );
  XOR U19829 ( .A(n19356), .B(n19355), .Z(n19357) );
  NANDN U19830 ( .A(n19309), .B(n19308), .Z(n19313) );
  NANDN U19831 ( .A(n19311), .B(n19310), .Z(n19312) );
  NAND U19832 ( .A(n19313), .B(n19312), .Z(n19358) );
  XOR U19833 ( .A(n19357), .B(n19358), .Z(n19325) );
  OR U19834 ( .A(n19315), .B(n19314), .Z(n19319) );
  NANDN U19835 ( .A(n19317), .B(n19316), .Z(n19318) );
  NAND U19836 ( .A(n19319), .B(n19318), .Z(n19326) );
  XNOR U19837 ( .A(n19325), .B(n19326), .Z(n19327) );
  XNOR U19838 ( .A(n19328), .B(n19327), .Z(n19361) );
  XNOR U19839 ( .A(n19361), .B(sreg[1485]), .Z(n19363) );
  NAND U19840 ( .A(n19320), .B(sreg[1484]), .Z(n19324) );
  OR U19841 ( .A(n19322), .B(n19321), .Z(n19323) );
  AND U19842 ( .A(n19324), .B(n19323), .Z(n19362) );
  XOR U19843 ( .A(n19363), .B(n19362), .Z(c[1485]) );
  NANDN U19844 ( .A(n19326), .B(n19325), .Z(n19330) );
  NAND U19845 ( .A(n19328), .B(n19327), .Z(n19329) );
  NAND U19846 ( .A(n19330), .B(n19329), .Z(n19369) );
  NAND U19847 ( .A(b[0]), .B(a[470]), .Z(n19331) );
  XNOR U19848 ( .A(b[1]), .B(n19331), .Z(n19333) );
  NAND U19849 ( .A(n82), .B(a[469]), .Z(n19332) );
  AND U19850 ( .A(n19333), .B(n19332), .Z(n19386) );
  XOR U19851 ( .A(a[466]), .B(n42197), .Z(n19375) );
  NANDN U19852 ( .A(n19375), .B(n42173), .Z(n19336) );
  NANDN U19853 ( .A(n19334), .B(n42172), .Z(n19335) );
  NAND U19854 ( .A(n19336), .B(n19335), .Z(n19384) );
  NAND U19855 ( .A(b[7]), .B(a[462]), .Z(n19385) );
  XNOR U19856 ( .A(n19384), .B(n19385), .Z(n19387) );
  XOR U19857 ( .A(n19386), .B(n19387), .Z(n19393) );
  NANDN U19858 ( .A(n19337), .B(n42093), .Z(n19339) );
  XOR U19859 ( .A(n42134), .B(a[468]), .Z(n19378) );
  NANDN U19860 ( .A(n19378), .B(n42095), .Z(n19338) );
  NAND U19861 ( .A(n19339), .B(n19338), .Z(n19391) );
  NANDN U19862 ( .A(n19340), .B(n42231), .Z(n19342) );
  XOR U19863 ( .A(n200), .B(a[464]), .Z(n19381) );
  NANDN U19864 ( .A(n19381), .B(n42234), .Z(n19341) );
  AND U19865 ( .A(n19342), .B(n19341), .Z(n19390) );
  XNOR U19866 ( .A(n19391), .B(n19390), .Z(n19392) );
  XNOR U19867 ( .A(n19393), .B(n19392), .Z(n19397) );
  NANDN U19868 ( .A(n19344), .B(n19343), .Z(n19348) );
  NAND U19869 ( .A(n19346), .B(n19345), .Z(n19347) );
  AND U19870 ( .A(n19348), .B(n19347), .Z(n19396) );
  XOR U19871 ( .A(n19397), .B(n19396), .Z(n19398) );
  NANDN U19872 ( .A(n19350), .B(n19349), .Z(n19354) );
  NANDN U19873 ( .A(n19352), .B(n19351), .Z(n19353) );
  NAND U19874 ( .A(n19354), .B(n19353), .Z(n19399) );
  XOR U19875 ( .A(n19398), .B(n19399), .Z(n19366) );
  OR U19876 ( .A(n19356), .B(n19355), .Z(n19360) );
  NANDN U19877 ( .A(n19358), .B(n19357), .Z(n19359) );
  NAND U19878 ( .A(n19360), .B(n19359), .Z(n19367) );
  XNOR U19879 ( .A(n19366), .B(n19367), .Z(n19368) );
  XNOR U19880 ( .A(n19369), .B(n19368), .Z(n19402) );
  XNOR U19881 ( .A(n19402), .B(sreg[1486]), .Z(n19404) );
  NAND U19882 ( .A(n19361), .B(sreg[1485]), .Z(n19365) );
  OR U19883 ( .A(n19363), .B(n19362), .Z(n19364) );
  AND U19884 ( .A(n19365), .B(n19364), .Z(n19403) );
  XOR U19885 ( .A(n19404), .B(n19403), .Z(c[1486]) );
  NANDN U19886 ( .A(n19367), .B(n19366), .Z(n19371) );
  NAND U19887 ( .A(n19369), .B(n19368), .Z(n19370) );
  NAND U19888 ( .A(n19371), .B(n19370), .Z(n19410) );
  NAND U19889 ( .A(b[0]), .B(a[471]), .Z(n19372) );
  XNOR U19890 ( .A(b[1]), .B(n19372), .Z(n19374) );
  NAND U19891 ( .A(n82), .B(a[470]), .Z(n19373) );
  AND U19892 ( .A(n19374), .B(n19373), .Z(n19427) );
  XOR U19893 ( .A(a[467]), .B(n42197), .Z(n19416) );
  NANDN U19894 ( .A(n19416), .B(n42173), .Z(n19377) );
  NANDN U19895 ( .A(n19375), .B(n42172), .Z(n19376) );
  NAND U19896 ( .A(n19377), .B(n19376), .Z(n19425) );
  NAND U19897 ( .A(b[7]), .B(a[463]), .Z(n19426) );
  XNOR U19898 ( .A(n19425), .B(n19426), .Z(n19428) );
  XOR U19899 ( .A(n19427), .B(n19428), .Z(n19434) );
  NANDN U19900 ( .A(n19378), .B(n42093), .Z(n19380) );
  XOR U19901 ( .A(n42134), .B(a[469]), .Z(n19419) );
  NANDN U19902 ( .A(n19419), .B(n42095), .Z(n19379) );
  NAND U19903 ( .A(n19380), .B(n19379), .Z(n19432) );
  NANDN U19904 ( .A(n19381), .B(n42231), .Z(n19383) );
  XOR U19905 ( .A(n200), .B(a[465]), .Z(n19422) );
  NANDN U19906 ( .A(n19422), .B(n42234), .Z(n19382) );
  AND U19907 ( .A(n19383), .B(n19382), .Z(n19431) );
  XNOR U19908 ( .A(n19432), .B(n19431), .Z(n19433) );
  XNOR U19909 ( .A(n19434), .B(n19433), .Z(n19438) );
  NANDN U19910 ( .A(n19385), .B(n19384), .Z(n19389) );
  NAND U19911 ( .A(n19387), .B(n19386), .Z(n19388) );
  AND U19912 ( .A(n19389), .B(n19388), .Z(n19437) );
  XOR U19913 ( .A(n19438), .B(n19437), .Z(n19439) );
  NANDN U19914 ( .A(n19391), .B(n19390), .Z(n19395) );
  NANDN U19915 ( .A(n19393), .B(n19392), .Z(n19394) );
  NAND U19916 ( .A(n19395), .B(n19394), .Z(n19440) );
  XOR U19917 ( .A(n19439), .B(n19440), .Z(n19407) );
  OR U19918 ( .A(n19397), .B(n19396), .Z(n19401) );
  NANDN U19919 ( .A(n19399), .B(n19398), .Z(n19400) );
  NAND U19920 ( .A(n19401), .B(n19400), .Z(n19408) );
  XNOR U19921 ( .A(n19407), .B(n19408), .Z(n19409) );
  XNOR U19922 ( .A(n19410), .B(n19409), .Z(n19443) );
  XNOR U19923 ( .A(n19443), .B(sreg[1487]), .Z(n19445) );
  NAND U19924 ( .A(n19402), .B(sreg[1486]), .Z(n19406) );
  OR U19925 ( .A(n19404), .B(n19403), .Z(n19405) );
  AND U19926 ( .A(n19406), .B(n19405), .Z(n19444) );
  XOR U19927 ( .A(n19445), .B(n19444), .Z(c[1487]) );
  NANDN U19928 ( .A(n19408), .B(n19407), .Z(n19412) );
  NAND U19929 ( .A(n19410), .B(n19409), .Z(n19411) );
  NAND U19930 ( .A(n19412), .B(n19411), .Z(n19451) );
  NAND U19931 ( .A(b[0]), .B(a[472]), .Z(n19413) );
  XNOR U19932 ( .A(b[1]), .B(n19413), .Z(n19415) );
  NAND U19933 ( .A(n82), .B(a[471]), .Z(n19414) );
  AND U19934 ( .A(n19415), .B(n19414), .Z(n19468) );
  XOR U19935 ( .A(a[468]), .B(n42197), .Z(n19457) );
  NANDN U19936 ( .A(n19457), .B(n42173), .Z(n19418) );
  NANDN U19937 ( .A(n19416), .B(n42172), .Z(n19417) );
  NAND U19938 ( .A(n19418), .B(n19417), .Z(n19466) );
  NAND U19939 ( .A(b[7]), .B(a[464]), .Z(n19467) );
  XNOR U19940 ( .A(n19466), .B(n19467), .Z(n19469) );
  XOR U19941 ( .A(n19468), .B(n19469), .Z(n19475) );
  NANDN U19942 ( .A(n19419), .B(n42093), .Z(n19421) );
  XOR U19943 ( .A(n42134), .B(a[470]), .Z(n19460) );
  NANDN U19944 ( .A(n19460), .B(n42095), .Z(n19420) );
  NAND U19945 ( .A(n19421), .B(n19420), .Z(n19473) );
  NANDN U19946 ( .A(n19422), .B(n42231), .Z(n19424) );
  XOR U19947 ( .A(n200), .B(a[466]), .Z(n19463) );
  NANDN U19948 ( .A(n19463), .B(n42234), .Z(n19423) );
  AND U19949 ( .A(n19424), .B(n19423), .Z(n19472) );
  XNOR U19950 ( .A(n19473), .B(n19472), .Z(n19474) );
  XNOR U19951 ( .A(n19475), .B(n19474), .Z(n19479) );
  NANDN U19952 ( .A(n19426), .B(n19425), .Z(n19430) );
  NAND U19953 ( .A(n19428), .B(n19427), .Z(n19429) );
  AND U19954 ( .A(n19430), .B(n19429), .Z(n19478) );
  XOR U19955 ( .A(n19479), .B(n19478), .Z(n19480) );
  NANDN U19956 ( .A(n19432), .B(n19431), .Z(n19436) );
  NANDN U19957 ( .A(n19434), .B(n19433), .Z(n19435) );
  NAND U19958 ( .A(n19436), .B(n19435), .Z(n19481) );
  XOR U19959 ( .A(n19480), .B(n19481), .Z(n19448) );
  OR U19960 ( .A(n19438), .B(n19437), .Z(n19442) );
  NANDN U19961 ( .A(n19440), .B(n19439), .Z(n19441) );
  NAND U19962 ( .A(n19442), .B(n19441), .Z(n19449) );
  XNOR U19963 ( .A(n19448), .B(n19449), .Z(n19450) );
  XNOR U19964 ( .A(n19451), .B(n19450), .Z(n19484) );
  XNOR U19965 ( .A(n19484), .B(sreg[1488]), .Z(n19486) );
  NAND U19966 ( .A(n19443), .B(sreg[1487]), .Z(n19447) );
  OR U19967 ( .A(n19445), .B(n19444), .Z(n19446) );
  AND U19968 ( .A(n19447), .B(n19446), .Z(n19485) );
  XOR U19969 ( .A(n19486), .B(n19485), .Z(c[1488]) );
  NANDN U19970 ( .A(n19449), .B(n19448), .Z(n19453) );
  NAND U19971 ( .A(n19451), .B(n19450), .Z(n19452) );
  NAND U19972 ( .A(n19453), .B(n19452), .Z(n19492) );
  NAND U19973 ( .A(b[0]), .B(a[473]), .Z(n19454) );
  XNOR U19974 ( .A(b[1]), .B(n19454), .Z(n19456) );
  NAND U19975 ( .A(n82), .B(a[472]), .Z(n19455) );
  AND U19976 ( .A(n19456), .B(n19455), .Z(n19509) );
  XOR U19977 ( .A(a[469]), .B(n42197), .Z(n19498) );
  NANDN U19978 ( .A(n19498), .B(n42173), .Z(n19459) );
  NANDN U19979 ( .A(n19457), .B(n42172), .Z(n19458) );
  NAND U19980 ( .A(n19459), .B(n19458), .Z(n19507) );
  NAND U19981 ( .A(b[7]), .B(a[465]), .Z(n19508) );
  XNOR U19982 ( .A(n19507), .B(n19508), .Z(n19510) );
  XOR U19983 ( .A(n19509), .B(n19510), .Z(n19516) );
  NANDN U19984 ( .A(n19460), .B(n42093), .Z(n19462) );
  XOR U19985 ( .A(n42134), .B(a[471]), .Z(n19501) );
  NANDN U19986 ( .A(n19501), .B(n42095), .Z(n19461) );
  NAND U19987 ( .A(n19462), .B(n19461), .Z(n19514) );
  NANDN U19988 ( .A(n19463), .B(n42231), .Z(n19465) );
  XOR U19989 ( .A(n201), .B(a[467]), .Z(n19504) );
  NANDN U19990 ( .A(n19504), .B(n42234), .Z(n19464) );
  AND U19991 ( .A(n19465), .B(n19464), .Z(n19513) );
  XNOR U19992 ( .A(n19514), .B(n19513), .Z(n19515) );
  XNOR U19993 ( .A(n19516), .B(n19515), .Z(n19520) );
  NANDN U19994 ( .A(n19467), .B(n19466), .Z(n19471) );
  NAND U19995 ( .A(n19469), .B(n19468), .Z(n19470) );
  AND U19996 ( .A(n19471), .B(n19470), .Z(n19519) );
  XOR U19997 ( .A(n19520), .B(n19519), .Z(n19521) );
  NANDN U19998 ( .A(n19473), .B(n19472), .Z(n19477) );
  NANDN U19999 ( .A(n19475), .B(n19474), .Z(n19476) );
  NAND U20000 ( .A(n19477), .B(n19476), .Z(n19522) );
  XOR U20001 ( .A(n19521), .B(n19522), .Z(n19489) );
  OR U20002 ( .A(n19479), .B(n19478), .Z(n19483) );
  NANDN U20003 ( .A(n19481), .B(n19480), .Z(n19482) );
  NAND U20004 ( .A(n19483), .B(n19482), .Z(n19490) );
  XNOR U20005 ( .A(n19489), .B(n19490), .Z(n19491) );
  XNOR U20006 ( .A(n19492), .B(n19491), .Z(n19525) );
  XNOR U20007 ( .A(n19525), .B(sreg[1489]), .Z(n19527) );
  NAND U20008 ( .A(n19484), .B(sreg[1488]), .Z(n19488) );
  OR U20009 ( .A(n19486), .B(n19485), .Z(n19487) );
  AND U20010 ( .A(n19488), .B(n19487), .Z(n19526) );
  XOR U20011 ( .A(n19527), .B(n19526), .Z(c[1489]) );
  NANDN U20012 ( .A(n19490), .B(n19489), .Z(n19494) );
  NAND U20013 ( .A(n19492), .B(n19491), .Z(n19493) );
  NAND U20014 ( .A(n19494), .B(n19493), .Z(n19533) );
  NAND U20015 ( .A(b[0]), .B(a[474]), .Z(n19495) );
  XNOR U20016 ( .A(b[1]), .B(n19495), .Z(n19497) );
  NAND U20017 ( .A(n82), .B(a[473]), .Z(n19496) );
  AND U20018 ( .A(n19497), .B(n19496), .Z(n19550) );
  XOR U20019 ( .A(a[470]), .B(n42197), .Z(n19539) );
  NANDN U20020 ( .A(n19539), .B(n42173), .Z(n19500) );
  NANDN U20021 ( .A(n19498), .B(n42172), .Z(n19499) );
  NAND U20022 ( .A(n19500), .B(n19499), .Z(n19548) );
  NAND U20023 ( .A(b[7]), .B(a[466]), .Z(n19549) );
  XNOR U20024 ( .A(n19548), .B(n19549), .Z(n19551) );
  XOR U20025 ( .A(n19550), .B(n19551), .Z(n19557) );
  NANDN U20026 ( .A(n19501), .B(n42093), .Z(n19503) );
  XOR U20027 ( .A(n42134), .B(a[472]), .Z(n19542) );
  NANDN U20028 ( .A(n19542), .B(n42095), .Z(n19502) );
  NAND U20029 ( .A(n19503), .B(n19502), .Z(n19555) );
  NANDN U20030 ( .A(n19504), .B(n42231), .Z(n19506) );
  XOR U20031 ( .A(n201), .B(a[468]), .Z(n19545) );
  NANDN U20032 ( .A(n19545), .B(n42234), .Z(n19505) );
  AND U20033 ( .A(n19506), .B(n19505), .Z(n19554) );
  XNOR U20034 ( .A(n19555), .B(n19554), .Z(n19556) );
  XNOR U20035 ( .A(n19557), .B(n19556), .Z(n19561) );
  NANDN U20036 ( .A(n19508), .B(n19507), .Z(n19512) );
  NAND U20037 ( .A(n19510), .B(n19509), .Z(n19511) );
  AND U20038 ( .A(n19512), .B(n19511), .Z(n19560) );
  XOR U20039 ( .A(n19561), .B(n19560), .Z(n19562) );
  NANDN U20040 ( .A(n19514), .B(n19513), .Z(n19518) );
  NANDN U20041 ( .A(n19516), .B(n19515), .Z(n19517) );
  NAND U20042 ( .A(n19518), .B(n19517), .Z(n19563) );
  XOR U20043 ( .A(n19562), .B(n19563), .Z(n19530) );
  OR U20044 ( .A(n19520), .B(n19519), .Z(n19524) );
  NANDN U20045 ( .A(n19522), .B(n19521), .Z(n19523) );
  NAND U20046 ( .A(n19524), .B(n19523), .Z(n19531) );
  XNOR U20047 ( .A(n19530), .B(n19531), .Z(n19532) );
  XNOR U20048 ( .A(n19533), .B(n19532), .Z(n19566) );
  XNOR U20049 ( .A(n19566), .B(sreg[1490]), .Z(n19568) );
  NAND U20050 ( .A(n19525), .B(sreg[1489]), .Z(n19529) );
  OR U20051 ( .A(n19527), .B(n19526), .Z(n19528) );
  AND U20052 ( .A(n19529), .B(n19528), .Z(n19567) );
  XOR U20053 ( .A(n19568), .B(n19567), .Z(c[1490]) );
  NANDN U20054 ( .A(n19531), .B(n19530), .Z(n19535) );
  NAND U20055 ( .A(n19533), .B(n19532), .Z(n19534) );
  NAND U20056 ( .A(n19535), .B(n19534), .Z(n19574) );
  NAND U20057 ( .A(b[0]), .B(a[475]), .Z(n19536) );
  XNOR U20058 ( .A(b[1]), .B(n19536), .Z(n19538) );
  NAND U20059 ( .A(n82), .B(a[474]), .Z(n19537) );
  AND U20060 ( .A(n19538), .B(n19537), .Z(n19591) );
  XOR U20061 ( .A(a[471]), .B(n42197), .Z(n19580) );
  NANDN U20062 ( .A(n19580), .B(n42173), .Z(n19541) );
  NANDN U20063 ( .A(n19539), .B(n42172), .Z(n19540) );
  NAND U20064 ( .A(n19541), .B(n19540), .Z(n19589) );
  NAND U20065 ( .A(b[7]), .B(a[467]), .Z(n19590) );
  XNOR U20066 ( .A(n19589), .B(n19590), .Z(n19592) );
  XOR U20067 ( .A(n19591), .B(n19592), .Z(n19598) );
  NANDN U20068 ( .A(n19542), .B(n42093), .Z(n19544) );
  XOR U20069 ( .A(n42134), .B(a[473]), .Z(n19583) );
  NANDN U20070 ( .A(n19583), .B(n42095), .Z(n19543) );
  NAND U20071 ( .A(n19544), .B(n19543), .Z(n19596) );
  NANDN U20072 ( .A(n19545), .B(n42231), .Z(n19547) );
  XOR U20073 ( .A(n201), .B(a[469]), .Z(n19586) );
  NANDN U20074 ( .A(n19586), .B(n42234), .Z(n19546) );
  AND U20075 ( .A(n19547), .B(n19546), .Z(n19595) );
  XNOR U20076 ( .A(n19596), .B(n19595), .Z(n19597) );
  XNOR U20077 ( .A(n19598), .B(n19597), .Z(n19602) );
  NANDN U20078 ( .A(n19549), .B(n19548), .Z(n19553) );
  NAND U20079 ( .A(n19551), .B(n19550), .Z(n19552) );
  AND U20080 ( .A(n19553), .B(n19552), .Z(n19601) );
  XOR U20081 ( .A(n19602), .B(n19601), .Z(n19603) );
  NANDN U20082 ( .A(n19555), .B(n19554), .Z(n19559) );
  NANDN U20083 ( .A(n19557), .B(n19556), .Z(n19558) );
  NAND U20084 ( .A(n19559), .B(n19558), .Z(n19604) );
  XOR U20085 ( .A(n19603), .B(n19604), .Z(n19571) );
  OR U20086 ( .A(n19561), .B(n19560), .Z(n19565) );
  NANDN U20087 ( .A(n19563), .B(n19562), .Z(n19564) );
  NAND U20088 ( .A(n19565), .B(n19564), .Z(n19572) );
  XNOR U20089 ( .A(n19571), .B(n19572), .Z(n19573) );
  XNOR U20090 ( .A(n19574), .B(n19573), .Z(n19607) );
  XNOR U20091 ( .A(n19607), .B(sreg[1491]), .Z(n19609) );
  NAND U20092 ( .A(n19566), .B(sreg[1490]), .Z(n19570) );
  OR U20093 ( .A(n19568), .B(n19567), .Z(n19569) );
  AND U20094 ( .A(n19570), .B(n19569), .Z(n19608) );
  XOR U20095 ( .A(n19609), .B(n19608), .Z(c[1491]) );
  NANDN U20096 ( .A(n19572), .B(n19571), .Z(n19576) );
  NAND U20097 ( .A(n19574), .B(n19573), .Z(n19575) );
  NAND U20098 ( .A(n19576), .B(n19575), .Z(n19615) );
  NAND U20099 ( .A(b[0]), .B(a[476]), .Z(n19577) );
  XNOR U20100 ( .A(b[1]), .B(n19577), .Z(n19579) );
  NAND U20101 ( .A(n83), .B(a[475]), .Z(n19578) );
  AND U20102 ( .A(n19579), .B(n19578), .Z(n19632) );
  XOR U20103 ( .A(a[472]), .B(n42197), .Z(n19621) );
  NANDN U20104 ( .A(n19621), .B(n42173), .Z(n19582) );
  NANDN U20105 ( .A(n19580), .B(n42172), .Z(n19581) );
  NAND U20106 ( .A(n19582), .B(n19581), .Z(n19630) );
  NAND U20107 ( .A(b[7]), .B(a[468]), .Z(n19631) );
  XNOR U20108 ( .A(n19630), .B(n19631), .Z(n19633) );
  XOR U20109 ( .A(n19632), .B(n19633), .Z(n19639) );
  NANDN U20110 ( .A(n19583), .B(n42093), .Z(n19585) );
  XOR U20111 ( .A(n42134), .B(a[474]), .Z(n19624) );
  NANDN U20112 ( .A(n19624), .B(n42095), .Z(n19584) );
  NAND U20113 ( .A(n19585), .B(n19584), .Z(n19637) );
  NANDN U20114 ( .A(n19586), .B(n42231), .Z(n19588) );
  XOR U20115 ( .A(n201), .B(a[470]), .Z(n19627) );
  NANDN U20116 ( .A(n19627), .B(n42234), .Z(n19587) );
  AND U20117 ( .A(n19588), .B(n19587), .Z(n19636) );
  XNOR U20118 ( .A(n19637), .B(n19636), .Z(n19638) );
  XNOR U20119 ( .A(n19639), .B(n19638), .Z(n19643) );
  NANDN U20120 ( .A(n19590), .B(n19589), .Z(n19594) );
  NAND U20121 ( .A(n19592), .B(n19591), .Z(n19593) );
  AND U20122 ( .A(n19594), .B(n19593), .Z(n19642) );
  XOR U20123 ( .A(n19643), .B(n19642), .Z(n19644) );
  NANDN U20124 ( .A(n19596), .B(n19595), .Z(n19600) );
  NANDN U20125 ( .A(n19598), .B(n19597), .Z(n19599) );
  NAND U20126 ( .A(n19600), .B(n19599), .Z(n19645) );
  XOR U20127 ( .A(n19644), .B(n19645), .Z(n19612) );
  OR U20128 ( .A(n19602), .B(n19601), .Z(n19606) );
  NANDN U20129 ( .A(n19604), .B(n19603), .Z(n19605) );
  NAND U20130 ( .A(n19606), .B(n19605), .Z(n19613) );
  XNOR U20131 ( .A(n19612), .B(n19613), .Z(n19614) );
  XNOR U20132 ( .A(n19615), .B(n19614), .Z(n19648) );
  XNOR U20133 ( .A(n19648), .B(sreg[1492]), .Z(n19650) );
  NAND U20134 ( .A(n19607), .B(sreg[1491]), .Z(n19611) );
  OR U20135 ( .A(n19609), .B(n19608), .Z(n19610) );
  AND U20136 ( .A(n19611), .B(n19610), .Z(n19649) );
  XOR U20137 ( .A(n19650), .B(n19649), .Z(c[1492]) );
  NANDN U20138 ( .A(n19613), .B(n19612), .Z(n19617) );
  NAND U20139 ( .A(n19615), .B(n19614), .Z(n19616) );
  NAND U20140 ( .A(n19617), .B(n19616), .Z(n19656) );
  NAND U20141 ( .A(b[0]), .B(a[477]), .Z(n19618) );
  XNOR U20142 ( .A(b[1]), .B(n19618), .Z(n19620) );
  NAND U20143 ( .A(n83), .B(a[476]), .Z(n19619) );
  AND U20144 ( .A(n19620), .B(n19619), .Z(n19673) );
  XOR U20145 ( .A(a[473]), .B(n42197), .Z(n19662) );
  NANDN U20146 ( .A(n19662), .B(n42173), .Z(n19623) );
  NANDN U20147 ( .A(n19621), .B(n42172), .Z(n19622) );
  NAND U20148 ( .A(n19623), .B(n19622), .Z(n19671) );
  NAND U20149 ( .A(b[7]), .B(a[469]), .Z(n19672) );
  XNOR U20150 ( .A(n19671), .B(n19672), .Z(n19674) );
  XOR U20151 ( .A(n19673), .B(n19674), .Z(n19680) );
  NANDN U20152 ( .A(n19624), .B(n42093), .Z(n19626) );
  XOR U20153 ( .A(n42134), .B(a[475]), .Z(n19665) );
  NANDN U20154 ( .A(n19665), .B(n42095), .Z(n19625) );
  NAND U20155 ( .A(n19626), .B(n19625), .Z(n19678) );
  NANDN U20156 ( .A(n19627), .B(n42231), .Z(n19629) );
  XOR U20157 ( .A(n201), .B(a[471]), .Z(n19668) );
  NANDN U20158 ( .A(n19668), .B(n42234), .Z(n19628) );
  AND U20159 ( .A(n19629), .B(n19628), .Z(n19677) );
  XNOR U20160 ( .A(n19678), .B(n19677), .Z(n19679) );
  XNOR U20161 ( .A(n19680), .B(n19679), .Z(n19684) );
  NANDN U20162 ( .A(n19631), .B(n19630), .Z(n19635) );
  NAND U20163 ( .A(n19633), .B(n19632), .Z(n19634) );
  AND U20164 ( .A(n19635), .B(n19634), .Z(n19683) );
  XOR U20165 ( .A(n19684), .B(n19683), .Z(n19685) );
  NANDN U20166 ( .A(n19637), .B(n19636), .Z(n19641) );
  NANDN U20167 ( .A(n19639), .B(n19638), .Z(n19640) );
  NAND U20168 ( .A(n19641), .B(n19640), .Z(n19686) );
  XOR U20169 ( .A(n19685), .B(n19686), .Z(n19653) );
  OR U20170 ( .A(n19643), .B(n19642), .Z(n19647) );
  NANDN U20171 ( .A(n19645), .B(n19644), .Z(n19646) );
  NAND U20172 ( .A(n19647), .B(n19646), .Z(n19654) );
  XNOR U20173 ( .A(n19653), .B(n19654), .Z(n19655) );
  XNOR U20174 ( .A(n19656), .B(n19655), .Z(n19689) );
  XNOR U20175 ( .A(n19689), .B(sreg[1493]), .Z(n19691) );
  NAND U20176 ( .A(n19648), .B(sreg[1492]), .Z(n19652) );
  OR U20177 ( .A(n19650), .B(n19649), .Z(n19651) );
  AND U20178 ( .A(n19652), .B(n19651), .Z(n19690) );
  XOR U20179 ( .A(n19691), .B(n19690), .Z(c[1493]) );
  NANDN U20180 ( .A(n19654), .B(n19653), .Z(n19658) );
  NAND U20181 ( .A(n19656), .B(n19655), .Z(n19657) );
  NAND U20182 ( .A(n19658), .B(n19657), .Z(n19697) );
  NAND U20183 ( .A(b[0]), .B(a[478]), .Z(n19659) );
  XNOR U20184 ( .A(b[1]), .B(n19659), .Z(n19661) );
  NAND U20185 ( .A(n83), .B(a[477]), .Z(n19660) );
  AND U20186 ( .A(n19661), .B(n19660), .Z(n19714) );
  XOR U20187 ( .A(a[474]), .B(n42197), .Z(n19703) );
  NANDN U20188 ( .A(n19703), .B(n42173), .Z(n19664) );
  NANDN U20189 ( .A(n19662), .B(n42172), .Z(n19663) );
  NAND U20190 ( .A(n19664), .B(n19663), .Z(n19712) );
  NAND U20191 ( .A(b[7]), .B(a[470]), .Z(n19713) );
  XNOR U20192 ( .A(n19712), .B(n19713), .Z(n19715) );
  XOR U20193 ( .A(n19714), .B(n19715), .Z(n19721) );
  NANDN U20194 ( .A(n19665), .B(n42093), .Z(n19667) );
  XOR U20195 ( .A(n42134), .B(a[476]), .Z(n19706) );
  NANDN U20196 ( .A(n19706), .B(n42095), .Z(n19666) );
  NAND U20197 ( .A(n19667), .B(n19666), .Z(n19719) );
  NANDN U20198 ( .A(n19668), .B(n42231), .Z(n19670) );
  XOR U20199 ( .A(n201), .B(a[472]), .Z(n19709) );
  NANDN U20200 ( .A(n19709), .B(n42234), .Z(n19669) );
  AND U20201 ( .A(n19670), .B(n19669), .Z(n19718) );
  XNOR U20202 ( .A(n19719), .B(n19718), .Z(n19720) );
  XNOR U20203 ( .A(n19721), .B(n19720), .Z(n19725) );
  NANDN U20204 ( .A(n19672), .B(n19671), .Z(n19676) );
  NAND U20205 ( .A(n19674), .B(n19673), .Z(n19675) );
  AND U20206 ( .A(n19676), .B(n19675), .Z(n19724) );
  XOR U20207 ( .A(n19725), .B(n19724), .Z(n19726) );
  NANDN U20208 ( .A(n19678), .B(n19677), .Z(n19682) );
  NANDN U20209 ( .A(n19680), .B(n19679), .Z(n19681) );
  NAND U20210 ( .A(n19682), .B(n19681), .Z(n19727) );
  XOR U20211 ( .A(n19726), .B(n19727), .Z(n19694) );
  OR U20212 ( .A(n19684), .B(n19683), .Z(n19688) );
  NANDN U20213 ( .A(n19686), .B(n19685), .Z(n19687) );
  NAND U20214 ( .A(n19688), .B(n19687), .Z(n19695) );
  XNOR U20215 ( .A(n19694), .B(n19695), .Z(n19696) );
  XNOR U20216 ( .A(n19697), .B(n19696), .Z(n19730) );
  XNOR U20217 ( .A(n19730), .B(sreg[1494]), .Z(n19732) );
  NAND U20218 ( .A(n19689), .B(sreg[1493]), .Z(n19693) );
  OR U20219 ( .A(n19691), .B(n19690), .Z(n19692) );
  AND U20220 ( .A(n19693), .B(n19692), .Z(n19731) );
  XOR U20221 ( .A(n19732), .B(n19731), .Z(c[1494]) );
  NANDN U20222 ( .A(n19695), .B(n19694), .Z(n19699) );
  NAND U20223 ( .A(n19697), .B(n19696), .Z(n19698) );
  NAND U20224 ( .A(n19699), .B(n19698), .Z(n19738) );
  NAND U20225 ( .A(b[0]), .B(a[479]), .Z(n19700) );
  XNOR U20226 ( .A(b[1]), .B(n19700), .Z(n19702) );
  NAND U20227 ( .A(n83), .B(a[478]), .Z(n19701) );
  AND U20228 ( .A(n19702), .B(n19701), .Z(n19755) );
  XOR U20229 ( .A(a[475]), .B(n42197), .Z(n19744) );
  NANDN U20230 ( .A(n19744), .B(n42173), .Z(n19705) );
  NANDN U20231 ( .A(n19703), .B(n42172), .Z(n19704) );
  NAND U20232 ( .A(n19705), .B(n19704), .Z(n19753) );
  NAND U20233 ( .A(b[7]), .B(a[471]), .Z(n19754) );
  XNOR U20234 ( .A(n19753), .B(n19754), .Z(n19756) );
  XOR U20235 ( .A(n19755), .B(n19756), .Z(n19762) );
  NANDN U20236 ( .A(n19706), .B(n42093), .Z(n19708) );
  XOR U20237 ( .A(n42134), .B(a[477]), .Z(n19747) );
  NANDN U20238 ( .A(n19747), .B(n42095), .Z(n19707) );
  NAND U20239 ( .A(n19708), .B(n19707), .Z(n19760) );
  NANDN U20240 ( .A(n19709), .B(n42231), .Z(n19711) );
  XOR U20241 ( .A(n201), .B(a[473]), .Z(n19750) );
  NANDN U20242 ( .A(n19750), .B(n42234), .Z(n19710) );
  AND U20243 ( .A(n19711), .B(n19710), .Z(n19759) );
  XNOR U20244 ( .A(n19760), .B(n19759), .Z(n19761) );
  XNOR U20245 ( .A(n19762), .B(n19761), .Z(n19766) );
  NANDN U20246 ( .A(n19713), .B(n19712), .Z(n19717) );
  NAND U20247 ( .A(n19715), .B(n19714), .Z(n19716) );
  AND U20248 ( .A(n19717), .B(n19716), .Z(n19765) );
  XOR U20249 ( .A(n19766), .B(n19765), .Z(n19767) );
  NANDN U20250 ( .A(n19719), .B(n19718), .Z(n19723) );
  NANDN U20251 ( .A(n19721), .B(n19720), .Z(n19722) );
  NAND U20252 ( .A(n19723), .B(n19722), .Z(n19768) );
  XOR U20253 ( .A(n19767), .B(n19768), .Z(n19735) );
  OR U20254 ( .A(n19725), .B(n19724), .Z(n19729) );
  NANDN U20255 ( .A(n19727), .B(n19726), .Z(n19728) );
  NAND U20256 ( .A(n19729), .B(n19728), .Z(n19736) );
  XNOR U20257 ( .A(n19735), .B(n19736), .Z(n19737) );
  XNOR U20258 ( .A(n19738), .B(n19737), .Z(n19771) );
  XNOR U20259 ( .A(n19771), .B(sreg[1495]), .Z(n19773) );
  NAND U20260 ( .A(n19730), .B(sreg[1494]), .Z(n19734) );
  OR U20261 ( .A(n19732), .B(n19731), .Z(n19733) );
  AND U20262 ( .A(n19734), .B(n19733), .Z(n19772) );
  XOR U20263 ( .A(n19773), .B(n19772), .Z(c[1495]) );
  NANDN U20264 ( .A(n19736), .B(n19735), .Z(n19740) );
  NAND U20265 ( .A(n19738), .B(n19737), .Z(n19739) );
  NAND U20266 ( .A(n19740), .B(n19739), .Z(n19779) );
  NAND U20267 ( .A(b[0]), .B(a[480]), .Z(n19741) );
  XNOR U20268 ( .A(b[1]), .B(n19741), .Z(n19743) );
  NAND U20269 ( .A(n83), .B(a[479]), .Z(n19742) );
  AND U20270 ( .A(n19743), .B(n19742), .Z(n19796) );
  XOR U20271 ( .A(a[476]), .B(n42197), .Z(n19785) );
  NANDN U20272 ( .A(n19785), .B(n42173), .Z(n19746) );
  NANDN U20273 ( .A(n19744), .B(n42172), .Z(n19745) );
  NAND U20274 ( .A(n19746), .B(n19745), .Z(n19794) );
  NAND U20275 ( .A(b[7]), .B(a[472]), .Z(n19795) );
  XNOR U20276 ( .A(n19794), .B(n19795), .Z(n19797) );
  XOR U20277 ( .A(n19796), .B(n19797), .Z(n19803) );
  NANDN U20278 ( .A(n19747), .B(n42093), .Z(n19749) );
  XOR U20279 ( .A(n42134), .B(a[478]), .Z(n19788) );
  NANDN U20280 ( .A(n19788), .B(n42095), .Z(n19748) );
  NAND U20281 ( .A(n19749), .B(n19748), .Z(n19801) );
  NANDN U20282 ( .A(n19750), .B(n42231), .Z(n19752) );
  XOR U20283 ( .A(n201), .B(a[474]), .Z(n19791) );
  NANDN U20284 ( .A(n19791), .B(n42234), .Z(n19751) );
  AND U20285 ( .A(n19752), .B(n19751), .Z(n19800) );
  XNOR U20286 ( .A(n19801), .B(n19800), .Z(n19802) );
  XNOR U20287 ( .A(n19803), .B(n19802), .Z(n19807) );
  NANDN U20288 ( .A(n19754), .B(n19753), .Z(n19758) );
  NAND U20289 ( .A(n19756), .B(n19755), .Z(n19757) );
  AND U20290 ( .A(n19758), .B(n19757), .Z(n19806) );
  XOR U20291 ( .A(n19807), .B(n19806), .Z(n19808) );
  NANDN U20292 ( .A(n19760), .B(n19759), .Z(n19764) );
  NANDN U20293 ( .A(n19762), .B(n19761), .Z(n19763) );
  NAND U20294 ( .A(n19764), .B(n19763), .Z(n19809) );
  XOR U20295 ( .A(n19808), .B(n19809), .Z(n19776) );
  OR U20296 ( .A(n19766), .B(n19765), .Z(n19770) );
  NANDN U20297 ( .A(n19768), .B(n19767), .Z(n19769) );
  NAND U20298 ( .A(n19770), .B(n19769), .Z(n19777) );
  XNOR U20299 ( .A(n19776), .B(n19777), .Z(n19778) );
  XNOR U20300 ( .A(n19779), .B(n19778), .Z(n19812) );
  XNOR U20301 ( .A(n19812), .B(sreg[1496]), .Z(n19814) );
  NAND U20302 ( .A(n19771), .B(sreg[1495]), .Z(n19775) );
  OR U20303 ( .A(n19773), .B(n19772), .Z(n19774) );
  AND U20304 ( .A(n19775), .B(n19774), .Z(n19813) );
  XOR U20305 ( .A(n19814), .B(n19813), .Z(c[1496]) );
  NANDN U20306 ( .A(n19777), .B(n19776), .Z(n19781) );
  NAND U20307 ( .A(n19779), .B(n19778), .Z(n19780) );
  NAND U20308 ( .A(n19781), .B(n19780), .Z(n19820) );
  NAND U20309 ( .A(b[0]), .B(a[481]), .Z(n19782) );
  XNOR U20310 ( .A(b[1]), .B(n19782), .Z(n19784) );
  NAND U20311 ( .A(n83), .B(a[480]), .Z(n19783) );
  AND U20312 ( .A(n19784), .B(n19783), .Z(n19837) );
  XOR U20313 ( .A(a[477]), .B(n42197), .Z(n19826) );
  NANDN U20314 ( .A(n19826), .B(n42173), .Z(n19787) );
  NANDN U20315 ( .A(n19785), .B(n42172), .Z(n19786) );
  NAND U20316 ( .A(n19787), .B(n19786), .Z(n19835) );
  NAND U20317 ( .A(b[7]), .B(a[473]), .Z(n19836) );
  XNOR U20318 ( .A(n19835), .B(n19836), .Z(n19838) );
  XOR U20319 ( .A(n19837), .B(n19838), .Z(n19844) );
  NANDN U20320 ( .A(n19788), .B(n42093), .Z(n19790) );
  XOR U20321 ( .A(n42134), .B(a[479]), .Z(n19829) );
  NANDN U20322 ( .A(n19829), .B(n42095), .Z(n19789) );
  NAND U20323 ( .A(n19790), .B(n19789), .Z(n19842) );
  NANDN U20324 ( .A(n19791), .B(n42231), .Z(n19793) );
  XOR U20325 ( .A(n201), .B(a[475]), .Z(n19832) );
  NANDN U20326 ( .A(n19832), .B(n42234), .Z(n19792) );
  AND U20327 ( .A(n19793), .B(n19792), .Z(n19841) );
  XNOR U20328 ( .A(n19842), .B(n19841), .Z(n19843) );
  XNOR U20329 ( .A(n19844), .B(n19843), .Z(n19848) );
  NANDN U20330 ( .A(n19795), .B(n19794), .Z(n19799) );
  NAND U20331 ( .A(n19797), .B(n19796), .Z(n19798) );
  AND U20332 ( .A(n19799), .B(n19798), .Z(n19847) );
  XOR U20333 ( .A(n19848), .B(n19847), .Z(n19849) );
  NANDN U20334 ( .A(n19801), .B(n19800), .Z(n19805) );
  NANDN U20335 ( .A(n19803), .B(n19802), .Z(n19804) );
  NAND U20336 ( .A(n19805), .B(n19804), .Z(n19850) );
  XOR U20337 ( .A(n19849), .B(n19850), .Z(n19817) );
  OR U20338 ( .A(n19807), .B(n19806), .Z(n19811) );
  NANDN U20339 ( .A(n19809), .B(n19808), .Z(n19810) );
  NAND U20340 ( .A(n19811), .B(n19810), .Z(n19818) );
  XNOR U20341 ( .A(n19817), .B(n19818), .Z(n19819) );
  XNOR U20342 ( .A(n19820), .B(n19819), .Z(n19853) );
  XNOR U20343 ( .A(n19853), .B(sreg[1497]), .Z(n19855) );
  NAND U20344 ( .A(n19812), .B(sreg[1496]), .Z(n19816) );
  OR U20345 ( .A(n19814), .B(n19813), .Z(n19815) );
  AND U20346 ( .A(n19816), .B(n19815), .Z(n19854) );
  XOR U20347 ( .A(n19855), .B(n19854), .Z(c[1497]) );
  NANDN U20348 ( .A(n19818), .B(n19817), .Z(n19822) );
  NAND U20349 ( .A(n19820), .B(n19819), .Z(n19821) );
  NAND U20350 ( .A(n19822), .B(n19821), .Z(n19861) );
  NAND U20351 ( .A(b[0]), .B(a[482]), .Z(n19823) );
  XNOR U20352 ( .A(b[1]), .B(n19823), .Z(n19825) );
  NAND U20353 ( .A(n83), .B(a[481]), .Z(n19824) );
  AND U20354 ( .A(n19825), .B(n19824), .Z(n19878) );
  XOR U20355 ( .A(a[478]), .B(n42197), .Z(n19867) );
  NANDN U20356 ( .A(n19867), .B(n42173), .Z(n19828) );
  NANDN U20357 ( .A(n19826), .B(n42172), .Z(n19827) );
  NAND U20358 ( .A(n19828), .B(n19827), .Z(n19876) );
  NAND U20359 ( .A(b[7]), .B(a[474]), .Z(n19877) );
  XNOR U20360 ( .A(n19876), .B(n19877), .Z(n19879) );
  XOR U20361 ( .A(n19878), .B(n19879), .Z(n19885) );
  NANDN U20362 ( .A(n19829), .B(n42093), .Z(n19831) );
  XOR U20363 ( .A(n42134), .B(a[480]), .Z(n19870) );
  NANDN U20364 ( .A(n19870), .B(n42095), .Z(n19830) );
  NAND U20365 ( .A(n19831), .B(n19830), .Z(n19883) );
  NANDN U20366 ( .A(n19832), .B(n42231), .Z(n19834) );
  XOR U20367 ( .A(n201), .B(a[476]), .Z(n19873) );
  NANDN U20368 ( .A(n19873), .B(n42234), .Z(n19833) );
  AND U20369 ( .A(n19834), .B(n19833), .Z(n19882) );
  XNOR U20370 ( .A(n19883), .B(n19882), .Z(n19884) );
  XNOR U20371 ( .A(n19885), .B(n19884), .Z(n19889) );
  NANDN U20372 ( .A(n19836), .B(n19835), .Z(n19840) );
  NAND U20373 ( .A(n19838), .B(n19837), .Z(n19839) );
  AND U20374 ( .A(n19840), .B(n19839), .Z(n19888) );
  XOR U20375 ( .A(n19889), .B(n19888), .Z(n19890) );
  NANDN U20376 ( .A(n19842), .B(n19841), .Z(n19846) );
  NANDN U20377 ( .A(n19844), .B(n19843), .Z(n19845) );
  NAND U20378 ( .A(n19846), .B(n19845), .Z(n19891) );
  XOR U20379 ( .A(n19890), .B(n19891), .Z(n19858) );
  OR U20380 ( .A(n19848), .B(n19847), .Z(n19852) );
  NANDN U20381 ( .A(n19850), .B(n19849), .Z(n19851) );
  NAND U20382 ( .A(n19852), .B(n19851), .Z(n19859) );
  XNOR U20383 ( .A(n19858), .B(n19859), .Z(n19860) );
  XNOR U20384 ( .A(n19861), .B(n19860), .Z(n19894) );
  XNOR U20385 ( .A(n19894), .B(sreg[1498]), .Z(n19896) );
  NAND U20386 ( .A(n19853), .B(sreg[1497]), .Z(n19857) );
  OR U20387 ( .A(n19855), .B(n19854), .Z(n19856) );
  AND U20388 ( .A(n19857), .B(n19856), .Z(n19895) );
  XOR U20389 ( .A(n19896), .B(n19895), .Z(c[1498]) );
  NANDN U20390 ( .A(n19859), .B(n19858), .Z(n19863) );
  NAND U20391 ( .A(n19861), .B(n19860), .Z(n19862) );
  NAND U20392 ( .A(n19863), .B(n19862), .Z(n19902) );
  NAND U20393 ( .A(b[0]), .B(a[483]), .Z(n19864) );
  XNOR U20394 ( .A(b[1]), .B(n19864), .Z(n19866) );
  NAND U20395 ( .A(n84), .B(a[482]), .Z(n19865) );
  AND U20396 ( .A(n19866), .B(n19865), .Z(n19919) );
  XOR U20397 ( .A(a[479]), .B(n42197), .Z(n19908) );
  NANDN U20398 ( .A(n19908), .B(n42173), .Z(n19869) );
  NANDN U20399 ( .A(n19867), .B(n42172), .Z(n19868) );
  NAND U20400 ( .A(n19869), .B(n19868), .Z(n19917) );
  NAND U20401 ( .A(b[7]), .B(a[475]), .Z(n19918) );
  XNOR U20402 ( .A(n19917), .B(n19918), .Z(n19920) );
  XOR U20403 ( .A(n19919), .B(n19920), .Z(n19926) );
  NANDN U20404 ( .A(n19870), .B(n42093), .Z(n19872) );
  XOR U20405 ( .A(n42134), .B(a[481]), .Z(n19911) );
  NANDN U20406 ( .A(n19911), .B(n42095), .Z(n19871) );
  NAND U20407 ( .A(n19872), .B(n19871), .Z(n19924) );
  NANDN U20408 ( .A(n19873), .B(n42231), .Z(n19875) );
  XOR U20409 ( .A(n201), .B(a[477]), .Z(n19914) );
  NANDN U20410 ( .A(n19914), .B(n42234), .Z(n19874) );
  AND U20411 ( .A(n19875), .B(n19874), .Z(n19923) );
  XNOR U20412 ( .A(n19924), .B(n19923), .Z(n19925) );
  XNOR U20413 ( .A(n19926), .B(n19925), .Z(n19930) );
  NANDN U20414 ( .A(n19877), .B(n19876), .Z(n19881) );
  NAND U20415 ( .A(n19879), .B(n19878), .Z(n19880) );
  AND U20416 ( .A(n19881), .B(n19880), .Z(n19929) );
  XOR U20417 ( .A(n19930), .B(n19929), .Z(n19931) );
  NANDN U20418 ( .A(n19883), .B(n19882), .Z(n19887) );
  NANDN U20419 ( .A(n19885), .B(n19884), .Z(n19886) );
  NAND U20420 ( .A(n19887), .B(n19886), .Z(n19932) );
  XOR U20421 ( .A(n19931), .B(n19932), .Z(n19899) );
  OR U20422 ( .A(n19889), .B(n19888), .Z(n19893) );
  NANDN U20423 ( .A(n19891), .B(n19890), .Z(n19892) );
  NAND U20424 ( .A(n19893), .B(n19892), .Z(n19900) );
  XNOR U20425 ( .A(n19899), .B(n19900), .Z(n19901) );
  XNOR U20426 ( .A(n19902), .B(n19901), .Z(n19935) );
  XNOR U20427 ( .A(n19935), .B(sreg[1499]), .Z(n19937) );
  NAND U20428 ( .A(n19894), .B(sreg[1498]), .Z(n19898) );
  OR U20429 ( .A(n19896), .B(n19895), .Z(n19897) );
  AND U20430 ( .A(n19898), .B(n19897), .Z(n19936) );
  XOR U20431 ( .A(n19937), .B(n19936), .Z(c[1499]) );
  NANDN U20432 ( .A(n19900), .B(n19899), .Z(n19904) );
  NAND U20433 ( .A(n19902), .B(n19901), .Z(n19903) );
  NAND U20434 ( .A(n19904), .B(n19903), .Z(n19943) );
  NAND U20435 ( .A(b[0]), .B(a[484]), .Z(n19905) );
  XNOR U20436 ( .A(b[1]), .B(n19905), .Z(n19907) );
  NAND U20437 ( .A(n84), .B(a[483]), .Z(n19906) );
  AND U20438 ( .A(n19907), .B(n19906), .Z(n19960) );
  XOR U20439 ( .A(a[480]), .B(n42197), .Z(n19949) );
  NANDN U20440 ( .A(n19949), .B(n42173), .Z(n19910) );
  NANDN U20441 ( .A(n19908), .B(n42172), .Z(n19909) );
  NAND U20442 ( .A(n19910), .B(n19909), .Z(n19958) );
  NAND U20443 ( .A(b[7]), .B(a[476]), .Z(n19959) );
  XNOR U20444 ( .A(n19958), .B(n19959), .Z(n19961) );
  XOR U20445 ( .A(n19960), .B(n19961), .Z(n19967) );
  NANDN U20446 ( .A(n19911), .B(n42093), .Z(n19913) );
  XOR U20447 ( .A(n42134), .B(a[482]), .Z(n19952) );
  NANDN U20448 ( .A(n19952), .B(n42095), .Z(n19912) );
  NAND U20449 ( .A(n19913), .B(n19912), .Z(n19965) );
  NANDN U20450 ( .A(n19914), .B(n42231), .Z(n19916) );
  XOR U20451 ( .A(n201), .B(a[478]), .Z(n19955) );
  NANDN U20452 ( .A(n19955), .B(n42234), .Z(n19915) );
  AND U20453 ( .A(n19916), .B(n19915), .Z(n19964) );
  XNOR U20454 ( .A(n19965), .B(n19964), .Z(n19966) );
  XNOR U20455 ( .A(n19967), .B(n19966), .Z(n19971) );
  NANDN U20456 ( .A(n19918), .B(n19917), .Z(n19922) );
  NAND U20457 ( .A(n19920), .B(n19919), .Z(n19921) );
  AND U20458 ( .A(n19922), .B(n19921), .Z(n19970) );
  XOR U20459 ( .A(n19971), .B(n19970), .Z(n19972) );
  NANDN U20460 ( .A(n19924), .B(n19923), .Z(n19928) );
  NANDN U20461 ( .A(n19926), .B(n19925), .Z(n19927) );
  NAND U20462 ( .A(n19928), .B(n19927), .Z(n19973) );
  XOR U20463 ( .A(n19972), .B(n19973), .Z(n19940) );
  OR U20464 ( .A(n19930), .B(n19929), .Z(n19934) );
  NANDN U20465 ( .A(n19932), .B(n19931), .Z(n19933) );
  NAND U20466 ( .A(n19934), .B(n19933), .Z(n19941) );
  XNOR U20467 ( .A(n19940), .B(n19941), .Z(n19942) );
  XNOR U20468 ( .A(n19943), .B(n19942), .Z(n19976) );
  XNOR U20469 ( .A(n19976), .B(sreg[1500]), .Z(n19978) );
  NAND U20470 ( .A(n19935), .B(sreg[1499]), .Z(n19939) );
  OR U20471 ( .A(n19937), .B(n19936), .Z(n19938) );
  AND U20472 ( .A(n19939), .B(n19938), .Z(n19977) );
  XOR U20473 ( .A(n19978), .B(n19977), .Z(c[1500]) );
  NANDN U20474 ( .A(n19941), .B(n19940), .Z(n19945) );
  NAND U20475 ( .A(n19943), .B(n19942), .Z(n19944) );
  NAND U20476 ( .A(n19945), .B(n19944), .Z(n19984) );
  NAND U20477 ( .A(b[0]), .B(a[485]), .Z(n19946) );
  XNOR U20478 ( .A(b[1]), .B(n19946), .Z(n19948) );
  NAND U20479 ( .A(n84), .B(a[484]), .Z(n19947) );
  AND U20480 ( .A(n19948), .B(n19947), .Z(n20001) );
  XOR U20481 ( .A(a[481]), .B(n42197), .Z(n19990) );
  NANDN U20482 ( .A(n19990), .B(n42173), .Z(n19951) );
  NANDN U20483 ( .A(n19949), .B(n42172), .Z(n19950) );
  NAND U20484 ( .A(n19951), .B(n19950), .Z(n19999) );
  NAND U20485 ( .A(b[7]), .B(a[477]), .Z(n20000) );
  XNOR U20486 ( .A(n19999), .B(n20000), .Z(n20002) );
  XOR U20487 ( .A(n20001), .B(n20002), .Z(n20008) );
  NANDN U20488 ( .A(n19952), .B(n42093), .Z(n19954) );
  XOR U20489 ( .A(n42134), .B(a[483]), .Z(n19993) );
  NANDN U20490 ( .A(n19993), .B(n42095), .Z(n19953) );
  NAND U20491 ( .A(n19954), .B(n19953), .Z(n20006) );
  NANDN U20492 ( .A(n19955), .B(n42231), .Z(n19957) );
  XOR U20493 ( .A(n202), .B(a[479]), .Z(n19996) );
  NANDN U20494 ( .A(n19996), .B(n42234), .Z(n19956) );
  AND U20495 ( .A(n19957), .B(n19956), .Z(n20005) );
  XNOR U20496 ( .A(n20006), .B(n20005), .Z(n20007) );
  XNOR U20497 ( .A(n20008), .B(n20007), .Z(n20012) );
  NANDN U20498 ( .A(n19959), .B(n19958), .Z(n19963) );
  NAND U20499 ( .A(n19961), .B(n19960), .Z(n19962) );
  AND U20500 ( .A(n19963), .B(n19962), .Z(n20011) );
  XOR U20501 ( .A(n20012), .B(n20011), .Z(n20013) );
  NANDN U20502 ( .A(n19965), .B(n19964), .Z(n19969) );
  NANDN U20503 ( .A(n19967), .B(n19966), .Z(n19968) );
  NAND U20504 ( .A(n19969), .B(n19968), .Z(n20014) );
  XOR U20505 ( .A(n20013), .B(n20014), .Z(n19981) );
  OR U20506 ( .A(n19971), .B(n19970), .Z(n19975) );
  NANDN U20507 ( .A(n19973), .B(n19972), .Z(n19974) );
  NAND U20508 ( .A(n19975), .B(n19974), .Z(n19982) );
  XNOR U20509 ( .A(n19981), .B(n19982), .Z(n19983) );
  XNOR U20510 ( .A(n19984), .B(n19983), .Z(n20017) );
  XNOR U20511 ( .A(n20017), .B(sreg[1501]), .Z(n20019) );
  NAND U20512 ( .A(n19976), .B(sreg[1500]), .Z(n19980) );
  OR U20513 ( .A(n19978), .B(n19977), .Z(n19979) );
  AND U20514 ( .A(n19980), .B(n19979), .Z(n20018) );
  XOR U20515 ( .A(n20019), .B(n20018), .Z(c[1501]) );
  NANDN U20516 ( .A(n19982), .B(n19981), .Z(n19986) );
  NAND U20517 ( .A(n19984), .B(n19983), .Z(n19985) );
  NAND U20518 ( .A(n19986), .B(n19985), .Z(n20025) );
  NAND U20519 ( .A(b[0]), .B(a[486]), .Z(n19987) );
  XNOR U20520 ( .A(b[1]), .B(n19987), .Z(n19989) );
  NAND U20521 ( .A(n84), .B(a[485]), .Z(n19988) );
  AND U20522 ( .A(n19989), .B(n19988), .Z(n20042) );
  XOR U20523 ( .A(a[482]), .B(n42197), .Z(n20031) );
  NANDN U20524 ( .A(n20031), .B(n42173), .Z(n19992) );
  NANDN U20525 ( .A(n19990), .B(n42172), .Z(n19991) );
  NAND U20526 ( .A(n19992), .B(n19991), .Z(n20040) );
  NAND U20527 ( .A(b[7]), .B(a[478]), .Z(n20041) );
  XNOR U20528 ( .A(n20040), .B(n20041), .Z(n20043) );
  XOR U20529 ( .A(n20042), .B(n20043), .Z(n20049) );
  NANDN U20530 ( .A(n19993), .B(n42093), .Z(n19995) );
  XOR U20531 ( .A(n42134), .B(a[484]), .Z(n20034) );
  NANDN U20532 ( .A(n20034), .B(n42095), .Z(n19994) );
  NAND U20533 ( .A(n19995), .B(n19994), .Z(n20047) );
  NANDN U20534 ( .A(n19996), .B(n42231), .Z(n19998) );
  XOR U20535 ( .A(n202), .B(a[480]), .Z(n20037) );
  NANDN U20536 ( .A(n20037), .B(n42234), .Z(n19997) );
  AND U20537 ( .A(n19998), .B(n19997), .Z(n20046) );
  XNOR U20538 ( .A(n20047), .B(n20046), .Z(n20048) );
  XNOR U20539 ( .A(n20049), .B(n20048), .Z(n20053) );
  NANDN U20540 ( .A(n20000), .B(n19999), .Z(n20004) );
  NAND U20541 ( .A(n20002), .B(n20001), .Z(n20003) );
  AND U20542 ( .A(n20004), .B(n20003), .Z(n20052) );
  XOR U20543 ( .A(n20053), .B(n20052), .Z(n20054) );
  NANDN U20544 ( .A(n20006), .B(n20005), .Z(n20010) );
  NANDN U20545 ( .A(n20008), .B(n20007), .Z(n20009) );
  NAND U20546 ( .A(n20010), .B(n20009), .Z(n20055) );
  XOR U20547 ( .A(n20054), .B(n20055), .Z(n20022) );
  OR U20548 ( .A(n20012), .B(n20011), .Z(n20016) );
  NANDN U20549 ( .A(n20014), .B(n20013), .Z(n20015) );
  NAND U20550 ( .A(n20016), .B(n20015), .Z(n20023) );
  XNOR U20551 ( .A(n20022), .B(n20023), .Z(n20024) );
  XNOR U20552 ( .A(n20025), .B(n20024), .Z(n20058) );
  XNOR U20553 ( .A(n20058), .B(sreg[1502]), .Z(n20060) );
  NAND U20554 ( .A(n20017), .B(sreg[1501]), .Z(n20021) );
  OR U20555 ( .A(n20019), .B(n20018), .Z(n20020) );
  AND U20556 ( .A(n20021), .B(n20020), .Z(n20059) );
  XOR U20557 ( .A(n20060), .B(n20059), .Z(c[1502]) );
  NANDN U20558 ( .A(n20023), .B(n20022), .Z(n20027) );
  NAND U20559 ( .A(n20025), .B(n20024), .Z(n20026) );
  NAND U20560 ( .A(n20027), .B(n20026), .Z(n20066) );
  NAND U20561 ( .A(b[0]), .B(a[487]), .Z(n20028) );
  XNOR U20562 ( .A(b[1]), .B(n20028), .Z(n20030) );
  NAND U20563 ( .A(n84), .B(a[486]), .Z(n20029) );
  AND U20564 ( .A(n20030), .B(n20029), .Z(n20083) );
  XOR U20565 ( .A(a[483]), .B(n42197), .Z(n20072) );
  NANDN U20566 ( .A(n20072), .B(n42173), .Z(n20033) );
  NANDN U20567 ( .A(n20031), .B(n42172), .Z(n20032) );
  NAND U20568 ( .A(n20033), .B(n20032), .Z(n20081) );
  NAND U20569 ( .A(b[7]), .B(a[479]), .Z(n20082) );
  XNOR U20570 ( .A(n20081), .B(n20082), .Z(n20084) );
  XOR U20571 ( .A(n20083), .B(n20084), .Z(n20090) );
  NANDN U20572 ( .A(n20034), .B(n42093), .Z(n20036) );
  XOR U20573 ( .A(n42134), .B(a[485]), .Z(n20075) );
  NANDN U20574 ( .A(n20075), .B(n42095), .Z(n20035) );
  NAND U20575 ( .A(n20036), .B(n20035), .Z(n20088) );
  NANDN U20576 ( .A(n20037), .B(n42231), .Z(n20039) );
  XOR U20577 ( .A(n202), .B(a[481]), .Z(n20078) );
  NANDN U20578 ( .A(n20078), .B(n42234), .Z(n20038) );
  AND U20579 ( .A(n20039), .B(n20038), .Z(n20087) );
  XNOR U20580 ( .A(n20088), .B(n20087), .Z(n20089) );
  XNOR U20581 ( .A(n20090), .B(n20089), .Z(n20094) );
  NANDN U20582 ( .A(n20041), .B(n20040), .Z(n20045) );
  NAND U20583 ( .A(n20043), .B(n20042), .Z(n20044) );
  AND U20584 ( .A(n20045), .B(n20044), .Z(n20093) );
  XOR U20585 ( .A(n20094), .B(n20093), .Z(n20095) );
  NANDN U20586 ( .A(n20047), .B(n20046), .Z(n20051) );
  NANDN U20587 ( .A(n20049), .B(n20048), .Z(n20050) );
  NAND U20588 ( .A(n20051), .B(n20050), .Z(n20096) );
  XOR U20589 ( .A(n20095), .B(n20096), .Z(n20063) );
  OR U20590 ( .A(n20053), .B(n20052), .Z(n20057) );
  NANDN U20591 ( .A(n20055), .B(n20054), .Z(n20056) );
  NAND U20592 ( .A(n20057), .B(n20056), .Z(n20064) );
  XNOR U20593 ( .A(n20063), .B(n20064), .Z(n20065) );
  XNOR U20594 ( .A(n20066), .B(n20065), .Z(n20099) );
  XNOR U20595 ( .A(n20099), .B(sreg[1503]), .Z(n20101) );
  NAND U20596 ( .A(n20058), .B(sreg[1502]), .Z(n20062) );
  OR U20597 ( .A(n20060), .B(n20059), .Z(n20061) );
  AND U20598 ( .A(n20062), .B(n20061), .Z(n20100) );
  XOR U20599 ( .A(n20101), .B(n20100), .Z(c[1503]) );
  NANDN U20600 ( .A(n20064), .B(n20063), .Z(n20068) );
  NAND U20601 ( .A(n20066), .B(n20065), .Z(n20067) );
  NAND U20602 ( .A(n20068), .B(n20067), .Z(n20107) );
  NAND U20603 ( .A(b[0]), .B(a[488]), .Z(n20069) );
  XNOR U20604 ( .A(b[1]), .B(n20069), .Z(n20071) );
  NAND U20605 ( .A(n84), .B(a[487]), .Z(n20070) );
  AND U20606 ( .A(n20071), .B(n20070), .Z(n20124) );
  XOR U20607 ( .A(a[484]), .B(n42197), .Z(n20113) );
  NANDN U20608 ( .A(n20113), .B(n42173), .Z(n20074) );
  NANDN U20609 ( .A(n20072), .B(n42172), .Z(n20073) );
  NAND U20610 ( .A(n20074), .B(n20073), .Z(n20122) );
  NAND U20611 ( .A(b[7]), .B(a[480]), .Z(n20123) );
  XNOR U20612 ( .A(n20122), .B(n20123), .Z(n20125) );
  XOR U20613 ( .A(n20124), .B(n20125), .Z(n20131) );
  NANDN U20614 ( .A(n20075), .B(n42093), .Z(n20077) );
  XOR U20615 ( .A(n42134), .B(a[486]), .Z(n20116) );
  NANDN U20616 ( .A(n20116), .B(n42095), .Z(n20076) );
  NAND U20617 ( .A(n20077), .B(n20076), .Z(n20129) );
  NANDN U20618 ( .A(n20078), .B(n42231), .Z(n20080) );
  XOR U20619 ( .A(n202), .B(a[482]), .Z(n20119) );
  NANDN U20620 ( .A(n20119), .B(n42234), .Z(n20079) );
  AND U20621 ( .A(n20080), .B(n20079), .Z(n20128) );
  XNOR U20622 ( .A(n20129), .B(n20128), .Z(n20130) );
  XNOR U20623 ( .A(n20131), .B(n20130), .Z(n20135) );
  NANDN U20624 ( .A(n20082), .B(n20081), .Z(n20086) );
  NAND U20625 ( .A(n20084), .B(n20083), .Z(n20085) );
  AND U20626 ( .A(n20086), .B(n20085), .Z(n20134) );
  XOR U20627 ( .A(n20135), .B(n20134), .Z(n20136) );
  NANDN U20628 ( .A(n20088), .B(n20087), .Z(n20092) );
  NANDN U20629 ( .A(n20090), .B(n20089), .Z(n20091) );
  NAND U20630 ( .A(n20092), .B(n20091), .Z(n20137) );
  XOR U20631 ( .A(n20136), .B(n20137), .Z(n20104) );
  OR U20632 ( .A(n20094), .B(n20093), .Z(n20098) );
  NANDN U20633 ( .A(n20096), .B(n20095), .Z(n20097) );
  NAND U20634 ( .A(n20098), .B(n20097), .Z(n20105) );
  XNOR U20635 ( .A(n20104), .B(n20105), .Z(n20106) );
  XNOR U20636 ( .A(n20107), .B(n20106), .Z(n20140) );
  XNOR U20637 ( .A(n20140), .B(sreg[1504]), .Z(n20142) );
  NAND U20638 ( .A(n20099), .B(sreg[1503]), .Z(n20103) );
  OR U20639 ( .A(n20101), .B(n20100), .Z(n20102) );
  AND U20640 ( .A(n20103), .B(n20102), .Z(n20141) );
  XOR U20641 ( .A(n20142), .B(n20141), .Z(c[1504]) );
  NANDN U20642 ( .A(n20105), .B(n20104), .Z(n20109) );
  NAND U20643 ( .A(n20107), .B(n20106), .Z(n20108) );
  NAND U20644 ( .A(n20109), .B(n20108), .Z(n20148) );
  NAND U20645 ( .A(b[0]), .B(a[489]), .Z(n20110) );
  XNOR U20646 ( .A(b[1]), .B(n20110), .Z(n20112) );
  NAND U20647 ( .A(n84), .B(a[488]), .Z(n20111) );
  AND U20648 ( .A(n20112), .B(n20111), .Z(n20165) );
  XOR U20649 ( .A(a[485]), .B(n42197), .Z(n20154) );
  NANDN U20650 ( .A(n20154), .B(n42173), .Z(n20115) );
  NANDN U20651 ( .A(n20113), .B(n42172), .Z(n20114) );
  NAND U20652 ( .A(n20115), .B(n20114), .Z(n20163) );
  NAND U20653 ( .A(b[7]), .B(a[481]), .Z(n20164) );
  XNOR U20654 ( .A(n20163), .B(n20164), .Z(n20166) );
  XOR U20655 ( .A(n20165), .B(n20166), .Z(n20172) );
  NANDN U20656 ( .A(n20116), .B(n42093), .Z(n20118) );
  XOR U20657 ( .A(n42134), .B(a[487]), .Z(n20157) );
  NANDN U20658 ( .A(n20157), .B(n42095), .Z(n20117) );
  NAND U20659 ( .A(n20118), .B(n20117), .Z(n20170) );
  NANDN U20660 ( .A(n20119), .B(n42231), .Z(n20121) );
  XOR U20661 ( .A(n202), .B(a[483]), .Z(n20160) );
  NANDN U20662 ( .A(n20160), .B(n42234), .Z(n20120) );
  AND U20663 ( .A(n20121), .B(n20120), .Z(n20169) );
  XNOR U20664 ( .A(n20170), .B(n20169), .Z(n20171) );
  XNOR U20665 ( .A(n20172), .B(n20171), .Z(n20176) );
  NANDN U20666 ( .A(n20123), .B(n20122), .Z(n20127) );
  NAND U20667 ( .A(n20125), .B(n20124), .Z(n20126) );
  AND U20668 ( .A(n20127), .B(n20126), .Z(n20175) );
  XOR U20669 ( .A(n20176), .B(n20175), .Z(n20177) );
  NANDN U20670 ( .A(n20129), .B(n20128), .Z(n20133) );
  NANDN U20671 ( .A(n20131), .B(n20130), .Z(n20132) );
  NAND U20672 ( .A(n20133), .B(n20132), .Z(n20178) );
  XOR U20673 ( .A(n20177), .B(n20178), .Z(n20145) );
  OR U20674 ( .A(n20135), .B(n20134), .Z(n20139) );
  NANDN U20675 ( .A(n20137), .B(n20136), .Z(n20138) );
  NAND U20676 ( .A(n20139), .B(n20138), .Z(n20146) );
  XNOR U20677 ( .A(n20145), .B(n20146), .Z(n20147) );
  XNOR U20678 ( .A(n20148), .B(n20147), .Z(n20181) );
  XNOR U20679 ( .A(n20181), .B(sreg[1505]), .Z(n20183) );
  NAND U20680 ( .A(n20140), .B(sreg[1504]), .Z(n20144) );
  OR U20681 ( .A(n20142), .B(n20141), .Z(n20143) );
  AND U20682 ( .A(n20144), .B(n20143), .Z(n20182) );
  XOR U20683 ( .A(n20183), .B(n20182), .Z(c[1505]) );
  NANDN U20684 ( .A(n20146), .B(n20145), .Z(n20150) );
  NAND U20685 ( .A(n20148), .B(n20147), .Z(n20149) );
  NAND U20686 ( .A(n20150), .B(n20149), .Z(n20189) );
  NAND U20687 ( .A(b[0]), .B(a[490]), .Z(n20151) );
  XNOR U20688 ( .A(b[1]), .B(n20151), .Z(n20153) );
  NAND U20689 ( .A(n85), .B(a[489]), .Z(n20152) );
  AND U20690 ( .A(n20153), .B(n20152), .Z(n20206) );
  XOR U20691 ( .A(a[486]), .B(n42197), .Z(n20195) );
  NANDN U20692 ( .A(n20195), .B(n42173), .Z(n20156) );
  NANDN U20693 ( .A(n20154), .B(n42172), .Z(n20155) );
  NAND U20694 ( .A(n20156), .B(n20155), .Z(n20204) );
  NAND U20695 ( .A(b[7]), .B(a[482]), .Z(n20205) );
  XNOR U20696 ( .A(n20204), .B(n20205), .Z(n20207) );
  XOR U20697 ( .A(n20206), .B(n20207), .Z(n20213) );
  NANDN U20698 ( .A(n20157), .B(n42093), .Z(n20159) );
  XOR U20699 ( .A(n42134), .B(a[488]), .Z(n20198) );
  NANDN U20700 ( .A(n20198), .B(n42095), .Z(n20158) );
  NAND U20701 ( .A(n20159), .B(n20158), .Z(n20211) );
  NANDN U20702 ( .A(n20160), .B(n42231), .Z(n20162) );
  XOR U20703 ( .A(n202), .B(a[484]), .Z(n20201) );
  NANDN U20704 ( .A(n20201), .B(n42234), .Z(n20161) );
  AND U20705 ( .A(n20162), .B(n20161), .Z(n20210) );
  XNOR U20706 ( .A(n20211), .B(n20210), .Z(n20212) );
  XNOR U20707 ( .A(n20213), .B(n20212), .Z(n20217) );
  NANDN U20708 ( .A(n20164), .B(n20163), .Z(n20168) );
  NAND U20709 ( .A(n20166), .B(n20165), .Z(n20167) );
  AND U20710 ( .A(n20168), .B(n20167), .Z(n20216) );
  XOR U20711 ( .A(n20217), .B(n20216), .Z(n20218) );
  NANDN U20712 ( .A(n20170), .B(n20169), .Z(n20174) );
  NANDN U20713 ( .A(n20172), .B(n20171), .Z(n20173) );
  NAND U20714 ( .A(n20174), .B(n20173), .Z(n20219) );
  XOR U20715 ( .A(n20218), .B(n20219), .Z(n20186) );
  OR U20716 ( .A(n20176), .B(n20175), .Z(n20180) );
  NANDN U20717 ( .A(n20178), .B(n20177), .Z(n20179) );
  NAND U20718 ( .A(n20180), .B(n20179), .Z(n20187) );
  XNOR U20719 ( .A(n20186), .B(n20187), .Z(n20188) );
  XNOR U20720 ( .A(n20189), .B(n20188), .Z(n20222) );
  XNOR U20721 ( .A(n20222), .B(sreg[1506]), .Z(n20224) );
  NAND U20722 ( .A(n20181), .B(sreg[1505]), .Z(n20185) );
  OR U20723 ( .A(n20183), .B(n20182), .Z(n20184) );
  AND U20724 ( .A(n20185), .B(n20184), .Z(n20223) );
  XOR U20725 ( .A(n20224), .B(n20223), .Z(c[1506]) );
  NANDN U20726 ( .A(n20187), .B(n20186), .Z(n20191) );
  NAND U20727 ( .A(n20189), .B(n20188), .Z(n20190) );
  NAND U20728 ( .A(n20191), .B(n20190), .Z(n20230) );
  NAND U20729 ( .A(b[0]), .B(a[491]), .Z(n20192) );
  XNOR U20730 ( .A(b[1]), .B(n20192), .Z(n20194) );
  NAND U20731 ( .A(n85), .B(a[490]), .Z(n20193) );
  AND U20732 ( .A(n20194), .B(n20193), .Z(n20247) );
  XOR U20733 ( .A(a[487]), .B(n42197), .Z(n20236) );
  NANDN U20734 ( .A(n20236), .B(n42173), .Z(n20197) );
  NANDN U20735 ( .A(n20195), .B(n42172), .Z(n20196) );
  NAND U20736 ( .A(n20197), .B(n20196), .Z(n20245) );
  NAND U20737 ( .A(b[7]), .B(a[483]), .Z(n20246) );
  XNOR U20738 ( .A(n20245), .B(n20246), .Z(n20248) );
  XOR U20739 ( .A(n20247), .B(n20248), .Z(n20254) );
  NANDN U20740 ( .A(n20198), .B(n42093), .Z(n20200) );
  XOR U20741 ( .A(n42134), .B(a[489]), .Z(n20239) );
  NANDN U20742 ( .A(n20239), .B(n42095), .Z(n20199) );
  NAND U20743 ( .A(n20200), .B(n20199), .Z(n20252) );
  NANDN U20744 ( .A(n20201), .B(n42231), .Z(n20203) );
  XOR U20745 ( .A(n202), .B(a[485]), .Z(n20242) );
  NANDN U20746 ( .A(n20242), .B(n42234), .Z(n20202) );
  AND U20747 ( .A(n20203), .B(n20202), .Z(n20251) );
  XNOR U20748 ( .A(n20252), .B(n20251), .Z(n20253) );
  XNOR U20749 ( .A(n20254), .B(n20253), .Z(n20258) );
  NANDN U20750 ( .A(n20205), .B(n20204), .Z(n20209) );
  NAND U20751 ( .A(n20207), .B(n20206), .Z(n20208) );
  AND U20752 ( .A(n20209), .B(n20208), .Z(n20257) );
  XOR U20753 ( .A(n20258), .B(n20257), .Z(n20259) );
  NANDN U20754 ( .A(n20211), .B(n20210), .Z(n20215) );
  NANDN U20755 ( .A(n20213), .B(n20212), .Z(n20214) );
  NAND U20756 ( .A(n20215), .B(n20214), .Z(n20260) );
  XOR U20757 ( .A(n20259), .B(n20260), .Z(n20227) );
  OR U20758 ( .A(n20217), .B(n20216), .Z(n20221) );
  NANDN U20759 ( .A(n20219), .B(n20218), .Z(n20220) );
  NAND U20760 ( .A(n20221), .B(n20220), .Z(n20228) );
  XNOR U20761 ( .A(n20227), .B(n20228), .Z(n20229) );
  XNOR U20762 ( .A(n20230), .B(n20229), .Z(n20263) );
  XNOR U20763 ( .A(n20263), .B(sreg[1507]), .Z(n20265) );
  NAND U20764 ( .A(n20222), .B(sreg[1506]), .Z(n20226) );
  OR U20765 ( .A(n20224), .B(n20223), .Z(n20225) );
  AND U20766 ( .A(n20226), .B(n20225), .Z(n20264) );
  XOR U20767 ( .A(n20265), .B(n20264), .Z(c[1507]) );
  NANDN U20768 ( .A(n20228), .B(n20227), .Z(n20232) );
  NAND U20769 ( .A(n20230), .B(n20229), .Z(n20231) );
  NAND U20770 ( .A(n20232), .B(n20231), .Z(n20271) );
  NAND U20771 ( .A(b[0]), .B(a[492]), .Z(n20233) );
  XNOR U20772 ( .A(b[1]), .B(n20233), .Z(n20235) );
  NAND U20773 ( .A(n85), .B(a[491]), .Z(n20234) );
  AND U20774 ( .A(n20235), .B(n20234), .Z(n20288) );
  XOR U20775 ( .A(a[488]), .B(n42197), .Z(n20277) );
  NANDN U20776 ( .A(n20277), .B(n42173), .Z(n20238) );
  NANDN U20777 ( .A(n20236), .B(n42172), .Z(n20237) );
  NAND U20778 ( .A(n20238), .B(n20237), .Z(n20286) );
  NAND U20779 ( .A(b[7]), .B(a[484]), .Z(n20287) );
  XNOR U20780 ( .A(n20286), .B(n20287), .Z(n20289) );
  XOR U20781 ( .A(n20288), .B(n20289), .Z(n20295) );
  NANDN U20782 ( .A(n20239), .B(n42093), .Z(n20241) );
  XOR U20783 ( .A(n42134), .B(a[490]), .Z(n20280) );
  NANDN U20784 ( .A(n20280), .B(n42095), .Z(n20240) );
  NAND U20785 ( .A(n20241), .B(n20240), .Z(n20293) );
  NANDN U20786 ( .A(n20242), .B(n42231), .Z(n20244) );
  XOR U20787 ( .A(n202), .B(a[486]), .Z(n20283) );
  NANDN U20788 ( .A(n20283), .B(n42234), .Z(n20243) );
  AND U20789 ( .A(n20244), .B(n20243), .Z(n20292) );
  XNOR U20790 ( .A(n20293), .B(n20292), .Z(n20294) );
  XNOR U20791 ( .A(n20295), .B(n20294), .Z(n20299) );
  NANDN U20792 ( .A(n20246), .B(n20245), .Z(n20250) );
  NAND U20793 ( .A(n20248), .B(n20247), .Z(n20249) );
  AND U20794 ( .A(n20250), .B(n20249), .Z(n20298) );
  XOR U20795 ( .A(n20299), .B(n20298), .Z(n20300) );
  NANDN U20796 ( .A(n20252), .B(n20251), .Z(n20256) );
  NANDN U20797 ( .A(n20254), .B(n20253), .Z(n20255) );
  NAND U20798 ( .A(n20256), .B(n20255), .Z(n20301) );
  XOR U20799 ( .A(n20300), .B(n20301), .Z(n20268) );
  OR U20800 ( .A(n20258), .B(n20257), .Z(n20262) );
  NANDN U20801 ( .A(n20260), .B(n20259), .Z(n20261) );
  NAND U20802 ( .A(n20262), .B(n20261), .Z(n20269) );
  XNOR U20803 ( .A(n20268), .B(n20269), .Z(n20270) );
  XNOR U20804 ( .A(n20271), .B(n20270), .Z(n20304) );
  XNOR U20805 ( .A(n20304), .B(sreg[1508]), .Z(n20306) );
  NAND U20806 ( .A(n20263), .B(sreg[1507]), .Z(n20267) );
  OR U20807 ( .A(n20265), .B(n20264), .Z(n20266) );
  AND U20808 ( .A(n20267), .B(n20266), .Z(n20305) );
  XOR U20809 ( .A(n20306), .B(n20305), .Z(c[1508]) );
  NANDN U20810 ( .A(n20269), .B(n20268), .Z(n20273) );
  NAND U20811 ( .A(n20271), .B(n20270), .Z(n20272) );
  NAND U20812 ( .A(n20273), .B(n20272), .Z(n20312) );
  NAND U20813 ( .A(b[0]), .B(a[493]), .Z(n20274) );
  XNOR U20814 ( .A(b[1]), .B(n20274), .Z(n20276) );
  NAND U20815 ( .A(n85), .B(a[492]), .Z(n20275) );
  AND U20816 ( .A(n20276), .B(n20275), .Z(n20329) );
  XOR U20817 ( .A(a[489]), .B(n42197), .Z(n20318) );
  NANDN U20818 ( .A(n20318), .B(n42173), .Z(n20279) );
  NANDN U20819 ( .A(n20277), .B(n42172), .Z(n20278) );
  NAND U20820 ( .A(n20279), .B(n20278), .Z(n20327) );
  NAND U20821 ( .A(b[7]), .B(a[485]), .Z(n20328) );
  XNOR U20822 ( .A(n20327), .B(n20328), .Z(n20330) );
  XOR U20823 ( .A(n20329), .B(n20330), .Z(n20336) );
  NANDN U20824 ( .A(n20280), .B(n42093), .Z(n20282) );
  XOR U20825 ( .A(n42134), .B(a[491]), .Z(n20321) );
  NANDN U20826 ( .A(n20321), .B(n42095), .Z(n20281) );
  NAND U20827 ( .A(n20282), .B(n20281), .Z(n20334) );
  NANDN U20828 ( .A(n20283), .B(n42231), .Z(n20285) );
  XOR U20829 ( .A(n202), .B(a[487]), .Z(n20324) );
  NANDN U20830 ( .A(n20324), .B(n42234), .Z(n20284) );
  AND U20831 ( .A(n20285), .B(n20284), .Z(n20333) );
  XNOR U20832 ( .A(n20334), .B(n20333), .Z(n20335) );
  XNOR U20833 ( .A(n20336), .B(n20335), .Z(n20340) );
  NANDN U20834 ( .A(n20287), .B(n20286), .Z(n20291) );
  NAND U20835 ( .A(n20289), .B(n20288), .Z(n20290) );
  AND U20836 ( .A(n20291), .B(n20290), .Z(n20339) );
  XOR U20837 ( .A(n20340), .B(n20339), .Z(n20341) );
  NANDN U20838 ( .A(n20293), .B(n20292), .Z(n20297) );
  NANDN U20839 ( .A(n20295), .B(n20294), .Z(n20296) );
  NAND U20840 ( .A(n20297), .B(n20296), .Z(n20342) );
  XOR U20841 ( .A(n20341), .B(n20342), .Z(n20309) );
  OR U20842 ( .A(n20299), .B(n20298), .Z(n20303) );
  NANDN U20843 ( .A(n20301), .B(n20300), .Z(n20302) );
  NAND U20844 ( .A(n20303), .B(n20302), .Z(n20310) );
  XNOR U20845 ( .A(n20309), .B(n20310), .Z(n20311) );
  XNOR U20846 ( .A(n20312), .B(n20311), .Z(n20345) );
  XNOR U20847 ( .A(n20345), .B(sreg[1509]), .Z(n20347) );
  NAND U20848 ( .A(n20304), .B(sreg[1508]), .Z(n20308) );
  OR U20849 ( .A(n20306), .B(n20305), .Z(n20307) );
  AND U20850 ( .A(n20308), .B(n20307), .Z(n20346) );
  XOR U20851 ( .A(n20347), .B(n20346), .Z(c[1509]) );
  NANDN U20852 ( .A(n20310), .B(n20309), .Z(n20314) );
  NAND U20853 ( .A(n20312), .B(n20311), .Z(n20313) );
  NAND U20854 ( .A(n20314), .B(n20313), .Z(n20353) );
  NAND U20855 ( .A(b[0]), .B(a[494]), .Z(n20315) );
  XNOR U20856 ( .A(b[1]), .B(n20315), .Z(n20317) );
  NAND U20857 ( .A(n85), .B(a[493]), .Z(n20316) );
  AND U20858 ( .A(n20317), .B(n20316), .Z(n20370) );
  XOR U20859 ( .A(a[490]), .B(n42197), .Z(n20359) );
  NANDN U20860 ( .A(n20359), .B(n42173), .Z(n20320) );
  NANDN U20861 ( .A(n20318), .B(n42172), .Z(n20319) );
  NAND U20862 ( .A(n20320), .B(n20319), .Z(n20368) );
  NAND U20863 ( .A(b[7]), .B(a[486]), .Z(n20369) );
  XNOR U20864 ( .A(n20368), .B(n20369), .Z(n20371) );
  XOR U20865 ( .A(n20370), .B(n20371), .Z(n20377) );
  NANDN U20866 ( .A(n20321), .B(n42093), .Z(n20323) );
  XOR U20867 ( .A(n42134), .B(a[492]), .Z(n20362) );
  NANDN U20868 ( .A(n20362), .B(n42095), .Z(n20322) );
  NAND U20869 ( .A(n20323), .B(n20322), .Z(n20375) );
  NANDN U20870 ( .A(n20324), .B(n42231), .Z(n20326) );
  XOR U20871 ( .A(n202), .B(a[488]), .Z(n20365) );
  NANDN U20872 ( .A(n20365), .B(n42234), .Z(n20325) );
  AND U20873 ( .A(n20326), .B(n20325), .Z(n20374) );
  XNOR U20874 ( .A(n20375), .B(n20374), .Z(n20376) );
  XNOR U20875 ( .A(n20377), .B(n20376), .Z(n20381) );
  NANDN U20876 ( .A(n20328), .B(n20327), .Z(n20332) );
  NAND U20877 ( .A(n20330), .B(n20329), .Z(n20331) );
  AND U20878 ( .A(n20332), .B(n20331), .Z(n20380) );
  XOR U20879 ( .A(n20381), .B(n20380), .Z(n20382) );
  NANDN U20880 ( .A(n20334), .B(n20333), .Z(n20338) );
  NANDN U20881 ( .A(n20336), .B(n20335), .Z(n20337) );
  NAND U20882 ( .A(n20338), .B(n20337), .Z(n20383) );
  XOR U20883 ( .A(n20382), .B(n20383), .Z(n20350) );
  OR U20884 ( .A(n20340), .B(n20339), .Z(n20344) );
  NANDN U20885 ( .A(n20342), .B(n20341), .Z(n20343) );
  NAND U20886 ( .A(n20344), .B(n20343), .Z(n20351) );
  XNOR U20887 ( .A(n20350), .B(n20351), .Z(n20352) );
  XNOR U20888 ( .A(n20353), .B(n20352), .Z(n20386) );
  XNOR U20889 ( .A(n20386), .B(sreg[1510]), .Z(n20388) );
  NAND U20890 ( .A(n20345), .B(sreg[1509]), .Z(n20349) );
  OR U20891 ( .A(n20347), .B(n20346), .Z(n20348) );
  AND U20892 ( .A(n20349), .B(n20348), .Z(n20387) );
  XOR U20893 ( .A(n20388), .B(n20387), .Z(c[1510]) );
  NANDN U20894 ( .A(n20351), .B(n20350), .Z(n20355) );
  NAND U20895 ( .A(n20353), .B(n20352), .Z(n20354) );
  NAND U20896 ( .A(n20355), .B(n20354), .Z(n20394) );
  NAND U20897 ( .A(b[0]), .B(a[495]), .Z(n20356) );
  XNOR U20898 ( .A(b[1]), .B(n20356), .Z(n20358) );
  NAND U20899 ( .A(n85), .B(a[494]), .Z(n20357) );
  AND U20900 ( .A(n20358), .B(n20357), .Z(n20411) );
  XOR U20901 ( .A(a[491]), .B(n42197), .Z(n20400) );
  NANDN U20902 ( .A(n20400), .B(n42173), .Z(n20361) );
  NANDN U20903 ( .A(n20359), .B(n42172), .Z(n20360) );
  NAND U20904 ( .A(n20361), .B(n20360), .Z(n20409) );
  NAND U20905 ( .A(b[7]), .B(a[487]), .Z(n20410) );
  XNOR U20906 ( .A(n20409), .B(n20410), .Z(n20412) );
  XOR U20907 ( .A(n20411), .B(n20412), .Z(n20418) );
  NANDN U20908 ( .A(n20362), .B(n42093), .Z(n20364) );
  XOR U20909 ( .A(n42134), .B(a[493]), .Z(n20403) );
  NANDN U20910 ( .A(n20403), .B(n42095), .Z(n20363) );
  NAND U20911 ( .A(n20364), .B(n20363), .Z(n20416) );
  NANDN U20912 ( .A(n20365), .B(n42231), .Z(n20367) );
  XOR U20913 ( .A(n202), .B(a[489]), .Z(n20406) );
  NANDN U20914 ( .A(n20406), .B(n42234), .Z(n20366) );
  AND U20915 ( .A(n20367), .B(n20366), .Z(n20415) );
  XNOR U20916 ( .A(n20416), .B(n20415), .Z(n20417) );
  XNOR U20917 ( .A(n20418), .B(n20417), .Z(n20422) );
  NANDN U20918 ( .A(n20369), .B(n20368), .Z(n20373) );
  NAND U20919 ( .A(n20371), .B(n20370), .Z(n20372) );
  AND U20920 ( .A(n20373), .B(n20372), .Z(n20421) );
  XOR U20921 ( .A(n20422), .B(n20421), .Z(n20423) );
  NANDN U20922 ( .A(n20375), .B(n20374), .Z(n20379) );
  NANDN U20923 ( .A(n20377), .B(n20376), .Z(n20378) );
  NAND U20924 ( .A(n20379), .B(n20378), .Z(n20424) );
  XOR U20925 ( .A(n20423), .B(n20424), .Z(n20391) );
  OR U20926 ( .A(n20381), .B(n20380), .Z(n20385) );
  NANDN U20927 ( .A(n20383), .B(n20382), .Z(n20384) );
  NAND U20928 ( .A(n20385), .B(n20384), .Z(n20392) );
  XNOR U20929 ( .A(n20391), .B(n20392), .Z(n20393) );
  XNOR U20930 ( .A(n20394), .B(n20393), .Z(n20427) );
  XNOR U20931 ( .A(n20427), .B(sreg[1511]), .Z(n20429) );
  NAND U20932 ( .A(n20386), .B(sreg[1510]), .Z(n20390) );
  OR U20933 ( .A(n20388), .B(n20387), .Z(n20389) );
  AND U20934 ( .A(n20390), .B(n20389), .Z(n20428) );
  XOR U20935 ( .A(n20429), .B(n20428), .Z(c[1511]) );
  NANDN U20936 ( .A(n20392), .B(n20391), .Z(n20396) );
  NAND U20937 ( .A(n20394), .B(n20393), .Z(n20395) );
  NAND U20938 ( .A(n20396), .B(n20395), .Z(n20435) );
  NAND U20939 ( .A(b[0]), .B(a[496]), .Z(n20397) );
  XNOR U20940 ( .A(b[1]), .B(n20397), .Z(n20399) );
  NAND U20941 ( .A(n85), .B(a[495]), .Z(n20398) );
  AND U20942 ( .A(n20399), .B(n20398), .Z(n20452) );
  XOR U20943 ( .A(a[492]), .B(n42197), .Z(n20441) );
  NANDN U20944 ( .A(n20441), .B(n42173), .Z(n20402) );
  NANDN U20945 ( .A(n20400), .B(n42172), .Z(n20401) );
  NAND U20946 ( .A(n20402), .B(n20401), .Z(n20450) );
  NAND U20947 ( .A(b[7]), .B(a[488]), .Z(n20451) );
  XNOR U20948 ( .A(n20450), .B(n20451), .Z(n20453) );
  XOR U20949 ( .A(n20452), .B(n20453), .Z(n20459) );
  NANDN U20950 ( .A(n20403), .B(n42093), .Z(n20405) );
  XOR U20951 ( .A(n42134), .B(a[494]), .Z(n20444) );
  NANDN U20952 ( .A(n20444), .B(n42095), .Z(n20404) );
  NAND U20953 ( .A(n20405), .B(n20404), .Z(n20457) );
  NANDN U20954 ( .A(n20406), .B(n42231), .Z(n20408) );
  XOR U20955 ( .A(n202), .B(a[490]), .Z(n20447) );
  NANDN U20956 ( .A(n20447), .B(n42234), .Z(n20407) );
  AND U20957 ( .A(n20408), .B(n20407), .Z(n20456) );
  XNOR U20958 ( .A(n20457), .B(n20456), .Z(n20458) );
  XNOR U20959 ( .A(n20459), .B(n20458), .Z(n20463) );
  NANDN U20960 ( .A(n20410), .B(n20409), .Z(n20414) );
  NAND U20961 ( .A(n20412), .B(n20411), .Z(n20413) );
  AND U20962 ( .A(n20414), .B(n20413), .Z(n20462) );
  XOR U20963 ( .A(n20463), .B(n20462), .Z(n20464) );
  NANDN U20964 ( .A(n20416), .B(n20415), .Z(n20420) );
  NANDN U20965 ( .A(n20418), .B(n20417), .Z(n20419) );
  NAND U20966 ( .A(n20420), .B(n20419), .Z(n20465) );
  XOR U20967 ( .A(n20464), .B(n20465), .Z(n20432) );
  OR U20968 ( .A(n20422), .B(n20421), .Z(n20426) );
  NANDN U20969 ( .A(n20424), .B(n20423), .Z(n20425) );
  NAND U20970 ( .A(n20426), .B(n20425), .Z(n20433) );
  XNOR U20971 ( .A(n20432), .B(n20433), .Z(n20434) );
  XNOR U20972 ( .A(n20435), .B(n20434), .Z(n20468) );
  XNOR U20973 ( .A(n20468), .B(sreg[1512]), .Z(n20470) );
  NAND U20974 ( .A(n20427), .B(sreg[1511]), .Z(n20431) );
  OR U20975 ( .A(n20429), .B(n20428), .Z(n20430) );
  AND U20976 ( .A(n20431), .B(n20430), .Z(n20469) );
  XOR U20977 ( .A(n20470), .B(n20469), .Z(c[1512]) );
  NANDN U20978 ( .A(n20433), .B(n20432), .Z(n20437) );
  NAND U20979 ( .A(n20435), .B(n20434), .Z(n20436) );
  NAND U20980 ( .A(n20437), .B(n20436), .Z(n20476) );
  NAND U20981 ( .A(b[0]), .B(a[497]), .Z(n20438) );
  XNOR U20982 ( .A(b[1]), .B(n20438), .Z(n20440) );
  NAND U20983 ( .A(n86), .B(a[496]), .Z(n20439) );
  AND U20984 ( .A(n20440), .B(n20439), .Z(n20493) );
  XOR U20985 ( .A(a[493]), .B(n42197), .Z(n20482) );
  NANDN U20986 ( .A(n20482), .B(n42173), .Z(n20443) );
  NANDN U20987 ( .A(n20441), .B(n42172), .Z(n20442) );
  NAND U20988 ( .A(n20443), .B(n20442), .Z(n20491) );
  NAND U20989 ( .A(b[7]), .B(a[489]), .Z(n20492) );
  XNOR U20990 ( .A(n20491), .B(n20492), .Z(n20494) );
  XOR U20991 ( .A(n20493), .B(n20494), .Z(n20500) );
  NANDN U20992 ( .A(n20444), .B(n42093), .Z(n20446) );
  XOR U20993 ( .A(n42134), .B(a[495]), .Z(n20485) );
  NANDN U20994 ( .A(n20485), .B(n42095), .Z(n20445) );
  NAND U20995 ( .A(n20446), .B(n20445), .Z(n20498) );
  NANDN U20996 ( .A(n20447), .B(n42231), .Z(n20449) );
  XOR U20997 ( .A(n203), .B(a[491]), .Z(n20488) );
  NANDN U20998 ( .A(n20488), .B(n42234), .Z(n20448) );
  AND U20999 ( .A(n20449), .B(n20448), .Z(n20497) );
  XNOR U21000 ( .A(n20498), .B(n20497), .Z(n20499) );
  XNOR U21001 ( .A(n20500), .B(n20499), .Z(n20504) );
  NANDN U21002 ( .A(n20451), .B(n20450), .Z(n20455) );
  NAND U21003 ( .A(n20453), .B(n20452), .Z(n20454) );
  AND U21004 ( .A(n20455), .B(n20454), .Z(n20503) );
  XOR U21005 ( .A(n20504), .B(n20503), .Z(n20505) );
  NANDN U21006 ( .A(n20457), .B(n20456), .Z(n20461) );
  NANDN U21007 ( .A(n20459), .B(n20458), .Z(n20460) );
  NAND U21008 ( .A(n20461), .B(n20460), .Z(n20506) );
  XOR U21009 ( .A(n20505), .B(n20506), .Z(n20473) );
  OR U21010 ( .A(n20463), .B(n20462), .Z(n20467) );
  NANDN U21011 ( .A(n20465), .B(n20464), .Z(n20466) );
  NAND U21012 ( .A(n20467), .B(n20466), .Z(n20474) );
  XNOR U21013 ( .A(n20473), .B(n20474), .Z(n20475) );
  XNOR U21014 ( .A(n20476), .B(n20475), .Z(n20509) );
  XNOR U21015 ( .A(n20509), .B(sreg[1513]), .Z(n20511) );
  NAND U21016 ( .A(n20468), .B(sreg[1512]), .Z(n20472) );
  OR U21017 ( .A(n20470), .B(n20469), .Z(n20471) );
  AND U21018 ( .A(n20472), .B(n20471), .Z(n20510) );
  XOR U21019 ( .A(n20511), .B(n20510), .Z(c[1513]) );
  NANDN U21020 ( .A(n20474), .B(n20473), .Z(n20478) );
  NAND U21021 ( .A(n20476), .B(n20475), .Z(n20477) );
  NAND U21022 ( .A(n20478), .B(n20477), .Z(n20517) );
  NAND U21023 ( .A(b[0]), .B(a[498]), .Z(n20479) );
  XNOR U21024 ( .A(b[1]), .B(n20479), .Z(n20481) );
  NAND U21025 ( .A(n86), .B(a[497]), .Z(n20480) );
  AND U21026 ( .A(n20481), .B(n20480), .Z(n20534) );
  XOR U21027 ( .A(a[494]), .B(n42197), .Z(n20523) );
  NANDN U21028 ( .A(n20523), .B(n42173), .Z(n20484) );
  NANDN U21029 ( .A(n20482), .B(n42172), .Z(n20483) );
  NAND U21030 ( .A(n20484), .B(n20483), .Z(n20532) );
  NAND U21031 ( .A(b[7]), .B(a[490]), .Z(n20533) );
  XNOR U21032 ( .A(n20532), .B(n20533), .Z(n20535) );
  XOR U21033 ( .A(n20534), .B(n20535), .Z(n20541) );
  NANDN U21034 ( .A(n20485), .B(n42093), .Z(n20487) );
  XOR U21035 ( .A(n42134), .B(a[496]), .Z(n20526) );
  NANDN U21036 ( .A(n20526), .B(n42095), .Z(n20486) );
  NAND U21037 ( .A(n20487), .B(n20486), .Z(n20539) );
  NANDN U21038 ( .A(n20488), .B(n42231), .Z(n20490) );
  XOR U21039 ( .A(n203), .B(a[492]), .Z(n20529) );
  NANDN U21040 ( .A(n20529), .B(n42234), .Z(n20489) );
  AND U21041 ( .A(n20490), .B(n20489), .Z(n20538) );
  XNOR U21042 ( .A(n20539), .B(n20538), .Z(n20540) );
  XNOR U21043 ( .A(n20541), .B(n20540), .Z(n20545) );
  NANDN U21044 ( .A(n20492), .B(n20491), .Z(n20496) );
  NAND U21045 ( .A(n20494), .B(n20493), .Z(n20495) );
  AND U21046 ( .A(n20496), .B(n20495), .Z(n20544) );
  XOR U21047 ( .A(n20545), .B(n20544), .Z(n20546) );
  NANDN U21048 ( .A(n20498), .B(n20497), .Z(n20502) );
  NANDN U21049 ( .A(n20500), .B(n20499), .Z(n20501) );
  NAND U21050 ( .A(n20502), .B(n20501), .Z(n20547) );
  XOR U21051 ( .A(n20546), .B(n20547), .Z(n20514) );
  OR U21052 ( .A(n20504), .B(n20503), .Z(n20508) );
  NANDN U21053 ( .A(n20506), .B(n20505), .Z(n20507) );
  NAND U21054 ( .A(n20508), .B(n20507), .Z(n20515) );
  XNOR U21055 ( .A(n20514), .B(n20515), .Z(n20516) );
  XNOR U21056 ( .A(n20517), .B(n20516), .Z(n20550) );
  XNOR U21057 ( .A(n20550), .B(sreg[1514]), .Z(n20552) );
  NAND U21058 ( .A(n20509), .B(sreg[1513]), .Z(n20513) );
  OR U21059 ( .A(n20511), .B(n20510), .Z(n20512) );
  AND U21060 ( .A(n20513), .B(n20512), .Z(n20551) );
  XOR U21061 ( .A(n20552), .B(n20551), .Z(c[1514]) );
  NANDN U21062 ( .A(n20515), .B(n20514), .Z(n20519) );
  NAND U21063 ( .A(n20517), .B(n20516), .Z(n20518) );
  NAND U21064 ( .A(n20519), .B(n20518), .Z(n20558) );
  NAND U21065 ( .A(b[0]), .B(a[499]), .Z(n20520) );
  XNOR U21066 ( .A(b[1]), .B(n20520), .Z(n20522) );
  NAND U21067 ( .A(n86), .B(a[498]), .Z(n20521) );
  AND U21068 ( .A(n20522), .B(n20521), .Z(n20575) );
  XOR U21069 ( .A(a[495]), .B(n42197), .Z(n20564) );
  NANDN U21070 ( .A(n20564), .B(n42173), .Z(n20525) );
  NANDN U21071 ( .A(n20523), .B(n42172), .Z(n20524) );
  NAND U21072 ( .A(n20525), .B(n20524), .Z(n20573) );
  NAND U21073 ( .A(b[7]), .B(a[491]), .Z(n20574) );
  XNOR U21074 ( .A(n20573), .B(n20574), .Z(n20576) );
  XOR U21075 ( .A(n20575), .B(n20576), .Z(n20582) );
  NANDN U21076 ( .A(n20526), .B(n42093), .Z(n20528) );
  XOR U21077 ( .A(n42134), .B(a[497]), .Z(n20567) );
  NANDN U21078 ( .A(n20567), .B(n42095), .Z(n20527) );
  NAND U21079 ( .A(n20528), .B(n20527), .Z(n20580) );
  NANDN U21080 ( .A(n20529), .B(n42231), .Z(n20531) );
  XOR U21081 ( .A(n203), .B(a[493]), .Z(n20570) );
  NANDN U21082 ( .A(n20570), .B(n42234), .Z(n20530) );
  AND U21083 ( .A(n20531), .B(n20530), .Z(n20579) );
  XNOR U21084 ( .A(n20580), .B(n20579), .Z(n20581) );
  XNOR U21085 ( .A(n20582), .B(n20581), .Z(n20586) );
  NANDN U21086 ( .A(n20533), .B(n20532), .Z(n20537) );
  NAND U21087 ( .A(n20535), .B(n20534), .Z(n20536) );
  AND U21088 ( .A(n20537), .B(n20536), .Z(n20585) );
  XOR U21089 ( .A(n20586), .B(n20585), .Z(n20587) );
  NANDN U21090 ( .A(n20539), .B(n20538), .Z(n20543) );
  NANDN U21091 ( .A(n20541), .B(n20540), .Z(n20542) );
  NAND U21092 ( .A(n20543), .B(n20542), .Z(n20588) );
  XOR U21093 ( .A(n20587), .B(n20588), .Z(n20555) );
  OR U21094 ( .A(n20545), .B(n20544), .Z(n20549) );
  NANDN U21095 ( .A(n20547), .B(n20546), .Z(n20548) );
  NAND U21096 ( .A(n20549), .B(n20548), .Z(n20556) );
  XNOR U21097 ( .A(n20555), .B(n20556), .Z(n20557) );
  XNOR U21098 ( .A(n20558), .B(n20557), .Z(n20591) );
  XNOR U21099 ( .A(n20591), .B(sreg[1515]), .Z(n20593) );
  NAND U21100 ( .A(n20550), .B(sreg[1514]), .Z(n20554) );
  OR U21101 ( .A(n20552), .B(n20551), .Z(n20553) );
  AND U21102 ( .A(n20554), .B(n20553), .Z(n20592) );
  XOR U21103 ( .A(n20593), .B(n20592), .Z(c[1515]) );
  NANDN U21104 ( .A(n20556), .B(n20555), .Z(n20560) );
  NAND U21105 ( .A(n20558), .B(n20557), .Z(n20559) );
  NAND U21106 ( .A(n20560), .B(n20559), .Z(n20599) );
  NAND U21107 ( .A(b[0]), .B(a[500]), .Z(n20561) );
  XNOR U21108 ( .A(b[1]), .B(n20561), .Z(n20563) );
  NAND U21109 ( .A(n86), .B(a[499]), .Z(n20562) );
  AND U21110 ( .A(n20563), .B(n20562), .Z(n20616) );
  XOR U21111 ( .A(a[496]), .B(n42197), .Z(n20605) );
  NANDN U21112 ( .A(n20605), .B(n42173), .Z(n20566) );
  NANDN U21113 ( .A(n20564), .B(n42172), .Z(n20565) );
  NAND U21114 ( .A(n20566), .B(n20565), .Z(n20614) );
  NAND U21115 ( .A(b[7]), .B(a[492]), .Z(n20615) );
  XNOR U21116 ( .A(n20614), .B(n20615), .Z(n20617) );
  XOR U21117 ( .A(n20616), .B(n20617), .Z(n20623) );
  NANDN U21118 ( .A(n20567), .B(n42093), .Z(n20569) );
  XOR U21119 ( .A(n42134), .B(a[498]), .Z(n20608) );
  NANDN U21120 ( .A(n20608), .B(n42095), .Z(n20568) );
  NAND U21121 ( .A(n20569), .B(n20568), .Z(n20621) );
  NANDN U21122 ( .A(n20570), .B(n42231), .Z(n20572) );
  XOR U21123 ( .A(n203), .B(a[494]), .Z(n20611) );
  NANDN U21124 ( .A(n20611), .B(n42234), .Z(n20571) );
  AND U21125 ( .A(n20572), .B(n20571), .Z(n20620) );
  XNOR U21126 ( .A(n20621), .B(n20620), .Z(n20622) );
  XNOR U21127 ( .A(n20623), .B(n20622), .Z(n20627) );
  NANDN U21128 ( .A(n20574), .B(n20573), .Z(n20578) );
  NAND U21129 ( .A(n20576), .B(n20575), .Z(n20577) );
  AND U21130 ( .A(n20578), .B(n20577), .Z(n20626) );
  XOR U21131 ( .A(n20627), .B(n20626), .Z(n20628) );
  NANDN U21132 ( .A(n20580), .B(n20579), .Z(n20584) );
  NANDN U21133 ( .A(n20582), .B(n20581), .Z(n20583) );
  NAND U21134 ( .A(n20584), .B(n20583), .Z(n20629) );
  XOR U21135 ( .A(n20628), .B(n20629), .Z(n20596) );
  OR U21136 ( .A(n20586), .B(n20585), .Z(n20590) );
  NANDN U21137 ( .A(n20588), .B(n20587), .Z(n20589) );
  NAND U21138 ( .A(n20590), .B(n20589), .Z(n20597) );
  XNOR U21139 ( .A(n20596), .B(n20597), .Z(n20598) );
  XNOR U21140 ( .A(n20599), .B(n20598), .Z(n20632) );
  XNOR U21141 ( .A(n20632), .B(sreg[1516]), .Z(n20634) );
  NAND U21142 ( .A(n20591), .B(sreg[1515]), .Z(n20595) );
  OR U21143 ( .A(n20593), .B(n20592), .Z(n20594) );
  AND U21144 ( .A(n20595), .B(n20594), .Z(n20633) );
  XOR U21145 ( .A(n20634), .B(n20633), .Z(c[1516]) );
  NANDN U21146 ( .A(n20597), .B(n20596), .Z(n20601) );
  NAND U21147 ( .A(n20599), .B(n20598), .Z(n20600) );
  NAND U21148 ( .A(n20601), .B(n20600), .Z(n20640) );
  NAND U21149 ( .A(b[0]), .B(a[501]), .Z(n20602) );
  XNOR U21150 ( .A(b[1]), .B(n20602), .Z(n20604) );
  NAND U21151 ( .A(n86), .B(a[500]), .Z(n20603) );
  AND U21152 ( .A(n20604), .B(n20603), .Z(n20657) );
  XOR U21153 ( .A(a[497]), .B(n42197), .Z(n20646) );
  NANDN U21154 ( .A(n20646), .B(n42173), .Z(n20607) );
  NANDN U21155 ( .A(n20605), .B(n42172), .Z(n20606) );
  NAND U21156 ( .A(n20607), .B(n20606), .Z(n20655) );
  NAND U21157 ( .A(b[7]), .B(a[493]), .Z(n20656) );
  XNOR U21158 ( .A(n20655), .B(n20656), .Z(n20658) );
  XOR U21159 ( .A(n20657), .B(n20658), .Z(n20664) );
  NANDN U21160 ( .A(n20608), .B(n42093), .Z(n20610) );
  XOR U21161 ( .A(n42134), .B(a[499]), .Z(n20649) );
  NANDN U21162 ( .A(n20649), .B(n42095), .Z(n20609) );
  NAND U21163 ( .A(n20610), .B(n20609), .Z(n20662) );
  NANDN U21164 ( .A(n20611), .B(n42231), .Z(n20613) );
  XOR U21165 ( .A(n203), .B(a[495]), .Z(n20652) );
  NANDN U21166 ( .A(n20652), .B(n42234), .Z(n20612) );
  AND U21167 ( .A(n20613), .B(n20612), .Z(n20661) );
  XNOR U21168 ( .A(n20662), .B(n20661), .Z(n20663) );
  XNOR U21169 ( .A(n20664), .B(n20663), .Z(n20668) );
  NANDN U21170 ( .A(n20615), .B(n20614), .Z(n20619) );
  NAND U21171 ( .A(n20617), .B(n20616), .Z(n20618) );
  AND U21172 ( .A(n20619), .B(n20618), .Z(n20667) );
  XOR U21173 ( .A(n20668), .B(n20667), .Z(n20669) );
  NANDN U21174 ( .A(n20621), .B(n20620), .Z(n20625) );
  NANDN U21175 ( .A(n20623), .B(n20622), .Z(n20624) );
  NAND U21176 ( .A(n20625), .B(n20624), .Z(n20670) );
  XOR U21177 ( .A(n20669), .B(n20670), .Z(n20637) );
  OR U21178 ( .A(n20627), .B(n20626), .Z(n20631) );
  NANDN U21179 ( .A(n20629), .B(n20628), .Z(n20630) );
  NAND U21180 ( .A(n20631), .B(n20630), .Z(n20638) );
  XNOR U21181 ( .A(n20637), .B(n20638), .Z(n20639) );
  XNOR U21182 ( .A(n20640), .B(n20639), .Z(n20673) );
  XNOR U21183 ( .A(n20673), .B(sreg[1517]), .Z(n20675) );
  NAND U21184 ( .A(n20632), .B(sreg[1516]), .Z(n20636) );
  OR U21185 ( .A(n20634), .B(n20633), .Z(n20635) );
  AND U21186 ( .A(n20636), .B(n20635), .Z(n20674) );
  XOR U21187 ( .A(n20675), .B(n20674), .Z(c[1517]) );
  NANDN U21188 ( .A(n20638), .B(n20637), .Z(n20642) );
  NAND U21189 ( .A(n20640), .B(n20639), .Z(n20641) );
  NAND U21190 ( .A(n20642), .B(n20641), .Z(n20681) );
  NAND U21191 ( .A(b[0]), .B(a[502]), .Z(n20643) );
  XNOR U21192 ( .A(b[1]), .B(n20643), .Z(n20645) );
  NAND U21193 ( .A(n86), .B(a[501]), .Z(n20644) );
  AND U21194 ( .A(n20645), .B(n20644), .Z(n20698) );
  XOR U21195 ( .A(a[498]), .B(n42197), .Z(n20687) );
  NANDN U21196 ( .A(n20687), .B(n42173), .Z(n20648) );
  NANDN U21197 ( .A(n20646), .B(n42172), .Z(n20647) );
  NAND U21198 ( .A(n20648), .B(n20647), .Z(n20696) );
  NAND U21199 ( .A(b[7]), .B(a[494]), .Z(n20697) );
  XNOR U21200 ( .A(n20696), .B(n20697), .Z(n20699) );
  XOR U21201 ( .A(n20698), .B(n20699), .Z(n20705) );
  NANDN U21202 ( .A(n20649), .B(n42093), .Z(n20651) );
  XOR U21203 ( .A(n42134), .B(a[500]), .Z(n20690) );
  NANDN U21204 ( .A(n20690), .B(n42095), .Z(n20650) );
  NAND U21205 ( .A(n20651), .B(n20650), .Z(n20703) );
  NANDN U21206 ( .A(n20652), .B(n42231), .Z(n20654) );
  XOR U21207 ( .A(n203), .B(a[496]), .Z(n20693) );
  NANDN U21208 ( .A(n20693), .B(n42234), .Z(n20653) );
  AND U21209 ( .A(n20654), .B(n20653), .Z(n20702) );
  XNOR U21210 ( .A(n20703), .B(n20702), .Z(n20704) );
  XNOR U21211 ( .A(n20705), .B(n20704), .Z(n20709) );
  NANDN U21212 ( .A(n20656), .B(n20655), .Z(n20660) );
  NAND U21213 ( .A(n20658), .B(n20657), .Z(n20659) );
  AND U21214 ( .A(n20660), .B(n20659), .Z(n20708) );
  XOR U21215 ( .A(n20709), .B(n20708), .Z(n20710) );
  NANDN U21216 ( .A(n20662), .B(n20661), .Z(n20666) );
  NANDN U21217 ( .A(n20664), .B(n20663), .Z(n20665) );
  NAND U21218 ( .A(n20666), .B(n20665), .Z(n20711) );
  XOR U21219 ( .A(n20710), .B(n20711), .Z(n20678) );
  OR U21220 ( .A(n20668), .B(n20667), .Z(n20672) );
  NANDN U21221 ( .A(n20670), .B(n20669), .Z(n20671) );
  NAND U21222 ( .A(n20672), .B(n20671), .Z(n20679) );
  XNOR U21223 ( .A(n20678), .B(n20679), .Z(n20680) );
  XNOR U21224 ( .A(n20681), .B(n20680), .Z(n20714) );
  XNOR U21225 ( .A(n20714), .B(sreg[1518]), .Z(n20716) );
  NAND U21226 ( .A(n20673), .B(sreg[1517]), .Z(n20677) );
  OR U21227 ( .A(n20675), .B(n20674), .Z(n20676) );
  AND U21228 ( .A(n20677), .B(n20676), .Z(n20715) );
  XOR U21229 ( .A(n20716), .B(n20715), .Z(c[1518]) );
  NANDN U21230 ( .A(n20679), .B(n20678), .Z(n20683) );
  NAND U21231 ( .A(n20681), .B(n20680), .Z(n20682) );
  NAND U21232 ( .A(n20683), .B(n20682), .Z(n20722) );
  NAND U21233 ( .A(b[0]), .B(a[503]), .Z(n20684) );
  XNOR U21234 ( .A(b[1]), .B(n20684), .Z(n20686) );
  NAND U21235 ( .A(n86), .B(a[502]), .Z(n20685) );
  AND U21236 ( .A(n20686), .B(n20685), .Z(n20739) );
  XOR U21237 ( .A(a[499]), .B(n42197), .Z(n20728) );
  NANDN U21238 ( .A(n20728), .B(n42173), .Z(n20689) );
  NANDN U21239 ( .A(n20687), .B(n42172), .Z(n20688) );
  NAND U21240 ( .A(n20689), .B(n20688), .Z(n20737) );
  NAND U21241 ( .A(b[7]), .B(a[495]), .Z(n20738) );
  XNOR U21242 ( .A(n20737), .B(n20738), .Z(n20740) );
  XOR U21243 ( .A(n20739), .B(n20740), .Z(n20746) );
  NANDN U21244 ( .A(n20690), .B(n42093), .Z(n20692) );
  XOR U21245 ( .A(n42134), .B(a[501]), .Z(n20731) );
  NANDN U21246 ( .A(n20731), .B(n42095), .Z(n20691) );
  NAND U21247 ( .A(n20692), .B(n20691), .Z(n20744) );
  NANDN U21248 ( .A(n20693), .B(n42231), .Z(n20695) );
  XOR U21249 ( .A(n203), .B(a[497]), .Z(n20734) );
  NANDN U21250 ( .A(n20734), .B(n42234), .Z(n20694) );
  AND U21251 ( .A(n20695), .B(n20694), .Z(n20743) );
  XNOR U21252 ( .A(n20744), .B(n20743), .Z(n20745) );
  XNOR U21253 ( .A(n20746), .B(n20745), .Z(n20750) );
  NANDN U21254 ( .A(n20697), .B(n20696), .Z(n20701) );
  NAND U21255 ( .A(n20699), .B(n20698), .Z(n20700) );
  AND U21256 ( .A(n20701), .B(n20700), .Z(n20749) );
  XOR U21257 ( .A(n20750), .B(n20749), .Z(n20751) );
  NANDN U21258 ( .A(n20703), .B(n20702), .Z(n20707) );
  NANDN U21259 ( .A(n20705), .B(n20704), .Z(n20706) );
  NAND U21260 ( .A(n20707), .B(n20706), .Z(n20752) );
  XOR U21261 ( .A(n20751), .B(n20752), .Z(n20719) );
  OR U21262 ( .A(n20709), .B(n20708), .Z(n20713) );
  NANDN U21263 ( .A(n20711), .B(n20710), .Z(n20712) );
  NAND U21264 ( .A(n20713), .B(n20712), .Z(n20720) );
  XNOR U21265 ( .A(n20719), .B(n20720), .Z(n20721) );
  XNOR U21266 ( .A(n20722), .B(n20721), .Z(n20755) );
  XNOR U21267 ( .A(n20755), .B(sreg[1519]), .Z(n20757) );
  NAND U21268 ( .A(n20714), .B(sreg[1518]), .Z(n20718) );
  OR U21269 ( .A(n20716), .B(n20715), .Z(n20717) );
  AND U21270 ( .A(n20718), .B(n20717), .Z(n20756) );
  XOR U21271 ( .A(n20757), .B(n20756), .Z(c[1519]) );
  NANDN U21272 ( .A(n20720), .B(n20719), .Z(n20724) );
  NAND U21273 ( .A(n20722), .B(n20721), .Z(n20723) );
  NAND U21274 ( .A(n20724), .B(n20723), .Z(n20763) );
  NAND U21275 ( .A(b[0]), .B(a[504]), .Z(n20725) );
  XNOR U21276 ( .A(b[1]), .B(n20725), .Z(n20727) );
  NAND U21277 ( .A(n87), .B(a[503]), .Z(n20726) );
  AND U21278 ( .A(n20727), .B(n20726), .Z(n20780) );
  XOR U21279 ( .A(a[500]), .B(n42197), .Z(n20769) );
  NANDN U21280 ( .A(n20769), .B(n42173), .Z(n20730) );
  NANDN U21281 ( .A(n20728), .B(n42172), .Z(n20729) );
  NAND U21282 ( .A(n20730), .B(n20729), .Z(n20778) );
  NAND U21283 ( .A(b[7]), .B(a[496]), .Z(n20779) );
  XNOR U21284 ( .A(n20778), .B(n20779), .Z(n20781) );
  XOR U21285 ( .A(n20780), .B(n20781), .Z(n20787) );
  NANDN U21286 ( .A(n20731), .B(n42093), .Z(n20733) );
  XOR U21287 ( .A(n42134), .B(a[502]), .Z(n20772) );
  NANDN U21288 ( .A(n20772), .B(n42095), .Z(n20732) );
  NAND U21289 ( .A(n20733), .B(n20732), .Z(n20785) );
  NANDN U21290 ( .A(n20734), .B(n42231), .Z(n20736) );
  XOR U21291 ( .A(n203), .B(a[498]), .Z(n20775) );
  NANDN U21292 ( .A(n20775), .B(n42234), .Z(n20735) );
  AND U21293 ( .A(n20736), .B(n20735), .Z(n20784) );
  XNOR U21294 ( .A(n20785), .B(n20784), .Z(n20786) );
  XNOR U21295 ( .A(n20787), .B(n20786), .Z(n20791) );
  NANDN U21296 ( .A(n20738), .B(n20737), .Z(n20742) );
  NAND U21297 ( .A(n20740), .B(n20739), .Z(n20741) );
  AND U21298 ( .A(n20742), .B(n20741), .Z(n20790) );
  XOR U21299 ( .A(n20791), .B(n20790), .Z(n20792) );
  NANDN U21300 ( .A(n20744), .B(n20743), .Z(n20748) );
  NANDN U21301 ( .A(n20746), .B(n20745), .Z(n20747) );
  NAND U21302 ( .A(n20748), .B(n20747), .Z(n20793) );
  XOR U21303 ( .A(n20792), .B(n20793), .Z(n20760) );
  OR U21304 ( .A(n20750), .B(n20749), .Z(n20754) );
  NANDN U21305 ( .A(n20752), .B(n20751), .Z(n20753) );
  NAND U21306 ( .A(n20754), .B(n20753), .Z(n20761) );
  XNOR U21307 ( .A(n20760), .B(n20761), .Z(n20762) );
  XNOR U21308 ( .A(n20763), .B(n20762), .Z(n20796) );
  XNOR U21309 ( .A(n20796), .B(sreg[1520]), .Z(n20798) );
  NAND U21310 ( .A(n20755), .B(sreg[1519]), .Z(n20759) );
  OR U21311 ( .A(n20757), .B(n20756), .Z(n20758) );
  AND U21312 ( .A(n20759), .B(n20758), .Z(n20797) );
  XOR U21313 ( .A(n20798), .B(n20797), .Z(c[1520]) );
  NANDN U21314 ( .A(n20761), .B(n20760), .Z(n20765) );
  NAND U21315 ( .A(n20763), .B(n20762), .Z(n20764) );
  NAND U21316 ( .A(n20765), .B(n20764), .Z(n20804) );
  NAND U21317 ( .A(b[0]), .B(a[505]), .Z(n20766) );
  XNOR U21318 ( .A(b[1]), .B(n20766), .Z(n20768) );
  NAND U21319 ( .A(n87), .B(a[504]), .Z(n20767) );
  AND U21320 ( .A(n20768), .B(n20767), .Z(n20821) );
  XOR U21321 ( .A(a[501]), .B(n42197), .Z(n20810) );
  NANDN U21322 ( .A(n20810), .B(n42173), .Z(n20771) );
  NANDN U21323 ( .A(n20769), .B(n42172), .Z(n20770) );
  NAND U21324 ( .A(n20771), .B(n20770), .Z(n20819) );
  NAND U21325 ( .A(b[7]), .B(a[497]), .Z(n20820) );
  XNOR U21326 ( .A(n20819), .B(n20820), .Z(n20822) );
  XOR U21327 ( .A(n20821), .B(n20822), .Z(n20828) );
  NANDN U21328 ( .A(n20772), .B(n42093), .Z(n20774) );
  XOR U21329 ( .A(n42134), .B(a[503]), .Z(n20813) );
  NANDN U21330 ( .A(n20813), .B(n42095), .Z(n20773) );
  NAND U21331 ( .A(n20774), .B(n20773), .Z(n20826) );
  NANDN U21332 ( .A(n20775), .B(n42231), .Z(n20777) );
  XOR U21333 ( .A(n203), .B(a[499]), .Z(n20816) );
  NANDN U21334 ( .A(n20816), .B(n42234), .Z(n20776) );
  AND U21335 ( .A(n20777), .B(n20776), .Z(n20825) );
  XNOR U21336 ( .A(n20826), .B(n20825), .Z(n20827) );
  XNOR U21337 ( .A(n20828), .B(n20827), .Z(n20832) );
  NANDN U21338 ( .A(n20779), .B(n20778), .Z(n20783) );
  NAND U21339 ( .A(n20781), .B(n20780), .Z(n20782) );
  AND U21340 ( .A(n20783), .B(n20782), .Z(n20831) );
  XOR U21341 ( .A(n20832), .B(n20831), .Z(n20833) );
  NANDN U21342 ( .A(n20785), .B(n20784), .Z(n20789) );
  NANDN U21343 ( .A(n20787), .B(n20786), .Z(n20788) );
  NAND U21344 ( .A(n20789), .B(n20788), .Z(n20834) );
  XOR U21345 ( .A(n20833), .B(n20834), .Z(n20801) );
  OR U21346 ( .A(n20791), .B(n20790), .Z(n20795) );
  NANDN U21347 ( .A(n20793), .B(n20792), .Z(n20794) );
  NAND U21348 ( .A(n20795), .B(n20794), .Z(n20802) );
  XNOR U21349 ( .A(n20801), .B(n20802), .Z(n20803) );
  XNOR U21350 ( .A(n20804), .B(n20803), .Z(n20837) );
  XNOR U21351 ( .A(n20837), .B(sreg[1521]), .Z(n20839) );
  NAND U21352 ( .A(n20796), .B(sreg[1520]), .Z(n20800) );
  OR U21353 ( .A(n20798), .B(n20797), .Z(n20799) );
  AND U21354 ( .A(n20800), .B(n20799), .Z(n20838) );
  XOR U21355 ( .A(n20839), .B(n20838), .Z(c[1521]) );
  NANDN U21356 ( .A(n20802), .B(n20801), .Z(n20806) );
  NAND U21357 ( .A(n20804), .B(n20803), .Z(n20805) );
  NAND U21358 ( .A(n20806), .B(n20805), .Z(n20845) );
  NAND U21359 ( .A(b[0]), .B(a[506]), .Z(n20807) );
  XNOR U21360 ( .A(b[1]), .B(n20807), .Z(n20809) );
  NAND U21361 ( .A(n87), .B(a[505]), .Z(n20808) );
  AND U21362 ( .A(n20809), .B(n20808), .Z(n20862) );
  XOR U21363 ( .A(a[502]), .B(n42197), .Z(n20851) );
  NANDN U21364 ( .A(n20851), .B(n42173), .Z(n20812) );
  NANDN U21365 ( .A(n20810), .B(n42172), .Z(n20811) );
  NAND U21366 ( .A(n20812), .B(n20811), .Z(n20860) );
  NAND U21367 ( .A(b[7]), .B(a[498]), .Z(n20861) );
  XNOR U21368 ( .A(n20860), .B(n20861), .Z(n20863) );
  XOR U21369 ( .A(n20862), .B(n20863), .Z(n20869) );
  NANDN U21370 ( .A(n20813), .B(n42093), .Z(n20815) );
  XOR U21371 ( .A(n42134), .B(a[504]), .Z(n20854) );
  NANDN U21372 ( .A(n20854), .B(n42095), .Z(n20814) );
  NAND U21373 ( .A(n20815), .B(n20814), .Z(n20867) );
  NANDN U21374 ( .A(n20816), .B(n42231), .Z(n20818) );
  XOR U21375 ( .A(n203), .B(a[500]), .Z(n20857) );
  NANDN U21376 ( .A(n20857), .B(n42234), .Z(n20817) );
  AND U21377 ( .A(n20818), .B(n20817), .Z(n20866) );
  XNOR U21378 ( .A(n20867), .B(n20866), .Z(n20868) );
  XNOR U21379 ( .A(n20869), .B(n20868), .Z(n20873) );
  NANDN U21380 ( .A(n20820), .B(n20819), .Z(n20824) );
  NAND U21381 ( .A(n20822), .B(n20821), .Z(n20823) );
  AND U21382 ( .A(n20824), .B(n20823), .Z(n20872) );
  XOR U21383 ( .A(n20873), .B(n20872), .Z(n20874) );
  NANDN U21384 ( .A(n20826), .B(n20825), .Z(n20830) );
  NANDN U21385 ( .A(n20828), .B(n20827), .Z(n20829) );
  NAND U21386 ( .A(n20830), .B(n20829), .Z(n20875) );
  XOR U21387 ( .A(n20874), .B(n20875), .Z(n20842) );
  OR U21388 ( .A(n20832), .B(n20831), .Z(n20836) );
  NANDN U21389 ( .A(n20834), .B(n20833), .Z(n20835) );
  NAND U21390 ( .A(n20836), .B(n20835), .Z(n20843) );
  XNOR U21391 ( .A(n20842), .B(n20843), .Z(n20844) );
  XNOR U21392 ( .A(n20845), .B(n20844), .Z(n20878) );
  XNOR U21393 ( .A(n20878), .B(sreg[1522]), .Z(n20880) );
  NAND U21394 ( .A(n20837), .B(sreg[1521]), .Z(n20841) );
  OR U21395 ( .A(n20839), .B(n20838), .Z(n20840) );
  AND U21396 ( .A(n20841), .B(n20840), .Z(n20879) );
  XOR U21397 ( .A(n20880), .B(n20879), .Z(c[1522]) );
  NANDN U21398 ( .A(n20843), .B(n20842), .Z(n20847) );
  NAND U21399 ( .A(n20845), .B(n20844), .Z(n20846) );
  NAND U21400 ( .A(n20847), .B(n20846), .Z(n20886) );
  NAND U21401 ( .A(b[0]), .B(a[507]), .Z(n20848) );
  XNOR U21402 ( .A(b[1]), .B(n20848), .Z(n20850) );
  NAND U21403 ( .A(n87), .B(a[506]), .Z(n20849) );
  AND U21404 ( .A(n20850), .B(n20849), .Z(n20903) );
  XOR U21405 ( .A(a[503]), .B(n42197), .Z(n20892) );
  NANDN U21406 ( .A(n20892), .B(n42173), .Z(n20853) );
  NANDN U21407 ( .A(n20851), .B(n42172), .Z(n20852) );
  NAND U21408 ( .A(n20853), .B(n20852), .Z(n20901) );
  NAND U21409 ( .A(b[7]), .B(a[499]), .Z(n20902) );
  XNOR U21410 ( .A(n20901), .B(n20902), .Z(n20904) );
  XOR U21411 ( .A(n20903), .B(n20904), .Z(n20910) );
  NANDN U21412 ( .A(n20854), .B(n42093), .Z(n20856) );
  XOR U21413 ( .A(n42134), .B(a[505]), .Z(n20895) );
  NANDN U21414 ( .A(n20895), .B(n42095), .Z(n20855) );
  NAND U21415 ( .A(n20856), .B(n20855), .Z(n20908) );
  NANDN U21416 ( .A(n20857), .B(n42231), .Z(n20859) );
  XOR U21417 ( .A(n203), .B(a[501]), .Z(n20898) );
  NANDN U21418 ( .A(n20898), .B(n42234), .Z(n20858) );
  AND U21419 ( .A(n20859), .B(n20858), .Z(n20907) );
  XNOR U21420 ( .A(n20908), .B(n20907), .Z(n20909) );
  XNOR U21421 ( .A(n20910), .B(n20909), .Z(n20914) );
  NANDN U21422 ( .A(n20861), .B(n20860), .Z(n20865) );
  NAND U21423 ( .A(n20863), .B(n20862), .Z(n20864) );
  AND U21424 ( .A(n20865), .B(n20864), .Z(n20913) );
  XOR U21425 ( .A(n20914), .B(n20913), .Z(n20915) );
  NANDN U21426 ( .A(n20867), .B(n20866), .Z(n20871) );
  NANDN U21427 ( .A(n20869), .B(n20868), .Z(n20870) );
  NAND U21428 ( .A(n20871), .B(n20870), .Z(n20916) );
  XOR U21429 ( .A(n20915), .B(n20916), .Z(n20883) );
  OR U21430 ( .A(n20873), .B(n20872), .Z(n20877) );
  NANDN U21431 ( .A(n20875), .B(n20874), .Z(n20876) );
  NAND U21432 ( .A(n20877), .B(n20876), .Z(n20884) );
  XNOR U21433 ( .A(n20883), .B(n20884), .Z(n20885) );
  XNOR U21434 ( .A(n20886), .B(n20885), .Z(n20919) );
  XNOR U21435 ( .A(n20919), .B(sreg[1523]), .Z(n20921) );
  NAND U21436 ( .A(n20878), .B(sreg[1522]), .Z(n20882) );
  OR U21437 ( .A(n20880), .B(n20879), .Z(n20881) );
  AND U21438 ( .A(n20882), .B(n20881), .Z(n20920) );
  XOR U21439 ( .A(n20921), .B(n20920), .Z(c[1523]) );
  NANDN U21440 ( .A(n20884), .B(n20883), .Z(n20888) );
  NAND U21441 ( .A(n20886), .B(n20885), .Z(n20887) );
  NAND U21442 ( .A(n20888), .B(n20887), .Z(n20927) );
  NAND U21443 ( .A(b[0]), .B(a[508]), .Z(n20889) );
  XNOR U21444 ( .A(b[1]), .B(n20889), .Z(n20891) );
  NAND U21445 ( .A(n87), .B(a[507]), .Z(n20890) );
  AND U21446 ( .A(n20891), .B(n20890), .Z(n20944) );
  XOR U21447 ( .A(a[504]), .B(n42197), .Z(n20933) );
  NANDN U21448 ( .A(n20933), .B(n42173), .Z(n20894) );
  NANDN U21449 ( .A(n20892), .B(n42172), .Z(n20893) );
  NAND U21450 ( .A(n20894), .B(n20893), .Z(n20942) );
  NAND U21451 ( .A(b[7]), .B(a[500]), .Z(n20943) );
  XNOR U21452 ( .A(n20942), .B(n20943), .Z(n20945) );
  XOR U21453 ( .A(n20944), .B(n20945), .Z(n20951) );
  NANDN U21454 ( .A(n20895), .B(n42093), .Z(n20897) );
  XOR U21455 ( .A(n42134), .B(a[506]), .Z(n20936) );
  NANDN U21456 ( .A(n20936), .B(n42095), .Z(n20896) );
  NAND U21457 ( .A(n20897), .B(n20896), .Z(n20949) );
  NANDN U21458 ( .A(n20898), .B(n42231), .Z(n20900) );
  XOR U21459 ( .A(n203), .B(a[502]), .Z(n20939) );
  NANDN U21460 ( .A(n20939), .B(n42234), .Z(n20899) );
  AND U21461 ( .A(n20900), .B(n20899), .Z(n20948) );
  XNOR U21462 ( .A(n20949), .B(n20948), .Z(n20950) );
  XNOR U21463 ( .A(n20951), .B(n20950), .Z(n20955) );
  NANDN U21464 ( .A(n20902), .B(n20901), .Z(n20906) );
  NAND U21465 ( .A(n20904), .B(n20903), .Z(n20905) );
  AND U21466 ( .A(n20906), .B(n20905), .Z(n20954) );
  XOR U21467 ( .A(n20955), .B(n20954), .Z(n20956) );
  NANDN U21468 ( .A(n20908), .B(n20907), .Z(n20912) );
  NANDN U21469 ( .A(n20910), .B(n20909), .Z(n20911) );
  NAND U21470 ( .A(n20912), .B(n20911), .Z(n20957) );
  XOR U21471 ( .A(n20956), .B(n20957), .Z(n20924) );
  OR U21472 ( .A(n20914), .B(n20913), .Z(n20918) );
  NANDN U21473 ( .A(n20916), .B(n20915), .Z(n20917) );
  NAND U21474 ( .A(n20918), .B(n20917), .Z(n20925) );
  XNOR U21475 ( .A(n20924), .B(n20925), .Z(n20926) );
  XNOR U21476 ( .A(n20927), .B(n20926), .Z(n20960) );
  XNOR U21477 ( .A(n20960), .B(sreg[1524]), .Z(n20962) );
  NAND U21478 ( .A(n20919), .B(sreg[1523]), .Z(n20923) );
  OR U21479 ( .A(n20921), .B(n20920), .Z(n20922) );
  AND U21480 ( .A(n20923), .B(n20922), .Z(n20961) );
  XOR U21481 ( .A(n20962), .B(n20961), .Z(c[1524]) );
  NANDN U21482 ( .A(n20925), .B(n20924), .Z(n20929) );
  NAND U21483 ( .A(n20927), .B(n20926), .Z(n20928) );
  NAND U21484 ( .A(n20929), .B(n20928), .Z(n20968) );
  NAND U21485 ( .A(b[0]), .B(a[509]), .Z(n20930) );
  XNOR U21486 ( .A(b[1]), .B(n20930), .Z(n20932) );
  NAND U21487 ( .A(n87), .B(a[508]), .Z(n20931) );
  AND U21488 ( .A(n20932), .B(n20931), .Z(n20985) );
  XOR U21489 ( .A(a[505]), .B(n42197), .Z(n20974) );
  NANDN U21490 ( .A(n20974), .B(n42173), .Z(n20935) );
  NANDN U21491 ( .A(n20933), .B(n42172), .Z(n20934) );
  NAND U21492 ( .A(n20935), .B(n20934), .Z(n20983) );
  NAND U21493 ( .A(b[7]), .B(a[501]), .Z(n20984) );
  XNOR U21494 ( .A(n20983), .B(n20984), .Z(n20986) );
  XOR U21495 ( .A(n20985), .B(n20986), .Z(n20992) );
  NANDN U21496 ( .A(n20936), .B(n42093), .Z(n20938) );
  XOR U21497 ( .A(n42134), .B(a[507]), .Z(n20977) );
  NANDN U21498 ( .A(n20977), .B(n42095), .Z(n20937) );
  NAND U21499 ( .A(n20938), .B(n20937), .Z(n20990) );
  NANDN U21500 ( .A(n20939), .B(n42231), .Z(n20941) );
  XOR U21501 ( .A(n204), .B(a[503]), .Z(n20980) );
  NANDN U21502 ( .A(n20980), .B(n42234), .Z(n20940) );
  AND U21503 ( .A(n20941), .B(n20940), .Z(n20989) );
  XNOR U21504 ( .A(n20990), .B(n20989), .Z(n20991) );
  XNOR U21505 ( .A(n20992), .B(n20991), .Z(n20996) );
  NANDN U21506 ( .A(n20943), .B(n20942), .Z(n20947) );
  NAND U21507 ( .A(n20945), .B(n20944), .Z(n20946) );
  AND U21508 ( .A(n20947), .B(n20946), .Z(n20995) );
  XOR U21509 ( .A(n20996), .B(n20995), .Z(n20997) );
  NANDN U21510 ( .A(n20949), .B(n20948), .Z(n20953) );
  NANDN U21511 ( .A(n20951), .B(n20950), .Z(n20952) );
  NAND U21512 ( .A(n20953), .B(n20952), .Z(n20998) );
  XOR U21513 ( .A(n20997), .B(n20998), .Z(n20965) );
  OR U21514 ( .A(n20955), .B(n20954), .Z(n20959) );
  NANDN U21515 ( .A(n20957), .B(n20956), .Z(n20958) );
  NAND U21516 ( .A(n20959), .B(n20958), .Z(n20966) );
  XNOR U21517 ( .A(n20965), .B(n20966), .Z(n20967) );
  XNOR U21518 ( .A(n20968), .B(n20967), .Z(n21001) );
  XNOR U21519 ( .A(n21001), .B(sreg[1525]), .Z(n21003) );
  NAND U21520 ( .A(n20960), .B(sreg[1524]), .Z(n20964) );
  OR U21521 ( .A(n20962), .B(n20961), .Z(n20963) );
  AND U21522 ( .A(n20964), .B(n20963), .Z(n21002) );
  XOR U21523 ( .A(n21003), .B(n21002), .Z(c[1525]) );
  NANDN U21524 ( .A(n20966), .B(n20965), .Z(n20970) );
  NAND U21525 ( .A(n20968), .B(n20967), .Z(n20969) );
  NAND U21526 ( .A(n20970), .B(n20969), .Z(n21009) );
  NAND U21527 ( .A(b[0]), .B(a[510]), .Z(n20971) );
  XNOR U21528 ( .A(b[1]), .B(n20971), .Z(n20973) );
  NAND U21529 ( .A(n87), .B(a[509]), .Z(n20972) );
  AND U21530 ( .A(n20973), .B(n20972), .Z(n21026) );
  XOR U21531 ( .A(a[506]), .B(n42197), .Z(n21015) );
  NANDN U21532 ( .A(n21015), .B(n42173), .Z(n20976) );
  NANDN U21533 ( .A(n20974), .B(n42172), .Z(n20975) );
  NAND U21534 ( .A(n20976), .B(n20975), .Z(n21024) );
  NAND U21535 ( .A(b[7]), .B(a[502]), .Z(n21025) );
  XNOR U21536 ( .A(n21024), .B(n21025), .Z(n21027) );
  XOR U21537 ( .A(n21026), .B(n21027), .Z(n21033) );
  NANDN U21538 ( .A(n20977), .B(n42093), .Z(n20979) );
  XOR U21539 ( .A(n42134), .B(a[508]), .Z(n21018) );
  NANDN U21540 ( .A(n21018), .B(n42095), .Z(n20978) );
  NAND U21541 ( .A(n20979), .B(n20978), .Z(n21031) );
  NANDN U21542 ( .A(n20980), .B(n42231), .Z(n20982) );
  XOR U21543 ( .A(n204), .B(a[504]), .Z(n21021) );
  NANDN U21544 ( .A(n21021), .B(n42234), .Z(n20981) );
  AND U21545 ( .A(n20982), .B(n20981), .Z(n21030) );
  XNOR U21546 ( .A(n21031), .B(n21030), .Z(n21032) );
  XNOR U21547 ( .A(n21033), .B(n21032), .Z(n21037) );
  NANDN U21548 ( .A(n20984), .B(n20983), .Z(n20988) );
  NAND U21549 ( .A(n20986), .B(n20985), .Z(n20987) );
  AND U21550 ( .A(n20988), .B(n20987), .Z(n21036) );
  XOR U21551 ( .A(n21037), .B(n21036), .Z(n21038) );
  NANDN U21552 ( .A(n20990), .B(n20989), .Z(n20994) );
  NANDN U21553 ( .A(n20992), .B(n20991), .Z(n20993) );
  NAND U21554 ( .A(n20994), .B(n20993), .Z(n21039) );
  XOR U21555 ( .A(n21038), .B(n21039), .Z(n21006) );
  OR U21556 ( .A(n20996), .B(n20995), .Z(n21000) );
  NANDN U21557 ( .A(n20998), .B(n20997), .Z(n20999) );
  NAND U21558 ( .A(n21000), .B(n20999), .Z(n21007) );
  XNOR U21559 ( .A(n21006), .B(n21007), .Z(n21008) );
  XNOR U21560 ( .A(n21009), .B(n21008), .Z(n21042) );
  XNOR U21561 ( .A(n21042), .B(sreg[1526]), .Z(n21044) );
  NAND U21562 ( .A(n21001), .B(sreg[1525]), .Z(n21005) );
  OR U21563 ( .A(n21003), .B(n21002), .Z(n21004) );
  AND U21564 ( .A(n21005), .B(n21004), .Z(n21043) );
  XOR U21565 ( .A(n21044), .B(n21043), .Z(c[1526]) );
  NANDN U21566 ( .A(n21007), .B(n21006), .Z(n21011) );
  NAND U21567 ( .A(n21009), .B(n21008), .Z(n21010) );
  NAND U21568 ( .A(n21011), .B(n21010), .Z(n21050) );
  NAND U21569 ( .A(b[0]), .B(a[511]), .Z(n21012) );
  XNOR U21570 ( .A(b[1]), .B(n21012), .Z(n21014) );
  NAND U21571 ( .A(n88), .B(a[510]), .Z(n21013) );
  AND U21572 ( .A(n21014), .B(n21013), .Z(n21067) );
  XOR U21573 ( .A(a[507]), .B(n42197), .Z(n21056) );
  NANDN U21574 ( .A(n21056), .B(n42173), .Z(n21017) );
  NANDN U21575 ( .A(n21015), .B(n42172), .Z(n21016) );
  NAND U21576 ( .A(n21017), .B(n21016), .Z(n21065) );
  NAND U21577 ( .A(b[7]), .B(a[503]), .Z(n21066) );
  XNOR U21578 ( .A(n21065), .B(n21066), .Z(n21068) );
  XOR U21579 ( .A(n21067), .B(n21068), .Z(n21074) );
  NANDN U21580 ( .A(n21018), .B(n42093), .Z(n21020) );
  XOR U21581 ( .A(n42134), .B(a[509]), .Z(n21059) );
  NANDN U21582 ( .A(n21059), .B(n42095), .Z(n21019) );
  NAND U21583 ( .A(n21020), .B(n21019), .Z(n21072) );
  NANDN U21584 ( .A(n21021), .B(n42231), .Z(n21023) );
  XOR U21585 ( .A(n204), .B(a[505]), .Z(n21062) );
  NANDN U21586 ( .A(n21062), .B(n42234), .Z(n21022) );
  AND U21587 ( .A(n21023), .B(n21022), .Z(n21071) );
  XNOR U21588 ( .A(n21072), .B(n21071), .Z(n21073) );
  XNOR U21589 ( .A(n21074), .B(n21073), .Z(n21078) );
  NANDN U21590 ( .A(n21025), .B(n21024), .Z(n21029) );
  NAND U21591 ( .A(n21027), .B(n21026), .Z(n21028) );
  AND U21592 ( .A(n21029), .B(n21028), .Z(n21077) );
  XOR U21593 ( .A(n21078), .B(n21077), .Z(n21079) );
  NANDN U21594 ( .A(n21031), .B(n21030), .Z(n21035) );
  NANDN U21595 ( .A(n21033), .B(n21032), .Z(n21034) );
  NAND U21596 ( .A(n21035), .B(n21034), .Z(n21080) );
  XOR U21597 ( .A(n21079), .B(n21080), .Z(n21047) );
  OR U21598 ( .A(n21037), .B(n21036), .Z(n21041) );
  NANDN U21599 ( .A(n21039), .B(n21038), .Z(n21040) );
  NAND U21600 ( .A(n21041), .B(n21040), .Z(n21048) );
  XNOR U21601 ( .A(n21047), .B(n21048), .Z(n21049) );
  XNOR U21602 ( .A(n21050), .B(n21049), .Z(n21083) );
  XNOR U21603 ( .A(n21083), .B(sreg[1527]), .Z(n21085) );
  NAND U21604 ( .A(n21042), .B(sreg[1526]), .Z(n21046) );
  OR U21605 ( .A(n21044), .B(n21043), .Z(n21045) );
  AND U21606 ( .A(n21046), .B(n21045), .Z(n21084) );
  XOR U21607 ( .A(n21085), .B(n21084), .Z(c[1527]) );
  NANDN U21608 ( .A(n21048), .B(n21047), .Z(n21052) );
  NAND U21609 ( .A(n21050), .B(n21049), .Z(n21051) );
  NAND U21610 ( .A(n21052), .B(n21051), .Z(n21091) );
  NAND U21611 ( .A(b[0]), .B(a[512]), .Z(n21053) );
  XNOR U21612 ( .A(b[1]), .B(n21053), .Z(n21055) );
  NAND U21613 ( .A(n88), .B(a[511]), .Z(n21054) );
  AND U21614 ( .A(n21055), .B(n21054), .Z(n21108) );
  XOR U21615 ( .A(a[508]), .B(n42197), .Z(n21097) );
  NANDN U21616 ( .A(n21097), .B(n42173), .Z(n21058) );
  NANDN U21617 ( .A(n21056), .B(n42172), .Z(n21057) );
  NAND U21618 ( .A(n21058), .B(n21057), .Z(n21106) );
  NAND U21619 ( .A(b[7]), .B(a[504]), .Z(n21107) );
  XNOR U21620 ( .A(n21106), .B(n21107), .Z(n21109) );
  XOR U21621 ( .A(n21108), .B(n21109), .Z(n21115) );
  NANDN U21622 ( .A(n21059), .B(n42093), .Z(n21061) );
  XOR U21623 ( .A(n42134), .B(a[510]), .Z(n21100) );
  NANDN U21624 ( .A(n21100), .B(n42095), .Z(n21060) );
  NAND U21625 ( .A(n21061), .B(n21060), .Z(n21113) );
  NANDN U21626 ( .A(n21062), .B(n42231), .Z(n21064) );
  XOR U21627 ( .A(n204), .B(a[506]), .Z(n21103) );
  NANDN U21628 ( .A(n21103), .B(n42234), .Z(n21063) );
  AND U21629 ( .A(n21064), .B(n21063), .Z(n21112) );
  XNOR U21630 ( .A(n21113), .B(n21112), .Z(n21114) );
  XNOR U21631 ( .A(n21115), .B(n21114), .Z(n21119) );
  NANDN U21632 ( .A(n21066), .B(n21065), .Z(n21070) );
  NAND U21633 ( .A(n21068), .B(n21067), .Z(n21069) );
  AND U21634 ( .A(n21070), .B(n21069), .Z(n21118) );
  XOR U21635 ( .A(n21119), .B(n21118), .Z(n21120) );
  NANDN U21636 ( .A(n21072), .B(n21071), .Z(n21076) );
  NANDN U21637 ( .A(n21074), .B(n21073), .Z(n21075) );
  NAND U21638 ( .A(n21076), .B(n21075), .Z(n21121) );
  XOR U21639 ( .A(n21120), .B(n21121), .Z(n21088) );
  OR U21640 ( .A(n21078), .B(n21077), .Z(n21082) );
  NANDN U21641 ( .A(n21080), .B(n21079), .Z(n21081) );
  NAND U21642 ( .A(n21082), .B(n21081), .Z(n21089) );
  XNOR U21643 ( .A(n21088), .B(n21089), .Z(n21090) );
  XNOR U21644 ( .A(n21091), .B(n21090), .Z(n21124) );
  XNOR U21645 ( .A(n21124), .B(sreg[1528]), .Z(n21126) );
  NAND U21646 ( .A(n21083), .B(sreg[1527]), .Z(n21087) );
  OR U21647 ( .A(n21085), .B(n21084), .Z(n21086) );
  AND U21648 ( .A(n21087), .B(n21086), .Z(n21125) );
  XOR U21649 ( .A(n21126), .B(n21125), .Z(c[1528]) );
  NANDN U21650 ( .A(n21089), .B(n21088), .Z(n21093) );
  NAND U21651 ( .A(n21091), .B(n21090), .Z(n21092) );
  NAND U21652 ( .A(n21093), .B(n21092), .Z(n21132) );
  NAND U21653 ( .A(b[0]), .B(a[513]), .Z(n21094) );
  XNOR U21654 ( .A(b[1]), .B(n21094), .Z(n21096) );
  NAND U21655 ( .A(n88), .B(a[512]), .Z(n21095) );
  AND U21656 ( .A(n21096), .B(n21095), .Z(n21149) );
  XOR U21657 ( .A(a[509]), .B(n42197), .Z(n21138) );
  NANDN U21658 ( .A(n21138), .B(n42173), .Z(n21099) );
  NANDN U21659 ( .A(n21097), .B(n42172), .Z(n21098) );
  NAND U21660 ( .A(n21099), .B(n21098), .Z(n21147) );
  NAND U21661 ( .A(b[7]), .B(a[505]), .Z(n21148) );
  XNOR U21662 ( .A(n21147), .B(n21148), .Z(n21150) );
  XOR U21663 ( .A(n21149), .B(n21150), .Z(n21156) );
  NANDN U21664 ( .A(n21100), .B(n42093), .Z(n21102) );
  XOR U21665 ( .A(n42134), .B(a[511]), .Z(n21141) );
  NANDN U21666 ( .A(n21141), .B(n42095), .Z(n21101) );
  NAND U21667 ( .A(n21102), .B(n21101), .Z(n21154) );
  NANDN U21668 ( .A(n21103), .B(n42231), .Z(n21105) );
  XOR U21669 ( .A(n204), .B(a[507]), .Z(n21144) );
  NANDN U21670 ( .A(n21144), .B(n42234), .Z(n21104) );
  AND U21671 ( .A(n21105), .B(n21104), .Z(n21153) );
  XNOR U21672 ( .A(n21154), .B(n21153), .Z(n21155) );
  XNOR U21673 ( .A(n21156), .B(n21155), .Z(n21160) );
  NANDN U21674 ( .A(n21107), .B(n21106), .Z(n21111) );
  NAND U21675 ( .A(n21109), .B(n21108), .Z(n21110) );
  AND U21676 ( .A(n21111), .B(n21110), .Z(n21159) );
  XOR U21677 ( .A(n21160), .B(n21159), .Z(n21161) );
  NANDN U21678 ( .A(n21113), .B(n21112), .Z(n21117) );
  NANDN U21679 ( .A(n21115), .B(n21114), .Z(n21116) );
  NAND U21680 ( .A(n21117), .B(n21116), .Z(n21162) );
  XOR U21681 ( .A(n21161), .B(n21162), .Z(n21129) );
  OR U21682 ( .A(n21119), .B(n21118), .Z(n21123) );
  NANDN U21683 ( .A(n21121), .B(n21120), .Z(n21122) );
  NAND U21684 ( .A(n21123), .B(n21122), .Z(n21130) );
  XNOR U21685 ( .A(n21129), .B(n21130), .Z(n21131) );
  XNOR U21686 ( .A(n21132), .B(n21131), .Z(n21165) );
  XNOR U21687 ( .A(n21165), .B(sreg[1529]), .Z(n21167) );
  NAND U21688 ( .A(n21124), .B(sreg[1528]), .Z(n21128) );
  OR U21689 ( .A(n21126), .B(n21125), .Z(n21127) );
  AND U21690 ( .A(n21128), .B(n21127), .Z(n21166) );
  XOR U21691 ( .A(n21167), .B(n21166), .Z(c[1529]) );
  NANDN U21692 ( .A(n21130), .B(n21129), .Z(n21134) );
  NAND U21693 ( .A(n21132), .B(n21131), .Z(n21133) );
  NAND U21694 ( .A(n21134), .B(n21133), .Z(n21173) );
  NAND U21695 ( .A(b[0]), .B(a[514]), .Z(n21135) );
  XNOR U21696 ( .A(b[1]), .B(n21135), .Z(n21137) );
  NAND U21697 ( .A(n88), .B(a[513]), .Z(n21136) );
  AND U21698 ( .A(n21137), .B(n21136), .Z(n21190) );
  XOR U21699 ( .A(a[510]), .B(n42197), .Z(n21179) );
  NANDN U21700 ( .A(n21179), .B(n42173), .Z(n21140) );
  NANDN U21701 ( .A(n21138), .B(n42172), .Z(n21139) );
  NAND U21702 ( .A(n21140), .B(n21139), .Z(n21188) );
  NAND U21703 ( .A(b[7]), .B(a[506]), .Z(n21189) );
  XNOR U21704 ( .A(n21188), .B(n21189), .Z(n21191) );
  XOR U21705 ( .A(n21190), .B(n21191), .Z(n21197) );
  NANDN U21706 ( .A(n21141), .B(n42093), .Z(n21143) );
  XOR U21707 ( .A(n42134), .B(a[512]), .Z(n21182) );
  NANDN U21708 ( .A(n21182), .B(n42095), .Z(n21142) );
  NAND U21709 ( .A(n21143), .B(n21142), .Z(n21195) );
  NANDN U21710 ( .A(n21144), .B(n42231), .Z(n21146) );
  XOR U21711 ( .A(n204), .B(a[508]), .Z(n21185) );
  NANDN U21712 ( .A(n21185), .B(n42234), .Z(n21145) );
  AND U21713 ( .A(n21146), .B(n21145), .Z(n21194) );
  XNOR U21714 ( .A(n21195), .B(n21194), .Z(n21196) );
  XNOR U21715 ( .A(n21197), .B(n21196), .Z(n21201) );
  NANDN U21716 ( .A(n21148), .B(n21147), .Z(n21152) );
  NAND U21717 ( .A(n21150), .B(n21149), .Z(n21151) );
  AND U21718 ( .A(n21152), .B(n21151), .Z(n21200) );
  XOR U21719 ( .A(n21201), .B(n21200), .Z(n21202) );
  NANDN U21720 ( .A(n21154), .B(n21153), .Z(n21158) );
  NANDN U21721 ( .A(n21156), .B(n21155), .Z(n21157) );
  NAND U21722 ( .A(n21158), .B(n21157), .Z(n21203) );
  XOR U21723 ( .A(n21202), .B(n21203), .Z(n21170) );
  OR U21724 ( .A(n21160), .B(n21159), .Z(n21164) );
  NANDN U21725 ( .A(n21162), .B(n21161), .Z(n21163) );
  NAND U21726 ( .A(n21164), .B(n21163), .Z(n21171) );
  XNOR U21727 ( .A(n21170), .B(n21171), .Z(n21172) );
  XNOR U21728 ( .A(n21173), .B(n21172), .Z(n21206) );
  XNOR U21729 ( .A(n21206), .B(sreg[1530]), .Z(n21208) );
  NAND U21730 ( .A(n21165), .B(sreg[1529]), .Z(n21169) );
  OR U21731 ( .A(n21167), .B(n21166), .Z(n21168) );
  AND U21732 ( .A(n21169), .B(n21168), .Z(n21207) );
  XOR U21733 ( .A(n21208), .B(n21207), .Z(c[1530]) );
  NANDN U21734 ( .A(n21171), .B(n21170), .Z(n21175) );
  NAND U21735 ( .A(n21173), .B(n21172), .Z(n21174) );
  NAND U21736 ( .A(n21175), .B(n21174), .Z(n21214) );
  NAND U21737 ( .A(b[0]), .B(a[515]), .Z(n21176) );
  XNOR U21738 ( .A(b[1]), .B(n21176), .Z(n21178) );
  NAND U21739 ( .A(n88), .B(a[514]), .Z(n21177) );
  AND U21740 ( .A(n21178), .B(n21177), .Z(n21231) );
  XOR U21741 ( .A(a[511]), .B(n42197), .Z(n21220) );
  NANDN U21742 ( .A(n21220), .B(n42173), .Z(n21181) );
  NANDN U21743 ( .A(n21179), .B(n42172), .Z(n21180) );
  NAND U21744 ( .A(n21181), .B(n21180), .Z(n21229) );
  NAND U21745 ( .A(b[7]), .B(a[507]), .Z(n21230) );
  XNOR U21746 ( .A(n21229), .B(n21230), .Z(n21232) );
  XOR U21747 ( .A(n21231), .B(n21232), .Z(n21238) );
  NANDN U21748 ( .A(n21182), .B(n42093), .Z(n21184) );
  XOR U21749 ( .A(n42134), .B(a[513]), .Z(n21223) );
  NANDN U21750 ( .A(n21223), .B(n42095), .Z(n21183) );
  NAND U21751 ( .A(n21184), .B(n21183), .Z(n21236) );
  NANDN U21752 ( .A(n21185), .B(n42231), .Z(n21187) );
  XOR U21753 ( .A(n204), .B(a[509]), .Z(n21226) );
  NANDN U21754 ( .A(n21226), .B(n42234), .Z(n21186) );
  AND U21755 ( .A(n21187), .B(n21186), .Z(n21235) );
  XNOR U21756 ( .A(n21236), .B(n21235), .Z(n21237) );
  XNOR U21757 ( .A(n21238), .B(n21237), .Z(n21242) );
  NANDN U21758 ( .A(n21189), .B(n21188), .Z(n21193) );
  NAND U21759 ( .A(n21191), .B(n21190), .Z(n21192) );
  AND U21760 ( .A(n21193), .B(n21192), .Z(n21241) );
  XOR U21761 ( .A(n21242), .B(n21241), .Z(n21243) );
  NANDN U21762 ( .A(n21195), .B(n21194), .Z(n21199) );
  NANDN U21763 ( .A(n21197), .B(n21196), .Z(n21198) );
  NAND U21764 ( .A(n21199), .B(n21198), .Z(n21244) );
  XOR U21765 ( .A(n21243), .B(n21244), .Z(n21211) );
  OR U21766 ( .A(n21201), .B(n21200), .Z(n21205) );
  NANDN U21767 ( .A(n21203), .B(n21202), .Z(n21204) );
  NAND U21768 ( .A(n21205), .B(n21204), .Z(n21212) );
  XNOR U21769 ( .A(n21211), .B(n21212), .Z(n21213) );
  XNOR U21770 ( .A(n21214), .B(n21213), .Z(n21247) );
  XNOR U21771 ( .A(n21247), .B(sreg[1531]), .Z(n21249) );
  NAND U21772 ( .A(n21206), .B(sreg[1530]), .Z(n21210) );
  OR U21773 ( .A(n21208), .B(n21207), .Z(n21209) );
  AND U21774 ( .A(n21210), .B(n21209), .Z(n21248) );
  XOR U21775 ( .A(n21249), .B(n21248), .Z(c[1531]) );
  NANDN U21776 ( .A(n21212), .B(n21211), .Z(n21216) );
  NAND U21777 ( .A(n21214), .B(n21213), .Z(n21215) );
  NAND U21778 ( .A(n21216), .B(n21215), .Z(n21255) );
  NAND U21779 ( .A(b[0]), .B(a[516]), .Z(n21217) );
  XNOR U21780 ( .A(b[1]), .B(n21217), .Z(n21219) );
  NAND U21781 ( .A(n88), .B(a[515]), .Z(n21218) );
  AND U21782 ( .A(n21219), .B(n21218), .Z(n21272) );
  XOR U21783 ( .A(a[512]), .B(n42197), .Z(n21261) );
  NANDN U21784 ( .A(n21261), .B(n42173), .Z(n21222) );
  NANDN U21785 ( .A(n21220), .B(n42172), .Z(n21221) );
  NAND U21786 ( .A(n21222), .B(n21221), .Z(n21270) );
  NAND U21787 ( .A(b[7]), .B(a[508]), .Z(n21271) );
  XNOR U21788 ( .A(n21270), .B(n21271), .Z(n21273) );
  XOR U21789 ( .A(n21272), .B(n21273), .Z(n21279) );
  NANDN U21790 ( .A(n21223), .B(n42093), .Z(n21225) );
  XOR U21791 ( .A(n42134), .B(a[514]), .Z(n21264) );
  NANDN U21792 ( .A(n21264), .B(n42095), .Z(n21224) );
  NAND U21793 ( .A(n21225), .B(n21224), .Z(n21277) );
  NANDN U21794 ( .A(n21226), .B(n42231), .Z(n21228) );
  XOR U21795 ( .A(n204), .B(a[510]), .Z(n21267) );
  NANDN U21796 ( .A(n21267), .B(n42234), .Z(n21227) );
  AND U21797 ( .A(n21228), .B(n21227), .Z(n21276) );
  XNOR U21798 ( .A(n21277), .B(n21276), .Z(n21278) );
  XNOR U21799 ( .A(n21279), .B(n21278), .Z(n21283) );
  NANDN U21800 ( .A(n21230), .B(n21229), .Z(n21234) );
  NAND U21801 ( .A(n21232), .B(n21231), .Z(n21233) );
  AND U21802 ( .A(n21234), .B(n21233), .Z(n21282) );
  XOR U21803 ( .A(n21283), .B(n21282), .Z(n21284) );
  NANDN U21804 ( .A(n21236), .B(n21235), .Z(n21240) );
  NANDN U21805 ( .A(n21238), .B(n21237), .Z(n21239) );
  NAND U21806 ( .A(n21240), .B(n21239), .Z(n21285) );
  XOR U21807 ( .A(n21284), .B(n21285), .Z(n21252) );
  OR U21808 ( .A(n21242), .B(n21241), .Z(n21246) );
  NANDN U21809 ( .A(n21244), .B(n21243), .Z(n21245) );
  NAND U21810 ( .A(n21246), .B(n21245), .Z(n21253) );
  XNOR U21811 ( .A(n21252), .B(n21253), .Z(n21254) );
  XNOR U21812 ( .A(n21255), .B(n21254), .Z(n21288) );
  XNOR U21813 ( .A(n21288), .B(sreg[1532]), .Z(n21290) );
  NAND U21814 ( .A(n21247), .B(sreg[1531]), .Z(n21251) );
  OR U21815 ( .A(n21249), .B(n21248), .Z(n21250) );
  AND U21816 ( .A(n21251), .B(n21250), .Z(n21289) );
  XOR U21817 ( .A(n21290), .B(n21289), .Z(c[1532]) );
  NANDN U21818 ( .A(n21253), .B(n21252), .Z(n21257) );
  NAND U21819 ( .A(n21255), .B(n21254), .Z(n21256) );
  NAND U21820 ( .A(n21257), .B(n21256), .Z(n21296) );
  NAND U21821 ( .A(b[0]), .B(a[517]), .Z(n21258) );
  XNOR U21822 ( .A(b[1]), .B(n21258), .Z(n21260) );
  NAND U21823 ( .A(n88), .B(a[516]), .Z(n21259) );
  AND U21824 ( .A(n21260), .B(n21259), .Z(n21313) );
  XOR U21825 ( .A(a[513]), .B(n42197), .Z(n21302) );
  NANDN U21826 ( .A(n21302), .B(n42173), .Z(n21263) );
  NANDN U21827 ( .A(n21261), .B(n42172), .Z(n21262) );
  NAND U21828 ( .A(n21263), .B(n21262), .Z(n21311) );
  NAND U21829 ( .A(b[7]), .B(a[509]), .Z(n21312) );
  XNOR U21830 ( .A(n21311), .B(n21312), .Z(n21314) );
  XOR U21831 ( .A(n21313), .B(n21314), .Z(n21320) );
  NANDN U21832 ( .A(n21264), .B(n42093), .Z(n21266) );
  XOR U21833 ( .A(n42134), .B(a[515]), .Z(n21305) );
  NANDN U21834 ( .A(n21305), .B(n42095), .Z(n21265) );
  NAND U21835 ( .A(n21266), .B(n21265), .Z(n21318) );
  NANDN U21836 ( .A(n21267), .B(n42231), .Z(n21269) );
  XOR U21837 ( .A(n204), .B(a[511]), .Z(n21308) );
  NANDN U21838 ( .A(n21308), .B(n42234), .Z(n21268) );
  AND U21839 ( .A(n21269), .B(n21268), .Z(n21317) );
  XNOR U21840 ( .A(n21318), .B(n21317), .Z(n21319) );
  XNOR U21841 ( .A(n21320), .B(n21319), .Z(n21324) );
  NANDN U21842 ( .A(n21271), .B(n21270), .Z(n21275) );
  NAND U21843 ( .A(n21273), .B(n21272), .Z(n21274) );
  AND U21844 ( .A(n21275), .B(n21274), .Z(n21323) );
  XOR U21845 ( .A(n21324), .B(n21323), .Z(n21325) );
  NANDN U21846 ( .A(n21277), .B(n21276), .Z(n21281) );
  NANDN U21847 ( .A(n21279), .B(n21278), .Z(n21280) );
  NAND U21848 ( .A(n21281), .B(n21280), .Z(n21326) );
  XOR U21849 ( .A(n21325), .B(n21326), .Z(n21293) );
  OR U21850 ( .A(n21283), .B(n21282), .Z(n21287) );
  NANDN U21851 ( .A(n21285), .B(n21284), .Z(n21286) );
  NAND U21852 ( .A(n21287), .B(n21286), .Z(n21294) );
  XNOR U21853 ( .A(n21293), .B(n21294), .Z(n21295) );
  XNOR U21854 ( .A(n21296), .B(n21295), .Z(n21329) );
  XNOR U21855 ( .A(n21329), .B(sreg[1533]), .Z(n21331) );
  NAND U21856 ( .A(n21288), .B(sreg[1532]), .Z(n21292) );
  OR U21857 ( .A(n21290), .B(n21289), .Z(n21291) );
  AND U21858 ( .A(n21292), .B(n21291), .Z(n21330) );
  XOR U21859 ( .A(n21331), .B(n21330), .Z(c[1533]) );
  NANDN U21860 ( .A(n21294), .B(n21293), .Z(n21298) );
  NAND U21861 ( .A(n21296), .B(n21295), .Z(n21297) );
  NAND U21862 ( .A(n21298), .B(n21297), .Z(n21337) );
  NAND U21863 ( .A(b[0]), .B(a[518]), .Z(n21299) );
  XNOR U21864 ( .A(b[1]), .B(n21299), .Z(n21301) );
  NAND U21865 ( .A(n89), .B(a[517]), .Z(n21300) );
  AND U21866 ( .A(n21301), .B(n21300), .Z(n21354) );
  XOR U21867 ( .A(a[514]), .B(n42197), .Z(n21343) );
  NANDN U21868 ( .A(n21343), .B(n42173), .Z(n21304) );
  NANDN U21869 ( .A(n21302), .B(n42172), .Z(n21303) );
  NAND U21870 ( .A(n21304), .B(n21303), .Z(n21352) );
  NAND U21871 ( .A(b[7]), .B(a[510]), .Z(n21353) );
  XNOR U21872 ( .A(n21352), .B(n21353), .Z(n21355) );
  XOR U21873 ( .A(n21354), .B(n21355), .Z(n21361) );
  NANDN U21874 ( .A(n21305), .B(n42093), .Z(n21307) );
  XOR U21875 ( .A(n42134), .B(a[516]), .Z(n21346) );
  NANDN U21876 ( .A(n21346), .B(n42095), .Z(n21306) );
  NAND U21877 ( .A(n21307), .B(n21306), .Z(n21359) );
  NANDN U21878 ( .A(n21308), .B(n42231), .Z(n21310) );
  XOR U21879 ( .A(n204), .B(a[512]), .Z(n21349) );
  NANDN U21880 ( .A(n21349), .B(n42234), .Z(n21309) );
  AND U21881 ( .A(n21310), .B(n21309), .Z(n21358) );
  XNOR U21882 ( .A(n21359), .B(n21358), .Z(n21360) );
  XNOR U21883 ( .A(n21361), .B(n21360), .Z(n21365) );
  NANDN U21884 ( .A(n21312), .B(n21311), .Z(n21316) );
  NAND U21885 ( .A(n21314), .B(n21313), .Z(n21315) );
  AND U21886 ( .A(n21316), .B(n21315), .Z(n21364) );
  XOR U21887 ( .A(n21365), .B(n21364), .Z(n21366) );
  NANDN U21888 ( .A(n21318), .B(n21317), .Z(n21322) );
  NANDN U21889 ( .A(n21320), .B(n21319), .Z(n21321) );
  NAND U21890 ( .A(n21322), .B(n21321), .Z(n21367) );
  XOR U21891 ( .A(n21366), .B(n21367), .Z(n21334) );
  OR U21892 ( .A(n21324), .B(n21323), .Z(n21328) );
  NANDN U21893 ( .A(n21326), .B(n21325), .Z(n21327) );
  NAND U21894 ( .A(n21328), .B(n21327), .Z(n21335) );
  XNOR U21895 ( .A(n21334), .B(n21335), .Z(n21336) );
  XNOR U21896 ( .A(n21337), .B(n21336), .Z(n21370) );
  XNOR U21897 ( .A(n21370), .B(sreg[1534]), .Z(n21372) );
  NAND U21898 ( .A(n21329), .B(sreg[1533]), .Z(n21333) );
  OR U21899 ( .A(n21331), .B(n21330), .Z(n21332) );
  AND U21900 ( .A(n21333), .B(n21332), .Z(n21371) );
  XOR U21901 ( .A(n21372), .B(n21371), .Z(c[1534]) );
  NANDN U21902 ( .A(n21335), .B(n21334), .Z(n21339) );
  NAND U21903 ( .A(n21337), .B(n21336), .Z(n21338) );
  NAND U21904 ( .A(n21339), .B(n21338), .Z(n21378) );
  NAND U21905 ( .A(b[0]), .B(a[519]), .Z(n21340) );
  XNOR U21906 ( .A(b[1]), .B(n21340), .Z(n21342) );
  NAND U21907 ( .A(n89), .B(a[518]), .Z(n21341) );
  AND U21908 ( .A(n21342), .B(n21341), .Z(n21395) );
  XOR U21909 ( .A(a[515]), .B(n42197), .Z(n21384) );
  NANDN U21910 ( .A(n21384), .B(n42173), .Z(n21345) );
  NANDN U21911 ( .A(n21343), .B(n42172), .Z(n21344) );
  NAND U21912 ( .A(n21345), .B(n21344), .Z(n21393) );
  NAND U21913 ( .A(b[7]), .B(a[511]), .Z(n21394) );
  XNOR U21914 ( .A(n21393), .B(n21394), .Z(n21396) );
  XOR U21915 ( .A(n21395), .B(n21396), .Z(n21402) );
  NANDN U21916 ( .A(n21346), .B(n42093), .Z(n21348) );
  XOR U21917 ( .A(n42134), .B(a[517]), .Z(n21387) );
  NANDN U21918 ( .A(n21387), .B(n42095), .Z(n21347) );
  NAND U21919 ( .A(n21348), .B(n21347), .Z(n21400) );
  NANDN U21920 ( .A(n21349), .B(n42231), .Z(n21351) );
  XOR U21921 ( .A(n204), .B(a[513]), .Z(n21390) );
  NANDN U21922 ( .A(n21390), .B(n42234), .Z(n21350) );
  AND U21923 ( .A(n21351), .B(n21350), .Z(n21399) );
  XNOR U21924 ( .A(n21400), .B(n21399), .Z(n21401) );
  XNOR U21925 ( .A(n21402), .B(n21401), .Z(n21406) );
  NANDN U21926 ( .A(n21353), .B(n21352), .Z(n21357) );
  NAND U21927 ( .A(n21355), .B(n21354), .Z(n21356) );
  AND U21928 ( .A(n21357), .B(n21356), .Z(n21405) );
  XOR U21929 ( .A(n21406), .B(n21405), .Z(n21407) );
  NANDN U21930 ( .A(n21359), .B(n21358), .Z(n21363) );
  NANDN U21931 ( .A(n21361), .B(n21360), .Z(n21362) );
  NAND U21932 ( .A(n21363), .B(n21362), .Z(n21408) );
  XOR U21933 ( .A(n21407), .B(n21408), .Z(n21375) );
  OR U21934 ( .A(n21365), .B(n21364), .Z(n21369) );
  NANDN U21935 ( .A(n21367), .B(n21366), .Z(n21368) );
  NAND U21936 ( .A(n21369), .B(n21368), .Z(n21376) );
  XNOR U21937 ( .A(n21375), .B(n21376), .Z(n21377) );
  XNOR U21938 ( .A(n21378), .B(n21377), .Z(n21411) );
  XNOR U21939 ( .A(n21411), .B(sreg[1535]), .Z(n21413) );
  NAND U21940 ( .A(n21370), .B(sreg[1534]), .Z(n21374) );
  OR U21941 ( .A(n21372), .B(n21371), .Z(n21373) );
  AND U21942 ( .A(n21374), .B(n21373), .Z(n21412) );
  XOR U21943 ( .A(n21413), .B(n21412), .Z(c[1535]) );
  NANDN U21944 ( .A(n21376), .B(n21375), .Z(n21380) );
  NAND U21945 ( .A(n21378), .B(n21377), .Z(n21379) );
  NAND U21946 ( .A(n21380), .B(n21379), .Z(n21419) );
  NAND U21947 ( .A(b[0]), .B(a[520]), .Z(n21381) );
  XNOR U21948 ( .A(b[1]), .B(n21381), .Z(n21383) );
  NAND U21949 ( .A(n89), .B(a[519]), .Z(n21382) );
  AND U21950 ( .A(n21383), .B(n21382), .Z(n21436) );
  XOR U21951 ( .A(a[516]), .B(n42197), .Z(n21425) );
  NANDN U21952 ( .A(n21425), .B(n42173), .Z(n21386) );
  NANDN U21953 ( .A(n21384), .B(n42172), .Z(n21385) );
  NAND U21954 ( .A(n21386), .B(n21385), .Z(n21434) );
  NAND U21955 ( .A(b[7]), .B(a[512]), .Z(n21435) );
  XNOR U21956 ( .A(n21434), .B(n21435), .Z(n21437) );
  XOR U21957 ( .A(n21436), .B(n21437), .Z(n21443) );
  NANDN U21958 ( .A(n21387), .B(n42093), .Z(n21389) );
  XOR U21959 ( .A(n42134), .B(a[518]), .Z(n21428) );
  NANDN U21960 ( .A(n21428), .B(n42095), .Z(n21388) );
  NAND U21961 ( .A(n21389), .B(n21388), .Z(n21441) );
  NANDN U21962 ( .A(n21390), .B(n42231), .Z(n21392) );
  XOR U21963 ( .A(n204), .B(a[514]), .Z(n21431) );
  NANDN U21964 ( .A(n21431), .B(n42234), .Z(n21391) );
  AND U21965 ( .A(n21392), .B(n21391), .Z(n21440) );
  XNOR U21966 ( .A(n21441), .B(n21440), .Z(n21442) );
  XNOR U21967 ( .A(n21443), .B(n21442), .Z(n21447) );
  NANDN U21968 ( .A(n21394), .B(n21393), .Z(n21398) );
  NAND U21969 ( .A(n21396), .B(n21395), .Z(n21397) );
  AND U21970 ( .A(n21398), .B(n21397), .Z(n21446) );
  XOR U21971 ( .A(n21447), .B(n21446), .Z(n21448) );
  NANDN U21972 ( .A(n21400), .B(n21399), .Z(n21404) );
  NANDN U21973 ( .A(n21402), .B(n21401), .Z(n21403) );
  NAND U21974 ( .A(n21404), .B(n21403), .Z(n21449) );
  XOR U21975 ( .A(n21448), .B(n21449), .Z(n21416) );
  OR U21976 ( .A(n21406), .B(n21405), .Z(n21410) );
  NANDN U21977 ( .A(n21408), .B(n21407), .Z(n21409) );
  NAND U21978 ( .A(n21410), .B(n21409), .Z(n21417) );
  XNOR U21979 ( .A(n21416), .B(n21417), .Z(n21418) );
  XNOR U21980 ( .A(n21419), .B(n21418), .Z(n21452) );
  XNOR U21981 ( .A(n21452), .B(sreg[1536]), .Z(n21454) );
  NAND U21982 ( .A(n21411), .B(sreg[1535]), .Z(n21415) );
  OR U21983 ( .A(n21413), .B(n21412), .Z(n21414) );
  AND U21984 ( .A(n21415), .B(n21414), .Z(n21453) );
  XOR U21985 ( .A(n21454), .B(n21453), .Z(c[1536]) );
  NANDN U21986 ( .A(n21417), .B(n21416), .Z(n21421) );
  NAND U21987 ( .A(n21419), .B(n21418), .Z(n21420) );
  NAND U21988 ( .A(n21421), .B(n21420), .Z(n21460) );
  NAND U21989 ( .A(b[0]), .B(a[521]), .Z(n21422) );
  XNOR U21990 ( .A(b[1]), .B(n21422), .Z(n21424) );
  NAND U21991 ( .A(n89), .B(a[520]), .Z(n21423) );
  AND U21992 ( .A(n21424), .B(n21423), .Z(n21477) );
  XOR U21993 ( .A(a[517]), .B(n42197), .Z(n21466) );
  NANDN U21994 ( .A(n21466), .B(n42173), .Z(n21427) );
  NANDN U21995 ( .A(n21425), .B(n42172), .Z(n21426) );
  NAND U21996 ( .A(n21427), .B(n21426), .Z(n21475) );
  NAND U21997 ( .A(b[7]), .B(a[513]), .Z(n21476) );
  XNOR U21998 ( .A(n21475), .B(n21476), .Z(n21478) );
  XOR U21999 ( .A(n21477), .B(n21478), .Z(n21484) );
  NANDN U22000 ( .A(n21428), .B(n42093), .Z(n21430) );
  XOR U22001 ( .A(n42134), .B(a[519]), .Z(n21469) );
  NANDN U22002 ( .A(n21469), .B(n42095), .Z(n21429) );
  NAND U22003 ( .A(n21430), .B(n21429), .Z(n21482) );
  NANDN U22004 ( .A(n21431), .B(n42231), .Z(n21433) );
  XOR U22005 ( .A(n205), .B(a[515]), .Z(n21472) );
  NANDN U22006 ( .A(n21472), .B(n42234), .Z(n21432) );
  AND U22007 ( .A(n21433), .B(n21432), .Z(n21481) );
  XNOR U22008 ( .A(n21482), .B(n21481), .Z(n21483) );
  XNOR U22009 ( .A(n21484), .B(n21483), .Z(n21488) );
  NANDN U22010 ( .A(n21435), .B(n21434), .Z(n21439) );
  NAND U22011 ( .A(n21437), .B(n21436), .Z(n21438) );
  AND U22012 ( .A(n21439), .B(n21438), .Z(n21487) );
  XOR U22013 ( .A(n21488), .B(n21487), .Z(n21489) );
  NANDN U22014 ( .A(n21441), .B(n21440), .Z(n21445) );
  NANDN U22015 ( .A(n21443), .B(n21442), .Z(n21444) );
  NAND U22016 ( .A(n21445), .B(n21444), .Z(n21490) );
  XOR U22017 ( .A(n21489), .B(n21490), .Z(n21457) );
  OR U22018 ( .A(n21447), .B(n21446), .Z(n21451) );
  NANDN U22019 ( .A(n21449), .B(n21448), .Z(n21450) );
  NAND U22020 ( .A(n21451), .B(n21450), .Z(n21458) );
  XNOR U22021 ( .A(n21457), .B(n21458), .Z(n21459) );
  XNOR U22022 ( .A(n21460), .B(n21459), .Z(n21493) );
  XNOR U22023 ( .A(n21493), .B(sreg[1537]), .Z(n21495) );
  NAND U22024 ( .A(n21452), .B(sreg[1536]), .Z(n21456) );
  OR U22025 ( .A(n21454), .B(n21453), .Z(n21455) );
  AND U22026 ( .A(n21456), .B(n21455), .Z(n21494) );
  XOR U22027 ( .A(n21495), .B(n21494), .Z(c[1537]) );
  NANDN U22028 ( .A(n21458), .B(n21457), .Z(n21462) );
  NAND U22029 ( .A(n21460), .B(n21459), .Z(n21461) );
  NAND U22030 ( .A(n21462), .B(n21461), .Z(n21501) );
  NAND U22031 ( .A(b[0]), .B(a[522]), .Z(n21463) );
  XNOR U22032 ( .A(b[1]), .B(n21463), .Z(n21465) );
  NAND U22033 ( .A(n89), .B(a[521]), .Z(n21464) );
  AND U22034 ( .A(n21465), .B(n21464), .Z(n21518) );
  XOR U22035 ( .A(a[518]), .B(n42197), .Z(n21507) );
  NANDN U22036 ( .A(n21507), .B(n42173), .Z(n21468) );
  NANDN U22037 ( .A(n21466), .B(n42172), .Z(n21467) );
  NAND U22038 ( .A(n21468), .B(n21467), .Z(n21516) );
  NAND U22039 ( .A(b[7]), .B(a[514]), .Z(n21517) );
  XNOR U22040 ( .A(n21516), .B(n21517), .Z(n21519) );
  XOR U22041 ( .A(n21518), .B(n21519), .Z(n21525) );
  NANDN U22042 ( .A(n21469), .B(n42093), .Z(n21471) );
  XOR U22043 ( .A(n42134), .B(a[520]), .Z(n21510) );
  NANDN U22044 ( .A(n21510), .B(n42095), .Z(n21470) );
  NAND U22045 ( .A(n21471), .B(n21470), .Z(n21523) );
  NANDN U22046 ( .A(n21472), .B(n42231), .Z(n21474) );
  XOR U22047 ( .A(n205), .B(a[516]), .Z(n21513) );
  NANDN U22048 ( .A(n21513), .B(n42234), .Z(n21473) );
  AND U22049 ( .A(n21474), .B(n21473), .Z(n21522) );
  XNOR U22050 ( .A(n21523), .B(n21522), .Z(n21524) );
  XNOR U22051 ( .A(n21525), .B(n21524), .Z(n21529) );
  NANDN U22052 ( .A(n21476), .B(n21475), .Z(n21480) );
  NAND U22053 ( .A(n21478), .B(n21477), .Z(n21479) );
  AND U22054 ( .A(n21480), .B(n21479), .Z(n21528) );
  XOR U22055 ( .A(n21529), .B(n21528), .Z(n21530) );
  NANDN U22056 ( .A(n21482), .B(n21481), .Z(n21486) );
  NANDN U22057 ( .A(n21484), .B(n21483), .Z(n21485) );
  NAND U22058 ( .A(n21486), .B(n21485), .Z(n21531) );
  XOR U22059 ( .A(n21530), .B(n21531), .Z(n21498) );
  OR U22060 ( .A(n21488), .B(n21487), .Z(n21492) );
  NANDN U22061 ( .A(n21490), .B(n21489), .Z(n21491) );
  NAND U22062 ( .A(n21492), .B(n21491), .Z(n21499) );
  XNOR U22063 ( .A(n21498), .B(n21499), .Z(n21500) );
  XNOR U22064 ( .A(n21501), .B(n21500), .Z(n21534) );
  XNOR U22065 ( .A(n21534), .B(sreg[1538]), .Z(n21536) );
  NAND U22066 ( .A(n21493), .B(sreg[1537]), .Z(n21497) );
  OR U22067 ( .A(n21495), .B(n21494), .Z(n21496) );
  AND U22068 ( .A(n21497), .B(n21496), .Z(n21535) );
  XOR U22069 ( .A(n21536), .B(n21535), .Z(c[1538]) );
  NANDN U22070 ( .A(n21499), .B(n21498), .Z(n21503) );
  NAND U22071 ( .A(n21501), .B(n21500), .Z(n21502) );
  NAND U22072 ( .A(n21503), .B(n21502), .Z(n21542) );
  NAND U22073 ( .A(b[0]), .B(a[523]), .Z(n21504) );
  XNOR U22074 ( .A(b[1]), .B(n21504), .Z(n21506) );
  NAND U22075 ( .A(n89), .B(a[522]), .Z(n21505) );
  AND U22076 ( .A(n21506), .B(n21505), .Z(n21559) );
  XOR U22077 ( .A(a[519]), .B(n42197), .Z(n21548) );
  NANDN U22078 ( .A(n21548), .B(n42173), .Z(n21509) );
  NANDN U22079 ( .A(n21507), .B(n42172), .Z(n21508) );
  NAND U22080 ( .A(n21509), .B(n21508), .Z(n21557) );
  NAND U22081 ( .A(b[7]), .B(a[515]), .Z(n21558) );
  XNOR U22082 ( .A(n21557), .B(n21558), .Z(n21560) );
  XOR U22083 ( .A(n21559), .B(n21560), .Z(n21566) );
  NANDN U22084 ( .A(n21510), .B(n42093), .Z(n21512) );
  XOR U22085 ( .A(n42134), .B(a[521]), .Z(n21551) );
  NANDN U22086 ( .A(n21551), .B(n42095), .Z(n21511) );
  NAND U22087 ( .A(n21512), .B(n21511), .Z(n21564) );
  NANDN U22088 ( .A(n21513), .B(n42231), .Z(n21515) );
  XOR U22089 ( .A(n205), .B(a[517]), .Z(n21554) );
  NANDN U22090 ( .A(n21554), .B(n42234), .Z(n21514) );
  AND U22091 ( .A(n21515), .B(n21514), .Z(n21563) );
  XNOR U22092 ( .A(n21564), .B(n21563), .Z(n21565) );
  XNOR U22093 ( .A(n21566), .B(n21565), .Z(n21570) );
  NANDN U22094 ( .A(n21517), .B(n21516), .Z(n21521) );
  NAND U22095 ( .A(n21519), .B(n21518), .Z(n21520) );
  AND U22096 ( .A(n21521), .B(n21520), .Z(n21569) );
  XOR U22097 ( .A(n21570), .B(n21569), .Z(n21571) );
  NANDN U22098 ( .A(n21523), .B(n21522), .Z(n21527) );
  NANDN U22099 ( .A(n21525), .B(n21524), .Z(n21526) );
  NAND U22100 ( .A(n21527), .B(n21526), .Z(n21572) );
  XOR U22101 ( .A(n21571), .B(n21572), .Z(n21539) );
  OR U22102 ( .A(n21529), .B(n21528), .Z(n21533) );
  NANDN U22103 ( .A(n21531), .B(n21530), .Z(n21532) );
  NAND U22104 ( .A(n21533), .B(n21532), .Z(n21540) );
  XNOR U22105 ( .A(n21539), .B(n21540), .Z(n21541) );
  XNOR U22106 ( .A(n21542), .B(n21541), .Z(n21575) );
  XNOR U22107 ( .A(n21575), .B(sreg[1539]), .Z(n21577) );
  NAND U22108 ( .A(n21534), .B(sreg[1538]), .Z(n21538) );
  OR U22109 ( .A(n21536), .B(n21535), .Z(n21537) );
  AND U22110 ( .A(n21538), .B(n21537), .Z(n21576) );
  XOR U22111 ( .A(n21577), .B(n21576), .Z(c[1539]) );
  NANDN U22112 ( .A(n21540), .B(n21539), .Z(n21544) );
  NAND U22113 ( .A(n21542), .B(n21541), .Z(n21543) );
  NAND U22114 ( .A(n21544), .B(n21543), .Z(n21583) );
  NAND U22115 ( .A(b[0]), .B(a[524]), .Z(n21545) );
  XNOR U22116 ( .A(b[1]), .B(n21545), .Z(n21547) );
  NAND U22117 ( .A(n89), .B(a[523]), .Z(n21546) );
  AND U22118 ( .A(n21547), .B(n21546), .Z(n21600) );
  XOR U22119 ( .A(a[520]), .B(n42197), .Z(n21589) );
  NANDN U22120 ( .A(n21589), .B(n42173), .Z(n21550) );
  NANDN U22121 ( .A(n21548), .B(n42172), .Z(n21549) );
  NAND U22122 ( .A(n21550), .B(n21549), .Z(n21598) );
  NAND U22123 ( .A(b[7]), .B(a[516]), .Z(n21599) );
  XNOR U22124 ( .A(n21598), .B(n21599), .Z(n21601) );
  XOR U22125 ( .A(n21600), .B(n21601), .Z(n21607) );
  NANDN U22126 ( .A(n21551), .B(n42093), .Z(n21553) );
  XOR U22127 ( .A(n42134), .B(a[522]), .Z(n21592) );
  NANDN U22128 ( .A(n21592), .B(n42095), .Z(n21552) );
  NAND U22129 ( .A(n21553), .B(n21552), .Z(n21605) );
  NANDN U22130 ( .A(n21554), .B(n42231), .Z(n21556) );
  XOR U22131 ( .A(n205), .B(a[518]), .Z(n21595) );
  NANDN U22132 ( .A(n21595), .B(n42234), .Z(n21555) );
  AND U22133 ( .A(n21556), .B(n21555), .Z(n21604) );
  XNOR U22134 ( .A(n21605), .B(n21604), .Z(n21606) );
  XNOR U22135 ( .A(n21607), .B(n21606), .Z(n21611) );
  NANDN U22136 ( .A(n21558), .B(n21557), .Z(n21562) );
  NAND U22137 ( .A(n21560), .B(n21559), .Z(n21561) );
  AND U22138 ( .A(n21562), .B(n21561), .Z(n21610) );
  XOR U22139 ( .A(n21611), .B(n21610), .Z(n21612) );
  NANDN U22140 ( .A(n21564), .B(n21563), .Z(n21568) );
  NANDN U22141 ( .A(n21566), .B(n21565), .Z(n21567) );
  NAND U22142 ( .A(n21568), .B(n21567), .Z(n21613) );
  XOR U22143 ( .A(n21612), .B(n21613), .Z(n21580) );
  OR U22144 ( .A(n21570), .B(n21569), .Z(n21574) );
  NANDN U22145 ( .A(n21572), .B(n21571), .Z(n21573) );
  NAND U22146 ( .A(n21574), .B(n21573), .Z(n21581) );
  XNOR U22147 ( .A(n21580), .B(n21581), .Z(n21582) );
  XNOR U22148 ( .A(n21583), .B(n21582), .Z(n21616) );
  XNOR U22149 ( .A(n21616), .B(sreg[1540]), .Z(n21618) );
  NAND U22150 ( .A(n21575), .B(sreg[1539]), .Z(n21579) );
  OR U22151 ( .A(n21577), .B(n21576), .Z(n21578) );
  AND U22152 ( .A(n21579), .B(n21578), .Z(n21617) );
  XOR U22153 ( .A(n21618), .B(n21617), .Z(c[1540]) );
  NANDN U22154 ( .A(n21581), .B(n21580), .Z(n21585) );
  NAND U22155 ( .A(n21583), .B(n21582), .Z(n21584) );
  NAND U22156 ( .A(n21585), .B(n21584), .Z(n21624) );
  NAND U22157 ( .A(b[0]), .B(a[525]), .Z(n21586) );
  XNOR U22158 ( .A(b[1]), .B(n21586), .Z(n21588) );
  NAND U22159 ( .A(n90), .B(a[524]), .Z(n21587) );
  AND U22160 ( .A(n21588), .B(n21587), .Z(n21641) );
  XOR U22161 ( .A(a[521]), .B(n42197), .Z(n21630) );
  NANDN U22162 ( .A(n21630), .B(n42173), .Z(n21591) );
  NANDN U22163 ( .A(n21589), .B(n42172), .Z(n21590) );
  NAND U22164 ( .A(n21591), .B(n21590), .Z(n21639) );
  NAND U22165 ( .A(b[7]), .B(a[517]), .Z(n21640) );
  XNOR U22166 ( .A(n21639), .B(n21640), .Z(n21642) );
  XOR U22167 ( .A(n21641), .B(n21642), .Z(n21648) );
  NANDN U22168 ( .A(n21592), .B(n42093), .Z(n21594) );
  XOR U22169 ( .A(n42134), .B(a[523]), .Z(n21633) );
  NANDN U22170 ( .A(n21633), .B(n42095), .Z(n21593) );
  NAND U22171 ( .A(n21594), .B(n21593), .Z(n21646) );
  NANDN U22172 ( .A(n21595), .B(n42231), .Z(n21597) );
  XOR U22173 ( .A(n205), .B(a[519]), .Z(n21636) );
  NANDN U22174 ( .A(n21636), .B(n42234), .Z(n21596) );
  AND U22175 ( .A(n21597), .B(n21596), .Z(n21645) );
  XNOR U22176 ( .A(n21646), .B(n21645), .Z(n21647) );
  XNOR U22177 ( .A(n21648), .B(n21647), .Z(n21652) );
  NANDN U22178 ( .A(n21599), .B(n21598), .Z(n21603) );
  NAND U22179 ( .A(n21601), .B(n21600), .Z(n21602) );
  AND U22180 ( .A(n21603), .B(n21602), .Z(n21651) );
  XOR U22181 ( .A(n21652), .B(n21651), .Z(n21653) );
  NANDN U22182 ( .A(n21605), .B(n21604), .Z(n21609) );
  NANDN U22183 ( .A(n21607), .B(n21606), .Z(n21608) );
  NAND U22184 ( .A(n21609), .B(n21608), .Z(n21654) );
  XOR U22185 ( .A(n21653), .B(n21654), .Z(n21621) );
  OR U22186 ( .A(n21611), .B(n21610), .Z(n21615) );
  NANDN U22187 ( .A(n21613), .B(n21612), .Z(n21614) );
  NAND U22188 ( .A(n21615), .B(n21614), .Z(n21622) );
  XNOR U22189 ( .A(n21621), .B(n21622), .Z(n21623) );
  XNOR U22190 ( .A(n21624), .B(n21623), .Z(n21657) );
  XNOR U22191 ( .A(n21657), .B(sreg[1541]), .Z(n21659) );
  NAND U22192 ( .A(n21616), .B(sreg[1540]), .Z(n21620) );
  OR U22193 ( .A(n21618), .B(n21617), .Z(n21619) );
  AND U22194 ( .A(n21620), .B(n21619), .Z(n21658) );
  XOR U22195 ( .A(n21659), .B(n21658), .Z(c[1541]) );
  NANDN U22196 ( .A(n21622), .B(n21621), .Z(n21626) );
  NAND U22197 ( .A(n21624), .B(n21623), .Z(n21625) );
  NAND U22198 ( .A(n21626), .B(n21625), .Z(n21665) );
  NAND U22199 ( .A(b[0]), .B(a[526]), .Z(n21627) );
  XNOR U22200 ( .A(b[1]), .B(n21627), .Z(n21629) );
  NAND U22201 ( .A(n90), .B(a[525]), .Z(n21628) );
  AND U22202 ( .A(n21629), .B(n21628), .Z(n21682) );
  XOR U22203 ( .A(a[522]), .B(n42197), .Z(n21671) );
  NANDN U22204 ( .A(n21671), .B(n42173), .Z(n21632) );
  NANDN U22205 ( .A(n21630), .B(n42172), .Z(n21631) );
  NAND U22206 ( .A(n21632), .B(n21631), .Z(n21680) );
  NAND U22207 ( .A(b[7]), .B(a[518]), .Z(n21681) );
  XNOR U22208 ( .A(n21680), .B(n21681), .Z(n21683) );
  XOR U22209 ( .A(n21682), .B(n21683), .Z(n21689) );
  NANDN U22210 ( .A(n21633), .B(n42093), .Z(n21635) );
  XOR U22211 ( .A(n42134), .B(a[524]), .Z(n21674) );
  NANDN U22212 ( .A(n21674), .B(n42095), .Z(n21634) );
  NAND U22213 ( .A(n21635), .B(n21634), .Z(n21687) );
  NANDN U22214 ( .A(n21636), .B(n42231), .Z(n21638) );
  XOR U22215 ( .A(n205), .B(a[520]), .Z(n21677) );
  NANDN U22216 ( .A(n21677), .B(n42234), .Z(n21637) );
  AND U22217 ( .A(n21638), .B(n21637), .Z(n21686) );
  XNOR U22218 ( .A(n21687), .B(n21686), .Z(n21688) );
  XNOR U22219 ( .A(n21689), .B(n21688), .Z(n21693) );
  NANDN U22220 ( .A(n21640), .B(n21639), .Z(n21644) );
  NAND U22221 ( .A(n21642), .B(n21641), .Z(n21643) );
  AND U22222 ( .A(n21644), .B(n21643), .Z(n21692) );
  XOR U22223 ( .A(n21693), .B(n21692), .Z(n21694) );
  NANDN U22224 ( .A(n21646), .B(n21645), .Z(n21650) );
  NANDN U22225 ( .A(n21648), .B(n21647), .Z(n21649) );
  NAND U22226 ( .A(n21650), .B(n21649), .Z(n21695) );
  XOR U22227 ( .A(n21694), .B(n21695), .Z(n21662) );
  OR U22228 ( .A(n21652), .B(n21651), .Z(n21656) );
  NANDN U22229 ( .A(n21654), .B(n21653), .Z(n21655) );
  NAND U22230 ( .A(n21656), .B(n21655), .Z(n21663) );
  XNOR U22231 ( .A(n21662), .B(n21663), .Z(n21664) );
  XNOR U22232 ( .A(n21665), .B(n21664), .Z(n21698) );
  XNOR U22233 ( .A(n21698), .B(sreg[1542]), .Z(n21700) );
  NAND U22234 ( .A(n21657), .B(sreg[1541]), .Z(n21661) );
  OR U22235 ( .A(n21659), .B(n21658), .Z(n21660) );
  AND U22236 ( .A(n21661), .B(n21660), .Z(n21699) );
  XOR U22237 ( .A(n21700), .B(n21699), .Z(c[1542]) );
  NANDN U22238 ( .A(n21663), .B(n21662), .Z(n21667) );
  NAND U22239 ( .A(n21665), .B(n21664), .Z(n21666) );
  NAND U22240 ( .A(n21667), .B(n21666), .Z(n21706) );
  NAND U22241 ( .A(b[0]), .B(a[527]), .Z(n21668) );
  XNOR U22242 ( .A(b[1]), .B(n21668), .Z(n21670) );
  NAND U22243 ( .A(n90), .B(a[526]), .Z(n21669) );
  AND U22244 ( .A(n21670), .B(n21669), .Z(n21723) );
  XOR U22245 ( .A(a[523]), .B(n42197), .Z(n21712) );
  NANDN U22246 ( .A(n21712), .B(n42173), .Z(n21673) );
  NANDN U22247 ( .A(n21671), .B(n42172), .Z(n21672) );
  NAND U22248 ( .A(n21673), .B(n21672), .Z(n21721) );
  NAND U22249 ( .A(b[7]), .B(a[519]), .Z(n21722) );
  XNOR U22250 ( .A(n21721), .B(n21722), .Z(n21724) );
  XOR U22251 ( .A(n21723), .B(n21724), .Z(n21730) );
  NANDN U22252 ( .A(n21674), .B(n42093), .Z(n21676) );
  XOR U22253 ( .A(n42134), .B(a[525]), .Z(n21715) );
  NANDN U22254 ( .A(n21715), .B(n42095), .Z(n21675) );
  NAND U22255 ( .A(n21676), .B(n21675), .Z(n21728) );
  NANDN U22256 ( .A(n21677), .B(n42231), .Z(n21679) );
  XOR U22257 ( .A(n205), .B(a[521]), .Z(n21718) );
  NANDN U22258 ( .A(n21718), .B(n42234), .Z(n21678) );
  AND U22259 ( .A(n21679), .B(n21678), .Z(n21727) );
  XNOR U22260 ( .A(n21728), .B(n21727), .Z(n21729) );
  XNOR U22261 ( .A(n21730), .B(n21729), .Z(n21734) );
  NANDN U22262 ( .A(n21681), .B(n21680), .Z(n21685) );
  NAND U22263 ( .A(n21683), .B(n21682), .Z(n21684) );
  AND U22264 ( .A(n21685), .B(n21684), .Z(n21733) );
  XOR U22265 ( .A(n21734), .B(n21733), .Z(n21735) );
  NANDN U22266 ( .A(n21687), .B(n21686), .Z(n21691) );
  NANDN U22267 ( .A(n21689), .B(n21688), .Z(n21690) );
  NAND U22268 ( .A(n21691), .B(n21690), .Z(n21736) );
  XOR U22269 ( .A(n21735), .B(n21736), .Z(n21703) );
  OR U22270 ( .A(n21693), .B(n21692), .Z(n21697) );
  NANDN U22271 ( .A(n21695), .B(n21694), .Z(n21696) );
  NAND U22272 ( .A(n21697), .B(n21696), .Z(n21704) );
  XNOR U22273 ( .A(n21703), .B(n21704), .Z(n21705) );
  XNOR U22274 ( .A(n21706), .B(n21705), .Z(n21739) );
  XNOR U22275 ( .A(n21739), .B(sreg[1543]), .Z(n21741) );
  NAND U22276 ( .A(n21698), .B(sreg[1542]), .Z(n21702) );
  OR U22277 ( .A(n21700), .B(n21699), .Z(n21701) );
  AND U22278 ( .A(n21702), .B(n21701), .Z(n21740) );
  XOR U22279 ( .A(n21741), .B(n21740), .Z(c[1543]) );
  NANDN U22280 ( .A(n21704), .B(n21703), .Z(n21708) );
  NAND U22281 ( .A(n21706), .B(n21705), .Z(n21707) );
  NAND U22282 ( .A(n21708), .B(n21707), .Z(n21747) );
  NAND U22283 ( .A(b[0]), .B(a[528]), .Z(n21709) );
  XNOR U22284 ( .A(b[1]), .B(n21709), .Z(n21711) );
  NAND U22285 ( .A(n90), .B(a[527]), .Z(n21710) );
  AND U22286 ( .A(n21711), .B(n21710), .Z(n21764) );
  XOR U22287 ( .A(a[524]), .B(n42197), .Z(n21753) );
  NANDN U22288 ( .A(n21753), .B(n42173), .Z(n21714) );
  NANDN U22289 ( .A(n21712), .B(n42172), .Z(n21713) );
  NAND U22290 ( .A(n21714), .B(n21713), .Z(n21762) );
  NAND U22291 ( .A(b[7]), .B(a[520]), .Z(n21763) );
  XNOR U22292 ( .A(n21762), .B(n21763), .Z(n21765) );
  XOR U22293 ( .A(n21764), .B(n21765), .Z(n21771) );
  NANDN U22294 ( .A(n21715), .B(n42093), .Z(n21717) );
  XOR U22295 ( .A(n42134), .B(a[526]), .Z(n21756) );
  NANDN U22296 ( .A(n21756), .B(n42095), .Z(n21716) );
  NAND U22297 ( .A(n21717), .B(n21716), .Z(n21769) );
  NANDN U22298 ( .A(n21718), .B(n42231), .Z(n21720) );
  XOR U22299 ( .A(n205), .B(a[522]), .Z(n21759) );
  NANDN U22300 ( .A(n21759), .B(n42234), .Z(n21719) );
  AND U22301 ( .A(n21720), .B(n21719), .Z(n21768) );
  XNOR U22302 ( .A(n21769), .B(n21768), .Z(n21770) );
  XNOR U22303 ( .A(n21771), .B(n21770), .Z(n21775) );
  NANDN U22304 ( .A(n21722), .B(n21721), .Z(n21726) );
  NAND U22305 ( .A(n21724), .B(n21723), .Z(n21725) );
  AND U22306 ( .A(n21726), .B(n21725), .Z(n21774) );
  XOR U22307 ( .A(n21775), .B(n21774), .Z(n21776) );
  NANDN U22308 ( .A(n21728), .B(n21727), .Z(n21732) );
  NANDN U22309 ( .A(n21730), .B(n21729), .Z(n21731) );
  NAND U22310 ( .A(n21732), .B(n21731), .Z(n21777) );
  XOR U22311 ( .A(n21776), .B(n21777), .Z(n21744) );
  OR U22312 ( .A(n21734), .B(n21733), .Z(n21738) );
  NANDN U22313 ( .A(n21736), .B(n21735), .Z(n21737) );
  NAND U22314 ( .A(n21738), .B(n21737), .Z(n21745) );
  XNOR U22315 ( .A(n21744), .B(n21745), .Z(n21746) );
  XNOR U22316 ( .A(n21747), .B(n21746), .Z(n21780) );
  XNOR U22317 ( .A(n21780), .B(sreg[1544]), .Z(n21782) );
  NAND U22318 ( .A(n21739), .B(sreg[1543]), .Z(n21743) );
  OR U22319 ( .A(n21741), .B(n21740), .Z(n21742) );
  AND U22320 ( .A(n21743), .B(n21742), .Z(n21781) );
  XOR U22321 ( .A(n21782), .B(n21781), .Z(c[1544]) );
  NANDN U22322 ( .A(n21745), .B(n21744), .Z(n21749) );
  NAND U22323 ( .A(n21747), .B(n21746), .Z(n21748) );
  NAND U22324 ( .A(n21749), .B(n21748), .Z(n21788) );
  NAND U22325 ( .A(b[0]), .B(a[529]), .Z(n21750) );
  XNOR U22326 ( .A(b[1]), .B(n21750), .Z(n21752) );
  NAND U22327 ( .A(n90), .B(a[528]), .Z(n21751) );
  AND U22328 ( .A(n21752), .B(n21751), .Z(n21805) );
  XOR U22329 ( .A(a[525]), .B(n42197), .Z(n21794) );
  NANDN U22330 ( .A(n21794), .B(n42173), .Z(n21755) );
  NANDN U22331 ( .A(n21753), .B(n42172), .Z(n21754) );
  NAND U22332 ( .A(n21755), .B(n21754), .Z(n21803) );
  NAND U22333 ( .A(b[7]), .B(a[521]), .Z(n21804) );
  XNOR U22334 ( .A(n21803), .B(n21804), .Z(n21806) );
  XOR U22335 ( .A(n21805), .B(n21806), .Z(n21812) );
  NANDN U22336 ( .A(n21756), .B(n42093), .Z(n21758) );
  XOR U22337 ( .A(n42134), .B(a[527]), .Z(n21797) );
  NANDN U22338 ( .A(n21797), .B(n42095), .Z(n21757) );
  NAND U22339 ( .A(n21758), .B(n21757), .Z(n21810) );
  NANDN U22340 ( .A(n21759), .B(n42231), .Z(n21761) );
  XOR U22341 ( .A(n205), .B(a[523]), .Z(n21800) );
  NANDN U22342 ( .A(n21800), .B(n42234), .Z(n21760) );
  AND U22343 ( .A(n21761), .B(n21760), .Z(n21809) );
  XNOR U22344 ( .A(n21810), .B(n21809), .Z(n21811) );
  XNOR U22345 ( .A(n21812), .B(n21811), .Z(n21816) );
  NANDN U22346 ( .A(n21763), .B(n21762), .Z(n21767) );
  NAND U22347 ( .A(n21765), .B(n21764), .Z(n21766) );
  AND U22348 ( .A(n21767), .B(n21766), .Z(n21815) );
  XOR U22349 ( .A(n21816), .B(n21815), .Z(n21817) );
  NANDN U22350 ( .A(n21769), .B(n21768), .Z(n21773) );
  NANDN U22351 ( .A(n21771), .B(n21770), .Z(n21772) );
  NAND U22352 ( .A(n21773), .B(n21772), .Z(n21818) );
  XOR U22353 ( .A(n21817), .B(n21818), .Z(n21785) );
  OR U22354 ( .A(n21775), .B(n21774), .Z(n21779) );
  NANDN U22355 ( .A(n21777), .B(n21776), .Z(n21778) );
  NAND U22356 ( .A(n21779), .B(n21778), .Z(n21786) );
  XNOR U22357 ( .A(n21785), .B(n21786), .Z(n21787) );
  XNOR U22358 ( .A(n21788), .B(n21787), .Z(n21821) );
  XNOR U22359 ( .A(n21821), .B(sreg[1545]), .Z(n21823) );
  NAND U22360 ( .A(n21780), .B(sreg[1544]), .Z(n21784) );
  OR U22361 ( .A(n21782), .B(n21781), .Z(n21783) );
  AND U22362 ( .A(n21784), .B(n21783), .Z(n21822) );
  XOR U22363 ( .A(n21823), .B(n21822), .Z(c[1545]) );
  NANDN U22364 ( .A(n21786), .B(n21785), .Z(n21790) );
  NAND U22365 ( .A(n21788), .B(n21787), .Z(n21789) );
  NAND U22366 ( .A(n21790), .B(n21789), .Z(n21829) );
  NAND U22367 ( .A(b[0]), .B(a[530]), .Z(n21791) );
  XNOR U22368 ( .A(b[1]), .B(n21791), .Z(n21793) );
  NAND U22369 ( .A(n90), .B(a[529]), .Z(n21792) );
  AND U22370 ( .A(n21793), .B(n21792), .Z(n21846) );
  XOR U22371 ( .A(a[526]), .B(n42197), .Z(n21835) );
  NANDN U22372 ( .A(n21835), .B(n42173), .Z(n21796) );
  NANDN U22373 ( .A(n21794), .B(n42172), .Z(n21795) );
  NAND U22374 ( .A(n21796), .B(n21795), .Z(n21844) );
  NAND U22375 ( .A(b[7]), .B(a[522]), .Z(n21845) );
  XNOR U22376 ( .A(n21844), .B(n21845), .Z(n21847) );
  XOR U22377 ( .A(n21846), .B(n21847), .Z(n21853) );
  NANDN U22378 ( .A(n21797), .B(n42093), .Z(n21799) );
  XOR U22379 ( .A(n42134), .B(a[528]), .Z(n21838) );
  NANDN U22380 ( .A(n21838), .B(n42095), .Z(n21798) );
  NAND U22381 ( .A(n21799), .B(n21798), .Z(n21851) );
  NANDN U22382 ( .A(n21800), .B(n42231), .Z(n21802) );
  XOR U22383 ( .A(n205), .B(a[524]), .Z(n21841) );
  NANDN U22384 ( .A(n21841), .B(n42234), .Z(n21801) );
  AND U22385 ( .A(n21802), .B(n21801), .Z(n21850) );
  XNOR U22386 ( .A(n21851), .B(n21850), .Z(n21852) );
  XNOR U22387 ( .A(n21853), .B(n21852), .Z(n21857) );
  NANDN U22388 ( .A(n21804), .B(n21803), .Z(n21808) );
  NAND U22389 ( .A(n21806), .B(n21805), .Z(n21807) );
  AND U22390 ( .A(n21808), .B(n21807), .Z(n21856) );
  XOR U22391 ( .A(n21857), .B(n21856), .Z(n21858) );
  NANDN U22392 ( .A(n21810), .B(n21809), .Z(n21814) );
  NANDN U22393 ( .A(n21812), .B(n21811), .Z(n21813) );
  NAND U22394 ( .A(n21814), .B(n21813), .Z(n21859) );
  XOR U22395 ( .A(n21858), .B(n21859), .Z(n21826) );
  OR U22396 ( .A(n21816), .B(n21815), .Z(n21820) );
  NANDN U22397 ( .A(n21818), .B(n21817), .Z(n21819) );
  NAND U22398 ( .A(n21820), .B(n21819), .Z(n21827) );
  XNOR U22399 ( .A(n21826), .B(n21827), .Z(n21828) );
  XNOR U22400 ( .A(n21829), .B(n21828), .Z(n21862) );
  XNOR U22401 ( .A(n21862), .B(sreg[1546]), .Z(n21864) );
  NAND U22402 ( .A(n21821), .B(sreg[1545]), .Z(n21825) );
  OR U22403 ( .A(n21823), .B(n21822), .Z(n21824) );
  AND U22404 ( .A(n21825), .B(n21824), .Z(n21863) );
  XOR U22405 ( .A(n21864), .B(n21863), .Z(c[1546]) );
  NANDN U22406 ( .A(n21827), .B(n21826), .Z(n21831) );
  NAND U22407 ( .A(n21829), .B(n21828), .Z(n21830) );
  NAND U22408 ( .A(n21831), .B(n21830), .Z(n21870) );
  NAND U22409 ( .A(b[0]), .B(a[531]), .Z(n21832) );
  XNOR U22410 ( .A(b[1]), .B(n21832), .Z(n21834) );
  NAND U22411 ( .A(n90), .B(a[530]), .Z(n21833) );
  AND U22412 ( .A(n21834), .B(n21833), .Z(n21887) );
  XOR U22413 ( .A(a[527]), .B(n42197), .Z(n21876) );
  NANDN U22414 ( .A(n21876), .B(n42173), .Z(n21837) );
  NANDN U22415 ( .A(n21835), .B(n42172), .Z(n21836) );
  NAND U22416 ( .A(n21837), .B(n21836), .Z(n21885) );
  NAND U22417 ( .A(b[7]), .B(a[523]), .Z(n21886) );
  XNOR U22418 ( .A(n21885), .B(n21886), .Z(n21888) );
  XOR U22419 ( .A(n21887), .B(n21888), .Z(n21894) );
  NANDN U22420 ( .A(n21838), .B(n42093), .Z(n21840) );
  XOR U22421 ( .A(n42134), .B(a[529]), .Z(n21879) );
  NANDN U22422 ( .A(n21879), .B(n42095), .Z(n21839) );
  NAND U22423 ( .A(n21840), .B(n21839), .Z(n21892) );
  NANDN U22424 ( .A(n21841), .B(n42231), .Z(n21843) );
  XOR U22425 ( .A(n205), .B(a[525]), .Z(n21882) );
  NANDN U22426 ( .A(n21882), .B(n42234), .Z(n21842) );
  AND U22427 ( .A(n21843), .B(n21842), .Z(n21891) );
  XNOR U22428 ( .A(n21892), .B(n21891), .Z(n21893) );
  XNOR U22429 ( .A(n21894), .B(n21893), .Z(n21898) );
  NANDN U22430 ( .A(n21845), .B(n21844), .Z(n21849) );
  NAND U22431 ( .A(n21847), .B(n21846), .Z(n21848) );
  AND U22432 ( .A(n21849), .B(n21848), .Z(n21897) );
  XOR U22433 ( .A(n21898), .B(n21897), .Z(n21899) );
  NANDN U22434 ( .A(n21851), .B(n21850), .Z(n21855) );
  NANDN U22435 ( .A(n21853), .B(n21852), .Z(n21854) );
  NAND U22436 ( .A(n21855), .B(n21854), .Z(n21900) );
  XOR U22437 ( .A(n21899), .B(n21900), .Z(n21867) );
  OR U22438 ( .A(n21857), .B(n21856), .Z(n21861) );
  NANDN U22439 ( .A(n21859), .B(n21858), .Z(n21860) );
  NAND U22440 ( .A(n21861), .B(n21860), .Z(n21868) );
  XNOR U22441 ( .A(n21867), .B(n21868), .Z(n21869) );
  XNOR U22442 ( .A(n21870), .B(n21869), .Z(n21903) );
  XNOR U22443 ( .A(n21903), .B(sreg[1547]), .Z(n21905) );
  NAND U22444 ( .A(n21862), .B(sreg[1546]), .Z(n21866) );
  OR U22445 ( .A(n21864), .B(n21863), .Z(n21865) );
  AND U22446 ( .A(n21866), .B(n21865), .Z(n21904) );
  XOR U22447 ( .A(n21905), .B(n21904), .Z(c[1547]) );
  NANDN U22448 ( .A(n21868), .B(n21867), .Z(n21872) );
  NAND U22449 ( .A(n21870), .B(n21869), .Z(n21871) );
  NAND U22450 ( .A(n21872), .B(n21871), .Z(n21911) );
  NAND U22451 ( .A(b[0]), .B(a[532]), .Z(n21873) );
  XNOR U22452 ( .A(b[1]), .B(n21873), .Z(n21875) );
  NAND U22453 ( .A(n91), .B(a[531]), .Z(n21874) );
  AND U22454 ( .A(n21875), .B(n21874), .Z(n21928) );
  XOR U22455 ( .A(a[528]), .B(n42197), .Z(n21917) );
  NANDN U22456 ( .A(n21917), .B(n42173), .Z(n21878) );
  NANDN U22457 ( .A(n21876), .B(n42172), .Z(n21877) );
  NAND U22458 ( .A(n21878), .B(n21877), .Z(n21926) );
  NAND U22459 ( .A(b[7]), .B(a[524]), .Z(n21927) );
  XNOR U22460 ( .A(n21926), .B(n21927), .Z(n21929) );
  XOR U22461 ( .A(n21928), .B(n21929), .Z(n21935) );
  NANDN U22462 ( .A(n21879), .B(n42093), .Z(n21881) );
  XOR U22463 ( .A(n42134), .B(a[530]), .Z(n21920) );
  NANDN U22464 ( .A(n21920), .B(n42095), .Z(n21880) );
  NAND U22465 ( .A(n21881), .B(n21880), .Z(n21933) );
  NANDN U22466 ( .A(n21882), .B(n42231), .Z(n21884) );
  XOR U22467 ( .A(n205), .B(a[526]), .Z(n21923) );
  NANDN U22468 ( .A(n21923), .B(n42234), .Z(n21883) );
  AND U22469 ( .A(n21884), .B(n21883), .Z(n21932) );
  XNOR U22470 ( .A(n21933), .B(n21932), .Z(n21934) );
  XNOR U22471 ( .A(n21935), .B(n21934), .Z(n21939) );
  NANDN U22472 ( .A(n21886), .B(n21885), .Z(n21890) );
  NAND U22473 ( .A(n21888), .B(n21887), .Z(n21889) );
  AND U22474 ( .A(n21890), .B(n21889), .Z(n21938) );
  XOR U22475 ( .A(n21939), .B(n21938), .Z(n21940) );
  NANDN U22476 ( .A(n21892), .B(n21891), .Z(n21896) );
  NANDN U22477 ( .A(n21894), .B(n21893), .Z(n21895) );
  NAND U22478 ( .A(n21896), .B(n21895), .Z(n21941) );
  XOR U22479 ( .A(n21940), .B(n21941), .Z(n21908) );
  OR U22480 ( .A(n21898), .B(n21897), .Z(n21902) );
  NANDN U22481 ( .A(n21900), .B(n21899), .Z(n21901) );
  NAND U22482 ( .A(n21902), .B(n21901), .Z(n21909) );
  XNOR U22483 ( .A(n21908), .B(n21909), .Z(n21910) );
  XNOR U22484 ( .A(n21911), .B(n21910), .Z(n21944) );
  XNOR U22485 ( .A(n21944), .B(sreg[1548]), .Z(n21946) );
  NAND U22486 ( .A(n21903), .B(sreg[1547]), .Z(n21907) );
  OR U22487 ( .A(n21905), .B(n21904), .Z(n21906) );
  AND U22488 ( .A(n21907), .B(n21906), .Z(n21945) );
  XOR U22489 ( .A(n21946), .B(n21945), .Z(c[1548]) );
  NANDN U22490 ( .A(n21909), .B(n21908), .Z(n21913) );
  NAND U22491 ( .A(n21911), .B(n21910), .Z(n21912) );
  NAND U22492 ( .A(n21913), .B(n21912), .Z(n21952) );
  NAND U22493 ( .A(b[0]), .B(a[533]), .Z(n21914) );
  XNOR U22494 ( .A(b[1]), .B(n21914), .Z(n21916) );
  NAND U22495 ( .A(n91), .B(a[532]), .Z(n21915) );
  AND U22496 ( .A(n21916), .B(n21915), .Z(n21969) );
  XOR U22497 ( .A(a[529]), .B(n42197), .Z(n21958) );
  NANDN U22498 ( .A(n21958), .B(n42173), .Z(n21919) );
  NANDN U22499 ( .A(n21917), .B(n42172), .Z(n21918) );
  NAND U22500 ( .A(n21919), .B(n21918), .Z(n21967) );
  NAND U22501 ( .A(b[7]), .B(a[525]), .Z(n21968) );
  XNOR U22502 ( .A(n21967), .B(n21968), .Z(n21970) );
  XOR U22503 ( .A(n21969), .B(n21970), .Z(n21976) );
  NANDN U22504 ( .A(n21920), .B(n42093), .Z(n21922) );
  XOR U22505 ( .A(n42134), .B(a[531]), .Z(n21961) );
  NANDN U22506 ( .A(n21961), .B(n42095), .Z(n21921) );
  NAND U22507 ( .A(n21922), .B(n21921), .Z(n21974) );
  NANDN U22508 ( .A(n21923), .B(n42231), .Z(n21925) );
  XOR U22509 ( .A(n206), .B(a[527]), .Z(n21964) );
  NANDN U22510 ( .A(n21964), .B(n42234), .Z(n21924) );
  AND U22511 ( .A(n21925), .B(n21924), .Z(n21973) );
  XNOR U22512 ( .A(n21974), .B(n21973), .Z(n21975) );
  XNOR U22513 ( .A(n21976), .B(n21975), .Z(n21980) );
  NANDN U22514 ( .A(n21927), .B(n21926), .Z(n21931) );
  NAND U22515 ( .A(n21929), .B(n21928), .Z(n21930) );
  AND U22516 ( .A(n21931), .B(n21930), .Z(n21979) );
  XOR U22517 ( .A(n21980), .B(n21979), .Z(n21981) );
  NANDN U22518 ( .A(n21933), .B(n21932), .Z(n21937) );
  NANDN U22519 ( .A(n21935), .B(n21934), .Z(n21936) );
  NAND U22520 ( .A(n21937), .B(n21936), .Z(n21982) );
  XOR U22521 ( .A(n21981), .B(n21982), .Z(n21949) );
  OR U22522 ( .A(n21939), .B(n21938), .Z(n21943) );
  NANDN U22523 ( .A(n21941), .B(n21940), .Z(n21942) );
  NAND U22524 ( .A(n21943), .B(n21942), .Z(n21950) );
  XNOR U22525 ( .A(n21949), .B(n21950), .Z(n21951) );
  XNOR U22526 ( .A(n21952), .B(n21951), .Z(n21985) );
  XNOR U22527 ( .A(n21985), .B(sreg[1549]), .Z(n21987) );
  NAND U22528 ( .A(n21944), .B(sreg[1548]), .Z(n21948) );
  OR U22529 ( .A(n21946), .B(n21945), .Z(n21947) );
  AND U22530 ( .A(n21948), .B(n21947), .Z(n21986) );
  XOR U22531 ( .A(n21987), .B(n21986), .Z(c[1549]) );
  NANDN U22532 ( .A(n21950), .B(n21949), .Z(n21954) );
  NAND U22533 ( .A(n21952), .B(n21951), .Z(n21953) );
  NAND U22534 ( .A(n21954), .B(n21953), .Z(n21993) );
  NAND U22535 ( .A(b[0]), .B(a[534]), .Z(n21955) );
  XNOR U22536 ( .A(b[1]), .B(n21955), .Z(n21957) );
  NAND U22537 ( .A(n91), .B(a[533]), .Z(n21956) );
  AND U22538 ( .A(n21957), .B(n21956), .Z(n22010) );
  XOR U22539 ( .A(a[530]), .B(n42197), .Z(n21999) );
  NANDN U22540 ( .A(n21999), .B(n42173), .Z(n21960) );
  NANDN U22541 ( .A(n21958), .B(n42172), .Z(n21959) );
  NAND U22542 ( .A(n21960), .B(n21959), .Z(n22008) );
  NAND U22543 ( .A(b[7]), .B(a[526]), .Z(n22009) );
  XNOR U22544 ( .A(n22008), .B(n22009), .Z(n22011) );
  XOR U22545 ( .A(n22010), .B(n22011), .Z(n22017) );
  NANDN U22546 ( .A(n21961), .B(n42093), .Z(n21963) );
  XOR U22547 ( .A(n42134), .B(a[532]), .Z(n22002) );
  NANDN U22548 ( .A(n22002), .B(n42095), .Z(n21962) );
  NAND U22549 ( .A(n21963), .B(n21962), .Z(n22015) );
  NANDN U22550 ( .A(n21964), .B(n42231), .Z(n21966) );
  XOR U22551 ( .A(n206), .B(a[528]), .Z(n22005) );
  NANDN U22552 ( .A(n22005), .B(n42234), .Z(n21965) );
  AND U22553 ( .A(n21966), .B(n21965), .Z(n22014) );
  XNOR U22554 ( .A(n22015), .B(n22014), .Z(n22016) );
  XNOR U22555 ( .A(n22017), .B(n22016), .Z(n22021) );
  NANDN U22556 ( .A(n21968), .B(n21967), .Z(n21972) );
  NAND U22557 ( .A(n21970), .B(n21969), .Z(n21971) );
  AND U22558 ( .A(n21972), .B(n21971), .Z(n22020) );
  XOR U22559 ( .A(n22021), .B(n22020), .Z(n22022) );
  NANDN U22560 ( .A(n21974), .B(n21973), .Z(n21978) );
  NANDN U22561 ( .A(n21976), .B(n21975), .Z(n21977) );
  NAND U22562 ( .A(n21978), .B(n21977), .Z(n22023) );
  XOR U22563 ( .A(n22022), .B(n22023), .Z(n21990) );
  OR U22564 ( .A(n21980), .B(n21979), .Z(n21984) );
  NANDN U22565 ( .A(n21982), .B(n21981), .Z(n21983) );
  NAND U22566 ( .A(n21984), .B(n21983), .Z(n21991) );
  XNOR U22567 ( .A(n21990), .B(n21991), .Z(n21992) );
  XNOR U22568 ( .A(n21993), .B(n21992), .Z(n22026) );
  XNOR U22569 ( .A(n22026), .B(sreg[1550]), .Z(n22028) );
  NAND U22570 ( .A(n21985), .B(sreg[1549]), .Z(n21989) );
  OR U22571 ( .A(n21987), .B(n21986), .Z(n21988) );
  AND U22572 ( .A(n21989), .B(n21988), .Z(n22027) );
  XOR U22573 ( .A(n22028), .B(n22027), .Z(c[1550]) );
  NANDN U22574 ( .A(n21991), .B(n21990), .Z(n21995) );
  NAND U22575 ( .A(n21993), .B(n21992), .Z(n21994) );
  NAND U22576 ( .A(n21995), .B(n21994), .Z(n22034) );
  NAND U22577 ( .A(b[0]), .B(a[535]), .Z(n21996) );
  XNOR U22578 ( .A(b[1]), .B(n21996), .Z(n21998) );
  NAND U22579 ( .A(n91), .B(a[534]), .Z(n21997) );
  AND U22580 ( .A(n21998), .B(n21997), .Z(n22051) );
  XOR U22581 ( .A(a[531]), .B(n42197), .Z(n22040) );
  NANDN U22582 ( .A(n22040), .B(n42173), .Z(n22001) );
  NANDN U22583 ( .A(n21999), .B(n42172), .Z(n22000) );
  NAND U22584 ( .A(n22001), .B(n22000), .Z(n22049) );
  NAND U22585 ( .A(b[7]), .B(a[527]), .Z(n22050) );
  XNOR U22586 ( .A(n22049), .B(n22050), .Z(n22052) );
  XOR U22587 ( .A(n22051), .B(n22052), .Z(n22058) );
  NANDN U22588 ( .A(n22002), .B(n42093), .Z(n22004) );
  XOR U22589 ( .A(n42134), .B(a[533]), .Z(n22043) );
  NANDN U22590 ( .A(n22043), .B(n42095), .Z(n22003) );
  NAND U22591 ( .A(n22004), .B(n22003), .Z(n22056) );
  NANDN U22592 ( .A(n22005), .B(n42231), .Z(n22007) );
  XOR U22593 ( .A(n206), .B(a[529]), .Z(n22046) );
  NANDN U22594 ( .A(n22046), .B(n42234), .Z(n22006) );
  AND U22595 ( .A(n22007), .B(n22006), .Z(n22055) );
  XNOR U22596 ( .A(n22056), .B(n22055), .Z(n22057) );
  XNOR U22597 ( .A(n22058), .B(n22057), .Z(n22062) );
  NANDN U22598 ( .A(n22009), .B(n22008), .Z(n22013) );
  NAND U22599 ( .A(n22011), .B(n22010), .Z(n22012) );
  AND U22600 ( .A(n22013), .B(n22012), .Z(n22061) );
  XOR U22601 ( .A(n22062), .B(n22061), .Z(n22063) );
  NANDN U22602 ( .A(n22015), .B(n22014), .Z(n22019) );
  NANDN U22603 ( .A(n22017), .B(n22016), .Z(n22018) );
  NAND U22604 ( .A(n22019), .B(n22018), .Z(n22064) );
  XOR U22605 ( .A(n22063), .B(n22064), .Z(n22031) );
  OR U22606 ( .A(n22021), .B(n22020), .Z(n22025) );
  NANDN U22607 ( .A(n22023), .B(n22022), .Z(n22024) );
  NAND U22608 ( .A(n22025), .B(n22024), .Z(n22032) );
  XNOR U22609 ( .A(n22031), .B(n22032), .Z(n22033) );
  XNOR U22610 ( .A(n22034), .B(n22033), .Z(n22067) );
  XNOR U22611 ( .A(n22067), .B(sreg[1551]), .Z(n22069) );
  NAND U22612 ( .A(n22026), .B(sreg[1550]), .Z(n22030) );
  OR U22613 ( .A(n22028), .B(n22027), .Z(n22029) );
  AND U22614 ( .A(n22030), .B(n22029), .Z(n22068) );
  XOR U22615 ( .A(n22069), .B(n22068), .Z(c[1551]) );
  NANDN U22616 ( .A(n22032), .B(n22031), .Z(n22036) );
  NAND U22617 ( .A(n22034), .B(n22033), .Z(n22035) );
  NAND U22618 ( .A(n22036), .B(n22035), .Z(n22075) );
  NAND U22619 ( .A(b[0]), .B(a[536]), .Z(n22037) );
  XNOR U22620 ( .A(b[1]), .B(n22037), .Z(n22039) );
  NAND U22621 ( .A(n91), .B(a[535]), .Z(n22038) );
  AND U22622 ( .A(n22039), .B(n22038), .Z(n22092) );
  XOR U22623 ( .A(a[532]), .B(n42197), .Z(n22081) );
  NANDN U22624 ( .A(n22081), .B(n42173), .Z(n22042) );
  NANDN U22625 ( .A(n22040), .B(n42172), .Z(n22041) );
  NAND U22626 ( .A(n22042), .B(n22041), .Z(n22090) );
  NAND U22627 ( .A(b[7]), .B(a[528]), .Z(n22091) );
  XNOR U22628 ( .A(n22090), .B(n22091), .Z(n22093) );
  XOR U22629 ( .A(n22092), .B(n22093), .Z(n22099) );
  NANDN U22630 ( .A(n22043), .B(n42093), .Z(n22045) );
  XOR U22631 ( .A(n42134), .B(a[534]), .Z(n22084) );
  NANDN U22632 ( .A(n22084), .B(n42095), .Z(n22044) );
  NAND U22633 ( .A(n22045), .B(n22044), .Z(n22097) );
  NANDN U22634 ( .A(n22046), .B(n42231), .Z(n22048) );
  XOR U22635 ( .A(n206), .B(a[530]), .Z(n22087) );
  NANDN U22636 ( .A(n22087), .B(n42234), .Z(n22047) );
  AND U22637 ( .A(n22048), .B(n22047), .Z(n22096) );
  XNOR U22638 ( .A(n22097), .B(n22096), .Z(n22098) );
  XNOR U22639 ( .A(n22099), .B(n22098), .Z(n22103) );
  NANDN U22640 ( .A(n22050), .B(n22049), .Z(n22054) );
  NAND U22641 ( .A(n22052), .B(n22051), .Z(n22053) );
  AND U22642 ( .A(n22054), .B(n22053), .Z(n22102) );
  XOR U22643 ( .A(n22103), .B(n22102), .Z(n22104) );
  NANDN U22644 ( .A(n22056), .B(n22055), .Z(n22060) );
  NANDN U22645 ( .A(n22058), .B(n22057), .Z(n22059) );
  NAND U22646 ( .A(n22060), .B(n22059), .Z(n22105) );
  XOR U22647 ( .A(n22104), .B(n22105), .Z(n22072) );
  OR U22648 ( .A(n22062), .B(n22061), .Z(n22066) );
  NANDN U22649 ( .A(n22064), .B(n22063), .Z(n22065) );
  NAND U22650 ( .A(n22066), .B(n22065), .Z(n22073) );
  XNOR U22651 ( .A(n22072), .B(n22073), .Z(n22074) );
  XNOR U22652 ( .A(n22075), .B(n22074), .Z(n22108) );
  XNOR U22653 ( .A(n22108), .B(sreg[1552]), .Z(n22110) );
  NAND U22654 ( .A(n22067), .B(sreg[1551]), .Z(n22071) );
  OR U22655 ( .A(n22069), .B(n22068), .Z(n22070) );
  AND U22656 ( .A(n22071), .B(n22070), .Z(n22109) );
  XOR U22657 ( .A(n22110), .B(n22109), .Z(c[1552]) );
  NANDN U22658 ( .A(n22073), .B(n22072), .Z(n22077) );
  NAND U22659 ( .A(n22075), .B(n22074), .Z(n22076) );
  NAND U22660 ( .A(n22077), .B(n22076), .Z(n22116) );
  NAND U22661 ( .A(b[0]), .B(a[537]), .Z(n22078) );
  XNOR U22662 ( .A(b[1]), .B(n22078), .Z(n22080) );
  NAND U22663 ( .A(n91), .B(a[536]), .Z(n22079) );
  AND U22664 ( .A(n22080), .B(n22079), .Z(n22133) );
  XOR U22665 ( .A(a[533]), .B(n42197), .Z(n22122) );
  NANDN U22666 ( .A(n22122), .B(n42173), .Z(n22083) );
  NANDN U22667 ( .A(n22081), .B(n42172), .Z(n22082) );
  NAND U22668 ( .A(n22083), .B(n22082), .Z(n22131) );
  NAND U22669 ( .A(b[7]), .B(a[529]), .Z(n22132) );
  XNOR U22670 ( .A(n22131), .B(n22132), .Z(n22134) );
  XOR U22671 ( .A(n22133), .B(n22134), .Z(n22140) );
  NANDN U22672 ( .A(n22084), .B(n42093), .Z(n22086) );
  XOR U22673 ( .A(n42134), .B(a[535]), .Z(n22125) );
  NANDN U22674 ( .A(n22125), .B(n42095), .Z(n22085) );
  NAND U22675 ( .A(n22086), .B(n22085), .Z(n22138) );
  NANDN U22676 ( .A(n22087), .B(n42231), .Z(n22089) );
  XOR U22677 ( .A(n206), .B(a[531]), .Z(n22128) );
  NANDN U22678 ( .A(n22128), .B(n42234), .Z(n22088) );
  AND U22679 ( .A(n22089), .B(n22088), .Z(n22137) );
  XNOR U22680 ( .A(n22138), .B(n22137), .Z(n22139) );
  XNOR U22681 ( .A(n22140), .B(n22139), .Z(n22144) );
  NANDN U22682 ( .A(n22091), .B(n22090), .Z(n22095) );
  NAND U22683 ( .A(n22093), .B(n22092), .Z(n22094) );
  AND U22684 ( .A(n22095), .B(n22094), .Z(n22143) );
  XOR U22685 ( .A(n22144), .B(n22143), .Z(n22145) );
  NANDN U22686 ( .A(n22097), .B(n22096), .Z(n22101) );
  NANDN U22687 ( .A(n22099), .B(n22098), .Z(n22100) );
  NAND U22688 ( .A(n22101), .B(n22100), .Z(n22146) );
  XOR U22689 ( .A(n22145), .B(n22146), .Z(n22113) );
  OR U22690 ( .A(n22103), .B(n22102), .Z(n22107) );
  NANDN U22691 ( .A(n22105), .B(n22104), .Z(n22106) );
  NAND U22692 ( .A(n22107), .B(n22106), .Z(n22114) );
  XNOR U22693 ( .A(n22113), .B(n22114), .Z(n22115) );
  XNOR U22694 ( .A(n22116), .B(n22115), .Z(n22149) );
  XNOR U22695 ( .A(n22149), .B(sreg[1553]), .Z(n22151) );
  NAND U22696 ( .A(n22108), .B(sreg[1552]), .Z(n22112) );
  OR U22697 ( .A(n22110), .B(n22109), .Z(n22111) );
  AND U22698 ( .A(n22112), .B(n22111), .Z(n22150) );
  XOR U22699 ( .A(n22151), .B(n22150), .Z(c[1553]) );
  NANDN U22700 ( .A(n22114), .B(n22113), .Z(n22118) );
  NAND U22701 ( .A(n22116), .B(n22115), .Z(n22117) );
  NAND U22702 ( .A(n22118), .B(n22117), .Z(n22157) );
  NAND U22703 ( .A(b[0]), .B(a[538]), .Z(n22119) );
  XNOR U22704 ( .A(b[1]), .B(n22119), .Z(n22121) );
  NAND U22705 ( .A(n91), .B(a[537]), .Z(n22120) );
  AND U22706 ( .A(n22121), .B(n22120), .Z(n22174) );
  XOR U22707 ( .A(a[534]), .B(n42197), .Z(n22163) );
  NANDN U22708 ( .A(n22163), .B(n42173), .Z(n22124) );
  NANDN U22709 ( .A(n22122), .B(n42172), .Z(n22123) );
  NAND U22710 ( .A(n22124), .B(n22123), .Z(n22172) );
  NAND U22711 ( .A(b[7]), .B(a[530]), .Z(n22173) );
  XNOR U22712 ( .A(n22172), .B(n22173), .Z(n22175) );
  XOR U22713 ( .A(n22174), .B(n22175), .Z(n22181) );
  NANDN U22714 ( .A(n22125), .B(n42093), .Z(n22127) );
  XOR U22715 ( .A(n42134), .B(a[536]), .Z(n22166) );
  NANDN U22716 ( .A(n22166), .B(n42095), .Z(n22126) );
  NAND U22717 ( .A(n22127), .B(n22126), .Z(n22179) );
  NANDN U22718 ( .A(n22128), .B(n42231), .Z(n22130) );
  XOR U22719 ( .A(n206), .B(a[532]), .Z(n22169) );
  NANDN U22720 ( .A(n22169), .B(n42234), .Z(n22129) );
  AND U22721 ( .A(n22130), .B(n22129), .Z(n22178) );
  XNOR U22722 ( .A(n22179), .B(n22178), .Z(n22180) );
  XNOR U22723 ( .A(n22181), .B(n22180), .Z(n22185) );
  NANDN U22724 ( .A(n22132), .B(n22131), .Z(n22136) );
  NAND U22725 ( .A(n22134), .B(n22133), .Z(n22135) );
  AND U22726 ( .A(n22136), .B(n22135), .Z(n22184) );
  XOR U22727 ( .A(n22185), .B(n22184), .Z(n22186) );
  NANDN U22728 ( .A(n22138), .B(n22137), .Z(n22142) );
  NANDN U22729 ( .A(n22140), .B(n22139), .Z(n22141) );
  NAND U22730 ( .A(n22142), .B(n22141), .Z(n22187) );
  XOR U22731 ( .A(n22186), .B(n22187), .Z(n22154) );
  OR U22732 ( .A(n22144), .B(n22143), .Z(n22148) );
  NANDN U22733 ( .A(n22146), .B(n22145), .Z(n22147) );
  NAND U22734 ( .A(n22148), .B(n22147), .Z(n22155) );
  XNOR U22735 ( .A(n22154), .B(n22155), .Z(n22156) );
  XNOR U22736 ( .A(n22157), .B(n22156), .Z(n22190) );
  XNOR U22737 ( .A(n22190), .B(sreg[1554]), .Z(n22192) );
  NAND U22738 ( .A(n22149), .B(sreg[1553]), .Z(n22153) );
  OR U22739 ( .A(n22151), .B(n22150), .Z(n22152) );
  AND U22740 ( .A(n22153), .B(n22152), .Z(n22191) );
  XOR U22741 ( .A(n22192), .B(n22191), .Z(c[1554]) );
  NANDN U22742 ( .A(n22155), .B(n22154), .Z(n22159) );
  NAND U22743 ( .A(n22157), .B(n22156), .Z(n22158) );
  NAND U22744 ( .A(n22159), .B(n22158), .Z(n22198) );
  NAND U22745 ( .A(b[0]), .B(a[539]), .Z(n22160) );
  XNOR U22746 ( .A(b[1]), .B(n22160), .Z(n22162) );
  NAND U22747 ( .A(n92), .B(a[538]), .Z(n22161) );
  AND U22748 ( .A(n22162), .B(n22161), .Z(n22215) );
  XOR U22749 ( .A(a[535]), .B(n42197), .Z(n22204) );
  NANDN U22750 ( .A(n22204), .B(n42173), .Z(n22165) );
  NANDN U22751 ( .A(n22163), .B(n42172), .Z(n22164) );
  NAND U22752 ( .A(n22165), .B(n22164), .Z(n22213) );
  NAND U22753 ( .A(b[7]), .B(a[531]), .Z(n22214) );
  XNOR U22754 ( .A(n22213), .B(n22214), .Z(n22216) );
  XOR U22755 ( .A(n22215), .B(n22216), .Z(n22222) );
  NANDN U22756 ( .A(n22166), .B(n42093), .Z(n22168) );
  XOR U22757 ( .A(n42134), .B(a[537]), .Z(n22207) );
  NANDN U22758 ( .A(n22207), .B(n42095), .Z(n22167) );
  NAND U22759 ( .A(n22168), .B(n22167), .Z(n22220) );
  NANDN U22760 ( .A(n22169), .B(n42231), .Z(n22171) );
  XOR U22761 ( .A(n206), .B(a[533]), .Z(n22210) );
  NANDN U22762 ( .A(n22210), .B(n42234), .Z(n22170) );
  AND U22763 ( .A(n22171), .B(n22170), .Z(n22219) );
  XNOR U22764 ( .A(n22220), .B(n22219), .Z(n22221) );
  XNOR U22765 ( .A(n22222), .B(n22221), .Z(n22226) );
  NANDN U22766 ( .A(n22173), .B(n22172), .Z(n22177) );
  NAND U22767 ( .A(n22175), .B(n22174), .Z(n22176) );
  AND U22768 ( .A(n22177), .B(n22176), .Z(n22225) );
  XOR U22769 ( .A(n22226), .B(n22225), .Z(n22227) );
  NANDN U22770 ( .A(n22179), .B(n22178), .Z(n22183) );
  NANDN U22771 ( .A(n22181), .B(n22180), .Z(n22182) );
  NAND U22772 ( .A(n22183), .B(n22182), .Z(n22228) );
  XOR U22773 ( .A(n22227), .B(n22228), .Z(n22195) );
  OR U22774 ( .A(n22185), .B(n22184), .Z(n22189) );
  NANDN U22775 ( .A(n22187), .B(n22186), .Z(n22188) );
  NAND U22776 ( .A(n22189), .B(n22188), .Z(n22196) );
  XNOR U22777 ( .A(n22195), .B(n22196), .Z(n22197) );
  XNOR U22778 ( .A(n22198), .B(n22197), .Z(n22231) );
  XNOR U22779 ( .A(n22231), .B(sreg[1555]), .Z(n22233) );
  NAND U22780 ( .A(n22190), .B(sreg[1554]), .Z(n22194) );
  OR U22781 ( .A(n22192), .B(n22191), .Z(n22193) );
  AND U22782 ( .A(n22194), .B(n22193), .Z(n22232) );
  XOR U22783 ( .A(n22233), .B(n22232), .Z(c[1555]) );
  NANDN U22784 ( .A(n22196), .B(n22195), .Z(n22200) );
  NAND U22785 ( .A(n22198), .B(n22197), .Z(n22199) );
  NAND U22786 ( .A(n22200), .B(n22199), .Z(n22239) );
  NAND U22787 ( .A(b[0]), .B(a[540]), .Z(n22201) );
  XNOR U22788 ( .A(b[1]), .B(n22201), .Z(n22203) );
  NAND U22789 ( .A(n92), .B(a[539]), .Z(n22202) );
  AND U22790 ( .A(n22203), .B(n22202), .Z(n22256) );
  XOR U22791 ( .A(a[536]), .B(n42197), .Z(n22245) );
  NANDN U22792 ( .A(n22245), .B(n42173), .Z(n22206) );
  NANDN U22793 ( .A(n22204), .B(n42172), .Z(n22205) );
  NAND U22794 ( .A(n22206), .B(n22205), .Z(n22254) );
  NAND U22795 ( .A(b[7]), .B(a[532]), .Z(n22255) );
  XNOR U22796 ( .A(n22254), .B(n22255), .Z(n22257) );
  XOR U22797 ( .A(n22256), .B(n22257), .Z(n22263) );
  NANDN U22798 ( .A(n22207), .B(n42093), .Z(n22209) );
  XOR U22799 ( .A(n42134), .B(a[538]), .Z(n22248) );
  NANDN U22800 ( .A(n22248), .B(n42095), .Z(n22208) );
  NAND U22801 ( .A(n22209), .B(n22208), .Z(n22261) );
  NANDN U22802 ( .A(n22210), .B(n42231), .Z(n22212) );
  XOR U22803 ( .A(n206), .B(a[534]), .Z(n22251) );
  NANDN U22804 ( .A(n22251), .B(n42234), .Z(n22211) );
  AND U22805 ( .A(n22212), .B(n22211), .Z(n22260) );
  XNOR U22806 ( .A(n22261), .B(n22260), .Z(n22262) );
  XNOR U22807 ( .A(n22263), .B(n22262), .Z(n22267) );
  NANDN U22808 ( .A(n22214), .B(n22213), .Z(n22218) );
  NAND U22809 ( .A(n22216), .B(n22215), .Z(n22217) );
  AND U22810 ( .A(n22218), .B(n22217), .Z(n22266) );
  XOR U22811 ( .A(n22267), .B(n22266), .Z(n22268) );
  NANDN U22812 ( .A(n22220), .B(n22219), .Z(n22224) );
  NANDN U22813 ( .A(n22222), .B(n22221), .Z(n22223) );
  NAND U22814 ( .A(n22224), .B(n22223), .Z(n22269) );
  XOR U22815 ( .A(n22268), .B(n22269), .Z(n22236) );
  OR U22816 ( .A(n22226), .B(n22225), .Z(n22230) );
  NANDN U22817 ( .A(n22228), .B(n22227), .Z(n22229) );
  NAND U22818 ( .A(n22230), .B(n22229), .Z(n22237) );
  XNOR U22819 ( .A(n22236), .B(n22237), .Z(n22238) );
  XNOR U22820 ( .A(n22239), .B(n22238), .Z(n22272) );
  XNOR U22821 ( .A(n22272), .B(sreg[1556]), .Z(n22274) );
  NAND U22822 ( .A(n22231), .B(sreg[1555]), .Z(n22235) );
  OR U22823 ( .A(n22233), .B(n22232), .Z(n22234) );
  AND U22824 ( .A(n22235), .B(n22234), .Z(n22273) );
  XOR U22825 ( .A(n22274), .B(n22273), .Z(c[1556]) );
  NANDN U22826 ( .A(n22237), .B(n22236), .Z(n22241) );
  NAND U22827 ( .A(n22239), .B(n22238), .Z(n22240) );
  NAND U22828 ( .A(n22241), .B(n22240), .Z(n22280) );
  NAND U22829 ( .A(b[0]), .B(a[541]), .Z(n22242) );
  XNOR U22830 ( .A(b[1]), .B(n22242), .Z(n22244) );
  NAND U22831 ( .A(n92), .B(a[540]), .Z(n22243) );
  AND U22832 ( .A(n22244), .B(n22243), .Z(n22297) );
  XOR U22833 ( .A(a[537]), .B(n42197), .Z(n22286) );
  NANDN U22834 ( .A(n22286), .B(n42173), .Z(n22247) );
  NANDN U22835 ( .A(n22245), .B(n42172), .Z(n22246) );
  NAND U22836 ( .A(n22247), .B(n22246), .Z(n22295) );
  NAND U22837 ( .A(b[7]), .B(a[533]), .Z(n22296) );
  XNOR U22838 ( .A(n22295), .B(n22296), .Z(n22298) );
  XOR U22839 ( .A(n22297), .B(n22298), .Z(n22304) );
  NANDN U22840 ( .A(n22248), .B(n42093), .Z(n22250) );
  XOR U22841 ( .A(n42134), .B(a[539]), .Z(n22289) );
  NANDN U22842 ( .A(n22289), .B(n42095), .Z(n22249) );
  NAND U22843 ( .A(n22250), .B(n22249), .Z(n22302) );
  NANDN U22844 ( .A(n22251), .B(n42231), .Z(n22253) );
  XOR U22845 ( .A(n206), .B(a[535]), .Z(n22292) );
  NANDN U22846 ( .A(n22292), .B(n42234), .Z(n22252) );
  AND U22847 ( .A(n22253), .B(n22252), .Z(n22301) );
  XNOR U22848 ( .A(n22302), .B(n22301), .Z(n22303) );
  XNOR U22849 ( .A(n22304), .B(n22303), .Z(n22308) );
  NANDN U22850 ( .A(n22255), .B(n22254), .Z(n22259) );
  NAND U22851 ( .A(n22257), .B(n22256), .Z(n22258) );
  AND U22852 ( .A(n22259), .B(n22258), .Z(n22307) );
  XOR U22853 ( .A(n22308), .B(n22307), .Z(n22309) );
  NANDN U22854 ( .A(n22261), .B(n22260), .Z(n22265) );
  NANDN U22855 ( .A(n22263), .B(n22262), .Z(n22264) );
  NAND U22856 ( .A(n22265), .B(n22264), .Z(n22310) );
  XOR U22857 ( .A(n22309), .B(n22310), .Z(n22277) );
  OR U22858 ( .A(n22267), .B(n22266), .Z(n22271) );
  NANDN U22859 ( .A(n22269), .B(n22268), .Z(n22270) );
  NAND U22860 ( .A(n22271), .B(n22270), .Z(n22278) );
  XNOR U22861 ( .A(n22277), .B(n22278), .Z(n22279) );
  XNOR U22862 ( .A(n22280), .B(n22279), .Z(n22313) );
  XNOR U22863 ( .A(n22313), .B(sreg[1557]), .Z(n22315) );
  NAND U22864 ( .A(n22272), .B(sreg[1556]), .Z(n22276) );
  OR U22865 ( .A(n22274), .B(n22273), .Z(n22275) );
  AND U22866 ( .A(n22276), .B(n22275), .Z(n22314) );
  XOR U22867 ( .A(n22315), .B(n22314), .Z(c[1557]) );
  NANDN U22868 ( .A(n22278), .B(n22277), .Z(n22282) );
  NAND U22869 ( .A(n22280), .B(n22279), .Z(n22281) );
  NAND U22870 ( .A(n22282), .B(n22281), .Z(n22321) );
  NAND U22871 ( .A(b[0]), .B(a[542]), .Z(n22283) );
  XNOR U22872 ( .A(b[1]), .B(n22283), .Z(n22285) );
  NAND U22873 ( .A(n92), .B(a[541]), .Z(n22284) );
  AND U22874 ( .A(n22285), .B(n22284), .Z(n22338) );
  XOR U22875 ( .A(a[538]), .B(n42197), .Z(n22327) );
  NANDN U22876 ( .A(n22327), .B(n42173), .Z(n22288) );
  NANDN U22877 ( .A(n22286), .B(n42172), .Z(n22287) );
  NAND U22878 ( .A(n22288), .B(n22287), .Z(n22336) );
  NAND U22879 ( .A(b[7]), .B(a[534]), .Z(n22337) );
  XNOR U22880 ( .A(n22336), .B(n22337), .Z(n22339) );
  XOR U22881 ( .A(n22338), .B(n22339), .Z(n22345) );
  NANDN U22882 ( .A(n22289), .B(n42093), .Z(n22291) );
  XOR U22883 ( .A(n42134), .B(a[540]), .Z(n22330) );
  NANDN U22884 ( .A(n22330), .B(n42095), .Z(n22290) );
  NAND U22885 ( .A(n22291), .B(n22290), .Z(n22343) );
  NANDN U22886 ( .A(n22292), .B(n42231), .Z(n22294) );
  XOR U22887 ( .A(n206), .B(a[536]), .Z(n22333) );
  NANDN U22888 ( .A(n22333), .B(n42234), .Z(n22293) );
  AND U22889 ( .A(n22294), .B(n22293), .Z(n22342) );
  XNOR U22890 ( .A(n22343), .B(n22342), .Z(n22344) );
  XNOR U22891 ( .A(n22345), .B(n22344), .Z(n22349) );
  NANDN U22892 ( .A(n22296), .B(n22295), .Z(n22300) );
  NAND U22893 ( .A(n22298), .B(n22297), .Z(n22299) );
  AND U22894 ( .A(n22300), .B(n22299), .Z(n22348) );
  XOR U22895 ( .A(n22349), .B(n22348), .Z(n22350) );
  NANDN U22896 ( .A(n22302), .B(n22301), .Z(n22306) );
  NANDN U22897 ( .A(n22304), .B(n22303), .Z(n22305) );
  NAND U22898 ( .A(n22306), .B(n22305), .Z(n22351) );
  XOR U22899 ( .A(n22350), .B(n22351), .Z(n22318) );
  OR U22900 ( .A(n22308), .B(n22307), .Z(n22312) );
  NANDN U22901 ( .A(n22310), .B(n22309), .Z(n22311) );
  NAND U22902 ( .A(n22312), .B(n22311), .Z(n22319) );
  XNOR U22903 ( .A(n22318), .B(n22319), .Z(n22320) );
  XNOR U22904 ( .A(n22321), .B(n22320), .Z(n22354) );
  XNOR U22905 ( .A(n22354), .B(sreg[1558]), .Z(n22356) );
  NAND U22906 ( .A(n22313), .B(sreg[1557]), .Z(n22317) );
  OR U22907 ( .A(n22315), .B(n22314), .Z(n22316) );
  AND U22908 ( .A(n22317), .B(n22316), .Z(n22355) );
  XOR U22909 ( .A(n22356), .B(n22355), .Z(c[1558]) );
  NANDN U22910 ( .A(n22319), .B(n22318), .Z(n22323) );
  NAND U22911 ( .A(n22321), .B(n22320), .Z(n22322) );
  NAND U22912 ( .A(n22323), .B(n22322), .Z(n22362) );
  NAND U22913 ( .A(b[0]), .B(a[543]), .Z(n22324) );
  XNOR U22914 ( .A(b[1]), .B(n22324), .Z(n22326) );
  NAND U22915 ( .A(n92), .B(a[542]), .Z(n22325) );
  AND U22916 ( .A(n22326), .B(n22325), .Z(n22379) );
  XOR U22917 ( .A(a[539]), .B(n42197), .Z(n22368) );
  NANDN U22918 ( .A(n22368), .B(n42173), .Z(n22329) );
  NANDN U22919 ( .A(n22327), .B(n42172), .Z(n22328) );
  NAND U22920 ( .A(n22329), .B(n22328), .Z(n22377) );
  NAND U22921 ( .A(b[7]), .B(a[535]), .Z(n22378) );
  XNOR U22922 ( .A(n22377), .B(n22378), .Z(n22380) );
  XOR U22923 ( .A(n22379), .B(n22380), .Z(n22386) );
  NANDN U22924 ( .A(n22330), .B(n42093), .Z(n22332) );
  XOR U22925 ( .A(n42134), .B(a[541]), .Z(n22371) );
  NANDN U22926 ( .A(n22371), .B(n42095), .Z(n22331) );
  NAND U22927 ( .A(n22332), .B(n22331), .Z(n22384) );
  NANDN U22928 ( .A(n22333), .B(n42231), .Z(n22335) );
  XOR U22929 ( .A(n206), .B(a[537]), .Z(n22374) );
  NANDN U22930 ( .A(n22374), .B(n42234), .Z(n22334) );
  AND U22931 ( .A(n22335), .B(n22334), .Z(n22383) );
  XNOR U22932 ( .A(n22384), .B(n22383), .Z(n22385) );
  XNOR U22933 ( .A(n22386), .B(n22385), .Z(n22390) );
  NANDN U22934 ( .A(n22337), .B(n22336), .Z(n22341) );
  NAND U22935 ( .A(n22339), .B(n22338), .Z(n22340) );
  AND U22936 ( .A(n22341), .B(n22340), .Z(n22389) );
  XOR U22937 ( .A(n22390), .B(n22389), .Z(n22391) );
  NANDN U22938 ( .A(n22343), .B(n22342), .Z(n22347) );
  NANDN U22939 ( .A(n22345), .B(n22344), .Z(n22346) );
  NAND U22940 ( .A(n22347), .B(n22346), .Z(n22392) );
  XOR U22941 ( .A(n22391), .B(n22392), .Z(n22359) );
  OR U22942 ( .A(n22349), .B(n22348), .Z(n22353) );
  NANDN U22943 ( .A(n22351), .B(n22350), .Z(n22352) );
  NAND U22944 ( .A(n22353), .B(n22352), .Z(n22360) );
  XNOR U22945 ( .A(n22359), .B(n22360), .Z(n22361) );
  XNOR U22946 ( .A(n22362), .B(n22361), .Z(n22395) );
  XNOR U22947 ( .A(n22395), .B(sreg[1559]), .Z(n22397) );
  NAND U22948 ( .A(n22354), .B(sreg[1558]), .Z(n22358) );
  OR U22949 ( .A(n22356), .B(n22355), .Z(n22357) );
  AND U22950 ( .A(n22358), .B(n22357), .Z(n22396) );
  XOR U22951 ( .A(n22397), .B(n22396), .Z(c[1559]) );
  NANDN U22952 ( .A(n22360), .B(n22359), .Z(n22364) );
  NAND U22953 ( .A(n22362), .B(n22361), .Z(n22363) );
  NAND U22954 ( .A(n22364), .B(n22363), .Z(n22403) );
  NAND U22955 ( .A(b[0]), .B(a[544]), .Z(n22365) );
  XNOR U22956 ( .A(b[1]), .B(n22365), .Z(n22367) );
  NAND U22957 ( .A(n92), .B(a[543]), .Z(n22366) );
  AND U22958 ( .A(n22367), .B(n22366), .Z(n22420) );
  XOR U22959 ( .A(a[540]), .B(n42197), .Z(n22409) );
  NANDN U22960 ( .A(n22409), .B(n42173), .Z(n22370) );
  NANDN U22961 ( .A(n22368), .B(n42172), .Z(n22369) );
  NAND U22962 ( .A(n22370), .B(n22369), .Z(n22418) );
  NAND U22963 ( .A(b[7]), .B(a[536]), .Z(n22419) );
  XNOR U22964 ( .A(n22418), .B(n22419), .Z(n22421) );
  XOR U22965 ( .A(n22420), .B(n22421), .Z(n22427) );
  NANDN U22966 ( .A(n22371), .B(n42093), .Z(n22373) );
  XOR U22967 ( .A(n42134), .B(a[542]), .Z(n22412) );
  NANDN U22968 ( .A(n22412), .B(n42095), .Z(n22372) );
  NAND U22969 ( .A(n22373), .B(n22372), .Z(n22425) );
  NANDN U22970 ( .A(n22374), .B(n42231), .Z(n22376) );
  XOR U22971 ( .A(n206), .B(a[538]), .Z(n22415) );
  NANDN U22972 ( .A(n22415), .B(n42234), .Z(n22375) );
  AND U22973 ( .A(n22376), .B(n22375), .Z(n22424) );
  XNOR U22974 ( .A(n22425), .B(n22424), .Z(n22426) );
  XNOR U22975 ( .A(n22427), .B(n22426), .Z(n22431) );
  NANDN U22976 ( .A(n22378), .B(n22377), .Z(n22382) );
  NAND U22977 ( .A(n22380), .B(n22379), .Z(n22381) );
  AND U22978 ( .A(n22382), .B(n22381), .Z(n22430) );
  XOR U22979 ( .A(n22431), .B(n22430), .Z(n22432) );
  NANDN U22980 ( .A(n22384), .B(n22383), .Z(n22388) );
  NANDN U22981 ( .A(n22386), .B(n22385), .Z(n22387) );
  NAND U22982 ( .A(n22388), .B(n22387), .Z(n22433) );
  XOR U22983 ( .A(n22432), .B(n22433), .Z(n22400) );
  OR U22984 ( .A(n22390), .B(n22389), .Z(n22394) );
  NANDN U22985 ( .A(n22392), .B(n22391), .Z(n22393) );
  NAND U22986 ( .A(n22394), .B(n22393), .Z(n22401) );
  XNOR U22987 ( .A(n22400), .B(n22401), .Z(n22402) );
  XNOR U22988 ( .A(n22403), .B(n22402), .Z(n22436) );
  XNOR U22989 ( .A(n22436), .B(sreg[1560]), .Z(n22438) );
  NAND U22990 ( .A(n22395), .B(sreg[1559]), .Z(n22399) );
  OR U22991 ( .A(n22397), .B(n22396), .Z(n22398) );
  AND U22992 ( .A(n22399), .B(n22398), .Z(n22437) );
  XOR U22993 ( .A(n22438), .B(n22437), .Z(c[1560]) );
  NANDN U22994 ( .A(n22401), .B(n22400), .Z(n22405) );
  NAND U22995 ( .A(n22403), .B(n22402), .Z(n22404) );
  NAND U22996 ( .A(n22405), .B(n22404), .Z(n22444) );
  NAND U22997 ( .A(b[0]), .B(a[545]), .Z(n22406) );
  XNOR U22998 ( .A(b[1]), .B(n22406), .Z(n22408) );
  NAND U22999 ( .A(n92), .B(a[544]), .Z(n22407) );
  AND U23000 ( .A(n22408), .B(n22407), .Z(n22461) );
  XOR U23001 ( .A(a[541]), .B(n42197), .Z(n22450) );
  NANDN U23002 ( .A(n22450), .B(n42173), .Z(n22411) );
  NANDN U23003 ( .A(n22409), .B(n42172), .Z(n22410) );
  NAND U23004 ( .A(n22411), .B(n22410), .Z(n22459) );
  NAND U23005 ( .A(b[7]), .B(a[537]), .Z(n22460) );
  XNOR U23006 ( .A(n22459), .B(n22460), .Z(n22462) );
  XOR U23007 ( .A(n22461), .B(n22462), .Z(n22468) );
  NANDN U23008 ( .A(n22412), .B(n42093), .Z(n22414) );
  XOR U23009 ( .A(n42134), .B(a[543]), .Z(n22453) );
  NANDN U23010 ( .A(n22453), .B(n42095), .Z(n22413) );
  NAND U23011 ( .A(n22414), .B(n22413), .Z(n22466) );
  NANDN U23012 ( .A(n22415), .B(n42231), .Z(n22417) );
  XOR U23013 ( .A(n207), .B(a[539]), .Z(n22456) );
  NANDN U23014 ( .A(n22456), .B(n42234), .Z(n22416) );
  AND U23015 ( .A(n22417), .B(n22416), .Z(n22465) );
  XNOR U23016 ( .A(n22466), .B(n22465), .Z(n22467) );
  XNOR U23017 ( .A(n22468), .B(n22467), .Z(n22472) );
  NANDN U23018 ( .A(n22419), .B(n22418), .Z(n22423) );
  NAND U23019 ( .A(n22421), .B(n22420), .Z(n22422) );
  AND U23020 ( .A(n22423), .B(n22422), .Z(n22471) );
  XOR U23021 ( .A(n22472), .B(n22471), .Z(n22473) );
  NANDN U23022 ( .A(n22425), .B(n22424), .Z(n22429) );
  NANDN U23023 ( .A(n22427), .B(n22426), .Z(n22428) );
  NAND U23024 ( .A(n22429), .B(n22428), .Z(n22474) );
  XOR U23025 ( .A(n22473), .B(n22474), .Z(n22441) );
  OR U23026 ( .A(n22431), .B(n22430), .Z(n22435) );
  NANDN U23027 ( .A(n22433), .B(n22432), .Z(n22434) );
  NAND U23028 ( .A(n22435), .B(n22434), .Z(n22442) );
  XNOR U23029 ( .A(n22441), .B(n22442), .Z(n22443) );
  XNOR U23030 ( .A(n22444), .B(n22443), .Z(n22477) );
  XNOR U23031 ( .A(n22477), .B(sreg[1561]), .Z(n22479) );
  NAND U23032 ( .A(n22436), .B(sreg[1560]), .Z(n22440) );
  OR U23033 ( .A(n22438), .B(n22437), .Z(n22439) );
  AND U23034 ( .A(n22440), .B(n22439), .Z(n22478) );
  XOR U23035 ( .A(n22479), .B(n22478), .Z(c[1561]) );
  NANDN U23036 ( .A(n22442), .B(n22441), .Z(n22446) );
  NAND U23037 ( .A(n22444), .B(n22443), .Z(n22445) );
  NAND U23038 ( .A(n22446), .B(n22445), .Z(n22485) );
  NAND U23039 ( .A(b[0]), .B(a[546]), .Z(n22447) );
  XNOR U23040 ( .A(b[1]), .B(n22447), .Z(n22449) );
  NAND U23041 ( .A(n93), .B(a[545]), .Z(n22448) );
  AND U23042 ( .A(n22449), .B(n22448), .Z(n22502) );
  XOR U23043 ( .A(a[542]), .B(n42197), .Z(n22491) );
  NANDN U23044 ( .A(n22491), .B(n42173), .Z(n22452) );
  NANDN U23045 ( .A(n22450), .B(n42172), .Z(n22451) );
  NAND U23046 ( .A(n22452), .B(n22451), .Z(n22500) );
  NAND U23047 ( .A(b[7]), .B(a[538]), .Z(n22501) );
  XNOR U23048 ( .A(n22500), .B(n22501), .Z(n22503) );
  XOR U23049 ( .A(n22502), .B(n22503), .Z(n22509) );
  NANDN U23050 ( .A(n22453), .B(n42093), .Z(n22455) );
  XOR U23051 ( .A(n42134), .B(a[544]), .Z(n22494) );
  NANDN U23052 ( .A(n22494), .B(n42095), .Z(n22454) );
  NAND U23053 ( .A(n22455), .B(n22454), .Z(n22507) );
  NANDN U23054 ( .A(n22456), .B(n42231), .Z(n22458) );
  XOR U23055 ( .A(n207), .B(a[540]), .Z(n22497) );
  NANDN U23056 ( .A(n22497), .B(n42234), .Z(n22457) );
  AND U23057 ( .A(n22458), .B(n22457), .Z(n22506) );
  XNOR U23058 ( .A(n22507), .B(n22506), .Z(n22508) );
  XNOR U23059 ( .A(n22509), .B(n22508), .Z(n22513) );
  NANDN U23060 ( .A(n22460), .B(n22459), .Z(n22464) );
  NAND U23061 ( .A(n22462), .B(n22461), .Z(n22463) );
  AND U23062 ( .A(n22464), .B(n22463), .Z(n22512) );
  XOR U23063 ( .A(n22513), .B(n22512), .Z(n22514) );
  NANDN U23064 ( .A(n22466), .B(n22465), .Z(n22470) );
  NANDN U23065 ( .A(n22468), .B(n22467), .Z(n22469) );
  NAND U23066 ( .A(n22470), .B(n22469), .Z(n22515) );
  XOR U23067 ( .A(n22514), .B(n22515), .Z(n22482) );
  OR U23068 ( .A(n22472), .B(n22471), .Z(n22476) );
  NANDN U23069 ( .A(n22474), .B(n22473), .Z(n22475) );
  NAND U23070 ( .A(n22476), .B(n22475), .Z(n22483) );
  XNOR U23071 ( .A(n22482), .B(n22483), .Z(n22484) );
  XNOR U23072 ( .A(n22485), .B(n22484), .Z(n22518) );
  XNOR U23073 ( .A(n22518), .B(sreg[1562]), .Z(n22520) );
  NAND U23074 ( .A(n22477), .B(sreg[1561]), .Z(n22481) );
  OR U23075 ( .A(n22479), .B(n22478), .Z(n22480) );
  AND U23076 ( .A(n22481), .B(n22480), .Z(n22519) );
  XOR U23077 ( .A(n22520), .B(n22519), .Z(c[1562]) );
  NANDN U23078 ( .A(n22483), .B(n22482), .Z(n22487) );
  NAND U23079 ( .A(n22485), .B(n22484), .Z(n22486) );
  NAND U23080 ( .A(n22487), .B(n22486), .Z(n22526) );
  NAND U23081 ( .A(b[0]), .B(a[547]), .Z(n22488) );
  XNOR U23082 ( .A(b[1]), .B(n22488), .Z(n22490) );
  NAND U23083 ( .A(n93), .B(a[546]), .Z(n22489) );
  AND U23084 ( .A(n22490), .B(n22489), .Z(n22543) );
  XOR U23085 ( .A(a[543]), .B(n42197), .Z(n22532) );
  NANDN U23086 ( .A(n22532), .B(n42173), .Z(n22493) );
  NANDN U23087 ( .A(n22491), .B(n42172), .Z(n22492) );
  NAND U23088 ( .A(n22493), .B(n22492), .Z(n22541) );
  NAND U23089 ( .A(b[7]), .B(a[539]), .Z(n22542) );
  XNOR U23090 ( .A(n22541), .B(n22542), .Z(n22544) );
  XOR U23091 ( .A(n22543), .B(n22544), .Z(n22550) );
  NANDN U23092 ( .A(n22494), .B(n42093), .Z(n22496) );
  XOR U23093 ( .A(n42134), .B(a[545]), .Z(n22535) );
  NANDN U23094 ( .A(n22535), .B(n42095), .Z(n22495) );
  NAND U23095 ( .A(n22496), .B(n22495), .Z(n22548) );
  NANDN U23096 ( .A(n22497), .B(n42231), .Z(n22499) );
  XOR U23097 ( .A(n207), .B(a[541]), .Z(n22538) );
  NANDN U23098 ( .A(n22538), .B(n42234), .Z(n22498) );
  AND U23099 ( .A(n22499), .B(n22498), .Z(n22547) );
  XNOR U23100 ( .A(n22548), .B(n22547), .Z(n22549) );
  XNOR U23101 ( .A(n22550), .B(n22549), .Z(n22554) );
  NANDN U23102 ( .A(n22501), .B(n22500), .Z(n22505) );
  NAND U23103 ( .A(n22503), .B(n22502), .Z(n22504) );
  AND U23104 ( .A(n22505), .B(n22504), .Z(n22553) );
  XOR U23105 ( .A(n22554), .B(n22553), .Z(n22555) );
  NANDN U23106 ( .A(n22507), .B(n22506), .Z(n22511) );
  NANDN U23107 ( .A(n22509), .B(n22508), .Z(n22510) );
  NAND U23108 ( .A(n22511), .B(n22510), .Z(n22556) );
  XOR U23109 ( .A(n22555), .B(n22556), .Z(n22523) );
  OR U23110 ( .A(n22513), .B(n22512), .Z(n22517) );
  NANDN U23111 ( .A(n22515), .B(n22514), .Z(n22516) );
  NAND U23112 ( .A(n22517), .B(n22516), .Z(n22524) );
  XNOR U23113 ( .A(n22523), .B(n22524), .Z(n22525) );
  XNOR U23114 ( .A(n22526), .B(n22525), .Z(n22559) );
  XNOR U23115 ( .A(n22559), .B(sreg[1563]), .Z(n22561) );
  NAND U23116 ( .A(n22518), .B(sreg[1562]), .Z(n22522) );
  OR U23117 ( .A(n22520), .B(n22519), .Z(n22521) );
  AND U23118 ( .A(n22522), .B(n22521), .Z(n22560) );
  XOR U23119 ( .A(n22561), .B(n22560), .Z(c[1563]) );
  NANDN U23120 ( .A(n22524), .B(n22523), .Z(n22528) );
  NAND U23121 ( .A(n22526), .B(n22525), .Z(n22527) );
  NAND U23122 ( .A(n22528), .B(n22527), .Z(n22567) );
  NAND U23123 ( .A(b[0]), .B(a[548]), .Z(n22529) );
  XNOR U23124 ( .A(b[1]), .B(n22529), .Z(n22531) );
  NAND U23125 ( .A(n93), .B(a[547]), .Z(n22530) );
  AND U23126 ( .A(n22531), .B(n22530), .Z(n22584) );
  XOR U23127 ( .A(a[544]), .B(n42197), .Z(n22573) );
  NANDN U23128 ( .A(n22573), .B(n42173), .Z(n22534) );
  NANDN U23129 ( .A(n22532), .B(n42172), .Z(n22533) );
  NAND U23130 ( .A(n22534), .B(n22533), .Z(n22582) );
  NAND U23131 ( .A(b[7]), .B(a[540]), .Z(n22583) );
  XNOR U23132 ( .A(n22582), .B(n22583), .Z(n22585) );
  XOR U23133 ( .A(n22584), .B(n22585), .Z(n22591) );
  NANDN U23134 ( .A(n22535), .B(n42093), .Z(n22537) );
  XOR U23135 ( .A(n42134), .B(a[546]), .Z(n22576) );
  NANDN U23136 ( .A(n22576), .B(n42095), .Z(n22536) );
  NAND U23137 ( .A(n22537), .B(n22536), .Z(n22589) );
  NANDN U23138 ( .A(n22538), .B(n42231), .Z(n22540) );
  XOR U23139 ( .A(n207), .B(a[542]), .Z(n22579) );
  NANDN U23140 ( .A(n22579), .B(n42234), .Z(n22539) );
  AND U23141 ( .A(n22540), .B(n22539), .Z(n22588) );
  XNOR U23142 ( .A(n22589), .B(n22588), .Z(n22590) );
  XNOR U23143 ( .A(n22591), .B(n22590), .Z(n22595) );
  NANDN U23144 ( .A(n22542), .B(n22541), .Z(n22546) );
  NAND U23145 ( .A(n22544), .B(n22543), .Z(n22545) );
  AND U23146 ( .A(n22546), .B(n22545), .Z(n22594) );
  XOR U23147 ( .A(n22595), .B(n22594), .Z(n22596) );
  NANDN U23148 ( .A(n22548), .B(n22547), .Z(n22552) );
  NANDN U23149 ( .A(n22550), .B(n22549), .Z(n22551) );
  NAND U23150 ( .A(n22552), .B(n22551), .Z(n22597) );
  XOR U23151 ( .A(n22596), .B(n22597), .Z(n22564) );
  OR U23152 ( .A(n22554), .B(n22553), .Z(n22558) );
  NANDN U23153 ( .A(n22556), .B(n22555), .Z(n22557) );
  NAND U23154 ( .A(n22558), .B(n22557), .Z(n22565) );
  XNOR U23155 ( .A(n22564), .B(n22565), .Z(n22566) );
  XNOR U23156 ( .A(n22567), .B(n22566), .Z(n22600) );
  XNOR U23157 ( .A(n22600), .B(sreg[1564]), .Z(n22602) );
  NAND U23158 ( .A(n22559), .B(sreg[1563]), .Z(n22563) );
  OR U23159 ( .A(n22561), .B(n22560), .Z(n22562) );
  AND U23160 ( .A(n22563), .B(n22562), .Z(n22601) );
  XOR U23161 ( .A(n22602), .B(n22601), .Z(c[1564]) );
  NANDN U23162 ( .A(n22565), .B(n22564), .Z(n22569) );
  NAND U23163 ( .A(n22567), .B(n22566), .Z(n22568) );
  NAND U23164 ( .A(n22569), .B(n22568), .Z(n22608) );
  NAND U23165 ( .A(b[0]), .B(a[549]), .Z(n22570) );
  XNOR U23166 ( .A(b[1]), .B(n22570), .Z(n22572) );
  NAND U23167 ( .A(n93), .B(a[548]), .Z(n22571) );
  AND U23168 ( .A(n22572), .B(n22571), .Z(n22625) );
  XOR U23169 ( .A(a[545]), .B(n42197), .Z(n22614) );
  NANDN U23170 ( .A(n22614), .B(n42173), .Z(n22575) );
  NANDN U23171 ( .A(n22573), .B(n42172), .Z(n22574) );
  NAND U23172 ( .A(n22575), .B(n22574), .Z(n22623) );
  NAND U23173 ( .A(b[7]), .B(a[541]), .Z(n22624) );
  XNOR U23174 ( .A(n22623), .B(n22624), .Z(n22626) );
  XOR U23175 ( .A(n22625), .B(n22626), .Z(n22632) );
  NANDN U23176 ( .A(n22576), .B(n42093), .Z(n22578) );
  XOR U23177 ( .A(n42134), .B(a[547]), .Z(n22617) );
  NANDN U23178 ( .A(n22617), .B(n42095), .Z(n22577) );
  NAND U23179 ( .A(n22578), .B(n22577), .Z(n22630) );
  NANDN U23180 ( .A(n22579), .B(n42231), .Z(n22581) );
  XOR U23181 ( .A(n207), .B(a[543]), .Z(n22620) );
  NANDN U23182 ( .A(n22620), .B(n42234), .Z(n22580) );
  AND U23183 ( .A(n22581), .B(n22580), .Z(n22629) );
  XNOR U23184 ( .A(n22630), .B(n22629), .Z(n22631) );
  XNOR U23185 ( .A(n22632), .B(n22631), .Z(n22636) );
  NANDN U23186 ( .A(n22583), .B(n22582), .Z(n22587) );
  NAND U23187 ( .A(n22585), .B(n22584), .Z(n22586) );
  AND U23188 ( .A(n22587), .B(n22586), .Z(n22635) );
  XOR U23189 ( .A(n22636), .B(n22635), .Z(n22637) );
  NANDN U23190 ( .A(n22589), .B(n22588), .Z(n22593) );
  NANDN U23191 ( .A(n22591), .B(n22590), .Z(n22592) );
  NAND U23192 ( .A(n22593), .B(n22592), .Z(n22638) );
  XOR U23193 ( .A(n22637), .B(n22638), .Z(n22605) );
  OR U23194 ( .A(n22595), .B(n22594), .Z(n22599) );
  NANDN U23195 ( .A(n22597), .B(n22596), .Z(n22598) );
  NAND U23196 ( .A(n22599), .B(n22598), .Z(n22606) );
  XNOR U23197 ( .A(n22605), .B(n22606), .Z(n22607) );
  XNOR U23198 ( .A(n22608), .B(n22607), .Z(n22641) );
  XNOR U23199 ( .A(n22641), .B(sreg[1565]), .Z(n22643) );
  NAND U23200 ( .A(n22600), .B(sreg[1564]), .Z(n22604) );
  OR U23201 ( .A(n22602), .B(n22601), .Z(n22603) );
  AND U23202 ( .A(n22604), .B(n22603), .Z(n22642) );
  XOR U23203 ( .A(n22643), .B(n22642), .Z(c[1565]) );
  NANDN U23204 ( .A(n22606), .B(n22605), .Z(n22610) );
  NAND U23205 ( .A(n22608), .B(n22607), .Z(n22609) );
  NAND U23206 ( .A(n22610), .B(n22609), .Z(n22649) );
  NAND U23207 ( .A(b[0]), .B(a[550]), .Z(n22611) );
  XNOR U23208 ( .A(b[1]), .B(n22611), .Z(n22613) );
  NAND U23209 ( .A(n93), .B(a[549]), .Z(n22612) );
  AND U23210 ( .A(n22613), .B(n22612), .Z(n22666) );
  XOR U23211 ( .A(a[546]), .B(n42197), .Z(n22655) );
  NANDN U23212 ( .A(n22655), .B(n42173), .Z(n22616) );
  NANDN U23213 ( .A(n22614), .B(n42172), .Z(n22615) );
  NAND U23214 ( .A(n22616), .B(n22615), .Z(n22664) );
  NAND U23215 ( .A(b[7]), .B(a[542]), .Z(n22665) );
  XNOR U23216 ( .A(n22664), .B(n22665), .Z(n22667) );
  XOR U23217 ( .A(n22666), .B(n22667), .Z(n22673) );
  NANDN U23218 ( .A(n22617), .B(n42093), .Z(n22619) );
  XOR U23219 ( .A(n42134), .B(a[548]), .Z(n22658) );
  NANDN U23220 ( .A(n22658), .B(n42095), .Z(n22618) );
  NAND U23221 ( .A(n22619), .B(n22618), .Z(n22671) );
  NANDN U23222 ( .A(n22620), .B(n42231), .Z(n22622) );
  XOR U23223 ( .A(n207), .B(a[544]), .Z(n22661) );
  NANDN U23224 ( .A(n22661), .B(n42234), .Z(n22621) );
  AND U23225 ( .A(n22622), .B(n22621), .Z(n22670) );
  XNOR U23226 ( .A(n22671), .B(n22670), .Z(n22672) );
  XNOR U23227 ( .A(n22673), .B(n22672), .Z(n22677) );
  NANDN U23228 ( .A(n22624), .B(n22623), .Z(n22628) );
  NAND U23229 ( .A(n22626), .B(n22625), .Z(n22627) );
  AND U23230 ( .A(n22628), .B(n22627), .Z(n22676) );
  XOR U23231 ( .A(n22677), .B(n22676), .Z(n22678) );
  NANDN U23232 ( .A(n22630), .B(n22629), .Z(n22634) );
  NANDN U23233 ( .A(n22632), .B(n22631), .Z(n22633) );
  NAND U23234 ( .A(n22634), .B(n22633), .Z(n22679) );
  XOR U23235 ( .A(n22678), .B(n22679), .Z(n22646) );
  OR U23236 ( .A(n22636), .B(n22635), .Z(n22640) );
  NANDN U23237 ( .A(n22638), .B(n22637), .Z(n22639) );
  NAND U23238 ( .A(n22640), .B(n22639), .Z(n22647) );
  XNOR U23239 ( .A(n22646), .B(n22647), .Z(n22648) );
  XNOR U23240 ( .A(n22649), .B(n22648), .Z(n22682) );
  XNOR U23241 ( .A(n22682), .B(sreg[1566]), .Z(n22684) );
  NAND U23242 ( .A(n22641), .B(sreg[1565]), .Z(n22645) );
  OR U23243 ( .A(n22643), .B(n22642), .Z(n22644) );
  AND U23244 ( .A(n22645), .B(n22644), .Z(n22683) );
  XOR U23245 ( .A(n22684), .B(n22683), .Z(c[1566]) );
  NANDN U23246 ( .A(n22647), .B(n22646), .Z(n22651) );
  NAND U23247 ( .A(n22649), .B(n22648), .Z(n22650) );
  NAND U23248 ( .A(n22651), .B(n22650), .Z(n22690) );
  NAND U23249 ( .A(b[0]), .B(a[551]), .Z(n22652) );
  XNOR U23250 ( .A(b[1]), .B(n22652), .Z(n22654) );
  NAND U23251 ( .A(n93), .B(a[550]), .Z(n22653) );
  AND U23252 ( .A(n22654), .B(n22653), .Z(n22707) );
  XOR U23253 ( .A(a[547]), .B(n42197), .Z(n22696) );
  NANDN U23254 ( .A(n22696), .B(n42173), .Z(n22657) );
  NANDN U23255 ( .A(n22655), .B(n42172), .Z(n22656) );
  NAND U23256 ( .A(n22657), .B(n22656), .Z(n22705) );
  NAND U23257 ( .A(b[7]), .B(a[543]), .Z(n22706) );
  XNOR U23258 ( .A(n22705), .B(n22706), .Z(n22708) );
  XOR U23259 ( .A(n22707), .B(n22708), .Z(n22714) );
  NANDN U23260 ( .A(n22658), .B(n42093), .Z(n22660) );
  XOR U23261 ( .A(n42134), .B(a[549]), .Z(n22699) );
  NANDN U23262 ( .A(n22699), .B(n42095), .Z(n22659) );
  NAND U23263 ( .A(n22660), .B(n22659), .Z(n22712) );
  NANDN U23264 ( .A(n22661), .B(n42231), .Z(n22663) );
  XOR U23265 ( .A(n207), .B(a[545]), .Z(n22702) );
  NANDN U23266 ( .A(n22702), .B(n42234), .Z(n22662) );
  AND U23267 ( .A(n22663), .B(n22662), .Z(n22711) );
  XNOR U23268 ( .A(n22712), .B(n22711), .Z(n22713) );
  XNOR U23269 ( .A(n22714), .B(n22713), .Z(n22718) );
  NANDN U23270 ( .A(n22665), .B(n22664), .Z(n22669) );
  NAND U23271 ( .A(n22667), .B(n22666), .Z(n22668) );
  AND U23272 ( .A(n22669), .B(n22668), .Z(n22717) );
  XOR U23273 ( .A(n22718), .B(n22717), .Z(n22719) );
  NANDN U23274 ( .A(n22671), .B(n22670), .Z(n22675) );
  NANDN U23275 ( .A(n22673), .B(n22672), .Z(n22674) );
  NAND U23276 ( .A(n22675), .B(n22674), .Z(n22720) );
  XOR U23277 ( .A(n22719), .B(n22720), .Z(n22687) );
  OR U23278 ( .A(n22677), .B(n22676), .Z(n22681) );
  NANDN U23279 ( .A(n22679), .B(n22678), .Z(n22680) );
  NAND U23280 ( .A(n22681), .B(n22680), .Z(n22688) );
  XNOR U23281 ( .A(n22687), .B(n22688), .Z(n22689) );
  XNOR U23282 ( .A(n22690), .B(n22689), .Z(n22723) );
  XNOR U23283 ( .A(n22723), .B(sreg[1567]), .Z(n22725) );
  NAND U23284 ( .A(n22682), .B(sreg[1566]), .Z(n22686) );
  OR U23285 ( .A(n22684), .B(n22683), .Z(n22685) );
  AND U23286 ( .A(n22686), .B(n22685), .Z(n22724) );
  XOR U23287 ( .A(n22725), .B(n22724), .Z(c[1567]) );
  NANDN U23288 ( .A(n22688), .B(n22687), .Z(n22692) );
  NAND U23289 ( .A(n22690), .B(n22689), .Z(n22691) );
  NAND U23290 ( .A(n22692), .B(n22691), .Z(n22731) );
  NAND U23291 ( .A(b[0]), .B(a[552]), .Z(n22693) );
  XNOR U23292 ( .A(b[1]), .B(n22693), .Z(n22695) );
  NAND U23293 ( .A(n93), .B(a[551]), .Z(n22694) );
  AND U23294 ( .A(n22695), .B(n22694), .Z(n22748) );
  XOR U23295 ( .A(a[548]), .B(n42197), .Z(n22737) );
  NANDN U23296 ( .A(n22737), .B(n42173), .Z(n22698) );
  NANDN U23297 ( .A(n22696), .B(n42172), .Z(n22697) );
  NAND U23298 ( .A(n22698), .B(n22697), .Z(n22746) );
  NAND U23299 ( .A(b[7]), .B(a[544]), .Z(n22747) );
  XNOR U23300 ( .A(n22746), .B(n22747), .Z(n22749) );
  XOR U23301 ( .A(n22748), .B(n22749), .Z(n22755) );
  NANDN U23302 ( .A(n22699), .B(n42093), .Z(n22701) );
  XOR U23303 ( .A(n42134), .B(a[550]), .Z(n22740) );
  NANDN U23304 ( .A(n22740), .B(n42095), .Z(n22700) );
  NAND U23305 ( .A(n22701), .B(n22700), .Z(n22753) );
  NANDN U23306 ( .A(n22702), .B(n42231), .Z(n22704) );
  XOR U23307 ( .A(n207), .B(a[546]), .Z(n22743) );
  NANDN U23308 ( .A(n22743), .B(n42234), .Z(n22703) );
  AND U23309 ( .A(n22704), .B(n22703), .Z(n22752) );
  XNOR U23310 ( .A(n22753), .B(n22752), .Z(n22754) );
  XNOR U23311 ( .A(n22755), .B(n22754), .Z(n22759) );
  NANDN U23312 ( .A(n22706), .B(n22705), .Z(n22710) );
  NAND U23313 ( .A(n22708), .B(n22707), .Z(n22709) );
  AND U23314 ( .A(n22710), .B(n22709), .Z(n22758) );
  XOR U23315 ( .A(n22759), .B(n22758), .Z(n22760) );
  NANDN U23316 ( .A(n22712), .B(n22711), .Z(n22716) );
  NANDN U23317 ( .A(n22714), .B(n22713), .Z(n22715) );
  NAND U23318 ( .A(n22716), .B(n22715), .Z(n22761) );
  XOR U23319 ( .A(n22760), .B(n22761), .Z(n22728) );
  OR U23320 ( .A(n22718), .B(n22717), .Z(n22722) );
  NANDN U23321 ( .A(n22720), .B(n22719), .Z(n22721) );
  NAND U23322 ( .A(n22722), .B(n22721), .Z(n22729) );
  XNOR U23323 ( .A(n22728), .B(n22729), .Z(n22730) );
  XNOR U23324 ( .A(n22731), .B(n22730), .Z(n22764) );
  XNOR U23325 ( .A(n22764), .B(sreg[1568]), .Z(n22766) );
  NAND U23326 ( .A(n22723), .B(sreg[1567]), .Z(n22727) );
  OR U23327 ( .A(n22725), .B(n22724), .Z(n22726) );
  AND U23328 ( .A(n22727), .B(n22726), .Z(n22765) );
  XOR U23329 ( .A(n22766), .B(n22765), .Z(c[1568]) );
  NANDN U23330 ( .A(n22729), .B(n22728), .Z(n22733) );
  NAND U23331 ( .A(n22731), .B(n22730), .Z(n22732) );
  NAND U23332 ( .A(n22733), .B(n22732), .Z(n22772) );
  NAND U23333 ( .A(b[0]), .B(a[553]), .Z(n22734) );
  XNOR U23334 ( .A(b[1]), .B(n22734), .Z(n22736) );
  NAND U23335 ( .A(n94), .B(a[552]), .Z(n22735) );
  AND U23336 ( .A(n22736), .B(n22735), .Z(n22789) );
  XOR U23337 ( .A(a[549]), .B(n42197), .Z(n22778) );
  NANDN U23338 ( .A(n22778), .B(n42173), .Z(n22739) );
  NANDN U23339 ( .A(n22737), .B(n42172), .Z(n22738) );
  NAND U23340 ( .A(n22739), .B(n22738), .Z(n22787) );
  NAND U23341 ( .A(b[7]), .B(a[545]), .Z(n22788) );
  XNOR U23342 ( .A(n22787), .B(n22788), .Z(n22790) );
  XOR U23343 ( .A(n22789), .B(n22790), .Z(n22796) );
  NANDN U23344 ( .A(n22740), .B(n42093), .Z(n22742) );
  XOR U23345 ( .A(n42134), .B(a[551]), .Z(n22781) );
  NANDN U23346 ( .A(n22781), .B(n42095), .Z(n22741) );
  NAND U23347 ( .A(n22742), .B(n22741), .Z(n22794) );
  NANDN U23348 ( .A(n22743), .B(n42231), .Z(n22745) );
  XOR U23349 ( .A(n207), .B(a[547]), .Z(n22784) );
  NANDN U23350 ( .A(n22784), .B(n42234), .Z(n22744) );
  AND U23351 ( .A(n22745), .B(n22744), .Z(n22793) );
  XNOR U23352 ( .A(n22794), .B(n22793), .Z(n22795) );
  XNOR U23353 ( .A(n22796), .B(n22795), .Z(n22800) );
  NANDN U23354 ( .A(n22747), .B(n22746), .Z(n22751) );
  NAND U23355 ( .A(n22749), .B(n22748), .Z(n22750) );
  AND U23356 ( .A(n22751), .B(n22750), .Z(n22799) );
  XOR U23357 ( .A(n22800), .B(n22799), .Z(n22801) );
  NANDN U23358 ( .A(n22753), .B(n22752), .Z(n22757) );
  NANDN U23359 ( .A(n22755), .B(n22754), .Z(n22756) );
  NAND U23360 ( .A(n22757), .B(n22756), .Z(n22802) );
  XOR U23361 ( .A(n22801), .B(n22802), .Z(n22769) );
  OR U23362 ( .A(n22759), .B(n22758), .Z(n22763) );
  NANDN U23363 ( .A(n22761), .B(n22760), .Z(n22762) );
  NAND U23364 ( .A(n22763), .B(n22762), .Z(n22770) );
  XNOR U23365 ( .A(n22769), .B(n22770), .Z(n22771) );
  XNOR U23366 ( .A(n22772), .B(n22771), .Z(n22805) );
  XNOR U23367 ( .A(n22805), .B(sreg[1569]), .Z(n22807) );
  NAND U23368 ( .A(n22764), .B(sreg[1568]), .Z(n22768) );
  OR U23369 ( .A(n22766), .B(n22765), .Z(n22767) );
  AND U23370 ( .A(n22768), .B(n22767), .Z(n22806) );
  XOR U23371 ( .A(n22807), .B(n22806), .Z(c[1569]) );
  NANDN U23372 ( .A(n22770), .B(n22769), .Z(n22774) );
  NAND U23373 ( .A(n22772), .B(n22771), .Z(n22773) );
  NAND U23374 ( .A(n22774), .B(n22773), .Z(n22813) );
  NAND U23375 ( .A(b[0]), .B(a[554]), .Z(n22775) );
  XNOR U23376 ( .A(b[1]), .B(n22775), .Z(n22777) );
  NAND U23377 ( .A(n94), .B(a[553]), .Z(n22776) );
  AND U23378 ( .A(n22777), .B(n22776), .Z(n22830) );
  XOR U23379 ( .A(a[550]), .B(n42197), .Z(n22819) );
  NANDN U23380 ( .A(n22819), .B(n42173), .Z(n22780) );
  NANDN U23381 ( .A(n22778), .B(n42172), .Z(n22779) );
  NAND U23382 ( .A(n22780), .B(n22779), .Z(n22828) );
  NAND U23383 ( .A(b[7]), .B(a[546]), .Z(n22829) );
  XNOR U23384 ( .A(n22828), .B(n22829), .Z(n22831) );
  XOR U23385 ( .A(n22830), .B(n22831), .Z(n22837) );
  NANDN U23386 ( .A(n22781), .B(n42093), .Z(n22783) );
  XOR U23387 ( .A(n42134), .B(a[552]), .Z(n22822) );
  NANDN U23388 ( .A(n22822), .B(n42095), .Z(n22782) );
  NAND U23389 ( .A(n22783), .B(n22782), .Z(n22835) );
  NANDN U23390 ( .A(n22784), .B(n42231), .Z(n22786) );
  XOR U23391 ( .A(n207), .B(a[548]), .Z(n22825) );
  NANDN U23392 ( .A(n22825), .B(n42234), .Z(n22785) );
  AND U23393 ( .A(n22786), .B(n22785), .Z(n22834) );
  XNOR U23394 ( .A(n22835), .B(n22834), .Z(n22836) );
  XNOR U23395 ( .A(n22837), .B(n22836), .Z(n22841) );
  NANDN U23396 ( .A(n22788), .B(n22787), .Z(n22792) );
  NAND U23397 ( .A(n22790), .B(n22789), .Z(n22791) );
  AND U23398 ( .A(n22792), .B(n22791), .Z(n22840) );
  XOR U23399 ( .A(n22841), .B(n22840), .Z(n22842) );
  NANDN U23400 ( .A(n22794), .B(n22793), .Z(n22798) );
  NANDN U23401 ( .A(n22796), .B(n22795), .Z(n22797) );
  NAND U23402 ( .A(n22798), .B(n22797), .Z(n22843) );
  XOR U23403 ( .A(n22842), .B(n22843), .Z(n22810) );
  OR U23404 ( .A(n22800), .B(n22799), .Z(n22804) );
  NANDN U23405 ( .A(n22802), .B(n22801), .Z(n22803) );
  NAND U23406 ( .A(n22804), .B(n22803), .Z(n22811) );
  XNOR U23407 ( .A(n22810), .B(n22811), .Z(n22812) );
  XNOR U23408 ( .A(n22813), .B(n22812), .Z(n22846) );
  XNOR U23409 ( .A(n22846), .B(sreg[1570]), .Z(n22848) );
  NAND U23410 ( .A(n22805), .B(sreg[1569]), .Z(n22809) );
  OR U23411 ( .A(n22807), .B(n22806), .Z(n22808) );
  AND U23412 ( .A(n22809), .B(n22808), .Z(n22847) );
  XOR U23413 ( .A(n22848), .B(n22847), .Z(c[1570]) );
  NANDN U23414 ( .A(n22811), .B(n22810), .Z(n22815) );
  NAND U23415 ( .A(n22813), .B(n22812), .Z(n22814) );
  NAND U23416 ( .A(n22815), .B(n22814), .Z(n22854) );
  NAND U23417 ( .A(b[0]), .B(a[555]), .Z(n22816) );
  XNOR U23418 ( .A(b[1]), .B(n22816), .Z(n22818) );
  NAND U23419 ( .A(n94), .B(a[554]), .Z(n22817) );
  AND U23420 ( .A(n22818), .B(n22817), .Z(n22871) );
  XOR U23421 ( .A(a[551]), .B(n42197), .Z(n22860) );
  NANDN U23422 ( .A(n22860), .B(n42173), .Z(n22821) );
  NANDN U23423 ( .A(n22819), .B(n42172), .Z(n22820) );
  NAND U23424 ( .A(n22821), .B(n22820), .Z(n22869) );
  NAND U23425 ( .A(b[7]), .B(a[547]), .Z(n22870) );
  XNOR U23426 ( .A(n22869), .B(n22870), .Z(n22872) );
  XOR U23427 ( .A(n22871), .B(n22872), .Z(n22878) );
  NANDN U23428 ( .A(n22822), .B(n42093), .Z(n22824) );
  XOR U23429 ( .A(n42134), .B(a[553]), .Z(n22863) );
  NANDN U23430 ( .A(n22863), .B(n42095), .Z(n22823) );
  NAND U23431 ( .A(n22824), .B(n22823), .Z(n22876) );
  NANDN U23432 ( .A(n22825), .B(n42231), .Z(n22827) );
  XOR U23433 ( .A(n207), .B(a[549]), .Z(n22866) );
  NANDN U23434 ( .A(n22866), .B(n42234), .Z(n22826) );
  AND U23435 ( .A(n22827), .B(n22826), .Z(n22875) );
  XNOR U23436 ( .A(n22876), .B(n22875), .Z(n22877) );
  XNOR U23437 ( .A(n22878), .B(n22877), .Z(n22882) );
  NANDN U23438 ( .A(n22829), .B(n22828), .Z(n22833) );
  NAND U23439 ( .A(n22831), .B(n22830), .Z(n22832) );
  AND U23440 ( .A(n22833), .B(n22832), .Z(n22881) );
  XOR U23441 ( .A(n22882), .B(n22881), .Z(n22883) );
  NANDN U23442 ( .A(n22835), .B(n22834), .Z(n22839) );
  NANDN U23443 ( .A(n22837), .B(n22836), .Z(n22838) );
  NAND U23444 ( .A(n22839), .B(n22838), .Z(n22884) );
  XOR U23445 ( .A(n22883), .B(n22884), .Z(n22851) );
  OR U23446 ( .A(n22841), .B(n22840), .Z(n22845) );
  NANDN U23447 ( .A(n22843), .B(n22842), .Z(n22844) );
  NAND U23448 ( .A(n22845), .B(n22844), .Z(n22852) );
  XNOR U23449 ( .A(n22851), .B(n22852), .Z(n22853) );
  XNOR U23450 ( .A(n22854), .B(n22853), .Z(n22887) );
  XNOR U23451 ( .A(n22887), .B(sreg[1571]), .Z(n22889) );
  NAND U23452 ( .A(n22846), .B(sreg[1570]), .Z(n22850) );
  OR U23453 ( .A(n22848), .B(n22847), .Z(n22849) );
  AND U23454 ( .A(n22850), .B(n22849), .Z(n22888) );
  XOR U23455 ( .A(n22889), .B(n22888), .Z(c[1571]) );
  NANDN U23456 ( .A(n22852), .B(n22851), .Z(n22856) );
  NAND U23457 ( .A(n22854), .B(n22853), .Z(n22855) );
  NAND U23458 ( .A(n22856), .B(n22855), .Z(n22895) );
  NAND U23459 ( .A(b[0]), .B(a[556]), .Z(n22857) );
  XNOR U23460 ( .A(b[1]), .B(n22857), .Z(n22859) );
  NAND U23461 ( .A(n94), .B(a[555]), .Z(n22858) );
  AND U23462 ( .A(n22859), .B(n22858), .Z(n22912) );
  XOR U23463 ( .A(a[552]), .B(n42197), .Z(n22901) );
  NANDN U23464 ( .A(n22901), .B(n42173), .Z(n22862) );
  NANDN U23465 ( .A(n22860), .B(n42172), .Z(n22861) );
  NAND U23466 ( .A(n22862), .B(n22861), .Z(n22910) );
  NAND U23467 ( .A(b[7]), .B(a[548]), .Z(n22911) );
  XNOR U23468 ( .A(n22910), .B(n22911), .Z(n22913) );
  XOR U23469 ( .A(n22912), .B(n22913), .Z(n22919) );
  NANDN U23470 ( .A(n22863), .B(n42093), .Z(n22865) );
  XOR U23471 ( .A(n42134), .B(a[554]), .Z(n22904) );
  NANDN U23472 ( .A(n22904), .B(n42095), .Z(n22864) );
  NAND U23473 ( .A(n22865), .B(n22864), .Z(n22917) );
  NANDN U23474 ( .A(n22866), .B(n42231), .Z(n22868) );
  XOR U23475 ( .A(n207), .B(a[550]), .Z(n22907) );
  NANDN U23476 ( .A(n22907), .B(n42234), .Z(n22867) );
  AND U23477 ( .A(n22868), .B(n22867), .Z(n22916) );
  XNOR U23478 ( .A(n22917), .B(n22916), .Z(n22918) );
  XNOR U23479 ( .A(n22919), .B(n22918), .Z(n22923) );
  NANDN U23480 ( .A(n22870), .B(n22869), .Z(n22874) );
  NAND U23481 ( .A(n22872), .B(n22871), .Z(n22873) );
  AND U23482 ( .A(n22874), .B(n22873), .Z(n22922) );
  XOR U23483 ( .A(n22923), .B(n22922), .Z(n22924) );
  NANDN U23484 ( .A(n22876), .B(n22875), .Z(n22880) );
  NANDN U23485 ( .A(n22878), .B(n22877), .Z(n22879) );
  NAND U23486 ( .A(n22880), .B(n22879), .Z(n22925) );
  XOR U23487 ( .A(n22924), .B(n22925), .Z(n22892) );
  OR U23488 ( .A(n22882), .B(n22881), .Z(n22886) );
  NANDN U23489 ( .A(n22884), .B(n22883), .Z(n22885) );
  NAND U23490 ( .A(n22886), .B(n22885), .Z(n22893) );
  XNOR U23491 ( .A(n22892), .B(n22893), .Z(n22894) );
  XNOR U23492 ( .A(n22895), .B(n22894), .Z(n22928) );
  XNOR U23493 ( .A(n22928), .B(sreg[1572]), .Z(n22930) );
  NAND U23494 ( .A(n22887), .B(sreg[1571]), .Z(n22891) );
  OR U23495 ( .A(n22889), .B(n22888), .Z(n22890) );
  AND U23496 ( .A(n22891), .B(n22890), .Z(n22929) );
  XOR U23497 ( .A(n22930), .B(n22929), .Z(c[1572]) );
  NANDN U23498 ( .A(n22893), .B(n22892), .Z(n22897) );
  NAND U23499 ( .A(n22895), .B(n22894), .Z(n22896) );
  NAND U23500 ( .A(n22897), .B(n22896), .Z(n22936) );
  NAND U23501 ( .A(b[0]), .B(a[557]), .Z(n22898) );
  XNOR U23502 ( .A(b[1]), .B(n22898), .Z(n22900) );
  NAND U23503 ( .A(n94), .B(a[556]), .Z(n22899) );
  AND U23504 ( .A(n22900), .B(n22899), .Z(n22953) );
  XOR U23505 ( .A(a[553]), .B(n42197), .Z(n22942) );
  NANDN U23506 ( .A(n22942), .B(n42173), .Z(n22903) );
  NANDN U23507 ( .A(n22901), .B(n42172), .Z(n22902) );
  NAND U23508 ( .A(n22903), .B(n22902), .Z(n22951) );
  NAND U23509 ( .A(b[7]), .B(a[549]), .Z(n22952) );
  XNOR U23510 ( .A(n22951), .B(n22952), .Z(n22954) );
  XOR U23511 ( .A(n22953), .B(n22954), .Z(n22960) );
  NANDN U23512 ( .A(n22904), .B(n42093), .Z(n22906) );
  XOR U23513 ( .A(n42134), .B(a[555]), .Z(n22945) );
  NANDN U23514 ( .A(n22945), .B(n42095), .Z(n22905) );
  NAND U23515 ( .A(n22906), .B(n22905), .Z(n22958) );
  NANDN U23516 ( .A(n22907), .B(n42231), .Z(n22909) );
  XOR U23517 ( .A(n208), .B(a[551]), .Z(n22948) );
  NANDN U23518 ( .A(n22948), .B(n42234), .Z(n22908) );
  AND U23519 ( .A(n22909), .B(n22908), .Z(n22957) );
  XNOR U23520 ( .A(n22958), .B(n22957), .Z(n22959) );
  XNOR U23521 ( .A(n22960), .B(n22959), .Z(n22964) );
  NANDN U23522 ( .A(n22911), .B(n22910), .Z(n22915) );
  NAND U23523 ( .A(n22913), .B(n22912), .Z(n22914) );
  AND U23524 ( .A(n22915), .B(n22914), .Z(n22963) );
  XOR U23525 ( .A(n22964), .B(n22963), .Z(n22965) );
  NANDN U23526 ( .A(n22917), .B(n22916), .Z(n22921) );
  NANDN U23527 ( .A(n22919), .B(n22918), .Z(n22920) );
  NAND U23528 ( .A(n22921), .B(n22920), .Z(n22966) );
  XOR U23529 ( .A(n22965), .B(n22966), .Z(n22933) );
  OR U23530 ( .A(n22923), .B(n22922), .Z(n22927) );
  NANDN U23531 ( .A(n22925), .B(n22924), .Z(n22926) );
  NAND U23532 ( .A(n22927), .B(n22926), .Z(n22934) );
  XNOR U23533 ( .A(n22933), .B(n22934), .Z(n22935) );
  XNOR U23534 ( .A(n22936), .B(n22935), .Z(n22969) );
  XNOR U23535 ( .A(n22969), .B(sreg[1573]), .Z(n22971) );
  NAND U23536 ( .A(n22928), .B(sreg[1572]), .Z(n22932) );
  OR U23537 ( .A(n22930), .B(n22929), .Z(n22931) );
  AND U23538 ( .A(n22932), .B(n22931), .Z(n22970) );
  XOR U23539 ( .A(n22971), .B(n22970), .Z(c[1573]) );
  NANDN U23540 ( .A(n22934), .B(n22933), .Z(n22938) );
  NAND U23541 ( .A(n22936), .B(n22935), .Z(n22937) );
  NAND U23542 ( .A(n22938), .B(n22937), .Z(n22977) );
  NAND U23543 ( .A(b[0]), .B(a[558]), .Z(n22939) );
  XNOR U23544 ( .A(b[1]), .B(n22939), .Z(n22941) );
  NAND U23545 ( .A(n94), .B(a[557]), .Z(n22940) );
  AND U23546 ( .A(n22941), .B(n22940), .Z(n22994) );
  XOR U23547 ( .A(a[554]), .B(n42197), .Z(n22983) );
  NANDN U23548 ( .A(n22983), .B(n42173), .Z(n22944) );
  NANDN U23549 ( .A(n22942), .B(n42172), .Z(n22943) );
  NAND U23550 ( .A(n22944), .B(n22943), .Z(n22992) );
  NAND U23551 ( .A(b[7]), .B(a[550]), .Z(n22993) );
  XNOR U23552 ( .A(n22992), .B(n22993), .Z(n22995) );
  XOR U23553 ( .A(n22994), .B(n22995), .Z(n23001) );
  NANDN U23554 ( .A(n22945), .B(n42093), .Z(n22947) );
  XOR U23555 ( .A(n42134), .B(a[556]), .Z(n22986) );
  NANDN U23556 ( .A(n22986), .B(n42095), .Z(n22946) );
  NAND U23557 ( .A(n22947), .B(n22946), .Z(n22999) );
  NANDN U23558 ( .A(n22948), .B(n42231), .Z(n22950) );
  XOR U23559 ( .A(n208), .B(a[552]), .Z(n22989) );
  NANDN U23560 ( .A(n22989), .B(n42234), .Z(n22949) );
  AND U23561 ( .A(n22950), .B(n22949), .Z(n22998) );
  XNOR U23562 ( .A(n22999), .B(n22998), .Z(n23000) );
  XNOR U23563 ( .A(n23001), .B(n23000), .Z(n23005) );
  NANDN U23564 ( .A(n22952), .B(n22951), .Z(n22956) );
  NAND U23565 ( .A(n22954), .B(n22953), .Z(n22955) );
  AND U23566 ( .A(n22956), .B(n22955), .Z(n23004) );
  XOR U23567 ( .A(n23005), .B(n23004), .Z(n23006) );
  NANDN U23568 ( .A(n22958), .B(n22957), .Z(n22962) );
  NANDN U23569 ( .A(n22960), .B(n22959), .Z(n22961) );
  NAND U23570 ( .A(n22962), .B(n22961), .Z(n23007) );
  XOR U23571 ( .A(n23006), .B(n23007), .Z(n22974) );
  OR U23572 ( .A(n22964), .B(n22963), .Z(n22968) );
  NANDN U23573 ( .A(n22966), .B(n22965), .Z(n22967) );
  NAND U23574 ( .A(n22968), .B(n22967), .Z(n22975) );
  XNOR U23575 ( .A(n22974), .B(n22975), .Z(n22976) );
  XNOR U23576 ( .A(n22977), .B(n22976), .Z(n23010) );
  XNOR U23577 ( .A(n23010), .B(sreg[1574]), .Z(n23012) );
  NAND U23578 ( .A(n22969), .B(sreg[1573]), .Z(n22973) );
  OR U23579 ( .A(n22971), .B(n22970), .Z(n22972) );
  AND U23580 ( .A(n22973), .B(n22972), .Z(n23011) );
  XOR U23581 ( .A(n23012), .B(n23011), .Z(c[1574]) );
  NANDN U23582 ( .A(n22975), .B(n22974), .Z(n22979) );
  NAND U23583 ( .A(n22977), .B(n22976), .Z(n22978) );
  NAND U23584 ( .A(n22979), .B(n22978), .Z(n23018) );
  NAND U23585 ( .A(b[0]), .B(a[559]), .Z(n22980) );
  XNOR U23586 ( .A(b[1]), .B(n22980), .Z(n22982) );
  NAND U23587 ( .A(n94), .B(a[558]), .Z(n22981) );
  AND U23588 ( .A(n22982), .B(n22981), .Z(n23035) );
  XOR U23589 ( .A(a[555]), .B(n42197), .Z(n23024) );
  NANDN U23590 ( .A(n23024), .B(n42173), .Z(n22985) );
  NANDN U23591 ( .A(n22983), .B(n42172), .Z(n22984) );
  NAND U23592 ( .A(n22985), .B(n22984), .Z(n23033) );
  NAND U23593 ( .A(b[7]), .B(a[551]), .Z(n23034) );
  XNOR U23594 ( .A(n23033), .B(n23034), .Z(n23036) );
  XOR U23595 ( .A(n23035), .B(n23036), .Z(n23042) );
  NANDN U23596 ( .A(n22986), .B(n42093), .Z(n22988) );
  XOR U23597 ( .A(n42134), .B(a[557]), .Z(n23027) );
  NANDN U23598 ( .A(n23027), .B(n42095), .Z(n22987) );
  NAND U23599 ( .A(n22988), .B(n22987), .Z(n23040) );
  NANDN U23600 ( .A(n22989), .B(n42231), .Z(n22991) );
  XOR U23601 ( .A(n208), .B(a[553]), .Z(n23030) );
  NANDN U23602 ( .A(n23030), .B(n42234), .Z(n22990) );
  AND U23603 ( .A(n22991), .B(n22990), .Z(n23039) );
  XNOR U23604 ( .A(n23040), .B(n23039), .Z(n23041) );
  XNOR U23605 ( .A(n23042), .B(n23041), .Z(n23046) );
  NANDN U23606 ( .A(n22993), .B(n22992), .Z(n22997) );
  NAND U23607 ( .A(n22995), .B(n22994), .Z(n22996) );
  AND U23608 ( .A(n22997), .B(n22996), .Z(n23045) );
  XOR U23609 ( .A(n23046), .B(n23045), .Z(n23047) );
  NANDN U23610 ( .A(n22999), .B(n22998), .Z(n23003) );
  NANDN U23611 ( .A(n23001), .B(n23000), .Z(n23002) );
  NAND U23612 ( .A(n23003), .B(n23002), .Z(n23048) );
  XOR U23613 ( .A(n23047), .B(n23048), .Z(n23015) );
  OR U23614 ( .A(n23005), .B(n23004), .Z(n23009) );
  NANDN U23615 ( .A(n23007), .B(n23006), .Z(n23008) );
  NAND U23616 ( .A(n23009), .B(n23008), .Z(n23016) );
  XNOR U23617 ( .A(n23015), .B(n23016), .Z(n23017) );
  XNOR U23618 ( .A(n23018), .B(n23017), .Z(n23051) );
  XNOR U23619 ( .A(n23051), .B(sreg[1575]), .Z(n23053) );
  NAND U23620 ( .A(n23010), .B(sreg[1574]), .Z(n23014) );
  OR U23621 ( .A(n23012), .B(n23011), .Z(n23013) );
  AND U23622 ( .A(n23014), .B(n23013), .Z(n23052) );
  XOR U23623 ( .A(n23053), .B(n23052), .Z(c[1575]) );
  NANDN U23624 ( .A(n23016), .B(n23015), .Z(n23020) );
  NAND U23625 ( .A(n23018), .B(n23017), .Z(n23019) );
  NAND U23626 ( .A(n23020), .B(n23019), .Z(n23059) );
  NAND U23627 ( .A(b[0]), .B(a[560]), .Z(n23021) );
  XNOR U23628 ( .A(b[1]), .B(n23021), .Z(n23023) );
  NAND U23629 ( .A(n95), .B(a[559]), .Z(n23022) );
  AND U23630 ( .A(n23023), .B(n23022), .Z(n23076) );
  XOR U23631 ( .A(a[556]), .B(n42197), .Z(n23065) );
  NANDN U23632 ( .A(n23065), .B(n42173), .Z(n23026) );
  NANDN U23633 ( .A(n23024), .B(n42172), .Z(n23025) );
  NAND U23634 ( .A(n23026), .B(n23025), .Z(n23074) );
  NAND U23635 ( .A(b[7]), .B(a[552]), .Z(n23075) );
  XNOR U23636 ( .A(n23074), .B(n23075), .Z(n23077) );
  XOR U23637 ( .A(n23076), .B(n23077), .Z(n23083) );
  NANDN U23638 ( .A(n23027), .B(n42093), .Z(n23029) );
  XOR U23639 ( .A(n42134), .B(a[558]), .Z(n23068) );
  NANDN U23640 ( .A(n23068), .B(n42095), .Z(n23028) );
  NAND U23641 ( .A(n23029), .B(n23028), .Z(n23081) );
  NANDN U23642 ( .A(n23030), .B(n42231), .Z(n23032) );
  XOR U23643 ( .A(n208), .B(a[554]), .Z(n23071) );
  NANDN U23644 ( .A(n23071), .B(n42234), .Z(n23031) );
  AND U23645 ( .A(n23032), .B(n23031), .Z(n23080) );
  XNOR U23646 ( .A(n23081), .B(n23080), .Z(n23082) );
  XNOR U23647 ( .A(n23083), .B(n23082), .Z(n23087) );
  NANDN U23648 ( .A(n23034), .B(n23033), .Z(n23038) );
  NAND U23649 ( .A(n23036), .B(n23035), .Z(n23037) );
  AND U23650 ( .A(n23038), .B(n23037), .Z(n23086) );
  XOR U23651 ( .A(n23087), .B(n23086), .Z(n23088) );
  NANDN U23652 ( .A(n23040), .B(n23039), .Z(n23044) );
  NANDN U23653 ( .A(n23042), .B(n23041), .Z(n23043) );
  NAND U23654 ( .A(n23044), .B(n23043), .Z(n23089) );
  XOR U23655 ( .A(n23088), .B(n23089), .Z(n23056) );
  OR U23656 ( .A(n23046), .B(n23045), .Z(n23050) );
  NANDN U23657 ( .A(n23048), .B(n23047), .Z(n23049) );
  NAND U23658 ( .A(n23050), .B(n23049), .Z(n23057) );
  XNOR U23659 ( .A(n23056), .B(n23057), .Z(n23058) );
  XNOR U23660 ( .A(n23059), .B(n23058), .Z(n23092) );
  XNOR U23661 ( .A(n23092), .B(sreg[1576]), .Z(n23094) );
  NAND U23662 ( .A(n23051), .B(sreg[1575]), .Z(n23055) );
  OR U23663 ( .A(n23053), .B(n23052), .Z(n23054) );
  AND U23664 ( .A(n23055), .B(n23054), .Z(n23093) );
  XOR U23665 ( .A(n23094), .B(n23093), .Z(c[1576]) );
  NANDN U23666 ( .A(n23057), .B(n23056), .Z(n23061) );
  NAND U23667 ( .A(n23059), .B(n23058), .Z(n23060) );
  NAND U23668 ( .A(n23061), .B(n23060), .Z(n23100) );
  NAND U23669 ( .A(b[0]), .B(a[561]), .Z(n23062) );
  XNOR U23670 ( .A(b[1]), .B(n23062), .Z(n23064) );
  NAND U23671 ( .A(n95), .B(a[560]), .Z(n23063) );
  AND U23672 ( .A(n23064), .B(n23063), .Z(n23117) );
  XOR U23673 ( .A(a[557]), .B(n42197), .Z(n23106) );
  NANDN U23674 ( .A(n23106), .B(n42173), .Z(n23067) );
  NANDN U23675 ( .A(n23065), .B(n42172), .Z(n23066) );
  NAND U23676 ( .A(n23067), .B(n23066), .Z(n23115) );
  NAND U23677 ( .A(b[7]), .B(a[553]), .Z(n23116) );
  XNOR U23678 ( .A(n23115), .B(n23116), .Z(n23118) );
  XOR U23679 ( .A(n23117), .B(n23118), .Z(n23124) );
  NANDN U23680 ( .A(n23068), .B(n42093), .Z(n23070) );
  XOR U23681 ( .A(n42134), .B(a[559]), .Z(n23109) );
  NANDN U23682 ( .A(n23109), .B(n42095), .Z(n23069) );
  NAND U23683 ( .A(n23070), .B(n23069), .Z(n23122) );
  NANDN U23684 ( .A(n23071), .B(n42231), .Z(n23073) );
  XOR U23685 ( .A(n208), .B(a[555]), .Z(n23112) );
  NANDN U23686 ( .A(n23112), .B(n42234), .Z(n23072) );
  AND U23687 ( .A(n23073), .B(n23072), .Z(n23121) );
  XNOR U23688 ( .A(n23122), .B(n23121), .Z(n23123) );
  XNOR U23689 ( .A(n23124), .B(n23123), .Z(n23128) );
  NANDN U23690 ( .A(n23075), .B(n23074), .Z(n23079) );
  NAND U23691 ( .A(n23077), .B(n23076), .Z(n23078) );
  AND U23692 ( .A(n23079), .B(n23078), .Z(n23127) );
  XOR U23693 ( .A(n23128), .B(n23127), .Z(n23129) );
  NANDN U23694 ( .A(n23081), .B(n23080), .Z(n23085) );
  NANDN U23695 ( .A(n23083), .B(n23082), .Z(n23084) );
  NAND U23696 ( .A(n23085), .B(n23084), .Z(n23130) );
  XOR U23697 ( .A(n23129), .B(n23130), .Z(n23097) );
  OR U23698 ( .A(n23087), .B(n23086), .Z(n23091) );
  NANDN U23699 ( .A(n23089), .B(n23088), .Z(n23090) );
  NAND U23700 ( .A(n23091), .B(n23090), .Z(n23098) );
  XNOR U23701 ( .A(n23097), .B(n23098), .Z(n23099) );
  XNOR U23702 ( .A(n23100), .B(n23099), .Z(n23133) );
  XNOR U23703 ( .A(n23133), .B(sreg[1577]), .Z(n23135) );
  NAND U23704 ( .A(n23092), .B(sreg[1576]), .Z(n23096) );
  OR U23705 ( .A(n23094), .B(n23093), .Z(n23095) );
  AND U23706 ( .A(n23096), .B(n23095), .Z(n23134) );
  XOR U23707 ( .A(n23135), .B(n23134), .Z(c[1577]) );
  NANDN U23708 ( .A(n23098), .B(n23097), .Z(n23102) );
  NAND U23709 ( .A(n23100), .B(n23099), .Z(n23101) );
  NAND U23710 ( .A(n23102), .B(n23101), .Z(n23141) );
  NAND U23711 ( .A(b[0]), .B(a[562]), .Z(n23103) );
  XNOR U23712 ( .A(b[1]), .B(n23103), .Z(n23105) );
  NAND U23713 ( .A(n95), .B(a[561]), .Z(n23104) );
  AND U23714 ( .A(n23105), .B(n23104), .Z(n23158) );
  XOR U23715 ( .A(a[558]), .B(n42197), .Z(n23147) );
  NANDN U23716 ( .A(n23147), .B(n42173), .Z(n23108) );
  NANDN U23717 ( .A(n23106), .B(n42172), .Z(n23107) );
  NAND U23718 ( .A(n23108), .B(n23107), .Z(n23156) );
  NAND U23719 ( .A(b[7]), .B(a[554]), .Z(n23157) );
  XNOR U23720 ( .A(n23156), .B(n23157), .Z(n23159) );
  XOR U23721 ( .A(n23158), .B(n23159), .Z(n23165) );
  NANDN U23722 ( .A(n23109), .B(n42093), .Z(n23111) );
  XOR U23723 ( .A(n42134), .B(a[560]), .Z(n23150) );
  NANDN U23724 ( .A(n23150), .B(n42095), .Z(n23110) );
  NAND U23725 ( .A(n23111), .B(n23110), .Z(n23163) );
  NANDN U23726 ( .A(n23112), .B(n42231), .Z(n23114) );
  XOR U23727 ( .A(n208), .B(a[556]), .Z(n23153) );
  NANDN U23728 ( .A(n23153), .B(n42234), .Z(n23113) );
  AND U23729 ( .A(n23114), .B(n23113), .Z(n23162) );
  XNOR U23730 ( .A(n23163), .B(n23162), .Z(n23164) );
  XNOR U23731 ( .A(n23165), .B(n23164), .Z(n23169) );
  NANDN U23732 ( .A(n23116), .B(n23115), .Z(n23120) );
  NAND U23733 ( .A(n23118), .B(n23117), .Z(n23119) );
  AND U23734 ( .A(n23120), .B(n23119), .Z(n23168) );
  XOR U23735 ( .A(n23169), .B(n23168), .Z(n23170) );
  NANDN U23736 ( .A(n23122), .B(n23121), .Z(n23126) );
  NANDN U23737 ( .A(n23124), .B(n23123), .Z(n23125) );
  NAND U23738 ( .A(n23126), .B(n23125), .Z(n23171) );
  XOR U23739 ( .A(n23170), .B(n23171), .Z(n23138) );
  OR U23740 ( .A(n23128), .B(n23127), .Z(n23132) );
  NANDN U23741 ( .A(n23130), .B(n23129), .Z(n23131) );
  NAND U23742 ( .A(n23132), .B(n23131), .Z(n23139) );
  XNOR U23743 ( .A(n23138), .B(n23139), .Z(n23140) );
  XNOR U23744 ( .A(n23141), .B(n23140), .Z(n23174) );
  XNOR U23745 ( .A(n23174), .B(sreg[1578]), .Z(n23176) );
  NAND U23746 ( .A(n23133), .B(sreg[1577]), .Z(n23137) );
  OR U23747 ( .A(n23135), .B(n23134), .Z(n23136) );
  AND U23748 ( .A(n23137), .B(n23136), .Z(n23175) );
  XOR U23749 ( .A(n23176), .B(n23175), .Z(c[1578]) );
  NANDN U23750 ( .A(n23139), .B(n23138), .Z(n23143) );
  NAND U23751 ( .A(n23141), .B(n23140), .Z(n23142) );
  NAND U23752 ( .A(n23143), .B(n23142), .Z(n23182) );
  NAND U23753 ( .A(b[0]), .B(a[563]), .Z(n23144) );
  XNOR U23754 ( .A(b[1]), .B(n23144), .Z(n23146) );
  NAND U23755 ( .A(n95), .B(a[562]), .Z(n23145) );
  AND U23756 ( .A(n23146), .B(n23145), .Z(n23199) );
  XOR U23757 ( .A(a[559]), .B(n42197), .Z(n23188) );
  NANDN U23758 ( .A(n23188), .B(n42173), .Z(n23149) );
  NANDN U23759 ( .A(n23147), .B(n42172), .Z(n23148) );
  NAND U23760 ( .A(n23149), .B(n23148), .Z(n23197) );
  NAND U23761 ( .A(b[7]), .B(a[555]), .Z(n23198) );
  XNOR U23762 ( .A(n23197), .B(n23198), .Z(n23200) );
  XOR U23763 ( .A(n23199), .B(n23200), .Z(n23206) );
  NANDN U23764 ( .A(n23150), .B(n42093), .Z(n23152) );
  XOR U23765 ( .A(n42134), .B(a[561]), .Z(n23191) );
  NANDN U23766 ( .A(n23191), .B(n42095), .Z(n23151) );
  NAND U23767 ( .A(n23152), .B(n23151), .Z(n23204) );
  NANDN U23768 ( .A(n23153), .B(n42231), .Z(n23155) );
  XOR U23769 ( .A(n208), .B(a[557]), .Z(n23194) );
  NANDN U23770 ( .A(n23194), .B(n42234), .Z(n23154) );
  AND U23771 ( .A(n23155), .B(n23154), .Z(n23203) );
  XNOR U23772 ( .A(n23204), .B(n23203), .Z(n23205) );
  XNOR U23773 ( .A(n23206), .B(n23205), .Z(n23210) );
  NANDN U23774 ( .A(n23157), .B(n23156), .Z(n23161) );
  NAND U23775 ( .A(n23159), .B(n23158), .Z(n23160) );
  AND U23776 ( .A(n23161), .B(n23160), .Z(n23209) );
  XOR U23777 ( .A(n23210), .B(n23209), .Z(n23211) );
  NANDN U23778 ( .A(n23163), .B(n23162), .Z(n23167) );
  NANDN U23779 ( .A(n23165), .B(n23164), .Z(n23166) );
  NAND U23780 ( .A(n23167), .B(n23166), .Z(n23212) );
  XOR U23781 ( .A(n23211), .B(n23212), .Z(n23179) );
  OR U23782 ( .A(n23169), .B(n23168), .Z(n23173) );
  NANDN U23783 ( .A(n23171), .B(n23170), .Z(n23172) );
  NAND U23784 ( .A(n23173), .B(n23172), .Z(n23180) );
  XNOR U23785 ( .A(n23179), .B(n23180), .Z(n23181) );
  XNOR U23786 ( .A(n23182), .B(n23181), .Z(n23215) );
  XNOR U23787 ( .A(n23215), .B(sreg[1579]), .Z(n23217) );
  NAND U23788 ( .A(n23174), .B(sreg[1578]), .Z(n23178) );
  OR U23789 ( .A(n23176), .B(n23175), .Z(n23177) );
  AND U23790 ( .A(n23178), .B(n23177), .Z(n23216) );
  XOR U23791 ( .A(n23217), .B(n23216), .Z(c[1579]) );
  NANDN U23792 ( .A(n23180), .B(n23179), .Z(n23184) );
  NAND U23793 ( .A(n23182), .B(n23181), .Z(n23183) );
  NAND U23794 ( .A(n23184), .B(n23183), .Z(n23223) );
  NAND U23795 ( .A(b[0]), .B(a[564]), .Z(n23185) );
  XNOR U23796 ( .A(b[1]), .B(n23185), .Z(n23187) );
  NAND U23797 ( .A(n95), .B(a[563]), .Z(n23186) );
  AND U23798 ( .A(n23187), .B(n23186), .Z(n23240) );
  XOR U23799 ( .A(a[560]), .B(n42197), .Z(n23229) );
  NANDN U23800 ( .A(n23229), .B(n42173), .Z(n23190) );
  NANDN U23801 ( .A(n23188), .B(n42172), .Z(n23189) );
  NAND U23802 ( .A(n23190), .B(n23189), .Z(n23238) );
  NAND U23803 ( .A(b[7]), .B(a[556]), .Z(n23239) );
  XNOR U23804 ( .A(n23238), .B(n23239), .Z(n23241) );
  XOR U23805 ( .A(n23240), .B(n23241), .Z(n23247) );
  NANDN U23806 ( .A(n23191), .B(n42093), .Z(n23193) );
  XOR U23807 ( .A(n42134), .B(a[562]), .Z(n23232) );
  NANDN U23808 ( .A(n23232), .B(n42095), .Z(n23192) );
  NAND U23809 ( .A(n23193), .B(n23192), .Z(n23245) );
  NANDN U23810 ( .A(n23194), .B(n42231), .Z(n23196) );
  XOR U23811 ( .A(n208), .B(a[558]), .Z(n23235) );
  NANDN U23812 ( .A(n23235), .B(n42234), .Z(n23195) );
  AND U23813 ( .A(n23196), .B(n23195), .Z(n23244) );
  XNOR U23814 ( .A(n23245), .B(n23244), .Z(n23246) );
  XNOR U23815 ( .A(n23247), .B(n23246), .Z(n23251) );
  NANDN U23816 ( .A(n23198), .B(n23197), .Z(n23202) );
  NAND U23817 ( .A(n23200), .B(n23199), .Z(n23201) );
  AND U23818 ( .A(n23202), .B(n23201), .Z(n23250) );
  XOR U23819 ( .A(n23251), .B(n23250), .Z(n23252) );
  NANDN U23820 ( .A(n23204), .B(n23203), .Z(n23208) );
  NANDN U23821 ( .A(n23206), .B(n23205), .Z(n23207) );
  NAND U23822 ( .A(n23208), .B(n23207), .Z(n23253) );
  XOR U23823 ( .A(n23252), .B(n23253), .Z(n23220) );
  OR U23824 ( .A(n23210), .B(n23209), .Z(n23214) );
  NANDN U23825 ( .A(n23212), .B(n23211), .Z(n23213) );
  NAND U23826 ( .A(n23214), .B(n23213), .Z(n23221) );
  XNOR U23827 ( .A(n23220), .B(n23221), .Z(n23222) );
  XNOR U23828 ( .A(n23223), .B(n23222), .Z(n23256) );
  XNOR U23829 ( .A(n23256), .B(sreg[1580]), .Z(n23258) );
  NAND U23830 ( .A(n23215), .B(sreg[1579]), .Z(n23219) );
  OR U23831 ( .A(n23217), .B(n23216), .Z(n23218) );
  AND U23832 ( .A(n23219), .B(n23218), .Z(n23257) );
  XOR U23833 ( .A(n23258), .B(n23257), .Z(c[1580]) );
  NANDN U23834 ( .A(n23221), .B(n23220), .Z(n23225) );
  NAND U23835 ( .A(n23223), .B(n23222), .Z(n23224) );
  NAND U23836 ( .A(n23225), .B(n23224), .Z(n23264) );
  NAND U23837 ( .A(b[0]), .B(a[565]), .Z(n23226) );
  XNOR U23838 ( .A(b[1]), .B(n23226), .Z(n23228) );
  NAND U23839 ( .A(n95), .B(a[564]), .Z(n23227) );
  AND U23840 ( .A(n23228), .B(n23227), .Z(n23281) );
  XOR U23841 ( .A(a[561]), .B(n42197), .Z(n23270) );
  NANDN U23842 ( .A(n23270), .B(n42173), .Z(n23231) );
  NANDN U23843 ( .A(n23229), .B(n42172), .Z(n23230) );
  NAND U23844 ( .A(n23231), .B(n23230), .Z(n23279) );
  NAND U23845 ( .A(b[7]), .B(a[557]), .Z(n23280) );
  XNOR U23846 ( .A(n23279), .B(n23280), .Z(n23282) );
  XOR U23847 ( .A(n23281), .B(n23282), .Z(n23288) );
  NANDN U23848 ( .A(n23232), .B(n42093), .Z(n23234) );
  XOR U23849 ( .A(n42134), .B(a[563]), .Z(n23273) );
  NANDN U23850 ( .A(n23273), .B(n42095), .Z(n23233) );
  NAND U23851 ( .A(n23234), .B(n23233), .Z(n23286) );
  NANDN U23852 ( .A(n23235), .B(n42231), .Z(n23237) );
  XOR U23853 ( .A(n208), .B(a[559]), .Z(n23276) );
  NANDN U23854 ( .A(n23276), .B(n42234), .Z(n23236) );
  AND U23855 ( .A(n23237), .B(n23236), .Z(n23285) );
  XNOR U23856 ( .A(n23286), .B(n23285), .Z(n23287) );
  XNOR U23857 ( .A(n23288), .B(n23287), .Z(n23292) );
  NANDN U23858 ( .A(n23239), .B(n23238), .Z(n23243) );
  NAND U23859 ( .A(n23241), .B(n23240), .Z(n23242) );
  AND U23860 ( .A(n23243), .B(n23242), .Z(n23291) );
  XOR U23861 ( .A(n23292), .B(n23291), .Z(n23293) );
  NANDN U23862 ( .A(n23245), .B(n23244), .Z(n23249) );
  NANDN U23863 ( .A(n23247), .B(n23246), .Z(n23248) );
  NAND U23864 ( .A(n23249), .B(n23248), .Z(n23294) );
  XOR U23865 ( .A(n23293), .B(n23294), .Z(n23261) );
  OR U23866 ( .A(n23251), .B(n23250), .Z(n23255) );
  NANDN U23867 ( .A(n23253), .B(n23252), .Z(n23254) );
  NAND U23868 ( .A(n23255), .B(n23254), .Z(n23262) );
  XNOR U23869 ( .A(n23261), .B(n23262), .Z(n23263) );
  XNOR U23870 ( .A(n23264), .B(n23263), .Z(n23297) );
  XNOR U23871 ( .A(n23297), .B(sreg[1581]), .Z(n23299) );
  NAND U23872 ( .A(n23256), .B(sreg[1580]), .Z(n23260) );
  OR U23873 ( .A(n23258), .B(n23257), .Z(n23259) );
  AND U23874 ( .A(n23260), .B(n23259), .Z(n23298) );
  XOR U23875 ( .A(n23299), .B(n23298), .Z(c[1581]) );
  NANDN U23876 ( .A(n23262), .B(n23261), .Z(n23266) );
  NAND U23877 ( .A(n23264), .B(n23263), .Z(n23265) );
  NAND U23878 ( .A(n23266), .B(n23265), .Z(n23305) );
  NAND U23879 ( .A(b[0]), .B(a[566]), .Z(n23267) );
  XNOR U23880 ( .A(b[1]), .B(n23267), .Z(n23269) );
  NAND U23881 ( .A(n95), .B(a[565]), .Z(n23268) );
  AND U23882 ( .A(n23269), .B(n23268), .Z(n23322) );
  XOR U23883 ( .A(a[562]), .B(n42197), .Z(n23311) );
  NANDN U23884 ( .A(n23311), .B(n42173), .Z(n23272) );
  NANDN U23885 ( .A(n23270), .B(n42172), .Z(n23271) );
  NAND U23886 ( .A(n23272), .B(n23271), .Z(n23320) );
  NAND U23887 ( .A(b[7]), .B(a[558]), .Z(n23321) );
  XNOR U23888 ( .A(n23320), .B(n23321), .Z(n23323) );
  XOR U23889 ( .A(n23322), .B(n23323), .Z(n23329) );
  NANDN U23890 ( .A(n23273), .B(n42093), .Z(n23275) );
  XOR U23891 ( .A(n42134), .B(a[564]), .Z(n23314) );
  NANDN U23892 ( .A(n23314), .B(n42095), .Z(n23274) );
  NAND U23893 ( .A(n23275), .B(n23274), .Z(n23327) );
  NANDN U23894 ( .A(n23276), .B(n42231), .Z(n23278) );
  XOR U23895 ( .A(n208), .B(a[560]), .Z(n23317) );
  NANDN U23896 ( .A(n23317), .B(n42234), .Z(n23277) );
  AND U23897 ( .A(n23278), .B(n23277), .Z(n23326) );
  XNOR U23898 ( .A(n23327), .B(n23326), .Z(n23328) );
  XNOR U23899 ( .A(n23329), .B(n23328), .Z(n23333) );
  NANDN U23900 ( .A(n23280), .B(n23279), .Z(n23284) );
  NAND U23901 ( .A(n23282), .B(n23281), .Z(n23283) );
  AND U23902 ( .A(n23284), .B(n23283), .Z(n23332) );
  XOR U23903 ( .A(n23333), .B(n23332), .Z(n23334) );
  NANDN U23904 ( .A(n23286), .B(n23285), .Z(n23290) );
  NANDN U23905 ( .A(n23288), .B(n23287), .Z(n23289) );
  NAND U23906 ( .A(n23290), .B(n23289), .Z(n23335) );
  XOR U23907 ( .A(n23334), .B(n23335), .Z(n23302) );
  OR U23908 ( .A(n23292), .B(n23291), .Z(n23296) );
  NANDN U23909 ( .A(n23294), .B(n23293), .Z(n23295) );
  NAND U23910 ( .A(n23296), .B(n23295), .Z(n23303) );
  XNOR U23911 ( .A(n23302), .B(n23303), .Z(n23304) );
  XNOR U23912 ( .A(n23305), .B(n23304), .Z(n23338) );
  XNOR U23913 ( .A(n23338), .B(sreg[1582]), .Z(n23340) );
  NAND U23914 ( .A(n23297), .B(sreg[1581]), .Z(n23301) );
  OR U23915 ( .A(n23299), .B(n23298), .Z(n23300) );
  AND U23916 ( .A(n23301), .B(n23300), .Z(n23339) );
  XOR U23917 ( .A(n23340), .B(n23339), .Z(c[1582]) );
  NANDN U23918 ( .A(n23303), .B(n23302), .Z(n23307) );
  NAND U23919 ( .A(n23305), .B(n23304), .Z(n23306) );
  NAND U23920 ( .A(n23307), .B(n23306), .Z(n23346) );
  NAND U23921 ( .A(b[0]), .B(a[567]), .Z(n23308) );
  XNOR U23922 ( .A(b[1]), .B(n23308), .Z(n23310) );
  NAND U23923 ( .A(n96), .B(a[566]), .Z(n23309) );
  AND U23924 ( .A(n23310), .B(n23309), .Z(n23363) );
  XOR U23925 ( .A(a[563]), .B(n42197), .Z(n23352) );
  NANDN U23926 ( .A(n23352), .B(n42173), .Z(n23313) );
  NANDN U23927 ( .A(n23311), .B(n42172), .Z(n23312) );
  NAND U23928 ( .A(n23313), .B(n23312), .Z(n23361) );
  NAND U23929 ( .A(b[7]), .B(a[559]), .Z(n23362) );
  XNOR U23930 ( .A(n23361), .B(n23362), .Z(n23364) );
  XOR U23931 ( .A(n23363), .B(n23364), .Z(n23370) );
  NANDN U23932 ( .A(n23314), .B(n42093), .Z(n23316) );
  XOR U23933 ( .A(n42134), .B(a[565]), .Z(n23355) );
  NANDN U23934 ( .A(n23355), .B(n42095), .Z(n23315) );
  NAND U23935 ( .A(n23316), .B(n23315), .Z(n23368) );
  NANDN U23936 ( .A(n23317), .B(n42231), .Z(n23319) );
  XOR U23937 ( .A(n208), .B(a[561]), .Z(n23358) );
  NANDN U23938 ( .A(n23358), .B(n42234), .Z(n23318) );
  AND U23939 ( .A(n23319), .B(n23318), .Z(n23367) );
  XNOR U23940 ( .A(n23368), .B(n23367), .Z(n23369) );
  XNOR U23941 ( .A(n23370), .B(n23369), .Z(n23374) );
  NANDN U23942 ( .A(n23321), .B(n23320), .Z(n23325) );
  NAND U23943 ( .A(n23323), .B(n23322), .Z(n23324) );
  AND U23944 ( .A(n23325), .B(n23324), .Z(n23373) );
  XOR U23945 ( .A(n23374), .B(n23373), .Z(n23375) );
  NANDN U23946 ( .A(n23327), .B(n23326), .Z(n23331) );
  NANDN U23947 ( .A(n23329), .B(n23328), .Z(n23330) );
  NAND U23948 ( .A(n23331), .B(n23330), .Z(n23376) );
  XOR U23949 ( .A(n23375), .B(n23376), .Z(n23343) );
  OR U23950 ( .A(n23333), .B(n23332), .Z(n23337) );
  NANDN U23951 ( .A(n23335), .B(n23334), .Z(n23336) );
  NAND U23952 ( .A(n23337), .B(n23336), .Z(n23344) );
  XNOR U23953 ( .A(n23343), .B(n23344), .Z(n23345) );
  XNOR U23954 ( .A(n23346), .B(n23345), .Z(n23379) );
  XNOR U23955 ( .A(n23379), .B(sreg[1583]), .Z(n23381) );
  NAND U23956 ( .A(n23338), .B(sreg[1582]), .Z(n23342) );
  OR U23957 ( .A(n23340), .B(n23339), .Z(n23341) );
  AND U23958 ( .A(n23342), .B(n23341), .Z(n23380) );
  XOR U23959 ( .A(n23381), .B(n23380), .Z(c[1583]) );
  NANDN U23960 ( .A(n23344), .B(n23343), .Z(n23348) );
  NAND U23961 ( .A(n23346), .B(n23345), .Z(n23347) );
  NAND U23962 ( .A(n23348), .B(n23347), .Z(n23387) );
  NAND U23963 ( .A(b[0]), .B(a[568]), .Z(n23349) );
  XNOR U23964 ( .A(b[1]), .B(n23349), .Z(n23351) );
  NAND U23965 ( .A(n96), .B(a[567]), .Z(n23350) );
  AND U23966 ( .A(n23351), .B(n23350), .Z(n23404) );
  XOR U23967 ( .A(a[564]), .B(n42197), .Z(n23393) );
  NANDN U23968 ( .A(n23393), .B(n42173), .Z(n23354) );
  NANDN U23969 ( .A(n23352), .B(n42172), .Z(n23353) );
  NAND U23970 ( .A(n23354), .B(n23353), .Z(n23402) );
  NAND U23971 ( .A(b[7]), .B(a[560]), .Z(n23403) );
  XNOR U23972 ( .A(n23402), .B(n23403), .Z(n23405) );
  XOR U23973 ( .A(n23404), .B(n23405), .Z(n23411) );
  NANDN U23974 ( .A(n23355), .B(n42093), .Z(n23357) );
  XOR U23975 ( .A(n42134), .B(a[566]), .Z(n23396) );
  NANDN U23976 ( .A(n23396), .B(n42095), .Z(n23356) );
  NAND U23977 ( .A(n23357), .B(n23356), .Z(n23409) );
  NANDN U23978 ( .A(n23358), .B(n42231), .Z(n23360) );
  XOR U23979 ( .A(n208), .B(a[562]), .Z(n23399) );
  NANDN U23980 ( .A(n23399), .B(n42234), .Z(n23359) );
  AND U23981 ( .A(n23360), .B(n23359), .Z(n23408) );
  XNOR U23982 ( .A(n23409), .B(n23408), .Z(n23410) );
  XNOR U23983 ( .A(n23411), .B(n23410), .Z(n23415) );
  NANDN U23984 ( .A(n23362), .B(n23361), .Z(n23366) );
  NAND U23985 ( .A(n23364), .B(n23363), .Z(n23365) );
  AND U23986 ( .A(n23366), .B(n23365), .Z(n23414) );
  XOR U23987 ( .A(n23415), .B(n23414), .Z(n23416) );
  NANDN U23988 ( .A(n23368), .B(n23367), .Z(n23372) );
  NANDN U23989 ( .A(n23370), .B(n23369), .Z(n23371) );
  NAND U23990 ( .A(n23372), .B(n23371), .Z(n23417) );
  XOR U23991 ( .A(n23416), .B(n23417), .Z(n23384) );
  OR U23992 ( .A(n23374), .B(n23373), .Z(n23378) );
  NANDN U23993 ( .A(n23376), .B(n23375), .Z(n23377) );
  NAND U23994 ( .A(n23378), .B(n23377), .Z(n23385) );
  XNOR U23995 ( .A(n23384), .B(n23385), .Z(n23386) );
  XNOR U23996 ( .A(n23387), .B(n23386), .Z(n23420) );
  XNOR U23997 ( .A(n23420), .B(sreg[1584]), .Z(n23422) );
  NAND U23998 ( .A(n23379), .B(sreg[1583]), .Z(n23383) );
  OR U23999 ( .A(n23381), .B(n23380), .Z(n23382) );
  AND U24000 ( .A(n23383), .B(n23382), .Z(n23421) );
  XOR U24001 ( .A(n23422), .B(n23421), .Z(c[1584]) );
  NANDN U24002 ( .A(n23385), .B(n23384), .Z(n23389) );
  NAND U24003 ( .A(n23387), .B(n23386), .Z(n23388) );
  NAND U24004 ( .A(n23389), .B(n23388), .Z(n23428) );
  NAND U24005 ( .A(b[0]), .B(a[569]), .Z(n23390) );
  XNOR U24006 ( .A(b[1]), .B(n23390), .Z(n23392) );
  NAND U24007 ( .A(n96), .B(a[568]), .Z(n23391) );
  AND U24008 ( .A(n23392), .B(n23391), .Z(n23445) );
  XOR U24009 ( .A(a[565]), .B(n42197), .Z(n23434) );
  NANDN U24010 ( .A(n23434), .B(n42173), .Z(n23395) );
  NANDN U24011 ( .A(n23393), .B(n42172), .Z(n23394) );
  NAND U24012 ( .A(n23395), .B(n23394), .Z(n23443) );
  NAND U24013 ( .A(b[7]), .B(a[561]), .Z(n23444) );
  XNOR U24014 ( .A(n23443), .B(n23444), .Z(n23446) );
  XOR U24015 ( .A(n23445), .B(n23446), .Z(n23452) );
  NANDN U24016 ( .A(n23396), .B(n42093), .Z(n23398) );
  XOR U24017 ( .A(n42134), .B(a[567]), .Z(n23437) );
  NANDN U24018 ( .A(n23437), .B(n42095), .Z(n23397) );
  NAND U24019 ( .A(n23398), .B(n23397), .Z(n23450) );
  NANDN U24020 ( .A(n23399), .B(n42231), .Z(n23401) );
  XOR U24021 ( .A(n209), .B(a[563]), .Z(n23440) );
  NANDN U24022 ( .A(n23440), .B(n42234), .Z(n23400) );
  AND U24023 ( .A(n23401), .B(n23400), .Z(n23449) );
  XNOR U24024 ( .A(n23450), .B(n23449), .Z(n23451) );
  XNOR U24025 ( .A(n23452), .B(n23451), .Z(n23456) );
  NANDN U24026 ( .A(n23403), .B(n23402), .Z(n23407) );
  NAND U24027 ( .A(n23405), .B(n23404), .Z(n23406) );
  AND U24028 ( .A(n23407), .B(n23406), .Z(n23455) );
  XOR U24029 ( .A(n23456), .B(n23455), .Z(n23457) );
  NANDN U24030 ( .A(n23409), .B(n23408), .Z(n23413) );
  NANDN U24031 ( .A(n23411), .B(n23410), .Z(n23412) );
  NAND U24032 ( .A(n23413), .B(n23412), .Z(n23458) );
  XOR U24033 ( .A(n23457), .B(n23458), .Z(n23425) );
  OR U24034 ( .A(n23415), .B(n23414), .Z(n23419) );
  NANDN U24035 ( .A(n23417), .B(n23416), .Z(n23418) );
  NAND U24036 ( .A(n23419), .B(n23418), .Z(n23426) );
  XNOR U24037 ( .A(n23425), .B(n23426), .Z(n23427) );
  XNOR U24038 ( .A(n23428), .B(n23427), .Z(n23461) );
  XNOR U24039 ( .A(n23461), .B(sreg[1585]), .Z(n23463) );
  NAND U24040 ( .A(n23420), .B(sreg[1584]), .Z(n23424) );
  OR U24041 ( .A(n23422), .B(n23421), .Z(n23423) );
  AND U24042 ( .A(n23424), .B(n23423), .Z(n23462) );
  XOR U24043 ( .A(n23463), .B(n23462), .Z(c[1585]) );
  NANDN U24044 ( .A(n23426), .B(n23425), .Z(n23430) );
  NAND U24045 ( .A(n23428), .B(n23427), .Z(n23429) );
  NAND U24046 ( .A(n23430), .B(n23429), .Z(n23469) );
  NAND U24047 ( .A(b[0]), .B(a[570]), .Z(n23431) );
  XNOR U24048 ( .A(b[1]), .B(n23431), .Z(n23433) );
  NAND U24049 ( .A(n96), .B(a[569]), .Z(n23432) );
  AND U24050 ( .A(n23433), .B(n23432), .Z(n23486) );
  XOR U24051 ( .A(a[566]), .B(n42197), .Z(n23475) );
  NANDN U24052 ( .A(n23475), .B(n42173), .Z(n23436) );
  NANDN U24053 ( .A(n23434), .B(n42172), .Z(n23435) );
  NAND U24054 ( .A(n23436), .B(n23435), .Z(n23484) );
  NAND U24055 ( .A(b[7]), .B(a[562]), .Z(n23485) );
  XNOR U24056 ( .A(n23484), .B(n23485), .Z(n23487) );
  XOR U24057 ( .A(n23486), .B(n23487), .Z(n23493) );
  NANDN U24058 ( .A(n23437), .B(n42093), .Z(n23439) );
  XOR U24059 ( .A(n42134), .B(a[568]), .Z(n23478) );
  NANDN U24060 ( .A(n23478), .B(n42095), .Z(n23438) );
  NAND U24061 ( .A(n23439), .B(n23438), .Z(n23491) );
  NANDN U24062 ( .A(n23440), .B(n42231), .Z(n23442) );
  XOR U24063 ( .A(n209), .B(a[564]), .Z(n23481) );
  NANDN U24064 ( .A(n23481), .B(n42234), .Z(n23441) );
  AND U24065 ( .A(n23442), .B(n23441), .Z(n23490) );
  XNOR U24066 ( .A(n23491), .B(n23490), .Z(n23492) );
  XNOR U24067 ( .A(n23493), .B(n23492), .Z(n23497) );
  NANDN U24068 ( .A(n23444), .B(n23443), .Z(n23448) );
  NAND U24069 ( .A(n23446), .B(n23445), .Z(n23447) );
  AND U24070 ( .A(n23448), .B(n23447), .Z(n23496) );
  XOR U24071 ( .A(n23497), .B(n23496), .Z(n23498) );
  NANDN U24072 ( .A(n23450), .B(n23449), .Z(n23454) );
  NANDN U24073 ( .A(n23452), .B(n23451), .Z(n23453) );
  NAND U24074 ( .A(n23454), .B(n23453), .Z(n23499) );
  XOR U24075 ( .A(n23498), .B(n23499), .Z(n23466) );
  OR U24076 ( .A(n23456), .B(n23455), .Z(n23460) );
  NANDN U24077 ( .A(n23458), .B(n23457), .Z(n23459) );
  NAND U24078 ( .A(n23460), .B(n23459), .Z(n23467) );
  XNOR U24079 ( .A(n23466), .B(n23467), .Z(n23468) );
  XNOR U24080 ( .A(n23469), .B(n23468), .Z(n23502) );
  XNOR U24081 ( .A(n23502), .B(sreg[1586]), .Z(n23504) );
  NAND U24082 ( .A(n23461), .B(sreg[1585]), .Z(n23465) );
  OR U24083 ( .A(n23463), .B(n23462), .Z(n23464) );
  AND U24084 ( .A(n23465), .B(n23464), .Z(n23503) );
  XOR U24085 ( .A(n23504), .B(n23503), .Z(c[1586]) );
  NANDN U24086 ( .A(n23467), .B(n23466), .Z(n23471) );
  NAND U24087 ( .A(n23469), .B(n23468), .Z(n23470) );
  NAND U24088 ( .A(n23471), .B(n23470), .Z(n23510) );
  NAND U24089 ( .A(b[0]), .B(a[571]), .Z(n23472) );
  XNOR U24090 ( .A(b[1]), .B(n23472), .Z(n23474) );
  NAND U24091 ( .A(n96), .B(a[570]), .Z(n23473) );
  AND U24092 ( .A(n23474), .B(n23473), .Z(n23527) );
  XOR U24093 ( .A(a[567]), .B(n42197), .Z(n23516) );
  NANDN U24094 ( .A(n23516), .B(n42173), .Z(n23477) );
  NANDN U24095 ( .A(n23475), .B(n42172), .Z(n23476) );
  NAND U24096 ( .A(n23477), .B(n23476), .Z(n23525) );
  NAND U24097 ( .A(b[7]), .B(a[563]), .Z(n23526) );
  XNOR U24098 ( .A(n23525), .B(n23526), .Z(n23528) );
  XOR U24099 ( .A(n23527), .B(n23528), .Z(n23534) );
  NANDN U24100 ( .A(n23478), .B(n42093), .Z(n23480) );
  XOR U24101 ( .A(n42134), .B(a[569]), .Z(n23519) );
  NANDN U24102 ( .A(n23519), .B(n42095), .Z(n23479) );
  NAND U24103 ( .A(n23480), .B(n23479), .Z(n23532) );
  NANDN U24104 ( .A(n23481), .B(n42231), .Z(n23483) );
  XOR U24105 ( .A(n209), .B(a[565]), .Z(n23522) );
  NANDN U24106 ( .A(n23522), .B(n42234), .Z(n23482) );
  AND U24107 ( .A(n23483), .B(n23482), .Z(n23531) );
  XNOR U24108 ( .A(n23532), .B(n23531), .Z(n23533) );
  XNOR U24109 ( .A(n23534), .B(n23533), .Z(n23538) );
  NANDN U24110 ( .A(n23485), .B(n23484), .Z(n23489) );
  NAND U24111 ( .A(n23487), .B(n23486), .Z(n23488) );
  AND U24112 ( .A(n23489), .B(n23488), .Z(n23537) );
  XOR U24113 ( .A(n23538), .B(n23537), .Z(n23539) );
  NANDN U24114 ( .A(n23491), .B(n23490), .Z(n23495) );
  NANDN U24115 ( .A(n23493), .B(n23492), .Z(n23494) );
  NAND U24116 ( .A(n23495), .B(n23494), .Z(n23540) );
  XOR U24117 ( .A(n23539), .B(n23540), .Z(n23507) );
  OR U24118 ( .A(n23497), .B(n23496), .Z(n23501) );
  NANDN U24119 ( .A(n23499), .B(n23498), .Z(n23500) );
  NAND U24120 ( .A(n23501), .B(n23500), .Z(n23508) );
  XNOR U24121 ( .A(n23507), .B(n23508), .Z(n23509) );
  XNOR U24122 ( .A(n23510), .B(n23509), .Z(n23543) );
  XNOR U24123 ( .A(n23543), .B(sreg[1587]), .Z(n23545) );
  NAND U24124 ( .A(n23502), .B(sreg[1586]), .Z(n23506) );
  OR U24125 ( .A(n23504), .B(n23503), .Z(n23505) );
  AND U24126 ( .A(n23506), .B(n23505), .Z(n23544) );
  XOR U24127 ( .A(n23545), .B(n23544), .Z(c[1587]) );
  NANDN U24128 ( .A(n23508), .B(n23507), .Z(n23512) );
  NAND U24129 ( .A(n23510), .B(n23509), .Z(n23511) );
  NAND U24130 ( .A(n23512), .B(n23511), .Z(n23551) );
  NAND U24131 ( .A(b[0]), .B(a[572]), .Z(n23513) );
  XNOR U24132 ( .A(b[1]), .B(n23513), .Z(n23515) );
  NAND U24133 ( .A(n96), .B(a[571]), .Z(n23514) );
  AND U24134 ( .A(n23515), .B(n23514), .Z(n23568) );
  XOR U24135 ( .A(a[568]), .B(n42197), .Z(n23557) );
  NANDN U24136 ( .A(n23557), .B(n42173), .Z(n23518) );
  NANDN U24137 ( .A(n23516), .B(n42172), .Z(n23517) );
  NAND U24138 ( .A(n23518), .B(n23517), .Z(n23566) );
  NAND U24139 ( .A(b[7]), .B(a[564]), .Z(n23567) );
  XNOR U24140 ( .A(n23566), .B(n23567), .Z(n23569) );
  XOR U24141 ( .A(n23568), .B(n23569), .Z(n23575) );
  NANDN U24142 ( .A(n23519), .B(n42093), .Z(n23521) );
  XOR U24143 ( .A(n42134), .B(a[570]), .Z(n23560) );
  NANDN U24144 ( .A(n23560), .B(n42095), .Z(n23520) );
  NAND U24145 ( .A(n23521), .B(n23520), .Z(n23573) );
  NANDN U24146 ( .A(n23522), .B(n42231), .Z(n23524) );
  XOR U24147 ( .A(n209), .B(a[566]), .Z(n23563) );
  NANDN U24148 ( .A(n23563), .B(n42234), .Z(n23523) );
  AND U24149 ( .A(n23524), .B(n23523), .Z(n23572) );
  XNOR U24150 ( .A(n23573), .B(n23572), .Z(n23574) );
  XNOR U24151 ( .A(n23575), .B(n23574), .Z(n23579) );
  NANDN U24152 ( .A(n23526), .B(n23525), .Z(n23530) );
  NAND U24153 ( .A(n23528), .B(n23527), .Z(n23529) );
  AND U24154 ( .A(n23530), .B(n23529), .Z(n23578) );
  XOR U24155 ( .A(n23579), .B(n23578), .Z(n23580) );
  NANDN U24156 ( .A(n23532), .B(n23531), .Z(n23536) );
  NANDN U24157 ( .A(n23534), .B(n23533), .Z(n23535) );
  NAND U24158 ( .A(n23536), .B(n23535), .Z(n23581) );
  XOR U24159 ( .A(n23580), .B(n23581), .Z(n23548) );
  OR U24160 ( .A(n23538), .B(n23537), .Z(n23542) );
  NANDN U24161 ( .A(n23540), .B(n23539), .Z(n23541) );
  NAND U24162 ( .A(n23542), .B(n23541), .Z(n23549) );
  XNOR U24163 ( .A(n23548), .B(n23549), .Z(n23550) );
  XNOR U24164 ( .A(n23551), .B(n23550), .Z(n23584) );
  XNOR U24165 ( .A(n23584), .B(sreg[1588]), .Z(n23586) );
  NAND U24166 ( .A(n23543), .B(sreg[1587]), .Z(n23547) );
  OR U24167 ( .A(n23545), .B(n23544), .Z(n23546) );
  AND U24168 ( .A(n23547), .B(n23546), .Z(n23585) );
  XOR U24169 ( .A(n23586), .B(n23585), .Z(c[1588]) );
  NANDN U24170 ( .A(n23549), .B(n23548), .Z(n23553) );
  NAND U24171 ( .A(n23551), .B(n23550), .Z(n23552) );
  NAND U24172 ( .A(n23553), .B(n23552), .Z(n23592) );
  NAND U24173 ( .A(b[0]), .B(a[573]), .Z(n23554) );
  XNOR U24174 ( .A(b[1]), .B(n23554), .Z(n23556) );
  NAND U24175 ( .A(n96), .B(a[572]), .Z(n23555) );
  AND U24176 ( .A(n23556), .B(n23555), .Z(n23609) );
  XOR U24177 ( .A(a[569]), .B(n42197), .Z(n23598) );
  NANDN U24178 ( .A(n23598), .B(n42173), .Z(n23559) );
  NANDN U24179 ( .A(n23557), .B(n42172), .Z(n23558) );
  NAND U24180 ( .A(n23559), .B(n23558), .Z(n23607) );
  NAND U24181 ( .A(b[7]), .B(a[565]), .Z(n23608) );
  XNOR U24182 ( .A(n23607), .B(n23608), .Z(n23610) );
  XOR U24183 ( .A(n23609), .B(n23610), .Z(n23616) );
  NANDN U24184 ( .A(n23560), .B(n42093), .Z(n23562) );
  XOR U24185 ( .A(n42134), .B(a[571]), .Z(n23601) );
  NANDN U24186 ( .A(n23601), .B(n42095), .Z(n23561) );
  NAND U24187 ( .A(n23562), .B(n23561), .Z(n23614) );
  NANDN U24188 ( .A(n23563), .B(n42231), .Z(n23565) );
  XOR U24189 ( .A(n209), .B(a[567]), .Z(n23604) );
  NANDN U24190 ( .A(n23604), .B(n42234), .Z(n23564) );
  AND U24191 ( .A(n23565), .B(n23564), .Z(n23613) );
  XNOR U24192 ( .A(n23614), .B(n23613), .Z(n23615) );
  XNOR U24193 ( .A(n23616), .B(n23615), .Z(n23620) );
  NANDN U24194 ( .A(n23567), .B(n23566), .Z(n23571) );
  NAND U24195 ( .A(n23569), .B(n23568), .Z(n23570) );
  AND U24196 ( .A(n23571), .B(n23570), .Z(n23619) );
  XOR U24197 ( .A(n23620), .B(n23619), .Z(n23621) );
  NANDN U24198 ( .A(n23573), .B(n23572), .Z(n23577) );
  NANDN U24199 ( .A(n23575), .B(n23574), .Z(n23576) );
  NAND U24200 ( .A(n23577), .B(n23576), .Z(n23622) );
  XOR U24201 ( .A(n23621), .B(n23622), .Z(n23589) );
  OR U24202 ( .A(n23579), .B(n23578), .Z(n23583) );
  NANDN U24203 ( .A(n23581), .B(n23580), .Z(n23582) );
  NAND U24204 ( .A(n23583), .B(n23582), .Z(n23590) );
  XNOR U24205 ( .A(n23589), .B(n23590), .Z(n23591) );
  XNOR U24206 ( .A(n23592), .B(n23591), .Z(n23625) );
  XNOR U24207 ( .A(n23625), .B(sreg[1589]), .Z(n23627) );
  NAND U24208 ( .A(n23584), .B(sreg[1588]), .Z(n23588) );
  OR U24209 ( .A(n23586), .B(n23585), .Z(n23587) );
  AND U24210 ( .A(n23588), .B(n23587), .Z(n23626) );
  XOR U24211 ( .A(n23627), .B(n23626), .Z(c[1589]) );
  NANDN U24212 ( .A(n23590), .B(n23589), .Z(n23594) );
  NAND U24213 ( .A(n23592), .B(n23591), .Z(n23593) );
  NAND U24214 ( .A(n23594), .B(n23593), .Z(n23633) );
  NAND U24215 ( .A(b[0]), .B(a[574]), .Z(n23595) );
  XNOR U24216 ( .A(b[1]), .B(n23595), .Z(n23597) );
  NAND U24217 ( .A(n97), .B(a[573]), .Z(n23596) );
  AND U24218 ( .A(n23597), .B(n23596), .Z(n23650) );
  XOR U24219 ( .A(a[570]), .B(n42197), .Z(n23639) );
  NANDN U24220 ( .A(n23639), .B(n42173), .Z(n23600) );
  NANDN U24221 ( .A(n23598), .B(n42172), .Z(n23599) );
  NAND U24222 ( .A(n23600), .B(n23599), .Z(n23648) );
  NAND U24223 ( .A(b[7]), .B(a[566]), .Z(n23649) );
  XNOR U24224 ( .A(n23648), .B(n23649), .Z(n23651) );
  XOR U24225 ( .A(n23650), .B(n23651), .Z(n23657) );
  NANDN U24226 ( .A(n23601), .B(n42093), .Z(n23603) );
  XOR U24227 ( .A(n42134), .B(a[572]), .Z(n23642) );
  NANDN U24228 ( .A(n23642), .B(n42095), .Z(n23602) );
  NAND U24229 ( .A(n23603), .B(n23602), .Z(n23655) );
  NANDN U24230 ( .A(n23604), .B(n42231), .Z(n23606) );
  XOR U24231 ( .A(n209), .B(a[568]), .Z(n23645) );
  NANDN U24232 ( .A(n23645), .B(n42234), .Z(n23605) );
  AND U24233 ( .A(n23606), .B(n23605), .Z(n23654) );
  XNOR U24234 ( .A(n23655), .B(n23654), .Z(n23656) );
  XNOR U24235 ( .A(n23657), .B(n23656), .Z(n23661) );
  NANDN U24236 ( .A(n23608), .B(n23607), .Z(n23612) );
  NAND U24237 ( .A(n23610), .B(n23609), .Z(n23611) );
  AND U24238 ( .A(n23612), .B(n23611), .Z(n23660) );
  XOR U24239 ( .A(n23661), .B(n23660), .Z(n23662) );
  NANDN U24240 ( .A(n23614), .B(n23613), .Z(n23618) );
  NANDN U24241 ( .A(n23616), .B(n23615), .Z(n23617) );
  NAND U24242 ( .A(n23618), .B(n23617), .Z(n23663) );
  XOR U24243 ( .A(n23662), .B(n23663), .Z(n23630) );
  OR U24244 ( .A(n23620), .B(n23619), .Z(n23624) );
  NANDN U24245 ( .A(n23622), .B(n23621), .Z(n23623) );
  NAND U24246 ( .A(n23624), .B(n23623), .Z(n23631) );
  XNOR U24247 ( .A(n23630), .B(n23631), .Z(n23632) );
  XNOR U24248 ( .A(n23633), .B(n23632), .Z(n23666) );
  XNOR U24249 ( .A(n23666), .B(sreg[1590]), .Z(n23668) );
  NAND U24250 ( .A(n23625), .B(sreg[1589]), .Z(n23629) );
  OR U24251 ( .A(n23627), .B(n23626), .Z(n23628) );
  AND U24252 ( .A(n23629), .B(n23628), .Z(n23667) );
  XOR U24253 ( .A(n23668), .B(n23667), .Z(c[1590]) );
  NANDN U24254 ( .A(n23631), .B(n23630), .Z(n23635) );
  NAND U24255 ( .A(n23633), .B(n23632), .Z(n23634) );
  NAND U24256 ( .A(n23635), .B(n23634), .Z(n23674) );
  NAND U24257 ( .A(b[0]), .B(a[575]), .Z(n23636) );
  XNOR U24258 ( .A(b[1]), .B(n23636), .Z(n23638) );
  NAND U24259 ( .A(n97), .B(a[574]), .Z(n23637) );
  AND U24260 ( .A(n23638), .B(n23637), .Z(n23691) );
  XOR U24261 ( .A(a[571]), .B(n42197), .Z(n23680) );
  NANDN U24262 ( .A(n23680), .B(n42173), .Z(n23641) );
  NANDN U24263 ( .A(n23639), .B(n42172), .Z(n23640) );
  NAND U24264 ( .A(n23641), .B(n23640), .Z(n23689) );
  NAND U24265 ( .A(b[7]), .B(a[567]), .Z(n23690) );
  XNOR U24266 ( .A(n23689), .B(n23690), .Z(n23692) );
  XOR U24267 ( .A(n23691), .B(n23692), .Z(n23698) );
  NANDN U24268 ( .A(n23642), .B(n42093), .Z(n23644) );
  XOR U24269 ( .A(n42134), .B(a[573]), .Z(n23683) );
  NANDN U24270 ( .A(n23683), .B(n42095), .Z(n23643) );
  NAND U24271 ( .A(n23644), .B(n23643), .Z(n23696) );
  NANDN U24272 ( .A(n23645), .B(n42231), .Z(n23647) );
  XOR U24273 ( .A(n209), .B(a[569]), .Z(n23686) );
  NANDN U24274 ( .A(n23686), .B(n42234), .Z(n23646) );
  AND U24275 ( .A(n23647), .B(n23646), .Z(n23695) );
  XNOR U24276 ( .A(n23696), .B(n23695), .Z(n23697) );
  XNOR U24277 ( .A(n23698), .B(n23697), .Z(n23702) );
  NANDN U24278 ( .A(n23649), .B(n23648), .Z(n23653) );
  NAND U24279 ( .A(n23651), .B(n23650), .Z(n23652) );
  AND U24280 ( .A(n23653), .B(n23652), .Z(n23701) );
  XOR U24281 ( .A(n23702), .B(n23701), .Z(n23703) );
  NANDN U24282 ( .A(n23655), .B(n23654), .Z(n23659) );
  NANDN U24283 ( .A(n23657), .B(n23656), .Z(n23658) );
  NAND U24284 ( .A(n23659), .B(n23658), .Z(n23704) );
  XOR U24285 ( .A(n23703), .B(n23704), .Z(n23671) );
  OR U24286 ( .A(n23661), .B(n23660), .Z(n23665) );
  NANDN U24287 ( .A(n23663), .B(n23662), .Z(n23664) );
  NAND U24288 ( .A(n23665), .B(n23664), .Z(n23672) );
  XNOR U24289 ( .A(n23671), .B(n23672), .Z(n23673) );
  XNOR U24290 ( .A(n23674), .B(n23673), .Z(n23707) );
  XNOR U24291 ( .A(n23707), .B(sreg[1591]), .Z(n23709) );
  NAND U24292 ( .A(n23666), .B(sreg[1590]), .Z(n23670) );
  OR U24293 ( .A(n23668), .B(n23667), .Z(n23669) );
  AND U24294 ( .A(n23670), .B(n23669), .Z(n23708) );
  XOR U24295 ( .A(n23709), .B(n23708), .Z(c[1591]) );
  NANDN U24296 ( .A(n23672), .B(n23671), .Z(n23676) );
  NAND U24297 ( .A(n23674), .B(n23673), .Z(n23675) );
  NAND U24298 ( .A(n23676), .B(n23675), .Z(n23715) );
  NAND U24299 ( .A(b[0]), .B(a[576]), .Z(n23677) );
  XNOR U24300 ( .A(b[1]), .B(n23677), .Z(n23679) );
  NAND U24301 ( .A(n97), .B(a[575]), .Z(n23678) );
  AND U24302 ( .A(n23679), .B(n23678), .Z(n23732) );
  XOR U24303 ( .A(a[572]), .B(n42197), .Z(n23721) );
  NANDN U24304 ( .A(n23721), .B(n42173), .Z(n23682) );
  NANDN U24305 ( .A(n23680), .B(n42172), .Z(n23681) );
  NAND U24306 ( .A(n23682), .B(n23681), .Z(n23730) );
  NAND U24307 ( .A(b[7]), .B(a[568]), .Z(n23731) );
  XNOR U24308 ( .A(n23730), .B(n23731), .Z(n23733) );
  XOR U24309 ( .A(n23732), .B(n23733), .Z(n23739) );
  NANDN U24310 ( .A(n23683), .B(n42093), .Z(n23685) );
  XOR U24311 ( .A(n42134), .B(a[574]), .Z(n23724) );
  NANDN U24312 ( .A(n23724), .B(n42095), .Z(n23684) );
  NAND U24313 ( .A(n23685), .B(n23684), .Z(n23737) );
  NANDN U24314 ( .A(n23686), .B(n42231), .Z(n23688) );
  XOR U24315 ( .A(n209), .B(a[570]), .Z(n23727) );
  NANDN U24316 ( .A(n23727), .B(n42234), .Z(n23687) );
  AND U24317 ( .A(n23688), .B(n23687), .Z(n23736) );
  XNOR U24318 ( .A(n23737), .B(n23736), .Z(n23738) );
  XNOR U24319 ( .A(n23739), .B(n23738), .Z(n23743) );
  NANDN U24320 ( .A(n23690), .B(n23689), .Z(n23694) );
  NAND U24321 ( .A(n23692), .B(n23691), .Z(n23693) );
  AND U24322 ( .A(n23694), .B(n23693), .Z(n23742) );
  XOR U24323 ( .A(n23743), .B(n23742), .Z(n23744) );
  NANDN U24324 ( .A(n23696), .B(n23695), .Z(n23700) );
  NANDN U24325 ( .A(n23698), .B(n23697), .Z(n23699) );
  NAND U24326 ( .A(n23700), .B(n23699), .Z(n23745) );
  XOR U24327 ( .A(n23744), .B(n23745), .Z(n23712) );
  OR U24328 ( .A(n23702), .B(n23701), .Z(n23706) );
  NANDN U24329 ( .A(n23704), .B(n23703), .Z(n23705) );
  NAND U24330 ( .A(n23706), .B(n23705), .Z(n23713) );
  XNOR U24331 ( .A(n23712), .B(n23713), .Z(n23714) );
  XNOR U24332 ( .A(n23715), .B(n23714), .Z(n23748) );
  XNOR U24333 ( .A(n23748), .B(sreg[1592]), .Z(n23750) );
  NAND U24334 ( .A(n23707), .B(sreg[1591]), .Z(n23711) );
  OR U24335 ( .A(n23709), .B(n23708), .Z(n23710) );
  AND U24336 ( .A(n23711), .B(n23710), .Z(n23749) );
  XOR U24337 ( .A(n23750), .B(n23749), .Z(c[1592]) );
  NANDN U24338 ( .A(n23713), .B(n23712), .Z(n23717) );
  NAND U24339 ( .A(n23715), .B(n23714), .Z(n23716) );
  NAND U24340 ( .A(n23717), .B(n23716), .Z(n23756) );
  NAND U24341 ( .A(b[0]), .B(a[577]), .Z(n23718) );
  XNOR U24342 ( .A(b[1]), .B(n23718), .Z(n23720) );
  NAND U24343 ( .A(n97), .B(a[576]), .Z(n23719) );
  AND U24344 ( .A(n23720), .B(n23719), .Z(n23773) );
  XOR U24345 ( .A(a[573]), .B(n42197), .Z(n23762) );
  NANDN U24346 ( .A(n23762), .B(n42173), .Z(n23723) );
  NANDN U24347 ( .A(n23721), .B(n42172), .Z(n23722) );
  NAND U24348 ( .A(n23723), .B(n23722), .Z(n23771) );
  NAND U24349 ( .A(b[7]), .B(a[569]), .Z(n23772) );
  XNOR U24350 ( .A(n23771), .B(n23772), .Z(n23774) );
  XOR U24351 ( .A(n23773), .B(n23774), .Z(n23780) );
  NANDN U24352 ( .A(n23724), .B(n42093), .Z(n23726) );
  XOR U24353 ( .A(n42134), .B(a[575]), .Z(n23765) );
  NANDN U24354 ( .A(n23765), .B(n42095), .Z(n23725) );
  NAND U24355 ( .A(n23726), .B(n23725), .Z(n23778) );
  NANDN U24356 ( .A(n23727), .B(n42231), .Z(n23729) );
  XOR U24357 ( .A(n209), .B(a[571]), .Z(n23768) );
  NANDN U24358 ( .A(n23768), .B(n42234), .Z(n23728) );
  AND U24359 ( .A(n23729), .B(n23728), .Z(n23777) );
  XNOR U24360 ( .A(n23778), .B(n23777), .Z(n23779) );
  XNOR U24361 ( .A(n23780), .B(n23779), .Z(n23784) );
  NANDN U24362 ( .A(n23731), .B(n23730), .Z(n23735) );
  NAND U24363 ( .A(n23733), .B(n23732), .Z(n23734) );
  AND U24364 ( .A(n23735), .B(n23734), .Z(n23783) );
  XOR U24365 ( .A(n23784), .B(n23783), .Z(n23785) );
  NANDN U24366 ( .A(n23737), .B(n23736), .Z(n23741) );
  NANDN U24367 ( .A(n23739), .B(n23738), .Z(n23740) );
  NAND U24368 ( .A(n23741), .B(n23740), .Z(n23786) );
  XOR U24369 ( .A(n23785), .B(n23786), .Z(n23753) );
  OR U24370 ( .A(n23743), .B(n23742), .Z(n23747) );
  NANDN U24371 ( .A(n23745), .B(n23744), .Z(n23746) );
  NAND U24372 ( .A(n23747), .B(n23746), .Z(n23754) );
  XNOR U24373 ( .A(n23753), .B(n23754), .Z(n23755) );
  XNOR U24374 ( .A(n23756), .B(n23755), .Z(n23789) );
  XNOR U24375 ( .A(n23789), .B(sreg[1593]), .Z(n23791) );
  NAND U24376 ( .A(n23748), .B(sreg[1592]), .Z(n23752) );
  OR U24377 ( .A(n23750), .B(n23749), .Z(n23751) );
  AND U24378 ( .A(n23752), .B(n23751), .Z(n23790) );
  XOR U24379 ( .A(n23791), .B(n23790), .Z(c[1593]) );
  NANDN U24380 ( .A(n23754), .B(n23753), .Z(n23758) );
  NAND U24381 ( .A(n23756), .B(n23755), .Z(n23757) );
  NAND U24382 ( .A(n23758), .B(n23757), .Z(n23797) );
  NAND U24383 ( .A(b[0]), .B(a[578]), .Z(n23759) );
  XNOR U24384 ( .A(b[1]), .B(n23759), .Z(n23761) );
  NAND U24385 ( .A(n97), .B(a[577]), .Z(n23760) );
  AND U24386 ( .A(n23761), .B(n23760), .Z(n23814) );
  XOR U24387 ( .A(a[574]), .B(n42197), .Z(n23803) );
  NANDN U24388 ( .A(n23803), .B(n42173), .Z(n23764) );
  NANDN U24389 ( .A(n23762), .B(n42172), .Z(n23763) );
  NAND U24390 ( .A(n23764), .B(n23763), .Z(n23812) );
  NAND U24391 ( .A(b[7]), .B(a[570]), .Z(n23813) );
  XNOR U24392 ( .A(n23812), .B(n23813), .Z(n23815) );
  XOR U24393 ( .A(n23814), .B(n23815), .Z(n23821) );
  NANDN U24394 ( .A(n23765), .B(n42093), .Z(n23767) );
  XOR U24395 ( .A(n42134), .B(a[576]), .Z(n23806) );
  NANDN U24396 ( .A(n23806), .B(n42095), .Z(n23766) );
  NAND U24397 ( .A(n23767), .B(n23766), .Z(n23819) );
  NANDN U24398 ( .A(n23768), .B(n42231), .Z(n23770) );
  XOR U24399 ( .A(n209), .B(a[572]), .Z(n23809) );
  NANDN U24400 ( .A(n23809), .B(n42234), .Z(n23769) );
  AND U24401 ( .A(n23770), .B(n23769), .Z(n23818) );
  XNOR U24402 ( .A(n23819), .B(n23818), .Z(n23820) );
  XNOR U24403 ( .A(n23821), .B(n23820), .Z(n23825) );
  NANDN U24404 ( .A(n23772), .B(n23771), .Z(n23776) );
  NAND U24405 ( .A(n23774), .B(n23773), .Z(n23775) );
  AND U24406 ( .A(n23776), .B(n23775), .Z(n23824) );
  XOR U24407 ( .A(n23825), .B(n23824), .Z(n23826) );
  NANDN U24408 ( .A(n23778), .B(n23777), .Z(n23782) );
  NANDN U24409 ( .A(n23780), .B(n23779), .Z(n23781) );
  NAND U24410 ( .A(n23782), .B(n23781), .Z(n23827) );
  XOR U24411 ( .A(n23826), .B(n23827), .Z(n23794) );
  OR U24412 ( .A(n23784), .B(n23783), .Z(n23788) );
  NANDN U24413 ( .A(n23786), .B(n23785), .Z(n23787) );
  NAND U24414 ( .A(n23788), .B(n23787), .Z(n23795) );
  XNOR U24415 ( .A(n23794), .B(n23795), .Z(n23796) );
  XNOR U24416 ( .A(n23797), .B(n23796), .Z(n23830) );
  XNOR U24417 ( .A(n23830), .B(sreg[1594]), .Z(n23832) );
  NAND U24418 ( .A(n23789), .B(sreg[1593]), .Z(n23793) );
  OR U24419 ( .A(n23791), .B(n23790), .Z(n23792) );
  AND U24420 ( .A(n23793), .B(n23792), .Z(n23831) );
  XOR U24421 ( .A(n23832), .B(n23831), .Z(c[1594]) );
  NANDN U24422 ( .A(n23795), .B(n23794), .Z(n23799) );
  NAND U24423 ( .A(n23797), .B(n23796), .Z(n23798) );
  NAND U24424 ( .A(n23799), .B(n23798), .Z(n23838) );
  NAND U24425 ( .A(b[0]), .B(a[579]), .Z(n23800) );
  XNOR U24426 ( .A(b[1]), .B(n23800), .Z(n23802) );
  NAND U24427 ( .A(n97), .B(a[578]), .Z(n23801) );
  AND U24428 ( .A(n23802), .B(n23801), .Z(n23855) );
  XOR U24429 ( .A(a[575]), .B(n42197), .Z(n23844) );
  NANDN U24430 ( .A(n23844), .B(n42173), .Z(n23805) );
  NANDN U24431 ( .A(n23803), .B(n42172), .Z(n23804) );
  NAND U24432 ( .A(n23805), .B(n23804), .Z(n23853) );
  NAND U24433 ( .A(b[7]), .B(a[571]), .Z(n23854) );
  XNOR U24434 ( .A(n23853), .B(n23854), .Z(n23856) );
  XOR U24435 ( .A(n23855), .B(n23856), .Z(n23862) );
  NANDN U24436 ( .A(n23806), .B(n42093), .Z(n23808) );
  XOR U24437 ( .A(n42134), .B(a[577]), .Z(n23847) );
  NANDN U24438 ( .A(n23847), .B(n42095), .Z(n23807) );
  NAND U24439 ( .A(n23808), .B(n23807), .Z(n23860) );
  NANDN U24440 ( .A(n23809), .B(n42231), .Z(n23811) );
  XOR U24441 ( .A(n209), .B(a[573]), .Z(n23850) );
  NANDN U24442 ( .A(n23850), .B(n42234), .Z(n23810) );
  AND U24443 ( .A(n23811), .B(n23810), .Z(n23859) );
  XNOR U24444 ( .A(n23860), .B(n23859), .Z(n23861) );
  XNOR U24445 ( .A(n23862), .B(n23861), .Z(n23866) );
  NANDN U24446 ( .A(n23813), .B(n23812), .Z(n23817) );
  NAND U24447 ( .A(n23815), .B(n23814), .Z(n23816) );
  AND U24448 ( .A(n23817), .B(n23816), .Z(n23865) );
  XOR U24449 ( .A(n23866), .B(n23865), .Z(n23867) );
  NANDN U24450 ( .A(n23819), .B(n23818), .Z(n23823) );
  NANDN U24451 ( .A(n23821), .B(n23820), .Z(n23822) );
  NAND U24452 ( .A(n23823), .B(n23822), .Z(n23868) );
  XOR U24453 ( .A(n23867), .B(n23868), .Z(n23835) );
  OR U24454 ( .A(n23825), .B(n23824), .Z(n23829) );
  NANDN U24455 ( .A(n23827), .B(n23826), .Z(n23828) );
  NAND U24456 ( .A(n23829), .B(n23828), .Z(n23836) );
  XNOR U24457 ( .A(n23835), .B(n23836), .Z(n23837) );
  XNOR U24458 ( .A(n23838), .B(n23837), .Z(n23871) );
  XNOR U24459 ( .A(n23871), .B(sreg[1595]), .Z(n23873) );
  NAND U24460 ( .A(n23830), .B(sreg[1594]), .Z(n23834) );
  OR U24461 ( .A(n23832), .B(n23831), .Z(n23833) );
  AND U24462 ( .A(n23834), .B(n23833), .Z(n23872) );
  XOR U24463 ( .A(n23873), .B(n23872), .Z(c[1595]) );
  NANDN U24464 ( .A(n23836), .B(n23835), .Z(n23840) );
  NAND U24465 ( .A(n23838), .B(n23837), .Z(n23839) );
  NAND U24466 ( .A(n23840), .B(n23839), .Z(n23879) );
  NAND U24467 ( .A(b[0]), .B(a[580]), .Z(n23841) );
  XNOR U24468 ( .A(b[1]), .B(n23841), .Z(n23843) );
  NAND U24469 ( .A(n97), .B(a[579]), .Z(n23842) );
  AND U24470 ( .A(n23843), .B(n23842), .Z(n23896) );
  XOR U24471 ( .A(a[576]), .B(n42197), .Z(n23885) );
  NANDN U24472 ( .A(n23885), .B(n42173), .Z(n23846) );
  NANDN U24473 ( .A(n23844), .B(n42172), .Z(n23845) );
  NAND U24474 ( .A(n23846), .B(n23845), .Z(n23894) );
  NAND U24475 ( .A(b[7]), .B(a[572]), .Z(n23895) );
  XNOR U24476 ( .A(n23894), .B(n23895), .Z(n23897) );
  XOR U24477 ( .A(n23896), .B(n23897), .Z(n23903) );
  NANDN U24478 ( .A(n23847), .B(n42093), .Z(n23849) );
  XOR U24479 ( .A(n42134), .B(a[578]), .Z(n23888) );
  NANDN U24480 ( .A(n23888), .B(n42095), .Z(n23848) );
  NAND U24481 ( .A(n23849), .B(n23848), .Z(n23901) );
  NANDN U24482 ( .A(n23850), .B(n42231), .Z(n23852) );
  XOR U24483 ( .A(n209), .B(a[574]), .Z(n23891) );
  NANDN U24484 ( .A(n23891), .B(n42234), .Z(n23851) );
  AND U24485 ( .A(n23852), .B(n23851), .Z(n23900) );
  XNOR U24486 ( .A(n23901), .B(n23900), .Z(n23902) );
  XNOR U24487 ( .A(n23903), .B(n23902), .Z(n23907) );
  NANDN U24488 ( .A(n23854), .B(n23853), .Z(n23858) );
  NAND U24489 ( .A(n23856), .B(n23855), .Z(n23857) );
  AND U24490 ( .A(n23858), .B(n23857), .Z(n23906) );
  XOR U24491 ( .A(n23907), .B(n23906), .Z(n23908) );
  NANDN U24492 ( .A(n23860), .B(n23859), .Z(n23864) );
  NANDN U24493 ( .A(n23862), .B(n23861), .Z(n23863) );
  NAND U24494 ( .A(n23864), .B(n23863), .Z(n23909) );
  XOR U24495 ( .A(n23908), .B(n23909), .Z(n23876) );
  OR U24496 ( .A(n23866), .B(n23865), .Z(n23870) );
  NANDN U24497 ( .A(n23868), .B(n23867), .Z(n23869) );
  NAND U24498 ( .A(n23870), .B(n23869), .Z(n23877) );
  XNOR U24499 ( .A(n23876), .B(n23877), .Z(n23878) );
  XNOR U24500 ( .A(n23879), .B(n23878), .Z(n23912) );
  XNOR U24501 ( .A(n23912), .B(sreg[1596]), .Z(n23914) );
  NAND U24502 ( .A(n23871), .B(sreg[1595]), .Z(n23875) );
  OR U24503 ( .A(n23873), .B(n23872), .Z(n23874) );
  AND U24504 ( .A(n23875), .B(n23874), .Z(n23913) );
  XOR U24505 ( .A(n23914), .B(n23913), .Z(c[1596]) );
  NANDN U24506 ( .A(n23877), .B(n23876), .Z(n23881) );
  NAND U24507 ( .A(n23879), .B(n23878), .Z(n23880) );
  NAND U24508 ( .A(n23881), .B(n23880), .Z(n23920) );
  NAND U24509 ( .A(b[0]), .B(a[581]), .Z(n23882) );
  XNOR U24510 ( .A(b[1]), .B(n23882), .Z(n23884) );
  NAND U24511 ( .A(n98), .B(a[580]), .Z(n23883) );
  AND U24512 ( .A(n23884), .B(n23883), .Z(n23937) );
  XOR U24513 ( .A(a[577]), .B(n42197), .Z(n23926) );
  NANDN U24514 ( .A(n23926), .B(n42173), .Z(n23887) );
  NANDN U24515 ( .A(n23885), .B(n42172), .Z(n23886) );
  NAND U24516 ( .A(n23887), .B(n23886), .Z(n23935) );
  NAND U24517 ( .A(b[7]), .B(a[573]), .Z(n23936) );
  XNOR U24518 ( .A(n23935), .B(n23936), .Z(n23938) );
  XOR U24519 ( .A(n23937), .B(n23938), .Z(n23944) );
  NANDN U24520 ( .A(n23888), .B(n42093), .Z(n23890) );
  XOR U24521 ( .A(n42134), .B(a[579]), .Z(n23929) );
  NANDN U24522 ( .A(n23929), .B(n42095), .Z(n23889) );
  NAND U24523 ( .A(n23890), .B(n23889), .Z(n23942) );
  NANDN U24524 ( .A(n23891), .B(n42231), .Z(n23893) );
  XOR U24525 ( .A(n210), .B(a[575]), .Z(n23932) );
  NANDN U24526 ( .A(n23932), .B(n42234), .Z(n23892) );
  AND U24527 ( .A(n23893), .B(n23892), .Z(n23941) );
  XNOR U24528 ( .A(n23942), .B(n23941), .Z(n23943) );
  XNOR U24529 ( .A(n23944), .B(n23943), .Z(n23948) );
  NANDN U24530 ( .A(n23895), .B(n23894), .Z(n23899) );
  NAND U24531 ( .A(n23897), .B(n23896), .Z(n23898) );
  AND U24532 ( .A(n23899), .B(n23898), .Z(n23947) );
  XOR U24533 ( .A(n23948), .B(n23947), .Z(n23949) );
  NANDN U24534 ( .A(n23901), .B(n23900), .Z(n23905) );
  NANDN U24535 ( .A(n23903), .B(n23902), .Z(n23904) );
  NAND U24536 ( .A(n23905), .B(n23904), .Z(n23950) );
  XOR U24537 ( .A(n23949), .B(n23950), .Z(n23917) );
  OR U24538 ( .A(n23907), .B(n23906), .Z(n23911) );
  NANDN U24539 ( .A(n23909), .B(n23908), .Z(n23910) );
  NAND U24540 ( .A(n23911), .B(n23910), .Z(n23918) );
  XNOR U24541 ( .A(n23917), .B(n23918), .Z(n23919) );
  XNOR U24542 ( .A(n23920), .B(n23919), .Z(n23953) );
  XNOR U24543 ( .A(n23953), .B(sreg[1597]), .Z(n23955) );
  NAND U24544 ( .A(n23912), .B(sreg[1596]), .Z(n23916) );
  OR U24545 ( .A(n23914), .B(n23913), .Z(n23915) );
  AND U24546 ( .A(n23916), .B(n23915), .Z(n23954) );
  XOR U24547 ( .A(n23955), .B(n23954), .Z(c[1597]) );
  NANDN U24548 ( .A(n23918), .B(n23917), .Z(n23922) );
  NAND U24549 ( .A(n23920), .B(n23919), .Z(n23921) );
  NAND U24550 ( .A(n23922), .B(n23921), .Z(n23961) );
  NAND U24551 ( .A(b[0]), .B(a[582]), .Z(n23923) );
  XNOR U24552 ( .A(b[1]), .B(n23923), .Z(n23925) );
  NAND U24553 ( .A(n98), .B(a[581]), .Z(n23924) );
  AND U24554 ( .A(n23925), .B(n23924), .Z(n23978) );
  XOR U24555 ( .A(a[578]), .B(n42197), .Z(n23967) );
  NANDN U24556 ( .A(n23967), .B(n42173), .Z(n23928) );
  NANDN U24557 ( .A(n23926), .B(n42172), .Z(n23927) );
  NAND U24558 ( .A(n23928), .B(n23927), .Z(n23976) );
  NAND U24559 ( .A(b[7]), .B(a[574]), .Z(n23977) );
  XNOR U24560 ( .A(n23976), .B(n23977), .Z(n23979) );
  XOR U24561 ( .A(n23978), .B(n23979), .Z(n23985) );
  NANDN U24562 ( .A(n23929), .B(n42093), .Z(n23931) );
  XOR U24563 ( .A(n42134), .B(a[580]), .Z(n23970) );
  NANDN U24564 ( .A(n23970), .B(n42095), .Z(n23930) );
  NAND U24565 ( .A(n23931), .B(n23930), .Z(n23983) );
  NANDN U24566 ( .A(n23932), .B(n42231), .Z(n23934) );
  XOR U24567 ( .A(n210), .B(a[576]), .Z(n23973) );
  NANDN U24568 ( .A(n23973), .B(n42234), .Z(n23933) );
  AND U24569 ( .A(n23934), .B(n23933), .Z(n23982) );
  XNOR U24570 ( .A(n23983), .B(n23982), .Z(n23984) );
  XNOR U24571 ( .A(n23985), .B(n23984), .Z(n23989) );
  NANDN U24572 ( .A(n23936), .B(n23935), .Z(n23940) );
  NAND U24573 ( .A(n23938), .B(n23937), .Z(n23939) );
  AND U24574 ( .A(n23940), .B(n23939), .Z(n23988) );
  XOR U24575 ( .A(n23989), .B(n23988), .Z(n23990) );
  NANDN U24576 ( .A(n23942), .B(n23941), .Z(n23946) );
  NANDN U24577 ( .A(n23944), .B(n23943), .Z(n23945) );
  NAND U24578 ( .A(n23946), .B(n23945), .Z(n23991) );
  XOR U24579 ( .A(n23990), .B(n23991), .Z(n23958) );
  OR U24580 ( .A(n23948), .B(n23947), .Z(n23952) );
  NANDN U24581 ( .A(n23950), .B(n23949), .Z(n23951) );
  NAND U24582 ( .A(n23952), .B(n23951), .Z(n23959) );
  XNOR U24583 ( .A(n23958), .B(n23959), .Z(n23960) );
  XNOR U24584 ( .A(n23961), .B(n23960), .Z(n23994) );
  XNOR U24585 ( .A(n23994), .B(sreg[1598]), .Z(n23996) );
  NAND U24586 ( .A(n23953), .B(sreg[1597]), .Z(n23957) );
  OR U24587 ( .A(n23955), .B(n23954), .Z(n23956) );
  AND U24588 ( .A(n23957), .B(n23956), .Z(n23995) );
  XOR U24589 ( .A(n23996), .B(n23995), .Z(c[1598]) );
  NANDN U24590 ( .A(n23959), .B(n23958), .Z(n23963) );
  NAND U24591 ( .A(n23961), .B(n23960), .Z(n23962) );
  NAND U24592 ( .A(n23963), .B(n23962), .Z(n24002) );
  NAND U24593 ( .A(b[0]), .B(a[583]), .Z(n23964) );
  XNOR U24594 ( .A(b[1]), .B(n23964), .Z(n23966) );
  NAND U24595 ( .A(n98), .B(a[582]), .Z(n23965) );
  AND U24596 ( .A(n23966), .B(n23965), .Z(n24019) );
  XOR U24597 ( .A(a[579]), .B(n42197), .Z(n24008) );
  NANDN U24598 ( .A(n24008), .B(n42173), .Z(n23969) );
  NANDN U24599 ( .A(n23967), .B(n42172), .Z(n23968) );
  NAND U24600 ( .A(n23969), .B(n23968), .Z(n24017) );
  NAND U24601 ( .A(b[7]), .B(a[575]), .Z(n24018) );
  XNOR U24602 ( .A(n24017), .B(n24018), .Z(n24020) );
  XOR U24603 ( .A(n24019), .B(n24020), .Z(n24026) );
  NANDN U24604 ( .A(n23970), .B(n42093), .Z(n23972) );
  XOR U24605 ( .A(n42134), .B(a[581]), .Z(n24011) );
  NANDN U24606 ( .A(n24011), .B(n42095), .Z(n23971) );
  NAND U24607 ( .A(n23972), .B(n23971), .Z(n24024) );
  NANDN U24608 ( .A(n23973), .B(n42231), .Z(n23975) );
  XOR U24609 ( .A(n210), .B(a[577]), .Z(n24014) );
  NANDN U24610 ( .A(n24014), .B(n42234), .Z(n23974) );
  AND U24611 ( .A(n23975), .B(n23974), .Z(n24023) );
  XNOR U24612 ( .A(n24024), .B(n24023), .Z(n24025) );
  XNOR U24613 ( .A(n24026), .B(n24025), .Z(n24030) );
  NANDN U24614 ( .A(n23977), .B(n23976), .Z(n23981) );
  NAND U24615 ( .A(n23979), .B(n23978), .Z(n23980) );
  AND U24616 ( .A(n23981), .B(n23980), .Z(n24029) );
  XOR U24617 ( .A(n24030), .B(n24029), .Z(n24031) );
  NANDN U24618 ( .A(n23983), .B(n23982), .Z(n23987) );
  NANDN U24619 ( .A(n23985), .B(n23984), .Z(n23986) );
  NAND U24620 ( .A(n23987), .B(n23986), .Z(n24032) );
  XOR U24621 ( .A(n24031), .B(n24032), .Z(n23999) );
  OR U24622 ( .A(n23989), .B(n23988), .Z(n23993) );
  NANDN U24623 ( .A(n23991), .B(n23990), .Z(n23992) );
  NAND U24624 ( .A(n23993), .B(n23992), .Z(n24000) );
  XNOR U24625 ( .A(n23999), .B(n24000), .Z(n24001) );
  XNOR U24626 ( .A(n24002), .B(n24001), .Z(n24035) );
  XNOR U24627 ( .A(n24035), .B(sreg[1599]), .Z(n24037) );
  NAND U24628 ( .A(n23994), .B(sreg[1598]), .Z(n23998) );
  OR U24629 ( .A(n23996), .B(n23995), .Z(n23997) );
  AND U24630 ( .A(n23998), .B(n23997), .Z(n24036) );
  XOR U24631 ( .A(n24037), .B(n24036), .Z(c[1599]) );
  NANDN U24632 ( .A(n24000), .B(n23999), .Z(n24004) );
  NAND U24633 ( .A(n24002), .B(n24001), .Z(n24003) );
  NAND U24634 ( .A(n24004), .B(n24003), .Z(n24043) );
  NAND U24635 ( .A(b[0]), .B(a[584]), .Z(n24005) );
  XNOR U24636 ( .A(b[1]), .B(n24005), .Z(n24007) );
  NAND U24637 ( .A(n98), .B(a[583]), .Z(n24006) );
  AND U24638 ( .A(n24007), .B(n24006), .Z(n24060) );
  XOR U24639 ( .A(a[580]), .B(n42197), .Z(n24049) );
  NANDN U24640 ( .A(n24049), .B(n42173), .Z(n24010) );
  NANDN U24641 ( .A(n24008), .B(n42172), .Z(n24009) );
  NAND U24642 ( .A(n24010), .B(n24009), .Z(n24058) );
  NAND U24643 ( .A(b[7]), .B(a[576]), .Z(n24059) );
  XNOR U24644 ( .A(n24058), .B(n24059), .Z(n24061) );
  XOR U24645 ( .A(n24060), .B(n24061), .Z(n24067) );
  NANDN U24646 ( .A(n24011), .B(n42093), .Z(n24013) );
  XOR U24647 ( .A(n42134), .B(a[582]), .Z(n24052) );
  NANDN U24648 ( .A(n24052), .B(n42095), .Z(n24012) );
  NAND U24649 ( .A(n24013), .B(n24012), .Z(n24065) );
  NANDN U24650 ( .A(n24014), .B(n42231), .Z(n24016) );
  XOR U24651 ( .A(n210), .B(a[578]), .Z(n24055) );
  NANDN U24652 ( .A(n24055), .B(n42234), .Z(n24015) );
  AND U24653 ( .A(n24016), .B(n24015), .Z(n24064) );
  XNOR U24654 ( .A(n24065), .B(n24064), .Z(n24066) );
  XNOR U24655 ( .A(n24067), .B(n24066), .Z(n24071) );
  NANDN U24656 ( .A(n24018), .B(n24017), .Z(n24022) );
  NAND U24657 ( .A(n24020), .B(n24019), .Z(n24021) );
  AND U24658 ( .A(n24022), .B(n24021), .Z(n24070) );
  XOR U24659 ( .A(n24071), .B(n24070), .Z(n24072) );
  NANDN U24660 ( .A(n24024), .B(n24023), .Z(n24028) );
  NANDN U24661 ( .A(n24026), .B(n24025), .Z(n24027) );
  NAND U24662 ( .A(n24028), .B(n24027), .Z(n24073) );
  XOR U24663 ( .A(n24072), .B(n24073), .Z(n24040) );
  OR U24664 ( .A(n24030), .B(n24029), .Z(n24034) );
  NANDN U24665 ( .A(n24032), .B(n24031), .Z(n24033) );
  NAND U24666 ( .A(n24034), .B(n24033), .Z(n24041) );
  XNOR U24667 ( .A(n24040), .B(n24041), .Z(n24042) );
  XNOR U24668 ( .A(n24043), .B(n24042), .Z(n24076) );
  XNOR U24669 ( .A(n24076), .B(sreg[1600]), .Z(n24078) );
  NAND U24670 ( .A(n24035), .B(sreg[1599]), .Z(n24039) );
  OR U24671 ( .A(n24037), .B(n24036), .Z(n24038) );
  AND U24672 ( .A(n24039), .B(n24038), .Z(n24077) );
  XOR U24673 ( .A(n24078), .B(n24077), .Z(c[1600]) );
  NANDN U24674 ( .A(n24041), .B(n24040), .Z(n24045) );
  NAND U24675 ( .A(n24043), .B(n24042), .Z(n24044) );
  NAND U24676 ( .A(n24045), .B(n24044), .Z(n24084) );
  NAND U24677 ( .A(b[0]), .B(a[585]), .Z(n24046) );
  XNOR U24678 ( .A(b[1]), .B(n24046), .Z(n24048) );
  NAND U24679 ( .A(n98), .B(a[584]), .Z(n24047) );
  AND U24680 ( .A(n24048), .B(n24047), .Z(n24101) );
  XOR U24681 ( .A(a[581]), .B(n42197), .Z(n24090) );
  NANDN U24682 ( .A(n24090), .B(n42173), .Z(n24051) );
  NANDN U24683 ( .A(n24049), .B(n42172), .Z(n24050) );
  NAND U24684 ( .A(n24051), .B(n24050), .Z(n24099) );
  NAND U24685 ( .A(b[7]), .B(a[577]), .Z(n24100) );
  XNOR U24686 ( .A(n24099), .B(n24100), .Z(n24102) );
  XOR U24687 ( .A(n24101), .B(n24102), .Z(n24108) );
  NANDN U24688 ( .A(n24052), .B(n42093), .Z(n24054) );
  XOR U24689 ( .A(n42134), .B(a[583]), .Z(n24093) );
  NANDN U24690 ( .A(n24093), .B(n42095), .Z(n24053) );
  NAND U24691 ( .A(n24054), .B(n24053), .Z(n24106) );
  NANDN U24692 ( .A(n24055), .B(n42231), .Z(n24057) );
  XOR U24693 ( .A(n210), .B(a[579]), .Z(n24096) );
  NANDN U24694 ( .A(n24096), .B(n42234), .Z(n24056) );
  AND U24695 ( .A(n24057), .B(n24056), .Z(n24105) );
  XNOR U24696 ( .A(n24106), .B(n24105), .Z(n24107) );
  XNOR U24697 ( .A(n24108), .B(n24107), .Z(n24112) );
  NANDN U24698 ( .A(n24059), .B(n24058), .Z(n24063) );
  NAND U24699 ( .A(n24061), .B(n24060), .Z(n24062) );
  AND U24700 ( .A(n24063), .B(n24062), .Z(n24111) );
  XOR U24701 ( .A(n24112), .B(n24111), .Z(n24113) );
  NANDN U24702 ( .A(n24065), .B(n24064), .Z(n24069) );
  NANDN U24703 ( .A(n24067), .B(n24066), .Z(n24068) );
  NAND U24704 ( .A(n24069), .B(n24068), .Z(n24114) );
  XOR U24705 ( .A(n24113), .B(n24114), .Z(n24081) );
  OR U24706 ( .A(n24071), .B(n24070), .Z(n24075) );
  NANDN U24707 ( .A(n24073), .B(n24072), .Z(n24074) );
  NAND U24708 ( .A(n24075), .B(n24074), .Z(n24082) );
  XNOR U24709 ( .A(n24081), .B(n24082), .Z(n24083) );
  XNOR U24710 ( .A(n24084), .B(n24083), .Z(n24117) );
  XNOR U24711 ( .A(n24117), .B(sreg[1601]), .Z(n24119) );
  NAND U24712 ( .A(n24076), .B(sreg[1600]), .Z(n24080) );
  OR U24713 ( .A(n24078), .B(n24077), .Z(n24079) );
  AND U24714 ( .A(n24080), .B(n24079), .Z(n24118) );
  XOR U24715 ( .A(n24119), .B(n24118), .Z(c[1601]) );
  NANDN U24716 ( .A(n24082), .B(n24081), .Z(n24086) );
  NAND U24717 ( .A(n24084), .B(n24083), .Z(n24085) );
  NAND U24718 ( .A(n24086), .B(n24085), .Z(n24125) );
  NAND U24719 ( .A(b[0]), .B(a[586]), .Z(n24087) );
  XNOR U24720 ( .A(b[1]), .B(n24087), .Z(n24089) );
  NAND U24721 ( .A(n98), .B(a[585]), .Z(n24088) );
  AND U24722 ( .A(n24089), .B(n24088), .Z(n24142) );
  XOR U24723 ( .A(a[582]), .B(n42197), .Z(n24131) );
  NANDN U24724 ( .A(n24131), .B(n42173), .Z(n24092) );
  NANDN U24725 ( .A(n24090), .B(n42172), .Z(n24091) );
  NAND U24726 ( .A(n24092), .B(n24091), .Z(n24140) );
  NAND U24727 ( .A(b[7]), .B(a[578]), .Z(n24141) );
  XNOR U24728 ( .A(n24140), .B(n24141), .Z(n24143) );
  XOR U24729 ( .A(n24142), .B(n24143), .Z(n24149) );
  NANDN U24730 ( .A(n24093), .B(n42093), .Z(n24095) );
  XOR U24731 ( .A(n42134), .B(a[584]), .Z(n24134) );
  NANDN U24732 ( .A(n24134), .B(n42095), .Z(n24094) );
  NAND U24733 ( .A(n24095), .B(n24094), .Z(n24147) );
  NANDN U24734 ( .A(n24096), .B(n42231), .Z(n24098) );
  XOR U24735 ( .A(n210), .B(a[580]), .Z(n24137) );
  NANDN U24736 ( .A(n24137), .B(n42234), .Z(n24097) );
  AND U24737 ( .A(n24098), .B(n24097), .Z(n24146) );
  XNOR U24738 ( .A(n24147), .B(n24146), .Z(n24148) );
  XNOR U24739 ( .A(n24149), .B(n24148), .Z(n24153) );
  NANDN U24740 ( .A(n24100), .B(n24099), .Z(n24104) );
  NAND U24741 ( .A(n24102), .B(n24101), .Z(n24103) );
  AND U24742 ( .A(n24104), .B(n24103), .Z(n24152) );
  XOR U24743 ( .A(n24153), .B(n24152), .Z(n24154) );
  NANDN U24744 ( .A(n24106), .B(n24105), .Z(n24110) );
  NANDN U24745 ( .A(n24108), .B(n24107), .Z(n24109) );
  NAND U24746 ( .A(n24110), .B(n24109), .Z(n24155) );
  XOR U24747 ( .A(n24154), .B(n24155), .Z(n24122) );
  OR U24748 ( .A(n24112), .B(n24111), .Z(n24116) );
  NANDN U24749 ( .A(n24114), .B(n24113), .Z(n24115) );
  NAND U24750 ( .A(n24116), .B(n24115), .Z(n24123) );
  XNOR U24751 ( .A(n24122), .B(n24123), .Z(n24124) );
  XNOR U24752 ( .A(n24125), .B(n24124), .Z(n24158) );
  XNOR U24753 ( .A(n24158), .B(sreg[1602]), .Z(n24160) );
  NAND U24754 ( .A(n24117), .B(sreg[1601]), .Z(n24121) );
  OR U24755 ( .A(n24119), .B(n24118), .Z(n24120) );
  AND U24756 ( .A(n24121), .B(n24120), .Z(n24159) );
  XOR U24757 ( .A(n24160), .B(n24159), .Z(c[1602]) );
  NANDN U24758 ( .A(n24123), .B(n24122), .Z(n24127) );
  NAND U24759 ( .A(n24125), .B(n24124), .Z(n24126) );
  NAND U24760 ( .A(n24127), .B(n24126), .Z(n24166) );
  NAND U24761 ( .A(b[0]), .B(a[587]), .Z(n24128) );
  XNOR U24762 ( .A(b[1]), .B(n24128), .Z(n24130) );
  NAND U24763 ( .A(n98), .B(a[586]), .Z(n24129) );
  AND U24764 ( .A(n24130), .B(n24129), .Z(n24183) );
  XOR U24765 ( .A(a[583]), .B(n42197), .Z(n24172) );
  NANDN U24766 ( .A(n24172), .B(n42173), .Z(n24133) );
  NANDN U24767 ( .A(n24131), .B(n42172), .Z(n24132) );
  NAND U24768 ( .A(n24133), .B(n24132), .Z(n24181) );
  NAND U24769 ( .A(b[7]), .B(a[579]), .Z(n24182) );
  XNOR U24770 ( .A(n24181), .B(n24182), .Z(n24184) );
  XOR U24771 ( .A(n24183), .B(n24184), .Z(n24190) );
  NANDN U24772 ( .A(n24134), .B(n42093), .Z(n24136) );
  XOR U24773 ( .A(n42134), .B(a[585]), .Z(n24175) );
  NANDN U24774 ( .A(n24175), .B(n42095), .Z(n24135) );
  NAND U24775 ( .A(n24136), .B(n24135), .Z(n24188) );
  NANDN U24776 ( .A(n24137), .B(n42231), .Z(n24139) );
  XOR U24777 ( .A(n210), .B(a[581]), .Z(n24178) );
  NANDN U24778 ( .A(n24178), .B(n42234), .Z(n24138) );
  AND U24779 ( .A(n24139), .B(n24138), .Z(n24187) );
  XNOR U24780 ( .A(n24188), .B(n24187), .Z(n24189) );
  XNOR U24781 ( .A(n24190), .B(n24189), .Z(n24194) );
  NANDN U24782 ( .A(n24141), .B(n24140), .Z(n24145) );
  NAND U24783 ( .A(n24143), .B(n24142), .Z(n24144) );
  AND U24784 ( .A(n24145), .B(n24144), .Z(n24193) );
  XOR U24785 ( .A(n24194), .B(n24193), .Z(n24195) );
  NANDN U24786 ( .A(n24147), .B(n24146), .Z(n24151) );
  NANDN U24787 ( .A(n24149), .B(n24148), .Z(n24150) );
  NAND U24788 ( .A(n24151), .B(n24150), .Z(n24196) );
  XOR U24789 ( .A(n24195), .B(n24196), .Z(n24163) );
  OR U24790 ( .A(n24153), .B(n24152), .Z(n24157) );
  NANDN U24791 ( .A(n24155), .B(n24154), .Z(n24156) );
  NAND U24792 ( .A(n24157), .B(n24156), .Z(n24164) );
  XNOR U24793 ( .A(n24163), .B(n24164), .Z(n24165) );
  XNOR U24794 ( .A(n24166), .B(n24165), .Z(n24199) );
  XNOR U24795 ( .A(n24199), .B(sreg[1603]), .Z(n24201) );
  NAND U24796 ( .A(n24158), .B(sreg[1602]), .Z(n24162) );
  OR U24797 ( .A(n24160), .B(n24159), .Z(n24161) );
  AND U24798 ( .A(n24162), .B(n24161), .Z(n24200) );
  XOR U24799 ( .A(n24201), .B(n24200), .Z(c[1603]) );
  NANDN U24800 ( .A(n24164), .B(n24163), .Z(n24168) );
  NAND U24801 ( .A(n24166), .B(n24165), .Z(n24167) );
  NAND U24802 ( .A(n24168), .B(n24167), .Z(n24207) );
  NAND U24803 ( .A(b[0]), .B(a[588]), .Z(n24169) );
  XNOR U24804 ( .A(b[1]), .B(n24169), .Z(n24171) );
  NAND U24805 ( .A(n99), .B(a[587]), .Z(n24170) );
  AND U24806 ( .A(n24171), .B(n24170), .Z(n24224) );
  XOR U24807 ( .A(a[584]), .B(n42197), .Z(n24213) );
  NANDN U24808 ( .A(n24213), .B(n42173), .Z(n24174) );
  NANDN U24809 ( .A(n24172), .B(n42172), .Z(n24173) );
  NAND U24810 ( .A(n24174), .B(n24173), .Z(n24222) );
  NAND U24811 ( .A(b[7]), .B(a[580]), .Z(n24223) );
  XNOR U24812 ( .A(n24222), .B(n24223), .Z(n24225) );
  XOR U24813 ( .A(n24224), .B(n24225), .Z(n24231) );
  NANDN U24814 ( .A(n24175), .B(n42093), .Z(n24177) );
  XOR U24815 ( .A(n42134), .B(a[586]), .Z(n24216) );
  NANDN U24816 ( .A(n24216), .B(n42095), .Z(n24176) );
  NAND U24817 ( .A(n24177), .B(n24176), .Z(n24229) );
  NANDN U24818 ( .A(n24178), .B(n42231), .Z(n24180) );
  XOR U24819 ( .A(n210), .B(a[582]), .Z(n24219) );
  NANDN U24820 ( .A(n24219), .B(n42234), .Z(n24179) );
  AND U24821 ( .A(n24180), .B(n24179), .Z(n24228) );
  XNOR U24822 ( .A(n24229), .B(n24228), .Z(n24230) );
  XNOR U24823 ( .A(n24231), .B(n24230), .Z(n24235) );
  NANDN U24824 ( .A(n24182), .B(n24181), .Z(n24186) );
  NAND U24825 ( .A(n24184), .B(n24183), .Z(n24185) );
  AND U24826 ( .A(n24186), .B(n24185), .Z(n24234) );
  XOR U24827 ( .A(n24235), .B(n24234), .Z(n24236) );
  NANDN U24828 ( .A(n24188), .B(n24187), .Z(n24192) );
  NANDN U24829 ( .A(n24190), .B(n24189), .Z(n24191) );
  NAND U24830 ( .A(n24192), .B(n24191), .Z(n24237) );
  XOR U24831 ( .A(n24236), .B(n24237), .Z(n24204) );
  OR U24832 ( .A(n24194), .B(n24193), .Z(n24198) );
  NANDN U24833 ( .A(n24196), .B(n24195), .Z(n24197) );
  NAND U24834 ( .A(n24198), .B(n24197), .Z(n24205) );
  XNOR U24835 ( .A(n24204), .B(n24205), .Z(n24206) );
  XNOR U24836 ( .A(n24207), .B(n24206), .Z(n24240) );
  XNOR U24837 ( .A(n24240), .B(sreg[1604]), .Z(n24242) );
  NAND U24838 ( .A(n24199), .B(sreg[1603]), .Z(n24203) );
  OR U24839 ( .A(n24201), .B(n24200), .Z(n24202) );
  AND U24840 ( .A(n24203), .B(n24202), .Z(n24241) );
  XOR U24841 ( .A(n24242), .B(n24241), .Z(c[1604]) );
  NANDN U24842 ( .A(n24205), .B(n24204), .Z(n24209) );
  NAND U24843 ( .A(n24207), .B(n24206), .Z(n24208) );
  NAND U24844 ( .A(n24209), .B(n24208), .Z(n24248) );
  NAND U24845 ( .A(b[0]), .B(a[589]), .Z(n24210) );
  XNOR U24846 ( .A(b[1]), .B(n24210), .Z(n24212) );
  NAND U24847 ( .A(n99), .B(a[588]), .Z(n24211) );
  AND U24848 ( .A(n24212), .B(n24211), .Z(n24265) );
  XOR U24849 ( .A(a[585]), .B(n42197), .Z(n24254) );
  NANDN U24850 ( .A(n24254), .B(n42173), .Z(n24215) );
  NANDN U24851 ( .A(n24213), .B(n42172), .Z(n24214) );
  NAND U24852 ( .A(n24215), .B(n24214), .Z(n24263) );
  NAND U24853 ( .A(b[7]), .B(a[581]), .Z(n24264) );
  XNOR U24854 ( .A(n24263), .B(n24264), .Z(n24266) );
  XOR U24855 ( .A(n24265), .B(n24266), .Z(n24272) );
  NANDN U24856 ( .A(n24216), .B(n42093), .Z(n24218) );
  XOR U24857 ( .A(n42134), .B(a[587]), .Z(n24257) );
  NANDN U24858 ( .A(n24257), .B(n42095), .Z(n24217) );
  NAND U24859 ( .A(n24218), .B(n24217), .Z(n24270) );
  NANDN U24860 ( .A(n24219), .B(n42231), .Z(n24221) );
  XOR U24861 ( .A(n210), .B(a[583]), .Z(n24260) );
  NANDN U24862 ( .A(n24260), .B(n42234), .Z(n24220) );
  AND U24863 ( .A(n24221), .B(n24220), .Z(n24269) );
  XNOR U24864 ( .A(n24270), .B(n24269), .Z(n24271) );
  XNOR U24865 ( .A(n24272), .B(n24271), .Z(n24276) );
  NANDN U24866 ( .A(n24223), .B(n24222), .Z(n24227) );
  NAND U24867 ( .A(n24225), .B(n24224), .Z(n24226) );
  AND U24868 ( .A(n24227), .B(n24226), .Z(n24275) );
  XOR U24869 ( .A(n24276), .B(n24275), .Z(n24277) );
  NANDN U24870 ( .A(n24229), .B(n24228), .Z(n24233) );
  NANDN U24871 ( .A(n24231), .B(n24230), .Z(n24232) );
  NAND U24872 ( .A(n24233), .B(n24232), .Z(n24278) );
  XOR U24873 ( .A(n24277), .B(n24278), .Z(n24245) );
  OR U24874 ( .A(n24235), .B(n24234), .Z(n24239) );
  NANDN U24875 ( .A(n24237), .B(n24236), .Z(n24238) );
  NAND U24876 ( .A(n24239), .B(n24238), .Z(n24246) );
  XNOR U24877 ( .A(n24245), .B(n24246), .Z(n24247) );
  XNOR U24878 ( .A(n24248), .B(n24247), .Z(n24281) );
  XNOR U24879 ( .A(n24281), .B(sreg[1605]), .Z(n24283) );
  NAND U24880 ( .A(n24240), .B(sreg[1604]), .Z(n24244) );
  OR U24881 ( .A(n24242), .B(n24241), .Z(n24243) );
  AND U24882 ( .A(n24244), .B(n24243), .Z(n24282) );
  XOR U24883 ( .A(n24283), .B(n24282), .Z(c[1605]) );
  NANDN U24884 ( .A(n24246), .B(n24245), .Z(n24250) );
  NAND U24885 ( .A(n24248), .B(n24247), .Z(n24249) );
  NAND U24886 ( .A(n24250), .B(n24249), .Z(n24289) );
  NAND U24887 ( .A(b[0]), .B(a[590]), .Z(n24251) );
  XNOR U24888 ( .A(b[1]), .B(n24251), .Z(n24253) );
  NAND U24889 ( .A(n99), .B(a[589]), .Z(n24252) );
  AND U24890 ( .A(n24253), .B(n24252), .Z(n24306) );
  XOR U24891 ( .A(a[586]), .B(n42197), .Z(n24295) );
  NANDN U24892 ( .A(n24295), .B(n42173), .Z(n24256) );
  NANDN U24893 ( .A(n24254), .B(n42172), .Z(n24255) );
  NAND U24894 ( .A(n24256), .B(n24255), .Z(n24304) );
  NAND U24895 ( .A(b[7]), .B(a[582]), .Z(n24305) );
  XNOR U24896 ( .A(n24304), .B(n24305), .Z(n24307) );
  XOR U24897 ( .A(n24306), .B(n24307), .Z(n24313) );
  NANDN U24898 ( .A(n24257), .B(n42093), .Z(n24259) );
  XOR U24899 ( .A(n42134), .B(a[588]), .Z(n24298) );
  NANDN U24900 ( .A(n24298), .B(n42095), .Z(n24258) );
  NAND U24901 ( .A(n24259), .B(n24258), .Z(n24311) );
  NANDN U24902 ( .A(n24260), .B(n42231), .Z(n24262) );
  XOR U24903 ( .A(n210), .B(a[584]), .Z(n24301) );
  NANDN U24904 ( .A(n24301), .B(n42234), .Z(n24261) );
  AND U24905 ( .A(n24262), .B(n24261), .Z(n24310) );
  XNOR U24906 ( .A(n24311), .B(n24310), .Z(n24312) );
  XNOR U24907 ( .A(n24313), .B(n24312), .Z(n24317) );
  NANDN U24908 ( .A(n24264), .B(n24263), .Z(n24268) );
  NAND U24909 ( .A(n24266), .B(n24265), .Z(n24267) );
  AND U24910 ( .A(n24268), .B(n24267), .Z(n24316) );
  XOR U24911 ( .A(n24317), .B(n24316), .Z(n24318) );
  NANDN U24912 ( .A(n24270), .B(n24269), .Z(n24274) );
  NANDN U24913 ( .A(n24272), .B(n24271), .Z(n24273) );
  NAND U24914 ( .A(n24274), .B(n24273), .Z(n24319) );
  XOR U24915 ( .A(n24318), .B(n24319), .Z(n24286) );
  OR U24916 ( .A(n24276), .B(n24275), .Z(n24280) );
  NANDN U24917 ( .A(n24278), .B(n24277), .Z(n24279) );
  NAND U24918 ( .A(n24280), .B(n24279), .Z(n24287) );
  XNOR U24919 ( .A(n24286), .B(n24287), .Z(n24288) );
  XNOR U24920 ( .A(n24289), .B(n24288), .Z(n24322) );
  XNOR U24921 ( .A(n24322), .B(sreg[1606]), .Z(n24324) );
  NAND U24922 ( .A(n24281), .B(sreg[1605]), .Z(n24285) );
  OR U24923 ( .A(n24283), .B(n24282), .Z(n24284) );
  AND U24924 ( .A(n24285), .B(n24284), .Z(n24323) );
  XOR U24925 ( .A(n24324), .B(n24323), .Z(c[1606]) );
  NANDN U24926 ( .A(n24287), .B(n24286), .Z(n24291) );
  NAND U24927 ( .A(n24289), .B(n24288), .Z(n24290) );
  NAND U24928 ( .A(n24291), .B(n24290), .Z(n24330) );
  NAND U24929 ( .A(b[0]), .B(a[591]), .Z(n24292) );
  XNOR U24930 ( .A(b[1]), .B(n24292), .Z(n24294) );
  NAND U24931 ( .A(n99), .B(a[590]), .Z(n24293) );
  AND U24932 ( .A(n24294), .B(n24293), .Z(n24347) );
  XOR U24933 ( .A(a[587]), .B(n42197), .Z(n24336) );
  NANDN U24934 ( .A(n24336), .B(n42173), .Z(n24297) );
  NANDN U24935 ( .A(n24295), .B(n42172), .Z(n24296) );
  NAND U24936 ( .A(n24297), .B(n24296), .Z(n24345) );
  NAND U24937 ( .A(b[7]), .B(a[583]), .Z(n24346) );
  XNOR U24938 ( .A(n24345), .B(n24346), .Z(n24348) );
  XOR U24939 ( .A(n24347), .B(n24348), .Z(n24354) );
  NANDN U24940 ( .A(n24298), .B(n42093), .Z(n24300) );
  XOR U24941 ( .A(n42134), .B(a[589]), .Z(n24339) );
  NANDN U24942 ( .A(n24339), .B(n42095), .Z(n24299) );
  NAND U24943 ( .A(n24300), .B(n24299), .Z(n24352) );
  NANDN U24944 ( .A(n24301), .B(n42231), .Z(n24303) );
  XOR U24945 ( .A(n210), .B(a[585]), .Z(n24342) );
  NANDN U24946 ( .A(n24342), .B(n42234), .Z(n24302) );
  AND U24947 ( .A(n24303), .B(n24302), .Z(n24351) );
  XNOR U24948 ( .A(n24352), .B(n24351), .Z(n24353) );
  XNOR U24949 ( .A(n24354), .B(n24353), .Z(n24358) );
  NANDN U24950 ( .A(n24305), .B(n24304), .Z(n24309) );
  NAND U24951 ( .A(n24307), .B(n24306), .Z(n24308) );
  AND U24952 ( .A(n24309), .B(n24308), .Z(n24357) );
  XOR U24953 ( .A(n24358), .B(n24357), .Z(n24359) );
  NANDN U24954 ( .A(n24311), .B(n24310), .Z(n24315) );
  NANDN U24955 ( .A(n24313), .B(n24312), .Z(n24314) );
  NAND U24956 ( .A(n24315), .B(n24314), .Z(n24360) );
  XOR U24957 ( .A(n24359), .B(n24360), .Z(n24327) );
  OR U24958 ( .A(n24317), .B(n24316), .Z(n24321) );
  NANDN U24959 ( .A(n24319), .B(n24318), .Z(n24320) );
  NAND U24960 ( .A(n24321), .B(n24320), .Z(n24328) );
  XNOR U24961 ( .A(n24327), .B(n24328), .Z(n24329) );
  XNOR U24962 ( .A(n24330), .B(n24329), .Z(n24363) );
  XNOR U24963 ( .A(n24363), .B(sreg[1607]), .Z(n24365) );
  NAND U24964 ( .A(n24322), .B(sreg[1606]), .Z(n24326) );
  OR U24965 ( .A(n24324), .B(n24323), .Z(n24325) );
  AND U24966 ( .A(n24326), .B(n24325), .Z(n24364) );
  XOR U24967 ( .A(n24365), .B(n24364), .Z(c[1607]) );
  NANDN U24968 ( .A(n24328), .B(n24327), .Z(n24332) );
  NAND U24969 ( .A(n24330), .B(n24329), .Z(n24331) );
  NAND U24970 ( .A(n24332), .B(n24331), .Z(n24371) );
  NAND U24971 ( .A(b[0]), .B(a[592]), .Z(n24333) );
  XNOR U24972 ( .A(b[1]), .B(n24333), .Z(n24335) );
  NAND U24973 ( .A(n99), .B(a[591]), .Z(n24334) );
  AND U24974 ( .A(n24335), .B(n24334), .Z(n24388) );
  XOR U24975 ( .A(a[588]), .B(n42197), .Z(n24377) );
  NANDN U24976 ( .A(n24377), .B(n42173), .Z(n24338) );
  NANDN U24977 ( .A(n24336), .B(n42172), .Z(n24337) );
  NAND U24978 ( .A(n24338), .B(n24337), .Z(n24386) );
  NAND U24979 ( .A(b[7]), .B(a[584]), .Z(n24387) );
  XNOR U24980 ( .A(n24386), .B(n24387), .Z(n24389) );
  XOR U24981 ( .A(n24388), .B(n24389), .Z(n24395) );
  NANDN U24982 ( .A(n24339), .B(n42093), .Z(n24341) );
  XOR U24983 ( .A(n42134), .B(a[590]), .Z(n24380) );
  NANDN U24984 ( .A(n24380), .B(n42095), .Z(n24340) );
  NAND U24985 ( .A(n24341), .B(n24340), .Z(n24393) );
  NANDN U24986 ( .A(n24342), .B(n42231), .Z(n24344) );
  XOR U24987 ( .A(n210), .B(a[586]), .Z(n24383) );
  NANDN U24988 ( .A(n24383), .B(n42234), .Z(n24343) );
  AND U24989 ( .A(n24344), .B(n24343), .Z(n24392) );
  XNOR U24990 ( .A(n24393), .B(n24392), .Z(n24394) );
  XNOR U24991 ( .A(n24395), .B(n24394), .Z(n24399) );
  NANDN U24992 ( .A(n24346), .B(n24345), .Z(n24350) );
  NAND U24993 ( .A(n24348), .B(n24347), .Z(n24349) );
  AND U24994 ( .A(n24350), .B(n24349), .Z(n24398) );
  XOR U24995 ( .A(n24399), .B(n24398), .Z(n24400) );
  NANDN U24996 ( .A(n24352), .B(n24351), .Z(n24356) );
  NANDN U24997 ( .A(n24354), .B(n24353), .Z(n24355) );
  NAND U24998 ( .A(n24356), .B(n24355), .Z(n24401) );
  XOR U24999 ( .A(n24400), .B(n24401), .Z(n24368) );
  OR U25000 ( .A(n24358), .B(n24357), .Z(n24362) );
  NANDN U25001 ( .A(n24360), .B(n24359), .Z(n24361) );
  NAND U25002 ( .A(n24362), .B(n24361), .Z(n24369) );
  XNOR U25003 ( .A(n24368), .B(n24369), .Z(n24370) );
  XNOR U25004 ( .A(n24371), .B(n24370), .Z(n24404) );
  XNOR U25005 ( .A(n24404), .B(sreg[1608]), .Z(n24406) );
  NAND U25006 ( .A(n24363), .B(sreg[1607]), .Z(n24367) );
  OR U25007 ( .A(n24365), .B(n24364), .Z(n24366) );
  AND U25008 ( .A(n24367), .B(n24366), .Z(n24405) );
  XOR U25009 ( .A(n24406), .B(n24405), .Z(c[1608]) );
  NANDN U25010 ( .A(n24369), .B(n24368), .Z(n24373) );
  NAND U25011 ( .A(n24371), .B(n24370), .Z(n24372) );
  NAND U25012 ( .A(n24373), .B(n24372), .Z(n24412) );
  NAND U25013 ( .A(b[0]), .B(a[593]), .Z(n24374) );
  XNOR U25014 ( .A(b[1]), .B(n24374), .Z(n24376) );
  NAND U25015 ( .A(n99), .B(a[592]), .Z(n24375) );
  AND U25016 ( .A(n24376), .B(n24375), .Z(n24429) );
  XOR U25017 ( .A(a[589]), .B(n42197), .Z(n24418) );
  NANDN U25018 ( .A(n24418), .B(n42173), .Z(n24379) );
  NANDN U25019 ( .A(n24377), .B(n42172), .Z(n24378) );
  NAND U25020 ( .A(n24379), .B(n24378), .Z(n24427) );
  NAND U25021 ( .A(b[7]), .B(a[585]), .Z(n24428) );
  XNOR U25022 ( .A(n24427), .B(n24428), .Z(n24430) );
  XOR U25023 ( .A(n24429), .B(n24430), .Z(n24436) );
  NANDN U25024 ( .A(n24380), .B(n42093), .Z(n24382) );
  XOR U25025 ( .A(n42134), .B(a[591]), .Z(n24421) );
  NANDN U25026 ( .A(n24421), .B(n42095), .Z(n24381) );
  NAND U25027 ( .A(n24382), .B(n24381), .Z(n24434) );
  NANDN U25028 ( .A(n24383), .B(n42231), .Z(n24385) );
  XOR U25029 ( .A(n211), .B(a[587]), .Z(n24424) );
  NANDN U25030 ( .A(n24424), .B(n42234), .Z(n24384) );
  AND U25031 ( .A(n24385), .B(n24384), .Z(n24433) );
  XNOR U25032 ( .A(n24434), .B(n24433), .Z(n24435) );
  XNOR U25033 ( .A(n24436), .B(n24435), .Z(n24440) );
  NANDN U25034 ( .A(n24387), .B(n24386), .Z(n24391) );
  NAND U25035 ( .A(n24389), .B(n24388), .Z(n24390) );
  AND U25036 ( .A(n24391), .B(n24390), .Z(n24439) );
  XOR U25037 ( .A(n24440), .B(n24439), .Z(n24441) );
  NANDN U25038 ( .A(n24393), .B(n24392), .Z(n24397) );
  NANDN U25039 ( .A(n24395), .B(n24394), .Z(n24396) );
  NAND U25040 ( .A(n24397), .B(n24396), .Z(n24442) );
  XOR U25041 ( .A(n24441), .B(n24442), .Z(n24409) );
  OR U25042 ( .A(n24399), .B(n24398), .Z(n24403) );
  NANDN U25043 ( .A(n24401), .B(n24400), .Z(n24402) );
  NAND U25044 ( .A(n24403), .B(n24402), .Z(n24410) );
  XNOR U25045 ( .A(n24409), .B(n24410), .Z(n24411) );
  XNOR U25046 ( .A(n24412), .B(n24411), .Z(n24445) );
  XNOR U25047 ( .A(n24445), .B(sreg[1609]), .Z(n24447) );
  NAND U25048 ( .A(n24404), .B(sreg[1608]), .Z(n24408) );
  OR U25049 ( .A(n24406), .B(n24405), .Z(n24407) );
  AND U25050 ( .A(n24408), .B(n24407), .Z(n24446) );
  XOR U25051 ( .A(n24447), .B(n24446), .Z(c[1609]) );
  NANDN U25052 ( .A(n24410), .B(n24409), .Z(n24414) );
  NAND U25053 ( .A(n24412), .B(n24411), .Z(n24413) );
  NAND U25054 ( .A(n24414), .B(n24413), .Z(n24453) );
  NAND U25055 ( .A(b[0]), .B(a[594]), .Z(n24415) );
  XNOR U25056 ( .A(b[1]), .B(n24415), .Z(n24417) );
  NAND U25057 ( .A(n99), .B(a[593]), .Z(n24416) );
  AND U25058 ( .A(n24417), .B(n24416), .Z(n24470) );
  XOR U25059 ( .A(a[590]), .B(n42197), .Z(n24459) );
  NANDN U25060 ( .A(n24459), .B(n42173), .Z(n24420) );
  NANDN U25061 ( .A(n24418), .B(n42172), .Z(n24419) );
  NAND U25062 ( .A(n24420), .B(n24419), .Z(n24468) );
  NAND U25063 ( .A(b[7]), .B(a[586]), .Z(n24469) );
  XNOR U25064 ( .A(n24468), .B(n24469), .Z(n24471) );
  XOR U25065 ( .A(n24470), .B(n24471), .Z(n24477) );
  NANDN U25066 ( .A(n24421), .B(n42093), .Z(n24423) );
  XOR U25067 ( .A(n42134), .B(a[592]), .Z(n24462) );
  NANDN U25068 ( .A(n24462), .B(n42095), .Z(n24422) );
  NAND U25069 ( .A(n24423), .B(n24422), .Z(n24475) );
  NANDN U25070 ( .A(n24424), .B(n42231), .Z(n24426) );
  XOR U25071 ( .A(n211), .B(a[588]), .Z(n24465) );
  NANDN U25072 ( .A(n24465), .B(n42234), .Z(n24425) );
  AND U25073 ( .A(n24426), .B(n24425), .Z(n24474) );
  XNOR U25074 ( .A(n24475), .B(n24474), .Z(n24476) );
  XNOR U25075 ( .A(n24477), .B(n24476), .Z(n24481) );
  NANDN U25076 ( .A(n24428), .B(n24427), .Z(n24432) );
  NAND U25077 ( .A(n24430), .B(n24429), .Z(n24431) );
  AND U25078 ( .A(n24432), .B(n24431), .Z(n24480) );
  XOR U25079 ( .A(n24481), .B(n24480), .Z(n24482) );
  NANDN U25080 ( .A(n24434), .B(n24433), .Z(n24438) );
  NANDN U25081 ( .A(n24436), .B(n24435), .Z(n24437) );
  NAND U25082 ( .A(n24438), .B(n24437), .Z(n24483) );
  XOR U25083 ( .A(n24482), .B(n24483), .Z(n24450) );
  OR U25084 ( .A(n24440), .B(n24439), .Z(n24444) );
  NANDN U25085 ( .A(n24442), .B(n24441), .Z(n24443) );
  NAND U25086 ( .A(n24444), .B(n24443), .Z(n24451) );
  XNOR U25087 ( .A(n24450), .B(n24451), .Z(n24452) );
  XNOR U25088 ( .A(n24453), .B(n24452), .Z(n24486) );
  XNOR U25089 ( .A(n24486), .B(sreg[1610]), .Z(n24488) );
  NAND U25090 ( .A(n24445), .B(sreg[1609]), .Z(n24449) );
  OR U25091 ( .A(n24447), .B(n24446), .Z(n24448) );
  AND U25092 ( .A(n24449), .B(n24448), .Z(n24487) );
  XOR U25093 ( .A(n24488), .B(n24487), .Z(c[1610]) );
  NANDN U25094 ( .A(n24451), .B(n24450), .Z(n24455) );
  NAND U25095 ( .A(n24453), .B(n24452), .Z(n24454) );
  NAND U25096 ( .A(n24455), .B(n24454), .Z(n24494) );
  NAND U25097 ( .A(b[0]), .B(a[595]), .Z(n24456) );
  XNOR U25098 ( .A(b[1]), .B(n24456), .Z(n24458) );
  NAND U25099 ( .A(n100), .B(a[594]), .Z(n24457) );
  AND U25100 ( .A(n24458), .B(n24457), .Z(n24511) );
  XOR U25101 ( .A(a[591]), .B(n42197), .Z(n24500) );
  NANDN U25102 ( .A(n24500), .B(n42173), .Z(n24461) );
  NANDN U25103 ( .A(n24459), .B(n42172), .Z(n24460) );
  NAND U25104 ( .A(n24461), .B(n24460), .Z(n24509) );
  NAND U25105 ( .A(b[7]), .B(a[587]), .Z(n24510) );
  XNOR U25106 ( .A(n24509), .B(n24510), .Z(n24512) );
  XOR U25107 ( .A(n24511), .B(n24512), .Z(n24518) );
  NANDN U25108 ( .A(n24462), .B(n42093), .Z(n24464) );
  XOR U25109 ( .A(n42134), .B(a[593]), .Z(n24503) );
  NANDN U25110 ( .A(n24503), .B(n42095), .Z(n24463) );
  NAND U25111 ( .A(n24464), .B(n24463), .Z(n24516) );
  NANDN U25112 ( .A(n24465), .B(n42231), .Z(n24467) );
  XOR U25113 ( .A(n211), .B(a[589]), .Z(n24506) );
  NANDN U25114 ( .A(n24506), .B(n42234), .Z(n24466) );
  AND U25115 ( .A(n24467), .B(n24466), .Z(n24515) );
  XNOR U25116 ( .A(n24516), .B(n24515), .Z(n24517) );
  XNOR U25117 ( .A(n24518), .B(n24517), .Z(n24522) );
  NANDN U25118 ( .A(n24469), .B(n24468), .Z(n24473) );
  NAND U25119 ( .A(n24471), .B(n24470), .Z(n24472) );
  AND U25120 ( .A(n24473), .B(n24472), .Z(n24521) );
  XOR U25121 ( .A(n24522), .B(n24521), .Z(n24523) );
  NANDN U25122 ( .A(n24475), .B(n24474), .Z(n24479) );
  NANDN U25123 ( .A(n24477), .B(n24476), .Z(n24478) );
  NAND U25124 ( .A(n24479), .B(n24478), .Z(n24524) );
  XOR U25125 ( .A(n24523), .B(n24524), .Z(n24491) );
  OR U25126 ( .A(n24481), .B(n24480), .Z(n24485) );
  NANDN U25127 ( .A(n24483), .B(n24482), .Z(n24484) );
  NAND U25128 ( .A(n24485), .B(n24484), .Z(n24492) );
  XNOR U25129 ( .A(n24491), .B(n24492), .Z(n24493) );
  XNOR U25130 ( .A(n24494), .B(n24493), .Z(n24527) );
  XNOR U25131 ( .A(n24527), .B(sreg[1611]), .Z(n24529) );
  NAND U25132 ( .A(n24486), .B(sreg[1610]), .Z(n24490) );
  OR U25133 ( .A(n24488), .B(n24487), .Z(n24489) );
  AND U25134 ( .A(n24490), .B(n24489), .Z(n24528) );
  XOR U25135 ( .A(n24529), .B(n24528), .Z(c[1611]) );
  NANDN U25136 ( .A(n24492), .B(n24491), .Z(n24496) );
  NAND U25137 ( .A(n24494), .B(n24493), .Z(n24495) );
  NAND U25138 ( .A(n24496), .B(n24495), .Z(n24535) );
  NAND U25139 ( .A(b[0]), .B(a[596]), .Z(n24497) );
  XNOR U25140 ( .A(b[1]), .B(n24497), .Z(n24499) );
  NAND U25141 ( .A(n100), .B(a[595]), .Z(n24498) );
  AND U25142 ( .A(n24499), .B(n24498), .Z(n24552) );
  XOR U25143 ( .A(a[592]), .B(n42197), .Z(n24541) );
  NANDN U25144 ( .A(n24541), .B(n42173), .Z(n24502) );
  NANDN U25145 ( .A(n24500), .B(n42172), .Z(n24501) );
  NAND U25146 ( .A(n24502), .B(n24501), .Z(n24550) );
  NAND U25147 ( .A(b[7]), .B(a[588]), .Z(n24551) );
  XNOR U25148 ( .A(n24550), .B(n24551), .Z(n24553) );
  XOR U25149 ( .A(n24552), .B(n24553), .Z(n24559) );
  NANDN U25150 ( .A(n24503), .B(n42093), .Z(n24505) );
  XOR U25151 ( .A(n42134), .B(a[594]), .Z(n24544) );
  NANDN U25152 ( .A(n24544), .B(n42095), .Z(n24504) );
  NAND U25153 ( .A(n24505), .B(n24504), .Z(n24557) );
  NANDN U25154 ( .A(n24506), .B(n42231), .Z(n24508) );
  XOR U25155 ( .A(n211), .B(a[590]), .Z(n24547) );
  NANDN U25156 ( .A(n24547), .B(n42234), .Z(n24507) );
  AND U25157 ( .A(n24508), .B(n24507), .Z(n24556) );
  XNOR U25158 ( .A(n24557), .B(n24556), .Z(n24558) );
  XNOR U25159 ( .A(n24559), .B(n24558), .Z(n24563) );
  NANDN U25160 ( .A(n24510), .B(n24509), .Z(n24514) );
  NAND U25161 ( .A(n24512), .B(n24511), .Z(n24513) );
  AND U25162 ( .A(n24514), .B(n24513), .Z(n24562) );
  XOR U25163 ( .A(n24563), .B(n24562), .Z(n24564) );
  NANDN U25164 ( .A(n24516), .B(n24515), .Z(n24520) );
  NANDN U25165 ( .A(n24518), .B(n24517), .Z(n24519) );
  NAND U25166 ( .A(n24520), .B(n24519), .Z(n24565) );
  XOR U25167 ( .A(n24564), .B(n24565), .Z(n24532) );
  OR U25168 ( .A(n24522), .B(n24521), .Z(n24526) );
  NANDN U25169 ( .A(n24524), .B(n24523), .Z(n24525) );
  NAND U25170 ( .A(n24526), .B(n24525), .Z(n24533) );
  XNOR U25171 ( .A(n24532), .B(n24533), .Z(n24534) );
  XNOR U25172 ( .A(n24535), .B(n24534), .Z(n24568) );
  XNOR U25173 ( .A(n24568), .B(sreg[1612]), .Z(n24570) );
  NAND U25174 ( .A(n24527), .B(sreg[1611]), .Z(n24531) );
  OR U25175 ( .A(n24529), .B(n24528), .Z(n24530) );
  AND U25176 ( .A(n24531), .B(n24530), .Z(n24569) );
  XOR U25177 ( .A(n24570), .B(n24569), .Z(c[1612]) );
  NANDN U25178 ( .A(n24533), .B(n24532), .Z(n24537) );
  NAND U25179 ( .A(n24535), .B(n24534), .Z(n24536) );
  NAND U25180 ( .A(n24537), .B(n24536), .Z(n24576) );
  NAND U25181 ( .A(b[0]), .B(a[597]), .Z(n24538) );
  XNOR U25182 ( .A(b[1]), .B(n24538), .Z(n24540) );
  NAND U25183 ( .A(n100), .B(a[596]), .Z(n24539) );
  AND U25184 ( .A(n24540), .B(n24539), .Z(n24593) );
  XOR U25185 ( .A(a[593]), .B(n42197), .Z(n24582) );
  NANDN U25186 ( .A(n24582), .B(n42173), .Z(n24543) );
  NANDN U25187 ( .A(n24541), .B(n42172), .Z(n24542) );
  NAND U25188 ( .A(n24543), .B(n24542), .Z(n24591) );
  NAND U25189 ( .A(b[7]), .B(a[589]), .Z(n24592) );
  XNOR U25190 ( .A(n24591), .B(n24592), .Z(n24594) );
  XOR U25191 ( .A(n24593), .B(n24594), .Z(n24600) );
  NANDN U25192 ( .A(n24544), .B(n42093), .Z(n24546) );
  XOR U25193 ( .A(n42134), .B(a[595]), .Z(n24585) );
  NANDN U25194 ( .A(n24585), .B(n42095), .Z(n24545) );
  NAND U25195 ( .A(n24546), .B(n24545), .Z(n24598) );
  NANDN U25196 ( .A(n24547), .B(n42231), .Z(n24549) );
  XOR U25197 ( .A(n211), .B(a[591]), .Z(n24588) );
  NANDN U25198 ( .A(n24588), .B(n42234), .Z(n24548) );
  AND U25199 ( .A(n24549), .B(n24548), .Z(n24597) );
  XNOR U25200 ( .A(n24598), .B(n24597), .Z(n24599) );
  XNOR U25201 ( .A(n24600), .B(n24599), .Z(n24604) );
  NANDN U25202 ( .A(n24551), .B(n24550), .Z(n24555) );
  NAND U25203 ( .A(n24553), .B(n24552), .Z(n24554) );
  AND U25204 ( .A(n24555), .B(n24554), .Z(n24603) );
  XOR U25205 ( .A(n24604), .B(n24603), .Z(n24605) );
  NANDN U25206 ( .A(n24557), .B(n24556), .Z(n24561) );
  NANDN U25207 ( .A(n24559), .B(n24558), .Z(n24560) );
  NAND U25208 ( .A(n24561), .B(n24560), .Z(n24606) );
  XOR U25209 ( .A(n24605), .B(n24606), .Z(n24573) );
  OR U25210 ( .A(n24563), .B(n24562), .Z(n24567) );
  NANDN U25211 ( .A(n24565), .B(n24564), .Z(n24566) );
  NAND U25212 ( .A(n24567), .B(n24566), .Z(n24574) );
  XNOR U25213 ( .A(n24573), .B(n24574), .Z(n24575) );
  XNOR U25214 ( .A(n24576), .B(n24575), .Z(n24609) );
  XNOR U25215 ( .A(n24609), .B(sreg[1613]), .Z(n24611) );
  NAND U25216 ( .A(n24568), .B(sreg[1612]), .Z(n24572) );
  OR U25217 ( .A(n24570), .B(n24569), .Z(n24571) );
  AND U25218 ( .A(n24572), .B(n24571), .Z(n24610) );
  XOR U25219 ( .A(n24611), .B(n24610), .Z(c[1613]) );
  NANDN U25220 ( .A(n24574), .B(n24573), .Z(n24578) );
  NAND U25221 ( .A(n24576), .B(n24575), .Z(n24577) );
  NAND U25222 ( .A(n24578), .B(n24577), .Z(n24617) );
  NAND U25223 ( .A(b[0]), .B(a[598]), .Z(n24579) );
  XNOR U25224 ( .A(b[1]), .B(n24579), .Z(n24581) );
  NAND U25225 ( .A(n100), .B(a[597]), .Z(n24580) );
  AND U25226 ( .A(n24581), .B(n24580), .Z(n24634) );
  XOR U25227 ( .A(a[594]), .B(n42197), .Z(n24623) );
  NANDN U25228 ( .A(n24623), .B(n42173), .Z(n24584) );
  NANDN U25229 ( .A(n24582), .B(n42172), .Z(n24583) );
  NAND U25230 ( .A(n24584), .B(n24583), .Z(n24632) );
  NAND U25231 ( .A(b[7]), .B(a[590]), .Z(n24633) );
  XNOR U25232 ( .A(n24632), .B(n24633), .Z(n24635) );
  XOR U25233 ( .A(n24634), .B(n24635), .Z(n24641) );
  NANDN U25234 ( .A(n24585), .B(n42093), .Z(n24587) );
  XOR U25235 ( .A(n42134), .B(a[596]), .Z(n24626) );
  NANDN U25236 ( .A(n24626), .B(n42095), .Z(n24586) );
  NAND U25237 ( .A(n24587), .B(n24586), .Z(n24639) );
  NANDN U25238 ( .A(n24588), .B(n42231), .Z(n24590) );
  XOR U25239 ( .A(n211), .B(a[592]), .Z(n24629) );
  NANDN U25240 ( .A(n24629), .B(n42234), .Z(n24589) );
  AND U25241 ( .A(n24590), .B(n24589), .Z(n24638) );
  XNOR U25242 ( .A(n24639), .B(n24638), .Z(n24640) );
  XNOR U25243 ( .A(n24641), .B(n24640), .Z(n24645) );
  NANDN U25244 ( .A(n24592), .B(n24591), .Z(n24596) );
  NAND U25245 ( .A(n24594), .B(n24593), .Z(n24595) );
  AND U25246 ( .A(n24596), .B(n24595), .Z(n24644) );
  XOR U25247 ( .A(n24645), .B(n24644), .Z(n24646) );
  NANDN U25248 ( .A(n24598), .B(n24597), .Z(n24602) );
  NANDN U25249 ( .A(n24600), .B(n24599), .Z(n24601) );
  NAND U25250 ( .A(n24602), .B(n24601), .Z(n24647) );
  XOR U25251 ( .A(n24646), .B(n24647), .Z(n24614) );
  OR U25252 ( .A(n24604), .B(n24603), .Z(n24608) );
  NANDN U25253 ( .A(n24606), .B(n24605), .Z(n24607) );
  NAND U25254 ( .A(n24608), .B(n24607), .Z(n24615) );
  XNOR U25255 ( .A(n24614), .B(n24615), .Z(n24616) );
  XNOR U25256 ( .A(n24617), .B(n24616), .Z(n24650) );
  XNOR U25257 ( .A(n24650), .B(sreg[1614]), .Z(n24652) );
  NAND U25258 ( .A(n24609), .B(sreg[1613]), .Z(n24613) );
  OR U25259 ( .A(n24611), .B(n24610), .Z(n24612) );
  AND U25260 ( .A(n24613), .B(n24612), .Z(n24651) );
  XOR U25261 ( .A(n24652), .B(n24651), .Z(c[1614]) );
  NANDN U25262 ( .A(n24615), .B(n24614), .Z(n24619) );
  NAND U25263 ( .A(n24617), .B(n24616), .Z(n24618) );
  NAND U25264 ( .A(n24619), .B(n24618), .Z(n24658) );
  NAND U25265 ( .A(b[0]), .B(a[599]), .Z(n24620) );
  XNOR U25266 ( .A(b[1]), .B(n24620), .Z(n24622) );
  NAND U25267 ( .A(n100), .B(a[598]), .Z(n24621) );
  AND U25268 ( .A(n24622), .B(n24621), .Z(n24675) );
  XOR U25269 ( .A(a[595]), .B(n42197), .Z(n24664) );
  NANDN U25270 ( .A(n24664), .B(n42173), .Z(n24625) );
  NANDN U25271 ( .A(n24623), .B(n42172), .Z(n24624) );
  NAND U25272 ( .A(n24625), .B(n24624), .Z(n24673) );
  NAND U25273 ( .A(b[7]), .B(a[591]), .Z(n24674) );
  XNOR U25274 ( .A(n24673), .B(n24674), .Z(n24676) );
  XOR U25275 ( .A(n24675), .B(n24676), .Z(n24682) );
  NANDN U25276 ( .A(n24626), .B(n42093), .Z(n24628) );
  XOR U25277 ( .A(n42134), .B(a[597]), .Z(n24667) );
  NANDN U25278 ( .A(n24667), .B(n42095), .Z(n24627) );
  NAND U25279 ( .A(n24628), .B(n24627), .Z(n24680) );
  NANDN U25280 ( .A(n24629), .B(n42231), .Z(n24631) );
  XOR U25281 ( .A(n211), .B(a[593]), .Z(n24670) );
  NANDN U25282 ( .A(n24670), .B(n42234), .Z(n24630) );
  AND U25283 ( .A(n24631), .B(n24630), .Z(n24679) );
  XNOR U25284 ( .A(n24680), .B(n24679), .Z(n24681) );
  XNOR U25285 ( .A(n24682), .B(n24681), .Z(n24686) );
  NANDN U25286 ( .A(n24633), .B(n24632), .Z(n24637) );
  NAND U25287 ( .A(n24635), .B(n24634), .Z(n24636) );
  AND U25288 ( .A(n24637), .B(n24636), .Z(n24685) );
  XOR U25289 ( .A(n24686), .B(n24685), .Z(n24687) );
  NANDN U25290 ( .A(n24639), .B(n24638), .Z(n24643) );
  NANDN U25291 ( .A(n24641), .B(n24640), .Z(n24642) );
  NAND U25292 ( .A(n24643), .B(n24642), .Z(n24688) );
  XOR U25293 ( .A(n24687), .B(n24688), .Z(n24655) );
  OR U25294 ( .A(n24645), .B(n24644), .Z(n24649) );
  NANDN U25295 ( .A(n24647), .B(n24646), .Z(n24648) );
  NAND U25296 ( .A(n24649), .B(n24648), .Z(n24656) );
  XNOR U25297 ( .A(n24655), .B(n24656), .Z(n24657) );
  XNOR U25298 ( .A(n24658), .B(n24657), .Z(n24691) );
  XNOR U25299 ( .A(n24691), .B(sreg[1615]), .Z(n24693) );
  NAND U25300 ( .A(n24650), .B(sreg[1614]), .Z(n24654) );
  OR U25301 ( .A(n24652), .B(n24651), .Z(n24653) );
  AND U25302 ( .A(n24654), .B(n24653), .Z(n24692) );
  XOR U25303 ( .A(n24693), .B(n24692), .Z(c[1615]) );
  NANDN U25304 ( .A(n24656), .B(n24655), .Z(n24660) );
  NAND U25305 ( .A(n24658), .B(n24657), .Z(n24659) );
  NAND U25306 ( .A(n24660), .B(n24659), .Z(n24699) );
  NAND U25307 ( .A(b[0]), .B(a[600]), .Z(n24661) );
  XNOR U25308 ( .A(b[1]), .B(n24661), .Z(n24663) );
  NAND U25309 ( .A(n100), .B(a[599]), .Z(n24662) );
  AND U25310 ( .A(n24663), .B(n24662), .Z(n24716) );
  XOR U25311 ( .A(a[596]), .B(n42197), .Z(n24705) );
  NANDN U25312 ( .A(n24705), .B(n42173), .Z(n24666) );
  NANDN U25313 ( .A(n24664), .B(n42172), .Z(n24665) );
  NAND U25314 ( .A(n24666), .B(n24665), .Z(n24714) );
  NAND U25315 ( .A(b[7]), .B(a[592]), .Z(n24715) );
  XNOR U25316 ( .A(n24714), .B(n24715), .Z(n24717) );
  XOR U25317 ( .A(n24716), .B(n24717), .Z(n24723) );
  NANDN U25318 ( .A(n24667), .B(n42093), .Z(n24669) );
  XOR U25319 ( .A(n42134), .B(a[598]), .Z(n24708) );
  NANDN U25320 ( .A(n24708), .B(n42095), .Z(n24668) );
  NAND U25321 ( .A(n24669), .B(n24668), .Z(n24721) );
  NANDN U25322 ( .A(n24670), .B(n42231), .Z(n24672) );
  XOR U25323 ( .A(n211), .B(a[594]), .Z(n24711) );
  NANDN U25324 ( .A(n24711), .B(n42234), .Z(n24671) );
  AND U25325 ( .A(n24672), .B(n24671), .Z(n24720) );
  XNOR U25326 ( .A(n24721), .B(n24720), .Z(n24722) );
  XNOR U25327 ( .A(n24723), .B(n24722), .Z(n24727) );
  NANDN U25328 ( .A(n24674), .B(n24673), .Z(n24678) );
  NAND U25329 ( .A(n24676), .B(n24675), .Z(n24677) );
  AND U25330 ( .A(n24678), .B(n24677), .Z(n24726) );
  XOR U25331 ( .A(n24727), .B(n24726), .Z(n24728) );
  NANDN U25332 ( .A(n24680), .B(n24679), .Z(n24684) );
  NANDN U25333 ( .A(n24682), .B(n24681), .Z(n24683) );
  NAND U25334 ( .A(n24684), .B(n24683), .Z(n24729) );
  XOR U25335 ( .A(n24728), .B(n24729), .Z(n24696) );
  OR U25336 ( .A(n24686), .B(n24685), .Z(n24690) );
  NANDN U25337 ( .A(n24688), .B(n24687), .Z(n24689) );
  NAND U25338 ( .A(n24690), .B(n24689), .Z(n24697) );
  XNOR U25339 ( .A(n24696), .B(n24697), .Z(n24698) );
  XNOR U25340 ( .A(n24699), .B(n24698), .Z(n24732) );
  XNOR U25341 ( .A(n24732), .B(sreg[1616]), .Z(n24734) );
  NAND U25342 ( .A(n24691), .B(sreg[1615]), .Z(n24695) );
  OR U25343 ( .A(n24693), .B(n24692), .Z(n24694) );
  AND U25344 ( .A(n24695), .B(n24694), .Z(n24733) );
  XOR U25345 ( .A(n24734), .B(n24733), .Z(c[1616]) );
  NANDN U25346 ( .A(n24697), .B(n24696), .Z(n24701) );
  NAND U25347 ( .A(n24699), .B(n24698), .Z(n24700) );
  NAND U25348 ( .A(n24701), .B(n24700), .Z(n24740) );
  NAND U25349 ( .A(b[0]), .B(a[601]), .Z(n24702) );
  XNOR U25350 ( .A(b[1]), .B(n24702), .Z(n24704) );
  NAND U25351 ( .A(n100), .B(a[600]), .Z(n24703) );
  AND U25352 ( .A(n24704), .B(n24703), .Z(n24757) );
  XOR U25353 ( .A(a[597]), .B(n42197), .Z(n24746) );
  NANDN U25354 ( .A(n24746), .B(n42173), .Z(n24707) );
  NANDN U25355 ( .A(n24705), .B(n42172), .Z(n24706) );
  NAND U25356 ( .A(n24707), .B(n24706), .Z(n24755) );
  NAND U25357 ( .A(b[7]), .B(a[593]), .Z(n24756) );
  XNOR U25358 ( .A(n24755), .B(n24756), .Z(n24758) );
  XOR U25359 ( .A(n24757), .B(n24758), .Z(n24764) );
  NANDN U25360 ( .A(n24708), .B(n42093), .Z(n24710) );
  XOR U25361 ( .A(n42134), .B(a[599]), .Z(n24749) );
  NANDN U25362 ( .A(n24749), .B(n42095), .Z(n24709) );
  NAND U25363 ( .A(n24710), .B(n24709), .Z(n24762) );
  NANDN U25364 ( .A(n24711), .B(n42231), .Z(n24713) );
  XOR U25365 ( .A(n211), .B(a[595]), .Z(n24752) );
  NANDN U25366 ( .A(n24752), .B(n42234), .Z(n24712) );
  AND U25367 ( .A(n24713), .B(n24712), .Z(n24761) );
  XNOR U25368 ( .A(n24762), .B(n24761), .Z(n24763) );
  XNOR U25369 ( .A(n24764), .B(n24763), .Z(n24768) );
  NANDN U25370 ( .A(n24715), .B(n24714), .Z(n24719) );
  NAND U25371 ( .A(n24717), .B(n24716), .Z(n24718) );
  AND U25372 ( .A(n24719), .B(n24718), .Z(n24767) );
  XOR U25373 ( .A(n24768), .B(n24767), .Z(n24769) );
  NANDN U25374 ( .A(n24721), .B(n24720), .Z(n24725) );
  NANDN U25375 ( .A(n24723), .B(n24722), .Z(n24724) );
  NAND U25376 ( .A(n24725), .B(n24724), .Z(n24770) );
  XOR U25377 ( .A(n24769), .B(n24770), .Z(n24737) );
  OR U25378 ( .A(n24727), .B(n24726), .Z(n24731) );
  NANDN U25379 ( .A(n24729), .B(n24728), .Z(n24730) );
  NAND U25380 ( .A(n24731), .B(n24730), .Z(n24738) );
  XNOR U25381 ( .A(n24737), .B(n24738), .Z(n24739) );
  XNOR U25382 ( .A(n24740), .B(n24739), .Z(n24773) );
  XNOR U25383 ( .A(n24773), .B(sreg[1617]), .Z(n24775) );
  NAND U25384 ( .A(n24732), .B(sreg[1616]), .Z(n24736) );
  OR U25385 ( .A(n24734), .B(n24733), .Z(n24735) );
  AND U25386 ( .A(n24736), .B(n24735), .Z(n24774) );
  XOR U25387 ( .A(n24775), .B(n24774), .Z(c[1617]) );
  NANDN U25388 ( .A(n24738), .B(n24737), .Z(n24742) );
  NAND U25389 ( .A(n24740), .B(n24739), .Z(n24741) );
  NAND U25390 ( .A(n24742), .B(n24741), .Z(n24781) );
  NAND U25391 ( .A(b[0]), .B(a[602]), .Z(n24743) );
  XNOR U25392 ( .A(b[1]), .B(n24743), .Z(n24745) );
  NAND U25393 ( .A(n101), .B(a[601]), .Z(n24744) );
  AND U25394 ( .A(n24745), .B(n24744), .Z(n24798) );
  XOR U25395 ( .A(a[598]), .B(n42197), .Z(n24787) );
  NANDN U25396 ( .A(n24787), .B(n42173), .Z(n24748) );
  NANDN U25397 ( .A(n24746), .B(n42172), .Z(n24747) );
  NAND U25398 ( .A(n24748), .B(n24747), .Z(n24796) );
  NAND U25399 ( .A(b[7]), .B(a[594]), .Z(n24797) );
  XNOR U25400 ( .A(n24796), .B(n24797), .Z(n24799) );
  XOR U25401 ( .A(n24798), .B(n24799), .Z(n24805) );
  NANDN U25402 ( .A(n24749), .B(n42093), .Z(n24751) );
  XOR U25403 ( .A(n42134), .B(a[600]), .Z(n24790) );
  NANDN U25404 ( .A(n24790), .B(n42095), .Z(n24750) );
  NAND U25405 ( .A(n24751), .B(n24750), .Z(n24803) );
  NANDN U25406 ( .A(n24752), .B(n42231), .Z(n24754) );
  XOR U25407 ( .A(n211), .B(a[596]), .Z(n24793) );
  NANDN U25408 ( .A(n24793), .B(n42234), .Z(n24753) );
  AND U25409 ( .A(n24754), .B(n24753), .Z(n24802) );
  XNOR U25410 ( .A(n24803), .B(n24802), .Z(n24804) );
  XNOR U25411 ( .A(n24805), .B(n24804), .Z(n24809) );
  NANDN U25412 ( .A(n24756), .B(n24755), .Z(n24760) );
  NAND U25413 ( .A(n24758), .B(n24757), .Z(n24759) );
  AND U25414 ( .A(n24760), .B(n24759), .Z(n24808) );
  XOR U25415 ( .A(n24809), .B(n24808), .Z(n24810) );
  NANDN U25416 ( .A(n24762), .B(n24761), .Z(n24766) );
  NANDN U25417 ( .A(n24764), .B(n24763), .Z(n24765) );
  NAND U25418 ( .A(n24766), .B(n24765), .Z(n24811) );
  XOR U25419 ( .A(n24810), .B(n24811), .Z(n24778) );
  OR U25420 ( .A(n24768), .B(n24767), .Z(n24772) );
  NANDN U25421 ( .A(n24770), .B(n24769), .Z(n24771) );
  NAND U25422 ( .A(n24772), .B(n24771), .Z(n24779) );
  XNOR U25423 ( .A(n24778), .B(n24779), .Z(n24780) );
  XNOR U25424 ( .A(n24781), .B(n24780), .Z(n24814) );
  XNOR U25425 ( .A(n24814), .B(sreg[1618]), .Z(n24816) );
  NAND U25426 ( .A(n24773), .B(sreg[1617]), .Z(n24777) );
  OR U25427 ( .A(n24775), .B(n24774), .Z(n24776) );
  AND U25428 ( .A(n24777), .B(n24776), .Z(n24815) );
  XOR U25429 ( .A(n24816), .B(n24815), .Z(c[1618]) );
  NANDN U25430 ( .A(n24779), .B(n24778), .Z(n24783) );
  NAND U25431 ( .A(n24781), .B(n24780), .Z(n24782) );
  NAND U25432 ( .A(n24783), .B(n24782), .Z(n24822) );
  NAND U25433 ( .A(b[0]), .B(a[603]), .Z(n24784) );
  XNOR U25434 ( .A(b[1]), .B(n24784), .Z(n24786) );
  NAND U25435 ( .A(n101), .B(a[602]), .Z(n24785) );
  AND U25436 ( .A(n24786), .B(n24785), .Z(n24839) );
  XOR U25437 ( .A(a[599]), .B(n42197), .Z(n24828) );
  NANDN U25438 ( .A(n24828), .B(n42173), .Z(n24789) );
  NANDN U25439 ( .A(n24787), .B(n42172), .Z(n24788) );
  NAND U25440 ( .A(n24789), .B(n24788), .Z(n24837) );
  NAND U25441 ( .A(b[7]), .B(a[595]), .Z(n24838) );
  XNOR U25442 ( .A(n24837), .B(n24838), .Z(n24840) );
  XOR U25443 ( .A(n24839), .B(n24840), .Z(n24846) );
  NANDN U25444 ( .A(n24790), .B(n42093), .Z(n24792) );
  XOR U25445 ( .A(n42134), .B(a[601]), .Z(n24831) );
  NANDN U25446 ( .A(n24831), .B(n42095), .Z(n24791) );
  NAND U25447 ( .A(n24792), .B(n24791), .Z(n24844) );
  NANDN U25448 ( .A(n24793), .B(n42231), .Z(n24795) );
  XOR U25449 ( .A(n211), .B(a[597]), .Z(n24834) );
  NANDN U25450 ( .A(n24834), .B(n42234), .Z(n24794) );
  AND U25451 ( .A(n24795), .B(n24794), .Z(n24843) );
  XNOR U25452 ( .A(n24844), .B(n24843), .Z(n24845) );
  XNOR U25453 ( .A(n24846), .B(n24845), .Z(n24850) );
  NANDN U25454 ( .A(n24797), .B(n24796), .Z(n24801) );
  NAND U25455 ( .A(n24799), .B(n24798), .Z(n24800) );
  AND U25456 ( .A(n24801), .B(n24800), .Z(n24849) );
  XOR U25457 ( .A(n24850), .B(n24849), .Z(n24851) );
  NANDN U25458 ( .A(n24803), .B(n24802), .Z(n24807) );
  NANDN U25459 ( .A(n24805), .B(n24804), .Z(n24806) );
  NAND U25460 ( .A(n24807), .B(n24806), .Z(n24852) );
  XOR U25461 ( .A(n24851), .B(n24852), .Z(n24819) );
  OR U25462 ( .A(n24809), .B(n24808), .Z(n24813) );
  NANDN U25463 ( .A(n24811), .B(n24810), .Z(n24812) );
  NAND U25464 ( .A(n24813), .B(n24812), .Z(n24820) );
  XNOR U25465 ( .A(n24819), .B(n24820), .Z(n24821) );
  XNOR U25466 ( .A(n24822), .B(n24821), .Z(n24855) );
  XNOR U25467 ( .A(n24855), .B(sreg[1619]), .Z(n24857) );
  NAND U25468 ( .A(n24814), .B(sreg[1618]), .Z(n24818) );
  OR U25469 ( .A(n24816), .B(n24815), .Z(n24817) );
  AND U25470 ( .A(n24818), .B(n24817), .Z(n24856) );
  XOR U25471 ( .A(n24857), .B(n24856), .Z(c[1619]) );
  NANDN U25472 ( .A(n24820), .B(n24819), .Z(n24824) );
  NAND U25473 ( .A(n24822), .B(n24821), .Z(n24823) );
  NAND U25474 ( .A(n24824), .B(n24823), .Z(n24863) );
  NAND U25475 ( .A(b[0]), .B(a[604]), .Z(n24825) );
  XNOR U25476 ( .A(b[1]), .B(n24825), .Z(n24827) );
  NAND U25477 ( .A(n101), .B(a[603]), .Z(n24826) );
  AND U25478 ( .A(n24827), .B(n24826), .Z(n24880) );
  XOR U25479 ( .A(a[600]), .B(n42197), .Z(n24869) );
  NANDN U25480 ( .A(n24869), .B(n42173), .Z(n24830) );
  NANDN U25481 ( .A(n24828), .B(n42172), .Z(n24829) );
  NAND U25482 ( .A(n24830), .B(n24829), .Z(n24878) );
  NAND U25483 ( .A(b[7]), .B(a[596]), .Z(n24879) );
  XNOR U25484 ( .A(n24878), .B(n24879), .Z(n24881) );
  XOR U25485 ( .A(n24880), .B(n24881), .Z(n24887) );
  NANDN U25486 ( .A(n24831), .B(n42093), .Z(n24833) );
  XOR U25487 ( .A(n42134), .B(a[602]), .Z(n24872) );
  NANDN U25488 ( .A(n24872), .B(n42095), .Z(n24832) );
  NAND U25489 ( .A(n24833), .B(n24832), .Z(n24885) );
  NANDN U25490 ( .A(n24834), .B(n42231), .Z(n24836) );
  XOR U25491 ( .A(n211), .B(a[598]), .Z(n24875) );
  NANDN U25492 ( .A(n24875), .B(n42234), .Z(n24835) );
  AND U25493 ( .A(n24836), .B(n24835), .Z(n24884) );
  XNOR U25494 ( .A(n24885), .B(n24884), .Z(n24886) );
  XNOR U25495 ( .A(n24887), .B(n24886), .Z(n24891) );
  NANDN U25496 ( .A(n24838), .B(n24837), .Z(n24842) );
  NAND U25497 ( .A(n24840), .B(n24839), .Z(n24841) );
  AND U25498 ( .A(n24842), .B(n24841), .Z(n24890) );
  XOR U25499 ( .A(n24891), .B(n24890), .Z(n24892) );
  NANDN U25500 ( .A(n24844), .B(n24843), .Z(n24848) );
  NANDN U25501 ( .A(n24846), .B(n24845), .Z(n24847) );
  NAND U25502 ( .A(n24848), .B(n24847), .Z(n24893) );
  XOR U25503 ( .A(n24892), .B(n24893), .Z(n24860) );
  OR U25504 ( .A(n24850), .B(n24849), .Z(n24854) );
  NANDN U25505 ( .A(n24852), .B(n24851), .Z(n24853) );
  NAND U25506 ( .A(n24854), .B(n24853), .Z(n24861) );
  XNOR U25507 ( .A(n24860), .B(n24861), .Z(n24862) );
  XNOR U25508 ( .A(n24863), .B(n24862), .Z(n24896) );
  XNOR U25509 ( .A(n24896), .B(sreg[1620]), .Z(n24898) );
  NAND U25510 ( .A(n24855), .B(sreg[1619]), .Z(n24859) );
  OR U25511 ( .A(n24857), .B(n24856), .Z(n24858) );
  AND U25512 ( .A(n24859), .B(n24858), .Z(n24897) );
  XOR U25513 ( .A(n24898), .B(n24897), .Z(c[1620]) );
  NANDN U25514 ( .A(n24861), .B(n24860), .Z(n24865) );
  NAND U25515 ( .A(n24863), .B(n24862), .Z(n24864) );
  NAND U25516 ( .A(n24865), .B(n24864), .Z(n24904) );
  NAND U25517 ( .A(b[0]), .B(a[605]), .Z(n24866) );
  XNOR U25518 ( .A(b[1]), .B(n24866), .Z(n24868) );
  NAND U25519 ( .A(n101), .B(a[604]), .Z(n24867) );
  AND U25520 ( .A(n24868), .B(n24867), .Z(n24921) );
  XOR U25521 ( .A(a[601]), .B(n42197), .Z(n24910) );
  NANDN U25522 ( .A(n24910), .B(n42173), .Z(n24871) );
  NANDN U25523 ( .A(n24869), .B(n42172), .Z(n24870) );
  NAND U25524 ( .A(n24871), .B(n24870), .Z(n24919) );
  NAND U25525 ( .A(b[7]), .B(a[597]), .Z(n24920) );
  XNOR U25526 ( .A(n24919), .B(n24920), .Z(n24922) );
  XOR U25527 ( .A(n24921), .B(n24922), .Z(n24928) );
  NANDN U25528 ( .A(n24872), .B(n42093), .Z(n24874) );
  XOR U25529 ( .A(n42134), .B(a[603]), .Z(n24913) );
  NANDN U25530 ( .A(n24913), .B(n42095), .Z(n24873) );
  NAND U25531 ( .A(n24874), .B(n24873), .Z(n24926) );
  NANDN U25532 ( .A(n24875), .B(n42231), .Z(n24877) );
  XOR U25533 ( .A(n212), .B(a[599]), .Z(n24916) );
  NANDN U25534 ( .A(n24916), .B(n42234), .Z(n24876) );
  AND U25535 ( .A(n24877), .B(n24876), .Z(n24925) );
  XNOR U25536 ( .A(n24926), .B(n24925), .Z(n24927) );
  XNOR U25537 ( .A(n24928), .B(n24927), .Z(n24932) );
  NANDN U25538 ( .A(n24879), .B(n24878), .Z(n24883) );
  NAND U25539 ( .A(n24881), .B(n24880), .Z(n24882) );
  AND U25540 ( .A(n24883), .B(n24882), .Z(n24931) );
  XOR U25541 ( .A(n24932), .B(n24931), .Z(n24933) );
  NANDN U25542 ( .A(n24885), .B(n24884), .Z(n24889) );
  NANDN U25543 ( .A(n24887), .B(n24886), .Z(n24888) );
  NAND U25544 ( .A(n24889), .B(n24888), .Z(n24934) );
  XOR U25545 ( .A(n24933), .B(n24934), .Z(n24901) );
  OR U25546 ( .A(n24891), .B(n24890), .Z(n24895) );
  NANDN U25547 ( .A(n24893), .B(n24892), .Z(n24894) );
  NAND U25548 ( .A(n24895), .B(n24894), .Z(n24902) );
  XNOR U25549 ( .A(n24901), .B(n24902), .Z(n24903) );
  XNOR U25550 ( .A(n24904), .B(n24903), .Z(n24937) );
  XNOR U25551 ( .A(n24937), .B(sreg[1621]), .Z(n24939) );
  NAND U25552 ( .A(n24896), .B(sreg[1620]), .Z(n24900) );
  OR U25553 ( .A(n24898), .B(n24897), .Z(n24899) );
  AND U25554 ( .A(n24900), .B(n24899), .Z(n24938) );
  XOR U25555 ( .A(n24939), .B(n24938), .Z(c[1621]) );
  NANDN U25556 ( .A(n24902), .B(n24901), .Z(n24906) );
  NAND U25557 ( .A(n24904), .B(n24903), .Z(n24905) );
  NAND U25558 ( .A(n24906), .B(n24905), .Z(n24945) );
  NAND U25559 ( .A(b[0]), .B(a[606]), .Z(n24907) );
  XNOR U25560 ( .A(b[1]), .B(n24907), .Z(n24909) );
  NAND U25561 ( .A(n101), .B(a[605]), .Z(n24908) );
  AND U25562 ( .A(n24909), .B(n24908), .Z(n24962) );
  XOR U25563 ( .A(a[602]), .B(n42197), .Z(n24951) );
  NANDN U25564 ( .A(n24951), .B(n42173), .Z(n24912) );
  NANDN U25565 ( .A(n24910), .B(n42172), .Z(n24911) );
  NAND U25566 ( .A(n24912), .B(n24911), .Z(n24960) );
  NAND U25567 ( .A(b[7]), .B(a[598]), .Z(n24961) );
  XNOR U25568 ( .A(n24960), .B(n24961), .Z(n24963) );
  XOR U25569 ( .A(n24962), .B(n24963), .Z(n24969) );
  NANDN U25570 ( .A(n24913), .B(n42093), .Z(n24915) );
  XOR U25571 ( .A(n42134), .B(a[604]), .Z(n24954) );
  NANDN U25572 ( .A(n24954), .B(n42095), .Z(n24914) );
  NAND U25573 ( .A(n24915), .B(n24914), .Z(n24967) );
  NANDN U25574 ( .A(n24916), .B(n42231), .Z(n24918) );
  XOR U25575 ( .A(n212), .B(a[600]), .Z(n24957) );
  NANDN U25576 ( .A(n24957), .B(n42234), .Z(n24917) );
  AND U25577 ( .A(n24918), .B(n24917), .Z(n24966) );
  XNOR U25578 ( .A(n24967), .B(n24966), .Z(n24968) );
  XNOR U25579 ( .A(n24969), .B(n24968), .Z(n24973) );
  NANDN U25580 ( .A(n24920), .B(n24919), .Z(n24924) );
  NAND U25581 ( .A(n24922), .B(n24921), .Z(n24923) );
  AND U25582 ( .A(n24924), .B(n24923), .Z(n24972) );
  XOR U25583 ( .A(n24973), .B(n24972), .Z(n24974) );
  NANDN U25584 ( .A(n24926), .B(n24925), .Z(n24930) );
  NANDN U25585 ( .A(n24928), .B(n24927), .Z(n24929) );
  NAND U25586 ( .A(n24930), .B(n24929), .Z(n24975) );
  XOR U25587 ( .A(n24974), .B(n24975), .Z(n24942) );
  OR U25588 ( .A(n24932), .B(n24931), .Z(n24936) );
  NANDN U25589 ( .A(n24934), .B(n24933), .Z(n24935) );
  NAND U25590 ( .A(n24936), .B(n24935), .Z(n24943) );
  XNOR U25591 ( .A(n24942), .B(n24943), .Z(n24944) );
  XNOR U25592 ( .A(n24945), .B(n24944), .Z(n24978) );
  XNOR U25593 ( .A(n24978), .B(sreg[1622]), .Z(n24980) );
  NAND U25594 ( .A(n24937), .B(sreg[1621]), .Z(n24941) );
  OR U25595 ( .A(n24939), .B(n24938), .Z(n24940) );
  AND U25596 ( .A(n24941), .B(n24940), .Z(n24979) );
  XOR U25597 ( .A(n24980), .B(n24979), .Z(c[1622]) );
  NANDN U25598 ( .A(n24943), .B(n24942), .Z(n24947) );
  NAND U25599 ( .A(n24945), .B(n24944), .Z(n24946) );
  NAND U25600 ( .A(n24947), .B(n24946), .Z(n24986) );
  NAND U25601 ( .A(b[0]), .B(a[607]), .Z(n24948) );
  XNOR U25602 ( .A(b[1]), .B(n24948), .Z(n24950) );
  NAND U25603 ( .A(n101), .B(a[606]), .Z(n24949) );
  AND U25604 ( .A(n24950), .B(n24949), .Z(n25003) );
  XOR U25605 ( .A(a[603]), .B(n42197), .Z(n24992) );
  NANDN U25606 ( .A(n24992), .B(n42173), .Z(n24953) );
  NANDN U25607 ( .A(n24951), .B(n42172), .Z(n24952) );
  NAND U25608 ( .A(n24953), .B(n24952), .Z(n25001) );
  NAND U25609 ( .A(b[7]), .B(a[599]), .Z(n25002) );
  XNOR U25610 ( .A(n25001), .B(n25002), .Z(n25004) );
  XOR U25611 ( .A(n25003), .B(n25004), .Z(n25010) );
  NANDN U25612 ( .A(n24954), .B(n42093), .Z(n24956) );
  XOR U25613 ( .A(n42134), .B(a[605]), .Z(n24995) );
  NANDN U25614 ( .A(n24995), .B(n42095), .Z(n24955) );
  NAND U25615 ( .A(n24956), .B(n24955), .Z(n25008) );
  NANDN U25616 ( .A(n24957), .B(n42231), .Z(n24959) );
  XOR U25617 ( .A(n212), .B(a[601]), .Z(n24998) );
  NANDN U25618 ( .A(n24998), .B(n42234), .Z(n24958) );
  AND U25619 ( .A(n24959), .B(n24958), .Z(n25007) );
  XNOR U25620 ( .A(n25008), .B(n25007), .Z(n25009) );
  XNOR U25621 ( .A(n25010), .B(n25009), .Z(n25014) );
  NANDN U25622 ( .A(n24961), .B(n24960), .Z(n24965) );
  NAND U25623 ( .A(n24963), .B(n24962), .Z(n24964) );
  AND U25624 ( .A(n24965), .B(n24964), .Z(n25013) );
  XOR U25625 ( .A(n25014), .B(n25013), .Z(n25015) );
  NANDN U25626 ( .A(n24967), .B(n24966), .Z(n24971) );
  NANDN U25627 ( .A(n24969), .B(n24968), .Z(n24970) );
  NAND U25628 ( .A(n24971), .B(n24970), .Z(n25016) );
  XOR U25629 ( .A(n25015), .B(n25016), .Z(n24983) );
  OR U25630 ( .A(n24973), .B(n24972), .Z(n24977) );
  NANDN U25631 ( .A(n24975), .B(n24974), .Z(n24976) );
  NAND U25632 ( .A(n24977), .B(n24976), .Z(n24984) );
  XNOR U25633 ( .A(n24983), .B(n24984), .Z(n24985) );
  XNOR U25634 ( .A(n24986), .B(n24985), .Z(n25019) );
  XNOR U25635 ( .A(n25019), .B(sreg[1623]), .Z(n25021) );
  NAND U25636 ( .A(n24978), .B(sreg[1622]), .Z(n24982) );
  OR U25637 ( .A(n24980), .B(n24979), .Z(n24981) );
  AND U25638 ( .A(n24982), .B(n24981), .Z(n25020) );
  XOR U25639 ( .A(n25021), .B(n25020), .Z(c[1623]) );
  NANDN U25640 ( .A(n24984), .B(n24983), .Z(n24988) );
  NAND U25641 ( .A(n24986), .B(n24985), .Z(n24987) );
  NAND U25642 ( .A(n24988), .B(n24987), .Z(n25027) );
  NAND U25643 ( .A(b[0]), .B(a[608]), .Z(n24989) );
  XNOR U25644 ( .A(b[1]), .B(n24989), .Z(n24991) );
  NAND U25645 ( .A(n101), .B(a[607]), .Z(n24990) );
  AND U25646 ( .A(n24991), .B(n24990), .Z(n25044) );
  XOR U25647 ( .A(a[604]), .B(n42197), .Z(n25033) );
  NANDN U25648 ( .A(n25033), .B(n42173), .Z(n24994) );
  NANDN U25649 ( .A(n24992), .B(n42172), .Z(n24993) );
  NAND U25650 ( .A(n24994), .B(n24993), .Z(n25042) );
  NAND U25651 ( .A(b[7]), .B(a[600]), .Z(n25043) );
  XNOR U25652 ( .A(n25042), .B(n25043), .Z(n25045) );
  XOR U25653 ( .A(n25044), .B(n25045), .Z(n25051) );
  NANDN U25654 ( .A(n24995), .B(n42093), .Z(n24997) );
  XOR U25655 ( .A(n42134), .B(a[606]), .Z(n25036) );
  NANDN U25656 ( .A(n25036), .B(n42095), .Z(n24996) );
  NAND U25657 ( .A(n24997), .B(n24996), .Z(n25049) );
  NANDN U25658 ( .A(n24998), .B(n42231), .Z(n25000) );
  XOR U25659 ( .A(n212), .B(a[602]), .Z(n25039) );
  NANDN U25660 ( .A(n25039), .B(n42234), .Z(n24999) );
  AND U25661 ( .A(n25000), .B(n24999), .Z(n25048) );
  XNOR U25662 ( .A(n25049), .B(n25048), .Z(n25050) );
  XNOR U25663 ( .A(n25051), .B(n25050), .Z(n25055) );
  NANDN U25664 ( .A(n25002), .B(n25001), .Z(n25006) );
  NAND U25665 ( .A(n25004), .B(n25003), .Z(n25005) );
  AND U25666 ( .A(n25006), .B(n25005), .Z(n25054) );
  XOR U25667 ( .A(n25055), .B(n25054), .Z(n25056) );
  NANDN U25668 ( .A(n25008), .B(n25007), .Z(n25012) );
  NANDN U25669 ( .A(n25010), .B(n25009), .Z(n25011) );
  NAND U25670 ( .A(n25012), .B(n25011), .Z(n25057) );
  XOR U25671 ( .A(n25056), .B(n25057), .Z(n25024) );
  OR U25672 ( .A(n25014), .B(n25013), .Z(n25018) );
  NANDN U25673 ( .A(n25016), .B(n25015), .Z(n25017) );
  NAND U25674 ( .A(n25018), .B(n25017), .Z(n25025) );
  XNOR U25675 ( .A(n25024), .B(n25025), .Z(n25026) );
  XNOR U25676 ( .A(n25027), .B(n25026), .Z(n25060) );
  XNOR U25677 ( .A(n25060), .B(sreg[1624]), .Z(n25062) );
  NAND U25678 ( .A(n25019), .B(sreg[1623]), .Z(n25023) );
  OR U25679 ( .A(n25021), .B(n25020), .Z(n25022) );
  AND U25680 ( .A(n25023), .B(n25022), .Z(n25061) );
  XOR U25681 ( .A(n25062), .B(n25061), .Z(c[1624]) );
  NANDN U25682 ( .A(n25025), .B(n25024), .Z(n25029) );
  NAND U25683 ( .A(n25027), .B(n25026), .Z(n25028) );
  NAND U25684 ( .A(n25029), .B(n25028), .Z(n25068) );
  NAND U25685 ( .A(b[0]), .B(a[609]), .Z(n25030) );
  XNOR U25686 ( .A(b[1]), .B(n25030), .Z(n25032) );
  NAND U25687 ( .A(n102), .B(a[608]), .Z(n25031) );
  AND U25688 ( .A(n25032), .B(n25031), .Z(n25085) );
  XOR U25689 ( .A(a[605]), .B(n42197), .Z(n25074) );
  NANDN U25690 ( .A(n25074), .B(n42173), .Z(n25035) );
  NANDN U25691 ( .A(n25033), .B(n42172), .Z(n25034) );
  NAND U25692 ( .A(n25035), .B(n25034), .Z(n25083) );
  NAND U25693 ( .A(b[7]), .B(a[601]), .Z(n25084) );
  XNOR U25694 ( .A(n25083), .B(n25084), .Z(n25086) );
  XOR U25695 ( .A(n25085), .B(n25086), .Z(n25092) );
  NANDN U25696 ( .A(n25036), .B(n42093), .Z(n25038) );
  XOR U25697 ( .A(n42134), .B(a[607]), .Z(n25077) );
  NANDN U25698 ( .A(n25077), .B(n42095), .Z(n25037) );
  NAND U25699 ( .A(n25038), .B(n25037), .Z(n25090) );
  NANDN U25700 ( .A(n25039), .B(n42231), .Z(n25041) );
  XOR U25701 ( .A(n212), .B(a[603]), .Z(n25080) );
  NANDN U25702 ( .A(n25080), .B(n42234), .Z(n25040) );
  AND U25703 ( .A(n25041), .B(n25040), .Z(n25089) );
  XNOR U25704 ( .A(n25090), .B(n25089), .Z(n25091) );
  XNOR U25705 ( .A(n25092), .B(n25091), .Z(n25096) );
  NANDN U25706 ( .A(n25043), .B(n25042), .Z(n25047) );
  NAND U25707 ( .A(n25045), .B(n25044), .Z(n25046) );
  AND U25708 ( .A(n25047), .B(n25046), .Z(n25095) );
  XOR U25709 ( .A(n25096), .B(n25095), .Z(n25097) );
  NANDN U25710 ( .A(n25049), .B(n25048), .Z(n25053) );
  NANDN U25711 ( .A(n25051), .B(n25050), .Z(n25052) );
  NAND U25712 ( .A(n25053), .B(n25052), .Z(n25098) );
  XOR U25713 ( .A(n25097), .B(n25098), .Z(n25065) );
  OR U25714 ( .A(n25055), .B(n25054), .Z(n25059) );
  NANDN U25715 ( .A(n25057), .B(n25056), .Z(n25058) );
  NAND U25716 ( .A(n25059), .B(n25058), .Z(n25066) );
  XNOR U25717 ( .A(n25065), .B(n25066), .Z(n25067) );
  XNOR U25718 ( .A(n25068), .B(n25067), .Z(n25101) );
  XNOR U25719 ( .A(n25101), .B(sreg[1625]), .Z(n25103) );
  NAND U25720 ( .A(n25060), .B(sreg[1624]), .Z(n25064) );
  OR U25721 ( .A(n25062), .B(n25061), .Z(n25063) );
  AND U25722 ( .A(n25064), .B(n25063), .Z(n25102) );
  XOR U25723 ( .A(n25103), .B(n25102), .Z(c[1625]) );
  NANDN U25724 ( .A(n25066), .B(n25065), .Z(n25070) );
  NAND U25725 ( .A(n25068), .B(n25067), .Z(n25069) );
  NAND U25726 ( .A(n25070), .B(n25069), .Z(n25109) );
  NAND U25727 ( .A(b[0]), .B(a[610]), .Z(n25071) );
  XNOR U25728 ( .A(b[1]), .B(n25071), .Z(n25073) );
  NAND U25729 ( .A(n102), .B(a[609]), .Z(n25072) );
  AND U25730 ( .A(n25073), .B(n25072), .Z(n25126) );
  XOR U25731 ( .A(a[606]), .B(n42197), .Z(n25115) );
  NANDN U25732 ( .A(n25115), .B(n42173), .Z(n25076) );
  NANDN U25733 ( .A(n25074), .B(n42172), .Z(n25075) );
  NAND U25734 ( .A(n25076), .B(n25075), .Z(n25124) );
  NAND U25735 ( .A(b[7]), .B(a[602]), .Z(n25125) );
  XNOR U25736 ( .A(n25124), .B(n25125), .Z(n25127) );
  XOR U25737 ( .A(n25126), .B(n25127), .Z(n25133) );
  NANDN U25738 ( .A(n25077), .B(n42093), .Z(n25079) );
  XOR U25739 ( .A(n42134), .B(a[608]), .Z(n25118) );
  NANDN U25740 ( .A(n25118), .B(n42095), .Z(n25078) );
  NAND U25741 ( .A(n25079), .B(n25078), .Z(n25131) );
  NANDN U25742 ( .A(n25080), .B(n42231), .Z(n25082) );
  XOR U25743 ( .A(n212), .B(a[604]), .Z(n25121) );
  NANDN U25744 ( .A(n25121), .B(n42234), .Z(n25081) );
  AND U25745 ( .A(n25082), .B(n25081), .Z(n25130) );
  XNOR U25746 ( .A(n25131), .B(n25130), .Z(n25132) );
  XNOR U25747 ( .A(n25133), .B(n25132), .Z(n25137) );
  NANDN U25748 ( .A(n25084), .B(n25083), .Z(n25088) );
  NAND U25749 ( .A(n25086), .B(n25085), .Z(n25087) );
  AND U25750 ( .A(n25088), .B(n25087), .Z(n25136) );
  XOR U25751 ( .A(n25137), .B(n25136), .Z(n25138) );
  NANDN U25752 ( .A(n25090), .B(n25089), .Z(n25094) );
  NANDN U25753 ( .A(n25092), .B(n25091), .Z(n25093) );
  NAND U25754 ( .A(n25094), .B(n25093), .Z(n25139) );
  XOR U25755 ( .A(n25138), .B(n25139), .Z(n25106) );
  OR U25756 ( .A(n25096), .B(n25095), .Z(n25100) );
  NANDN U25757 ( .A(n25098), .B(n25097), .Z(n25099) );
  NAND U25758 ( .A(n25100), .B(n25099), .Z(n25107) );
  XNOR U25759 ( .A(n25106), .B(n25107), .Z(n25108) );
  XNOR U25760 ( .A(n25109), .B(n25108), .Z(n25142) );
  XNOR U25761 ( .A(n25142), .B(sreg[1626]), .Z(n25144) );
  NAND U25762 ( .A(n25101), .B(sreg[1625]), .Z(n25105) );
  OR U25763 ( .A(n25103), .B(n25102), .Z(n25104) );
  AND U25764 ( .A(n25105), .B(n25104), .Z(n25143) );
  XOR U25765 ( .A(n25144), .B(n25143), .Z(c[1626]) );
  NANDN U25766 ( .A(n25107), .B(n25106), .Z(n25111) );
  NAND U25767 ( .A(n25109), .B(n25108), .Z(n25110) );
  NAND U25768 ( .A(n25111), .B(n25110), .Z(n25150) );
  NAND U25769 ( .A(b[0]), .B(a[611]), .Z(n25112) );
  XNOR U25770 ( .A(b[1]), .B(n25112), .Z(n25114) );
  NAND U25771 ( .A(n102), .B(a[610]), .Z(n25113) );
  AND U25772 ( .A(n25114), .B(n25113), .Z(n25167) );
  XOR U25773 ( .A(a[607]), .B(n42197), .Z(n25156) );
  NANDN U25774 ( .A(n25156), .B(n42173), .Z(n25117) );
  NANDN U25775 ( .A(n25115), .B(n42172), .Z(n25116) );
  NAND U25776 ( .A(n25117), .B(n25116), .Z(n25165) );
  NAND U25777 ( .A(b[7]), .B(a[603]), .Z(n25166) );
  XNOR U25778 ( .A(n25165), .B(n25166), .Z(n25168) );
  XOR U25779 ( .A(n25167), .B(n25168), .Z(n25174) );
  NANDN U25780 ( .A(n25118), .B(n42093), .Z(n25120) );
  XOR U25781 ( .A(n42134), .B(a[609]), .Z(n25159) );
  NANDN U25782 ( .A(n25159), .B(n42095), .Z(n25119) );
  NAND U25783 ( .A(n25120), .B(n25119), .Z(n25172) );
  NANDN U25784 ( .A(n25121), .B(n42231), .Z(n25123) );
  XOR U25785 ( .A(n212), .B(a[605]), .Z(n25162) );
  NANDN U25786 ( .A(n25162), .B(n42234), .Z(n25122) );
  AND U25787 ( .A(n25123), .B(n25122), .Z(n25171) );
  XNOR U25788 ( .A(n25172), .B(n25171), .Z(n25173) );
  XNOR U25789 ( .A(n25174), .B(n25173), .Z(n25178) );
  NANDN U25790 ( .A(n25125), .B(n25124), .Z(n25129) );
  NAND U25791 ( .A(n25127), .B(n25126), .Z(n25128) );
  AND U25792 ( .A(n25129), .B(n25128), .Z(n25177) );
  XOR U25793 ( .A(n25178), .B(n25177), .Z(n25179) );
  NANDN U25794 ( .A(n25131), .B(n25130), .Z(n25135) );
  NANDN U25795 ( .A(n25133), .B(n25132), .Z(n25134) );
  NAND U25796 ( .A(n25135), .B(n25134), .Z(n25180) );
  XOR U25797 ( .A(n25179), .B(n25180), .Z(n25147) );
  OR U25798 ( .A(n25137), .B(n25136), .Z(n25141) );
  NANDN U25799 ( .A(n25139), .B(n25138), .Z(n25140) );
  NAND U25800 ( .A(n25141), .B(n25140), .Z(n25148) );
  XNOR U25801 ( .A(n25147), .B(n25148), .Z(n25149) );
  XNOR U25802 ( .A(n25150), .B(n25149), .Z(n25183) );
  XNOR U25803 ( .A(n25183), .B(sreg[1627]), .Z(n25185) );
  NAND U25804 ( .A(n25142), .B(sreg[1626]), .Z(n25146) );
  OR U25805 ( .A(n25144), .B(n25143), .Z(n25145) );
  AND U25806 ( .A(n25146), .B(n25145), .Z(n25184) );
  XOR U25807 ( .A(n25185), .B(n25184), .Z(c[1627]) );
  NANDN U25808 ( .A(n25148), .B(n25147), .Z(n25152) );
  NAND U25809 ( .A(n25150), .B(n25149), .Z(n25151) );
  NAND U25810 ( .A(n25152), .B(n25151), .Z(n25191) );
  NAND U25811 ( .A(b[0]), .B(a[612]), .Z(n25153) );
  XNOR U25812 ( .A(b[1]), .B(n25153), .Z(n25155) );
  NAND U25813 ( .A(n102), .B(a[611]), .Z(n25154) );
  AND U25814 ( .A(n25155), .B(n25154), .Z(n25208) );
  XOR U25815 ( .A(a[608]), .B(n42197), .Z(n25197) );
  NANDN U25816 ( .A(n25197), .B(n42173), .Z(n25158) );
  NANDN U25817 ( .A(n25156), .B(n42172), .Z(n25157) );
  NAND U25818 ( .A(n25158), .B(n25157), .Z(n25206) );
  NAND U25819 ( .A(b[7]), .B(a[604]), .Z(n25207) );
  XNOR U25820 ( .A(n25206), .B(n25207), .Z(n25209) );
  XOR U25821 ( .A(n25208), .B(n25209), .Z(n25215) );
  NANDN U25822 ( .A(n25159), .B(n42093), .Z(n25161) );
  XOR U25823 ( .A(n42134), .B(a[610]), .Z(n25200) );
  NANDN U25824 ( .A(n25200), .B(n42095), .Z(n25160) );
  NAND U25825 ( .A(n25161), .B(n25160), .Z(n25213) );
  NANDN U25826 ( .A(n25162), .B(n42231), .Z(n25164) );
  XOR U25827 ( .A(n212), .B(a[606]), .Z(n25203) );
  NANDN U25828 ( .A(n25203), .B(n42234), .Z(n25163) );
  AND U25829 ( .A(n25164), .B(n25163), .Z(n25212) );
  XNOR U25830 ( .A(n25213), .B(n25212), .Z(n25214) );
  XNOR U25831 ( .A(n25215), .B(n25214), .Z(n25219) );
  NANDN U25832 ( .A(n25166), .B(n25165), .Z(n25170) );
  NAND U25833 ( .A(n25168), .B(n25167), .Z(n25169) );
  AND U25834 ( .A(n25170), .B(n25169), .Z(n25218) );
  XOR U25835 ( .A(n25219), .B(n25218), .Z(n25220) );
  NANDN U25836 ( .A(n25172), .B(n25171), .Z(n25176) );
  NANDN U25837 ( .A(n25174), .B(n25173), .Z(n25175) );
  NAND U25838 ( .A(n25176), .B(n25175), .Z(n25221) );
  XOR U25839 ( .A(n25220), .B(n25221), .Z(n25188) );
  OR U25840 ( .A(n25178), .B(n25177), .Z(n25182) );
  NANDN U25841 ( .A(n25180), .B(n25179), .Z(n25181) );
  NAND U25842 ( .A(n25182), .B(n25181), .Z(n25189) );
  XNOR U25843 ( .A(n25188), .B(n25189), .Z(n25190) );
  XNOR U25844 ( .A(n25191), .B(n25190), .Z(n25224) );
  XNOR U25845 ( .A(n25224), .B(sreg[1628]), .Z(n25226) );
  NAND U25846 ( .A(n25183), .B(sreg[1627]), .Z(n25187) );
  OR U25847 ( .A(n25185), .B(n25184), .Z(n25186) );
  AND U25848 ( .A(n25187), .B(n25186), .Z(n25225) );
  XOR U25849 ( .A(n25226), .B(n25225), .Z(c[1628]) );
  NANDN U25850 ( .A(n25189), .B(n25188), .Z(n25193) );
  NAND U25851 ( .A(n25191), .B(n25190), .Z(n25192) );
  NAND U25852 ( .A(n25193), .B(n25192), .Z(n25232) );
  NAND U25853 ( .A(b[0]), .B(a[613]), .Z(n25194) );
  XNOR U25854 ( .A(b[1]), .B(n25194), .Z(n25196) );
  NAND U25855 ( .A(n102), .B(a[612]), .Z(n25195) );
  AND U25856 ( .A(n25196), .B(n25195), .Z(n25249) );
  XOR U25857 ( .A(a[609]), .B(n42197), .Z(n25238) );
  NANDN U25858 ( .A(n25238), .B(n42173), .Z(n25199) );
  NANDN U25859 ( .A(n25197), .B(n42172), .Z(n25198) );
  NAND U25860 ( .A(n25199), .B(n25198), .Z(n25247) );
  NAND U25861 ( .A(b[7]), .B(a[605]), .Z(n25248) );
  XNOR U25862 ( .A(n25247), .B(n25248), .Z(n25250) );
  XOR U25863 ( .A(n25249), .B(n25250), .Z(n25256) );
  NANDN U25864 ( .A(n25200), .B(n42093), .Z(n25202) );
  XOR U25865 ( .A(n42134), .B(a[611]), .Z(n25241) );
  NANDN U25866 ( .A(n25241), .B(n42095), .Z(n25201) );
  NAND U25867 ( .A(n25202), .B(n25201), .Z(n25254) );
  NANDN U25868 ( .A(n25203), .B(n42231), .Z(n25205) );
  XOR U25869 ( .A(n212), .B(a[607]), .Z(n25244) );
  NANDN U25870 ( .A(n25244), .B(n42234), .Z(n25204) );
  AND U25871 ( .A(n25205), .B(n25204), .Z(n25253) );
  XNOR U25872 ( .A(n25254), .B(n25253), .Z(n25255) );
  XNOR U25873 ( .A(n25256), .B(n25255), .Z(n25260) );
  NANDN U25874 ( .A(n25207), .B(n25206), .Z(n25211) );
  NAND U25875 ( .A(n25209), .B(n25208), .Z(n25210) );
  AND U25876 ( .A(n25211), .B(n25210), .Z(n25259) );
  XOR U25877 ( .A(n25260), .B(n25259), .Z(n25261) );
  NANDN U25878 ( .A(n25213), .B(n25212), .Z(n25217) );
  NANDN U25879 ( .A(n25215), .B(n25214), .Z(n25216) );
  NAND U25880 ( .A(n25217), .B(n25216), .Z(n25262) );
  XOR U25881 ( .A(n25261), .B(n25262), .Z(n25229) );
  OR U25882 ( .A(n25219), .B(n25218), .Z(n25223) );
  NANDN U25883 ( .A(n25221), .B(n25220), .Z(n25222) );
  NAND U25884 ( .A(n25223), .B(n25222), .Z(n25230) );
  XNOR U25885 ( .A(n25229), .B(n25230), .Z(n25231) );
  XNOR U25886 ( .A(n25232), .B(n25231), .Z(n25265) );
  XNOR U25887 ( .A(n25265), .B(sreg[1629]), .Z(n25267) );
  NAND U25888 ( .A(n25224), .B(sreg[1628]), .Z(n25228) );
  OR U25889 ( .A(n25226), .B(n25225), .Z(n25227) );
  AND U25890 ( .A(n25228), .B(n25227), .Z(n25266) );
  XOR U25891 ( .A(n25267), .B(n25266), .Z(c[1629]) );
  NANDN U25892 ( .A(n25230), .B(n25229), .Z(n25234) );
  NAND U25893 ( .A(n25232), .B(n25231), .Z(n25233) );
  NAND U25894 ( .A(n25234), .B(n25233), .Z(n25273) );
  NAND U25895 ( .A(b[0]), .B(a[614]), .Z(n25235) );
  XNOR U25896 ( .A(b[1]), .B(n25235), .Z(n25237) );
  NAND U25897 ( .A(n102), .B(a[613]), .Z(n25236) );
  AND U25898 ( .A(n25237), .B(n25236), .Z(n25290) );
  XOR U25899 ( .A(a[610]), .B(n42197), .Z(n25279) );
  NANDN U25900 ( .A(n25279), .B(n42173), .Z(n25240) );
  NANDN U25901 ( .A(n25238), .B(n42172), .Z(n25239) );
  NAND U25902 ( .A(n25240), .B(n25239), .Z(n25288) );
  NAND U25903 ( .A(b[7]), .B(a[606]), .Z(n25289) );
  XNOR U25904 ( .A(n25288), .B(n25289), .Z(n25291) );
  XOR U25905 ( .A(n25290), .B(n25291), .Z(n25297) );
  NANDN U25906 ( .A(n25241), .B(n42093), .Z(n25243) );
  XOR U25907 ( .A(n42134), .B(a[612]), .Z(n25282) );
  NANDN U25908 ( .A(n25282), .B(n42095), .Z(n25242) );
  NAND U25909 ( .A(n25243), .B(n25242), .Z(n25295) );
  NANDN U25910 ( .A(n25244), .B(n42231), .Z(n25246) );
  XOR U25911 ( .A(n212), .B(a[608]), .Z(n25285) );
  NANDN U25912 ( .A(n25285), .B(n42234), .Z(n25245) );
  AND U25913 ( .A(n25246), .B(n25245), .Z(n25294) );
  XNOR U25914 ( .A(n25295), .B(n25294), .Z(n25296) );
  XNOR U25915 ( .A(n25297), .B(n25296), .Z(n25301) );
  NANDN U25916 ( .A(n25248), .B(n25247), .Z(n25252) );
  NAND U25917 ( .A(n25250), .B(n25249), .Z(n25251) );
  AND U25918 ( .A(n25252), .B(n25251), .Z(n25300) );
  XOR U25919 ( .A(n25301), .B(n25300), .Z(n25302) );
  NANDN U25920 ( .A(n25254), .B(n25253), .Z(n25258) );
  NANDN U25921 ( .A(n25256), .B(n25255), .Z(n25257) );
  NAND U25922 ( .A(n25258), .B(n25257), .Z(n25303) );
  XOR U25923 ( .A(n25302), .B(n25303), .Z(n25270) );
  OR U25924 ( .A(n25260), .B(n25259), .Z(n25264) );
  NANDN U25925 ( .A(n25262), .B(n25261), .Z(n25263) );
  NAND U25926 ( .A(n25264), .B(n25263), .Z(n25271) );
  XNOR U25927 ( .A(n25270), .B(n25271), .Z(n25272) );
  XNOR U25928 ( .A(n25273), .B(n25272), .Z(n25306) );
  XNOR U25929 ( .A(n25306), .B(sreg[1630]), .Z(n25308) );
  NAND U25930 ( .A(n25265), .B(sreg[1629]), .Z(n25269) );
  OR U25931 ( .A(n25267), .B(n25266), .Z(n25268) );
  AND U25932 ( .A(n25269), .B(n25268), .Z(n25307) );
  XOR U25933 ( .A(n25308), .B(n25307), .Z(c[1630]) );
  NANDN U25934 ( .A(n25271), .B(n25270), .Z(n25275) );
  NAND U25935 ( .A(n25273), .B(n25272), .Z(n25274) );
  NAND U25936 ( .A(n25275), .B(n25274), .Z(n25314) );
  NAND U25937 ( .A(b[0]), .B(a[615]), .Z(n25276) );
  XNOR U25938 ( .A(b[1]), .B(n25276), .Z(n25278) );
  NAND U25939 ( .A(n102), .B(a[614]), .Z(n25277) );
  AND U25940 ( .A(n25278), .B(n25277), .Z(n25331) );
  XOR U25941 ( .A(a[611]), .B(n42197), .Z(n25320) );
  NANDN U25942 ( .A(n25320), .B(n42173), .Z(n25281) );
  NANDN U25943 ( .A(n25279), .B(n42172), .Z(n25280) );
  NAND U25944 ( .A(n25281), .B(n25280), .Z(n25329) );
  NAND U25945 ( .A(b[7]), .B(a[607]), .Z(n25330) );
  XNOR U25946 ( .A(n25329), .B(n25330), .Z(n25332) );
  XOR U25947 ( .A(n25331), .B(n25332), .Z(n25338) );
  NANDN U25948 ( .A(n25282), .B(n42093), .Z(n25284) );
  XOR U25949 ( .A(n42134), .B(a[613]), .Z(n25323) );
  NANDN U25950 ( .A(n25323), .B(n42095), .Z(n25283) );
  NAND U25951 ( .A(n25284), .B(n25283), .Z(n25336) );
  NANDN U25952 ( .A(n25285), .B(n42231), .Z(n25287) );
  XOR U25953 ( .A(n212), .B(a[609]), .Z(n25326) );
  NANDN U25954 ( .A(n25326), .B(n42234), .Z(n25286) );
  AND U25955 ( .A(n25287), .B(n25286), .Z(n25335) );
  XNOR U25956 ( .A(n25336), .B(n25335), .Z(n25337) );
  XNOR U25957 ( .A(n25338), .B(n25337), .Z(n25342) );
  NANDN U25958 ( .A(n25289), .B(n25288), .Z(n25293) );
  NAND U25959 ( .A(n25291), .B(n25290), .Z(n25292) );
  AND U25960 ( .A(n25293), .B(n25292), .Z(n25341) );
  XOR U25961 ( .A(n25342), .B(n25341), .Z(n25343) );
  NANDN U25962 ( .A(n25295), .B(n25294), .Z(n25299) );
  NANDN U25963 ( .A(n25297), .B(n25296), .Z(n25298) );
  NAND U25964 ( .A(n25299), .B(n25298), .Z(n25344) );
  XOR U25965 ( .A(n25343), .B(n25344), .Z(n25311) );
  OR U25966 ( .A(n25301), .B(n25300), .Z(n25305) );
  NANDN U25967 ( .A(n25303), .B(n25302), .Z(n25304) );
  NAND U25968 ( .A(n25305), .B(n25304), .Z(n25312) );
  XNOR U25969 ( .A(n25311), .B(n25312), .Z(n25313) );
  XNOR U25970 ( .A(n25314), .B(n25313), .Z(n25347) );
  XNOR U25971 ( .A(n25347), .B(sreg[1631]), .Z(n25349) );
  NAND U25972 ( .A(n25306), .B(sreg[1630]), .Z(n25310) );
  OR U25973 ( .A(n25308), .B(n25307), .Z(n25309) );
  AND U25974 ( .A(n25310), .B(n25309), .Z(n25348) );
  XOR U25975 ( .A(n25349), .B(n25348), .Z(c[1631]) );
  NANDN U25976 ( .A(n25312), .B(n25311), .Z(n25316) );
  NAND U25977 ( .A(n25314), .B(n25313), .Z(n25315) );
  NAND U25978 ( .A(n25316), .B(n25315), .Z(n25355) );
  NAND U25979 ( .A(b[0]), .B(a[616]), .Z(n25317) );
  XNOR U25980 ( .A(b[1]), .B(n25317), .Z(n25319) );
  NAND U25981 ( .A(n103), .B(a[615]), .Z(n25318) );
  AND U25982 ( .A(n25319), .B(n25318), .Z(n25372) );
  XOR U25983 ( .A(a[612]), .B(n42197), .Z(n25361) );
  NANDN U25984 ( .A(n25361), .B(n42173), .Z(n25322) );
  NANDN U25985 ( .A(n25320), .B(n42172), .Z(n25321) );
  NAND U25986 ( .A(n25322), .B(n25321), .Z(n25370) );
  NAND U25987 ( .A(b[7]), .B(a[608]), .Z(n25371) );
  XNOR U25988 ( .A(n25370), .B(n25371), .Z(n25373) );
  XOR U25989 ( .A(n25372), .B(n25373), .Z(n25379) );
  NANDN U25990 ( .A(n25323), .B(n42093), .Z(n25325) );
  XOR U25991 ( .A(n42134), .B(a[614]), .Z(n25364) );
  NANDN U25992 ( .A(n25364), .B(n42095), .Z(n25324) );
  NAND U25993 ( .A(n25325), .B(n25324), .Z(n25377) );
  NANDN U25994 ( .A(n25326), .B(n42231), .Z(n25328) );
  XOR U25995 ( .A(n212), .B(a[610]), .Z(n25367) );
  NANDN U25996 ( .A(n25367), .B(n42234), .Z(n25327) );
  AND U25997 ( .A(n25328), .B(n25327), .Z(n25376) );
  XNOR U25998 ( .A(n25377), .B(n25376), .Z(n25378) );
  XNOR U25999 ( .A(n25379), .B(n25378), .Z(n25383) );
  NANDN U26000 ( .A(n25330), .B(n25329), .Z(n25334) );
  NAND U26001 ( .A(n25332), .B(n25331), .Z(n25333) );
  AND U26002 ( .A(n25334), .B(n25333), .Z(n25382) );
  XOR U26003 ( .A(n25383), .B(n25382), .Z(n25384) );
  NANDN U26004 ( .A(n25336), .B(n25335), .Z(n25340) );
  NANDN U26005 ( .A(n25338), .B(n25337), .Z(n25339) );
  NAND U26006 ( .A(n25340), .B(n25339), .Z(n25385) );
  XOR U26007 ( .A(n25384), .B(n25385), .Z(n25352) );
  OR U26008 ( .A(n25342), .B(n25341), .Z(n25346) );
  NANDN U26009 ( .A(n25344), .B(n25343), .Z(n25345) );
  NAND U26010 ( .A(n25346), .B(n25345), .Z(n25353) );
  XNOR U26011 ( .A(n25352), .B(n25353), .Z(n25354) );
  XNOR U26012 ( .A(n25355), .B(n25354), .Z(n25388) );
  XNOR U26013 ( .A(n25388), .B(sreg[1632]), .Z(n25390) );
  NAND U26014 ( .A(n25347), .B(sreg[1631]), .Z(n25351) );
  OR U26015 ( .A(n25349), .B(n25348), .Z(n25350) );
  AND U26016 ( .A(n25351), .B(n25350), .Z(n25389) );
  XOR U26017 ( .A(n25390), .B(n25389), .Z(c[1632]) );
  NANDN U26018 ( .A(n25353), .B(n25352), .Z(n25357) );
  NAND U26019 ( .A(n25355), .B(n25354), .Z(n25356) );
  NAND U26020 ( .A(n25357), .B(n25356), .Z(n25396) );
  NAND U26021 ( .A(b[0]), .B(a[617]), .Z(n25358) );
  XNOR U26022 ( .A(b[1]), .B(n25358), .Z(n25360) );
  NAND U26023 ( .A(n103), .B(a[616]), .Z(n25359) );
  AND U26024 ( .A(n25360), .B(n25359), .Z(n25413) );
  XOR U26025 ( .A(a[613]), .B(n42197), .Z(n25402) );
  NANDN U26026 ( .A(n25402), .B(n42173), .Z(n25363) );
  NANDN U26027 ( .A(n25361), .B(n42172), .Z(n25362) );
  NAND U26028 ( .A(n25363), .B(n25362), .Z(n25411) );
  NAND U26029 ( .A(b[7]), .B(a[609]), .Z(n25412) );
  XNOR U26030 ( .A(n25411), .B(n25412), .Z(n25414) );
  XOR U26031 ( .A(n25413), .B(n25414), .Z(n25420) );
  NANDN U26032 ( .A(n25364), .B(n42093), .Z(n25366) );
  XOR U26033 ( .A(n42134), .B(a[615]), .Z(n25405) );
  NANDN U26034 ( .A(n25405), .B(n42095), .Z(n25365) );
  NAND U26035 ( .A(n25366), .B(n25365), .Z(n25418) );
  NANDN U26036 ( .A(n25367), .B(n42231), .Z(n25369) );
  XOR U26037 ( .A(n213), .B(a[611]), .Z(n25408) );
  NANDN U26038 ( .A(n25408), .B(n42234), .Z(n25368) );
  AND U26039 ( .A(n25369), .B(n25368), .Z(n25417) );
  XNOR U26040 ( .A(n25418), .B(n25417), .Z(n25419) );
  XNOR U26041 ( .A(n25420), .B(n25419), .Z(n25424) );
  NANDN U26042 ( .A(n25371), .B(n25370), .Z(n25375) );
  NAND U26043 ( .A(n25373), .B(n25372), .Z(n25374) );
  AND U26044 ( .A(n25375), .B(n25374), .Z(n25423) );
  XOR U26045 ( .A(n25424), .B(n25423), .Z(n25425) );
  NANDN U26046 ( .A(n25377), .B(n25376), .Z(n25381) );
  NANDN U26047 ( .A(n25379), .B(n25378), .Z(n25380) );
  NAND U26048 ( .A(n25381), .B(n25380), .Z(n25426) );
  XOR U26049 ( .A(n25425), .B(n25426), .Z(n25393) );
  OR U26050 ( .A(n25383), .B(n25382), .Z(n25387) );
  NANDN U26051 ( .A(n25385), .B(n25384), .Z(n25386) );
  NAND U26052 ( .A(n25387), .B(n25386), .Z(n25394) );
  XNOR U26053 ( .A(n25393), .B(n25394), .Z(n25395) );
  XNOR U26054 ( .A(n25396), .B(n25395), .Z(n25429) );
  XNOR U26055 ( .A(n25429), .B(sreg[1633]), .Z(n25431) );
  NAND U26056 ( .A(n25388), .B(sreg[1632]), .Z(n25392) );
  OR U26057 ( .A(n25390), .B(n25389), .Z(n25391) );
  AND U26058 ( .A(n25392), .B(n25391), .Z(n25430) );
  XOR U26059 ( .A(n25431), .B(n25430), .Z(c[1633]) );
  NANDN U26060 ( .A(n25394), .B(n25393), .Z(n25398) );
  NAND U26061 ( .A(n25396), .B(n25395), .Z(n25397) );
  NAND U26062 ( .A(n25398), .B(n25397), .Z(n25437) );
  NAND U26063 ( .A(b[0]), .B(a[618]), .Z(n25399) );
  XNOR U26064 ( .A(b[1]), .B(n25399), .Z(n25401) );
  NAND U26065 ( .A(n103), .B(a[617]), .Z(n25400) );
  AND U26066 ( .A(n25401), .B(n25400), .Z(n25454) );
  XOR U26067 ( .A(a[614]), .B(n42197), .Z(n25443) );
  NANDN U26068 ( .A(n25443), .B(n42173), .Z(n25404) );
  NANDN U26069 ( .A(n25402), .B(n42172), .Z(n25403) );
  NAND U26070 ( .A(n25404), .B(n25403), .Z(n25452) );
  NAND U26071 ( .A(b[7]), .B(a[610]), .Z(n25453) );
  XNOR U26072 ( .A(n25452), .B(n25453), .Z(n25455) );
  XOR U26073 ( .A(n25454), .B(n25455), .Z(n25461) );
  NANDN U26074 ( .A(n25405), .B(n42093), .Z(n25407) );
  XOR U26075 ( .A(n42134), .B(a[616]), .Z(n25446) );
  NANDN U26076 ( .A(n25446), .B(n42095), .Z(n25406) );
  NAND U26077 ( .A(n25407), .B(n25406), .Z(n25459) );
  NANDN U26078 ( .A(n25408), .B(n42231), .Z(n25410) );
  XOR U26079 ( .A(n213), .B(a[612]), .Z(n25449) );
  NANDN U26080 ( .A(n25449), .B(n42234), .Z(n25409) );
  AND U26081 ( .A(n25410), .B(n25409), .Z(n25458) );
  XNOR U26082 ( .A(n25459), .B(n25458), .Z(n25460) );
  XNOR U26083 ( .A(n25461), .B(n25460), .Z(n25465) );
  NANDN U26084 ( .A(n25412), .B(n25411), .Z(n25416) );
  NAND U26085 ( .A(n25414), .B(n25413), .Z(n25415) );
  AND U26086 ( .A(n25416), .B(n25415), .Z(n25464) );
  XOR U26087 ( .A(n25465), .B(n25464), .Z(n25466) );
  NANDN U26088 ( .A(n25418), .B(n25417), .Z(n25422) );
  NANDN U26089 ( .A(n25420), .B(n25419), .Z(n25421) );
  NAND U26090 ( .A(n25422), .B(n25421), .Z(n25467) );
  XOR U26091 ( .A(n25466), .B(n25467), .Z(n25434) );
  OR U26092 ( .A(n25424), .B(n25423), .Z(n25428) );
  NANDN U26093 ( .A(n25426), .B(n25425), .Z(n25427) );
  NAND U26094 ( .A(n25428), .B(n25427), .Z(n25435) );
  XNOR U26095 ( .A(n25434), .B(n25435), .Z(n25436) );
  XNOR U26096 ( .A(n25437), .B(n25436), .Z(n25470) );
  XNOR U26097 ( .A(n25470), .B(sreg[1634]), .Z(n25472) );
  NAND U26098 ( .A(n25429), .B(sreg[1633]), .Z(n25433) );
  OR U26099 ( .A(n25431), .B(n25430), .Z(n25432) );
  AND U26100 ( .A(n25433), .B(n25432), .Z(n25471) );
  XOR U26101 ( .A(n25472), .B(n25471), .Z(c[1634]) );
  NANDN U26102 ( .A(n25435), .B(n25434), .Z(n25439) );
  NAND U26103 ( .A(n25437), .B(n25436), .Z(n25438) );
  NAND U26104 ( .A(n25439), .B(n25438), .Z(n25478) );
  NAND U26105 ( .A(b[0]), .B(a[619]), .Z(n25440) );
  XNOR U26106 ( .A(b[1]), .B(n25440), .Z(n25442) );
  NAND U26107 ( .A(n103), .B(a[618]), .Z(n25441) );
  AND U26108 ( .A(n25442), .B(n25441), .Z(n25495) );
  XOR U26109 ( .A(a[615]), .B(n42197), .Z(n25484) );
  NANDN U26110 ( .A(n25484), .B(n42173), .Z(n25445) );
  NANDN U26111 ( .A(n25443), .B(n42172), .Z(n25444) );
  NAND U26112 ( .A(n25445), .B(n25444), .Z(n25493) );
  NAND U26113 ( .A(b[7]), .B(a[611]), .Z(n25494) );
  XNOR U26114 ( .A(n25493), .B(n25494), .Z(n25496) );
  XOR U26115 ( .A(n25495), .B(n25496), .Z(n25502) );
  NANDN U26116 ( .A(n25446), .B(n42093), .Z(n25448) );
  XOR U26117 ( .A(n42134), .B(a[617]), .Z(n25487) );
  NANDN U26118 ( .A(n25487), .B(n42095), .Z(n25447) );
  NAND U26119 ( .A(n25448), .B(n25447), .Z(n25500) );
  NANDN U26120 ( .A(n25449), .B(n42231), .Z(n25451) );
  XOR U26121 ( .A(n213), .B(a[613]), .Z(n25490) );
  NANDN U26122 ( .A(n25490), .B(n42234), .Z(n25450) );
  AND U26123 ( .A(n25451), .B(n25450), .Z(n25499) );
  XNOR U26124 ( .A(n25500), .B(n25499), .Z(n25501) );
  XNOR U26125 ( .A(n25502), .B(n25501), .Z(n25506) );
  NANDN U26126 ( .A(n25453), .B(n25452), .Z(n25457) );
  NAND U26127 ( .A(n25455), .B(n25454), .Z(n25456) );
  AND U26128 ( .A(n25457), .B(n25456), .Z(n25505) );
  XOR U26129 ( .A(n25506), .B(n25505), .Z(n25507) );
  NANDN U26130 ( .A(n25459), .B(n25458), .Z(n25463) );
  NANDN U26131 ( .A(n25461), .B(n25460), .Z(n25462) );
  NAND U26132 ( .A(n25463), .B(n25462), .Z(n25508) );
  XOR U26133 ( .A(n25507), .B(n25508), .Z(n25475) );
  OR U26134 ( .A(n25465), .B(n25464), .Z(n25469) );
  NANDN U26135 ( .A(n25467), .B(n25466), .Z(n25468) );
  NAND U26136 ( .A(n25469), .B(n25468), .Z(n25476) );
  XNOR U26137 ( .A(n25475), .B(n25476), .Z(n25477) );
  XNOR U26138 ( .A(n25478), .B(n25477), .Z(n25511) );
  XNOR U26139 ( .A(n25511), .B(sreg[1635]), .Z(n25513) );
  NAND U26140 ( .A(n25470), .B(sreg[1634]), .Z(n25474) );
  OR U26141 ( .A(n25472), .B(n25471), .Z(n25473) );
  AND U26142 ( .A(n25474), .B(n25473), .Z(n25512) );
  XOR U26143 ( .A(n25513), .B(n25512), .Z(c[1635]) );
  NANDN U26144 ( .A(n25476), .B(n25475), .Z(n25480) );
  NAND U26145 ( .A(n25478), .B(n25477), .Z(n25479) );
  NAND U26146 ( .A(n25480), .B(n25479), .Z(n25519) );
  NAND U26147 ( .A(b[0]), .B(a[620]), .Z(n25481) );
  XNOR U26148 ( .A(b[1]), .B(n25481), .Z(n25483) );
  NAND U26149 ( .A(n103), .B(a[619]), .Z(n25482) );
  AND U26150 ( .A(n25483), .B(n25482), .Z(n25536) );
  XOR U26151 ( .A(a[616]), .B(n42197), .Z(n25525) );
  NANDN U26152 ( .A(n25525), .B(n42173), .Z(n25486) );
  NANDN U26153 ( .A(n25484), .B(n42172), .Z(n25485) );
  NAND U26154 ( .A(n25486), .B(n25485), .Z(n25534) );
  NAND U26155 ( .A(b[7]), .B(a[612]), .Z(n25535) );
  XNOR U26156 ( .A(n25534), .B(n25535), .Z(n25537) );
  XOR U26157 ( .A(n25536), .B(n25537), .Z(n25543) );
  NANDN U26158 ( .A(n25487), .B(n42093), .Z(n25489) );
  XOR U26159 ( .A(n42134), .B(a[618]), .Z(n25528) );
  NANDN U26160 ( .A(n25528), .B(n42095), .Z(n25488) );
  NAND U26161 ( .A(n25489), .B(n25488), .Z(n25541) );
  NANDN U26162 ( .A(n25490), .B(n42231), .Z(n25492) );
  XOR U26163 ( .A(n213), .B(a[614]), .Z(n25531) );
  NANDN U26164 ( .A(n25531), .B(n42234), .Z(n25491) );
  AND U26165 ( .A(n25492), .B(n25491), .Z(n25540) );
  XNOR U26166 ( .A(n25541), .B(n25540), .Z(n25542) );
  XNOR U26167 ( .A(n25543), .B(n25542), .Z(n25547) );
  NANDN U26168 ( .A(n25494), .B(n25493), .Z(n25498) );
  NAND U26169 ( .A(n25496), .B(n25495), .Z(n25497) );
  AND U26170 ( .A(n25498), .B(n25497), .Z(n25546) );
  XOR U26171 ( .A(n25547), .B(n25546), .Z(n25548) );
  NANDN U26172 ( .A(n25500), .B(n25499), .Z(n25504) );
  NANDN U26173 ( .A(n25502), .B(n25501), .Z(n25503) );
  NAND U26174 ( .A(n25504), .B(n25503), .Z(n25549) );
  XOR U26175 ( .A(n25548), .B(n25549), .Z(n25516) );
  OR U26176 ( .A(n25506), .B(n25505), .Z(n25510) );
  NANDN U26177 ( .A(n25508), .B(n25507), .Z(n25509) );
  NAND U26178 ( .A(n25510), .B(n25509), .Z(n25517) );
  XNOR U26179 ( .A(n25516), .B(n25517), .Z(n25518) );
  XNOR U26180 ( .A(n25519), .B(n25518), .Z(n25552) );
  XNOR U26181 ( .A(n25552), .B(sreg[1636]), .Z(n25554) );
  NAND U26182 ( .A(n25511), .B(sreg[1635]), .Z(n25515) );
  OR U26183 ( .A(n25513), .B(n25512), .Z(n25514) );
  AND U26184 ( .A(n25515), .B(n25514), .Z(n25553) );
  XOR U26185 ( .A(n25554), .B(n25553), .Z(c[1636]) );
  NANDN U26186 ( .A(n25517), .B(n25516), .Z(n25521) );
  NAND U26187 ( .A(n25519), .B(n25518), .Z(n25520) );
  NAND U26188 ( .A(n25521), .B(n25520), .Z(n25560) );
  NAND U26189 ( .A(b[0]), .B(a[621]), .Z(n25522) );
  XNOR U26190 ( .A(b[1]), .B(n25522), .Z(n25524) );
  NAND U26191 ( .A(n103), .B(a[620]), .Z(n25523) );
  AND U26192 ( .A(n25524), .B(n25523), .Z(n25577) );
  XOR U26193 ( .A(a[617]), .B(n42197), .Z(n25566) );
  NANDN U26194 ( .A(n25566), .B(n42173), .Z(n25527) );
  NANDN U26195 ( .A(n25525), .B(n42172), .Z(n25526) );
  NAND U26196 ( .A(n25527), .B(n25526), .Z(n25575) );
  NAND U26197 ( .A(b[7]), .B(a[613]), .Z(n25576) );
  XNOR U26198 ( .A(n25575), .B(n25576), .Z(n25578) );
  XOR U26199 ( .A(n25577), .B(n25578), .Z(n25584) );
  NANDN U26200 ( .A(n25528), .B(n42093), .Z(n25530) );
  XOR U26201 ( .A(n42134), .B(a[619]), .Z(n25569) );
  NANDN U26202 ( .A(n25569), .B(n42095), .Z(n25529) );
  NAND U26203 ( .A(n25530), .B(n25529), .Z(n25582) );
  NANDN U26204 ( .A(n25531), .B(n42231), .Z(n25533) );
  XOR U26205 ( .A(n213), .B(a[615]), .Z(n25572) );
  NANDN U26206 ( .A(n25572), .B(n42234), .Z(n25532) );
  AND U26207 ( .A(n25533), .B(n25532), .Z(n25581) );
  XNOR U26208 ( .A(n25582), .B(n25581), .Z(n25583) );
  XNOR U26209 ( .A(n25584), .B(n25583), .Z(n25588) );
  NANDN U26210 ( .A(n25535), .B(n25534), .Z(n25539) );
  NAND U26211 ( .A(n25537), .B(n25536), .Z(n25538) );
  AND U26212 ( .A(n25539), .B(n25538), .Z(n25587) );
  XOR U26213 ( .A(n25588), .B(n25587), .Z(n25589) );
  NANDN U26214 ( .A(n25541), .B(n25540), .Z(n25545) );
  NANDN U26215 ( .A(n25543), .B(n25542), .Z(n25544) );
  NAND U26216 ( .A(n25545), .B(n25544), .Z(n25590) );
  XOR U26217 ( .A(n25589), .B(n25590), .Z(n25557) );
  OR U26218 ( .A(n25547), .B(n25546), .Z(n25551) );
  NANDN U26219 ( .A(n25549), .B(n25548), .Z(n25550) );
  NAND U26220 ( .A(n25551), .B(n25550), .Z(n25558) );
  XNOR U26221 ( .A(n25557), .B(n25558), .Z(n25559) );
  XNOR U26222 ( .A(n25560), .B(n25559), .Z(n25593) );
  XNOR U26223 ( .A(n25593), .B(sreg[1637]), .Z(n25595) );
  NAND U26224 ( .A(n25552), .B(sreg[1636]), .Z(n25556) );
  OR U26225 ( .A(n25554), .B(n25553), .Z(n25555) );
  AND U26226 ( .A(n25556), .B(n25555), .Z(n25594) );
  XOR U26227 ( .A(n25595), .B(n25594), .Z(c[1637]) );
  NANDN U26228 ( .A(n25558), .B(n25557), .Z(n25562) );
  NAND U26229 ( .A(n25560), .B(n25559), .Z(n25561) );
  NAND U26230 ( .A(n25562), .B(n25561), .Z(n25601) );
  NAND U26231 ( .A(b[0]), .B(a[622]), .Z(n25563) );
  XNOR U26232 ( .A(b[1]), .B(n25563), .Z(n25565) );
  NAND U26233 ( .A(n103), .B(a[621]), .Z(n25564) );
  AND U26234 ( .A(n25565), .B(n25564), .Z(n25618) );
  XOR U26235 ( .A(a[618]), .B(n42197), .Z(n25607) );
  NANDN U26236 ( .A(n25607), .B(n42173), .Z(n25568) );
  NANDN U26237 ( .A(n25566), .B(n42172), .Z(n25567) );
  NAND U26238 ( .A(n25568), .B(n25567), .Z(n25616) );
  NAND U26239 ( .A(b[7]), .B(a[614]), .Z(n25617) );
  XNOR U26240 ( .A(n25616), .B(n25617), .Z(n25619) );
  XOR U26241 ( .A(n25618), .B(n25619), .Z(n25625) );
  NANDN U26242 ( .A(n25569), .B(n42093), .Z(n25571) );
  XOR U26243 ( .A(n42134), .B(a[620]), .Z(n25610) );
  NANDN U26244 ( .A(n25610), .B(n42095), .Z(n25570) );
  NAND U26245 ( .A(n25571), .B(n25570), .Z(n25623) );
  NANDN U26246 ( .A(n25572), .B(n42231), .Z(n25574) );
  XOR U26247 ( .A(n213), .B(a[616]), .Z(n25613) );
  NANDN U26248 ( .A(n25613), .B(n42234), .Z(n25573) );
  AND U26249 ( .A(n25574), .B(n25573), .Z(n25622) );
  XNOR U26250 ( .A(n25623), .B(n25622), .Z(n25624) );
  XNOR U26251 ( .A(n25625), .B(n25624), .Z(n25629) );
  NANDN U26252 ( .A(n25576), .B(n25575), .Z(n25580) );
  NAND U26253 ( .A(n25578), .B(n25577), .Z(n25579) );
  AND U26254 ( .A(n25580), .B(n25579), .Z(n25628) );
  XOR U26255 ( .A(n25629), .B(n25628), .Z(n25630) );
  NANDN U26256 ( .A(n25582), .B(n25581), .Z(n25586) );
  NANDN U26257 ( .A(n25584), .B(n25583), .Z(n25585) );
  NAND U26258 ( .A(n25586), .B(n25585), .Z(n25631) );
  XOR U26259 ( .A(n25630), .B(n25631), .Z(n25598) );
  OR U26260 ( .A(n25588), .B(n25587), .Z(n25592) );
  NANDN U26261 ( .A(n25590), .B(n25589), .Z(n25591) );
  NAND U26262 ( .A(n25592), .B(n25591), .Z(n25599) );
  XNOR U26263 ( .A(n25598), .B(n25599), .Z(n25600) );
  XNOR U26264 ( .A(n25601), .B(n25600), .Z(n25634) );
  XNOR U26265 ( .A(n25634), .B(sreg[1638]), .Z(n25636) );
  NAND U26266 ( .A(n25593), .B(sreg[1637]), .Z(n25597) );
  OR U26267 ( .A(n25595), .B(n25594), .Z(n25596) );
  AND U26268 ( .A(n25597), .B(n25596), .Z(n25635) );
  XOR U26269 ( .A(n25636), .B(n25635), .Z(c[1638]) );
  NANDN U26270 ( .A(n25599), .B(n25598), .Z(n25603) );
  NAND U26271 ( .A(n25601), .B(n25600), .Z(n25602) );
  NAND U26272 ( .A(n25603), .B(n25602), .Z(n25642) );
  NAND U26273 ( .A(b[0]), .B(a[623]), .Z(n25604) );
  XNOR U26274 ( .A(b[1]), .B(n25604), .Z(n25606) );
  NAND U26275 ( .A(n104), .B(a[622]), .Z(n25605) );
  AND U26276 ( .A(n25606), .B(n25605), .Z(n25659) );
  XOR U26277 ( .A(a[619]), .B(n42197), .Z(n25648) );
  NANDN U26278 ( .A(n25648), .B(n42173), .Z(n25609) );
  NANDN U26279 ( .A(n25607), .B(n42172), .Z(n25608) );
  NAND U26280 ( .A(n25609), .B(n25608), .Z(n25657) );
  NAND U26281 ( .A(b[7]), .B(a[615]), .Z(n25658) );
  XNOR U26282 ( .A(n25657), .B(n25658), .Z(n25660) );
  XOR U26283 ( .A(n25659), .B(n25660), .Z(n25666) );
  NANDN U26284 ( .A(n25610), .B(n42093), .Z(n25612) );
  XOR U26285 ( .A(n42134), .B(a[621]), .Z(n25651) );
  NANDN U26286 ( .A(n25651), .B(n42095), .Z(n25611) );
  NAND U26287 ( .A(n25612), .B(n25611), .Z(n25664) );
  NANDN U26288 ( .A(n25613), .B(n42231), .Z(n25615) );
  XOR U26289 ( .A(n213), .B(a[617]), .Z(n25654) );
  NANDN U26290 ( .A(n25654), .B(n42234), .Z(n25614) );
  AND U26291 ( .A(n25615), .B(n25614), .Z(n25663) );
  XNOR U26292 ( .A(n25664), .B(n25663), .Z(n25665) );
  XNOR U26293 ( .A(n25666), .B(n25665), .Z(n25670) );
  NANDN U26294 ( .A(n25617), .B(n25616), .Z(n25621) );
  NAND U26295 ( .A(n25619), .B(n25618), .Z(n25620) );
  AND U26296 ( .A(n25621), .B(n25620), .Z(n25669) );
  XOR U26297 ( .A(n25670), .B(n25669), .Z(n25671) );
  NANDN U26298 ( .A(n25623), .B(n25622), .Z(n25627) );
  NANDN U26299 ( .A(n25625), .B(n25624), .Z(n25626) );
  NAND U26300 ( .A(n25627), .B(n25626), .Z(n25672) );
  XOR U26301 ( .A(n25671), .B(n25672), .Z(n25639) );
  OR U26302 ( .A(n25629), .B(n25628), .Z(n25633) );
  NANDN U26303 ( .A(n25631), .B(n25630), .Z(n25632) );
  NAND U26304 ( .A(n25633), .B(n25632), .Z(n25640) );
  XNOR U26305 ( .A(n25639), .B(n25640), .Z(n25641) );
  XNOR U26306 ( .A(n25642), .B(n25641), .Z(n25675) );
  XNOR U26307 ( .A(n25675), .B(sreg[1639]), .Z(n25677) );
  NAND U26308 ( .A(n25634), .B(sreg[1638]), .Z(n25638) );
  OR U26309 ( .A(n25636), .B(n25635), .Z(n25637) );
  AND U26310 ( .A(n25638), .B(n25637), .Z(n25676) );
  XOR U26311 ( .A(n25677), .B(n25676), .Z(c[1639]) );
  NANDN U26312 ( .A(n25640), .B(n25639), .Z(n25644) );
  NAND U26313 ( .A(n25642), .B(n25641), .Z(n25643) );
  NAND U26314 ( .A(n25644), .B(n25643), .Z(n25683) );
  NAND U26315 ( .A(b[0]), .B(a[624]), .Z(n25645) );
  XNOR U26316 ( .A(b[1]), .B(n25645), .Z(n25647) );
  NAND U26317 ( .A(n104), .B(a[623]), .Z(n25646) );
  AND U26318 ( .A(n25647), .B(n25646), .Z(n25700) );
  XOR U26319 ( .A(a[620]), .B(n42197), .Z(n25689) );
  NANDN U26320 ( .A(n25689), .B(n42173), .Z(n25650) );
  NANDN U26321 ( .A(n25648), .B(n42172), .Z(n25649) );
  NAND U26322 ( .A(n25650), .B(n25649), .Z(n25698) );
  NAND U26323 ( .A(b[7]), .B(a[616]), .Z(n25699) );
  XNOR U26324 ( .A(n25698), .B(n25699), .Z(n25701) );
  XOR U26325 ( .A(n25700), .B(n25701), .Z(n25707) );
  NANDN U26326 ( .A(n25651), .B(n42093), .Z(n25653) );
  XOR U26327 ( .A(n42134), .B(a[622]), .Z(n25692) );
  NANDN U26328 ( .A(n25692), .B(n42095), .Z(n25652) );
  NAND U26329 ( .A(n25653), .B(n25652), .Z(n25705) );
  NANDN U26330 ( .A(n25654), .B(n42231), .Z(n25656) );
  XOR U26331 ( .A(n213), .B(a[618]), .Z(n25695) );
  NANDN U26332 ( .A(n25695), .B(n42234), .Z(n25655) );
  AND U26333 ( .A(n25656), .B(n25655), .Z(n25704) );
  XNOR U26334 ( .A(n25705), .B(n25704), .Z(n25706) );
  XNOR U26335 ( .A(n25707), .B(n25706), .Z(n25711) );
  NANDN U26336 ( .A(n25658), .B(n25657), .Z(n25662) );
  NAND U26337 ( .A(n25660), .B(n25659), .Z(n25661) );
  AND U26338 ( .A(n25662), .B(n25661), .Z(n25710) );
  XOR U26339 ( .A(n25711), .B(n25710), .Z(n25712) );
  NANDN U26340 ( .A(n25664), .B(n25663), .Z(n25668) );
  NANDN U26341 ( .A(n25666), .B(n25665), .Z(n25667) );
  NAND U26342 ( .A(n25668), .B(n25667), .Z(n25713) );
  XOR U26343 ( .A(n25712), .B(n25713), .Z(n25680) );
  OR U26344 ( .A(n25670), .B(n25669), .Z(n25674) );
  NANDN U26345 ( .A(n25672), .B(n25671), .Z(n25673) );
  NAND U26346 ( .A(n25674), .B(n25673), .Z(n25681) );
  XNOR U26347 ( .A(n25680), .B(n25681), .Z(n25682) );
  XNOR U26348 ( .A(n25683), .B(n25682), .Z(n25716) );
  XNOR U26349 ( .A(n25716), .B(sreg[1640]), .Z(n25718) );
  NAND U26350 ( .A(n25675), .B(sreg[1639]), .Z(n25679) );
  OR U26351 ( .A(n25677), .B(n25676), .Z(n25678) );
  AND U26352 ( .A(n25679), .B(n25678), .Z(n25717) );
  XOR U26353 ( .A(n25718), .B(n25717), .Z(c[1640]) );
  NANDN U26354 ( .A(n25681), .B(n25680), .Z(n25685) );
  NAND U26355 ( .A(n25683), .B(n25682), .Z(n25684) );
  NAND U26356 ( .A(n25685), .B(n25684), .Z(n25724) );
  NAND U26357 ( .A(b[0]), .B(a[625]), .Z(n25686) );
  XNOR U26358 ( .A(b[1]), .B(n25686), .Z(n25688) );
  NAND U26359 ( .A(n104), .B(a[624]), .Z(n25687) );
  AND U26360 ( .A(n25688), .B(n25687), .Z(n25741) );
  XOR U26361 ( .A(a[621]), .B(n42197), .Z(n25730) );
  NANDN U26362 ( .A(n25730), .B(n42173), .Z(n25691) );
  NANDN U26363 ( .A(n25689), .B(n42172), .Z(n25690) );
  NAND U26364 ( .A(n25691), .B(n25690), .Z(n25739) );
  NAND U26365 ( .A(b[7]), .B(a[617]), .Z(n25740) );
  XNOR U26366 ( .A(n25739), .B(n25740), .Z(n25742) );
  XOR U26367 ( .A(n25741), .B(n25742), .Z(n25748) );
  NANDN U26368 ( .A(n25692), .B(n42093), .Z(n25694) );
  XOR U26369 ( .A(n42134), .B(a[623]), .Z(n25733) );
  NANDN U26370 ( .A(n25733), .B(n42095), .Z(n25693) );
  NAND U26371 ( .A(n25694), .B(n25693), .Z(n25746) );
  NANDN U26372 ( .A(n25695), .B(n42231), .Z(n25697) );
  XOR U26373 ( .A(n213), .B(a[619]), .Z(n25736) );
  NANDN U26374 ( .A(n25736), .B(n42234), .Z(n25696) );
  AND U26375 ( .A(n25697), .B(n25696), .Z(n25745) );
  XNOR U26376 ( .A(n25746), .B(n25745), .Z(n25747) );
  XNOR U26377 ( .A(n25748), .B(n25747), .Z(n25752) );
  NANDN U26378 ( .A(n25699), .B(n25698), .Z(n25703) );
  NAND U26379 ( .A(n25701), .B(n25700), .Z(n25702) );
  AND U26380 ( .A(n25703), .B(n25702), .Z(n25751) );
  XOR U26381 ( .A(n25752), .B(n25751), .Z(n25753) );
  NANDN U26382 ( .A(n25705), .B(n25704), .Z(n25709) );
  NANDN U26383 ( .A(n25707), .B(n25706), .Z(n25708) );
  NAND U26384 ( .A(n25709), .B(n25708), .Z(n25754) );
  XOR U26385 ( .A(n25753), .B(n25754), .Z(n25721) );
  OR U26386 ( .A(n25711), .B(n25710), .Z(n25715) );
  NANDN U26387 ( .A(n25713), .B(n25712), .Z(n25714) );
  NAND U26388 ( .A(n25715), .B(n25714), .Z(n25722) );
  XNOR U26389 ( .A(n25721), .B(n25722), .Z(n25723) );
  XNOR U26390 ( .A(n25724), .B(n25723), .Z(n25757) );
  XNOR U26391 ( .A(n25757), .B(sreg[1641]), .Z(n25759) );
  NAND U26392 ( .A(n25716), .B(sreg[1640]), .Z(n25720) );
  OR U26393 ( .A(n25718), .B(n25717), .Z(n25719) );
  AND U26394 ( .A(n25720), .B(n25719), .Z(n25758) );
  XOR U26395 ( .A(n25759), .B(n25758), .Z(c[1641]) );
  NANDN U26396 ( .A(n25722), .B(n25721), .Z(n25726) );
  NAND U26397 ( .A(n25724), .B(n25723), .Z(n25725) );
  NAND U26398 ( .A(n25726), .B(n25725), .Z(n25765) );
  NAND U26399 ( .A(b[0]), .B(a[626]), .Z(n25727) );
  XNOR U26400 ( .A(b[1]), .B(n25727), .Z(n25729) );
  NAND U26401 ( .A(n104), .B(a[625]), .Z(n25728) );
  AND U26402 ( .A(n25729), .B(n25728), .Z(n25782) );
  XOR U26403 ( .A(a[622]), .B(n42197), .Z(n25771) );
  NANDN U26404 ( .A(n25771), .B(n42173), .Z(n25732) );
  NANDN U26405 ( .A(n25730), .B(n42172), .Z(n25731) );
  NAND U26406 ( .A(n25732), .B(n25731), .Z(n25780) );
  NAND U26407 ( .A(b[7]), .B(a[618]), .Z(n25781) );
  XNOR U26408 ( .A(n25780), .B(n25781), .Z(n25783) );
  XOR U26409 ( .A(n25782), .B(n25783), .Z(n25789) );
  NANDN U26410 ( .A(n25733), .B(n42093), .Z(n25735) );
  XOR U26411 ( .A(n42134), .B(a[624]), .Z(n25774) );
  NANDN U26412 ( .A(n25774), .B(n42095), .Z(n25734) );
  NAND U26413 ( .A(n25735), .B(n25734), .Z(n25787) );
  NANDN U26414 ( .A(n25736), .B(n42231), .Z(n25738) );
  XOR U26415 ( .A(n213), .B(a[620]), .Z(n25777) );
  NANDN U26416 ( .A(n25777), .B(n42234), .Z(n25737) );
  AND U26417 ( .A(n25738), .B(n25737), .Z(n25786) );
  XNOR U26418 ( .A(n25787), .B(n25786), .Z(n25788) );
  XNOR U26419 ( .A(n25789), .B(n25788), .Z(n25793) );
  NANDN U26420 ( .A(n25740), .B(n25739), .Z(n25744) );
  NAND U26421 ( .A(n25742), .B(n25741), .Z(n25743) );
  AND U26422 ( .A(n25744), .B(n25743), .Z(n25792) );
  XOR U26423 ( .A(n25793), .B(n25792), .Z(n25794) );
  NANDN U26424 ( .A(n25746), .B(n25745), .Z(n25750) );
  NANDN U26425 ( .A(n25748), .B(n25747), .Z(n25749) );
  NAND U26426 ( .A(n25750), .B(n25749), .Z(n25795) );
  XOR U26427 ( .A(n25794), .B(n25795), .Z(n25762) );
  OR U26428 ( .A(n25752), .B(n25751), .Z(n25756) );
  NANDN U26429 ( .A(n25754), .B(n25753), .Z(n25755) );
  NAND U26430 ( .A(n25756), .B(n25755), .Z(n25763) );
  XNOR U26431 ( .A(n25762), .B(n25763), .Z(n25764) );
  XNOR U26432 ( .A(n25765), .B(n25764), .Z(n25798) );
  XNOR U26433 ( .A(n25798), .B(sreg[1642]), .Z(n25800) );
  NAND U26434 ( .A(n25757), .B(sreg[1641]), .Z(n25761) );
  OR U26435 ( .A(n25759), .B(n25758), .Z(n25760) );
  AND U26436 ( .A(n25761), .B(n25760), .Z(n25799) );
  XOR U26437 ( .A(n25800), .B(n25799), .Z(c[1642]) );
  NANDN U26438 ( .A(n25763), .B(n25762), .Z(n25767) );
  NAND U26439 ( .A(n25765), .B(n25764), .Z(n25766) );
  NAND U26440 ( .A(n25767), .B(n25766), .Z(n25806) );
  NAND U26441 ( .A(b[0]), .B(a[627]), .Z(n25768) );
  XNOR U26442 ( .A(b[1]), .B(n25768), .Z(n25770) );
  NAND U26443 ( .A(n104), .B(a[626]), .Z(n25769) );
  AND U26444 ( .A(n25770), .B(n25769), .Z(n25823) );
  XOR U26445 ( .A(a[623]), .B(n42197), .Z(n25812) );
  NANDN U26446 ( .A(n25812), .B(n42173), .Z(n25773) );
  NANDN U26447 ( .A(n25771), .B(n42172), .Z(n25772) );
  NAND U26448 ( .A(n25773), .B(n25772), .Z(n25821) );
  NAND U26449 ( .A(b[7]), .B(a[619]), .Z(n25822) );
  XNOR U26450 ( .A(n25821), .B(n25822), .Z(n25824) );
  XOR U26451 ( .A(n25823), .B(n25824), .Z(n25830) );
  NANDN U26452 ( .A(n25774), .B(n42093), .Z(n25776) );
  XOR U26453 ( .A(n42134), .B(a[625]), .Z(n25815) );
  NANDN U26454 ( .A(n25815), .B(n42095), .Z(n25775) );
  NAND U26455 ( .A(n25776), .B(n25775), .Z(n25828) );
  NANDN U26456 ( .A(n25777), .B(n42231), .Z(n25779) );
  XOR U26457 ( .A(n213), .B(a[621]), .Z(n25818) );
  NANDN U26458 ( .A(n25818), .B(n42234), .Z(n25778) );
  AND U26459 ( .A(n25779), .B(n25778), .Z(n25827) );
  XNOR U26460 ( .A(n25828), .B(n25827), .Z(n25829) );
  XNOR U26461 ( .A(n25830), .B(n25829), .Z(n25834) );
  NANDN U26462 ( .A(n25781), .B(n25780), .Z(n25785) );
  NAND U26463 ( .A(n25783), .B(n25782), .Z(n25784) );
  AND U26464 ( .A(n25785), .B(n25784), .Z(n25833) );
  XOR U26465 ( .A(n25834), .B(n25833), .Z(n25835) );
  NANDN U26466 ( .A(n25787), .B(n25786), .Z(n25791) );
  NANDN U26467 ( .A(n25789), .B(n25788), .Z(n25790) );
  NAND U26468 ( .A(n25791), .B(n25790), .Z(n25836) );
  XOR U26469 ( .A(n25835), .B(n25836), .Z(n25803) );
  OR U26470 ( .A(n25793), .B(n25792), .Z(n25797) );
  NANDN U26471 ( .A(n25795), .B(n25794), .Z(n25796) );
  NAND U26472 ( .A(n25797), .B(n25796), .Z(n25804) );
  XNOR U26473 ( .A(n25803), .B(n25804), .Z(n25805) );
  XNOR U26474 ( .A(n25806), .B(n25805), .Z(n25839) );
  XNOR U26475 ( .A(n25839), .B(sreg[1643]), .Z(n25841) );
  NAND U26476 ( .A(n25798), .B(sreg[1642]), .Z(n25802) );
  OR U26477 ( .A(n25800), .B(n25799), .Z(n25801) );
  AND U26478 ( .A(n25802), .B(n25801), .Z(n25840) );
  XOR U26479 ( .A(n25841), .B(n25840), .Z(c[1643]) );
  NANDN U26480 ( .A(n25804), .B(n25803), .Z(n25808) );
  NAND U26481 ( .A(n25806), .B(n25805), .Z(n25807) );
  NAND U26482 ( .A(n25808), .B(n25807), .Z(n25847) );
  NAND U26483 ( .A(b[0]), .B(a[628]), .Z(n25809) );
  XNOR U26484 ( .A(b[1]), .B(n25809), .Z(n25811) );
  NAND U26485 ( .A(n104), .B(a[627]), .Z(n25810) );
  AND U26486 ( .A(n25811), .B(n25810), .Z(n25864) );
  XOR U26487 ( .A(a[624]), .B(n42197), .Z(n25853) );
  NANDN U26488 ( .A(n25853), .B(n42173), .Z(n25814) );
  NANDN U26489 ( .A(n25812), .B(n42172), .Z(n25813) );
  NAND U26490 ( .A(n25814), .B(n25813), .Z(n25862) );
  NAND U26491 ( .A(b[7]), .B(a[620]), .Z(n25863) );
  XNOR U26492 ( .A(n25862), .B(n25863), .Z(n25865) );
  XOR U26493 ( .A(n25864), .B(n25865), .Z(n25871) );
  NANDN U26494 ( .A(n25815), .B(n42093), .Z(n25817) );
  XOR U26495 ( .A(n42134), .B(a[626]), .Z(n25856) );
  NANDN U26496 ( .A(n25856), .B(n42095), .Z(n25816) );
  NAND U26497 ( .A(n25817), .B(n25816), .Z(n25869) );
  NANDN U26498 ( .A(n25818), .B(n42231), .Z(n25820) );
  XOR U26499 ( .A(n213), .B(a[622]), .Z(n25859) );
  NANDN U26500 ( .A(n25859), .B(n42234), .Z(n25819) );
  AND U26501 ( .A(n25820), .B(n25819), .Z(n25868) );
  XNOR U26502 ( .A(n25869), .B(n25868), .Z(n25870) );
  XNOR U26503 ( .A(n25871), .B(n25870), .Z(n25875) );
  NANDN U26504 ( .A(n25822), .B(n25821), .Z(n25826) );
  NAND U26505 ( .A(n25824), .B(n25823), .Z(n25825) );
  AND U26506 ( .A(n25826), .B(n25825), .Z(n25874) );
  XOR U26507 ( .A(n25875), .B(n25874), .Z(n25876) );
  NANDN U26508 ( .A(n25828), .B(n25827), .Z(n25832) );
  NANDN U26509 ( .A(n25830), .B(n25829), .Z(n25831) );
  NAND U26510 ( .A(n25832), .B(n25831), .Z(n25877) );
  XOR U26511 ( .A(n25876), .B(n25877), .Z(n25844) );
  OR U26512 ( .A(n25834), .B(n25833), .Z(n25838) );
  NANDN U26513 ( .A(n25836), .B(n25835), .Z(n25837) );
  NAND U26514 ( .A(n25838), .B(n25837), .Z(n25845) );
  XNOR U26515 ( .A(n25844), .B(n25845), .Z(n25846) );
  XNOR U26516 ( .A(n25847), .B(n25846), .Z(n25880) );
  XNOR U26517 ( .A(n25880), .B(sreg[1644]), .Z(n25882) );
  NAND U26518 ( .A(n25839), .B(sreg[1643]), .Z(n25843) );
  OR U26519 ( .A(n25841), .B(n25840), .Z(n25842) );
  AND U26520 ( .A(n25843), .B(n25842), .Z(n25881) );
  XOR U26521 ( .A(n25882), .B(n25881), .Z(c[1644]) );
  NANDN U26522 ( .A(n25845), .B(n25844), .Z(n25849) );
  NAND U26523 ( .A(n25847), .B(n25846), .Z(n25848) );
  NAND U26524 ( .A(n25849), .B(n25848), .Z(n25888) );
  NAND U26525 ( .A(b[0]), .B(a[629]), .Z(n25850) );
  XNOR U26526 ( .A(b[1]), .B(n25850), .Z(n25852) );
  NAND U26527 ( .A(n104), .B(a[628]), .Z(n25851) );
  AND U26528 ( .A(n25852), .B(n25851), .Z(n25905) );
  XOR U26529 ( .A(a[625]), .B(n42197), .Z(n25894) );
  NANDN U26530 ( .A(n25894), .B(n42173), .Z(n25855) );
  NANDN U26531 ( .A(n25853), .B(n42172), .Z(n25854) );
  NAND U26532 ( .A(n25855), .B(n25854), .Z(n25903) );
  NAND U26533 ( .A(b[7]), .B(a[621]), .Z(n25904) );
  XNOR U26534 ( .A(n25903), .B(n25904), .Z(n25906) );
  XOR U26535 ( .A(n25905), .B(n25906), .Z(n25912) );
  NANDN U26536 ( .A(n25856), .B(n42093), .Z(n25858) );
  XOR U26537 ( .A(n42134), .B(a[627]), .Z(n25897) );
  NANDN U26538 ( .A(n25897), .B(n42095), .Z(n25857) );
  NAND U26539 ( .A(n25858), .B(n25857), .Z(n25910) );
  NANDN U26540 ( .A(n25859), .B(n42231), .Z(n25861) );
  XOR U26541 ( .A(n214), .B(a[623]), .Z(n25900) );
  NANDN U26542 ( .A(n25900), .B(n42234), .Z(n25860) );
  AND U26543 ( .A(n25861), .B(n25860), .Z(n25909) );
  XNOR U26544 ( .A(n25910), .B(n25909), .Z(n25911) );
  XNOR U26545 ( .A(n25912), .B(n25911), .Z(n25916) );
  NANDN U26546 ( .A(n25863), .B(n25862), .Z(n25867) );
  NAND U26547 ( .A(n25865), .B(n25864), .Z(n25866) );
  AND U26548 ( .A(n25867), .B(n25866), .Z(n25915) );
  XOR U26549 ( .A(n25916), .B(n25915), .Z(n25917) );
  NANDN U26550 ( .A(n25869), .B(n25868), .Z(n25873) );
  NANDN U26551 ( .A(n25871), .B(n25870), .Z(n25872) );
  NAND U26552 ( .A(n25873), .B(n25872), .Z(n25918) );
  XOR U26553 ( .A(n25917), .B(n25918), .Z(n25885) );
  OR U26554 ( .A(n25875), .B(n25874), .Z(n25879) );
  NANDN U26555 ( .A(n25877), .B(n25876), .Z(n25878) );
  NAND U26556 ( .A(n25879), .B(n25878), .Z(n25886) );
  XNOR U26557 ( .A(n25885), .B(n25886), .Z(n25887) );
  XNOR U26558 ( .A(n25888), .B(n25887), .Z(n25921) );
  XNOR U26559 ( .A(n25921), .B(sreg[1645]), .Z(n25923) );
  NAND U26560 ( .A(n25880), .B(sreg[1644]), .Z(n25884) );
  OR U26561 ( .A(n25882), .B(n25881), .Z(n25883) );
  AND U26562 ( .A(n25884), .B(n25883), .Z(n25922) );
  XOR U26563 ( .A(n25923), .B(n25922), .Z(c[1645]) );
  NANDN U26564 ( .A(n25886), .B(n25885), .Z(n25890) );
  NAND U26565 ( .A(n25888), .B(n25887), .Z(n25889) );
  NAND U26566 ( .A(n25890), .B(n25889), .Z(n25929) );
  NAND U26567 ( .A(b[0]), .B(a[630]), .Z(n25891) );
  XNOR U26568 ( .A(b[1]), .B(n25891), .Z(n25893) );
  NAND U26569 ( .A(n105), .B(a[629]), .Z(n25892) );
  AND U26570 ( .A(n25893), .B(n25892), .Z(n25946) );
  XOR U26571 ( .A(a[626]), .B(n42197), .Z(n25935) );
  NANDN U26572 ( .A(n25935), .B(n42173), .Z(n25896) );
  NANDN U26573 ( .A(n25894), .B(n42172), .Z(n25895) );
  NAND U26574 ( .A(n25896), .B(n25895), .Z(n25944) );
  NAND U26575 ( .A(b[7]), .B(a[622]), .Z(n25945) );
  XNOR U26576 ( .A(n25944), .B(n25945), .Z(n25947) );
  XOR U26577 ( .A(n25946), .B(n25947), .Z(n25953) );
  NANDN U26578 ( .A(n25897), .B(n42093), .Z(n25899) );
  XOR U26579 ( .A(n42134), .B(a[628]), .Z(n25938) );
  NANDN U26580 ( .A(n25938), .B(n42095), .Z(n25898) );
  NAND U26581 ( .A(n25899), .B(n25898), .Z(n25951) );
  NANDN U26582 ( .A(n25900), .B(n42231), .Z(n25902) );
  XOR U26583 ( .A(n214), .B(a[624]), .Z(n25941) );
  NANDN U26584 ( .A(n25941), .B(n42234), .Z(n25901) );
  AND U26585 ( .A(n25902), .B(n25901), .Z(n25950) );
  XNOR U26586 ( .A(n25951), .B(n25950), .Z(n25952) );
  XNOR U26587 ( .A(n25953), .B(n25952), .Z(n25957) );
  NANDN U26588 ( .A(n25904), .B(n25903), .Z(n25908) );
  NAND U26589 ( .A(n25906), .B(n25905), .Z(n25907) );
  AND U26590 ( .A(n25908), .B(n25907), .Z(n25956) );
  XOR U26591 ( .A(n25957), .B(n25956), .Z(n25958) );
  NANDN U26592 ( .A(n25910), .B(n25909), .Z(n25914) );
  NANDN U26593 ( .A(n25912), .B(n25911), .Z(n25913) );
  NAND U26594 ( .A(n25914), .B(n25913), .Z(n25959) );
  XOR U26595 ( .A(n25958), .B(n25959), .Z(n25926) );
  OR U26596 ( .A(n25916), .B(n25915), .Z(n25920) );
  NANDN U26597 ( .A(n25918), .B(n25917), .Z(n25919) );
  NAND U26598 ( .A(n25920), .B(n25919), .Z(n25927) );
  XNOR U26599 ( .A(n25926), .B(n25927), .Z(n25928) );
  XNOR U26600 ( .A(n25929), .B(n25928), .Z(n25962) );
  XNOR U26601 ( .A(n25962), .B(sreg[1646]), .Z(n25964) );
  NAND U26602 ( .A(n25921), .B(sreg[1645]), .Z(n25925) );
  OR U26603 ( .A(n25923), .B(n25922), .Z(n25924) );
  AND U26604 ( .A(n25925), .B(n25924), .Z(n25963) );
  XOR U26605 ( .A(n25964), .B(n25963), .Z(c[1646]) );
  NANDN U26606 ( .A(n25927), .B(n25926), .Z(n25931) );
  NAND U26607 ( .A(n25929), .B(n25928), .Z(n25930) );
  NAND U26608 ( .A(n25931), .B(n25930), .Z(n25970) );
  NAND U26609 ( .A(b[0]), .B(a[631]), .Z(n25932) );
  XNOR U26610 ( .A(b[1]), .B(n25932), .Z(n25934) );
  NAND U26611 ( .A(n105), .B(a[630]), .Z(n25933) );
  AND U26612 ( .A(n25934), .B(n25933), .Z(n25987) );
  XOR U26613 ( .A(a[627]), .B(n42197), .Z(n25976) );
  NANDN U26614 ( .A(n25976), .B(n42173), .Z(n25937) );
  NANDN U26615 ( .A(n25935), .B(n42172), .Z(n25936) );
  NAND U26616 ( .A(n25937), .B(n25936), .Z(n25985) );
  NAND U26617 ( .A(b[7]), .B(a[623]), .Z(n25986) );
  XNOR U26618 ( .A(n25985), .B(n25986), .Z(n25988) );
  XOR U26619 ( .A(n25987), .B(n25988), .Z(n25994) );
  NANDN U26620 ( .A(n25938), .B(n42093), .Z(n25940) );
  XOR U26621 ( .A(n42134), .B(a[629]), .Z(n25979) );
  NANDN U26622 ( .A(n25979), .B(n42095), .Z(n25939) );
  NAND U26623 ( .A(n25940), .B(n25939), .Z(n25992) );
  NANDN U26624 ( .A(n25941), .B(n42231), .Z(n25943) );
  XOR U26625 ( .A(n214), .B(a[625]), .Z(n25982) );
  NANDN U26626 ( .A(n25982), .B(n42234), .Z(n25942) );
  AND U26627 ( .A(n25943), .B(n25942), .Z(n25991) );
  XNOR U26628 ( .A(n25992), .B(n25991), .Z(n25993) );
  XNOR U26629 ( .A(n25994), .B(n25993), .Z(n25998) );
  NANDN U26630 ( .A(n25945), .B(n25944), .Z(n25949) );
  NAND U26631 ( .A(n25947), .B(n25946), .Z(n25948) );
  AND U26632 ( .A(n25949), .B(n25948), .Z(n25997) );
  XOR U26633 ( .A(n25998), .B(n25997), .Z(n25999) );
  NANDN U26634 ( .A(n25951), .B(n25950), .Z(n25955) );
  NANDN U26635 ( .A(n25953), .B(n25952), .Z(n25954) );
  NAND U26636 ( .A(n25955), .B(n25954), .Z(n26000) );
  XOR U26637 ( .A(n25999), .B(n26000), .Z(n25967) );
  OR U26638 ( .A(n25957), .B(n25956), .Z(n25961) );
  NANDN U26639 ( .A(n25959), .B(n25958), .Z(n25960) );
  NAND U26640 ( .A(n25961), .B(n25960), .Z(n25968) );
  XNOR U26641 ( .A(n25967), .B(n25968), .Z(n25969) );
  XNOR U26642 ( .A(n25970), .B(n25969), .Z(n26003) );
  XNOR U26643 ( .A(n26003), .B(sreg[1647]), .Z(n26005) );
  NAND U26644 ( .A(n25962), .B(sreg[1646]), .Z(n25966) );
  OR U26645 ( .A(n25964), .B(n25963), .Z(n25965) );
  AND U26646 ( .A(n25966), .B(n25965), .Z(n26004) );
  XOR U26647 ( .A(n26005), .B(n26004), .Z(c[1647]) );
  NANDN U26648 ( .A(n25968), .B(n25967), .Z(n25972) );
  NAND U26649 ( .A(n25970), .B(n25969), .Z(n25971) );
  NAND U26650 ( .A(n25972), .B(n25971), .Z(n26011) );
  NAND U26651 ( .A(b[0]), .B(a[632]), .Z(n25973) );
  XNOR U26652 ( .A(b[1]), .B(n25973), .Z(n25975) );
  NAND U26653 ( .A(n105), .B(a[631]), .Z(n25974) );
  AND U26654 ( .A(n25975), .B(n25974), .Z(n26028) );
  XOR U26655 ( .A(a[628]), .B(n42197), .Z(n26017) );
  NANDN U26656 ( .A(n26017), .B(n42173), .Z(n25978) );
  NANDN U26657 ( .A(n25976), .B(n42172), .Z(n25977) );
  NAND U26658 ( .A(n25978), .B(n25977), .Z(n26026) );
  NAND U26659 ( .A(b[7]), .B(a[624]), .Z(n26027) );
  XNOR U26660 ( .A(n26026), .B(n26027), .Z(n26029) );
  XOR U26661 ( .A(n26028), .B(n26029), .Z(n26035) );
  NANDN U26662 ( .A(n25979), .B(n42093), .Z(n25981) );
  XOR U26663 ( .A(n42134), .B(a[630]), .Z(n26020) );
  NANDN U26664 ( .A(n26020), .B(n42095), .Z(n25980) );
  NAND U26665 ( .A(n25981), .B(n25980), .Z(n26033) );
  NANDN U26666 ( .A(n25982), .B(n42231), .Z(n25984) );
  XOR U26667 ( .A(n214), .B(a[626]), .Z(n26023) );
  NANDN U26668 ( .A(n26023), .B(n42234), .Z(n25983) );
  AND U26669 ( .A(n25984), .B(n25983), .Z(n26032) );
  XNOR U26670 ( .A(n26033), .B(n26032), .Z(n26034) );
  XNOR U26671 ( .A(n26035), .B(n26034), .Z(n26039) );
  NANDN U26672 ( .A(n25986), .B(n25985), .Z(n25990) );
  NAND U26673 ( .A(n25988), .B(n25987), .Z(n25989) );
  AND U26674 ( .A(n25990), .B(n25989), .Z(n26038) );
  XOR U26675 ( .A(n26039), .B(n26038), .Z(n26040) );
  NANDN U26676 ( .A(n25992), .B(n25991), .Z(n25996) );
  NANDN U26677 ( .A(n25994), .B(n25993), .Z(n25995) );
  NAND U26678 ( .A(n25996), .B(n25995), .Z(n26041) );
  XOR U26679 ( .A(n26040), .B(n26041), .Z(n26008) );
  OR U26680 ( .A(n25998), .B(n25997), .Z(n26002) );
  NANDN U26681 ( .A(n26000), .B(n25999), .Z(n26001) );
  NAND U26682 ( .A(n26002), .B(n26001), .Z(n26009) );
  XNOR U26683 ( .A(n26008), .B(n26009), .Z(n26010) );
  XNOR U26684 ( .A(n26011), .B(n26010), .Z(n26044) );
  XNOR U26685 ( .A(n26044), .B(sreg[1648]), .Z(n26046) );
  NAND U26686 ( .A(n26003), .B(sreg[1647]), .Z(n26007) );
  OR U26687 ( .A(n26005), .B(n26004), .Z(n26006) );
  AND U26688 ( .A(n26007), .B(n26006), .Z(n26045) );
  XOR U26689 ( .A(n26046), .B(n26045), .Z(c[1648]) );
  NANDN U26690 ( .A(n26009), .B(n26008), .Z(n26013) );
  NAND U26691 ( .A(n26011), .B(n26010), .Z(n26012) );
  NAND U26692 ( .A(n26013), .B(n26012), .Z(n26052) );
  NAND U26693 ( .A(b[0]), .B(a[633]), .Z(n26014) );
  XNOR U26694 ( .A(b[1]), .B(n26014), .Z(n26016) );
  NAND U26695 ( .A(n105), .B(a[632]), .Z(n26015) );
  AND U26696 ( .A(n26016), .B(n26015), .Z(n26069) );
  XOR U26697 ( .A(a[629]), .B(n42197), .Z(n26058) );
  NANDN U26698 ( .A(n26058), .B(n42173), .Z(n26019) );
  NANDN U26699 ( .A(n26017), .B(n42172), .Z(n26018) );
  NAND U26700 ( .A(n26019), .B(n26018), .Z(n26067) );
  NAND U26701 ( .A(b[7]), .B(a[625]), .Z(n26068) );
  XNOR U26702 ( .A(n26067), .B(n26068), .Z(n26070) );
  XOR U26703 ( .A(n26069), .B(n26070), .Z(n26076) );
  NANDN U26704 ( .A(n26020), .B(n42093), .Z(n26022) );
  XOR U26705 ( .A(n42134), .B(a[631]), .Z(n26061) );
  NANDN U26706 ( .A(n26061), .B(n42095), .Z(n26021) );
  NAND U26707 ( .A(n26022), .B(n26021), .Z(n26074) );
  NANDN U26708 ( .A(n26023), .B(n42231), .Z(n26025) );
  XOR U26709 ( .A(n214), .B(a[627]), .Z(n26064) );
  NANDN U26710 ( .A(n26064), .B(n42234), .Z(n26024) );
  AND U26711 ( .A(n26025), .B(n26024), .Z(n26073) );
  XNOR U26712 ( .A(n26074), .B(n26073), .Z(n26075) );
  XNOR U26713 ( .A(n26076), .B(n26075), .Z(n26080) );
  NANDN U26714 ( .A(n26027), .B(n26026), .Z(n26031) );
  NAND U26715 ( .A(n26029), .B(n26028), .Z(n26030) );
  AND U26716 ( .A(n26031), .B(n26030), .Z(n26079) );
  XOR U26717 ( .A(n26080), .B(n26079), .Z(n26081) );
  NANDN U26718 ( .A(n26033), .B(n26032), .Z(n26037) );
  NANDN U26719 ( .A(n26035), .B(n26034), .Z(n26036) );
  NAND U26720 ( .A(n26037), .B(n26036), .Z(n26082) );
  XOR U26721 ( .A(n26081), .B(n26082), .Z(n26049) );
  OR U26722 ( .A(n26039), .B(n26038), .Z(n26043) );
  NANDN U26723 ( .A(n26041), .B(n26040), .Z(n26042) );
  NAND U26724 ( .A(n26043), .B(n26042), .Z(n26050) );
  XNOR U26725 ( .A(n26049), .B(n26050), .Z(n26051) );
  XNOR U26726 ( .A(n26052), .B(n26051), .Z(n26085) );
  XNOR U26727 ( .A(n26085), .B(sreg[1649]), .Z(n26087) );
  NAND U26728 ( .A(n26044), .B(sreg[1648]), .Z(n26048) );
  OR U26729 ( .A(n26046), .B(n26045), .Z(n26047) );
  AND U26730 ( .A(n26048), .B(n26047), .Z(n26086) );
  XOR U26731 ( .A(n26087), .B(n26086), .Z(c[1649]) );
  NANDN U26732 ( .A(n26050), .B(n26049), .Z(n26054) );
  NAND U26733 ( .A(n26052), .B(n26051), .Z(n26053) );
  NAND U26734 ( .A(n26054), .B(n26053), .Z(n26093) );
  NAND U26735 ( .A(b[0]), .B(a[634]), .Z(n26055) );
  XNOR U26736 ( .A(b[1]), .B(n26055), .Z(n26057) );
  NAND U26737 ( .A(n105), .B(a[633]), .Z(n26056) );
  AND U26738 ( .A(n26057), .B(n26056), .Z(n26110) );
  XOR U26739 ( .A(a[630]), .B(n42197), .Z(n26099) );
  NANDN U26740 ( .A(n26099), .B(n42173), .Z(n26060) );
  NANDN U26741 ( .A(n26058), .B(n42172), .Z(n26059) );
  NAND U26742 ( .A(n26060), .B(n26059), .Z(n26108) );
  NAND U26743 ( .A(b[7]), .B(a[626]), .Z(n26109) );
  XNOR U26744 ( .A(n26108), .B(n26109), .Z(n26111) );
  XOR U26745 ( .A(n26110), .B(n26111), .Z(n26117) );
  NANDN U26746 ( .A(n26061), .B(n42093), .Z(n26063) );
  XOR U26747 ( .A(n42134), .B(a[632]), .Z(n26102) );
  NANDN U26748 ( .A(n26102), .B(n42095), .Z(n26062) );
  NAND U26749 ( .A(n26063), .B(n26062), .Z(n26115) );
  NANDN U26750 ( .A(n26064), .B(n42231), .Z(n26066) );
  XOR U26751 ( .A(n214), .B(a[628]), .Z(n26105) );
  NANDN U26752 ( .A(n26105), .B(n42234), .Z(n26065) );
  AND U26753 ( .A(n26066), .B(n26065), .Z(n26114) );
  XNOR U26754 ( .A(n26115), .B(n26114), .Z(n26116) );
  XNOR U26755 ( .A(n26117), .B(n26116), .Z(n26121) );
  NANDN U26756 ( .A(n26068), .B(n26067), .Z(n26072) );
  NAND U26757 ( .A(n26070), .B(n26069), .Z(n26071) );
  AND U26758 ( .A(n26072), .B(n26071), .Z(n26120) );
  XOR U26759 ( .A(n26121), .B(n26120), .Z(n26122) );
  NANDN U26760 ( .A(n26074), .B(n26073), .Z(n26078) );
  NANDN U26761 ( .A(n26076), .B(n26075), .Z(n26077) );
  NAND U26762 ( .A(n26078), .B(n26077), .Z(n26123) );
  XOR U26763 ( .A(n26122), .B(n26123), .Z(n26090) );
  OR U26764 ( .A(n26080), .B(n26079), .Z(n26084) );
  NANDN U26765 ( .A(n26082), .B(n26081), .Z(n26083) );
  NAND U26766 ( .A(n26084), .B(n26083), .Z(n26091) );
  XNOR U26767 ( .A(n26090), .B(n26091), .Z(n26092) );
  XNOR U26768 ( .A(n26093), .B(n26092), .Z(n26126) );
  XNOR U26769 ( .A(n26126), .B(sreg[1650]), .Z(n26128) );
  NAND U26770 ( .A(n26085), .B(sreg[1649]), .Z(n26089) );
  OR U26771 ( .A(n26087), .B(n26086), .Z(n26088) );
  AND U26772 ( .A(n26089), .B(n26088), .Z(n26127) );
  XOR U26773 ( .A(n26128), .B(n26127), .Z(c[1650]) );
  NANDN U26774 ( .A(n26091), .B(n26090), .Z(n26095) );
  NAND U26775 ( .A(n26093), .B(n26092), .Z(n26094) );
  NAND U26776 ( .A(n26095), .B(n26094), .Z(n26134) );
  NAND U26777 ( .A(b[0]), .B(a[635]), .Z(n26096) );
  XNOR U26778 ( .A(b[1]), .B(n26096), .Z(n26098) );
  NAND U26779 ( .A(n105), .B(a[634]), .Z(n26097) );
  AND U26780 ( .A(n26098), .B(n26097), .Z(n26151) );
  XOR U26781 ( .A(a[631]), .B(n42197), .Z(n26140) );
  NANDN U26782 ( .A(n26140), .B(n42173), .Z(n26101) );
  NANDN U26783 ( .A(n26099), .B(n42172), .Z(n26100) );
  NAND U26784 ( .A(n26101), .B(n26100), .Z(n26149) );
  NAND U26785 ( .A(b[7]), .B(a[627]), .Z(n26150) );
  XNOR U26786 ( .A(n26149), .B(n26150), .Z(n26152) );
  XOR U26787 ( .A(n26151), .B(n26152), .Z(n26158) );
  NANDN U26788 ( .A(n26102), .B(n42093), .Z(n26104) );
  XOR U26789 ( .A(n42134), .B(a[633]), .Z(n26143) );
  NANDN U26790 ( .A(n26143), .B(n42095), .Z(n26103) );
  NAND U26791 ( .A(n26104), .B(n26103), .Z(n26156) );
  NANDN U26792 ( .A(n26105), .B(n42231), .Z(n26107) );
  XOR U26793 ( .A(n214), .B(a[629]), .Z(n26146) );
  NANDN U26794 ( .A(n26146), .B(n42234), .Z(n26106) );
  AND U26795 ( .A(n26107), .B(n26106), .Z(n26155) );
  XNOR U26796 ( .A(n26156), .B(n26155), .Z(n26157) );
  XNOR U26797 ( .A(n26158), .B(n26157), .Z(n26162) );
  NANDN U26798 ( .A(n26109), .B(n26108), .Z(n26113) );
  NAND U26799 ( .A(n26111), .B(n26110), .Z(n26112) );
  AND U26800 ( .A(n26113), .B(n26112), .Z(n26161) );
  XOR U26801 ( .A(n26162), .B(n26161), .Z(n26163) );
  NANDN U26802 ( .A(n26115), .B(n26114), .Z(n26119) );
  NANDN U26803 ( .A(n26117), .B(n26116), .Z(n26118) );
  NAND U26804 ( .A(n26119), .B(n26118), .Z(n26164) );
  XOR U26805 ( .A(n26163), .B(n26164), .Z(n26131) );
  OR U26806 ( .A(n26121), .B(n26120), .Z(n26125) );
  NANDN U26807 ( .A(n26123), .B(n26122), .Z(n26124) );
  NAND U26808 ( .A(n26125), .B(n26124), .Z(n26132) );
  XNOR U26809 ( .A(n26131), .B(n26132), .Z(n26133) );
  XNOR U26810 ( .A(n26134), .B(n26133), .Z(n26167) );
  XNOR U26811 ( .A(n26167), .B(sreg[1651]), .Z(n26169) );
  NAND U26812 ( .A(n26126), .B(sreg[1650]), .Z(n26130) );
  OR U26813 ( .A(n26128), .B(n26127), .Z(n26129) );
  AND U26814 ( .A(n26130), .B(n26129), .Z(n26168) );
  XOR U26815 ( .A(n26169), .B(n26168), .Z(c[1651]) );
  NANDN U26816 ( .A(n26132), .B(n26131), .Z(n26136) );
  NAND U26817 ( .A(n26134), .B(n26133), .Z(n26135) );
  NAND U26818 ( .A(n26136), .B(n26135), .Z(n26175) );
  NAND U26819 ( .A(b[0]), .B(a[636]), .Z(n26137) );
  XNOR U26820 ( .A(b[1]), .B(n26137), .Z(n26139) );
  NAND U26821 ( .A(n105), .B(a[635]), .Z(n26138) );
  AND U26822 ( .A(n26139), .B(n26138), .Z(n26192) );
  XOR U26823 ( .A(a[632]), .B(n42197), .Z(n26181) );
  NANDN U26824 ( .A(n26181), .B(n42173), .Z(n26142) );
  NANDN U26825 ( .A(n26140), .B(n42172), .Z(n26141) );
  NAND U26826 ( .A(n26142), .B(n26141), .Z(n26190) );
  NAND U26827 ( .A(b[7]), .B(a[628]), .Z(n26191) );
  XNOR U26828 ( .A(n26190), .B(n26191), .Z(n26193) );
  XOR U26829 ( .A(n26192), .B(n26193), .Z(n26199) );
  NANDN U26830 ( .A(n26143), .B(n42093), .Z(n26145) );
  XOR U26831 ( .A(n42134), .B(a[634]), .Z(n26184) );
  NANDN U26832 ( .A(n26184), .B(n42095), .Z(n26144) );
  NAND U26833 ( .A(n26145), .B(n26144), .Z(n26197) );
  NANDN U26834 ( .A(n26146), .B(n42231), .Z(n26148) );
  XOR U26835 ( .A(n214), .B(a[630]), .Z(n26187) );
  NANDN U26836 ( .A(n26187), .B(n42234), .Z(n26147) );
  AND U26837 ( .A(n26148), .B(n26147), .Z(n26196) );
  XNOR U26838 ( .A(n26197), .B(n26196), .Z(n26198) );
  XNOR U26839 ( .A(n26199), .B(n26198), .Z(n26203) );
  NANDN U26840 ( .A(n26150), .B(n26149), .Z(n26154) );
  NAND U26841 ( .A(n26152), .B(n26151), .Z(n26153) );
  AND U26842 ( .A(n26154), .B(n26153), .Z(n26202) );
  XOR U26843 ( .A(n26203), .B(n26202), .Z(n26204) );
  NANDN U26844 ( .A(n26156), .B(n26155), .Z(n26160) );
  NANDN U26845 ( .A(n26158), .B(n26157), .Z(n26159) );
  NAND U26846 ( .A(n26160), .B(n26159), .Z(n26205) );
  XOR U26847 ( .A(n26204), .B(n26205), .Z(n26172) );
  OR U26848 ( .A(n26162), .B(n26161), .Z(n26166) );
  NANDN U26849 ( .A(n26164), .B(n26163), .Z(n26165) );
  NAND U26850 ( .A(n26166), .B(n26165), .Z(n26173) );
  XNOR U26851 ( .A(n26172), .B(n26173), .Z(n26174) );
  XNOR U26852 ( .A(n26175), .B(n26174), .Z(n26208) );
  XNOR U26853 ( .A(n26208), .B(sreg[1652]), .Z(n26210) );
  NAND U26854 ( .A(n26167), .B(sreg[1651]), .Z(n26171) );
  OR U26855 ( .A(n26169), .B(n26168), .Z(n26170) );
  AND U26856 ( .A(n26171), .B(n26170), .Z(n26209) );
  XOR U26857 ( .A(n26210), .B(n26209), .Z(c[1652]) );
  NANDN U26858 ( .A(n26173), .B(n26172), .Z(n26177) );
  NAND U26859 ( .A(n26175), .B(n26174), .Z(n26176) );
  NAND U26860 ( .A(n26177), .B(n26176), .Z(n26216) );
  NAND U26861 ( .A(b[0]), .B(a[637]), .Z(n26178) );
  XNOR U26862 ( .A(b[1]), .B(n26178), .Z(n26180) );
  NAND U26863 ( .A(n106), .B(a[636]), .Z(n26179) );
  AND U26864 ( .A(n26180), .B(n26179), .Z(n26233) );
  XOR U26865 ( .A(a[633]), .B(n42197), .Z(n26222) );
  NANDN U26866 ( .A(n26222), .B(n42173), .Z(n26183) );
  NANDN U26867 ( .A(n26181), .B(n42172), .Z(n26182) );
  NAND U26868 ( .A(n26183), .B(n26182), .Z(n26231) );
  NAND U26869 ( .A(b[7]), .B(a[629]), .Z(n26232) );
  XNOR U26870 ( .A(n26231), .B(n26232), .Z(n26234) );
  XOR U26871 ( .A(n26233), .B(n26234), .Z(n26240) );
  NANDN U26872 ( .A(n26184), .B(n42093), .Z(n26186) );
  XOR U26873 ( .A(n42134), .B(a[635]), .Z(n26225) );
  NANDN U26874 ( .A(n26225), .B(n42095), .Z(n26185) );
  NAND U26875 ( .A(n26186), .B(n26185), .Z(n26238) );
  NANDN U26876 ( .A(n26187), .B(n42231), .Z(n26189) );
  XOR U26877 ( .A(n214), .B(a[631]), .Z(n26228) );
  NANDN U26878 ( .A(n26228), .B(n42234), .Z(n26188) );
  AND U26879 ( .A(n26189), .B(n26188), .Z(n26237) );
  XNOR U26880 ( .A(n26238), .B(n26237), .Z(n26239) );
  XNOR U26881 ( .A(n26240), .B(n26239), .Z(n26244) );
  NANDN U26882 ( .A(n26191), .B(n26190), .Z(n26195) );
  NAND U26883 ( .A(n26193), .B(n26192), .Z(n26194) );
  AND U26884 ( .A(n26195), .B(n26194), .Z(n26243) );
  XOR U26885 ( .A(n26244), .B(n26243), .Z(n26245) );
  NANDN U26886 ( .A(n26197), .B(n26196), .Z(n26201) );
  NANDN U26887 ( .A(n26199), .B(n26198), .Z(n26200) );
  NAND U26888 ( .A(n26201), .B(n26200), .Z(n26246) );
  XOR U26889 ( .A(n26245), .B(n26246), .Z(n26213) );
  OR U26890 ( .A(n26203), .B(n26202), .Z(n26207) );
  NANDN U26891 ( .A(n26205), .B(n26204), .Z(n26206) );
  NAND U26892 ( .A(n26207), .B(n26206), .Z(n26214) );
  XNOR U26893 ( .A(n26213), .B(n26214), .Z(n26215) );
  XNOR U26894 ( .A(n26216), .B(n26215), .Z(n26249) );
  XNOR U26895 ( .A(n26249), .B(sreg[1653]), .Z(n26251) );
  NAND U26896 ( .A(n26208), .B(sreg[1652]), .Z(n26212) );
  OR U26897 ( .A(n26210), .B(n26209), .Z(n26211) );
  AND U26898 ( .A(n26212), .B(n26211), .Z(n26250) );
  XOR U26899 ( .A(n26251), .B(n26250), .Z(c[1653]) );
  NANDN U26900 ( .A(n26214), .B(n26213), .Z(n26218) );
  NAND U26901 ( .A(n26216), .B(n26215), .Z(n26217) );
  NAND U26902 ( .A(n26218), .B(n26217), .Z(n26257) );
  NAND U26903 ( .A(b[0]), .B(a[638]), .Z(n26219) );
  XNOR U26904 ( .A(b[1]), .B(n26219), .Z(n26221) );
  NAND U26905 ( .A(n106), .B(a[637]), .Z(n26220) );
  AND U26906 ( .A(n26221), .B(n26220), .Z(n26274) );
  XOR U26907 ( .A(a[634]), .B(n42197), .Z(n26263) );
  NANDN U26908 ( .A(n26263), .B(n42173), .Z(n26224) );
  NANDN U26909 ( .A(n26222), .B(n42172), .Z(n26223) );
  NAND U26910 ( .A(n26224), .B(n26223), .Z(n26272) );
  NAND U26911 ( .A(b[7]), .B(a[630]), .Z(n26273) );
  XNOR U26912 ( .A(n26272), .B(n26273), .Z(n26275) );
  XOR U26913 ( .A(n26274), .B(n26275), .Z(n26281) );
  NANDN U26914 ( .A(n26225), .B(n42093), .Z(n26227) );
  XOR U26915 ( .A(n42134), .B(a[636]), .Z(n26266) );
  NANDN U26916 ( .A(n26266), .B(n42095), .Z(n26226) );
  NAND U26917 ( .A(n26227), .B(n26226), .Z(n26279) );
  NANDN U26918 ( .A(n26228), .B(n42231), .Z(n26230) );
  XOR U26919 ( .A(n214), .B(a[632]), .Z(n26269) );
  NANDN U26920 ( .A(n26269), .B(n42234), .Z(n26229) );
  AND U26921 ( .A(n26230), .B(n26229), .Z(n26278) );
  XNOR U26922 ( .A(n26279), .B(n26278), .Z(n26280) );
  XNOR U26923 ( .A(n26281), .B(n26280), .Z(n26285) );
  NANDN U26924 ( .A(n26232), .B(n26231), .Z(n26236) );
  NAND U26925 ( .A(n26234), .B(n26233), .Z(n26235) );
  AND U26926 ( .A(n26236), .B(n26235), .Z(n26284) );
  XOR U26927 ( .A(n26285), .B(n26284), .Z(n26286) );
  NANDN U26928 ( .A(n26238), .B(n26237), .Z(n26242) );
  NANDN U26929 ( .A(n26240), .B(n26239), .Z(n26241) );
  NAND U26930 ( .A(n26242), .B(n26241), .Z(n26287) );
  XOR U26931 ( .A(n26286), .B(n26287), .Z(n26254) );
  OR U26932 ( .A(n26244), .B(n26243), .Z(n26248) );
  NANDN U26933 ( .A(n26246), .B(n26245), .Z(n26247) );
  NAND U26934 ( .A(n26248), .B(n26247), .Z(n26255) );
  XNOR U26935 ( .A(n26254), .B(n26255), .Z(n26256) );
  XNOR U26936 ( .A(n26257), .B(n26256), .Z(n26290) );
  XNOR U26937 ( .A(n26290), .B(sreg[1654]), .Z(n26292) );
  NAND U26938 ( .A(n26249), .B(sreg[1653]), .Z(n26253) );
  OR U26939 ( .A(n26251), .B(n26250), .Z(n26252) );
  AND U26940 ( .A(n26253), .B(n26252), .Z(n26291) );
  XOR U26941 ( .A(n26292), .B(n26291), .Z(c[1654]) );
  NANDN U26942 ( .A(n26255), .B(n26254), .Z(n26259) );
  NAND U26943 ( .A(n26257), .B(n26256), .Z(n26258) );
  NAND U26944 ( .A(n26259), .B(n26258), .Z(n26298) );
  NAND U26945 ( .A(b[0]), .B(a[639]), .Z(n26260) );
  XNOR U26946 ( .A(b[1]), .B(n26260), .Z(n26262) );
  NAND U26947 ( .A(n106), .B(a[638]), .Z(n26261) );
  AND U26948 ( .A(n26262), .B(n26261), .Z(n26315) );
  XOR U26949 ( .A(a[635]), .B(n42197), .Z(n26304) );
  NANDN U26950 ( .A(n26304), .B(n42173), .Z(n26265) );
  NANDN U26951 ( .A(n26263), .B(n42172), .Z(n26264) );
  NAND U26952 ( .A(n26265), .B(n26264), .Z(n26313) );
  NAND U26953 ( .A(b[7]), .B(a[631]), .Z(n26314) );
  XNOR U26954 ( .A(n26313), .B(n26314), .Z(n26316) );
  XOR U26955 ( .A(n26315), .B(n26316), .Z(n26322) );
  NANDN U26956 ( .A(n26266), .B(n42093), .Z(n26268) );
  XOR U26957 ( .A(n42134), .B(a[637]), .Z(n26307) );
  NANDN U26958 ( .A(n26307), .B(n42095), .Z(n26267) );
  NAND U26959 ( .A(n26268), .B(n26267), .Z(n26320) );
  NANDN U26960 ( .A(n26269), .B(n42231), .Z(n26271) );
  XOR U26961 ( .A(n214), .B(a[633]), .Z(n26310) );
  NANDN U26962 ( .A(n26310), .B(n42234), .Z(n26270) );
  AND U26963 ( .A(n26271), .B(n26270), .Z(n26319) );
  XNOR U26964 ( .A(n26320), .B(n26319), .Z(n26321) );
  XNOR U26965 ( .A(n26322), .B(n26321), .Z(n26326) );
  NANDN U26966 ( .A(n26273), .B(n26272), .Z(n26277) );
  NAND U26967 ( .A(n26275), .B(n26274), .Z(n26276) );
  AND U26968 ( .A(n26277), .B(n26276), .Z(n26325) );
  XOR U26969 ( .A(n26326), .B(n26325), .Z(n26327) );
  NANDN U26970 ( .A(n26279), .B(n26278), .Z(n26283) );
  NANDN U26971 ( .A(n26281), .B(n26280), .Z(n26282) );
  NAND U26972 ( .A(n26283), .B(n26282), .Z(n26328) );
  XOR U26973 ( .A(n26327), .B(n26328), .Z(n26295) );
  OR U26974 ( .A(n26285), .B(n26284), .Z(n26289) );
  NANDN U26975 ( .A(n26287), .B(n26286), .Z(n26288) );
  NAND U26976 ( .A(n26289), .B(n26288), .Z(n26296) );
  XNOR U26977 ( .A(n26295), .B(n26296), .Z(n26297) );
  XNOR U26978 ( .A(n26298), .B(n26297), .Z(n26331) );
  XNOR U26979 ( .A(n26331), .B(sreg[1655]), .Z(n26333) );
  NAND U26980 ( .A(n26290), .B(sreg[1654]), .Z(n26294) );
  OR U26981 ( .A(n26292), .B(n26291), .Z(n26293) );
  AND U26982 ( .A(n26294), .B(n26293), .Z(n26332) );
  XOR U26983 ( .A(n26333), .B(n26332), .Z(c[1655]) );
  NANDN U26984 ( .A(n26296), .B(n26295), .Z(n26300) );
  NAND U26985 ( .A(n26298), .B(n26297), .Z(n26299) );
  NAND U26986 ( .A(n26300), .B(n26299), .Z(n26339) );
  NAND U26987 ( .A(b[0]), .B(a[640]), .Z(n26301) );
  XNOR U26988 ( .A(b[1]), .B(n26301), .Z(n26303) );
  NAND U26989 ( .A(n106), .B(a[639]), .Z(n26302) );
  AND U26990 ( .A(n26303), .B(n26302), .Z(n26356) );
  XOR U26991 ( .A(a[636]), .B(n42197), .Z(n26345) );
  NANDN U26992 ( .A(n26345), .B(n42173), .Z(n26306) );
  NANDN U26993 ( .A(n26304), .B(n42172), .Z(n26305) );
  NAND U26994 ( .A(n26306), .B(n26305), .Z(n26354) );
  NAND U26995 ( .A(b[7]), .B(a[632]), .Z(n26355) );
  XNOR U26996 ( .A(n26354), .B(n26355), .Z(n26357) );
  XOR U26997 ( .A(n26356), .B(n26357), .Z(n26363) );
  NANDN U26998 ( .A(n26307), .B(n42093), .Z(n26309) );
  XOR U26999 ( .A(n42134), .B(a[638]), .Z(n26348) );
  NANDN U27000 ( .A(n26348), .B(n42095), .Z(n26308) );
  NAND U27001 ( .A(n26309), .B(n26308), .Z(n26361) );
  NANDN U27002 ( .A(n26310), .B(n42231), .Z(n26312) );
  XOR U27003 ( .A(n214), .B(a[634]), .Z(n26351) );
  NANDN U27004 ( .A(n26351), .B(n42234), .Z(n26311) );
  AND U27005 ( .A(n26312), .B(n26311), .Z(n26360) );
  XNOR U27006 ( .A(n26361), .B(n26360), .Z(n26362) );
  XNOR U27007 ( .A(n26363), .B(n26362), .Z(n26367) );
  NANDN U27008 ( .A(n26314), .B(n26313), .Z(n26318) );
  NAND U27009 ( .A(n26316), .B(n26315), .Z(n26317) );
  AND U27010 ( .A(n26318), .B(n26317), .Z(n26366) );
  XOR U27011 ( .A(n26367), .B(n26366), .Z(n26368) );
  NANDN U27012 ( .A(n26320), .B(n26319), .Z(n26324) );
  NANDN U27013 ( .A(n26322), .B(n26321), .Z(n26323) );
  NAND U27014 ( .A(n26324), .B(n26323), .Z(n26369) );
  XOR U27015 ( .A(n26368), .B(n26369), .Z(n26336) );
  OR U27016 ( .A(n26326), .B(n26325), .Z(n26330) );
  NANDN U27017 ( .A(n26328), .B(n26327), .Z(n26329) );
  NAND U27018 ( .A(n26330), .B(n26329), .Z(n26337) );
  XNOR U27019 ( .A(n26336), .B(n26337), .Z(n26338) );
  XNOR U27020 ( .A(n26339), .B(n26338), .Z(n26372) );
  XNOR U27021 ( .A(n26372), .B(sreg[1656]), .Z(n26374) );
  NAND U27022 ( .A(n26331), .B(sreg[1655]), .Z(n26335) );
  OR U27023 ( .A(n26333), .B(n26332), .Z(n26334) );
  AND U27024 ( .A(n26335), .B(n26334), .Z(n26373) );
  XOR U27025 ( .A(n26374), .B(n26373), .Z(c[1656]) );
  NANDN U27026 ( .A(n26337), .B(n26336), .Z(n26341) );
  NAND U27027 ( .A(n26339), .B(n26338), .Z(n26340) );
  NAND U27028 ( .A(n26341), .B(n26340), .Z(n26380) );
  NAND U27029 ( .A(b[0]), .B(a[641]), .Z(n26342) );
  XNOR U27030 ( .A(b[1]), .B(n26342), .Z(n26344) );
  NAND U27031 ( .A(n106), .B(a[640]), .Z(n26343) );
  AND U27032 ( .A(n26344), .B(n26343), .Z(n26397) );
  XOR U27033 ( .A(a[637]), .B(n42197), .Z(n26386) );
  NANDN U27034 ( .A(n26386), .B(n42173), .Z(n26347) );
  NANDN U27035 ( .A(n26345), .B(n42172), .Z(n26346) );
  NAND U27036 ( .A(n26347), .B(n26346), .Z(n26395) );
  NAND U27037 ( .A(b[7]), .B(a[633]), .Z(n26396) );
  XNOR U27038 ( .A(n26395), .B(n26396), .Z(n26398) );
  XOR U27039 ( .A(n26397), .B(n26398), .Z(n26404) );
  NANDN U27040 ( .A(n26348), .B(n42093), .Z(n26350) );
  XOR U27041 ( .A(n42134), .B(a[639]), .Z(n26389) );
  NANDN U27042 ( .A(n26389), .B(n42095), .Z(n26349) );
  NAND U27043 ( .A(n26350), .B(n26349), .Z(n26402) );
  NANDN U27044 ( .A(n26351), .B(n42231), .Z(n26353) );
  XOR U27045 ( .A(n215), .B(a[635]), .Z(n26392) );
  NANDN U27046 ( .A(n26392), .B(n42234), .Z(n26352) );
  AND U27047 ( .A(n26353), .B(n26352), .Z(n26401) );
  XNOR U27048 ( .A(n26402), .B(n26401), .Z(n26403) );
  XNOR U27049 ( .A(n26404), .B(n26403), .Z(n26408) );
  NANDN U27050 ( .A(n26355), .B(n26354), .Z(n26359) );
  NAND U27051 ( .A(n26357), .B(n26356), .Z(n26358) );
  AND U27052 ( .A(n26359), .B(n26358), .Z(n26407) );
  XOR U27053 ( .A(n26408), .B(n26407), .Z(n26409) );
  NANDN U27054 ( .A(n26361), .B(n26360), .Z(n26365) );
  NANDN U27055 ( .A(n26363), .B(n26362), .Z(n26364) );
  NAND U27056 ( .A(n26365), .B(n26364), .Z(n26410) );
  XOR U27057 ( .A(n26409), .B(n26410), .Z(n26377) );
  OR U27058 ( .A(n26367), .B(n26366), .Z(n26371) );
  NANDN U27059 ( .A(n26369), .B(n26368), .Z(n26370) );
  NAND U27060 ( .A(n26371), .B(n26370), .Z(n26378) );
  XNOR U27061 ( .A(n26377), .B(n26378), .Z(n26379) );
  XNOR U27062 ( .A(n26380), .B(n26379), .Z(n26413) );
  XNOR U27063 ( .A(n26413), .B(sreg[1657]), .Z(n26415) );
  NAND U27064 ( .A(n26372), .B(sreg[1656]), .Z(n26376) );
  OR U27065 ( .A(n26374), .B(n26373), .Z(n26375) );
  AND U27066 ( .A(n26376), .B(n26375), .Z(n26414) );
  XOR U27067 ( .A(n26415), .B(n26414), .Z(c[1657]) );
  NANDN U27068 ( .A(n26378), .B(n26377), .Z(n26382) );
  NAND U27069 ( .A(n26380), .B(n26379), .Z(n26381) );
  NAND U27070 ( .A(n26382), .B(n26381), .Z(n26421) );
  NAND U27071 ( .A(b[0]), .B(a[642]), .Z(n26383) );
  XNOR U27072 ( .A(b[1]), .B(n26383), .Z(n26385) );
  NAND U27073 ( .A(n106), .B(a[641]), .Z(n26384) );
  AND U27074 ( .A(n26385), .B(n26384), .Z(n26438) );
  XOR U27075 ( .A(a[638]), .B(n42197), .Z(n26427) );
  NANDN U27076 ( .A(n26427), .B(n42173), .Z(n26388) );
  NANDN U27077 ( .A(n26386), .B(n42172), .Z(n26387) );
  NAND U27078 ( .A(n26388), .B(n26387), .Z(n26436) );
  NAND U27079 ( .A(b[7]), .B(a[634]), .Z(n26437) );
  XNOR U27080 ( .A(n26436), .B(n26437), .Z(n26439) );
  XOR U27081 ( .A(n26438), .B(n26439), .Z(n26445) );
  NANDN U27082 ( .A(n26389), .B(n42093), .Z(n26391) );
  XOR U27083 ( .A(n42134), .B(a[640]), .Z(n26430) );
  NANDN U27084 ( .A(n26430), .B(n42095), .Z(n26390) );
  NAND U27085 ( .A(n26391), .B(n26390), .Z(n26443) );
  NANDN U27086 ( .A(n26392), .B(n42231), .Z(n26394) );
  XOR U27087 ( .A(n215), .B(a[636]), .Z(n26433) );
  NANDN U27088 ( .A(n26433), .B(n42234), .Z(n26393) );
  AND U27089 ( .A(n26394), .B(n26393), .Z(n26442) );
  XNOR U27090 ( .A(n26443), .B(n26442), .Z(n26444) );
  XNOR U27091 ( .A(n26445), .B(n26444), .Z(n26449) );
  NANDN U27092 ( .A(n26396), .B(n26395), .Z(n26400) );
  NAND U27093 ( .A(n26398), .B(n26397), .Z(n26399) );
  AND U27094 ( .A(n26400), .B(n26399), .Z(n26448) );
  XOR U27095 ( .A(n26449), .B(n26448), .Z(n26450) );
  NANDN U27096 ( .A(n26402), .B(n26401), .Z(n26406) );
  NANDN U27097 ( .A(n26404), .B(n26403), .Z(n26405) );
  NAND U27098 ( .A(n26406), .B(n26405), .Z(n26451) );
  XOR U27099 ( .A(n26450), .B(n26451), .Z(n26418) );
  OR U27100 ( .A(n26408), .B(n26407), .Z(n26412) );
  NANDN U27101 ( .A(n26410), .B(n26409), .Z(n26411) );
  NAND U27102 ( .A(n26412), .B(n26411), .Z(n26419) );
  XNOR U27103 ( .A(n26418), .B(n26419), .Z(n26420) );
  XNOR U27104 ( .A(n26421), .B(n26420), .Z(n26454) );
  XNOR U27105 ( .A(n26454), .B(sreg[1658]), .Z(n26456) );
  NAND U27106 ( .A(n26413), .B(sreg[1657]), .Z(n26417) );
  OR U27107 ( .A(n26415), .B(n26414), .Z(n26416) );
  AND U27108 ( .A(n26417), .B(n26416), .Z(n26455) );
  XOR U27109 ( .A(n26456), .B(n26455), .Z(c[1658]) );
  NANDN U27110 ( .A(n26419), .B(n26418), .Z(n26423) );
  NAND U27111 ( .A(n26421), .B(n26420), .Z(n26422) );
  NAND U27112 ( .A(n26423), .B(n26422), .Z(n26462) );
  NAND U27113 ( .A(b[0]), .B(a[643]), .Z(n26424) );
  XNOR U27114 ( .A(b[1]), .B(n26424), .Z(n26426) );
  NAND U27115 ( .A(n106), .B(a[642]), .Z(n26425) );
  AND U27116 ( .A(n26426), .B(n26425), .Z(n26479) );
  XOR U27117 ( .A(a[639]), .B(n42197), .Z(n26468) );
  NANDN U27118 ( .A(n26468), .B(n42173), .Z(n26429) );
  NANDN U27119 ( .A(n26427), .B(n42172), .Z(n26428) );
  NAND U27120 ( .A(n26429), .B(n26428), .Z(n26477) );
  NAND U27121 ( .A(b[7]), .B(a[635]), .Z(n26478) );
  XNOR U27122 ( .A(n26477), .B(n26478), .Z(n26480) );
  XOR U27123 ( .A(n26479), .B(n26480), .Z(n26486) );
  NANDN U27124 ( .A(n26430), .B(n42093), .Z(n26432) );
  XOR U27125 ( .A(n42134), .B(a[641]), .Z(n26471) );
  NANDN U27126 ( .A(n26471), .B(n42095), .Z(n26431) );
  NAND U27127 ( .A(n26432), .B(n26431), .Z(n26484) );
  NANDN U27128 ( .A(n26433), .B(n42231), .Z(n26435) );
  XOR U27129 ( .A(n215), .B(a[637]), .Z(n26474) );
  NANDN U27130 ( .A(n26474), .B(n42234), .Z(n26434) );
  AND U27131 ( .A(n26435), .B(n26434), .Z(n26483) );
  XNOR U27132 ( .A(n26484), .B(n26483), .Z(n26485) );
  XNOR U27133 ( .A(n26486), .B(n26485), .Z(n26490) );
  NANDN U27134 ( .A(n26437), .B(n26436), .Z(n26441) );
  NAND U27135 ( .A(n26439), .B(n26438), .Z(n26440) );
  AND U27136 ( .A(n26441), .B(n26440), .Z(n26489) );
  XOR U27137 ( .A(n26490), .B(n26489), .Z(n26491) );
  NANDN U27138 ( .A(n26443), .B(n26442), .Z(n26447) );
  NANDN U27139 ( .A(n26445), .B(n26444), .Z(n26446) );
  NAND U27140 ( .A(n26447), .B(n26446), .Z(n26492) );
  XOR U27141 ( .A(n26491), .B(n26492), .Z(n26459) );
  OR U27142 ( .A(n26449), .B(n26448), .Z(n26453) );
  NANDN U27143 ( .A(n26451), .B(n26450), .Z(n26452) );
  NAND U27144 ( .A(n26453), .B(n26452), .Z(n26460) );
  XNOR U27145 ( .A(n26459), .B(n26460), .Z(n26461) );
  XNOR U27146 ( .A(n26462), .B(n26461), .Z(n26495) );
  XNOR U27147 ( .A(n26495), .B(sreg[1659]), .Z(n26497) );
  NAND U27148 ( .A(n26454), .B(sreg[1658]), .Z(n26458) );
  OR U27149 ( .A(n26456), .B(n26455), .Z(n26457) );
  AND U27150 ( .A(n26458), .B(n26457), .Z(n26496) );
  XOR U27151 ( .A(n26497), .B(n26496), .Z(c[1659]) );
  NANDN U27152 ( .A(n26460), .B(n26459), .Z(n26464) );
  NAND U27153 ( .A(n26462), .B(n26461), .Z(n26463) );
  NAND U27154 ( .A(n26464), .B(n26463), .Z(n26503) );
  NAND U27155 ( .A(b[0]), .B(a[644]), .Z(n26465) );
  XNOR U27156 ( .A(b[1]), .B(n26465), .Z(n26467) );
  NAND U27157 ( .A(n107), .B(a[643]), .Z(n26466) );
  AND U27158 ( .A(n26467), .B(n26466), .Z(n26520) );
  XOR U27159 ( .A(a[640]), .B(n42197), .Z(n26509) );
  NANDN U27160 ( .A(n26509), .B(n42173), .Z(n26470) );
  NANDN U27161 ( .A(n26468), .B(n42172), .Z(n26469) );
  NAND U27162 ( .A(n26470), .B(n26469), .Z(n26518) );
  NAND U27163 ( .A(b[7]), .B(a[636]), .Z(n26519) );
  XNOR U27164 ( .A(n26518), .B(n26519), .Z(n26521) );
  XOR U27165 ( .A(n26520), .B(n26521), .Z(n26527) );
  NANDN U27166 ( .A(n26471), .B(n42093), .Z(n26473) );
  XOR U27167 ( .A(n42134), .B(a[642]), .Z(n26512) );
  NANDN U27168 ( .A(n26512), .B(n42095), .Z(n26472) );
  NAND U27169 ( .A(n26473), .B(n26472), .Z(n26525) );
  NANDN U27170 ( .A(n26474), .B(n42231), .Z(n26476) );
  XOR U27171 ( .A(n215), .B(a[638]), .Z(n26515) );
  NANDN U27172 ( .A(n26515), .B(n42234), .Z(n26475) );
  AND U27173 ( .A(n26476), .B(n26475), .Z(n26524) );
  XNOR U27174 ( .A(n26525), .B(n26524), .Z(n26526) );
  XNOR U27175 ( .A(n26527), .B(n26526), .Z(n26531) );
  NANDN U27176 ( .A(n26478), .B(n26477), .Z(n26482) );
  NAND U27177 ( .A(n26480), .B(n26479), .Z(n26481) );
  AND U27178 ( .A(n26482), .B(n26481), .Z(n26530) );
  XOR U27179 ( .A(n26531), .B(n26530), .Z(n26532) );
  NANDN U27180 ( .A(n26484), .B(n26483), .Z(n26488) );
  NANDN U27181 ( .A(n26486), .B(n26485), .Z(n26487) );
  NAND U27182 ( .A(n26488), .B(n26487), .Z(n26533) );
  XOR U27183 ( .A(n26532), .B(n26533), .Z(n26500) );
  OR U27184 ( .A(n26490), .B(n26489), .Z(n26494) );
  NANDN U27185 ( .A(n26492), .B(n26491), .Z(n26493) );
  NAND U27186 ( .A(n26494), .B(n26493), .Z(n26501) );
  XNOR U27187 ( .A(n26500), .B(n26501), .Z(n26502) );
  XNOR U27188 ( .A(n26503), .B(n26502), .Z(n26536) );
  XNOR U27189 ( .A(n26536), .B(sreg[1660]), .Z(n26538) );
  NAND U27190 ( .A(n26495), .B(sreg[1659]), .Z(n26499) );
  OR U27191 ( .A(n26497), .B(n26496), .Z(n26498) );
  AND U27192 ( .A(n26499), .B(n26498), .Z(n26537) );
  XOR U27193 ( .A(n26538), .B(n26537), .Z(c[1660]) );
  NANDN U27194 ( .A(n26501), .B(n26500), .Z(n26505) );
  NAND U27195 ( .A(n26503), .B(n26502), .Z(n26504) );
  NAND U27196 ( .A(n26505), .B(n26504), .Z(n26544) );
  NAND U27197 ( .A(b[0]), .B(a[645]), .Z(n26506) );
  XNOR U27198 ( .A(b[1]), .B(n26506), .Z(n26508) );
  NAND U27199 ( .A(n107), .B(a[644]), .Z(n26507) );
  AND U27200 ( .A(n26508), .B(n26507), .Z(n26561) );
  XOR U27201 ( .A(a[641]), .B(n42197), .Z(n26550) );
  NANDN U27202 ( .A(n26550), .B(n42173), .Z(n26511) );
  NANDN U27203 ( .A(n26509), .B(n42172), .Z(n26510) );
  NAND U27204 ( .A(n26511), .B(n26510), .Z(n26559) );
  NAND U27205 ( .A(b[7]), .B(a[637]), .Z(n26560) );
  XNOR U27206 ( .A(n26559), .B(n26560), .Z(n26562) );
  XOR U27207 ( .A(n26561), .B(n26562), .Z(n26568) );
  NANDN U27208 ( .A(n26512), .B(n42093), .Z(n26514) );
  XOR U27209 ( .A(n42134), .B(a[643]), .Z(n26553) );
  NANDN U27210 ( .A(n26553), .B(n42095), .Z(n26513) );
  NAND U27211 ( .A(n26514), .B(n26513), .Z(n26566) );
  NANDN U27212 ( .A(n26515), .B(n42231), .Z(n26517) );
  XOR U27213 ( .A(n215), .B(a[639]), .Z(n26556) );
  NANDN U27214 ( .A(n26556), .B(n42234), .Z(n26516) );
  AND U27215 ( .A(n26517), .B(n26516), .Z(n26565) );
  XNOR U27216 ( .A(n26566), .B(n26565), .Z(n26567) );
  XNOR U27217 ( .A(n26568), .B(n26567), .Z(n26572) );
  NANDN U27218 ( .A(n26519), .B(n26518), .Z(n26523) );
  NAND U27219 ( .A(n26521), .B(n26520), .Z(n26522) );
  AND U27220 ( .A(n26523), .B(n26522), .Z(n26571) );
  XOR U27221 ( .A(n26572), .B(n26571), .Z(n26573) );
  NANDN U27222 ( .A(n26525), .B(n26524), .Z(n26529) );
  NANDN U27223 ( .A(n26527), .B(n26526), .Z(n26528) );
  NAND U27224 ( .A(n26529), .B(n26528), .Z(n26574) );
  XOR U27225 ( .A(n26573), .B(n26574), .Z(n26541) );
  OR U27226 ( .A(n26531), .B(n26530), .Z(n26535) );
  NANDN U27227 ( .A(n26533), .B(n26532), .Z(n26534) );
  NAND U27228 ( .A(n26535), .B(n26534), .Z(n26542) );
  XNOR U27229 ( .A(n26541), .B(n26542), .Z(n26543) );
  XNOR U27230 ( .A(n26544), .B(n26543), .Z(n26577) );
  XNOR U27231 ( .A(n26577), .B(sreg[1661]), .Z(n26579) );
  NAND U27232 ( .A(n26536), .B(sreg[1660]), .Z(n26540) );
  OR U27233 ( .A(n26538), .B(n26537), .Z(n26539) );
  AND U27234 ( .A(n26540), .B(n26539), .Z(n26578) );
  XOR U27235 ( .A(n26579), .B(n26578), .Z(c[1661]) );
  NANDN U27236 ( .A(n26542), .B(n26541), .Z(n26546) );
  NAND U27237 ( .A(n26544), .B(n26543), .Z(n26545) );
  NAND U27238 ( .A(n26546), .B(n26545), .Z(n26585) );
  NAND U27239 ( .A(b[0]), .B(a[646]), .Z(n26547) );
  XNOR U27240 ( .A(b[1]), .B(n26547), .Z(n26549) );
  NAND U27241 ( .A(n107), .B(a[645]), .Z(n26548) );
  AND U27242 ( .A(n26549), .B(n26548), .Z(n26602) );
  XOR U27243 ( .A(a[642]), .B(n42197), .Z(n26591) );
  NANDN U27244 ( .A(n26591), .B(n42173), .Z(n26552) );
  NANDN U27245 ( .A(n26550), .B(n42172), .Z(n26551) );
  NAND U27246 ( .A(n26552), .B(n26551), .Z(n26600) );
  NAND U27247 ( .A(b[7]), .B(a[638]), .Z(n26601) );
  XNOR U27248 ( .A(n26600), .B(n26601), .Z(n26603) );
  XOR U27249 ( .A(n26602), .B(n26603), .Z(n26609) );
  NANDN U27250 ( .A(n26553), .B(n42093), .Z(n26555) );
  XOR U27251 ( .A(n42134), .B(a[644]), .Z(n26594) );
  NANDN U27252 ( .A(n26594), .B(n42095), .Z(n26554) );
  NAND U27253 ( .A(n26555), .B(n26554), .Z(n26607) );
  NANDN U27254 ( .A(n26556), .B(n42231), .Z(n26558) );
  XOR U27255 ( .A(n215), .B(a[640]), .Z(n26597) );
  NANDN U27256 ( .A(n26597), .B(n42234), .Z(n26557) );
  AND U27257 ( .A(n26558), .B(n26557), .Z(n26606) );
  XNOR U27258 ( .A(n26607), .B(n26606), .Z(n26608) );
  XNOR U27259 ( .A(n26609), .B(n26608), .Z(n26613) );
  NANDN U27260 ( .A(n26560), .B(n26559), .Z(n26564) );
  NAND U27261 ( .A(n26562), .B(n26561), .Z(n26563) );
  AND U27262 ( .A(n26564), .B(n26563), .Z(n26612) );
  XOR U27263 ( .A(n26613), .B(n26612), .Z(n26614) );
  NANDN U27264 ( .A(n26566), .B(n26565), .Z(n26570) );
  NANDN U27265 ( .A(n26568), .B(n26567), .Z(n26569) );
  NAND U27266 ( .A(n26570), .B(n26569), .Z(n26615) );
  XOR U27267 ( .A(n26614), .B(n26615), .Z(n26582) );
  OR U27268 ( .A(n26572), .B(n26571), .Z(n26576) );
  NANDN U27269 ( .A(n26574), .B(n26573), .Z(n26575) );
  NAND U27270 ( .A(n26576), .B(n26575), .Z(n26583) );
  XNOR U27271 ( .A(n26582), .B(n26583), .Z(n26584) );
  XNOR U27272 ( .A(n26585), .B(n26584), .Z(n26618) );
  XNOR U27273 ( .A(n26618), .B(sreg[1662]), .Z(n26620) );
  NAND U27274 ( .A(n26577), .B(sreg[1661]), .Z(n26581) );
  OR U27275 ( .A(n26579), .B(n26578), .Z(n26580) );
  AND U27276 ( .A(n26581), .B(n26580), .Z(n26619) );
  XOR U27277 ( .A(n26620), .B(n26619), .Z(c[1662]) );
  NANDN U27278 ( .A(n26583), .B(n26582), .Z(n26587) );
  NAND U27279 ( .A(n26585), .B(n26584), .Z(n26586) );
  NAND U27280 ( .A(n26587), .B(n26586), .Z(n26626) );
  NAND U27281 ( .A(b[0]), .B(a[647]), .Z(n26588) );
  XNOR U27282 ( .A(b[1]), .B(n26588), .Z(n26590) );
  NAND U27283 ( .A(n107), .B(a[646]), .Z(n26589) );
  AND U27284 ( .A(n26590), .B(n26589), .Z(n26643) );
  XOR U27285 ( .A(a[643]), .B(n42197), .Z(n26632) );
  NANDN U27286 ( .A(n26632), .B(n42173), .Z(n26593) );
  NANDN U27287 ( .A(n26591), .B(n42172), .Z(n26592) );
  NAND U27288 ( .A(n26593), .B(n26592), .Z(n26641) );
  NAND U27289 ( .A(b[7]), .B(a[639]), .Z(n26642) );
  XNOR U27290 ( .A(n26641), .B(n26642), .Z(n26644) );
  XOR U27291 ( .A(n26643), .B(n26644), .Z(n26650) );
  NANDN U27292 ( .A(n26594), .B(n42093), .Z(n26596) );
  XOR U27293 ( .A(n42134), .B(a[645]), .Z(n26635) );
  NANDN U27294 ( .A(n26635), .B(n42095), .Z(n26595) );
  NAND U27295 ( .A(n26596), .B(n26595), .Z(n26648) );
  NANDN U27296 ( .A(n26597), .B(n42231), .Z(n26599) );
  XOR U27297 ( .A(n215), .B(a[641]), .Z(n26638) );
  NANDN U27298 ( .A(n26638), .B(n42234), .Z(n26598) );
  AND U27299 ( .A(n26599), .B(n26598), .Z(n26647) );
  XNOR U27300 ( .A(n26648), .B(n26647), .Z(n26649) );
  XNOR U27301 ( .A(n26650), .B(n26649), .Z(n26654) );
  NANDN U27302 ( .A(n26601), .B(n26600), .Z(n26605) );
  NAND U27303 ( .A(n26603), .B(n26602), .Z(n26604) );
  AND U27304 ( .A(n26605), .B(n26604), .Z(n26653) );
  XOR U27305 ( .A(n26654), .B(n26653), .Z(n26655) );
  NANDN U27306 ( .A(n26607), .B(n26606), .Z(n26611) );
  NANDN U27307 ( .A(n26609), .B(n26608), .Z(n26610) );
  NAND U27308 ( .A(n26611), .B(n26610), .Z(n26656) );
  XOR U27309 ( .A(n26655), .B(n26656), .Z(n26623) );
  OR U27310 ( .A(n26613), .B(n26612), .Z(n26617) );
  NANDN U27311 ( .A(n26615), .B(n26614), .Z(n26616) );
  NAND U27312 ( .A(n26617), .B(n26616), .Z(n26624) );
  XNOR U27313 ( .A(n26623), .B(n26624), .Z(n26625) );
  XNOR U27314 ( .A(n26626), .B(n26625), .Z(n26659) );
  XNOR U27315 ( .A(n26659), .B(sreg[1663]), .Z(n26661) );
  NAND U27316 ( .A(n26618), .B(sreg[1662]), .Z(n26622) );
  OR U27317 ( .A(n26620), .B(n26619), .Z(n26621) );
  AND U27318 ( .A(n26622), .B(n26621), .Z(n26660) );
  XOR U27319 ( .A(n26661), .B(n26660), .Z(c[1663]) );
  NANDN U27320 ( .A(n26624), .B(n26623), .Z(n26628) );
  NAND U27321 ( .A(n26626), .B(n26625), .Z(n26627) );
  NAND U27322 ( .A(n26628), .B(n26627), .Z(n26667) );
  NAND U27323 ( .A(b[0]), .B(a[648]), .Z(n26629) );
  XNOR U27324 ( .A(b[1]), .B(n26629), .Z(n26631) );
  NAND U27325 ( .A(n107), .B(a[647]), .Z(n26630) );
  AND U27326 ( .A(n26631), .B(n26630), .Z(n26684) );
  XOR U27327 ( .A(a[644]), .B(n42197), .Z(n26673) );
  NANDN U27328 ( .A(n26673), .B(n42173), .Z(n26634) );
  NANDN U27329 ( .A(n26632), .B(n42172), .Z(n26633) );
  NAND U27330 ( .A(n26634), .B(n26633), .Z(n26682) );
  NAND U27331 ( .A(b[7]), .B(a[640]), .Z(n26683) );
  XNOR U27332 ( .A(n26682), .B(n26683), .Z(n26685) );
  XOR U27333 ( .A(n26684), .B(n26685), .Z(n26691) );
  NANDN U27334 ( .A(n26635), .B(n42093), .Z(n26637) );
  XOR U27335 ( .A(n42134), .B(a[646]), .Z(n26676) );
  NANDN U27336 ( .A(n26676), .B(n42095), .Z(n26636) );
  NAND U27337 ( .A(n26637), .B(n26636), .Z(n26689) );
  NANDN U27338 ( .A(n26638), .B(n42231), .Z(n26640) );
  XOR U27339 ( .A(n215), .B(a[642]), .Z(n26679) );
  NANDN U27340 ( .A(n26679), .B(n42234), .Z(n26639) );
  AND U27341 ( .A(n26640), .B(n26639), .Z(n26688) );
  XNOR U27342 ( .A(n26689), .B(n26688), .Z(n26690) );
  XNOR U27343 ( .A(n26691), .B(n26690), .Z(n26695) );
  NANDN U27344 ( .A(n26642), .B(n26641), .Z(n26646) );
  NAND U27345 ( .A(n26644), .B(n26643), .Z(n26645) );
  AND U27346 ( .A(n26646), .B(n26645), .Z(n26694) );
  XOR U27347 ( .A(n26695), .B(n26694), .Z(n26696) );
  NANDN U27348 ( .A(n26648), .B(n26647), .Z(n26652) );
  NANDN U27349 ( .A(n26650), .B(n26649), .Z(n26651) );
  NAND U27350 ( .A(n26652), .B(n26651), .Z(n26697) );
  XOR U27351 ( .A(n26696), .B(n26697), .Z(n26664) );
  OR U27352 ( .A(n26654), .B(n26653), .Z(n26658) );
  NANDN U27353 ( .A(n26656), .B(n26655), .Z(n26657) );
  NAND U27354 ( .A(n26658), .B(n26657), .Z(n26665) );
  XNOR U27355 ( .A(n26664), .B(n26665), .Z(n26666) );
  XNOR U27356 ( .A(n26667), .B(n26666), .Z(n26700) );
  XNOR U27357 ( .A(n26700), .B(sreg[1664]), .Z(n26702) );
  NAND U27358 ( .A(n26659), .B(sreg[1663]), .Z(n26663) );
  OR U27359 ( .A(n26661), .B(n26660), .Z(n26662) );
  AND U27360 ( .A(n26663), .B(n26662), .Z(n26701) );
  XOR U27361 ( .A(n26702), .B(n26701), .Z(c[1664]) );
  NANDN U27362 ( .A(n26665), .B(n26664), .Z(n26669) );
  NAND U27363 ( .A(n26667), .B(n26666), .Z(n26668) );
  NAND U27364 ( .A(n26669), .B(n26668), .Z(n26708) );
  NAND U27365 ( .A(b[0]), .B(a[649]), .Z(n26670) );
  XNOR U27366 ( .A(b[1]), .B(n26670), .Z(n26672) );
  NAND U27367 ( .A(n107), .B(a[648]), .Z(n26671) );
  AND U27368 ( .A(n26672), .B(n26671), .Z(n26725) );
  XOR U27369 ( .A(a[645]), .B(n42197), .Z(n26714) );
  NANDN U27370 ( .A(n26714), .B(n42173), .Z(n26675) );
  NANDN U27371 ( .A(n26673), .B(n42172), .Z(n26674) );
  NAND U27372 ( .A(n26675), .B(n26674), .Z(n26723) );
  NAND U27373 ( .A(b[7]), .B(a[641]), .Z(n26724) );
  XNOR U27374 ( .A(n26723), .B(n26724), .Z(n26726) );
  XOR U27375 ( .A(n26725), .B(n26726), .Z(n26732) );
  NANDN U27376 ( .A(n26676), .B(n42093), .Z(n26678) );
  XOR U27377 ( .A(n42134), .B(a[647]), .Z(n26717) );
  NANDN U27378 ( .A(n26717), .B(n42095), .Z(n26677) );
  NAND U27379 ( .A(n26678), .B(n26677), .Z(n26730) );
  NANDN U27380 ( .A(n26679), .B(n42231), .Z(n26681) );
  XOR U27381 ( .A(n215), .B(a[643]), .Z(n26720) );
  NANDN U27382 ( .A(n26720), .B(n42234), .Z(n26680) );
  AND U27383 ( .A(n26681), .B(n26680), .Z(n26729) );
  XNOR U27384 ( .A(n26730), .B(n26729), .Z(n26731) );
  XNOR U27385 ( .A(n26732), .B(n26731), .Z(n26736) );
  NANDN U27386 ( .A(n26683), .B(n26682), .Z(n26687) );
  NAND U27387 ( .A(n26685), .B(n26684), .Z(n26686) );
  AND U27388 ( .A(n26687), .B(n26686), .Z(n26735) );
  XOR U27389 ( .A(n26736), .B(n26735), .Z(n26737) );
  NANDN U27390 ( .A(n26689), .B(n26688), .Z(n26693) );
  NANDN U27391 ( .A(n26691), .B(n26690), .Z(n26692) );
  NAND U27392 ( .A(n26693), .B(n26692), .Z(n26738) );
  XOR U27393 ( .A(n26737), .B(n26738), .Z(n26705) );
  OR U27394 ( .A(n26695), .B(n26694), .Z(n26699) );
  NANDN U27395 ( .A(n26697), .B(n26696), .Z(n26698) );
  NAND U27396 ( .A(n26699), .B(n26698), .Z(n26706) );
  XNOR U27397 ( .A(n26705), .B(n26706), .Z(n26707) );
  XNOR U27398 ( .A(n26708), .B(n26707), .Z(n26741) );
  XNOR U27399 ( .A(n26741), .B(sreg[1665]), .Z(n26743) );
  NAND U27400 ( .A(n26700), .B(sreg[1664]), .Z(n26704) );
  OR U27401 ( .A(n26702), .B(n26701), .Z(n26703) );
  AND U27402 ( .A(n26704), .B(n26703), .Z(n26742) );
  XOR U27403 ( .A(n26743), .B(n26742), .Z(c[1665]) );
  NANDN U27404 ( .A(n26706), .B(n26705), .Z(n26710) );
  NAND U27405 ( .A(n26708), .B(n26707), .Z(n26709) );
  NAND U27406 ( .A(n26710), .B(n26709), .Z(n26749) );
  NAND U27407 ( .A(b[0]), .B(a[650]), .Z(n26711) );
  XNOR U27408 ( .A(b[1]), .B(n26711), .Z(n26713) );
  NAND U27409 ( .A(n107), .B(a[649]), .Z(n26712) );
  AND U27410 ( .A(n26713), .B(n26712), .Z(n26766) );
  XOR U27411 ( .A(a[646]), .B(n42197), .Z(n26755) );
  NANDN U27412 ( .A(n26755), .B(n42173), .Z(n26716) );
  NANDN U27413 ( .A(n26714), .B(n42172), .Z(n26715) );
  NAND U27414 ( .A(n26716), .B(n26715), .Z(n26764) );
  NAND U27415 ( .A(b[7]), .B(a[642]), .Z(n26765) );
  XNOR U27416 ( .A(n26764), .B(n26765), .Z(n26767) );
  XOR U27417 ( .A(n26766), .B(n26767), .Z(n26773) );
  NANDN U27418 ( .A(n26717), .B(n42093), .Z(n26719) );
  XOR U27419 ( .A(n42134), .B(a[648]), .Z(n26758) );
  NANDN U27420 ( .A(n26758), .B(n42095), .Z(n26718) );
  NAND U27421 ( .A(n26719), .B(n26718), .Z(n26771) );
  NANDN U27422 ( .A(n26720), .B(n42231), .Z(n26722) );
  XOR U27423 ( .A(n215), .B(a[644]), .Z(n26761) );
  NANDN U27424 ( .A(n26761), .B(n42234), .Z(n26721) );
  AND U27425 ( .A(n26722), .B(n26721), .Z(n26770) );
  XNOR U27426 ( .A(n26771), .B(n26770), .Z(n26772) );
  XNOR U27427 ( .A(n26773), .B(n26772), .Z(n26777) );
  NANDN U27428 ( .A(n26724), .B(n26723), .Z(n26728) );
  NAND U27429 ( .A(n26726), .B(n26725), .Z(n26727) );
  AND U27430 ( .A(n26728), .B(n26727), .Z(n26776) );
  XOR U27431 ( .A(n26777), .B(n26776), .Z(n26778) );
  NANDN U27432 ( .A(n26730), .B(n26729), .Z(n26734) );
  NANDN U27433 ( .A(n26732), .B(n26731), .Z(n26733) );
  NAND U27434 ( .A(n26734), .B(n26733), .Z(n26779) );
  XOR U27435 ( .A(n26778), .B(n26779), .Z(n26746) );
  OR U27436 ( .A(n26736), .B(n26735), .Z(n26740) );
  NANDN U27437 ( .A(n26738), .B(n26737), .Z(n26739) );
  NAND U27438 ( .A(n26740), .B(n26739), .Z(n26747) );
  XNOR U27439 ( .A(n26746), .B(n26747), .Z(n26748) );
  XNOR U27440 ( .A(n26749), .B(n26748), .Z(n26782) );
  XNOR U27441 ( .A(n26782), .B(sreg[1666]), .Z(n26784) );
  NAND U27442 ( .A(n26741), .B(sreg[1665]), .Z(n26745) );
  OR U27443 ( .A(n26743), .B(n26742), .Z(n26744) );
  AND U27444 ( .A(n26745), .B(n26744), .Z(n26783) );
  XOR U27445 ( .A(n26784), .B(n26783), .Z(c[1666]) );
  NANDN U27446 ( .A(n26747), .B(n26746), .Z(n26751) );
  NAND U27447 ( .A(n26749), .B(n26748), .Z(n26750) );
  NAND U27448 ( .A(n26751), .B(n26750), .Z(n26790) );
  NAND U27449 ( .A(b[0]), .B(a[651]), .Z(n26752) );
  XNOR U27450 ( .A(b[1]), .B(n26752), .Z(n26754) );
  NAND U27451 ( .A(n108), .B(a[650]), .Z(n26753) );
  AND U27452 ( .A(n26754), .B(n26753), .Z(n26807) );
  XOR U27453 ( .A(a[647]), .B(n42197), .Z(n26796) );
  NANDN U27454 ( .A(n26796), .B(n42173), .Z(n26757) );
  NANDN U27455 ( .A(n26755), .B(n42172), .Z(n26756) );
  NAND U27456 ( .A(n26757), .B(n26756), .Z(n26805) );
  NAND U27457 ( .A(b[7]), .B(a[643]), .Z(n26806) );
  XNOR U27458 ( .A(n26805), .B(n26806), .Z(n26808) );
  XOR U27459 ( .A(n26807), .B(n26808), .Z(n26814) );
  NANDN U27460 ( .A(n26758), .B(n42093), .Z(n26760) );
  XOR U27461 ( .A(n42134), .B(a[649]), .Z(n26799) );
  NANDN U27462 ( .A(n26799), .B(n42095), .Z(n26759) );
  NAND U27463 ( .A(n26760), .B(n26759), .Z(n26812) );
  NANDN U27464 ( .A(n26761), .B(n42231), .Z(n26763) );
  XOR U27465 ( .A(n215), .B(a[645]), .Z(n26802) );
  NANDN U27466 ( .A(n26802), .B(n42234), .Z(n26762) );
  AND U27467 ( .A(n26763), .B(n26762), .Z(n26811) );
  XNOR U27468 ( .A(n26812), .B(n26811), .Z(n26813) );
  XNOR U27469 ( .A(n26814), .B(n26813), .Z(n26818) );
  NANDN U27470 ( .A(n26765), .B(n26764), .Z(n26769) );
  NAND U27471 ( .A(n26767), .B(n26766), .Z(n26768) );
  AND U27472 ( .A(n26769), .B(n26768), .Z(n26817) );
  XOR U27473 ( .A(n26818), .B(n26817), .Z(n26819) );
  NANDN U27474 ( .A(n26771), .B(n26770), .Z(n26775) );
  NANDN U27475 ( .A(n26773), .B(n26772), .Z(n26774) );
  NAND U27476 ( .A(n26775), .B(n26774), .Z(n26820) );
  XOR U27477 ( .A(n26819), .B(n26820), .Z(n26787) );
  OR U27478 ( .A(n26777), .B(n26776), .Z(n26781) );
  NANDN U27479 ( .A(n26779), .B(n26778), .Z(n26780) );
  NAND U27480 ( .A(n26781), .B(n26780), .Z(n26788) );
  XNOR U27481 ( .A(n26787), .B(n26788), .Z(n26789) );
  XNOR U27482 ( .A(n26790), .B(n26789), .Z(n26823) );
  XNOR U27483 ( .A(n26823), .B(sreg[1667]), .Z(n26825) );
  NAND U27484 ( .A(n26782), .B(sreg[1666]), .Z(n26786) );
  OR U27485 ( .A(n26784), .B(n26783), .Z(n26785) );
  AND U27486 ( .A(n26786), .B(n26785), .Z(n26824) );
  XOR U27487 ( .A(n26825), .B(n26824), .Z(c[1667]) );
  NANDN U27488 ( .A(n26788), .B(n26787), .Z(n26792) );
  NAND U27489 ( .A(n26790), .B(n26789), .Z(n26791) );
  NAND U27490 ( .A(n26792), .B(n26791), .Z(n26831) );
  NAND U27491 ( .A(b[0]), .B(a[652]), .Z(n26793) );
  XNOR U27492 ( .A(b[1]), .B(n26793), .Z(n26795) );
  NAND U27493 ( .A(n108), .B(a[651]), .Z(n26794) );
  AND U27494 ( .A(n26795), .B(n26794), .Z(n26848) );
  XOR U27495 ( .A(a[648]), .B(n42197), .Z(n26837) );
  NANDN U27496 ( .A(n26837), .B(n42173), .Z(n26798) );
  NANDN U27497 ( .A(n26796), .B(n42172), .Z(n26797) );
  NAND U27498 ( .A(n26798), .B(n26797), .Z(n26846) );
  NAND U27499 ( .A(b[7]), .B(a[644]), .Z(n26847) );
  XNOR U27500 ( .A(n26846), .B(n26847), .Z(n26849) );
  XOR U27501 ( .A(n26848), .B(n26849), .Z(n26855) );
  NANDN U27502 ( .A(n26799), .B(n42093), .Z(n26801) );
  XOR U27503 ( .A(n42134), .B(a[650]), .Z(n26840) );
  NANDN U27504 ( .A(n26840), .B(n42095), .Z(n26800) );
  NAND U27505 ( .A(n26801), .B(n26800), .Z(n26853) );
  NANDN U27506 ( .A(n26802), .B(n42231), .Z(n26804) );
  XOR U27507 ( .A(n215), .B(a[646]), .Z(n26843) );
  NANDN U27508 ( .A(n26843), .B(n42234), .Z(n26803) );
  AND U27509 ( .A(n26804), .B(n26803), .Z(n26852) );
  XNOR U27510 ( .A(n26853), .B(n26852), .Z(n26854) );
  XNOR U27511 ( .A(n26855), .B(n26854), .Z(n26859) );
  NANDN U27512 ( .A(n26806), .B(n26805), .Z(n26810) );
  NAND U27513 ( .A(n26808), .B(n26807), .Z(n26809) );
  AND U27514 ( .A(n26810), .B(n26809), .Z(n26858) );
  XOR U27515 ( .A(n26859), .B(n26858), .Z(n26860) );
  NANDN U27516 ( .A(n26812), .B(n26811), .Z(n26816) );
  NANDN U27517 ( .A(n26814), .B(n26813), .Z(n26815) );
  NAND U27518 ( .A(n26816), .B(n26815), .Z(n26861) );
  XOR U27519 ( .A(n26860), .B(n26861), .Z(n26828) );
  OR U27520 ( .A(n26818), .B(n26817), .Z(n26822) );
  NANDN U27521 ( .A(n26820), .B(n26819), .Z(n26821) );
  NAND U27522 ( .A(n26822), .B(n26821), .Z(n26829) );
  XNOR U27523 ( .A(n26828), .B(n26829), .Z(n26830) );
  XNOR U27524 ( .A(n26831), .B(n26830), .Z(n26864) );
  XNOR U27525 ( .A(n26864), .B(sreg[1668]), .Z(n26866) );
  NAND U27526 ( .A(n26823), .B(sreg[1667]), .Z(n26827) );
  OR U27527 ( .A(n26825), .B(n26824), .Z(n26826) );
  AND U27528 ( .A(n26827), .B(n26826), .Z(n26865) );
  XOR U27529 ( .A(n26866), .B(n26865), .Z(c[1668]) );
  NANDN U27530 ( .A(n26829), .B(n26828), .Z(n26833) );
  NAND U27531 ( .A(n26831), .B(n26830), .Z(n26832) );
  NAND U27532 ( .A(n26833), .B(n26832), .Z(n26872) );
  NAND U27533 ( .A(b[0]), .B(a[653]), .Z(n26834) );
  XNOR U27534 ( .A(b[1]), .B(n26834), .Z(n26836) );
  NAND U27535 ( .A(n108), .B(a[652]), .Z(n26835) );
  AND U27536 ( .A(n26836), .B(n26835), .Z(n26889) );
  XOR U27537 ( .A(a[649]), .B(n42197), .Z(n26878) );
  NANDN U27538 ( .A(n26878), .B(n42173), .Z(n26839) );
  NANDN U27539 ( .A(n26837), .B(n42172), .Z(n26838) );
  NAND U27540 ( .A(n26839), .B(n26838), .Z(n26887) );
  NAND U27541 ( .A(b[7]), .B(a[645]), .Z(n26888) );
  XNOR U27542 ( .A(n26887), .B(n26888), .Z(n26890) );
  XOR U27543 ( .A(n26889), .B(n26890), .Z(n26896) );
  NANDN U27544 ( .A(n26840), .B(n42093), .Z(n26842) );
  XOR U27545 ( .A(n42134), .B(a[651]), .Z(n26881) );
  NANDN U27546 ( .A(n26881), .B(n42095), .Z(n26841) );
  NAND U27547 ( .A(n26842), .B(n26841), .Z(n26894) );
  NANDN U27548 ( .A(n26843), .B(n42231), .Z(n26845) );
  XOR U27549 ( .A(n216), .B(a[647]), .Z(n26884) );
  NANDN U27550 ( .A(n26884), .B(n42234), .Z(n26844) );
  AND U27551 ( .A(n26845), .B(n26844), .Z(n26893) );
  XNOR U27552 ( .A(n26894), .B(n26893), .Z(n26895) );
  XNOR U27553 ( .A(n26896), .B(n26895), .Z(n26900) );
  NANDN U27554 ( .A(n26847), .B(n26846), .Z(n26851) );
  NAND U27555 ( .A(n26849), .B(n26848), .Z(n26850) );
  AND U27556 ( .A(n26851), .B(n26850), .Z(n26899) );
  XOR U27557 ( .A(n26900), .B(n26899), .Z(n26901) );
  NANDN U27558 ( .A(n26853), .B(n26852), .Z(n26857) );
  NANDN U27559 ( .A(n26855), .B(n26854), .Z(n26856) );
  NAND U27560 ( .A(n26857), .B(n26856), .Z(n26902) );
  XOR U27561 ( .A(n26901), .B(n26902), .Z(n26869) );
  OR U27562 ( .A(n26859), .B(n26858), .Z(n26863) );
  NANDN U27563 ( .A(n26861), .B(n26860), .Z(n26862) );
  NAND U27564 ( .A(n26863), .B(n26862), .Z(n26870) );
  XNOR U27565 ( .A(n26869), .B(n26870), .Z(n26871) );
  XNOR U27566 ( .A(n26872), .B(n26871), .Z(n26905) );
  XNOR U27567 ( .A(n26905), .B(sreg[1669]), .Z(n26907) );
  NAND U27568 ( .A(n26864), .B(sreg[1668]), .Z(n26868) );
  OR U27569 ( .A(n26866), .B(n26865), .Z(n26867) );
  AND U27570 ( .A(n26868), .B(n26867), .Z(n26906) );
  XOR U27571 ( .A(n26907), .B(n26906), .Z(c[1669]) );
  NANDN U27572 ( .A(n26870), .B(n26869), .Z(n26874) );
  NAND U27573 ( .A(n26872), .B(n26871), .Z(n26873) );
  NAND U27574 ( .A(n26874), .B(n26873), .Z(n26913) );
  NAND U27575 ( .A(b[0]), .B(a[654]), .Z(n26875) );
  XNOR U27576 ( .A(b[1]), .B(n26875), .Z(n26877) );
  NAND U27577 ( .A(n108), .B(a[653]), .Z(n26876) );
  AND U27578 ( .A(n26877), .B(n26876), .Z(n26930) );
  XOR U27579 ( .A(a[650]), .B(n42197), .Z(n26919) );
  NANDN U27580 ( .A(n26919), .B(n42173), .Z(n26880) );
  NANDN U27581 ( .A(n26878), .B(n42172), .Z(n26879) );
  NAND U27582 ( .A(n26880), .B(n26879), .Z(n26928) );
  NAND U27583 ( .A(b[7]), .B(a[646]), .Z(n26929) );
  XNOR U27584 ( .A(n26928), .B(n26929), .Z(n26931) );
  XOR U27585 ( .A(n26930), .B(n26931), .Z(n26937) );
  NANDN U27586 ( .A(n26881), .B(n42093), .Z(n26883) );
  XOR U27587 ( .A(n42134), .B(a[652]), .Z(n26922) );
  NANDN U27588 ( .A(n26922), .B(n42095), .Z(n26882) );
  NAND U27589 ( .A(n26883), .B(n26882), .Z(n26935) );
  NANDN U27590 ( .A(n26884), .B(n42231), .Z(n26886) );
  XOR U27591 ( .A(n216), .B(a[648]), .Z(n26925) );
  NANDN U27592 ( .A(n26925), .B(n42234), .Z(n26885) );
  AND U27593 ( .A(n26886), .B(n26885), .Z(n26934) );
  XNOR U27594 ( .A(n26935), .B(n26934), .Z(n26936) );
  XNOR U27595 ( .A(n26937), .B(n26936), .Z(n26941) );
  NANDN U27596 ( .A(n26888), .B(n26887), .Z(n26892) );
  NAND U27597 ( .A(n26890), .B(n26889), .Z(n26891) );
  AND U27598 ( .A(n26892), .B(n26891), .Z(n26940) );
  XOR U27599 ( .A(n26941), .B(n26940), .Z(n26942) );
  NANDN U27600 ( .A(n26894), .B(n26893), .Z(n26898) );
  NANDN U27601 ( .A(n26896), .B(n26895), .Z(n26897) );
  NAND U27602 ( .A(n26898), .B(n26897), .Z(n26943) );
  XOR U27603 ( .A(n26942), .B(n26943), .Z(n26910) );
  OR U27604 ( .A(n26900), .B(n26899), .Z(n26904) );
  NANDN U27605 ( .A(n26902), .B(n26901), .Z(n26903) );
  NAND U27606 ( .A(n26904), .B(n26903), .Z(n26911) );
  XNOR U27607 ( .A(n26910), .B(n26911), .Z(n26912) );
  XNOR U27608 ( .A(n26913), .B(n26912), .Z(n26946) );
  XNOR U27609 ( .A(n26946), .B(sreg[1670]), .Z(n26948) );
  NAND U27610 ( .A(n26905), .B(sreg[1669]), .Z(n26909) );
  OR U27611 ( .A(n26907), .B(n26906), .Z(n26908) );
  AND U27612 ( .A(n26909), .B(n26908), .Z(n26947) );
  XOR U27613 ( .A(n26948), .B(n26947), .Z(c[1670]) );
  NANDN U27614 ( .A(n26911), .B(n26910), .Z(n26915) );
  NAND U27615 ( .A(n26913), .B(n26912), .Z(n26914) );
  NAND U27616 ( .A(n26915), .B(n26914), .Z(n26954) );
  NAND U27617 ( .A(b[0]), .B(a[655]), .Z(n26916) );
  XNOR U27618 ( .A(b[1]), .B(n26916), .Z(n26918) );
  NAND U27619 ( .A(n108), .B(a[654]), .Z(n26917) );
  AND U27620 ( .A(n26918), .B(n26917), .Z(n26971) );
  XOR U27621 ( .A(a[651]), .B(n42197), .Z(n26960) );
  NANDN U27622 ( .A(n26960), .B(n42173), .Z(n26921) );
  NANDN U27623 ( .A(n26919), .B(n42172), .Z(n26920) );
  NAND U27624 ( .A(n26921), .B(n26920), .Z(n26969) );
  NAND U27625 ( .A(b[7]), .B(a[647]), .Z(n26970) );
  XNOR U27626 ( .A(n26969), .B(n26970), .Z(n26972) );
  XOR U27627 ( .A(n26971), .B(n26972), .Z(n26978) );
  NANDN U27628 ( .A(n26922), .B(n42093), .Z(n26924) );
  XOR U27629 ( .A(n42134), .B(a[653]), .Z(n26963) );
  NANDN U27630 ( .A(n26963), .B(n42095), .Z(n26923) );
  NAND U27631 ( .A(n26924), .B(n26923), .Z(n26976) );
  NANDN U27632 ( .A(n26925), .B(n42231), .Z(n26927) );
  XOR U27633 ( .A(n216), .B(a[649]), .Z(n26966) );
  NANDN U27634 ( .A(n26966), .B(n42234), .Z(n26926) );
  AND U27635 ( .A(n26927), .B(n26926), .Z(n26975) );
  XNOR U27636 ( .A(n26976), .B(n26975), .Z(n26977) );
  XNOR U27637 ( .A(n26978), .B(n26977), .Z(n26982) );
  NANDN U27638 ( .A(n26929), .B(n26928), .Z(n26933) );
  NAND U27639 ( .A(n26931), .B(n26930), .Z(n26932) );
  AND U27640 ( .A(n26933), .B(n26932), .Z(n26981) );
  XOR U27641 ( .A(n26982), .B(n26981), .Z(n26983) );
  NANDN U27642 ( .A(n26935), .B(n26934), .Z(n26939) );
  NANDN U27643 ( .A(n26937), .B(n26936), .Z(n26938) );
  NAND U27644 ( .A(n26939), .B(n26938), .Z(n26984) );
  XOR U27645 ( .A(n26983), .B(n26984), .Z(n26951) );
  OR U27646 ( .A(n26941), .B(n26940), .Z(n26945) );
  NANDN U27647 ( .A(n26943), .B(n26942), .Z(n26944) );
  NAND U27648 ( .A(n26945), .B(n26944), .Z(n26952) );
  XNOR U27649 ( .A(n26951), .B(n26952), .Z(n26953) );
  XNOR U27650 ( .A(n26954), .B(n26953), .Z(n26987) );
  XNOR U27651 ( .A(n26987), .B(sreg[1671]), .Z(n26989) );
  NAND U27652 ( .A(n26946), .B(sreg[1670]), .Z(n26950) );
  OR U27653 ( .A(n26948), .B(n26947), .Z(n26949) );
  AND U27654 ( .A(n26950), .B(n26949), .Z(n26988) );
  XOR U27655 ( .A(n26989), .B(n26988), .Z(c[1671]) );
  NANDN U27656 ( .A(n26952), .B(n26951), .Z(n26956) );
  NAND U27657 ( .A(n26954), .B(n26953), .Z(n26955) );
  NAND U27658 ( .A(n26956), .B(n26955), .Z(n26995) );
  NAND U27659 ( .A(b[0]), .B(a[656]), .Z(n26957) );
  XNOR U27660 ( .A(b[1]), .B(n26957), .Z(n26959) );
  NAND U27661 ( .A(n108), .B(a[655]), .Z(n26958) );
  AND U27662 ( .A(n26959), .B(n26958), .Z(n27012) );
  XOR U27663 ( .A(a[652]), .B(n42197), .Z(n27001) );
  NANDN U27664 ( .A(n27001), .B(n42173), .Z(n26962) );
  NANDN U27665 ( .A(n26960), .B(n42172), .Z(n26961) );
  NAND U27666 ( .A(n26962), .B(n26961), .Z(n27010) );
  NAND U27667 ( .A(b[7]), .B(a[648]), .Z(n27011) );
  XNOR U27668 ( .A(n27010), .B(n27011), .Z(n27013) );
  XOR U27669 ( .A(n27012), .B(n27013), .Z(n27019) );
  NANDN U27670 ( .A(n26963), .B(n42093), .Z(n26965) );
  XOR U27671 ( .A(n42134), .B(a[654]), .Z(n27004) );
  NANDN U27672 ( .A(n27004), .B(n42095), .Z(n26964) );
  NAND U27673 ( .A(n26965), .B(n26964), .Z(n27017) );
  NANDN U27674 ( .A(n26966), .B(n42231), .Z(n26968) );
  XOR U27675 ( .A(n216), .B(a[650]), .Z(n27007) );
  NANDN U27676 ( .A(n27007), .B(n42234), .Z(n26967) );
  AND U27677 ( .A(n26968), .B(n26967), .Z(n27016) );
  XNOR U27678 ( .A(n27017), .B(n27016), .Z(n27018) );
  XNOR U27679 ( .A(n27019), .B(n27018), .Z(n27023) );
  NANDN U27680 ( .A(n26970), .B(n26969), .Z(n26974) );
  NAND U27681 ( .A(n26972), .B(n26971), .Z(n26973) );
  AND U27682 ( .A(n26974), .B(n26973), .Z(n27022) );
  XOR U27683 ( .A(n27023), .B(n27022), .Z(n27024) );
  NANDN U27684 ( .A(n26976), .B(n26975), .Z(n26980) );
  NANDN U27685 ( .A(n26978), .B(n26977), .Z(n26979) );
  NAND U27686 ( .A(n26980), .B(n26979), .Z(n27025) );
  XOR U27687 ( .A(n27024), .B(n27025), .Z(n26992) );
  OR U27688 ( .A(n26982), .B(n26981), .Z(n26986) );
  NANDN U27689 ( .A(n26984), .B(n26983), .Z(n26985) );
  NAND U27690 ( .A(n26986), .B(n26985), .Z(n26993) );
  XNOR U27691 ( .A(n26992), .B(n26993), .Z(n26994) );
  XNOR U27692 ( .A(n26995), .B(n26994), .Z(n27028) );
  XNOR U27693 ( .A(n27028), .B(sreg[1672]), .Z(n27030) );
  NAND U27694 ( .A(n26987), .B(sreg[1671]), .Z(n26991) );
  OR U27695 ( .A(n26989), .B(n26988), .Z(n26990) );
  AND U27696 ( .A(n26991), .B(n26990), .Z(n27029) );
  XOR U27697 ( .A(n27030), .B(n27029), .Z(c[1672]) );
  NANDN U27698 ( .A(n26993), .B(n26992), .Z(n26997) );
  NAND U27699 ( .A(n26995), .B(n26994), .Z(n26996) );
  NAND U27700 ( .A(n26997), .B(n26996), .Z(n27036) );
  NAND U27701 ( .A(b[0]), .B(a[657]), .Z(n26998) );
  XNOR U27702 ( .A(b[1]), .B(n26998), .Z(n27000) );
  NAND U27703 ( .A(n108), .B(a[656]), .Z(n26999) );
  AND U27704 ( .A(n27000), .B(n26999), .Z(n27053) );
  XOR U27705 ( .A(a[653]), .B(n42197), .Z(n27042) );
  NANDN U27706 ( .A(n27042), .B(n42173), .Z(n27003) );
  NANDN U27707 ( .A(n27001), .B(n42172), .Z(n27002) );
  NAND U27708 ( .A(n27003), .B(n27002), .Z(n27051) );
  NAND U27709 ( .A(b[7]), .B(a[649]), .Z(n27052) );
  XNOR U27710 ( .A(n27051), .B(n27052), .Z(n27054) );
  XOR U27711 ( .A(n27053), .B(n27054), .Z(n27060) );
  NANDN U27712 ( .A(n27004), .B(n42093), .Z(n27006) );
  XOR U27713 ( .A(n42134), .B(a[655]), .Z(n27045) );
  NANDN U27714 ( .A(n27045), .B(n42095), .Z(n27005) );
  NAND U27715 ( .A(n27006), .B(n27005), .Z(n27058) );
  NANDN U27716 ( .A(n27007), .B(n42231), .Z(n27009) );
  XOR U27717 ( .A(n216), .B(a[651]), .Z(n27048) );
  NANDN U27718 ( .A(n27048), .B(n42234), .Z(n27008) );
  AND U27719 ( .A(n27009), .B(n27008), .Z(n27057) );
  XNOR U27720 ( .A(n27058), .B(n27057), .Z(n27059) );
  XNOR U27721 ( .A(n27060), .B(n27059), .Z(n27064) );
  NANDN U27722 ( .A(n27011), .B(n27010), .Z(n27015) );
  NAND U27723 ( .A(n27013), .B(n27012), .Z(n27014) );
  AND U27724 ( .A(n27015), .B(n27014), .Z(n27063) );
  XOR U27725 ( .A(n27064), .B(n27063), .Z(n27065) );
  NANDN U27726 ( .A(n27017), .B(n27016), .Z(n27021) );
  NANDN U27727 ( .A(n27019), .B(n27018), .Z(n27020) );
  NAND U27728 ( .A(n27021), .B(n27020), .Z(n27066) );
  XOR U27729 ( .A(n27065), .B(n27066), .Z(n27033) );
  OR U27730 ( .A(n27023), .B(n27022), .Z(n27027) );
  NANDN U27731 ( .A(n27025), .B(n27024), .Z(n27026) );
  NAND U27732 ( .A(n27027), .B(n27026), .Z(n27034) );
  XNOR U27733 ( .A(n27033), .B(n27034), .Z(n27035) );
  XNOR U27734 ( .A(n27036), .B(n27035), .Z(n27069) );
  XNOR U27735 ( .A(n27069), .B(sreg[1673]), .Z(n27071) );
  NAND U27736 ( .A(n27028), .B(sreg[1672]), .Z(n27032) );
  OR U27737 ( .A(n27030), .B(n27029), .Z(n27031) );
  AND U27738 ( .A(n27032), .B(n27031), .Z(n27070) );
  XOR U27739 ( .A(n27071), .B(n27070), .Z(c[1673]) );
  NANDN U27740 ( .A(n27034), .B(n27033), .Z(n27038) );
  NAND U27741 ( .A(n27036), .B(n27035), .Z(n27037) );
  NAND U27742 ( .A(n27038), .B(n27037), .Z(n27077) );
  NAND U27743 ( .A(b[0]), .B(a[658]), .Z(n27039) );
  XNOR U27744 ( .A(b[1]), .B(n27039), .Z(n27041) );
  NAND U27745 ( .A(n109), .B(a[657]), .Z(n27040) );
  AND U27746 ( .A(n27041), .B(n27040), .Z(n27094) );
  XOR U27747 ( .A(a[654]), .B(n42197), .Z(n27083) );
  NANDN U27748 ( .A(n27083), .B(n42173), .Z(n27044) );
  NANDN U27749 ( .A(n27042), .B(n42172), .Z(n27043) );
  NAND U27750 ( .A(n27044), .B(n27043), .Z(n27092) );
  NAND U27751 ( .A(b[7]), .B(a[650]), .Z(n27093) );
  XNOR U27752 ( .A(n27092), .B(n27093), .Z(n27095) );
  XOR U27753 ( .A(n27094), .B(n27095), .Z(n27101) );
  NANDN U27754 ( .A(n27045), .B(n42093), .Z(n27047) );
  XOR U27755 ( .A(n42134), .B(a[656]), .Z(n27086) );
  NANDN U27756 ( .A(n27086), .B(n42095), .Z(n27046) );
  NAND U27757 ( .A(n27047), .B(n27046), .Z(n27099) );
  NANDN U27758 ( .A(n27048), .B(n42231), .Z(n27050) );
  XOR U27759 ( .A(n216), .B(a[652]), .Z(n27089) );
  NANDN U27760 ( .A(n27089), .B(n42234), .Z(n27049) );
  AND U27761 ( .A(n27050), .B(n27049), .Z(n27098) );
  XNOR U27762 ( .A(n27099), .B(n27098), .Z(n27100) );
  XNOR U27763 ( .A(n27101), .B(n27100), .Z(n27105) );
  NANDN U27764 ( .A(n27052), .B(n27051), .Z(n27056) );
  NAND U27765 ( .A(n27054), .B(n27053), .Z(n27055) );
  AND U27766 ( .A(n27056), .B(n27055), .Z(n27104) );
  XOR U27767 ( .A(n27105), .B(n27104), .Z(n27106) );
  NANDN U27768 ( .A(n27058), .B(n27057), .Z(n27062) );
  NANDN U27769 ( .A(n27060), .B(n27059), .Z(n27061) );
  NAND U27770 ( .A(n27062), .B(n27061), .Z(n27107) );
  XOR U27771 ( .A(n27106), .B(n27107), .Z(n27074) );
  OR U27772 ( .A(n27064), .B(n27063), .Z(n27068) );
  NANDN U27773 ( .A(n27066), .B(n27065), .Z(n27067) );
  NAND U27774 ( .A(n27068), .B(n27067), .Z(n27075) );
  XNOR U27775 ( .A(n27074), .B(n27075), .Z(n27076) );
  XNOR U27776 ( .A(n27077), .B(n27076), .Z(n27110) );
  XNOR U27777 ( .A(n27110), .B(sreg[1674]), .Z(n27112) );
  NAND U27778 ( .A(n27069), .B(sreg[1673]), .Z(n27073) );
  OR U27779 ( .A(n27071), .B(n27070), .Z(n27072) );
  AND U27780 ( .A(n27073), .B(n27072), .Z(n27111) );
  XOR U27781 ( .A(n27112), .B(n27111), .Z(c[1674]) );
  NANDN U27782 ( .A(n27075), .B(n27074), .Z(n27079) );
  NAND U27783 ( .A(n27077), .B(n27076), .Z(n27078) );
  NAND U27784 ( .A(n27079), .B(n27078), .Z(n27118) );
  NAND U27785 ( .A(b[0]), .B(a[659]), .Z(n27080) );
  XNOR U27786 ( .A(b[1]), .B(n27080), .Z(n27082) );
  NAND U27787 ( .A(n109), .B(a[658]), .Z(n27081) );
  AND U27788 ( .A(n27082), .B(n27081), .Z(n27135) );
  XOR U27789 ( .A(a[655]), .B(n42197), .Z(n27124) );
  NANDN U27790 ( .A(n27124), .B(n42173), .Z(n27085) );
  NANDN U27791 ( .A(n27083), .B(n42172), .Z(n27084) );
  NAND U27792 ( .A(n27085), .B(n27084), .Z(n27133) );
  NAND U27793 ( .A(b[7]), .B(a[651]), .Z(n27134) );
  XNOR U27794 ( .A(n27133), .B(n27134), .Z(n27136) );
  XOR U27795 ( .A(n27135), .B(n27136), .Z(n27142) );
  NANDN U27796 ( .A(n27086), .B(n42093), .Z(n27088) );
  XOR U27797 ( .A(n42134), .B(a[657]), .Z(n27127) );
  NANDN U27798 ( .A(n27127), .B(n42095), .Z(n27087) );
  NAND U27799 ( .A(n27088), .B(n27087), .Z(n27140) );
  NANDN U27800 ( .A(n27089), .B(n42231), .Z(n27091) );
  XOR U27801 ( .A(n216), .B(a[653]), .Z(n27130) );
  NANDN U27802 ( .A(n27130), .B(n42234), .Z(n27090) );
  AND U27803 ( .A(n27091), .B(n27090), .Z(n27139) );
  XNOR U27804 ( .A(n27140), .B(n27139), .Z(n27141) );
  XNOR U27805 ( .A(n27142), .B(n27141), .Z(n27146) );
  NANDN U27806 ( .A(n27093), .B(n27092), .Z(n27097) );
  NAND U27807 ( .A(n27095), .B(n27094), .Z(n27096) );
  AND U27808 ( .A(n27097), .B(n27096), .Z(n27145) );
  XOR U27809 ( .A(n27146), .B(n27145), .Z(n27147) );
  NANDN U27810 ( .A(n27099), .B(n27098), .Z(n27103) );
  NANDN U27811 ( .A(n27101), .B(n27100), .Z(n27102) );
  NAND U27812 ( .A(n27103), .B(n27102), .Z(n27148) );
  XOR U27813 ( .A(n27147), .B(n27148), .Z(n27115) );
  OR U27814 ( .A(n27105), .B(n27104), .Z(n27109) );
  NANDN U27815 ( .A(n27107), .B(n27106), .Z(n27108) );
  NAND U27816 ( .A(n27109), .B(n27108), .Z(n27116) );
  XNOR U27817 ( .A(n27115), .B(n27116), .Z(n27117) );
  XNOR U27818 ( .A(n27118), .B(n27117), .Z(n27151) );
  XNOR U27819 ( .A(n27151), .B(sreg[1675]), .Z(n27153) );
  NAND U27820 ( .A(n27110), .B(sreg[1674]), .Z(n27114) );
  OR U27821 ( .A(n27112), .B(n27111), .Z(n27113) );
  AND U27822 ( .A(n27114), .B(n27113), .Z(n27152) );
  XOR U27823 ( .A(n27153), .B(n27152), .Z(c[1675]) );
  NANDN U27824 ( .A(n27116), .B(n27115), .Z(n27120) );
  NAND U27825 ( .A(n27118), .B(n27117), .Z(n27119) );
  NAND U27826 ( .A(n27120), .B(n27119), .Z(n27159) );
  NAND U27827 ( .A(b[0]), .B(a[660]), .Z(n27121) );
  XNOR U27828 ( .A(b[1]), .B(n27121), .Z(n27123) );
  NAND U27829 ( .A(n109), .B(a[659]), .Z(n27122) );
  AND U27830 ( .A(n27123), .B(n27122), .Z(n27176) );
  XOR U27831 ( .A(a[656]), .B(n42197), .Z(n27165) );
  NANDN U27832 ( .A(n27165), .B(n42173), .Z(n27126) );
  NANDN U27833 ( .A(n27124), .B(n42172), .Z(n27125) );
  NAND U27834 ( .A(n27126), .B(n27125), .Z(n27174) );
  NAND U27835 ( .A(b[7]), .B(a[652]), .Z(n27175) );
  XNOR U27836 ( .A(n27174), .B(n27175), .Z(n27177) );
  XOR U27837 ( .A(n27176), .B(n27177), .Z(n27183) );
  NANDN U27838 ( .A(n27127), .B(n42093), .Z(n27129) );
  XOR U27839 ( .A(n42134), .B(a[658]), .Z(n27168) );
  NANDN U27840 ( .A(n27168), .B(n42095), .Z(n27128) );
  NAND U27841 ( .A(n27129), .B(n27128), .Z(n27181) );
  NANDN U27842 ( .A(n27130), .B(n42231), .Z(n27132) );
  XOR U27843 ( .A(n216), .B(a[654]), .Z(n27171) );
  NANDN U27844 ( .A(n27171), .B(n42234), .Z(n27131) );
  AND U27845 ( .A(n27132), .B(n27131), .Z(n27180) );
  XNOR U27846 ( .A(n27181), .B(n27180), .Z(n27182) );
  XNOR U27847 ( .A(n27183), .B(n27182), .Z(n27187) );
  NANDN U27848 ( .A(n27134), .B(n27133), .Z(n27138) );
  NAND U27849 ( .A(n27136), .B(n27135), .Z(n27137) );
  AND U27850 ( .A(n27138), .B(n27137), .Z(n27186) );
  XOR U27851 ( .A(n27187), .B(n27186), .Z(n27188) );
  NANDN U27852 ( .A(n27140), .B(n27139), .Z(n27144) );
  NANDN U27853 ( .A(n27142), .B(n27141), .Z(n27143) );
  NAND U27854 ( .A(n27144), .B(n27143), .Z(n27189) );
  XOR U27855 ( .A(n27188), .B(n27189), .Z(n27156) );
  OR U27856 ( .A(n27146), .B(n27145), .Z(n27150) );
  NANDN U27857 ( .A(n27148), .B(n27147), .Z(n27149) );
  NAND U27858 ( .A(n27150), .B(n27149), .Z(n27157) );
  XNOR U27859 ( .A(n27156), .B(n27157), .Z(n27158) );
  XNOR U27860 ( .A(n27159), .B(n27158), .Z(n27192) );
  XNOR U27861 ( .A(n27192), .B(sreg[1676]), .Z(n27194) );
  NAND U27862 ( .A(n27151), .B(sreg[1675]), .Z(n27155) );
  OR U27863 ( .A(n27153), .B(n27152), .Z(n27154) );
  AND U27864 ( .A(n27155), .B(n27154), .Z(n27193) );
  XOR U27865 ( .A(n27194), .B(n27193), .Z(c[1676]) );
  NANDN U27866 ( .A(n27157), .B(n27156), .Z(n27161) );
  NAND U27867 ( .A(n27159), .B(n27158), .Z(n27160) );
  NAND U27868 ( .A(n27161), .B(n27160), .Z(n27200) );
  NAND U27869 ( .A(b[0]), .B(a[661]), .Z(n27162) );
  XNOR U27870 ( .A(b[1]), .B(n27162), .Z(n27164) );
  NAND U27871 ( .A(n109), .B(a[660]), .Z(n27163) );
  AND U27872 ( .A(n27164), .B(n27163), .Z(n27217) );
  XOR U27873 ( .A(a[657]), .B(n42197), .Z(n27206) );
  NANDN U27874 ( .A(n27206), .B(n42173), .Z(n27167) );
  NANDN U27875 ( .A(n27165), .B(n42172), .Z(n27166) );
  NAND U27876 ( .A(n27167), .B(n27166), .Z(n27215) );
  NAND U27877 ( .A(b[7]), .B(a[653]), .Z(n27216) );
  XNOR U27878 ( .A(n27215), .B(n27216), .Z(n27218) );
  XOR U27879 ( .A(n27217), .B(n27218), .Z(n27224) );
  NANDN U27880 ( .A(n27168), .B(n42093), .Z(n27170) );
  XOR U27881 ( .A(n42134), .B(a[659]), .Z(n27209) );
  NANDN U27882 ( .A(n27209), .B(n42095), .Z(n27169) );
  NAND U27883 ( .A(n27170), .B(n27169), .Z(n27222) );
  NANDN U27884 ( .A(n27171), .B(n42231), .Z(n27173) );
  XOR U27885 ( .A(n216), .B(a[655]), .Z(n27212) );
  NANDN U27886 ( .A(n27212), .B(n42234), .Z(n27172) );
  AND U27887 ( .A(n27173), .B(n27172), .Z(n27221) );
  XNOR U27888 ( .A(n27222), .B(n27221), .Z(n27223) );
  XNOR U27889 ( .A(n27224), .B(n27223), .Z(n27228) );
  NANDN U27890 ( .A(n27175), .B(n27174), .Z(n27179) );
  NAND U27891 ( .A(n27177), .B(n27176), .Z(n27178) );
  AND U27892 ( .A(n27179), .B(n27178), .Z(n27227) );
  XOR U27893 ( .A(n27228), .B(n27227), .Z(n27229) );
  NANDN U27894 ( .A(n27181), .B(n27180), .Z(n27185) );
  NANDN U27895 ( .A(n27183), .B(n27182), .Z(n27184) );
  NAND U27896 ( .A(n27185), .B(n27184), .Z(n27230) );
  XOR U27897 ( .A(n27229), .B(n27230), .Z(n27197) );
  OR U27898 ( .A(n27187), .B(n27186), .Z(n27191) );
  NANDN U27899 ( .A(n27189), .B(n27188), .Z(n27190) );
  NAND U27900 ( .A(n27191), .B(n27190), .Z(n27198) );
  XNOR U27901 ( .A(n27197), .B(n27198), .Z(n27199) );
  XNOR U27902 ( .A(n27200), .B(n27199), .Z(n27233) );
  XNOR U27903 ( .A(n27233), .B(sreg[1677]), .Z(n27235) );
  NAND U27904 ( .A(n27192), .B(sreg[1676]), .Z(n27196) );
  OR U27905 ( .A(n27194), .B(n27193), .Z(n27195) );
  AND U27906 ( .A(n27196), .B(n27195), .Z(n27234) );
  XOR U27907 ( .A(n27235), .B(n27234), .Z(c[1677]) );
  NANDN U27908 ( .A(n27198), .B(n27197), .Z(n27202) );
  NAND U27909 ( .A(n27200), .B(n27199), .Z(n27201) );
  NAND U27910 ( .A(n27202), .B(n27201), .Z(n27241) );
  NAND U27911 ( .A(b[0]), .B(a[662]), .Z(n27203) );
  XNOR U27912 ( .A(b[1]), .B(n27203), .Z(n27205) );
  NAND U27913 ( .A(n109), .B(a[661]), .Z(n27204) );
  AND U27914 ( .A(n27205), .B(n27204), .Z(n27258) );
  XOR U27915 ( .A(a[658]), .B(n42197), .Z(n27247) );
  NANDN U27916 ( .A(n27247), .B(n42173), .Z(n27208) );
  NANDN U27917 ( .A(n27206), .B(n42172), .Z(n27207) );
  NAND U27918 ( .A(n27208), .B(n27207), .Z(n27256) );
  NAND U27919 ( .A(b[7]), .B(a[654]), .Z(n27257) );
  XNOR U27920 ( .A(n27256), .B(n27257), .Z(n27259) );
  XOR U27921 ( .A(n27258), .B(n27259), .Z(n27265) );
  NANDN U27922 ( .A(n27209), .B(n42093), .Z(n27211) );
  XOR U27923 ( .A(n42134), .B(a[660]), .Z(n27250) );
  NANDN U27924 ( .A(n27250), .B(n42095), .Z(n27210) );
  NAND U27925 ( .A(n27211), .B(n27210), .Z(n27263) );
  NANDN U27926 ( .A(n27212), .B(n42231), .Z(n27214) );
  XOR U27927 ( .A(n216), .B(a[656]), .Z(n27253) );
  NANDN U27928 ( .A(n27253), .B(n42234), .Z(n27213) );
  AND U27929 ( .A(n27214), .B(n27213), .Z(n27262) );
  XNOR U27930 ( .A(n27263), .B(n27262), .Z(n27264) );
  XNOR U27931 ( .A(n27265), .B(n27264), .Z(n27269) );
  NANDN U27932 ( .A(n27216), .B(n27215), .Z(n27220) );
  NAND U27933 ( .A(n27218), .B(n27217), .Z(n27219) );
  AND U27934 ( .A(n27220), .B(n27219), .Z(n27268) );
  XOR U27935 ( .A(n27269), .B(n27268), .Z(n27270) );
  NANDN U27936 ( .A(n27222), .B(n27221), .Z(n27226) );
  NANDN U27937 ( .A(n27224), .B(n27223), .Z(n27225) );
  NAND U27938 ( .A(n27226), .B(n27225), .Z(n27271) );
  XOR U27939 ( .A(n27270), .B(n27271), .Z(n27238) );
  OR U27940 ( .A(n27228), .B(n27227), .Z(n27232) );
  NANDN U27941 ( .A(n27230), .B(n27229), .Z(n27231) );
  NAND U27942 ( .A(n27232), .B(n27231), .Z(n27239) );
  XNOR U27943 ( .A(n27238), .B(n27239), .Z(n27240) );
  XNOR U27944 ( .A(n27241), .B(n27240), .Z(n27274) );
  XNOR U27945 ( .A(n27274), .B(sreg[1678]), .Z(n27276) );
  NAND U27946 ( .A(n27233), .B(sreg[1677]), .Z(n27237) );
  OR U27947 ( .A(n27235), .B(n27234), .Z(n27236) );
  AND U27948 ( .A(n27237), .B(n27236), .Z(n27275) );
  XOR U27949 ( .A(n27276), .B(n27275), .Z(c[1678]) );
  NANDN U27950 ( .A(n27239), .B(n27238), .Z(n27243) );
  NAND U27951 ( .A(n27241), .B(n27240), .Z(n27242) );
  NAND U27952 ( .A(n27243), .B(n27242), .Z(n27282) );
  NAND U27953 ( .A(b[0]), .B(a[663]), .Z(n27244) );
  XNOR U27954 ( .A(b[1]), .B(n27244), .Z(n27246) );
  NAND U27955 ( .A(n109), .B(a[662]), .Z(n27245) );
  AND U27956 ( .A(n27246), .B(n27245), .Z(n27299) );
  XOR U27957 ( .A(a[659]), .B(n42197), .Z(n27288) );
  NANDN U27958 ( .A(n27288), .B(n42173), .Z(n27249) );
  NANDN U27959 ( .A(n27247), .B(n42172), .Z(n27248) );
  NAND U27960 ( .A(n27249), .B(n27248), .Z(n27297) );
  NAND U27961 ( .A(b[7]), .B(a[655]), .Z(n27298) );
  XNOR U27962 ( .A(n27297), .B(n27298), .Z(n27300) );
  XOR U27963 ( .A(n27299), .B(n27300), .Z(n27306) );
  NANDN U27964 ( .A(n27250), .B(n42093), .Z(n27252) );
  XOR U27965 ( .A(n42134), .B(a[661]), .Z(n27291) );
  NANDN U27966 ( .A(n27291), .B(n42095), .Z(n27251) );
  NAND U27967 ( .A(n27252), .B(n27251), .Z(n27304) );
  NANDN U27968 ( .A(n27253), .B(n42231), .Z(n27255) );
  XOR U27969 ( .A(n216), .B(a[657]), .Z(n27294) );
  NANDN U27970 ( .A(n27294), .B(n42234), .Z(n27254) );
  AND U27971 ( .A(n27255), .B(n27254), .Z(n27303) );
  XNOR U27972 ( .A(n27304), .B(n27303), .Z(n27305) );
  XNOR U27973 ( .A(n27306), .B(n27305), .Z(n27310) );
  NANDN U27974 ( .A(n27257), .B(n27256), .Z(n27261) );
  NAND U27975 ( .A(n27259), .B(n27258), .Z(n27260) );
  AND U27976 ( .A(n27261), .B(n27260), .Z(n27309) );
  XOR U27977 ( .A(n27310), .B(n27309), .Z(n27311) );
  NANDN U27978 ( .A(n27263), .B(n27262), .Z(n27267) );
  NANDN U27979 ( .A(n27265), .B(n27264), .Z(n27266) );
  NAND U27980 ( .A(n27267), .B(n27266), .Z(n27312) );
  XOR U27981 ( .A(n27311), .B(n27312), .Z(n27279) );
  OR U27982 ( .A(n27269), .B(n27268), .Z(n27273) );
  NANDN U27983 ( .A(n27271), .B(n27270), .Z(n27272) );
  NAND U27984 ( .A(n27273), .B(n27272), .Z(n27280) );
  XNOR U27985 ( .A(n27279), .B(n27280), .Z(n27281) );
  XNOR U27986 ( .A(n27282), .B(n27281), .Z(n27315) );
  XNOR U27987 ( .A(n27315), .B(sreg[1679]), .Z(n27317) );
  NAND U27988 ( .A(n27274), .B(sreg[1678]), .Z(n27278) );
  OR U27989 ( .A(n27276), .B(n27275), .Z(n27277) );
  AND U27990 ( .A(n27278), .B(n27277), .Z(n27316) );
  XOR U27991 ( .A(n27317), .B(n27316), .Z(c[1679]) );
  NANDN U27992 ( .A(n27280), .B(n27279), .Z(n27284) );
  NAND U27993 ( .A(n27282), .B(n27281), .Z(n27283) );
  NAND U27994 ( .A(n27284), .B(n27283), .Z(n27323) );
  NAND U27995 ( .A(b[0]), .B(a[664]), .Z(n27285) );
  XNOR U27996 ( .A(b[1]), .B(n27285), .Z(n27287) );
  NAND U27997 ( .A(n109), .B(a[663]), .Z(n27286) );
  AND U27998 ( .A(n27287), .B(n27286), .Z(n27340) );
  XOR U27999 ( .A(a[660]), .B(n42197), .Z(n27329) );
  NANDN U28000 ( .A(n27329), .B(n42173), .Z(n27290) );
  NANDN U28001 ( .A(n27288), .B(n42172), .Z(n27289) );
  NAND U28002 ( .A(n27290), .B(n27289), .Z(n27338) );
  NAND U28003 ( .A(b[7]), .B(a[656]), .Z(n27339) );
  XNOR U28004 ( .A(n27338), .B(n27339), .Z(n27341) );
  XOR U28005 ( .A(n27340), .B(n27341), .Z(n27347) );
  NANDN U28006 ( .A(n27291), .B(n42093), .Z(n27293) );
  XOR U28007 ( .A(n42134), .B(a[662]), .Z(n27332) );
  NANDN U28008 ( .A(n27332), .B(n42095), .Z(n27292) );
  NAND U28009 ( .A(n27293), .B(n27292), .Z(n27345) );
  NANDN U28010 ( .A(n27294), .B(n42231), .Z(n27296) );
  XOR U28011 ( .A(n216), .B(a[658]), .Z(n27335) );
  NANDN U28012 ( .A(n27335), .B(n42234), .Z(n27295) );
  AND U28013 ( .A(n27296), .B(n27295), .Z(n27344) );
  XNOR U28014 ( .A(n27345), .B(n27344), .Z(n27346) );
  XNOR U28015 ( .A(n27347), .B(n27346), .Z(n27351) );
  NANDN U28016 ( .A(n27298), .B(n27297), .Z(n27302) );
  NAND U28017 ( .A(n27300), .B(n27299), .Z(n27301) );
  AND U28018 ( .A(n27302), .B(n27301), .Z(n27350) );
  XOR U28019 ( .A(n27351), .B(n27350), .Z(n27352) );
  NANDN U28020 ( .A(n27304), .B(n27303), .Z(n27308) );
  NANDN U28021 ( .A(n27306), .B(n27305), .Z(n27307) );
  NAND U28022 ( .A(n27308), .B(n27307), .Z(n27353) );
  XOR U28023 ( .A(n27352), .B(n27353), .Z(n27320) );
  OR U28024 ( .A(n27310), .B(n27309), .Z(n27314) );
  NANDN U28025 ( .A(n27312), .B(n27311), .Z(n27313) );
  NAND U28026 ( .A(n27314), .B(n27313), .Z(n27321) );
  XNOR U28027 ( .A(n27320), .B(n27321), .Z(n27322) );
  XNOR U28028 ( .A(n27323), .B(n27322), .Z(n27356) );
  XNOR U28029 ( .A(n27356), .B(sreg[1680]), .Z(n27358) );
  NAND U28030 ( .A(n27315), .B(sreg[1679]), .Z(n27319) );
  OR U28031 ( .A(n27317), .B(n27316), .Z(n27318) );
  AND U28032 ( .A(n27319), .B(n27318), .Z(n27357) );
  XOR U28033 ( .A(n27358), .B(n27357), .Z(c[1680]) );
  NANDN U28034 ( .A(n27321), .B(n27320), .Z(n27325) );
  NAND U28035 ( .A(n27323), .B(n27322), .Z(n27324) );
  NAND U28036 ( .A(n27325), .B(n27324), .Z(n27364) );
  NAND U28037 ( .A(b[0]), .B(a[665]), .Z(n27326) );
  XNOR U28038 ( .A(b[1]), .B(n27326), .Z(n27328) );
  NAND U28039 ( .A(n110), .B(a[664]), .Z(n27327) );
  AND U28040 ( .A(n27328), .B(n27327), .Z(n27381) );
  XOR U28041 ( .A(a[661]), .B(n42197), .Z(n27370) );
  NANDN U28042 ( .A(n27370), .B(n42173), .Z(n27331) );
  NANDN U28043 ( .A(n27329), .B(n42172), .Z(n27330) );
  NAND U28044 ( .A(n27331), .B(n27330), .Z(n27379) );
  NAND U28045 ( .A(b[7]), .B(a[657]), .Z(n27380) );
  XNOR U28046 ( .A(n27379), .B(n27380), .Z(n27382) );
  XOR U28047 ( .A(n27381), .B(n27382), .Z(n27388) );
  NANDN U28048 ( .A(n27332), .B(n42093), .Z(n27334) );
  XOR U28049 ( .A(n42134), .B(a[663]), .Z(n27373) );
  NANDN U28050 ( .A(n27373), .B(n42095), .Z(n27333) );
  NAND U28051 ( .A(n27334), .B(n27333), .Z(n27386) );
  NANDN U28052 ( .A(n27335), .B(n42231), .Z(n27337) );
  XOR U28053 ( .A(n217), .B(a[659]), .Z(n27376) );
  NANDN U28054 ( .A(n27376), .B(n42234), .Z(n27336) );
  AND U28055 ( .A(n27337), .B(n27336), .Z(n27385) );
  XNOR U28056 ( .A(n27386), .B(n27385), .Z(n27387) );
  XNOR U28057 ( .A(n27388), .B(n27387), .Z(n27392) );
  NANDN U28058 ( .A(n27339), .B(n27338), .Z(n27343) );
  NAND U28059 ( .A(n27341), .B(n27340), .Z(n27342) );
  AND U28060 ( .A(n27343), .B(n27342), .Z(n27391) );
  XOR U28061 ( .A(n27392), .B(n27391), .Z(n27393) );
  NANDN U28062 ( .A(n27345), .B(n27344), .Z(n27349) );
  NANDN U28063 ( .A(n27347), .B(n27346), .Z(n27348) );
  NAND U28064 ( .A(n27349), .B(n27348), .Z(n27394) );
  XOR U28065 ( .A(n27393), .B(n27394), .Z(n27361) );
  OR U28066 ( .A(n27351), .B(n27350), .Z(n27355) );
  NANDN U28067 ( .A(n27353), .B(n27352), .Z(n27354) );
  NAND U28068 ( .A(n27355), .B(n27354), .Z(n27362) );
  XNOR U28069 ( .A(n27361), .B(n27362), .Z(n27363) );
  XNOR U28070 ( .A(n27364), .B(n27363), .Z(n27397) );
  XNOR U28071 ( .A(n27397), .B(sreg[1681]), .Z(n27399) );
  NAND U28072 ( .A(n27356), .B(sreg[1680]), .Z(n27360) );
  OR U28073 ( .A(n27358), .B(n27357), .Z(n27359) );
  AND U28074 ( .A(n27360), .B(n27359), .Z(n27398) );
  XOR U28075 ( .A(n27399), .B(n27398), .Z(c[1681]) );
  NANDN U28076 ( .A(n27362), .B(n27361), .Z(n27366) );
  NAND U28077 ( .A(n27364), .B(n27363), .Z(n27365) );
  NAND U28078 ( .A(n27366), .B(n27365), .Z(n27405) );
  NAND U28079 ( .A(b[0]), .B(a[666]), .Z(n27367) );
  XNOR U28080 ( .A(b[1]), .B(n27367), .Z(n27369) );
  NAND U28081 ( .A(n110), .B(a[665]), .Z(n27368) );
  AND U28082 ( .A(n27369), .B(n27368), .Z(n27422) );
  XOR U28083 ( .A(a[662]), .B(n42197), .Z(n27411) );
  NANDN U28084 ( .A(n27411), .B(n42173), .Z(n27372) );
  NANDN U28085 ( .A(n27370), .B(n42172), .Z(n27371) );
  NAND U28086 ( .A(n27372), .B(n27371), .Z(n27420) );
  NAND U28087 ( .A(b[7]), .B(a[658]), .Z(n27421) );
  XNOR U28088 ( .A(n27420), .B(n27421), .Z(n27423) );
  XOR U28089 ( .A(n27422), .B(n27423), .Z(n27429) );
  NANDN U28090 ( .A(n27373), .B(n42093), .Z(n27375) );
  XOR U28091 ( .A(n42134), .B(a[664]), .Z(n27414) );
  NANDN U28092 ( .A(n27414), .B(n42095), .Z(n27374) );
  NAND U28093 ( .A(n27375), .B(n27374), .Z(n27427) );
  NANDN U28094 ( .A(n27376), .B(n42231), .Z(n27378) );
  XOR U28095 ( .A(n217), .B(a[660]), .Z(n27417) );
  NANDN U28096 ( .A(n27417), .B(n42234), .Z(n27377) );
  AND U28097 ( .A(n27378), .B(n27377), .Z(n27426) );
  XNOR U28098 ( .A(n27427), .B(n27426), .Z(n27428) );
  XNOR U28099 ( .A(n27429), .B(n27428), .Z(n27433) );
  NANDN U28100 ( .A(n27380), .B(n27379), .Z(n27384) );
  NAND U28101 ( .A(n27382), .B(n27381), .Z(n27383) );
  AND U28102 ( .A(n27384), .B(n27383), .Z(n27432) );
  XOR U28103 ( .A(n27433), .B(n27432), .Z(n27434) );
  NANDN U28104 ( .A(n27386), .B(n27385), .Z(n27390) );
  NANDN U28105 ( .A(n27388), .B(n27387), .Z(n27389) );
  NAND U28106 ( .A(n27390), .B(n27389), .Z(n27435) );
  XOR U28107 ( .A(n27434), .B(n27435), .Z(n27402) );
  OR U28108 ( .A(n27392), .B(n27391), .Z(n27396) );
  NANDN U28109 ( .A(n27394), .B(n27393), .Z(n27395) );
  NAND U28110 ( .A(n27396), .B(n27395), .Z(n27403) );
  XNOR U28111 ( .A(n27402), .B(n27403), .Z(n27404) );
  XNOR U28112 ( .A(n27405), .B(n27404), .Z(n27438) );
  XNOR U28113 ( .A(n27438), .B(sreg[1682]), .Z(n27440) );
  NAND U28114 ( .A(n27397), .B(sreg[1681]), .Z(n27401) );
  OR U28115 ( .A(n27399), .B(n27398), .Z(n27400) );
  AND U28116 ( .A(n27401), .B(n27400), .Z(n27439) );
  XOR U28117 ( .A(n27440), .B(n27439), .Z(c[1682]) );
  NANDN U28118 ( .A(n27403), .B(n27402), .Z(n27407) );
  NAND U28119 ( .A(n27405), .B(n27404), .Z(n27406) );
  NAND U28120 ( .A(n27407), .B(n27406), .Z(n27446) );
  NAND U28121 ( .A(b[0]), .B(a[667]), .Z(n27408) );
  XNOR U28122 ( .A(b[1]), .B(n27408), .Z(n27410) );
  NAND U28123 ( .A(n110), .B(a[666]), .Z(n27409) );
  AND U28124 ( .A(n27410), .B(n27409), .Z(n27463) );
  XOR U28125 ( .A(a[663]), .B(n42197), .Z(n27452) );
  NANDN U28126 ( .A(n27452), .B(n42173), .Z(n27413) );
  NANDN U28127 ( .A(n27411), .B(n42172), .Z(n27412) );
  NAND U28128 ( .A(n27413), .B(n27412), .Z(n27461) );
  NAND U28129 ( .A(b[7]), .B(a[659]), .Z(n27462) );
  XNOR U28130 ( .A(n27461), .B(n27462), .Z(n27464) );
  XOR U28131 ( .A(n27463), .B(n27464), .Z(n27470) );
  NANDN U28132 ( .A(n27414), .B(n42093), .Z(n27416) );
  XOR U28133 ( .A(n42134), .B(a[665]), .Z(n27455) );
  NANDN U28134 ( .A(n27455), .B(n42095), .Z(n27415) );
  NAND U28135 ( .A(n27416), .B(n27415), .Z(n27468) );
  NANDN U28136 ( .A(n27417), .B(n42231), .Z(n27419) );
  XOR U28137 ( .A(n217), .B(a[661]), .Z(n27458) );
  NANDN U28138 ( .A(n27458), .B(n42234), .Z(n27418) );
  AND U28139 ( .A(n27419), .B(n27418), .Z(n27467) );
  XNOR U28140 ( .A(n27468), .B(n27467), .Z(n27469) );
  XNOR U28141 ( .A(n27470), .B(n27469), .Z(n27474) );
  NANDN U28142 ( .A(n27421), .B(n27420), .Z(n27425) );
  NAND U28143 ( .A(n27423), .B(n27422), .Z(n27424) );
  AND U28144 ( .A(n27425), .B(n27424), .Z(n27473) );
  XOR U28145 ( .A(n27474), .B(n27473), .Z(n27475) );
  NANDN U28146 ( .A(n27427), .B(n27426), .Z(n27431) );
  NANDN U28147 ( .A(n27429), .B(n27428), .Z(n27430) );
  NAND U28148 ( .A(n27431), .B(n27430), .Z(n27476) );
  XOR U28149 ( .A(n27475), .B(n27476), .Z(n27443) );
  OR U28150 ( .A(n27433), .B(n27432), .Z(n27437) );
  NANDN U28151 ( .A(n27435), .B(n27434), .Z(n27436) );
  NAND U28152 ( .A(n27437), .B(n27436), .Z(n27444) );
  XNOR U28153 ( .A(n27443), .B(n27444), .Z(n27445) );
  XNOR U28154 ( .A(n27446), .B(n27445), .Z(n27479) );
  XNOR U28155 ( .A(n27479), .B(sreg[1683]), .Z(n27481) );
  NAND U28156 ( .A(n27438), .B(sreg[1682]), .Z(n27442) );
  OR U28157 ( .A(n27440), .B(n27439), .Z(n27441) );
  AND U28158 ( .A(n27442), .B(n27441), .Z(n27480) );
  XOR U28159 ( .A(n27481), .B(n27480), .Z(c[1683]) );
  NANDN U28160 ( .A(n27444), .B(n27443), .Z(n27448) );
  NAND U28161 ( .A(n27446), .B(n27445), .Z(n27447) );
  NAND U28162 ( .A(n27448), .B(n27447), .Z(n27487) );
  NAND U28163 ( .A(b[0]), .B(a[668]), .Z(n27449) );
  XNOR U28164 ( .A(b[1]), .B(n27449), .Z(n27451) );
  NAND U28165 ( .A(n110), .B(a[667]), .Z(n27450) );
  AND U28166 ( .A(n27451), .B(n27450), .Z(n27504) );
  XOR U28167 ( .A(a[664]), .B(n42197), .Z(n27493) );
  NANDN U28168 ( .A(n27493), .B(n42173), .Z(n27454) );
  NANDN U28169 ( .A(n27452), .B(n42172), .Z(n27453) );
  NAND U28170 ( .A(n27454), .B(n27453), .Z(n27502) );
  NAND U28171 ( .A(b[7]), .B(a[660]), .Z(n27503) );
  XNOR U28172 ( .A(n27502), .B(n27503), .Z(n27505) );
  XOR U28173 ( .A(n27504), .B(n27505), .Z(n27511) );
  NANDN U28174 ( .A(n27455), .B(n42093), .Z(n27457) );
  XOR U28175 ( .A(n42134), .B(a[666]), .Z(n27496) );
  NANDN U28176 ( .A(n27496), .B(n42095), .Z(n27456) );
  NAND U28177 ( .A(n27457), .B(n27456), .Z(n27509) );
  NANDN U28178 ( .A(n27458), .B(n42231), .Z(n27460) );
  XOR U28179 ( .A(n217), .B(a[662]), .Z(n27499) );
  NANDN U28180 ( .A(n27499), .B(n42234), .Z(n27459) );
  AND U28181 ( .A(n27460), .B(n27459), .Z(n27508) );
  XNOR U28182 ( .A(n27509), .B(n27508), .Z(n27510) );
  XNOR U28183 ( .A(n27511), .B(n27510), .Z(n27515) );
  NANDN U28184 ( .A(n27462), .B(n27461), .Z(n27466) );
  NAND U28185 ( .A(n27464), .B(n27463), .Z(n27465) );
  AND U28186 ( .A(n27466), .B(n27465), .Z(n27514) );
  XOR U28187 ( .A(n27515), .B(n27514), .Z(n27516) );
  NANDN U28188 ( .A(n27468), .B(n27467), .Z(n27472) );
  NANDN U28189 ( .A(n27470), .B(n27469), .Z(n27471) );
  NAND U28190 ( .A(n27472), .B(n27471), .Z(n27517) );
  XOR U28191 ( .A(n27516), .B(n27517), .Z(n27484) );
  OR U28192 ( .A(n27474), .B(n27473), .Z(n27478) );
  NANDN U28193 ( .A(n27476), .B(n27475), .Z(n27477) );
  NAND U28194 ( .A(n27478), .B(n27477), .Z(n27485) );
  XNOR U28195 ( .A(n27484), .B(n27485), .Z(n27486) );
  XNOR U28196 ( .A(n27487), .B(n27486), .Z(n27520) );
  XNOR U28197 ( .A(n27520), .B(sreg[1684]), .Z(n27522) );
  NAND U28198 ( .A(n27479), .B(sreg[1683]), .Z(n27483) );
  OR U28199 ( .A(n27481), .B(n27480), .Z(n27482) );
  AND U28200 ( .A(n27483), .B(n27482), .Z(n27521) );
  XOR U28201 ( .A(n27522), .B(n27521), .Z(c[1684]) );
  NANDN U28202 ( .A(n27485), .B(n27484), .Z(n27489) );
  NAND U28203 ( .A(n27487), .B(n27486), .Z(n27488) );
  NAND U28204 ( .A(n27489), .B(n27488), .Z(n27528) );
  NAND U28205 ( .A(b[0]), .B(a[669]), .Z(n27490) );
  XNOR U28206 ( .A(b[1]), .B(n27490), .Z(n27492) );
  NAND U28207 ( .A(n110), .B(a[668]), .Z(n27491) );
  AND U28208 ( .A(n27492), .B(n27491), .Z(n27545) );
  XOR U28209 ( .A(a[665]), .B(n42197), .Z(n27534) );
  NANDN U28210 ( .A(n27534), .B(n42173), .Z(n27495) );
  NANDN U28211 ( .A(n27493), .B(n42172), .Z(n27494) );
  NAND U28212 ( .A(n27495), .B(n27494), .Z(n27543) );
  NAND U28213 ( .A(b[7]), .B(a[661]), .Z(n27544) );
  XNOR U28214 ( .A(n27543), .B(n27544), .Z(n27546) );
  XOR U28215 ( .A(n27545), .B(n27546), .Z(n27552) );
  NANDN U28216 ( .A(n27496), .B(n42093), .Z(n27498) );
  XOR U28217 ( .A(n42134), .B(a[667]), .Z(n27537) );
  NANDN U28218 ( .A(n27537), .B(n42095), .Z(n27497) );
  NAND U28219 ( .A(n27498), .B(n27497), .Z(n27550) );
  NANDN U28220 ( .A(n27499), .B(n42231), .Z(n27501) );
  XOR U28221 ( .A(n217), .B(a[663]), .Z(n27540) );
  NANDN U28222 ( .A(n27540), .B(n42234), .Z(n27500) );
  AND U28223 ( .A(n27501), .B(n27500), .Z(n27549) );
  XNOR U28224 ( .A(n27550), .B(n27549), .Z(n27551) );
  XNOR U28225 ( .A(n27552), .B(n27551), .Z(n27556) );
  NANDN U28226 ( .A(n27503), .B(n27502), .Z(n27507) );
  NAND U28227 ( .A(n27505), .B(n27504), .Z(n27506) );
  AND U28228 ( .A(n27507), .B(n27506), .Z(n27555) );
  XOR U28229 ( .A(n27556), .B(n27555), .Z(n27557) );
  NANDN U28230 ( .A(n27509), .B(n27508), .Z(n27513) );
  NANDN U28231 ( .A(n27511), .B(n27510), .Z(n27512) );
  NAND U28232 ( .A(n27513), .B(n27512), .Z(n27558) );
  XOR U28233 ( .A(n27557), .B(n27558), .Z(n27525) );
  OR U28234 ( .A(n27515), .B(n27514), .Z(n27519) );
  NANDN U28235 ( .A(n27517), .B(n27516), .Z(n27518) );
  NAND U28236 ( .A(n27519), .B(n27518), .Z(n27526) );
  XNOR U28237 ( .A(n27525), .B(n27526), .Z(n27527) );
  XNOR U28238 ( .A(n27528), .B(n27527), .Z(n27561) );
  XNOR U28239 ( .A(n27561), .B(sreg[1685]), .Z(n27563) );
  NAND U28240 ( .A(n27520), .B(sreg[1684]), .Z(n27524) );
  OR U28241 ( .A(n27522), .B(n27521), .Z(n27523) );
  AND U28242 ( .A(n27524), .B(n27523), .Z(n27562) );
  XOR U28243 ( .A(n27563), .B(n27562), .Z(c[1685]) );
  NANDN U28244 ( .A(n27526), .B(n27525), .Z(n27530) );
  NAND U28245 ( .A(n27528), .B(n27527), .Z(n27529) );
  NAND U28246 ( .A(n27530), .B(n27529), .Z(n27569) );
  NAND U28247 ( .A(b[0]), .B(a[670]), .Z(n27531) );
  XNOR U28248 ( .A(b[1]), .B(n27531), .Z(n27533) );
  NAND U28249 ( .A(n110), .B(a[669]), .Z(n27532) );
  AND U28250 ( .A(n27533), .B(n27532), .Z(n27586) );
  XOR U28251 ( .A(a[666]), .B(n42197), .Z(n27575) );
  NANDN U28252 ( .A(n27575), .B(n42173), .Z(n27536) );
  NANDN U28253 ( .A(n27534), .B(n42172), .Z(n27535) );
  NAND U28254 ( .A(n27536), .B(n27535), .Z(n27584) );
  NAND U28255 ( .A(b[7]), .B(a[662]), .Z(n27585) );
  XNOR U28256 ( .A(n27584), .B(n27585), .Z(n27587) );
  XOR U28257 ( .A(n27586), .B(n27587), .Z(n27593) );
  NANDN U28258 ( .A(n27537), .B(n42093), .Z(n27539) );
  XOR U28259 ( .A(n42134), .B(a[668]), .Z(n27578) );
  NANDN U28260 ( .A(n27578), .B(n42095), .Z(n27538) );
  NAND U28261 ( .A(n27539), .B(n27538), .Z(n27591) );
  NANDN U28262 ( .A(n27540), .B(n42231), .Z(n27542) );
  XOR U28263 ( .A(n217), .B(a[664]), .Z(n27581) );
  NANDN U28264 ( .A(n27581), .B(n42234), .Z(n27541) );
  AND U28265 ( .A(n27542), .B(n27541), .Z(n27590) );
  XNOR U28266 ( .A(n27591), .B(n27590), .Z(n27592) );
  XNOR U28267 ( .A(n27593), .B(n27592), .Z(n27597) );
  NANDN U28268 ( .A(n27544), .B(n27543), .Z(n27548) );
  NAND U28269 ( .A(n27546), .B(n27545), .Z(n27547) );
  AND U28270 ( .A(n27548), .B(n27547), .Z(n27596) );
  XOR U28271 ( .A(n27597), .B(n27596), .Z(n27598) );
  NANDN U28272 ( .A(n27550), .B(n27549), .Z(n27554) );
  NANDN U28273 ( .A(n27552), .B(n27551), .Z(n27553) );
  NAND U28274 ( .A(n27554), .B(n27553), .Z(n27599) );
  XOR U28275 ( .A(n27598), .B(n27599), .Z(n27566) );
  OR U28276 ( .A(n27556), .B(n27555), .Z(n27560) );
  NANDN U28277 ( .A(n27558), .B(n27557), .Z(n27559) );
  NAND U28278 ( .A(n27560), .B(n27559), .Z(n27567) );
  XNOR U28279 ( .A(n27566), .B(n27567), .Z(n27568) );
  XNOR U28280 ( .A(n27569), .B(n27568), .Z(n27602) );
  XNOR U28281 ( .A(n27602), .B(sreg[1686]), .Z(n27604) );
  NAND U28282 ( .A(n27561), .B(sreg[1685]), .Z(n27565) );
  OR U28283 ( .A(n27563), .B(n27562), .Z(n27564) );
  AND U28284 ( .A(n27565), .B(n27564), .Z(n27603) );
  XOR U28285 ( .A(n27604), .B(n27603), .Z(c[1686]) );
  NANDN U28286 ( .A(n27567), .B(n27566), .Z(n27571) );
  NAND U28287 ( .A(n27569), .B(n27568), .Z(n27570) );
  NAND U28288 ( .A(n27571), .B(n27570), .Z(n27610) );
  NAND U28289 ( .A(b[0]), .B(a[671]), .Z(n27572) );
  XNOR U28290 ( .A(b[1]), .B(n27572), .Z(n27574) );
  NAND U28291 ( .A(n110), .B(a[670]), .Z(n27573) );
  AND U28292 ( .A(n27574), .B(n27573), .Z(n27627) );
  XOR U28293 ( .A(a[667]), .B(n42197), .Z(n27616) );
  NANDN U28294 ( .A(n27616), .B(n42173), .Z(n27577) );
  NANDN U28295 ( .A(n27575), .B(n42172), .Z(n27576) );
  NAND U28296 ( .A(n27577), .B(n27576), .Z(n27625) );
  NAND U28297 ( .A(b[7]), .B(a[663]), .Z(n27626) );
  XNOR U28298 ( .A(n27625), .B(n27626), .Z(n27628) );
  XOR U28299 ( .A(n27627), .B(n27628), .Z(n27634) );
  NANDN U28300 ( .A(n27578), .B(n42093), .Z(n27580) );
  XOR U28301 ( .A(n42134), .B(a[669]), .Z(n27619) );
  NANDN U28302 ( .A(n27619), .B(n42095), .Z(n27579) );
  NAND U28303 ( .A(n27580), .B(n27579), .Z(n27632) );
  NANDN U28304 ( .A(n27581), .B(n42231), .Z(n27583) );
  XOR U28305 ( .A(n217), .B(a[665]), .Z(n27622) );
  NANDN U28306 ( .A(n27622), .B(n42234), .Z(n27582) );
  AND U28307 ( .A(n27583), .B(n27582), .Z(n27631) );
  XNOR U28308 ( .A(n27632), .B(n27631), .Z(n27633) );
  XNOR U28309 ( .A(n27634), .B(n27633), .Z(n27638) );
  NANDN U28310 ( .A(n27585), .B(n27584), .Z(n27589) );
  NAND U28311 ( .A(n27587), .B(n27586), .Z(n27588) );
  AND U28312 ( .A(n27589), .B(n27588), .Z(n27637) );
  XOR U28313 ( .A(n27638), .B(n27637), .Z(n27639) );
  NANDN U28314 ( .A(n27591), .B(n27590), .Z(n27595) );
  NANDN U28315 ( .A(n27593), .B(n27592), .Z(n27594) );
  NAND U28316 ( .A(n27595), .B(n27594), .Z(n27640) );
  XOR U28317 ( .A(n27639), .B(n27640), .Z(n27607) );
  OR U28318 ( .A(n27597), .B(n27596), .Z(n27601) );
  NANDN U28319 ( .A(n27599), .B(n27598), .Z(n27600) );
  NAND U28320 ( .A(n27601), .B(n27600), .Z(n27608) );
  XNOR U28321 ( .A(n27607), .B(n27608), .Z(n27609) );
  XNOR U28322 ( .A(n27610), .B(n27609), .Z(n27643) );
  XNOR U28323 ( .A(n27643), .B(sreg[1687]), .Z(n27645) );
  NAND U28324 ( .A(n27602), .B(sreg[1686]), .Z(n27606) );
  OR U28325 ( .A(n27604), .B(n27603), .Z(n27605) );
  AND U28326 ( .A(n27606), .B(n27605), .Z(n27644) );
  XOR U28327 ( .A(n27645), .B(n27644), .Z(c[1687]) );
  NANDN U28328 ( .A(n27608), .B(n27607), .Z(n27612) );
  NAND U28329 ( .A(n27610), .B(n27609), .Z(n27611) );
  NAND U28330 ( .A(n27612), .B(n27611), .Z(n27651) );
  NAND U28331 ( .A(b[0]), .B(a[672]), .Z(n27613) );
  XNOR U28332 ( .A(b[1]), .B(n27613), .Z(n27615) );
  NAND U28333 ( .A(n111), .B(a[671]), .Z(n27614) );
  AND U28334 ( .A(n27615), .B(n27614), .Z(n27668) );
  XOR U28335 ( .A(a[668]), .B(n42197), .Z(n27657) );
  NANDN U28336 ( .A(n27657), .B(n42173), .Z(n27618) );
  NANDN U28337 ( .A(n27616), .B(n42172), .Z(n27617) );
  NAND U28338 ( .A(n27618), .B(n27617), .Z(n27666) );
  NAND U28339 ( .A(b[7]), .B(a[664]), .Z(n27667) );
  XNOR U28340 ( .A(n27666), .B(n27667), .Z(n27669) );
  XOR U28341 ( .A(n27668), .B(n27669), .Z(n27675) );
  NANDN U28342 ( .A(n27619), .B(n42093), .Z(n27621) );
  XOR U28343 ( .A(n42134), .B(a[670]), .Z(n27660) );
  NANDN U28344 ( .A(n27660), .B(n42095), .Z(n27620) );
  NAND U28345 ( .A(n27621), .B(n27620), .Z(n27673) );
  NANDN U28346 ( .A(n27622), .B(n42231), .Z(n27624) );
  XOR U28347 ( .A(n217), .B(a[666]), .Z(n27663) );
  NANDN U28348 ( .A(n27663), .B(n42234), .Z(n27623) );
  AND U28349 ( .A(n27624), .B(n27623), .Z(n27672) );
  XNOR U28350 ( .A(n27673), .B(n27672), .Z(n27674) );
  XNOR U28351 ( .A(n27675), .B(n27674), .Z(n27679) );
  NANDN U28352 ( .A(n27626), .B(n27625), .Z(n27630) );
  NAND U28353 ( .A(n27628), .B(n27627), .Z(n27629) );
  AND U28354 ( .A(n27630), .B(n27629), .Z(n27678) );
  XOR U28355 ( .A(n27679), .B(n27678), .Z(n27680) );
  NANDN U28356 ( .A(n27632), .B(n27631), .Z(n27636) );
  NANDN U28357 ( .A(n27634), .B(n27633), .Z(n27635) );
  NAND U28358 ( .A(n27636), .B(n27635), .Z(n27681) );
  XOR U28359 ( .A(n27680), .B(n27681), .Z(n27648) );
  OR U28360 ( .A(n27638), .B(n27637), .Z(n27642) );
  NANDN U28361 ( .A(n27640), .B(n27639), .Z(n27641) );
  NAND U28362 ( .A(n27642), .B(n27641), .Z(n27649) );
  XNOR U28363 ( .A(n27648), .B(n27649), .Z(n27650) );
  XNOR U28364 ( .A(n27651), .B(n27650), .Z(n27684) );
  XNOR U28365 ( .A(n27684), .B(sreg[1688]), .Z(n27686) );
  NAND U28366 ( .A(n27643), .B(sreg[1687]), .Z(n27647) );
  OR U28367 ( .A(n27645), .B(n27644), .Z(n27646) );
  AND U28368 ( .A(n27647), .B(n27646), .Z(n27685) );
  XOR U28369 ( .A(n27686), .B(n27685), .Z(c[1688]) );
  NANDN U28370 ( .A(n27649), .B(n27648), .Z(n27653) );
  NAND U28371 ( .A(n27651), .B(n27650), .Z(n27652) );
  NAND U28372 ( .A(n27653), .B(n27652), .Z(n27692) );
  NAND U28373 ( .A(b[0]), .B(a[673]), .Z(n27654) );
  XNOR U28374 ( .A(b[1]), .B(n27654), .Z(n27656) );
  NAND U28375 ( .A(n111), .B(a[672]), .Z(n27655) );
  AND U28376 ( .A(n27656), .B(n27655), .Z(n27709) );
  XOR U28377 ( .A(a[669]), .B(n42197), .Z(n27698) );
  NANDN U28378 ( .A(n27698), .B(n42173), .Z(n27659) );
  NANDN U28379 ( .A(n27657), .B(n42172), .Z(n27658) );
  NAND U28380 ( .A(n27659), .B(n27658), .Z(n27707) );
  NAND U28381 ( .A(b[7]), .B(a[665]), .Z(n27708) );
  XNOR U28382 ( .A(n27707), .B(n27708), .Z(n27710) );
  XOR U28383 ( .A(n27709), .B(n27710), .Z(n27716) );
  NANDN U28384 ( .A(n27660), .B(n42093), .Z(n27662) );
  XOR U28385 ( .A(n42134), .B(a[671]), .Z(n27701) );
  NANDN U28386 ( .A(n27701), .B(n42095), .Z(n27661) );
  NAND U28387 ( .A(n27662), .B(n27661), .Z(n27714) );
  NANDN U28388 ( .A(n27663), .B(n42231), .Z(n27665) );
  XOR U28389 ( .A(n217), .B(a[667]), .Z(n27704) );
  NANDN U28390 ( .A(n27704), .B(n42234), .Z(n27664) );
  AND U28391 ( .A(n27665), .B(n27664), .Z(n27713) );
  XNOR U28392 ( .A(n27714), .B(n27713), .Z(n27715) );
  XNOR U28393 ( .A(n27716), .B(n27715), .Z(n27720) );
  NANDN U28394 ( .A(n27667), .B(n27666), .Z(n27671) );
  NAND U28395 ( .A(n27669), .B(n27668), .Z(n27670) );
  AND U28396 ( .A(n27671), .B(n27670), .Z(n27719) );
  XOR U28397 ( .A(n27720), .B(n27719), .Z(n27721) );
  NANDN U28398 ( .A(n27673), .B(n27672), .Z(n27677) );
  NANDN U28399 ( .A(n27675), .B(n27674), .Z(n27676) );
  NAND U28400 ( .A(n27677), .B(n27676), .Z(n27722) );
  XOR U28401 ( .A(n27721), .B(n27722), .Z(n27689) );
  OR U28402 ( .A(n27679), .B(n27678), .Z(n27683) );
  NANDN U28403 ( .A(n27681), .B(n27680), .Z(n27682) );
  NAND U28404 ( .A(n27683), .B(n27682), .Z(n27690) );
  XNOR U28405 ( .A(n27689), .B(n27690), .Z(n27691) );
  XNOR U28406 ( .A(n27692), .B(n27691), .Z(n27725) );
  XNOR U28407 ( .A(n27725), .B(sreg[1689]), .Z(n27727) );
  NAND U28408 ( .A(n27684), .B(sreg[1688]), .Z(n27688) );
  OR U28409 ( .A(n27686), .B(n27685), .Z(n27687) );
  AND U28410 ( .A(n27688), .B(n27687), .Z(n27726) );
  XOR U28411 ( .A(n27727), .B(n27726), .Z(c[1689]) );
  NANDN U28412 ( .A(n27690), .B(n27689), .Z(n27694) );
  NAND U28413 ( .A(n27692), .B(n27691), .Z(n27693) );
  NAND U28414 ( .A(n27694), .B(n27693), .Z(n27733) );
  NAND U28415 ( .A(b[0]), .B(a[674]), .Z(n27695) );
  XNOR U28416 ( .A(b[1]), .B(n27695), .Z(n27697) );
  NAND U28417 ( .A(n111), .B(a[673]), .Z(n27696) );
  AND U28418 ( .A(n27697), .B(n27696), .Z(n27750) );
  XOR U28419 ( .A(a[670]), .B(n42197), .Z(n27739) );
  NANDN U28420 ( .A(n27739), .B(n42173), .Z(n27700) );
  NANDN U28421 ( .A(n27698), .B(n42172), .Z(n27699) );
  NAND U28422 ( .A(n27700), .B(n27699), .Z(n27748) );
  NAND U28423 ( .A(b[7]), .B(a[666]), .Z(n27749) );
  XNOR U28424 ( .A(n27748), .B(n27749), .Z(n27751) );
  XOR U28425 ( .A(n27750), .B(n27751), .Z(n27757) );
  NANDN U28426 ( .A(n27701), .B(n42093), .Z(n27703) );
  XOR U28427 ( .A(n42134), .B(a[672]), .Z(n27742) );
  NANDN U28428 ( .A(n27742), .B(n42095), .Z(n27702) );
  NAND U28429 ( .A(n27703), .B(n27702), .Z(n27755) );
  NANDN U28430 ( .A(n27704), .B(n42231), .Z(n27706) );
  XOR U28431 ( .A(n217), .B(a[668]), .Z(n27745) );
  NANDN U28432 ( .A(n27745), .B(n42234), .Z(n27705) );
  AND U28433 ( .A(n27706), .B(n27705), .Z(n27754) );
  XNOR U28434 ( .A(n27755), .B(n27754), .Z(n27756) );
  XNOR U28435 ( .A(n27757), .B(n27756), .Z(n27761) );
  NANDN U28436 ( .A(n27708), .B(n27707), .Z(n27712) );
  NAND U28437 ( .A(n27710), .B(n27709), .Z(n27711) );
  AND U28438 ( .A(n27712), .B(n27711), .Z(n27760) );
  XOR U28439 ( .A(n27761), .B(n27760), .Z(n27762) );
  NANDN U28440 ( .A(n27714), .B(n27713), .Z(n27718) );
  NANDN U28441 ( .A(n27716), .B(n27715), .Z(n27717) );
  NAND U28442 ( .A(n27718), .B(n27717), .Z(n27763) );
  XOR U28443 ( .A(n27762), .B(n27763), .Z(n27730) );
  OR U28444 ( .A(n27720), .B(n27719), .Z(n27724) );
  NANDN U28445 ( .A(n27722), .B(n27721), .Z(n27723) );
  NAND U28446 ( .A(n27724), .B(n27723), .Z(n27731) );
  XNOR U28447 ( .A(n27730), .B(n27731), .Z(n27732) );
  XNOR U28448 ( .A(n27733), .B(n27732), .Z(n27766) );
  XNOR U28449 ( .A(n27766), .B(sreg[1690]), .Z(n27768) );
  NAND U28450 ( .A(n27725), .B(sreg[1689]), .Z(n27729) );
  OR U28451 ( .A(n27727), .B(n27726), .Z(n27728) );
  AND U28452 ( .A(n27729), .B(n27728), .Z(n27767) );
  XOR U28453 ( .A(n27768), .B(n27767), .Z(c[1690]) );
  NANDN U28454 ( .A(n27731), .B(n27730), .Z(n27735) );
  NAND U28455 ( .A(n27733), .B(n27732), .Z(n27734) );
  NAND U28456 ( .A(n27735), .B(n27734), .Z(n27774) );
  NAND U28457 ( .A(b[0]), .B(a[675]), .Z(n27736) );
  XNOR U28458 ( .A(b[1]), .B(n27736), .Z(n27738) );
  NAND U28459 ( .A(n111), .B(a[674]), .Z(n27737) );
  AND U28460 ( .A(n27738), .B(n27737), .Z(n27791) );
  XOR U28461 ( .A(a[671]), .B(n42197), .Z(n27780) );
  NANDN U28462 ( .A(n27780), .B(n42173), .Z(n27741) );
  NANDN U28463 ( .A(n27739), .B(n42172), .Z(n27740) );
  NAND U28464 ( .A(n27741), .B(n27740), .Z(n27789) );
  NAND U28465 ( .A(b[7]), .B(a[667]), .Z(n27790) );
  XNOR U28466 ( .A(n27789), .B(n27790), .Z(n27792) );
  XOR U28467 ( .A(n27791), .B(n27792), .Z(n27798) );
  NANDN U28468 ( .A(n27742), .B(n42093), .Z(n27744) );
  XOR U28469 ( .A(n42134), .B(a[673]), .Z(n27783) );
  NANDN U28470 ( .A(n27783), .B(n42095), .Z(n27743) );
  NAND U28471 ( .A(n27744), .B(n27743), .Z(n27796) );
  NANDN U28472 ( .A(n27745), .B(n42231), .Z(n27747) );
  XOR U28473 ( .A(n217), .B(a[669]), .Z(n27786) );
  NANDN U28474 ( .A(n27786), .B(n42234), .Z(n27746) );
  AND U28475 ( .A(n27747), .B(n27746), .Z(n27795) );
  XNOR U28476 ( .A(n27796), .B(n27795), .Z(n27797) );
  XNOR U28477 ( .A(n27798), .B(n27797), .Z(n27802) );
  NANDN U28478 ( .A(n27749), .B(n27748), .Z(n27753) );
  NAND U28479 ( .A(n27751), .B(n27750), .Z(n27752) );
  AND U28480 ( .A(n27753), .B(n27752), .Z(n27801) );
  XOR U28481 ( .A(n27802), .B(n27801), .Z(n27803) );
  NANDN U28482 ( .A(n27755), .B(n27754), .Z(n27759) );
  NANDN U28483 ( .A(n27757), .B(n27756), .Z(n27758) );
  NAND U28484 ( .A(n27759), .B(n27758), .Z(n27804) );
  XOR U28485 ( .A(n27803), .B(n27804), .Z(n27771) );
  OR U28486 ( .A(n27761), .B(n27760), .Z(n27765) );
  NANDN U28487 ( .A(n27763), .B(n27762), .Z(n27764) );
  NAND U28488 ( .A(n27765), .B(n27764), .Z(n27772) );
  XNOR U28489 ( .A(n27771), .B(n27772), .Z(n27773) );
  XNOR U28490 ( .A(n27774), .B(n27773), .Z(n27807) );
  XNOR U28491 ( .A(n27807), .B(sreg[1691]), .Z(n27809) );
  NAND U28492 ( .A(n27766), .B(sreg[1690]), .Z(n27770) );
  OR U28493 ( .A(n27768), .B(n27767), .Z(n27769) );
  AND U28494 ( .A(n27770), .B(n27769), .Z(n27808) );
  XOR U28495 ( .A(n27809), .B(n27808), .Z(c[1691]) );
  NANDN U28496 ( .A(n27772), .B(n27771), .Z(n27776) );
  NAND U28497 ( .A(n27774), .B(n27773), .Z(n27775) );
  NAND U28498 ( .A(n27776), .B(n27775), .Z(n27815) );
  NAND U28499 ( .A(b[0]), .B(a[676]), .Z(n27777) );
  XNOR U28500 ( .A(b[1]), .B(n27777), .Z(n27779) );
  NAND U28501 ( .A(n111), .B(a[675]), .Z(n27778) );
  AND U28502 ( .A(n27779), .B(n27778), .Z(n27832) );
  XOR U28503 ( .A(a[672]), .B(n42197), .Z(n27821) );
  NANDN U28504 ( .A(n27821), .B(n42173), .Z(n27782) );
  NANDN U28505 ( .A(n27780), .B(n42172), .Z(n27781) );
  NAND U28506 ( .A(n27782), .B(n27781), .Z(n27830) );
  NAND U28507 ( .A(b[7]), .B(a[668]), .Z(n27831) );
  XNOR U28508 ( .A(n27830), .B(n27831), .Z(n27833) );
  XOR U28509 ( .A(n27832), .B(n27833), .Z(n27839) );
  NANDN U28510 ( .A(n27783), .B(n42093), .Z(n27785) );
  XOR U28511 ( .A(n42134), .B(a[674]), .Z(n27824) );
  NANDN U28512 ( .A(n27824), .B(n42095), .Z(n27784) );
  NAND U28513 ( .A(n27785), .B(n27784), .Z(n27837) );
  NANDN U28514 ( .A(n27786), .B(n42231), .Z(n27788) );
  XOR U28515 ( .A(n217), .B(a[670]), .Z(n27827) );
  NANDN U28516 ( .A(n27827), .B(n42234), .Z(n27787) );
  AND U28517 ( .A(n27788), .B(n27787), .Z(n27836) );
  XNOR U28518 ( .A(n27837), .B(n27836), .Z(n27838) );
  XNOR U28519 ( .A(n27839), .B(n27838), .Z(n27843) );
  NANDN U28520 ( .A(n27790), .B(n27789), .Z(n27794) );
  NAND U28521 ( .A(n27792), .B(n27791), .Z(n27793) );
  AND U28522 ( .A(n27794), .B(n27793), .Z(n27842) );
  XOR U28523 ( .A(n27843), .B(n27842), .Z(n27844) );
  NANDN U28524 ( .A(n27796), .B(n27795), .Z(n27800) );
  NANDN U28525 ( .A(n27798), .B(n27797), .Z(n27799) );
  NAND U28526 ( .A(n27800), .B(n27799), .Z(n27845) );
  XOR U28527 ( .A(n27844), .B(n27845), .Z(n27812) );
  OR U28528 ( .A(n27802), .B(n27801), .Z(n27806) );
  NANDN U28529 ( .A(n27804), .B(n27803), .Z(n27805) );
  NAND U28530 ( .A(n27806), .B(n27805), .Z(n27813) );
  XNOR U28531 ( .A(n27812), .B(n27813), .Z(n27814) );
  XNOR U28532 ( .A(n27815), .B(n27814), .Z(n27848) );
  XNOR U28533 ( .A(n27848), .B(sreg[1692]), .Z(n27850) );
  NAND U28534 ( .A(n27807), .B(sreg[1691]), .Z(n27811) );
  OR U28535 ( .A(n27809), .B(n27808), .Z(n27810) );
  AND U28536 ( .A(n27811), .B(n27810), .Z(n27849) );
  XOR U28537 ( .A(n27850), .B(n27849), .Z(c[1692]) );
  NANDN U28538 ( .A(n27813), .B(n27812), .Z(n27817) );
  NAND U28539 ( .A(n27815), .B(n27814), .Z(n27816) );
  NAND U28540 ( .A(n27817), .B(n27816), .Z(n27856) );
  NAND U28541 ( .A(b[0]), .B(a[677]), .Z(n27818) );
  XNOR U28542 ( .A(b[1]), .B(n27818), .Z(n27820) );
  NAND U28543 ( .A(n111), .B(a[676]), .Z(n27819) );
  AND U28544 ( .A(n27820), .B(n27819), .Z(n27873) );
  XOR U28545 ( .A(a[673]), .B(n42197), .Z(n27862) );
  NANDN U28546 ( .A(n27862), .B(n42173), .Z(n27823) );
  NANDN U28547 ( .A(n27821), .B(n42172), .Z(n27822) );
  NAND U28548 ( .A(n27823), .B(n27822), .Z(n27871) );
  NAND U28549 ( .A(b[7]), .B(a[669]), .Z(n27872) );
  XNOR U28550 ( .A(n27871), .B(n27872), .Z(n27874) );
  XOR U28551 ( .A(n27873), .B(n27874), .Z(n27880) );
  NANDN U28552 ( .A(n27824), .B(n42093), .Z(n27826) );
  XOR U28553 ( .A(n42134), .B(a[675]), .Z(n27865) );
  NANDN U28554 ( .A(n27865), .B(n42095), .Z(n27825) );
  NAND U28555 ( .A(n27826), .B(n27825), .Z(n27878) );
  NANDN U28556 ( .A(n27827), .B(n42231), .Z(n27829) );
  XOR U28557 ( .A(n218), .B(a[671]), .Z(n27868) );
  NANDN U28558 ( .A(n27868), .B(n42234), .Z(n27828) );
  AND U28559 ( .A(n27829), .B(n27828), .Z(n27877) );
  XNOR U28560 ( .A(n27878), .B(n27877), .Z(n27879) );
  XNOR U28561 ( .A(n27880), .B(n27879), .Z(n27884) );
  NANDN U28562 ( .A(n27831), .B(n27830), .Z(n27835) );
  NAND U28563 ( .A(n27833), .B(n27832), .Z(n27834) );
  AND U28564 ( .A(n27835), .B(n27834), .Z(n27883) );
  XOR U28565 ( .A(n27884), .B(n27883), .Z(n27885) );
  NANDN U28566 ( .A(n27837), .B(n27836), .Z(n27841) );
  NANDN U28567 ( .A(n27839), .B(n27838), .Z(n27840) );
  NAND U28568 ( .A(n27841), .B(n27840), .Z(n27886) );
  XOR U28569 ( .A(n27885), .B(n27886), .Z(n27853) );
  OR U28570 ( .A(n27843), .B(n27842), .Z(n27847) );
  NANDN U28571 ( .A(n27845), .B(n27844), .Z(n27846) );
  NAND U28572 ( .A(n27847), .B(n27846), .Z(n27854) );
  XNOR U28573 ( .A(n27853), .B(n27854), .Z(n27855) );
  XNOR U28574 ( .A(n27856), .B(n27855), .Z(n27889) );
  XNOR U28575 ( .A(n27889), .B(sreg[1693]), .Z(n27891) );
  NAND U28576 ( .A(n27848), .B(sreg[1692]), .Z(n27852) );
  OR U28577 ( .A(n27850), .B(n27849), .Z(n27851) );
  AND U28578 ( .A(n27852), .B(n27851), .Z(n27890) );
  XOR U28579 ( .A(n27891), .B(n27890), .Z(c[1693]) );
  NANDN U28580 ( .A(n27854), .B(n27853), .Z(n27858) );
  NAND U28581 ( .A(n27856), .B(n27855), .Z(n27857) );
  NAND U28582 ( .A(n27858), .B(n27857), .Z(n27897) );
  NAND U28583 ( .A(b[0]), .B(a[678]), .Z(n27859) );
  XNOR U28584 ( .A(b[1]), .B(n27859), .Z(n27861) );
  NAND U28585 ( .A(n111), .B(a[677]), .Z(n27860) );
  AND U28586 ( .A(n27861), .B(n27860), .Z(n27914) );
  XOR U28587 ( .A(a[674]), .B(n42197), .Z(n27903) );
  NANDN U28588 ( .A(n27903), .B(n42173), .Z(n27864) );
  NANDN U28589 ( .A(n27862), .B(n42172), .Z(n27863) );
  NAND U28590 ( .A(n27864), .B(n27863), .Z(n27912) );
  NAND U28591 ( .A(b[7]), .B(a[670]), .Z(n27913) );
  XNOR U28592 ( .A(n27912), .B(n27913), .Z(n27915) );
  XOR U28593 ( .A(n27914), .B(n27915), .Z(n27921) );
  NANDN U28594 ( .A(n27865), .B(n42093), .Z(n27867) );
  XOR U28595 ( .A(n42134), .B(a[676]), .Z(n27906) );
  NANDN U28596 ( .A(n27906), .B(n42095), .Z(n27866) );
  NAND U28597 ( .A(n27867), .B(n27866), .Z(n27919) );
  NANDN U28598 ( .A(n27868), .B(n42231), .Z(n27870) );
  XOR U28599 ( .A(n218), .B(a[672]), .Z(n27909) );
  NANDN U28600 ( .A(n27909), .B(n42234), .Z(n27869) );
  AND U28601 ( .A(n27870), .B(n27869), .Z(n27918) );
  XNOR U28602 ( .A(n27919), .B(n27918), .Z(n27920) );
  XNOR U28603 ( .A(n27921), .B(n27920), .Z(n27925) );
  NANDN U28604 ( .A(n27872), .B(n27871), .Z(n27876) );
  NAND U28605 ( .A(n27874), .B(n27873), .Z(n27875) );
  AND U28606 ( .A(n27876), .B(n27875), .Z(n27924) );
  XOR U28607 ( .A(n27925), .B(n27924), .Z(n27926) );
  NANDN U28608 ( .A(n27878), .B(n27877), .Z(n27882) );
  NANDN U28609 ( .A(n27880), .B(n27879), .Z(n27881) );
  NAND U28610 ( .A(n27882), .B(n27881), .Z(n27927) );
  XOR U28611 ( .A(n27926), .B(n27927), .Z(n27894) );
  OR U28612 ( .A(n27884), .B(n27883), .Z(n27888) );
  NANDN U28613 ( .A(n27886), .B(n27885), .Z(n27887) );
  NAND U28614 ( .A(n27888), .B(n27887), .Z(n27895) );
  XNOR U28615 ( .A(n27894), .B(n27895), .Z(n27896) );
  XNOR U28616 ( .A(n27897), .B(n27896), .Z(n27930) );
  XNOR U28617 ( .A(n27930), .B(sreg[1694]), .Z(n27932) );
  NAND U28618 ( .A(n27889), .B(sreg[1693]), .Z(n27893) );
  OR U28619 ( .A(n27891), .B(n27890), .Z(n27892) );
  AND U28620 ( .A(n27893), .B(n27892), .Z(n27931) );
  XOR U28621 ( .A(n27932), .B(n27931), .Z(c[1694]) );
  NANDN U28622 ( .A(n27895), .B(n27894), .Z(n27899) );
  NAND U28623 ( .A(n27897), .B(n27896), .Z(n27898) );
  NAND U28624 ( .A(n27899), .B(n27898), .Z(n27938) );
  NAND U28625 ( .A(b[0]), .B(a[679]), .Z(n27900) );
  XNOR U28626 ( .A(b[1]), .B(n27900), .Z(n27902) );
  NAND U28627 ( .A(n112), .B(a[678]), .Z(n27901) );
  AND U28628 ( .A(n27902), .B(n27901), .Z(n27955) );
  XOR U28629 ( .A(a[675]), .B(n42197), .Z(n27944) );
  NANDN U28630 ( .A(n27944), .B(n42173), .Z(n27905) );
  NANDN U28631 ( .A(n27903), .B(n42172), .Z(n27904) );
  NAND U28632 ( .A(n27905), .B(n27904), .Z(n27953) );
  NAND U28633 ( .A(b[7]), .B(a[671]), .Z(n27954) );
  XNOR U28634 ( .A(n27953), .B(n27954), .Z(n27956) );
  XOR U28635 ( .A(n27955), .B(n27956), .Z(n27962) );
  NANDN U28636 ( .A(n27906), .B(n42093), .Z(n27908) );
  XOR U28637 ( .A(n42134), .B(a[677]), .Z(n27947) );
  NANDN U28638 ( .A(n27947), .B(n42095), .Z(n27907) );
  NAND U28639 ( .A(n27908), .B(n27907), .Z(n27960) );
  NANDN U28640 ( .A(n27909), .B(n42231), .Z(n27911) );
  XOR U28641 ( .A(n218), .B(a[673]), .Z(n27950) );
  NANDN U28642 ( .A(n27950), .B(n42234), .Z(n27910) );
  AND U28643 ( .A(n27911), .B(n27910), .Z(n27959) );
  XNOR U28644 ( .A(n27960), .B(n27959), .Z(n27961) );
  XNOR U28645 ( .A(n27962), .B(n27961), .Z(n27966) );
  NANDN U28646 ( .A(n27913), .B(n27912), .Z(n27917) );
  NAND U28647 ( .A(n27915), .B(n27914), .Z(n27916) );
  AND U28648 ( .A(n27917), .B(n27916), .Z(n27965) );
  XOR U28649 ( .A(n27966), .B(n27965), .Z(n27967) );
  NANDN U28650 ( .A(n27919), .B(n27918), .Z(n27923) );
  NANDN U28651 ( .A(n27921), .B(n27920), .Z(n27922) );
  NAND U28652 ( .A(n27923), .B(n27922), .Z(n27968) );
  XOR U28653 ( .A(n27967), .B(n27968), .Z(n27935) );
  OR U28654 ( .A(n27925), .B(n27924), .Z(n27929) );
  NANDN U28655 ( .A(n27927), .B(n27926), .Z(n27928) );
  NAND U28656 ( .A(n27929), .B(n27928), .Z(n27936) );
  XNOR U28657 ( .A(n27935), .B(n27936), .Z(n27937) );
  XNOR U28658 ( .A(n27938), .B(n27937), .Z(n27971) );
  XNOR U28659 ( .A(n27971), .B(sreg[1695]), .Z(n27973) );
  NAND U28660 ( .A(n27930), .B(sreg[1694]), .Z(n27934) );
  OR U28661 ( .A(n27932), .B(n27931), .Z(n27933) );
  AND U28662 ( .A(n27934), .B(n27933), .Z(n27972) );
  XOR U28663 ( .A(n27973), .B(n27972), .Z(c[1695]) );
  NANDN U28664 ( .A(n27936), .B(n27935), .Z(n27940) );
  NAND U28665 ( .A(n27938), .B(n27937), .Z(n27939) );
  NAND U28666 ( .A(n27940), .B(n27939), .Z(n27979) );
  NAND U28667 ( .A(b[0]), .B(a[680]), .Z(n27941) );
  XNOR U28668 ( .A(b[1]), .B(n27941), .Z(n27943) );
  NAND U28669 ( .A(n112), .B(a[679]), .Z(n27942) );
  AND U28670 ( .A(n27943), .B(n27942), .Z(n27996) );
  XOR U28671 ( .A(a[676]), .B(n42197), .Z(n27985) );
  NANDN U28672 ( .A(n27985), .B(n42173), .Z(n27946) );
  NANDN U28673 ( .A(n27944), .B(n42172), .Z(n27945) );
  NAND U28674 ( .A(n27946), .B(n27945), .Z(n27994) );
  NAND U28675 ( .A(b[7]), .B(a[672]), .Z(n27995) );
  XNOR U28676 ( .A(n27994), .B(n27995), .Z(n27997) );
  XOR U28677 ( .A(n27996), .B(n27997), .Z(n28003) );
  NANDN U28678 ( .A(n27947), .B(n42093), .Z(n27949) );
  XOR U28679 ( .A(n42134), .B(a[678]), .Z(n27988) );
  NANDN U28680 ( .A(n27988), .B(n42095), .Z(n27948) );
  NAND U28681 ( .A(n27949), .B(n27948), .Z(n28001) );
  NANDN U28682 ( .A(n27950), .B(n42231), .Z(n27952) );
  XOR U28683 ( .A(n218), .B(a[674]), .Z(n27991) );
  NANDN U28684 ( .A(n27991), .B(n42234), .Z(n27951) );
  AND U28685 ( .A(n27952), .B(n27951), .Z(n28000) );
  XNOR U28686 ( .A(n28001), .B(n28000), .Z(n28002) );
  XNOR U28687 ( .A(n28003), .B(n28002), .Z(n28007) );
  NANDN U28688 ( .A(n27954), .B(n27953), .Z(n27958) );
  NAND U28689 ( .A(n27956), .B(n27955), .Z(n27957) );
  AND U28690 ( .A(n27958), .B(n27957), .Z(n28006) );
  XOR U28691 ( .A(n28007), .B(n28006), .Z(n28008) );
  NANDN U28692 ( .A(n27960), .B(n27959), .Z(n27964) );
  NANDN U28693 ( .A(n27962), .B(n27961), .Z(n27963) );
  NAND U28694 ( .A(n27964), .B(n27963), .Z(n28009) );
  XOR U28695 ( .A(n28008), .B(n28009), .Z(n27976) );
  OR U28696 ( .A(n27966), .B(n27965), .Z(n27970) );
  NANDN U28697 ( .A(n27968), .B(n27967), .Z(n27969) );
  NAND U28698 ( .A(n27970), .B(n27969), .Z(n27977) );
  XNOR U28699 ( .A(n27976), .B(n27977), .Z(n27978) );
  XNOR U28700 ( .A(n27979), .B(n27978), .Z(n28012) );
  XNOR U28701 ( .A(n28012), .B(sreg[1696]), .Z(n28014) );
  NAND U28702 ( .A(n27971), .B(sreg[1695]), .Z(n27975) );
  OR U28703 ( .A(n27973), .B(n27972), .Z(n27974) );
  AND U28704 ( .A(n27975), .B(n27974), .Z(n28013) );
  XOR U28705 ( .A(n28014), .B(n28013), .Z(c[1696]) );
  NANDN U28706 ( .A(n27977), .B(n27976), .Z(n27981) );
  NAND U28707 ( .A(n27979), .B(n27978), .Z(n27980) );
  NAND U28708 ( .A(n27981), .B(n27980), .Z(n28020) );
  NAND U28709 ( .A(b[0]), .B(a[681]), .Z(n27982) );
  XNOR U28710 ( .A(b[1]), .B(n27982), .Z(n27984) );
  NAND U28711 ( .A(n112), .B(a[680]), .Z(n27983) );
  AND U28712 ( .A(n27984), .B(n27983), .Z(n28037) );
  XOR U28713 ( .A(a[677]), .B(n42197), .Z(n28026) );
  NANDN U28714 ( .A(n28026), .B(n42173), .Z(n27987) );
  NANDN U28715 ( .A(n27985), .B(n42172), .Z(n27986) );
  NAND U28716 ( .A(n27987), .B(n27986), .Z(n28035) );
  NAND U28717 ( .A(b[7]), .B(a[673]), .Z(n28036) );
  XNOR U28718 ( .A(n28035), .B(n28036), .Z(n28038) );
  XOR U28719 ( .A(n28037), .B(n28038), .Z(n28044) );
  NANDN U28720 ( .A(n27988), .B(n42093), .Z(n27990) );
  XOR U28721 ( .A(n42134), .B(a[679]), .Z(n28029) );
  NANDN U28722 ( .A(n28029), .B(n42095), .Z(n27989) );
  NAND U28723 ( .A(n27990), .B(n27989), .Z(n28042) );
  NANDN U28724 ( .A(n27991), .B(n42231), .Z(n27993) );
  XOR U28725 ( .A(n218), .B(a[675]), .Z(n28032) );
  NANDN U28726 ( .A(n28032), .B(n42234), .Z(n27992) );
  AND U28727 ( .A(n27993), .B(n27992), .Z(n28041) );
  XNOR U28728 ( .A(n28042), .B(n28041), .Z(n28043) );
  XNOR U28729 ( .A(n28044), .B(n28043), .Z(n28048) );
  NANDN U28730 ( .A(n27995), .B(n27994), .Z(n27999) );
  NAND U28731 ( .A(n27997), .B(n27996), .Z(n27998) );
  AND U28732 ( .A(n27999), .B(n27998), .Z(n28047) );
  XOR U28733 ( .A(n28048), .B(n28047), .Z(n28049) );
  NANDN U28734 ( .A(n28001), .B(n28000), .Z(n28005) );
  NANDN U28735 ( .A(n28003), .B(n28002), .Z(n28004) );
  NAND U28736 ( .A(n28005), .B(n28004), .Z(n28050) );
  XOR U28737 ( .A(n28049), .B(n28050), .Z(n28017) );
  OR U28738 ( .A(n28007), .B(n28006), .Z(n28011) );
  NANDN U28739 ( .A(n28009), .B(n28008), .Z(n28010) );
  NAND U28740 ( .A(n28011), .B(n28010), .Z(n28018) );
  XNOR U28741 ( .A(n28017), .B(n28018), .Z(n28019) );
  XNOR U28742 ( .A(n28020), .B(n28019), .Z(n28053) );
  XNOR U28743 ( .A(n28053), .B(sreg[1697]), .Z(n28055) );
  NAND U28744 ( .A(n28012), .B(sreg[1696]), .Z(n28016) );
  OR U28745 ( .A(n28014), .B(n28013), .Z(n28015) );
  AND U28746 ( .A(n28016), .B(n28015), .Z(n28054) );
  XOR U28747 ( .A(n28055), .B(n28054), .Z(c[1697]) );
  NANDN U28748 ( .A(n28018), .B(n28017), .Z(n28022) );
  NAND U28749 ( .A(n28020), .B(n28019), .Z(n28021) );
  NAND U28750 ( .A(n28022), .B(n28021), .Z(n28061) );
  NAND U28751 ( .A(b[0]), .B(a[682]), .Z(n28023) );
  XNOR U28752 ( .A(b[1]), .B(n28023), .Z(n28025) );
  NAND U28753 ( .A(n112), .B(a[681]), .Z(n28024) );
  AND U28754 ( .A(n28025), .B(n28024), .Z(n28078) );
  XOR U28755 ( .A(a[678]), .B(n42197), .Z(n28067) );
  NANDN U28756 ( .A(n28067), .B(n42173), .Z(n28028) );
  NANDN U28757 ( .A(n28026), .B(n42172), .Z(n28027) );
  NAND U28758 ( .A(n28028), .B(n28027), .Z(n28076) );
  NAND U28759 ( .A(b[7]), .B(a[674]), .Z(n28077) );
  XNOR U28760 ( .A(n28076), .B(n28077), .Z(n28079) );
  XOR U28761 ( .A(n28078), .B(n28079), .Z(n28085) );
  NANDN U28762 ( .A(n28029), .B(n42093), .Z(n28031) );
  XOR U28763 ( .A(n42134), .B(a[680]), .Z(n28070) );
  NANDN U28764 ( .A(n28070), .B(n42095), .Z(n28030) );
  NAND U28765 ( .A(n28031), .B(n28030), .Z(n28083) );
  NANDN U28766 ( .A(n28032), .B(n42231), .Z(n28034) );
  XOR U28767 ( .A(n218), .B(a[676]), .Z(n28073) );
  NANDN U28768 ( .A(n28073), .B(n42234), .Z(n28033) );
  AND U28769 ( .A(n28034), .B(n28033), .Z(n28082) );
  XNOR U28770 ( .A(n28083), .B(n28082), .Z(n28084) );
  XNOR U28771 ( .A(n28085), .B(n28084), .Z(n28089) );
  NANDN U28772 ( .A(n28036), .B(n28035), .Z(n28040) );
  NAND U28773 ( .A(n28038), .B(n28037), .Z(n28039) );
  AND U28774 ( .A(n28040), .B(n28039), .Z(n28088) );
  XOR U28775 ( .A(n28089), .B(n28088), .Z(n28090) );
  NANDN U28776 ( .A(n28042), .B(n28041), .Z(n28046) );
  NANDN U28777 ( .A(n28044), .B(n28043), .Z(n28045) );
  NAND U28778 ( .A(n28046), .B(n28045), .Z(n28091) );
  XOR U28779 ( .A(n28090), .B(n28091), .Z(n28058) );
  OR U28780 ( .A(n28048), .B(n28047), .Z(n28052) );
  NANDN U28781 ( .A(n28050), .B(n28049), .Z(n28051) );
  NAND U28782 ( .A(n28052), .B(n28051), .Z(n28059) );
  XNOR U28783 ( .A(n28058), .B(n28059), .Z(n28060) );
  XNOR U28784 ( .A(n28061), .B(n28060), .Z(n28094) );
  XNOR U28785 ( .A(n28094), .B(sreg[1698]), .Z(n28096) );
  NAND U28786 ( .A(n28053), .B(sreg[1697]), .Z(n28057) );
  OR U28787 ( .A(n28055), .B(n28054), .Z(n28056) );
  AND U28788 ( .A(n28057), .B(n28056), .Z(n28095) );
  XOR U28789 ( .A(n28096), .B(n28095), .Z(c[1698]) );
  NANDN U28790 ( .A(n28059), .B(n28058), .Z(n28063) );
  NAND U28791 ( .A(n28061), .B(n28060), .Z(n28062) );
  NAND U28792 ( .A(n28063), .B(n28062), .Z(n28102) );
  NAND U28793 ( .A(b[0]), .B(a[683]), .Z(n28064) );
  XNOR U28794 ( .A(b[1]), .B(n28064), .Z(n28066) );
  NAND U28795 ( .A(n112), .B(a[682]), .Z(n28065) );
  AND U28796 ( .A(n28066), .B(n28065), .Z(n28119) );
  XOR U28797 ( .A(a[679]), .B(n42197), .Z(n28108) );
  NANDN U28798 ( .A(n28108), .B(n42173), .Z(n28069) );
  NANDN U28799 ( .A(n28067), .B(n42172), .Z(n28068) );
  NAND U28800 ( .A(n28069), .B(n28068), .Z(n28117) );
  NAND U28801 ( .A(b[7]), .B(a[675]), .Z(n28118) );
  XNOR U28802 ( .A(n28117), .B(n28118), .Z(n28120) );
  XOR U28803 ( .A(n28119), .B(n28120), .Z(n28126) );
  NANDN U28804 ( .A(n28070), .B(n42093), .Z(n28072) );
  XOR U28805 ( .A(n42134), .B(a[681]), .Z(n28111) );
  NANDN U28806 ( .A(n28111), .B(n42095), .Z(n28071) );
  NAND U28807 ( .A(n28072), .B(n28071), .Z(n28124) );
  NANDN U28808 ( .A(n28073), .B(n42231), .Z(n28075) );
  XOR U28809 ( .A(n218), .B(a[677]), .Z(n28114) );
  NANDN U28810 ( .A(n28114), .B(n42234), .Z(n28074) );
  AND U28811 ( .A(n28075), .B(n28074), .Z(n28123) );
  XNOR U28812 ( .A(n28124), .B(n28123), .Z(n28125) );
  XNOR U28813 ( .A(n28126), .B(n28125), .Z(n28130) );
  NANDN U28814 ( .A(n28077), .B(n28076), .Z(n28081) );
  NAND U28815 ( .A(n28079), .B(n28078), .Z(n28080) );
  AND U28816 ( .A(n28081), .B(n28080), .Z(n28129) );
  XOR U28817 ( .A(n28130), .B(n28129), .Z(n28131) );
  NANDN U28818 ( .A(n28083), .B(n28082), .Z(n28087) );
  NANDN U28819 ( .A(n28085), .B(n28084), .Z(n28086) );
  NAND U28820 ( .A(n28087), .B(n28086), .Z(n28132) );
  XOR U28821 ( .A(n28131), .B(n28132), .Z(n28099) );
  OR U28822 ( .A(n28089), .B(n28088), .Z(n28093) );
  NANDN U28823 ( .A(n28091), .B(n28090), .Z(n28092) );
  NAND U28824 ( .A(n28093), .B(n28092), .Z(n28100) );
  XNOR U28825 ( .A(n28099), .B(n28100), .Z(n28101) );
  XNOR U28826 ( .A(n28102), .B(n28101), .Z(n28135) );
  XNOR U28827 ( .A(n28135), .B(sreg[1699]), .Z(n28137) );
  NAND U28828 ( .A(n28094), .B(sreg[1698]), .Z(n28098) );
  OR U28829 ( .A(n28096), .B(n28095), .Z(n28097) );
  AND U28830 ( .A(n28098), .B(n28097), .Z(n28136) );
  XOR U28831 ( .A(n28137), .B(n28136), .Z(c[1699]) );
  NANDN U28832 ( .A(n28100), .B(n28099), .Z(n28104) );
  NAND U28833 ( .A(n28102), .B(n28101), .Z(n28103) );
  NAND U28834 ( .A(n28104), .B(n28103), .Z(n28143) );
  NAND U28835 ( .A(b[0]), .B(a[684]), .Z(n28105) );
  XNOR U28836 ( .A(b[1]), .B(n28105), .Z(n28107) );
  NAND U28837 ( .A(n112), .B(a[683]), .Z(n28106) );
  AND U28838 ( .A(n28107), .B(n28106), .Z(n28160) );
  XOR U28839 ( .A(a[680]), .B(n42197), .Z(n28149) );
  NANDN U28840 ( .A(n28149), .B(n42173), .Z(n28110) );
  NANDN U28841 ( .A(n28108), .B(n42172), .Z(n28109) );
  NAND U28842 ( .A(n28110), .B(n28109), .Z(n28158) );
  NAND U28843 ( .A(b[7]), .B(a[676]), .Z(n28159) );
  XNOR U28844 ( .A(n28158), .B(n28159), .Z(n28161) );
  XOR U28845 ( .A(n28160), .B(n28161), .Z(n28167) );
  NANDN U28846 ( .A(n28111), .B(n42093), .Z(n28113) );
  XOR U28847 ( .A(n42134), .B(a[682]), .Z(n28152) );
  NANDN U28848 ( .A(n28152), .B(n42095), .Z(n28112) );
  NAND U28849 ( .A(n28113), .B(n28112), .Z(n28165) );
  NANDN U28850 ( .A(n28114), .B(n42231), .Z(n28116) );
  XOR U28851 ( .A(n218), .B(a[678]), .Z(n28155) );
  NANDN U28852 ( .A(n28155), .B(n42234), .Z(n28115) );
  AND U28853 ( .A(n28116), .B(n28115), .Z(n28164) );
  XNOR U28854 ( .A(n28165), .B(n28164), .Z(n28166) );
  XNOR U28855 ( .A(n28167), .B(n28166), .Z(n28171) );
  NANDN U28856 ( .A(n28118), .B(n28117), .Z(n28122) );
  NAND U28857 ( .A(n28120), .B(n28119), .Z(n28121) );
  AND U28858 ( .A(n28122), .B(n28121), .Z(n28170) );
  XOR U28859 ( .A(n28171), .B(n28170), .Z(n28172) );
  NANDN U28860 ( .A(n28124), .B(n28123), .Z(n28128) );
  NANDN U28861 ( .A(n28126), .B(n28125), .Z(n28127) );
  NAND U28862 ( .A(n28128), .B(n28127), .Z(n28173) );
  XOR U28863 ( .A(n28172), .B(n28173), .Z(n28140) );
  OR U28864 ( .A(n28130), .B(n28129), .Z(n28134) );
  NANDN U28865 ( .A(n28132), .B(n28131), .Z(n28133) );
  NAND U28866 ( .A(n28134), .B(n28133), .Z(n28141) );
  XNOR U28867 ( .A(n28140), .B(n28141), .Z(n28142) );
  XNOR U28868 ( .A(n28143), .B(n28142), .Z(n28176) );
  XNOR U28869 ( .A(n28176), .B(sreg[1700]), .Z(n28178) );
  NAND U28870 ( .A(n28135), .B(sreg[1699]), .Z(n28139) );
  OR U28871 ( .A(n28137), .B(n28136), .Z(n28138) );
  AND U28872 ( .A(n28139), .B(n28138), .Z(n28177) );
  XOR U28873 ( .A(n28178), .B(n28177), .Z(c[1700]) );
  NANDN U28874 ( .A(n28141), .B(n28140), .Z(n28145) );
  NAND U28875 ( .A(n28143), .B(n28142), .Z(n28144) );
  NAND U28876 ( .A(n28145), .B(n28144), .Z(n28184) );
  NAND U28877 ( .A(b[0]), .B(a[685]), .Z(n28146) );
  XNOR U28878 ( .A(b[1]), .B(n28146), .Z(n28148) );
  NAND U28879 ( .A(n112), .B(a[684]), .Z(n28147) );
  AND U28880 ( .A(n28148), .B(n28147), .Z(n28201) );
  XOR U28881 ( .A(a[681]), .B(n42197), .Z(n28190) );
  NANDN U28882 ( .A(n28190), .B(n42173), .Z(n28151) );
  NANDN U28883 ( .A(n28149), .B(n42172), .Z(n28150) );
  NAND U28884 ( .A(n28151), .B(n28150), .Z(n28199) );
  NAND U28885 ( .A(b[7]), .B(a[677]), .Z(n28200) );
  XNOR U28886 ( .A(n28199), .B(n28200), .Z(n28202) );
  XOR U28887 ( .A(n28201), .B(n28202), .Z(n28208) );
  NANDN U28888 ( .A(n28152), .B(n42093), .Z(n28154) );
  XOR U28889 ( .A(n42134), .B(a[683]), .Z(n28193) );
  NANDN U28890 ( .A(n28193), .B(n42095), .Z(n28153) );
  NAND U28891 ( .A(n28154), .B(n28153), .Z(n28206) );
  NANDN U28892 ( .A(n28155), .B(n42231), .Z(n28157) );
  XOR U28893 ( .A(n218), .B(a[679]), .Z(n28196) );
  NANDN U28894 ( .A(n28196), .B(n42234), .Z(n28156) );
  AND U28895 ( .A(n28157), .B(n28156), .Z(n28205) );
  XNOR U28896 ( .A(n28206), .B(n28205), .Z(n28207) );
  XNOR U28897 ( .A(n28208), .B(n28207), .Z(n28212) );
  NANDN U28898 ( .A(n28159), .B(n28158), .Z(n28163) );
  NAND U28899 ( .A(n28161), .B(n28160), .Z(n28162) );
  AND U28900 ( .A(n28163), .B(n28162), .Z(n28211) );
  XOR U28901 ( .A(n28212), .B(n28211), .Z(n28213) );
  NANDN U28902 ( .A(n28165), .B(n28164), .Z(n28169) );
  NANDN U28903 ( .A(n28167), .B(n28166), .Z(n28168) );
  NAND U28904 ( .A(n28169), .B(n28168), .Z(n28214) );
  XOR U28905 ( .A(n28213), .B(n28214), .Z(n28181) );
  OR U28906 ( .A(n28171), .B(n28170), .Z(n28175) );
  NANDN U28907 ( .A(n28173), .B(n28172), .Z(n28174) );
  NAND U28908 ( .A(n28175), .B(n28174), .Z(n28182) );
  XNOR U28909 ( .A(n28181), .B(n28182), .Z(n28183) );
  XNOR U28910 ( .A(n28184), .B(n28183), .Z(n28217) );
  XNOR U28911 ( .A(n28217), .B(sreg[1701]), .Z(n28219) );
  NAND U28912 ( .A(n28176), .B(sreg[1700]), .Z(n28180) );
  OR U28913 ( .A(n28178), .B(n28177), .Z(n28179) );
  AND U28914 ( .A(n28180), .B(n28179), .Z(n28218) );
  XOR U28915 ( .A(n28219), .B(n28218), .Z(c[1701]) );
  NANDN U28916 ( .A(n28182), .B(n28181), .Z(n28186) );
  NAND U28917 ( .A(n28184), .B(n28183), .Z(n28185) );
  NAND U28918 ( .A(n28186), .B(n28185), .Z(n28225) );
  NAND U28919 ( .A(b[0]), .B(a[686]), .Z(n28187) );
  XNOR U28920 ( .A(b[1]), .B(n28187), .Z(n28189) );
  NAND U28921 ( .A(n113), .B(a[685]), .Z(n28188) );
  AND U28922 ( .A(n28189), .B(n28188), .Z(n28242) );
  XOR U28923 ( .A(a[682]), .B(n42197), .Z(n28231) );
  NANDN U28924 ( .A(n28231), .B(n42173), .Z(n28192) );
  NANDN U28925 ( .A(n28190), .B(n42172), .Z(n28191) );
  NAND U28926 ( .A(n28192), .B(n28191), .Z(n28240) );
  NAND U28927 ( .A(b[7]), .B(a[678]), .Z(n28241) );
  XNOR U28928 ( .A(n28240), .B(n28241), .Z(n28243) );
  XOR U28929 ( .A(n28242), .B(n28243), .Z(n28249) );
  NANDN U28930 ( .A(n28193), .B(n42093), .Z(n28195) );
  XOR U28931 ( .A(n42134), .B(a[684]), .Z(n28234) );
  NANDN U28932 ( .A(n28234), .B(n42095), .Z(n28194) );
  NAND U28933 ( .A(n28195), .B(n28194), .Z(n28247) );
  NANDN U28934 ( .A(n28196), .B(n42231), .Z(n28198) );
  XOR U28935 ( .A(n218), .B(a[680]), .Z(n28237) );
  NANDN U28936 ( .A(n28237), .B(n42234), .Z(n28197) );
  AND U28937 ( .A(n28198), .B(n28197), .Z(n28246) );
  XNOR U28938 ( .A(n28247), .B(n28246), .Z(n28248) );
  XNOR U28939 ( .A(n28249), .B(n28248), .Z(n28253) );
  NANDN U28940 ( .A(n28200), .B(n28199), .Z(n28204) );
  NAND U28941 ( .A(n28202), .B(n28201), .Z(n28203) );
  AND U28942 ( .A(n28204), .B(n28203), .Z(n28252) );
  XOR U28943 ( .A(n28253), .B(n28252), .Z(n28254) );
  NANDN U28944 ( .A(n28206), .B(n28205), .Z(n28210) );
  NANDN U28945 ( .A(n28208), .B(n28207), .Z(n28209) );
  NAND U28946 ( .A(n28210), .B(n28209), .Z(n28255) );
  XOR U28947 ( .A(n28254), .B(n28255), .Z(n28222) );
  OR U28948 ( .A(n28212), .B(n28211), .Z(n28216) );
  NANDN U28949 ( .A(n28214), .B(n28213), .Z(n28215) );
  NAND U28950 ( .A(n28216), .B(n28215), .Z(n28223) );
  XNOR U28951 ( .A(n28222), .B(n28223), .Z(n28224) );
  XNOR U28952 ( .A(n28225), .B(n28224), .Z(n28258) );
  XNOR U28953 ( .A(n28258), .B(sreg[1702]), .Z(n28260) );
  NAND U28954 ( .A(n28217), .B(sreg[1701]), .Z(n28221) );
  OR U28955 ( .A(n28219), .B(n28218), .Z(n28220) );
  AND U28956 ( .A(n28221), .B(n28220), .Z(n28259) );
  XOR U28957 ( .A(n28260), .B(n28259), .Z(c[1702]) );
  NANDN U28958 ( .A(n28223), .B(n28222), .Z(n28227) );
  NAND U28959 ( .A(n28225), .B(n28224), .Z(n28226) );
  NAND U28960 ( .A(n28227), .B(n28226), .Z(n28266) );
  NAND U28961 ( .A(b[0]), .B(a[687]), .Z(n28228) );
  XNOR U28962 ( .A(b[1]), .B(n28228), .Z(n28230) );
  NAND U28963 ( .A(n113), .B(a[686]), .Z(n28229) );
  AND U28964 ( .A(n28230), .B(n28229), .Z(n28283) );
  XOR U28965 ( .A(a[683]), .B(n42197), .Z(n28272) );
  NANDN U28966 ( .A(n28272), .B(n42173), .Z(n28233) );
  NANDN U28967 ( .A(n28231), .B(n42172), .Z(n28232) );
  NAND U28968 ( .A(n28233), .B(n28232), .Z(n28281) );
  NAND U28969 ( .A(b[7]), .B(a[679]), .Z(n28282) );
  XNOR U28970 ( .A(n28281), .B(n28282), .Z(n28284) );
  XOR U28971 ( .A(n28283), .B(n28284), .Z(n28290) );
  NANDN U28972 ( .A(n28234), .B(n42093), .Z(n28236) );
  XOR U28973 ( .A(n42134), .B(a[685]), .Z(n28275) );
  NANDN U28974 ( .A(n28275), .B(n42095), .Z(n28235) );
  NAND U28975 ( .A(n28236), .B(n28235), .Z(n28288) );
  NANDN U28976 ( .A(n28237), .B(n42231), .Z(n28239) );
  XOR U28977 ( .A(n218), .B(a[681]), .Z(n28278) );
  NANDN U28978 ( .A(n28278), .B(n42234), .Z(n28238) );
  AND U28979 ( .A(n28239), .B(n28238), .Z(n28287) );
  XNOR U28980 ( .A(n28288), .B(n28287), .Z(n28289) );
  XNOR U28981 ( .A(n28290), .B(n28289), .Z(n28294) );
  NANDN U28982 ( .A(n28241), .B(n28240), .Z(n28245) );
  NAND U28983 ( .A(n28243), .B(n28242), .Z(n28244) );
  AND U28984 ( .A(n28245), .B(n28244), .Z(n28293) );
  XOR U28985 ( .A(n28294), .B(n28293), .Z(n28295) );
  NANDN U28986 ( .A(n28247), .B(n28246), .Z(n28251) );
  NANDN U28987 ( .A(n28249), .B(n28248), .Z(n28250) );
  NAND U28988 ( .A(n28251), .B(n28250), .Z(n28296) );
  XOR U28989 ( .A(n28295), .B(n28296), .Z(n28263) );
  OR U28990 ( .A(n28253), .B(n28252), .Z(n28257) );
  NANDN U28991 ( .A(n28255), .B(n28254), .Z(n28256) );
  NAND U28992 ( .A(n28257), .B(n28256), .Z(n28264) );
  XNOR U28993 ( .A(n28263), .B(n28264), .Z(n28265) );
  XNOR U28994 ( .A(n28266), .B(n28265), .Z(n28299) );
  XNOR U28995 ( .A(n28299), .B(sreg[1703]), .Z(n28301) );
  NAND U28996 ( .A(n28258), .B(sreg[1702]), .Z(n28262) );
  OR U28997 ( .A(n28260), .B(n28259), .Z(n28261) );
  AND U28998 ( .A(n28262), .B(n28261), .Z(n28300) );
  XOR U28999 ( .A(n28301), .B(n28300), .Z(c[1703]) );
  NANDN U29000 ( .A(n28264), .B(n28263), .Z(n28268) );
  NAND U29001 ( .A(n28266), .B(n28265), .Z(n28267) );
  NAND U29002 ( .A(n28268), .B(n28267), .Z(n28307) );
  NAND U29003 ( .A(b[0]), .B(a[688]), .Z(n28269) );
  XNOR U29004 ( .A(b[1]), .B(n28269), .Z(n28271) );
  NAND U29005 ( .A(n113), .B(a[687]), .Z(n28270) );
  AND U29006 ( .A(n28271), .B(n28270), .Z(n28324) );
  XOR U29007 ( .A(a[684]), .B(n42197), .Z(n28313) );
  NANDN U29008 ( .A(n28313), .B(n42173), .Z(n28274) );
  NANDN U29009 ( .A(n28272), .B(n42172), .Z(n28273) );
  NAND U29010 ( .A(n28274), .B(n28273), .Z(n28322) );
  NAND U29011 ( .A(b[7]), .B(a[680]), .Z(n28323) );
  XNOR U29012 ( .A(n28322), .B(n28323), .Z(n28325) );
  XOR U29013 ( .A(n28324), .B(n28325), .Z(n28331) );
  NANDN U29014 ( .A(n28275), .B(n42093), .Z(n28277) );
  XOR U29015 ( .A(n42134), .B(a[686]), .Z(n28316) );
  NANDN U29016 ( .A(n28316), .B(n42095), .Z(n28276) );
  NAND U29017 ( .A(n28277), .B(n28276), .Z(n28329) );
  NANDN U29018 ( .A(n28278), .B(n42231), .Z(n28280) );
  XOR U29019 ( .A(n218), .B(a[682]), .Z(n28319) );
  NANDN U29020 ( .A(n28319), .B(n42234), .Z(n28279) );
  AND U29021 ( .A(n28280), .B(n28279), .Z(n28328) );
  XNOR U29022 ( .A(n28329), .B(n28328), .Z(n28330) );
  XNOR U29023 ( .A(n28331), .B(n28330), .Z(n28335) );
  NANDN U29024 ( .A(n28282), .B(n28281), .Z(n28286) );
  NAND U29025 ( .A(n28284), .B(n28283), .Z(n28285) );
  AND U29026 ( .A(n28286), .B(n28285), .Z(n28334) );
  XOR U29027 ( .A(n28335), .B(n28334), .Z(n28336) );
  NANDN U29028 ( .A(n28288), .B(n28287), .Z(n28292) );
  NANDN U29029 ( .A(n28290), .B(n28289), .Z(n28291) );
  NAND U29030 ( .A(n28292), .B(n28291), .Z(n28337) );
  XOR U29031 ( .A(n28336), .B(n28337), .Z(n28304) );
  OR U29032 ( .A(n28294), .B(n28293), .Z(n28298) );
  NANDN U29033 ( .A(n28296), .B(n28295), .Z(n28297) );
  NAND U29034 ( .A(n28298), .B(n28297), .Z(n28305) );
  XNOR U29035 ( .A(n28304), .B(n28305), .Z(n28306) );
  XNOR U29036 ( .A(n28307), .B(n28306), .Z(n28340) );
  XNOR U29037 ( .A(n28340), .B(sreg[1704]), .Z(n28342) );
  NAND U29038 ( .A(n28299), .B(sreg[1703]), .Z(n28303) );
  OR U29039 ( .A(n28301), .B(n28300), .Z(n28302) );
  AND U29040 ( .A(n28303), .B(n28302), .Z(n28341) );
  XOR U29041 ( .A(n28342), .B(n28341), .Z(c[1704]) );
  NANDN U29042 ( .A(n28305), .B(n28304), .Z(n28309) );
  NAND U29043 ( .A(n28307), .B(n28306), .Z(n28308) );
  NAND U29044 ( .A(n28309), .B(n28308), .Z(n28348) );
  NAND U29045 ( .A(b[0]), .B(a[689]), .Z(n28310) );
  XNOR U29046 ( .A(b[1]), .B(n28310), .Z(n28312) );
  NAND U29047 ( .A(n113), .B(a[688]), .Z(n28311) );
  AND U29048 ( .A(n28312), .B(n28311), .Z(n28365) );
  XOR U29049 ( .A(a[685]), .B(n42197), .Z(n28354) );
  NANDN U29050 ( .A(n28354), .B(n42173), .Z(n28315) );
  NANDN U29051 ( .A(n28313), .B(n42172), .Z(n28314) );
  NAND U29052 ( .A(n28315), .B(n28314), .Z(n28363) );
  NAND U29053 ( .A(b[7]), .B(a[681]), .Z(n28364) );
  XNOR U29054 ( .A(n28363), .B(n28364), .Z(n28366) );
  XOR U29055 ( .A(n28365), .B(n28366), .Z(n28372) );
  NANDN U29056 ( .A(n28316), .B(n42093), .Z(n28318) );
  XOR U29057 ( .A(n42134), .B(a[687]), .Z(n28357) );
  NANDN U29058 ( .A(n28357), .B(n42095), .Z(n28317) );
  NAND U29059 ( .A(n28318), .B(n28317), .Z(n28370) );
  NANDN U29060 ( .A(n28319), .B(n42231), .Z(n28321) );
  XOR U29061 ( .A(n219), .B(a[683]), .Z(n28360) );
  NANDN U29062 ( .A(n28360), .B(n42234), .Z(n28320) );
  AND U29063 ( .A(n28321), .B(n28320), .Z(n28369) );
  XNOR U29064 ( .A(n28370), .B(n28369), .Z(n28371) );
  XNOR U29065 ( .A(n28372), .B(n28371), .Z(n28376) );
  NANDN U29066 ( .A(n28323), .B(n28322), .Z(n28327) );
  NAND U29067 ( .A(n28325), .B(n28324), .Z(n28326) );
  AND U29068 ( .A(n28327), .B(n28326), .Z(n28375) );
  XOR U29069 ( .A(n28376), .B(n28375), .Z(n28377) );
  NANDN U29070 ( .A(n28329), .B(n28328), .Z(n28333) );
  NANDN U29071 ( .A(n28331), .B(n28330), .Z(n28332) );
  NAND U29072 ( .A(n28333), .B(n28332), .Z(n28378) );
  XOR U29073 ( .A(n28377), .B(n28378), .Z(n28345) );
  OR U29074 ( .A(n28335), .B(n28334), .Z(n28339) );
  NANDN U29075 ( .A(n28337), .B(n28336), .Z(n28338) );
  NAND U29076 ( .A(n28339), .B(n28338), .Z(n28346) );
  XNOR U29077 ( .A(n28345), .B(n28346), .Z(n28347) );
  XNOR U29078 ( .A(n28348), .B(n28347), .Z(n28381) );
  XNOR U29079 ( .A(n28381), .B(sreg[1705]), .Z(n28383) );
  NAND U29080 ( .A(n28340), .B(sreg[1704]), .Z(n28344) );
  OR U29081 ( .A(n28342), .B(n28341), .Z(n28343) );
  AND U29082 ( .A(n28344), .B(n28343), .Z(n28382) );
  XOR U29083 ( .A(n28383), .B(n28382), .Z(c[1705]) );
  NANDN U29084 ( .A(n28346), .B(n28345), .Z(n28350) );
  NAND U29085 ( .A(n28348), .B(n28347), .Z(n28349) );
  NAND U29086 ( .A(n28350), .B(n28349), .Z(n28389) );
  NAND U29087 ( .A(b[0]), .B(a[690]), .Z(n28351) );
  XNOR U29088 ( .A(b[1]), .B(n28351), .Z(n28353) );
  NAND U29089 ( .A(n113), .B(a[689]), .Z(n28352) );
  AND U29090 ( .A(n28353), .B(n28352), .Z(n28406) );
  XOR U29091 ( .A(a[686]), .B(n42197), .Z(n28395) );
  NANDN U29092 ( .A(n28395), .B(n42173), .Z(n28356) );
  NANDN U29093 ( .A(n28354), .B(n42172), .Z(n28355) );
  NAND U29094 ( .A(n28356), .B(n28355), .Z(n28404) );
  NAND U29095 ( .A(b[7]), .B(a[682]), .Z(n28405) );
  XNOR U29096 ( .A(n28404), .B(n28405), .Z(n28407) );
  XOR U29097 ( .A(n28406), .B(n28407), .Z(n28413) );
  NANDN U29098 ( .A(n28357), .B(n42093), .Z(n28359) );
  XOR U29099 ( .A(n42134), .B(a[688]), .Z(n28398) );
  NANDN U29100 ( .A(n28398), .B(n42095), .Z(n28358) );
  NAND U29101 ( .A(n28359), .B(n28358), .Z(n28411) );
  NANDN U29102 ( .A(n28360), .B(n42231), .Z(n28362) );
  XOR U29103 ( .A(n219), .B(a[684]), .Z(n28401) );
  NANDN U29104 ( .A(n28401), .B(n42234), .Z(n28361) );
  AND U29105 ( .A(n28362), .B(n28361), .Z(n28410) );
  XNOR U29106 ( .A(n28411), .B(n28410), .Z(n28412) );
  XNOR U29107 ( .A(n28413), .B(n28412), .Z(n28417) );
  NANDN U29108 ( .A(n28364), .B(n28363), .Z(n28368) );
  NAND U29109 ( .A(n28366), .B(n28365), .Z(n28367) );
  AND U29110 ( .A(n28368), .B(n28367), .Z(n28416) );
  XOR U29111 ( .A(n28417), .B(n28416), .Z(n28418) );
  NANDN U29112 ( .A(n28370), .B(n28369), .Z(n28374) );
  NANDN U29113 ( .A(n28372), .B(n28371), .Z(n28373) );
  NAND U29114 ( .A(n28374), .B(n28373), .Z(n28419) );
  XOR U29115 ( .A(n28418), .B(n28419), .Z(n28386) );
  OR U29116 ( .A(n28376), .B(n28375), .Z(n28380) );
  NANDN U29117 ( .A(n28378), .B(n28377), .Z(n28379) );
  NAND U29118 ( .A(n28380), .B(n28379), .Z(n28387) );
  XNOR U29119 ( .A(n28386), .B(n28387), .Z(n28388) );
  XNOR U29120 ( .A(n28389), .B(n28388), .Z(n28422) );
  XNOR U29121 ( .A(n28422), .B(sreg[1706]), .Z(n28424) );
  NAND U29122 ( .A(n28381), .B(sreg[1705]), .Z(n28385) );
  OR U29123 ( .A(n28383), .B(n28382), .Z(n28384) );
  AND U29124 ( .A(n28385), .B(n28384), .Z(n28423) );
  XOR U29125 ( .A(n28424), .B(n28423), .Z(c[1706]) );
  NANDN U29126 ( .A(n28387), .B(n28386), .Z(n28391) );
  NAND U29127 ( .A(n28389), .B(n28388), .Z(n28390) );
  NAND U29128 ( .A(n28391), .B(n28390), .Z(n28430) );
  NAND U29129 ( .A(b[0]), .B(a[691]), .Z(n28392) );
  XNOR U29130 ( .A(b[1]), .B(n28392), .Z(n28394) );
  NAND U29131 ( .A(n113), .B(a[690]), .Z(n28393) );
  AND U29132 ( .A(n28394), .B(n28393), .Z(n28447) );
  XOR U29133 ( .A(a[687]), .B(n42197), .Z(n28436) );
  NANDN U29134 ( .A(n28436), .B(n42173), .Z(n28397) );
  NANDN U29135 ( .A(n28395), .B(n42172), .Z(n28396) );
  NAND U29136 ( .A(n28397), .B(n28396), .Z(n28445) );
  NAND U29137 ( .A(b[7]), .B(a[683]), .Z(n28446) );
  XNOR U29138 ( .A(n28445), .B(n28446), .Z(n28448) );
  XOR U29139 ( .A(n28447), .B(n28448), .Z(n28454) );
  NANDN U29140 ( .A(n28398), .B(n42093), .Z(n28400) );
  XOR U29141 ( .A(n42134), .B(a[689]), .Z(n28439) );
  NANDN U29142 ( .A(n28439), .B(n42095), .Z(n28399) );
  NAND U29143 ( .A(n28400), .B(n28399), .Z(n28452) );
  NANDN U29144 ( .A(n28401), .B(n42231), .Z(n28403) );
  XOR U29145 ( .A(n219), .B(a[685]), .Z(n28442) );
  NANDN U29146 ( .A(n28442), .B(n42234), .Z(n28402) );
  AND U29147 ( .A(n28403), .B(n28402), .Z(n28451) );
  XNOR U29148 ( .A(n28452), .B(n28451), .Z(n28453) );
  XNOR U29149 ( .A(n28454), .B(n28453), .Z(n28458) );
  NANDN U29150 ( .A(n28405), .B(n28404), .Z(n28409) );
  NAND U29151 ( .A(n28407), .B(n28406), .Z(n28408) );
  AND U29152 ( .A(n28409), .B(n28408), .Z(n28457) );
  XOR U29153 ( .A(n28458), .B(n28457), .Z(n28459) );
  NANDN U29154 ( .A(n28411), .B(n28410), .Z(n28415) );
  NANDN U29155 ( .A(n28413), .B(n28412), .Z(n28414) );
  NAND U29156 ( .A(n28415), .B(n28414), .Z(n28460) );
  XOR U29157 ( .A(n28459), .B(n28460), .Z(n28427) );
  OR U29158 ( .A(n28417), .B(n28416), .Z(n28421) );
  NANDN U29159 ( .A(n28419), .B(n28418), .Z(n28420) );
  NAND U29160 ( .A(n28421), .B(n28420), .Z(n28428) );
  XNOR U29161 ( .A(n28427), .B(n28428), .Z(n28429) );
  XNOR U29162 ( .A(n28430), .B(n28429), .Z(n28463) );
  XNOR U29163 ( .A(n28463), .B(sreg[1707]), .Z(n28465) );
  NAND U29164 ( .A(n28422), .B(sreg[1706]), .Z(n28426) );
  OR U29165 ( .A(n28424), .B(n28423), .Z(n28425) );
  AND U29166 ( .A(n28426), .B(n28425), .Z(n28464) );
  XOR U29167 ( .A(n28465), .B(n28464), .Z(c[1707]) );
  NANDN U29168 ( .A(n28428), .B(n28427), .Z(n28432) );
  NAND U29169 ( .A(n28430), .B(n28429), .Z(n28431) );
  NAND U29170 ( .A(n28432), .B(n28431), .Z(n28471) );
  NAND U29171 ( .A(b[0]), .B(a[692]), .Z(n28433) );
  XNOR U29172 ( .A(b[1]), .B(n28433), .Z(n28435) );
  NAND U29173 ( .A(n113), .B(a[691]), .Z(n28434) );
  AND U29174 ( .A(n28435), .B(n28434), .Z(n28488) );
  XOR U29175 ( .A(a[688]), .B(n42197), .Z(n28477) );
  NANDN U29176 ( .A(n28477), .B(n42173), .Z(n28438) );
  NANDN U29177 ( .A(n28436), .B(n42172), .Z(n28437) );
  NAND U29178 ( .A(n28438), .B(n28437), .Z(n28486) );
  NAND U29179 ( .A(b[7]), .B(a[684]), .Z(n28487) );
  XNOR U29180 ( .A(n28486), .B(n28487), .Z(n28489) );
  XOR U29181 ( .A(n28488), .B(n28489), .Z(n28495) );
  NANDN U29182 ( .A(n28439), .B(n42093), .Z(n28441) );
  XOR U29183 ( .A(n42134), .B(a[690]), .Z(n28480) );
  NANDN U29184 ( .A(n28480), .B(n42095), .Z(n28440) );
  NAND U29185 ( .A(n28441), .B(n28440), .Z(n28493) );
  NANDN U29186 ( .A(n28442), .B(n42231), .Z(n28444) );
  XOR U29187 ( .A(n219), .B(a[686]), .Z(n28483) );
  NANDN U29188 ( .A(n28483), .B(n42234), .Z(n28443) );
  AND U29189 ( .A(n28444), .B(n28443), .Z(n28492) );
  XNOR U29190 ( .A(n28493), .B(n28492), .Z(n28494) );
  XNOR U29191 ( .A(n28495), .B(n28494), .Z(n28499) );
  NANDN U29192 ( .A(n28446), .B(n28445), .Z(n28450) );
  NAND U29193 ( .A(n28448), .B(n28447), .Z(n28449) );
  AND U29194 ( .A(n28450), .B(n28449), .Z(n28498) );
  XOR U29195 ( .A(n28499), .B(n28498), .Z(n28500) );
  NANDN U29196 ( .A(n28452), .B(n28451), .Z(n28456) );
  NANDN U29197 ( .A(n28454), .B(n28453), .Z(n28455) );
  NAND U29198 ( .A(n28456), .B(n28455), .Z(n28501) );
  XOR U29199 ( .A(n28500), .B(n28501), .Z(n28468) );
  OR U29200 ( .A(n28458), .B(n28457), .Z(n28462) );
  NANDN U29201 ( .A(n28460), .B(n28459), .Z(n28461) );
  NAND U29202 ( .A(n28462), .B(n28461), .Z(n28469) );
  XNOR U29203 ( .A(n28468), .B(n28469), .Z(n28470) );
  XNOR U29204 ( .A(n28471), .B(n28470), .Z(n28504) );
  XNOR U29205 ( .A(n28504), .B(sreg[1708]), .Z(n28506) );
  NAND U29206 ( .A(n28463), .B(sreg[1707]), .Z(n28467) );
  OR U29207 ( .A(n28465), .B(n28464), .Z(n28466) );
  AND U29208 ( .A(n28467), .B(n28466), .Z(n28505) );
  XOR U29209 ( .A(n28506), .B(n28505), .Z(c[1708]) );
  NANDN U29210 ( .A(n28469), .B(n28468), .Z(n28473) );
  NAND U29211 ( .A(n28471), .B(n28470), .Z(n28472) );
  NAND U29212 ( .A(n28473), .B(n28472), .Z(n28512) );
  NAND U29213 ( .A(b[0]), .B(a[693]), .Z(n28474) );
  XNOR U29214 ( .A(b[1]), .B(n28474), .Z(n28476) );
  NAND U29215 ( .A(n114), .B(a[692]), .Z(n28475) );
  AND U29216 ( .A(n28476), .B(n28475), .Z(n28529) );
  XOR U29217 ( .A(a[689]), .B(n42197), .Z(n28518) );
  NANDN U29218 ( .A(n28518), .B(n42173), .Z(n28479) );
  NANDN U29219 ( .A(n28477), .B(n42172), .Z(n28478) );
  NAND U29220 ( .A(n28479), .B(n28478), .Z(n28527) );
  NAND U29221 ( .A(b[7]), .B(a[685]), .Z(n28528) );
  XNOR U29222 ( .A(n28527), .B(n28528), .Z(n28530) );
  XOR U29223 ( .A(n28529), .B(n28530), .Z(n28536) );
  NANDN U29224 ( .A(n28480), .B(n42093), .Z(n28482) );
  XOR U29225 ( .A(n42134), .B(a[691]), .Z(n28521) );
  NANDN U29226 ( .A(n28521), .B(n42095), .Z(n28481) );
  NAND U29227 ( .A(n28482), .B(n28481), .Z(n28534) );
  NANDN U29228 ( .A(n28483), .B(n42231), .Z(n28485) );
  XOR U29229 ( .A(n219), .B(a[687]), .Z(n28524) );
  NANDN U29230 ( .A(n28524), .B(n42234), .Z(n28484) );
  AND U29231 ( .A(n28485), .B(n28484), .Z(n28533) );
  XNOR U29232 ( .A(n28534), .B(n28533), .Z(n28535) );
  XNOR U29233 ( .A(n28536), .B(n28535), .Z(n28540) );
  NANDN U29234 ( .A(n28487), .B(n28486), .Z(n28491) );
  NAND U29235 ( .A(n28489), .B(n28488), .Z(n28490) );
  AND U29236 ( .A(n28491), .B(n28490), .Z(n28539) );
  XOR U29237 ( .A(n28540), .B(n28539), .Z(n28541) );
  NANDN U29238 ( .A(n28493), .B(n28492), .Z(n28497) );
  NANDN U29239 ( .A(n28495), .B(n28494), .Z(n28496) );
  NAND U29240 ( .A(n28497), .B(n28496), .Z(n28542) );
  XOR U29241 ( .A(n28541), .B(n28542), .Z(n28509) );
  OR U29242 ( .A(n28499), .B(n28498), .Z(n28503) );
  NANDN U29243 ( .A(n28501), .B(n28500), .Z(n28502) );
  NAND U29244 ( .A(n28503), .B(n28502), .Z(n28510) );
  XNOR U29245 ( .A(n28509), .B(n28510), .Z(n28511) );
  XNOR U29246 ( .A(n28512), .B(n28511), .Z(n28545) );
  XNOR U29247 ( .A(n28545), .B(sreg[1709]), .Z(n28547) );
  NAND U29248 ( .A(n28504), .B(sreg[1708]), .Z(n28508) );
  OR U29249 ( .A(n28506), .B(n28505), .Z(n28507) );
  AND U29250 ( .A(n28508), .B(n28507), .Z(n28546) );
  XOR U29251 ( .A(n28547), .B(n28546), .Z(c[1709]) );
  NANDN U29252 ( .A(n28510), .B(n28509), .Z(n28514) );
  NAND U29253 ( .A(n28512), .B(n28511), .Z(n28513) );
  NAND U29254 ( .A(n28514), .B(n28513), .Z(n28553) );
  NAND U29255 ( .A(b[0]), .B(a[694]), .Z(n28515) );
  XNOR U29256 ( .A(b[1]), .B(n28515), .Z(n28517) );
  NAND U29257 ( .A(n114), .B(a[693]), .Z(n28516) );
  AND U29258 ( .A(n28517), .B(n28516), .Z(n28570) );
  XOR U29259 ( .A(a[690]), .B(n42197), .Z(n28559) );
  NANDN U29260 ( .A(n28559), .B(n42173), .Z(n28520) );
  NANDN U29261 ( .A(n28518), .B(n42172), .Z(n28519) );
  NAND U29262 ( .A(n28520), .B(n28519), .Z(n28568) );
  NAND U29263 ( .A(b[7]), .B(a[686]), .Z(n28569) );
  XNOR U29264 ( .A(n28568), .B(n28569), .Z(n28571) );
  XOR U29265 ( .A(n28570), .B(n28571), .Z(n28577) );
  NANDN U29266 ( .A(n28521), .B(n42093), .Z(n28523) );
  XOR U29267 ( .A(n42134), .B(a[692]), .Z(n28562) );
  NANDN U29268 ( .A(n28562), .B(n42095), .Z(n28522) );
  NAND U29269 ( .A(n28523), .B(n28522), .Z(n28575) );
  NANDN U29270 ( .A(n28524), .B(n42231), .Z(n28526) );
  XOR U29271 ( .A(n219), .B(a[688]), .Z(n28565) );
  NANDN U29272 ( .A(n28565), .B(n42234), .Z(n28525) );
  AND U29273 ( .A(n28526), .B(n28525), .Z(n28574) );
  XNOR U29274 ( .A(n28575), .B(n28574), .Z(n28576) );
  XNOR U29275 ( .A(n28577), .B(n28576), .Z(n28581) );
  NANDN U29276 ( .A(n28528), .B(n28527), .Z(n28532) );
  NAND U29277 ( .A(n28530), .B(n28529), .Z(n28531) );
  AND U29278 ( .A(n28532), .B(n28531), .Z(n28580) );
  XOR U29279 ( .A(n28581), .B(n28580), .Z(n28582) );
  NANDN U29280 ( .A(n28534), .B(n28533), .Z(n28538) );
  NANDN U29281 ( .A(n28536), .B(n28535), .Z(n28537) );
  NAND U29282 ( .A(n28538), .B(n28537), .Z(n28583) );
  XOR U29283 ( .A(n28582), .B(n28583), .Z(n28550) );
  OR U29284 ( .A(n28540), .B(n28539), .Z(n28544) );
  NANDN U29285 ( .A(n28542), .B(n28541), .Z(n28543) );
  NAND U29286 ( .A(n28544), .B(n28543), .Z(n28551) );
  XNOR U29287 ( .A(n28550), .B(n28551), .Z(n28552) );
  XNOR U29288 ( .A(n28553), .B(n28552), .Z(n28586) );
  XNOR U29289 ( .A(n28586), .B(sreg[1710]), .Z(n28588) );
  NAND U29290 ( .A(n28545), .B(sreg[1709]), .Z(n28549) );
  OR U29291 ( .A(n28547), .B(n28546), .Z(n28548) );
  AND U29292 ( .A(n28549), .B(n28548), .Z(n28587) );
  XOR U29293 ( .A(n28588), .B(n28587), .Z(c[1710]) );
  NANDN U29294 ( .A(n28551), .B(n28550), .Z(n28555) );
  NAND U29295 ( .A(n28553), .B(n28552), .Z(n28554) );
  NAND U29296 ( .A(n28555), .B(n28554), .Z(n28594) );
  NAND U29297 ( .A(b[0]), .B(a[695]), .Z(n28556) );
  XNOR U29298 ( .A(b[1]), .B(n28556), .Z(n28558) );
  NAND U29299 ( .A(n114), .B(a[694]), .Z(n28557) );
  AND U29300 ( .A(n28558), .B(n28557), .Z(n28611) );
  XOR U29301 ( .A(a[691]), .B(n42197), .Z(n28600) );
  NANDN U29302 ( .A(n28600), .B(n42173), .Z(n28561) );
  NANDN U29303 ( .A(n28559), .B(n42172), .Z(n28560) );
  NAND U29304 ( .A(n28561), .B(n28560), .Z(n28609) );
  NAND U29305 ( .A(b[7]), .B(a[687]), .Z(n28610) );
  XNOR U29306 ( .A(n28609), .B(n28610), .Z(n28612) );
  XOR U29307 ( .A(n28611), .B(n28612), .Z(n28618) );
  NANDN U29308 ( .A(n28562), .B(n42093), .Z(n28564) );
  XOR U29309 ( .A(n42134), .B(a[693]), .Z(n28603) );
  NANDN U29310 ( .A(n28603), .B(n42095), .Z(n28563) );
  NAND U29311 ( .A(n28564), .B(n28563), .Z(n28616) );
  NANDN U29312 ( .A(n28565), .B(n42231), .Z(n28567) );
  XOR U29313 ( .A(n219), .B(a[689]), .Z(n28606) );
  NANDN U29314 ( .A(n28606), .B(n42234), .Z(n28566) );
  AND U29315 ( .A(n28567), .B(n28566), .Z(n28615) );
  XNOR U29316 ( .A(n28616), .B(n28615), .Z(n28617) );
  XNOR U29317 ( .A(n28618), .B(n28617), .Z(n28622) );
  NANDN U29318 ( .A(n28569), .B(n28568), .Z(n28573) );
  NAND U29319 ( .A(n28571), .B(n28570), .Z(n28572) );
  AND U29320 ( .A(n28573), .B(n28572), .Z(n28621) );
  XOR U29321 ( .A(n28622), .B(n28621), .Z(n28623) );
  NANDN U29322 ( .A(n28575), .B(n28574), .Z(n28579) );
  NANDN U29323 ( .A(n28577), .B(n28576), .Z(n28578) );
  NAND U29324 ( .A(n28579), .B(n28578), .Z(n28624) );
  XOR U29325 ( .A(n28623), .B(n28624), .Z(n28591) );
  OR U29326 ( .A(n28581), .B(n28580), .Z(n28585) );
  NANDN U29327 ( .A(n28583), .B(n28582), .Z(n28584) );
  NAND U29328 ( .A(n28585), .B(n28584), .Z(n28592) );
  XNOR U29329 ( .A(n28591), .B(n28592), .Z(n28593) );
  XNOR U29330 ( .A(n28594), .B(n28593), .Z(n28627) );
  XNOR U29331 ( .A(n28627), .B(sreg[1711]), .Z(n28629) );
  NAND U29332 ( .A(n28586), .B(sreg[1710]), .Z(n28590) );
  OR U29333 ( .A(n28588), .B(n28587), .Z(n28589) );
  AND U29334 ( .A(n28590), .B(n28589), .Z(n28628) );
  XOR U29335 ( .A(n28629), .B(n28628), .Z(c[1711]) );
  NANDN U29336 ( .A(n28592), .B(n28591), .Z(n28596) );
  NAND U29337 ( .A(n28594), .B(n28593), .Z(n28595) );
  NAND U29338 ( .A(n28596), .B(n28595), .Z(n28635) );
  NAND U29339 ( .A(b[0]), .B(a[696]), .Z(n28597) );
  XNOR U29340 ( .A(b[1]), .B(n28597), .Z(n28599) );
  NAND U29341 ( .A(n114), .B(a[695]), .Z(n28598) );
  AND U29342 ( .A(n28599), .B(n28598), .Z(n28652) );
  XOR U29343 ( .A(a[692]), .B(n42197), .Z(n28641) );
  NANDN U29344 ( .A(n28641), .B(n42173), .Z(n28602) );
  NANDN U29345 ( .A(n28600), .B(n42172), .Z(n28601) );
  NAND U29346 ( .A(n28602), .B(n28601), .Z(n28650) );
  NAND U29347 ( .A(b[7]), .B(a[688]), .Z(n28651) );
  XNOR U29348 ( .A(n28650), .B(n28651), .Z(n28653) );
  XOR U29349 ( .A(n28652), .B(n28653), .Z(n28659) );
  NANDN U29350 ( .A(n28603), .B(n42093), .Z(n28605) );
  XOR U29351 ( .A(n42134), .B(a[694]), .Z(n28644) );
  NANDN U29352 ( .A(n28644), .B(n42095), .Z(n28604) );
  NAND U29353 ( .A(n28605), .B(n28604), .Z(n28657) );
  NANDN U29354 ( .A(n28606), .B(n42231), .Z(n28608) );
  XOR U29355 ( .A(n219), .B(a[690]), .Z(n28647) );
  NANDN U29356 ( .A(n28647), .B(n42234), .Z(n28607) );
  AND U29357 ( .A(n28608), .B(n28607), .Z(n28656) );
  XNOR U29358 ( .A(n28657), .B(n28656), .Z(n28658) );
  XNOR U29359 ( .A(n28659), .B(n28658), .Z(n28663) );
  NANDN U29360 ( .A(n28610), .B(n28609), .Z(n28614) );
  NAND U29361 ( .A(n28612), .B(n28611), .Z(n28613) );
  AND U29362 ( .A(n28614), .B(n28613), .Z(n28662) );
  XOR U29363 ( .A(n28663), .B(n28662), .Z(n28664) );
  NANDN U29364 ( .A(n28616), .B(n28615), .Z(n28620) );
  NANDN U29365 ( .A(n28618), .B(n28617), .Z(n28619) );
  NAND U29366 ( .A(n28620), .B(n28619), .Z(n28665) );
  XOR U29367 ( .A(n28664), .B(n28665), .Z(n28632) );
  OR U29368 ( .A(n28622), .B(n28621), .Z(n28626) );
  NANDN U29369 ( .A(n28624), .B(n28623), .Z(n28625) );
  NAND U29370 ( .A(n28626), .B(n28625), .Z(n28633) );
  XNOR U29371 ( .A(n28632), .B(n28633), .Z(n28634) );
  XNOR U29372 ( .A(n28635), .B(n28634), .Z(n28668) );
  XNOR U29373 ( .A(n28668), .B(sreg[1712]), .Z(n28670) );
  NAND U29374 ( .A(n28627), .B(sreg[1711]), .Z(n28631) );
  OR U29375 ( .A(n28629), .B(n28628), .Z(n28630) );
  AND U29376 ( .A(n28631), .B(n28630), .Z(n28669) );
  XOR U29377 ( .A(n28670), .B(n28669), .Z(c[1712]) );
  NANDN U29378 ( .A(n28633), .B(n28632), .Z(n28637) );
  NAND U29379 ( .A(n28635), .B(n28634), .Z(n28636) );
  NAND U29380 ( .A(n28637), .B(n28636), .Z(n28676) );
  NAND U29381 ( .A(b[0]), .B(a[697]), .Z(n28638) );
  XNOR U29382 ( .A(b[1]), .B(n28638), .Z(n28640) );
  NAND U29383 ( .A(n114), .B(a[696]), .Z(n28639) );
  AND U29384 ( .A(n28640), .B(n28639), .Z(n28693) );
  XOR U29385 ( .A(a[693]), .B(n42197), .Z(n28682) );
  NANDN U29386 ( .A(n28682), .B(n42173), .Z(n28643) );
  NANDN U29387 ( .A(n28641), .B(n42172), .Z(n28642) );
  NAND U29388 ( .A(n28643), .B(n28642), .Z(n28691) );
  NAND U29389 ( .A(b[7]), .B(a[689]), .Z(n28692) );
  XNOR U29390 ( .A(n28691), .B(n28692), .Z(n28694) );
  XOR U29391 ( .A(n28693), .B(n28694), .Z(n28700) );
  NANDN U29392 ( .A(n28644), .B(n42093), .Z(n28646) );
  XOR U29393 ( .A(n42134), .B(a[695]), .Z(n28685) );
  NANDN U29394 ( .A(n28685), .B(n42095), .Z(n28645) );
  NAND U29395 ( .A(n28646), .B(n28645), .Z(n28698) );
  NANDN U29396 ( .A(n28647), .B(n42231), .Z(n28649) );
  XOR U29397 ( .A(n219), .B(a[691]), .Z(n28688) );
  NANDN U29398 ( .A(n28688), .B(n42234), .Z(n28648) );
  AND U29399 ( .A(n28649), .B(n28648), .Z(n28697) );
  XNOR U29400 ( .A(n28698), .B(n28697), .Z(n28699) );
  XNOR U29401 ( .A(n28700), .B(n28699), .Z(n28704) );
  NANDN U29402 ( .A(n28651), .B(n28650), .Z(n28655) );
  NAND U29403 ( .A(n28653), .B(n28652), .Z(n28654) );
  AND U29404 ( .A(n28655), .B(n28654), .Z(n28703) );
  XOR U29405 ( .A(n28704), .B(n28703), .Z(n28705) );
  NANDN U29406 ( .A(n28657), .B(n28656), .Z(n28661) );
  NANDN U29407 ( .A(n28659), .B(n28658), .Z(n28660) );
  NAND U29408 ( .A(n28661), .B(n28660), .Z(n28706) );
  XOR U29409 ( .A(n28705), .B(n28706), .Z(n28673) );
  OR U29410 ( .A(n28663), .B(n28662), .Z(n28667) );
  NANDN U29411 ( .A(n28665), .B(n28664), .Z(n28666) );
  NAND U29412 ( .A(n28667), .B(n28666), .Z(n28674) );
  XNOR U29413 ( .A(n28673), .B(n28674), .Z(n28675) );
  XNOR U29414 ( .A(n28676), .B(n28675), .Z(n28709) );
  XNOR U29415 ( .A(n28709), .B(sreg[1713]), .Z(n28711) );
  NAND U29416 ( .A(n28668), .B(sreg[1712]), .Z(n28672) );
  OR U29417 ( .A(n28670), .B(n28669), .Z(n28671) );
  AND U29418 ( .A(n28672), .B(n28671), .Z(n28710) );
  XOR U29419 ( .A(n28711), .B(n28710), .Z(c[1713]) );
  NANDN U29420 ( .A(n28674), .B(n28673), .Z(n28678) );
  NAND U29421 ( .A(n28676), .B(n28675), .Z(n28677) );
  NAND U29422 ( .A(n28678), .B(n28677), .Z(n28717) );
  NAND U29423 ( .A(b[0]), .B(a[698]), .Z(n28679) );
  XNOR U29424 ( .A(b[1]), .B(n28679), .Z(n28681) );
  NAND U29425 ( .A(n114), .B(a[697]), .Z(n28680) );
  AND U29426 ( .A(n28681), .B(n28680), .Z(n28734) );
  XOR U29427 ( .A(a[694]), .B(n42197), .Z(n28723) );
  NANDN U29428 ( .A(n28723), .B(n42173), .Z(n28684) );
  NANDN U29429 ( .A(n28682), .B(n42172), .Z(n28683) );
  NAND U29430 ( .A(n28684), .B(n28683), .Z(n28732) );
  NAND U29431 ( .A(b[7]), .B(a[690]), .Z(n28733) );
  XNOR U29432 ( .A(n28732), .B(n28733), .Z(n28735) );
  XOR U29433 ( .A(n28734), .B(n28735), .Z(n28741) );
  NANDN U29434 ( .A(n28685), .B(n42093), .Z(n28687) );
  XOR U29435 ( .A(n42134), .B(a[696]), .Z(n28726) );
  NANDN U29436 ( .A(n28726), .B(n42095), .Z(n28686) );
  NAND U29437 ( .A(n28687), .B(n28686), .Z(n28739) );
  NANDN U29438 ( .A(n28688), .B(n42231), .Z(n28690) );
  XOR U29439 ( .A(n219), .B(a[692]), .Z(n28729) );
  NANDN U29440 ( .A(n28729), .B(n42234), .Z(n28689) );
  AND U29441 ( .A(n28690), .B(n28689), .Z(n28738) );
  XNOR U29442 ( .A(n28739), .B(n28738), .Z(n28740) );
  XNOR U29443 ( .A(n28741), .B(n28740), .Z(n28745) );
  NANDN U29444 ( .A(n28692), .B(n28691), .Z(n28696) );
  NAND U29445 ( .A(n28694), .B(n28693), .Z(n28695) );
  AND U29446 ( .A(n28696), .B(n28695), .Z(n28744) );
  XOR U29447 ( .A(n28745), .B(n28744), .Z(n28746) );
  NANDN U29448 ( .A(n28698), .B(n28697), .Z(n28702) );
  NANDN U29449 ( .A(n28700), .B(n28699), .Z(n28701) );
  NAND U29450 ( .A(n28702), .B(n28701), .Z(n28747) );
  XOR U29451 ( .A(n28746), .B(n28747), .Z(n28714) );
  OR U29452 ( .A(n28704), .B(n28703), .Z(n28708) );
  NANDN U29453 ( .A(n28706), .B(n28705), .Z(n28707) );
  NAND U29454 ( .A(n28708), .B(n28707), .Z(n28715) );
  XNOR U29455 ( .A(n28714), .B(n28715), .Z(n28716) );
  XNOR U29456 ( .A(n28717), .B(n28716), .Z(n28750) );
  XNOR U29457 ( .A(n28750), .B(sreg[1714]), .Z(n28752) );
  NAND U29458 ( .A(n28709), .B(sreg[1713]), .Z(n28713) );
  OR U29459 ( .A(n28711), .B(n28710), .Z(n28712) );
  AND U29460 ( .A(n28713), .B(n28712), .Z(n28751) );
  XOR U29461 ( .A(n28752), .B(n28751), .Z(c[1714]) );
  NANDN U29462 ( .A(n28715), .B(n28714), .Z(n28719) );
  NAND U29463 ( .A(n28717), .B(n28716), .Z(n28718) );
  NAND U29464 ( .A(n28719), .B(n28718), .Z(n28758) );
  NAND U29465 ( .A(b[0]), .B(a[699]), .Z(n28720) );
  XNOR U29466 ( .A(b[1]), .B(n28720), .Z(n28722) );
  NAND U29467 ( .A(n114), .B(a[698]), .Z(n28721) );
  AND U29468 ( .A(n28722), .B(n28721), .Z(n28775) );
  XOR U29469 ( .A(a[695]), .B(n42197), .Z(n28764) );
  NANDN U29470 ( .A(n28764), .B(n42173), .Z(n28725) );
  NANDN U29471 ( .A(n28723), .B(n42172), .Z(n28724) );
  NAND U29472 ( .A(n28725), .B(n28724), .Z(n28773) );
  NAND U29473 ( .A(b[7]), .B(a[691]), .Z(n28774) );
  XNOR U29474 ( .A(n28773), .B(n28774), .Z(n28776) );
  XOR U29475 ( .A(n28775), .B(n28776), .Z(n28782) );
  NANDN U29476 ( .A(n28726), .B(n42093), .Z(n28728) );
  XOR U29477 ( .A(n42134), .B(a[697]), .Z(n28767) );
  NANDN U29478 ( .A(n28767), .B(n42095), .Z(n28727) );
  NAND U29479 ( .A(n28728), .B(n28727), .Z(n28780) );
  NANDN U29480 ( .A(n28729), .B(n42231), .Z(n28731) );
  XOR U29481 ( .A(n219), .B(a[693]), .Z(n28770) );
  NANDN U29482 ( .A(n28770), .B(n42234), .Z(n28730) );
  AND U29483 ( .A(n28731), .B(n28730), .Z(n28779) );
  XNOR U29484 ( .A(n28780), .B(n28779), .Z(n28781) );
  XNOR U29485 ( .A(n28782), .B(n28781), .Z(n28786) );
  NANDN U29486 ( .A(n28733), .B(n28732), .Z(n28737) );
  NAND U29487 ( .A(n28735), .B(n28734), .Z(n28736) );
  AND U29488 ( .A(n28737), .B(n28736), .Z(n28785) );
  XOR U29489 ( .A(n28786), .B(n28785), .Z(n28787) );
  NANDN U29490 ( .A(n28739), .B(n28738), .Z(n28743) );
  NANDN U29491 ( .A(n28741), .B(n28740), .Z(n28742) );
  NAND U29492 ( .A(n28743), .B(n28742), .Z(n28788) );
  XOR U29493 ( .A(n28787), .B(n28788), .Z(n28755) );
  OR U29494 ( .A(n28745), .B(n28744), .Z(n28749) );
  NANDN U29495 ( .A(n28747), .B(n28746), .Z(n28748) );
  NAND U29496 ( .A(n28749), .B(n28748), .Z(n28756) );
  XNOR U29497 ( .A(n28755), .B(n28756), .Z(n28757) );
  XNOR U29498 ( .A(n28758), .B(n28757), .Z(n28791) );
  XNOR U29499 ( .A(n28791), .B(sreg[1715]), .Z(n28793) );
  NAND U29500 ( .A(n28750), .B(sreg[1714]), .Z(n28754) );
  OR U29501 ( .A(n28752), .B(n28751), .Z(n28753) );
  AND U29502 ( .A(n28754), .B(n28753), .Z(n28792) );
  XOR U29503 ( .A(n28793), .B(n28792), .Z(c[1715]) );
  NANDN U29504 ( .A(n28756), .B(n28755), .Z(n28760) );
  NAND U29505 ( .A(n28758), .B(n28757), .Z(n28759) );
  NAND U29506 ( .A(n28760), .B(n28759), .Z(n28799) );
  NAND U29507 ( .A(b[0]), .B(a[700]), .Z(n28761) );
  XNOR U29508 ( .A(b[1]), .B(n28761), .Z(n28763) );
  NAND U29509 ( .A(n115), .B(a[699]), .Z(n28762) );
  AND U29510 ( .A(n28763), .B(n28762), .Z(n28816) );
  XOR U29511 ( .A(a[696]), .B(n42197), .Z(n28805) );
  NANDN U29512 ( .A(n28805), .B(n42173), .Z(n28766) );
  NANDN U29513 ( .A(n28764), .B(n42172), .Z(n28765) );
  NAND U29514 ( .A(n28766), .B(n28765), .Z(n28814) );
  NAND U29515 ( .A(b[7]), .B(a[692]), .Z(n28815) );
  XNOR U29516 ( .A(n28814), .B(n28815), .Z(n28817) );
  XOR U29517 ( .A(n28816), .B(n28817), .Z(n28823) );
  NANDN U29518 ( .A(n28767), .B(n42093), .Z(n28769) );
  XOR U29519 ( .A(n42134), .B(a[698]), .Z(n28808) );
  NANDN U29520 ( .A(n28808), .B(n42095), .Z(n28768) );
  NAND U29521 ( .A(n28769), .B(n28768), .Z(n28821) );
  NANDN U29522 ( .A(n28770), .B(n42231), .Z(n28772) );
  XOR U29523 ( .A(n219), .B(a[694]), .Z(n28811) );
  NANDN U29524 ( .A(n28811), .B(n42234), .Z(n28771) );
  AND U29525 ( .A(n28772), .B(n28771), .Z(n28820) );
  XNOR U29526 ( .A(n28821), .B(n28820), .Z(n28822) );
  XNOR U29527 ( .A(n28823), .B(n28822), .Z(n28827) );
  NANDN U29528 ( .A(n28774), .B(n28773), .Z(n28778) );
  NAND U29529 ( .A(n28776), .B(n28775), .Z(n28777) );
  AND U29530 ( .A(n28778), .B(n28777), .Z(n28826) );
  XOR U29531 ( .A(n28827), .B(n28826), .Z(n28828) );
  NANDN U29532 ( .A(n28780), .B(n28779), .Z(n28784) );
  NANDN U29533 ( .A(n28782), .B(n28781), .Z(n28783) );
  NAND U29534 ( .A(n28784), .B(n28783), .Z(n28829) );
  XOR U29535 ( .A(n28828), .B(n28829), .Z(n28796) );
  OR U29536 ( .A(n28786), .B(n28785), .Z(n28790) );
  NANDN U29537 ( .A(n28788), .B(n28787), .Z(n28789) );
  NAND U29538 ( .A(n28790), .B(n28789), .Z(n28797) );
  XNOR U29539 ( .A(n28796), .B(n28797), .Z(n28798) );
  XNOR U29540 ( .A(n28799), .B(n28798), .Z(n28832) );
  XNOR U29541 ( .A(n28832), .B(sreg[1716]), .Z(n28834) );
  NAND U29542 ( .A(n28791), .B(sreg[1715]), .Z(n28795) );
  OR U29543 ( .A(n28793), .B(n28792), .Z(n28794) );
  AND U29544 ( .A(n28795), .B(n28794), .Z(n28833) );
  XOR U29545 ( .A(n28834), .B(n28833), .Z(c[1716]) );
  NANDN U29546 ( .A(n28797), .B(n28796), .Z(n28801) );
  NAND U29547 ( .A(n28799), .B(n28798), .Z(n28800) );
  NAND U29548 ( .A(n28801), .B(n28800), .Z(n28840) );
  NAND U29549 ( .A(b[0]), .B(a[701]), .Z(n28802) );
  XNOR U29550 ( .A(b[1]), .B(n28802), .Z(n28804) );
  NAND U29551 ( .A(n115), .B(a[700]), .Z(n28803) );
  AND U29552 ( .A(n28804), .B(n28803), .Z(n28857) );
  XOR U29553 ( .A(a[697]), .B(n42197), .Z(n28846) );
  NANDN U29554 ( .A(n28846), .B(n42173), .Z(n28807) );
  NANDN U29555 ( .A(n28805), .B(n42172), .Z(n28806) );
  NAND U29556 ( .A(n28807), .B(n28806), .Z(n28855) );
  NAND U29557 ( .A(b[7]), .B(a[693]), .Z(n28856) );
  XNOR U29558 ( .A(n28855), .B(n28856), .Z(n28858) );
  XOR U29559 ( .A(n28857), .B(n28858), .Z(n28864) );
  NANDN U29560 ( .A(n28808), .B(n42093), .Z(n28810) );
  XOR U29561 ( .A(n42134), .B(a[699]), .Z(n28849) );
  NANDN U29562 ( .A(n28849), .B(n42095), .Z(n28809) );
  NAND U29563 ( .A(n28810), .B(n28809), .Z(n28862) );
  NANDN U29564 ( .A(n28811), .B(n42231), .Z(n28813) );
  XOR U29565 ( .A(n220), .B(a[695]), .Z(n28852) );
  NANDN U29566 ( .A(n28852), .B(n42234), .Z(n28812) );
  AND U29567 ( .A(n28813), .B(n28812), .Z(n28861) );
  XNOR U29568 ( .A(n28862), .B(n28861), .Z(n28863) );
  XNOR U29569 ( .A(n28864), .B(n28863), .Z(n28868) );
  NANDN U29570 ( .A(n28815), .B(n28814), .Z(n28819) );
  NAND U29571 ( .A(n28817), .B(n28816), .Z(n28818) );
  AND U29572 ( .A(n28819), .B(n28818), .Z(n28867) );
  XOR U29573 ( .A(n28868), .B(n28867), .Z(n28869) );
  NANDN U29574 ( .A(n28821), .B(n28820), .Z(n28825) );
  NANDN U29575 ( .A(n28823), .B(n28822), .Z(n28824) );
  NAND U29576 ( .A(n28825), .B(n28824), .Z(n28870) );
  XOR U29577 ( .A(n28869), .B(n28870), .Z(n28837) );
  OR U29578 ( .A(n28827), .B(n28826), .Z(n28831) );
  NANDN U29579 ( .A(n28829), .B(n28828), .Z(n28830) );
  NAND U29580 ( .A(n28831), .B(n28830), .Z(n28838) );
  XNOR U29581 ( .A(n28837), .B(n28838), .Z(n28839) );
  XNOR U29582 ( .A(n28840), .B(n28839), .Z(n28873) );
  XNOR U29583 ( .A(n28873), .B(sreg[1717]), .Z(n28875) );
  NAND U29584 ( .A(n28832), .B(sreg[1716]), .Z(n28836) );
  OR U29585 ( .A(n28834), .B(n28833), .Z(n28835) );
  AND U29586 ( .A(n28836), .B(n28835), .Z(n28874) );
  XOR U29587 ( .A(n28875), .B(n28874), .Z(c[1717]) );
  NANDN U29588 ( .A(n28838), .B(n28837), .Z(n28842) );
  NAND U29589 ( .A(n28840), .B(n28839), .Z(n28841) );
  NAND U29590 ( .A(n28842), .B(n28841), .Z(n28881) );
  NAND U29591 ( .A(b[0]), .B(a[702]), .Z(n28843) );
  XNOR U29592 ( .A(b[1]), .B(n28843), .Z(n28845) );
  NAND U29593 ( .A(n115), .B(a[701]), .Z(n28844) );
  AND U29594 ( .A(n28845), .B(n28844), .Z(n28898) );
  XOR U29595 ( .A(a[698]), .B(n42197), .Z(n28887) );
  NANDN U29596 ( .A(n28887), .B(n42173), .Z(n28848) );
  NANDN U29597 ( .A(n28846), .B(n42172), .Z(n28847) );
  NAND U29598 ( .A(n28848), .B(n28847), .Z(n28896) );
  NAND U29599 ( .A(b[7]), .B(a[694]), .Z(n28897) );
  XNOR U29600 ( .A(n28896), .B(n28897), .Z(n28899) );
  XOR U29601 ( .A(n28898), .B(n28899), .Z(n28905) );
  NANDN U29602 ( .A(n28849), .B(n42093), .Z(n28851) );
  XOR U29603 ( .A(n42134), .B(a[700]), .Z(n28890) );
  NANDN U29604 ( .A(n28890), .B(n42095), .Z(n28850) );
  NAND U29605 ( .A(n28851), .B(n28850), .Z(n28903) );
  NANDN U29606 ( .A(n28852), .B(n42231), .Z(n28854) );
  XOR U29607 ( .A(n220), .B(a[696]), .Z(n28893) );
  NANDN U29608 ( .A(n28893), .B(n42234), .Z(n28853) );
  AND U29609 ( .A(n28854), .B(n28853), .Z(n28902) );
  XNOR U29610 ( .A(n28903), .B(n28902), .Z(n28904) );
  XNOR U29611 ( .A(n28905), .B(n28904), .Z(n28909) );
  NANDN U29612 ( .A(n28856), .B(n28855), .Z(n28860) );
  NAND U29613 ( .A(n28858), .B(n28857), .Z(n28859) );
  AND U29614 ( .A(n28860), .B(n28859), .Z(n28908) );
  XOR U29615 ( .A(n28909), .B(n28908), .Z(n28910) );
  NANDN U29616 ( .A(n28862), .B(n28861), .Z(n28866) );
  NANDN U29617 ( .A(n28864), .B(n28863), .Z(n28865) );
  NAND U29618 ( .A(n28866), .B(n28865), .Z(n28911) );
  XOR U29619 ( .A(n28910), .B(n28911), .Z(n28878) );
  OR U29620 ( .A(n28868), .B(n28867), .Z(n28872) );
  NANDN U29621 ( .A(n28870), .B(n28869), .Z(n28871) );
  NAND U29622 ( .A(n28872), .B(n28871), .Z(n28879) );
  XNOR U29623 ( .A(n28878), .B(n28879), .Z(n28880) );
  XNOR U29624 ( .A(n28881), .B(n28880), .Z(n28914) );
  XNOR U29625 ( .A(n28914), .B(sreg[1718]), .Z(n28916) );
  NAND U29626 ( .A(n28873), .B(sreg[1717]), .Z(n28877) );
  OR U29627 ( .A(n28875), .B(n28874), .Z(n28876) );
  AND U29628 ( .A(n28877), .B(n28876), .Z(n28915) );
  XOR U29629 ( .A(n28916), .B(n28915), .Z(c[1718]) );
  NANDN U29630 ( .A(n28879), .B(n28878), .Z(n28883) );
  NAND U29631 ( .A(n28881), .B(n28880), .Z(n28882) );
  NAND U29632 ( .A(n28883), .B(n28882), .Z(n28922) );
  NAND U29633 ( .A(b[0]), .B(a[703]), .Z(n28884) );
  XNOR U29634 ( .A(b[1]), .B(n28884), .Z(n28886) );
  NAND U29635 ( .A(n115), .B(a[702]), .Z(n28885) );
  AND U29636 ( .A(n28886), .B(n28885), .Z(n28939) );
  XOR U29637 ( .A(a[699]), .B(n42197), .Z(n28928) );
  NANDN U29638 ( .A(n28928), .B(n42173), .Z(n28889) );
  NANDN U29639 ( .A(n28887), .B(n42172), .Z(n28888) );
  NAND U29640 ( .A(n28889), .B(n28888), .Z(n28937) );
  NAND U29641 ( .A(b[7]), .B(a[695]), .Z(n28938) );
  XNOR U29642 ( .A(n28937), .B(n28938), .Z(n28940) );
  XOR U29643 ( .A(n28939), .B(n28940), .Z(n28946) );
  NANDN U29644 ( .A(n28890), .B(n42093), .Z(n28892) );
  XOR U29645 ( .A(n42134), .B(a[701]), .Z(n28931) );
  NANDN U29646 ( .A(n28931), .B(n42095), .Z(n28891) );
  NAND U29647 ( .A(n28892), .B(n28891), .Z(n28944) );
  NANDN U29648 ( .A(n28893), .B(n42231), .Z(n28895) );
  XOR U29649 ( .A(n220), .B(a[697]), .Z(n28934) );
  NANDN U29650 ( .A(n28934), .B(n42234), .Z(n28894) );
  AND U29651 ( .A(n28895), .B(n28894), .Z(n28943) );
  XNOR U29652 ( .A(n28944), .B(n28943), .Z(n28945) );
  XNOR U29653 ( .A(n28946), .B(n28945), .Z(n28950) );
  NANDN U29654 ( .A(n28897), .B(n28896), .Z(n28901) );
  NAND U29655 ( .A(n28899), .B(n28898), .Z(n28900) );
  AND U29656 ( .A(n28901), .B(n28900), .Z(n28949) );
  XOR U29657 ( .A(n28950), .B(n28949), .Z(n28951) );
  NANDN U29658 ( .A(n28903), .B(n28902), .Z(n28907) );
  NANDN U29659 ( .A(n28905), .B(n28904), .Z(n28906) );
  NAND U29660 ( .A(n28907), .B(n28906), .Z(n28952) );
  XOR U29661 ( .A(n28951), .B(n28952), .Z(n28919) );
  OR U29662 ( .A(n28909), .B(n28908), .Z(n28913) );
  NANDN U29663 ( .A(n28911), .B(n28910), .Z(n28912) );
  NAND U29664 ( .A(n28913), .B(n28912), .Z(n28920) );
  XNOR U29665 ( .A(n28919), .B(n28920), .Z(n28921) );
  XNOR U29666 ( .A(n28922), .B(n28921), .Z(n28955) );
  XNOR U29667 ( .A(n28955), .B(sreg[1719]), .Z(n28957) );
  NAND U29668 ( .A(n28914), .B(sreg[1718]), .Z(n28918) );
  OR U29669 ( .A(n28916), .B(n28915), .Z(n28917) );
  AND U29670 ( .A(n28918), .B(n28917), .Z(n28956) );
  XOR U29671 ( .A(n28957), .B(n28956), .Z(c[1719]) );
  NANDN U29672 ( .A(n28920), .B(n28919), .Z(n28924) );
  NAND U29673 ( .A(n28922), .B(n28921), .Z(n28923) );
  NAND U29674 ( .A(n28924), .B(n28923), .Z(n28963) );
  NAND U29675 ( .A(b[0]), .B(a[704]), .Z(n28925) );
  XNOR U29676 ( .A(b[1]), .B(n28925), .Z(n28927) );
  NAND U29677 ( .A(n115), .B(a[703]), .Z(n28926) );
  AND U29678 ( .A(n28927), .B(n28926), .Z(n28980) );
  XOR U29679 ( .A(a[700]), .B(n42197), .Z(n28969) );
  NANDN U29680 ( .A(n28969), .B(n42173), .Z(n28930) );
  NANDN U29681 ( .A(n28928), .B(n42172), .Z(n28929) );
  NAND U29682 ( .A(n28930), .B(n28929), .Z(n28978) );
  NAND U29683 ( .A(b[7]), .B(a[696]), .Z(n28979) );
  XNOR U29684 ( .A(n28978), .B(n28979), .Z(n28981) );
  XOR U29685 ( .A(n28980), .B(n28981), .Z(n28987) );
  NANDN U29686 ( .A(n28931), .B(n42093), .Z(n28933) );
  XOR U29687 ( .A(n42134), .B(a[702]), .Z(n28972) );
  NANDN U29688 ( .A(n28972), .B(n42095), .Z(n28932) );
  NAND U29689 ( .A(n28933), .B(n28932), .Z(n28985) );
  NANDN U29690 ( .A(n28934), .B(n42231), .Z(n28936) );
  XOR U29691 ( .A(n220), .B(a[698]), .Z(n28975) );
  NANDN U29692 ( .A(n28975), .B(n42234), .Z(n28935) );
  AND U29693 ( .A(n28936), .B(n28935), .Z(n28984) );
  XNOR U29694 ( .A(n28985), .B(n28984), .Z(n28986) );
  XNOR U29695 ( .A(n28987), .B(n28986), .Z(n28991) );
  NANDN U29696 ( .A(n28938), .B(n28937), .Z(n28942) );
  NAND U29697 ( .A(n28940), .B(n28939), .Z(n28941) );
  AND U29698 ( .A(n28942), .B(n28941), .Z(n28990) );
  XOR U29699 ( .A(n28991), .B(n28990), .Z(n28992) );
  NANDN U29700 ( .A(n28944), .B(n28943), .Z(n28948) );
  NANDN U29701 ( .A(n28946), .B(n28945), .Z(n28947) );
  NAND U29702 ( .A(n28948), .B(n28947), .Z(n28993) );
  XOR U29703 ( .A(n28992), .B(n28993), .Z(n28960) );
  OR U29704 ( .A(n28950), .B(n28949), .Z(n28954) );
  NANDN U29705 ( .A(n28952), .B(n28951), .Z(n28953) );
  NAND U29706 ( .A(n28954), .B(n28953), .Z(n28961) );
  XNOR U29707 ( .A(n28960), .B(n28961), .Z(n28962) );
  XNOR U29708 ( .A(n28963), .B(n28962), .Z(n28996) );
  XNOR U29709 ( .A(n28996), .B(sreg[1720]), .Z(n28998) );
  NAND U29710 ( .A(n28955), .B(sreg[1719]), .Z(n28959) );
  OR U29711 ( .A(n28957), .B(n28956), .Z(n28958) );
  AND U29712 ( .A(n28959), .B(n28958), .Z(n28997) );
  XOR U29713 ( .A(n28998), .B(n28997), .Z(c[1720]) );
  NANDN U29714 ( .A(n28961), .B(n28960), .Z(n28965) );
  NAND U29715 ( .A(n28963), .B(n28962), .Z(n28964) );
  NAND U29716 ( .A(n28965), .B(n28964), .Z(n29004) );
  NAND U29717 ( .A(b[0]), .B(a[705]), .Z(n28966) );
  XNOR U29718 ( .A(b[1]), .B(n28966), .Z(n28968) );
  NAND U29719 ( .A(n115), .B(a[704]), .Z(n28967) );
  AND U29720 ( .A(n28968), .B(n28967), .Z(n29021) );
  XOR U29721 ( .A(a[701]), .B(n42197), .Z(n29010) );
  NANDN U29722 ( .A(n29010), .B(n42173), .Z(n28971) );
  NANDN U29723 ( .A(n28969), .B(n42172), .Z(n28970) );
  NAND U29724 ( .A(n28971), .B(n28970), .Z(n29019) );
  NAND U29725 ( .A(b[7]), .B(a[697]), .Z(n29020) );
  XNOR U29726 ( .A(n29019), .B(n29020), .Z(n29022) );
  XOR U29727 ( .A(n29021), .B(n29022), .Z(n29028) );
  NANDN U29728 ( .A(n28972), .B(n42093), .Z(n28974) );
  XOR U29729 ( .A(n42134), .B(a[703]), .Z(n29013) );
  NANDN U29730 ( .A(n29013), .B(n42095), .Z(n28973) );
  NAND U29731 ( .A(n28974), .B(n28973), .Z(n29026) );
  NANDN U29732 ( .A(n28975), .B(n42231), .Z(n28977) );
  XOR U29733 ( .A(n220), .B(a[699]), .Z(n29016) );
  NANDN U29734 ( .A(n29016), .B(n42234), .Z(n28976) );
  AND U29735 ( .A(n28977), .B(n28976), .Z(n29025) );
  XNOR U29736 ( .A(n29026), .B(n29025), .Z(n29027) );
  XNOR U29737 ( .A(n29028), .B(n29027), .Z(n29032) );
  NANDN U29738 ( .A(n28979), .B(n28978), .Z(n28983) );
  NAND U29739 ( .A(n28981), .B(n28980), .Z(n28982) );
  AND U29740 ( .A(n28983), .B(n28982), .Z(n29031) );
  XOR U29741 ( .A(n29032), .B(n29031), .Z(n29033) );
  NANDN U29742 ( .A(n28985), .B(n28984), .Z(n28989) );
  NANDN U29743 ( .A(n28987), .B(n28986), .Z(n28988) );
  NAND U29744 ( .A(n28989), .B(n28988), .Z(n29034) );
  XOR U29745 ( .A(n29033), .B(n29034), .Z(n29001) );
  OR U29746 ( .A(n28991), .B(n28990), .Z(n28995) );
  NANDN U29747 ( .A(n28993), .B(n28992), .Z(n28994) );
  NAND U29748 ( .A(n28995), .B(n28994), .Z(n29002) );
  XNOR U29749 ( .A(n29001), .B(n29002), .Z(n29003) );
  XNOR U29750 ( .A(n29004), .B(n29003), .Z(n29037) );
  XNOR U29751 ( .A(n29037), .B(sreg[1721]), .Z(n29039) );
  NAND U29752 ( .A(n28996), .B(sreg[1720]), .Z(n29000) );
  OR U29753 ( .A(n28998), .B(n28997), .Z(n28999) );
  AND U29754 ( .A(n29000), .B(n28999), .Z(n29038) );
  XOR U29755 ( .A(n29039), .B(n29038), .Z(c[1721]) );
  NANDN U29756 ( .A(n29002), .B(n29001), .Z(n29006) );
  NAND U29757 ( .A(n29004), .B(n29003), .Z(n29005) );
  NAND U29758 ( .A(n29006), .B(n29005), .Z(n29045) );
  NAND U29759 ( .A(b[0]), .B(a[706]), .Z(n29007) );
  XNOR U29760 ( .A(b[1]), .B(n29007), .Z(n29009) );
  NAND U29761 ( .A(n115), .B(a[705]), .Z(n29008) );
  AND U29762 ( .A(n29009), .B(n29008), .Z(n29062) );
  XOR U29763 ( .A(a[702]), .B(n42197), .Z(n29051) );
  NANDN U29764 ( .A(n29051), .B(n42173), .Z(n29012) );
  NANDN U29765 ( .A(n29010), .B(n42172), .Z(n29011) );
  NAND U29766 ( .A(n29012), .B(n29011), .Z(n29060) );
  NAND U29767 ( .A(b[7]), .B(a[698]), .Z(n29061) );
  XNOR U29768 ( .A(n29060), .B(n29061), .Z(n29063) );
  XOR U29769 ( .A(n29062), .B(n29063), .Z(n29069) );
  NANDN U29770 ( .A(n29013), .B(n42093), .Z(n29015) );
  XOR U29771 ( .A(n42134), .B(a[704]), .Z(n29054) );
  NANDN U29772 ( .A(n29054), .B(n42095), .Z(n29014) );
  NAND U29773 ( .A(n29015), .B(n29014), .Z(n29067) );
  NANDN U29774 ( .A(n29016), .B(n42231), .Z(n29018) );
  XOR U29775 ( .A(n220), .B(a[700]), .Z(n29057) );
  NANDN U29776 ( .A(n29057), .B(n42234), .Z(n29017) );
  AND U29777 ( .A(n29018), .B(n29017), .Z(n29066) );
  XNOR U29778 ( .A(n29067), .B(n29066), .Z(n29068) );
  XNOR U29779 ( .A(n29069), .B(n29068), .Z(n29073) );
  NANDN U29780 ( .A(n29020), .B(n29019), .Z(n29024) );
  NAND U29781 ( .A(n29022), .B(n29021), .Z(n29023) );
  AND U29782 ( .A(n29024), .B(n29023), .Z(n29072) );
  XOR U29783 ( .A(n29073), .B(n29072), .Z(n29074) );
  NANDN U29784 ( .A(n29026), .B(n29025), .Z(n29030) );
  NANDN U29785 ( .A(n29028), .B(n29027), .Z(n29029) );
  NAND U29786 ( .A(n29030), .B(n29029), .Z(n29075) );
  XOR U29787 ( .A(n29074), .B(n29075), .Z(n29042) );
  OR U29788 ( .A(n29032), .B(n29031), .Z(n29036) );
  NANDN U29789 ( .A(n29034), .B(n29033), .Z(n29035) );
  NAND U29790 ( .A(n29036), .B(n29035), .Z(n29043) );
  XNOR U29791 ( .A(n29042), .B(n29043), .Z(n29044) );
  XNOR U29792 ( .A(n29045), .B(n29044), .Z(n29078) );
  XNOR U29793 ( .A(n29078), .B(sreg[1722]), .Z(n29080) );
  NAND U29794 ( .A(n29037), .B(sreg[1721]), .Z(n29041) );
  OR U29795 ( .A(n29039), .B(n29038), .Z(n29040) );
  AND U29796 ( .A(n29041), .B(n29040), .Z(n29079) );
  XOR U29797 ( .A(n29080), .B(n29079), .Z(c[1722]) );
  NANDN U29798 ( .A(n29043), .B(n29042), .Z(n29047) );
  NAND U29799 ( .A(n29045), .B(n29044), .Z(n29046) );
  NAND U29800 ( .A(n29047), .B(n29046), .Z(n29086) );
  NAND U29801 ( .A(b[0]), .B(a[707]), .Z(n29048) );
  XNOR U29802 ( .A(b[1]), .B(n29048), .Z(n29050) );
  NAND U29803 ( .A(n116), .B(a[706]), .Z(n29049) );
  AND U29804 ( .A(n29050), .B(n29049), .Z(n29103) );
  XOR U29805 ( .A(a[703]), .B(n42197), .Z(n29092) );
  NANDN U29806 ( .A(n29092), .B(n42173), .Z(n29053) );
  NANDN U29807 ( .A(n29051), .B(n42172), .Z(n29052) );
  NAND U29808 ( .A(n29053), .B(n29052), .Z(n29101) );
  NAND U29809 ( .A(b[7]), .B(a[699]), .Z(n29102) );
  XNOR U29810 ( .A(n29101), .B(n29102), .Z(n29104) );
  XOR U29811 ( .A(n29103), .B(n29104), .Z(n29110) );
  NANDN U29812 ( .A(n29054), .B(n42093), .Z(n29056) );
  XOR U29813 ( .A(n42134), .B(a[705]), .Z(n29095) );
  NANDN U29814 ( .A(n29095), .B(n42095), .Z(n29055) );
  NAND U29815 ( .A(n29056), .B(n29055), .Z(n29108) );
  NANDN U29816 ( .A(n29057), .B(n42231), .Z(n29059) );
  XOR U29817 ( .A(n220), .B(a[701]), .Z(n29098) );
  NANDN U29818 ( .A(n29098), .B(n42234), .Z(n29058) );
  AND U29819 ( .A(n29059), .B(n29058), .Z(n29107) );
  XNOR U29820 ( .A(n29108), .B(n29107), .Z(n29109) );
  XNOR U29821 ( .A(n29110), .B(n29109), .Z(n29114) );
  NANDN U29822 ( .A(n29061), .B(n29060), .Z(n29065) );
  NAND U29823 ( .A(n29063), .B(n29062), .Z(n29064) );
  AND U29824 ( .A(n29065), .B(n29064), .Z(n29113) );
  XOR U29825 ( .A(n29114), .B(n29113), .Z(n29115) );
  NANDN U29826 ( .A(n29067), .B(n29066), .Z(n29071) );
  NANDN U29827 ( .A(n29069), .B(n29068), .Z(n29070) );
  NAND U29828 ( .A(n29071), .B(n29070), .Z(n29116) );
  XOR U29829 ( .A(n29115), .B(n29116), .Z(n29083) );
  OR U29830 ( .A(n29073), .B(n29072), .Z(n29077) );
  NANDN U29831 ( .A(n29075), .B(n29074), .Z(n29076) );
  NAND U29832 ( .A(n29077), .B(n29076), .Z(n29084) );
  XNOR U29833 ( .A(n29083), .B(n29084), .Z(n29085) );
  XNOR U29834 ( .A(n29086), .B(n29085), .Z(n29119) );
  XNOR U29835 ( .A(n29119), .B(sreg[1723]), .Z(n29121) );
  NAND U29836 ( .A(n29078), .B(sreg[1722]), .Z(n29082) );
  OR U29837 ( .A(n29080), .B(n29079), .Z(n29081) );
  AND U29838 ( .A(n29082), .B(n29081), .Z(n29120) );
  XOR U29839 ( .A(n29121), .B(n29120), .Z(c[1723]) );
  NANDN U29840 ( .A(n29084), .B(n29083), .Z(n29088) );
  NAND U29841 ( .A(n29086), .B(n29085), .Z(n29087) );
  NAND U29842 ( .A(n29088), .B(n29087), .Z(n29127) );
  NAND U29843 ( .A(b[0]), .B(a[708]), .Z(n29089) );
  XNOR U29844 ( .A(b[1]), .B(n29089), .Z(n29091) );
  NAND U29845 ( .A(n116), .B(a[707]), .Z(n29090) );
  AND U29846 ( .A(n29091), .B(n29090), .Z(n29144) );
  XOR U29847 ( .A(a[704]), .B(n42197), .Z(n29133) );
  NANDN U29848 ( .A(n29133), .B(n42173), .Z(n29094) );
  NANDN U29849 ( .A(n29092), .B(n42172), .Z(n29093) );
  NAND U29850 ( .A(n29094), .B(n29093), .Z(n29142) );
  NAND U29851 ( .A(b[7]), .B(a[700]), .Z(n29143) );
  XNOR U29852 ( .A(n29142), .B(n29143), .Z(n29145) );
  XOR U29853 ( .A(n29144), .B(n29145), .Z(n29151) );
  NANDN U29854 ( .A(n29095), .B(n42093), .Z(n29097) );
  XOR U29855 ( .A(n42134), .B(a[706]), .Z(n29136) );
  NANDN U29856 ( .A(n29136), .B(n42095), .Z(n29096) );
  NAND U29857 ( .A(n29097), .B(n29096), .Z(n29149) );
  NANDN U29858 ( .A(n29098), .B(n42231), .Z(n29100) );
  XOR U29859 ( .A(n220), .B(a[702]), .Z(n29139) );
  NANDN U29860 ( .A(n29139), .B(n42234), .Z(n29099) );
  AND U29861 ( .A(n29100), .B(n29099), .Z(n29148) );
  XNOR U29862 ( .A(n29149), .B(n29148), .Z(n29150) );
  XNOR U29863 ( .A(n29151), .B(n29150), .Z(n29155) );
  NANDN U29864 ( .A(n29102), .B(n29101), .Z(n29106) );
  NAND U29865 ( .A(n29104), .B(n29103), .Z(n29105) );
  AND U29866 ( .A(n29106), .B(n29105), .Z(n29154) );
  XOR U29867 ( .A(n29155), .B(n29154), .Z(n29156) );
  NANDN U29868 ( .A(n29108), .B(n29107), .Z(n29112) );
  NANDN U29869 ( .A(n29110), .B(n29109), .Z(n29111) );
  NAND U29870 ( .A(n29112), .B(n29111), .Z(n29157) );
  XOR U29871 ( .A(n29156), .B(n29157), .Z(n29124) );
  OR U29872 ( .A(n29114), .B(n29113), .Z(n29118) );
  NANDN U29873 ( .A(n29116), .B(n29115), .Z(n29117) );
  NAND U29874 ( .A(n29118), .B(n29117), .Z(n29125) );
  XNOR U29875 ( .A(n29124), .B(n29125), .Z(n29126) );
  XNOR U29876 ( .A(n29127), .B(n29126), .Z(n29160) );
  XNOR U29877 ( .A(n29160), .B(sreg[1724]), .Z(n29162) );
  NAND U29878 ( .A(n29119), .B(sreg[1723]), .Z(n29123) );
  OR U29879 ( .A(n29121), .B(n29120), .Z(n29122) );
  AND U29880 ( .A(n29123), .B(n29122), .Z(n29161) );
  XOR U29881 ( .A(n29162), .B(n29161), .Z(c[1724]) );
  NANDN U29882 ( .A(n29125), .B(n29124), .Z(n29129) );
  NAND U29883 ( .A(n29127), .B(n29126), .Z(n29128) );
  NAND U29884 ( .A(n29129), .B(n29128), .Z(n29168) );
  NAND U29885 ( .A(b[0]), .B(a[709]), .Z(n29130) );
  XNOR U29886 ( .A(b[1]), .B(n29130), .Z(n29132) );
  NAND U29887 ( .A(n116), .B(a[708]), .Z(n29131) );
  AND U29888 ( .A(n29132), .B(n29131), .Z(n29185) );
  XOR U29889 ( .A(a[705]), .B(n42197), .Z(n29174) );
  NANDN U29890 ( .A(n29174), .B(n42173), .Z(n29135) );
  NANDN U29891 ( .A(n29133), .B(n42172), .Z(n29134) );
  NAND U29892 ( .A(n29135), .B(n29134), .Z(n29183) );
  NAND U29893 ( .A(b[7]), .B(a[701]), .Z(n29184) );
  XNOR U29894 ( .A(n29183), .B(n29184), .Z(n29186) );
  XOR U29895 ( .A(n29185), .B(n29186), .Z(n29192) );
  NANDN U29896 ( .A(n29136), .B(n42093), .Z(n29138) );
  XOR U29897 ( .A(n42134), .B(a[707]), .Z(n29177) );
  NANDN U29898 ( .A(n29177), .B(n42095), .Z(n29137) );
  NAND U29899 ( .A(n29138), .B(n29137), .Z(n29190) );
  NANDN U29900 ( .A(n29139), .B(n42231), .Z(n29141) );
  XOR U29901 ( .A(n220), .B(a[703]), .Z(n29180) );
  NANDN U29902 ( .A(n29180), .B(n42234), .Z(n29140) );
  AND U29903 ( .A(n29141), .B(n29140), .Z(n29189) );
  XNOR U29904 ( .A(n29190), .B(n29189), .Z(n29191) );
  XNOR U29905 ( .A(n29192), .B(n29191), .Z(n29196) );
  NANDN U29906 ( .A(n29143), .B(n29142), .Z(n29147) );
  NAND U29907 ( .A(n29145), .B(n29144), .Z(n29146) );
  AND U29908 ( .A(n29147), .B(n29146), .Z(n29195) );
  XOR U29909 ( .A(n29196), .B(n29195), .Z(n29197) );
  NANDN U29910 ( .A(n29149), .B(n29148), .Z(n29153) );
  NANDN U29911 ( .A(n29151), .B(n29150), .Z(n29152) );
  NAND U29912 ( .A(n29153), .B(n29152), .Z(n29198) );
  XOR U29913 ( .A(n29197), .B(n29198), .Z(n29165) );
  OR U29914 ( .A(n29155), .B(n29154), .Z(n29159) );
  NANDN U29915 ( .A(n29157), .B(n29156), .Z(n29158) );
  NAND U29916 ( .A(n29159), .B(n29158), .Z(n29166) );
  XNOR U29917 ( .A(n29165), .B(n29166), .Z(n29167) );
  XNOR U29918 ( .A(n29168), .B(n29167), .Z(n29201) );
  XNOR U29919 ( .A(n29201), .B(sreg[1725]), .Z(n29203) );
  NAND U29920 ( .A(n29160), .B(sreg[1724]), .Z(n29164) );
  OR U29921 ( .A(n29162), .B(n29161), .Z(n29163) );
  AND U29922 ( .A(n29164), .B(n29163), .Z(n29202) );
  XOR U29923 ( .A(n29203), .B(n29202), .Z(c[1725]) );
  NANDN U29924 ( .A(n29166), .B(n29165), .Z(n29170) );
  NAND U29925 ( .A(n29168), .B(n29167), .Z(n29169) );
  NAND U29926 ( .A(n29170), .B(n29169), .Z(n29209) );
  NAND U29927 ( .A(b[0]), .B(a[710]), .Z(n29171) );
  XNOR U29928 ( .A(b[1]), .B(n29171), .Z(n29173) );
  NAND U29929 ( .A(n116), .B(a[709]), .Z(n29172) );
  AND U29930 ( .A(n29173), .B(n29172), .Z(n29226) );
  XOR U29931 ( .A(a[706]), .B(n42197), .Z(n29215) );
  NANDN U29932 ( .A(n29215), .B(n42173), .Z(n29176) );
  NANDN U29933 ( .A(n29174), .B(n42172), .Z(n29175) );
  NAND U29934 ( .A(n29176), .B(n29175), .Z(n29224) );
  NAND U29935 ( .A(b[7]), .B(a[702]), .Z(n29225) );
  XNOR U29936 ( .A(n29224), .B(n29225), .Z(n29227) );
  XOR U29937 ( .A(n29226), .B(n29227), .Z(n29233) );
  NANDN U29938 ( .A(n29177), .B(n42093), .Z(n29179) );
  XOR U29939 ( .A(n42134), .B(a[708]), .Z(n29218) );
  NANDN U29940 ( .A(n29218), .B(n42095), .Z(n29178) );
  NAND U29941 ( .A(n29179), .B(n29178), .Z(n29231) );
  NANDN U29942 ( .A(n29180), .B(n42231), .Z(n29182) );
  XOR U29943 ( .A(n220), .B(a[704]), .Z(n29221) );
  NANDN U29944 ( .A(n29221), .B(n42234), .Z(n29181) );
  AND U29945 ( .A(n29182), .B(n29181), .Z(n29230) );
  XNOR U29946 ( .A(n29231), .B(n29230), .Z(n29232) );
  XNOR U29947 ( .A(n29233), .B(n29232), .Z(n29237) );
  NANDN U29948 ( .A(n29184), .B(n29183), .Z(n29188) );
  NAND U29949 ( .A(n29186), .B(n29185), .Z(n29187) );
  AND U29950 ( .A(n29188), .B(n29187), .Z(n29236) );
  XOR U29951 ( .A(n29237), .B(n29236), .Z(n29238) );
  NANDN U29952 ( .A(n29190), .B(n29189), .Z(n29194) );
  NANDN U29953 ( .A(n29192), .B(n29191), .Z(n29193) );
  NAND U29954 ( .A(n29194), .B(n29193), .Z(n29239) );
  XOR U29955 ( .A(n29238), .B(n29239), .Z(n29206) );
  OR U29956 ( .A(n29196), .B(n29195), .Z(n29200) );
  NANDN U29957 ( .A(n29198), .B(n29197), .Z(n29199) );
  NAND U29958 ( .A(n29200), .B(n29199), .Z(n29207) );
  XNOR U29959 ( .A(n29206), .B(n29207), .Z(n29208) );
  XNOR U29960 ( .A(n29209), .B(n29208), .Z(n29242) );
  XNOR U29961 ( .A(n29242), .B(sreg[1726]), .Z(n29244) );
  NAND U29962 ( .A(n29201), .B(sreg[1725]), .Z(n29205) );
  OR U29963 ( .A(n29203), .B(n29202), .Z(n29204) );
  AND U29964 ( .A(n29205), .B(n29204), .Z(n29243) );
  XOR U29965 ( .A(n29244), .B(n29243), .Z(c[1726]) );
  NANDN U29966 ( .A(n29207), .B(n29206), .Z(n29211) );
  NAND U29967 ( .A(n29209), .B(n29208), .Z(n29210) );
  NAND U29968 ( .A(n29211), .B(n29210), .Z(n29250) );
  NAND U29969 ( .A(b[0]), .B(a[711]), .Z(n29212) );
  XNOR U29970 ( .A(b[1]), .B(n29212), .Z(n29214) );
  NAND U29971 ( .A(n116), .B(a[710]), .Z(n29213) );
  AND U29972 ( .A(n29214), .B(n29213), .Z(n29267) );
  XOR U29973 ( .A(a[707]), .B(n42197), .Z(n29256) );
  NANDN U29974 ( .A(n29256), .B(n42173), .Z(n29217) );
  NANDN U29975 ( .A(n29215), .B(n42172), .Z(n29216) );
  NAND U29976 ( .A(n29217), .B(n29216), .Z(n29265) );
  NAND U29977 ( .A(b[7]), .B(a[703]), .Z(n29266) );
  XNOR U29978 ( .A(n29265), .B(n29266), .Z(n29268) );
  XOR U29979 ( .A(n29267), .B(n29268), .Z(n29274) );
  NANDN U29980 ( .A(n29218), .B(n42093), .Z(n29220) );
  XOR U29981 ( .A(n42134), .B(a[709]), .Z(n29259) );
  NANDN U29982 ( .A(n29259), .B(n42095), .Z(n29219) );
  NAND U29983 ( .A(n29220), .B(n29219), .Z(n29272) );
  NANDN U29984 ( .A(n29221), .B(n42231), .Z(n29223) );
  XOR U29985 ( .A(n220), .B(a[705]), .Z(n29262) );
  NANDN U29986 ( .A(n29262), .B(n42234), .Z(n29222) );
  AND U29987 ( .A(n29223), .B(n29222), .Z(n29271) );
  XNOR U29988 ( .A(n29272), .B(n29271), .Z(n29273) );
  XNOR U29989 ( .A(n29274), .B(n29273), .Z(n29278) );
  NANDN U29990 ( .A(n29225), .B(n29224), .Z(n29229) );
  NAND U29991 ( .A(n29227), .B(n29226), .Z(n29228) );
  AND U29992 ( .A(n29229), .B(n29228), .Z(n29277) );
  XOR U29993 ( .A(n29278), .B(n29277), .Z(n29279) );
  NANDN U29994 ( .A(n29231), .B(n29230), .Z(n29235) );
  NANDN U29995 ( .A(n29233), .B(n29232), .Z(n29234) );
  NAND U29996 ( .A(n29235), .B(n29234), .Z(n29280) );
  XOR U29997 ( .A(n29279), .B(n29280), .Z(n29247) );
  OR U29998 ( .A(n29237), .B(n29236), .Z(n29241) );
  NANDN U29999 ( .A(n29239), .B(n29238), .Z(n29240) );
  NAND U30000 ( .A(n29241), .B(n29240), .Z(n29248) );
  XNOR U30001 ( .A(n29247), .B(n29248), .Z(n29249) );
  XNOR U30002 ( .A(n29250), .B(n29249), .Z(n29283) );
  XNOR U30003 ( .A(n29283), .B(sreg[1727]), .Z(n29285) );
  NAND U30004 ( .A(n29242), .B(sreg[1726]), .Z(n29246) );
  OR U30005 ( .A(n29244), .B(n29243), .Z(n29245) );
  AND U30006 ( .A(n29246), .B(n29245), .Z(n29284) );
  XOR U30007 ( .A(n29285), .B(n29284), .Z(c[1727]) );
  NANDN U30008 ( .A(n29248), .B(n29247), .Z(n29252) );
  NAND U30009 ( .A(n29250), .B(n29249), .Z(n29251) );
  NAND U30010 ( .A(n29252), .B(n29251), .Z(n29291) );
  NAND U30011 ( .A(b[0]), .B(a[712]), .Z(n29253) );
  XNOR U30012 ( .A(b[1]), .B(n29253), .Z(n29255) );
  NAND U30013 ( .A(n116), .B(a[711]), .Z(n29254) );
  AND U30014 ( .A(n29255), .B(n29254), .Z(n29308) );
  XOR U30015 ( .A(a[708]), .B(n42197), .Z(n29297) );
  NANDN U30016 ( .A(n29297), .B(n42173), .Z(n29258) );
  NANDN U30017 ( .A(n29256), .B(n42172), .Z(n29257) );
  NAND U30018 ( .A(n29258), .B(n29257), .Z(n29306) );
  NAND U30019 ( .A(b[7]), .B(a[704]), .Z(n29307) );
  XNOR U30020 ( .A(n29306), .B(n29307), .Z(n29309) );
  XOR U30021 ( .A(n29308), .B(n29309), .Z(n29315) );
  NANDN U30022 ( .A(n29259), .B(n42093), .Z(n29261) );
  XOR U30023 ( .A(n42134), .B(a[710]), .Z(n29300) );
  NANDN U30024 ( .A(n29300), .B(n42095), .Z(n29260) );
  NAND U30025 ( .A(n29261), .B(n29260), .Z(n29313) );
  NANDN U30026 ( .A(n29262), .B(n42231), .Z(n29264) );
  XOR U30027 ( .A(n220), .B(a[706]), .Z(n29303) );
  NANDN U30028 ( .A(n29303), .B(n42234), .Z(n29263) );
  AND U30029 ( .A(n29264), .B(n29263), .Z(n29312) );
  XNOR U30030 ( .A(n29313), .B(n29312), .Z(n29314) );
  XNOR U30031 ( .A(n29315), .B(n29314), .Z(n29319) );
  NANDN U30032 ( .A(n29266), .B(n29265), .Z(n29270) );
  NAND U30033 ( .A(n29268), .B(n29267), .Z(n29269) );
  AND U30034 ( .A(n29270), .B(n29269), .Z(n29318) );
  XOR U30035 ( .A(n29319), .B(n29318), .Z(n29320) );
  NANDN U30036 ( .A(n29272), .B(n29271), .Z(n29276) );
  NANDN U30037 ( .A(n29274), .B(n29273), .Z(n29275) );
  NAND U30038 ( .A(n29276), .B(n29275), .Z(n29321) );
  XOR U30039 ( .A(n29320), .B(n29321), .Z(n29288) );
  OR U30040 ( .A(n29278), .B(n29277), .Z(n29282) );
  NANDN U30041 ( .A(n29280), .B(n29279), .Z(n29281) );
  NAND U30042 ( .A(n29282), .B(n29281), .Z(n29289) );
  XNOR U30043 ( .A(n29288), .B(n29289), .Z(n29290) );
  XNOR U30044 ( .A(n29291), .B(n29290), .Z(n29324) );
  XNOR U30045 ( .A(n29324), .B(sreg[1728]), .Z(n29326) );
  NAND U30046 ( .A(n29283), .B(sreg[1727]), .Z(n29287) );
  OR U30047 ( .A(n29285), .B(n29284), .Z(n29286) );
  AND U30048 ( .A(n29287), .B(n29286), .Z(n29325) );
  XOR U30049 ( .A(n29326), .B(n29325), .Z(c[1728]) );
  NANDN U30050 ( .A(n29289), .B(n29288), .Z(n29293) );
  NAND U30051 ( .A(n29291), .B(n29290), .Z(n29292) );
  NAND U30052 ( .A(n29293), .B(n29292), .Z(n29332) );
  NAND U30053 ( .A(b[0]), .B(a[713]), .Z(n29294) );
  XNOR U30054 ( .A(b[1]), .B(n29294), .Z(n29296) );
  NAND U30055 ( .A(n116), .B(a[712]), .Z(n29295) );
  AND U30056 ( .A(n29296), .B(n29295), .Z(n29349) );
  XOR U30057 ( .A(a[709]), .B(n42197), .Z(n29338) );
  NANDN U30058 ( .A(n29338), .B(n42173), .Z(n29299) );
  NANDN U30059 ( .A(n29297), .B(n42172), .Z(n29298) );
  NAND U30060 ( .A(n29299), .B(n29298), .Z(n29347) );
  NAND U30061 ( .A(b[7]), .B(a[705]), .Z(n29348) );
  XNOR U30062 ( .A(n29347), .B(n29348), .Z(n29350) );
  XOR U30063 ( .A(n29349), .B(n29350), .Z(n29356) );
  NANDN U30064 ( .A(n29300), .B(n42093), .Z(n29302) );
  XOR U30065 ( .A(n42134), .B(a[711]), .Z(n29341) );
  NANDN U30066 ( .A(n29341), .B(n42095), .Z(n29301) );
  NAND U30067 ( .A(n29302), .B(n29301), .Z(n29354) );
  NANDN U30068 ( .A(n29303), .B(n42231), .Z(n29305) );
  XOR U30069 ( .A(n221), .B(a[707]), .Z(n29344) );
  NANDN U30070 ( .A(n29344), .B(n42234), .Z(n29304) );
  AND U30071 ( .A(n29305), .B(n29304), .Z(n29353) );
  XNOR U30072 ( .A(n29354), .B(n29353), .Z(n29355) );
  XNOR U30073 ( .A(n29356), .B(n29355), .Z(n29360) );
  NANDN U30074 ( .A(n29307), .B(n29306), .Z(n29311) );
  NAND U30075 ( .A(n29309), .B(n29308), .Z(n29310) );
  AND U30076 ( .A(n29311), .B(n29310), .Z(n29359) );
  XOR U30077 ( .A(n29360), .B(n29359), .Z(n29361) );
  NANDN U30078 ( .A(n29313), .B(n29312), .Z(n29317) );
  NANDN U30079 ( .A(n29315), .B(n29314), .Z(n29316) );
  NAND U30080 ( .A(n29317), .B(n29316), .Z(n29362) );
  XOR U30081 ( .A(n29361), .B(n29362), .Z(n29329) );
  OR U30082 ( .A(n29319), .B(n29318), .Z(n29323) );
  NANDN U30083 ( .A(n29321), .B(n29320), .Z(n29322) );
  NAND U30084 ( .A(n29323), .B(n29322), .Z(n29330) );
  XNOR U30085 ( .A(n29329), .B(n29330), .Z(n29331) );
  XNOR U30086 ( .A(n29332), .B(n29331), .Z(n29365) );
  XNOR U30087 ( .A(n29365), .B(sreg[1729]), .Z(n29367) );
  NAND U30088 ( .A(n29324), .B(sreg[1728]), .Z(n29328) );
  OR U30089 ( .A(n29326), .B(n29325), .Z(n29327) );
  AND U30090 ( .A(n29328), .B(n29327), .Z(n29366) );
  XOR U30091 ( .A(n29367), .B(n29366), .Z(c[1729]) );
  NANDN U30092 ( .A(n29330), .B(n29329), .Z(n29334) );
  NAND U30093 ( .A(n29332), .B(n29331), .Z(n29333) );
  NAND U30094 ( .A(n29334), .B(n29333), .Z(n29373) );
  NAND U30095 ( .A(b[0]), .B(a[714]), .Z(n29335) );
  XNOR U30096 ( .A(b[1]), .B(n29335), .Z(n29337) );
  NAND U30097 ( .A(n117), .B(a[713]), .Z(n29336) );
  AND U30098 ( .A(n29337), .B(n29336), .Z(n29390) );
  XOR U30099 ( .A(a[710]), .B(n42197), .Z(n29379) );
  NANDN U30100 ( .A(n29379), .B(n42173), .Z(n29340) );
  NANDN U30101 ( .A(n29338), .B(n42172), .Z(n29339) );
  NAND U30102 ( .A(n29340), .B(n29339), .Z(n29388) );
  NAND U30103 ( .A(b[7]), .B(a[706]), .Z(n29389) );
  XNOR U30104 ( .A(n29388), .B(n29389), .Z(n29391) );
  XOR U30105 ( .A(n29390), .B(n29391), .Z(n29397) );
  NANDN U30106 ( .A(n29341), .B(n42093), .Z(n29343) );
  XOR U30107 ( .A(n42134), .B(a[712]), .Z(n29382) );
  NANDN U30108 ( .A(n29382), .B(n42095), .Z(n29342) );
  NAND U30109 ( .A(n29343), .B(n29342), .Z(n29395) );
  NANDN U30110 ( .A(n29344), .B(n42231), .Z(n29346) );
  XOR U30111 ( .A(n221), .B(a[708]), .Z(n29385) );
  NANDN U30112 ( .A(n29385), .B(n42234), .Z(n29345) );
  AND U30113 ( .A(n29346), .B(n29345), .Z(n29394) );
  XNOR U30114 ( .A(n29395), .B(n29394), .Z(n29396) );
  XNOR U30115 ( .A(n29397), .B(n29396), .Z(n29401) );
  NANDN U30116 ( .A(n29348), .B(n29347), .Z(n29352) );
  NAND U30117 ( .A(n29350), .B(n29349), .Z(n29351) );
  AND U30118 ( .A(n29352), .B(n29351), .Z(n29400) );
  XOR U30119 ( .A(n29401), .B(n29400), .Z(n29402) );
  NANDN U30120 ( .A(n29354), .B(n29353), .Z(n29358) );
  NANDN U30121 ( .A(n29356), .B(n29355), .Z(n29357) );
  NAND U30122 ( .A(n29358), .B(n29357), .Z(n29403) );
  XOR U30123 ( .A(n29402), .B(n29403), .Z(n29370) );
  OR U30124 ( .A(n29360), .B(n29359), .Z(n29364) );
  NANDN U30125 ( .A(n29362), .B(n29361), .Z(n29363) );
  NAND U30126 ( .A(n29364), .B(n29363), .Z(n29371) );
  XNOR U30127 ( .A(n29370), .B(n29371), .Z(n29372) );
  XNOR U30128 ( .A(n29373), .B(n29372), .Z(n29406) );
  XNOR U30129 ( .A(n29406), .B(sreg[1730]), .Z(n29408) );
  NAND U30130 ( .A(n29365), .B(sreg[1729]), .Z(n29369) );
  OR U30131 ( .A(n29367), .B(n29366), .Z(n29368) );
  AND U30132 ( .A(n29369), .B(n29368), .Z(n29407) );
  XOR U30133 ( .A(n29408), .B(n29407), .Z(c[1730]) );
  NANDN U30134 ( .A(n29371), .B(n29370), .Z(n29375) );
  NAND U30135 ( .A(n29373), .B(n29372), .Z(n29374) );
  NAND U30136 ( .A(n29375), .B(n29374), .Z(n29414) );
  NAND U30137 ( .A(b[0]), .B(a[715]), .Z(n29376) );
  XNOR U30138 ( .A(b[1]), .B(n29376), .Z(n29378) );
  NAND U30139 ( .A(n117), .B(a[714]), .Z(n29377) );
  AND U30140 ( .A(n29378), .B(n29377), .Z(n29431) );
  XOR U30141 ( .A(a[711]), .B(n42197), .Z(n29420) );
  NANDN U30142 ( .A(n29420), .B(n42173), .Z(n29381) );
  NANDN U30143 ( .A(n29379), .B(n42172), .Z(n29380) );
  NAND U30144 ( .A(n29381), .B(n29380), .Z(n29429) );
  NAND U30145 ( .A(b[7]), .B(a[707]), .Z(n29430) );
  XNOR U30146 ( .A(n29429), .B(n29430), .Z(n29432) );
  XOR U30147 ( .A(n29431), .B(n29432), .Z(n29438) );
  NANDN U30148 ( .A(n29382), .B(n42093), .Z(n29384) );
  XOR U30149 ( .A(n42134), .B(a[713]), .Z(n29423) );
  NANDN U30150 ( .A(n29423), .B(n42095), .Z(n29383) );
  NAND U30151 ( .A(n29384), .B(n29383), .Z(n29436) );
  NANDN U30152 ( .A(n29385), .B(n42231), .Z(n29387) );
  XOR U30153 ( .A(n221), .B(a[709]), .Z(n29426) );
  NANDN U30154 ( .A(n29426), .B(n42234), .Z(n29386) );
  AND U30155 ( .A(n29387), .B(n29386), .Z(n29435) );
  XNOR U30156 ( .A(n29436), .B(n29435), .Z(n29437) );
  XNOR U30157 ( .A(n29438), .B(n29437), .Z(n29442) );
  NANDN U30158 ( .A(n29389), .B(n29388), .Z(n29393) );
  NAND U30159 ( .A(n29391), .B(n29390), .Z(n29392) );
  AND U30160 ( .A(n29393), .B(n29392), .Z(n29441) );
  XOR U30161 ( .A(n29442), .B(n29441), .Z(n29443) );
  NANDN U30162 ( .A(n29395), .B(n29394), .Z(n29399) );
  NANDN U30163 ( .A(n29397), .B(n29396), .Z(n29398) );
  NAND U30164 ( .A(n29399), .B(n29398), .Z(n29444) );
  XOR U30165 ( .A(n29443), .B(n29444), .Z(n29411) );
  OR U30166 ( .A(n29401), .B(n29400), .Z(n29405) );
  NANDN U30167 ( .A(n29403), .B(n29402), .Z(n29404) );
  NAND U30168 ( .A(n29405), .B(n29404), .Z(n29412) );
  XNOR U30169 ( .A(n29411), .B(n29412), .Z(n29413) );
  XNOR U30170 ( .A(n29414), .B(n29413), .Z(n29447) );
  XNOR U30171 ( .A(n29447), .B(sreg[1731]), .Z(n29449) );
  NAND U30172 ( .A(n29406), .B(sreg[1730]), .Z(n29410) );
  OR U30173 ( .A(n29408), .B(n29407), .Z(n29409) );
  AND U30174 ( .A(n29410), .B(n29409), .Z(n29448) );
  XOR U30175 ( .A(n29449), .B(n29448), .Z(c[1731]) );
  NANDN U30176 ( .A(n29412), .B(n29411), .Z(n29416) );
  NAND U30177 ( .A(n29414), .B(n29413), .Z(n29415) );
  NAND U30178 ( .A(n29416), .B(n29415), .Z(n29455) );
  NAND U30179 ( .A(b[0]), .B(a[716]), .Z(n29417) );
  XNOR U30180 ( .A(b[1]), .B(n29417), .Z(n29419) );
  NAND U30181 ( .A(n117), .B(a[715]), .Z(n29418) );
  AND U30182 ( .A(n29419), .B(n29418), .Z(n29472) );
  XOR U30183 ( .A(a[712]), .B(n42197), .Z(n29461) );
  NANDN U30184 ( .A(n29461), .B(n42173), .Z(n29422) );
  NANDN U30185 ( .A(n29420), .B(n42172), .Z(n29421) );
  NAND U30186 ( .A(n29422), .B(n29421), .Z(n29470) );
  NAND U30187 ( .A(b[7]), .B(a[708]), .Z(n29471) );
  XNOR U30188 ( .A(n29470), .B(n29471), .Z(n29473) );
  XOR U30189 ( .A(n29472), .B(n29473), .Z(n29479) );
  NANDN U30190 ( .A(n29423), .B(n42093), .Z(n29425) );
  XOR U30191 ( .A(n42134), .B(a[714]), .Z(n29464) );
  NANDN U30192 ( .A(n29464), .B(n42095), .Z(n29424) );
  NAND U30193 ( .A(n29425), .B(n29424), .Z(n29477) );
  NANDN U30194 ( .A(n29426), .B(n42231), .Z(n29428) );
  XOR U30195 ( .A(n221), .B(a[710]), .Z(n29467) );
  NANDN U30196 ( .A(n29467), .B(n42234), .Z(n29427) );
  AND U30197 ( .A(n29428), .B(n29427), .Z(n29476) );
  XNOR U30198 ( .A(n29477), .B(n29476), .Z(n29478) );
  XNOR U30199 ( .A(n29479), .B(n29478), .Z(n29483) );
  NANDN U30200 ( .A(n29430), .B(n29429), .Z(n29434) );
  NAND U30201 ( .A(n29432), .B(n29431), .Z(n29433) );
  AND U30202 ( .A(n29434), .B(n29433), .Z(n29482) );
  XOR U30203 ( .A(n29483), .B(n29482), .Z(n29484) );
  NANDN U30204 ( .A(n29436), .B(n29435), .Z(n29440) );
  NANDN U30205 ( .A(n29438), .B(n29437), .Z(n29439) );
  NAND U30206 ( .A(n29440), .B(n29439), .Z(n29485) );
  XOR U30207 ( .A(n29484), .B(n29485), .Z(n29452) );
  OR U30208 ( .A(n29442), .B(n29441), .Z(n29446) );
  NANDN U30209 ( .A(n29444), .B(n29443), .Z(n29445) );
  NAND U30210 ( .A(n29446), .B(n29445), .Z(n29453) );
  XNOR U30211 ( .A(n29452), .B(n29453), .Z(n29454) );
  XNOR U30212 ( .A(n29455), .B(n29454), .Z(n29488) );
  XNOR U30213 ( .A(n29488), .B(sreg[1732]), .Z(n29490) );
  NAND U30214 ( .A(n29447), .B(sreg[1731]), .Z(n29451) );
  OR U30215 ( .A(n29449), .B(n29448), .Z(n29450) );
  AND U30216 ( .A(n29451), .B(n29450), .Z(n29489) );
  XOR U30217 ( .A(n29490), .B(n29489), .Z(c[1732]) );
  NANDN U30218 ( .A(n29453), .B(n29452), .Z(n29457) );
  NAND U30219 ( .A(n29455), .B(n29454), .Z(n29456) );
  NAND U30220 ( .A(n29457), .B(n29456), .Z(n29496) );
  NAND U30221 ( .A(b[0]), .B(a[717]), .Z(n29458) );
  XNOR U30222 ( .A(b[1]), .B(n29458), .Z(n29460) );
  NAND U30223 ( .A(n117), .B(a[716]), .Z(n29459) );
  AND U30224 ( .A(n29460), .B(n29459), .Z(n29513) );
  XOR U30225 ( .A(a[713]), .B(n42197), .Z(n29502) );
  NANDN U30226 ( .A(n29502), .B(n42173), .Z(n29463) );
  NANDN U30227 ( .A(n29461), .B(n42172), .Z(n29462) );
  NAND U30228 ( .A(n29463), .B(n29462), .Z(n29511) );
  NAND U30229 ( .A(b[7]), .B(a[709]), .Z(n29512) );
  XNOR U30230 ( .A(n29511), .B(n29512), .Z(n29514) );
  XOR U30231 ( .A(n29513), .B(n29514), .Z(n29520) );
  NANDN U30232 ( .A(n29464), .B(n42093), .Z(n29466) );
  XOR U30233 ( .A(n42134), .B(a[715]), .Z(n29505) );
  NANDN U30234 ( .A(n29505), .B(n42095), .Z(n29465) );
  NAND U30235 ( .A(n29466), .B(n29465), .Z(n29518) );
  NANDN U30236 ( .A(n29467), .B(n42231), .Z(n29469) );
  XOR U30237 ( .A(n221), .B(a[711]), .Z(n29508) );
  NANDN U30238 ( .A(n29508), .B(n42234), .Z(n29468) );
  AND U30239 ( .A(n29469), .B(n29468), .Z(n29517) );
  XNOR U30240 ( .A(n29518), .B(n29517), .Z(n29519) );
  XNOR U30241 ( .A(n29520), .B(n29519), .Z(n29524) );
  NANDN U30242 ( .A(n29471), .B(n29470), .Z(n29475) );
  NAND U30243 ( .A(n29473), .B(n29472), .Z(n29474) );
  AND U30244 ( .A(n29475), .B(n29474), .Z(n29523) );
  XOR U30245 ( .A(n29524), .B(n29523), .Z(n29525) );
  NANDN U30246 ( .A(n29477), .B(n29476), .Z(n29481) );
  NANDN U30247 ( .A(n29479), .B(n29478), .Z(n29480) );
  NAND U30248 ( .A(n29481), .B(n29480), .Z(n29526) );
  XOR U30249 ( .A(n29525), .B(n29526), .Z(n29493) );
  OR U30250 ( .A(n29483), .B(n29482), .Z(n29487) );
  NANDN U30251 ( .A(n29485), .B(n29484), .Z(n29486) );
  NAND U30252 ( .A(n29487), .B(n29486), .Z(n29494) );
  XNOR U30253 ( .A(n29493), .B(n29494), .Z(n29495) );
  XNOR U30254 ( .A(n29496), .B(n29495), .Z(n29529) );
  XNOR U30255 ( .A(n29529), .B(sreg[1733]), .Z(n29531) );
  NAND U30256 ( .A(n29488), .B(sreg[1732]), .Z(n29492) );
  OR U30257 ( .A(n29490), .B(n29489), .Z(n29491) );
  AND U30258 ( .A(n29492), .B(n29491), .Z(n29530) );
  XOR U30259 ( .A(n29531), .B(n29530), .Z(c[1733]) );
  NANDN U30260 ( .A(n29494), .B(n29493), .Z(n29498) );
  NAND U30261 ( .A(n29496), .B(n29495), .Z(n29497) );
  NAND U30262 ( .A(n29498), .B(n29497), .Z(n29537) );
  NAND U30263 ( .A(b[0]), .B(a[718]), .Z(n29499) );
  XNOR U30264 ( .A(b[1]), .B(n29499), .Z(n29501) );
  NAND U30265 ( .A(n117), .B(a[717]), .Z(n29500) );
  AND U30266 ( .A(n29501), .B(n29500), .Z(n29554) );
  XOR U30267 ( .A(a[714]), .B(n42197), .Z(n29543) );
  NANDN U30268 ( .A(n29543), .B(n42173), .Z(n29504) );
  NANDN U30269 ( .A(n29502), .B(n42172), .Z(n29503) );
  NAND U30270 ( .A(n29504), .B(n29503), .Z(n29552) );
  NAND U30271 ( .A(b[7]), .B(a[710]), .Z(n29553) );
  XNOR U30272 ( .A(n29552), .B(n29553), .Z(n29555) );
  XOR U30273 ( .A(n29554), .B(n29555), .Z(n29561) );
  NANDN U30274 ( .A(n29505), .B(n42093), .Z(n29507) );
  XOR U30275 ( .A(n42134), .B(a[716]), .Z(n29546) );
  NANDN U30276 ( .A(n29546), .B(n42095), .Z(n29506) );
  NAND U30277 ( .A(n29507), .B(n29506), .Z(n29559) );
  NANDN U30278 ( .A(n29508), .B(n42231), .Z(n29510) );
  XOR U30279 ( .A(n221), .B(a[712]), .Z(n29549) );
  NANDN U30280 ( .A(n29549), .B(n42234), .Z(n29509) );
  AND U30281 ( .A(n29510), .B(n29509), .Z(n29558) );
  XNOR U30282 ( .A(n29559), .B(n29558), .Z(n29560) );
  XNOR U30283 ( .A(n29561), .B(n29560), .Z(n29565) );
  NANDN U30284 ( .A(n29512), .B(n29511), .Z(n29516) );
  NAND U30285 ( .A(n29514), .B(n29513), .Z(n29515) );
  AND U30286 ( .A(n29516), .B(n29515), .Z(n29564) );
  XOR U30287 ( .A(n29565), .B(n29564), .Z(n29566) );
  NANDN U30288 ( .A(n29518), .B(n29517), .Z(n29522) );
  NANDN U30289 ( .A(n29520), .B(n29519), .Z(n29521) );
  NAND U30290 ( .A(n29522), .B(n29521), .Z(n29567) );
  XOR U30291 ( .A(n29566), .B(n29567), .Z(n29534) );
  OR U30292 ( .A(n29524), .B(n29523), .Z(n29528) );
  NANDN U30293 ( .A(n29526), .B(n29525), .Z(n29527) );
  NAND U30294 ( .A(n29528), .B(n29527), .Z(n29535) );
  XNOR U30295 ( .A(n29534), .B(n29535), .Z(n29536) );
  XNOR U30296 ( .A(n29537), .B(n29536), .Z(n29570) );
  XNOR U30297 ( .A(n29570), .B(sreg[1734]), .Z(n29572) );
  NAND U30298 ( .A(n29529), .B(sreg[1733]), .Z(n29533) );
  OR U30299 ( .A(n29531), .B(n29530), .Z(n29532) );
  AND U30300 ( .A(n29533), .B(n29532), .Z(n29571) );
  XOR U30301 ( .A(n29572), .B(n29571), .Z(c[1734]) );
  NANDN U30302 ( .A(n29535), .B(n29534), .Z(n29539) );
  NAND U30303 ( .A(n29537), .B(n29536), .Z(n29538) );
  NAND U30304 ( .A(n29539), .B(n29538), .Z(n29578) );
  NAND U30305 ( .A(b[0]), .B(a[719]), .Z(n29540) );
  XNOR U30306 ( .A(b[1]), .B(n29540), .Z(n29542) );
  NAND U30307 ( .A(n117), .B(a[718]), .Z(n29541) );
  AND U30308 ( .A(n29542), .B(n29541), .Z(n29595) );
  XOR U30309 ( .A(a[715]), .B(n42197), .Z(n29584) );
  NANDN U30310 ( .A(n29584), .B(n42173), .Z(n29545) );
  NANDN U30311 ( .A(n29543), .B(n42172), .Z(n29544) );
  NAND U30312 ( .A(n29545), .B(n29544), .Z(n29593) );
  NAND U30313 ( .A(b[7]), .B(a[711]), .Z(n29594) );
  XNOR U30314 ( .A(n29593), .B(n29594), .Z(n29596) );
  XOR U30315 ( .A(n29595), .B(n29596), .Z(n29602) );
  NANDN U30316 ( .A(n29546), .B(n42093), .Z(n29548) );
  XOR U30317 ( .A(n42134), .B(a[717]), .Z(n29587) );
  NANDN U30318 ( .A(n29587), .B(n42095), .Z(n29547) );
  NAND U30319 ( .A(n29548), .B(n29547), .Z(n29600) );
  NANDN U30320 ( .A(n29549), .B(n42231), .Z(n29551) );
  XOR U30321 ( .A(n221), .B(a[713]), .Z(n29590) );
  NANDN U30322 ( .A(n29590), .B(n42234), .Z(n29550) );
  AND U30323 ( .A(n29551), .B(n29550), .Z(n29599) );
  XNOR U30324 ( .A(n29600), .B(n29599), .Z(n29601) );
  XNOR U30325 ( .A(n29602), .B(n29601), .Z(n29606) );
  NANDN U30326 ( .A(n29553), .B(n29552), .Z(n29557) );
  NAND U30327 ( .A(n29555), .B(n29554), .Z(n29556) );
  AND U30328 ( .A(n29557), .B(n29556), .Z(n29605) );
  XOR U30329 ( .A(n29606), .B(n29605), .Z(n29607) );
  NANDN U30330 ( .A(n29559), .B(n29558), .Z(n29563) );
  NANDN U30331 ( .A(n29561), .B(n29560), .Z(n29562) );
  NAND U30332 ( .A(n29563), .B(n29562), .Z(n29608) );
  XOR U30333 ( .A(n29607), .B(n29608), .Z(n29575) );
  OR U30334 ( .A(n29565), .B(n29564), .Z(n29569) );
  NANDN U30335 ( .A(n29567), .B(n29566), .Z(n29568) );
  NAND U30336 ( .A(n29569), .B(n29568), .Z(n29576) );
  XNOR U30337 ( .A(n29575), .B(n29576), .Z(n29577) );
  XNOR U30338 ( .A(n29578), .B(n29577), .Z(n29611) );
  XNOR U30339 ( .A(n29611), .B(sreg[1735]), .Z(n29613) );
  NAND U30340 ( .A(n29570), .B(sreg[1734]), .Z(n29574) );
  OR U30341 ( .A(n29572), .B(n29571), .Z(n29573) );
  AND U30342 ( .A(n29574), .B(n29573), .Z(n29612) );
  XOR U30343 ( .A(n29613), .B(n29612), .Z(c[1735]) );
  NANDN U30344 ( .A(n29576), .B(n29575), .Z(n29580) );
  NAND U30345 ( .A(n29578), .B(n29577), .Z(n29579) );
  NAND U30346 ( .A(n29580), .B(n29579), .Z(n29619) );
  NAND U30347 ( .A(b[0]), .B(a[720]), .Z(n29581) );
  XNOR U30348 ( .A(b[1]), .B(n29581), .Z(n29583) );
  NAND U30349 ( .A(n117), .B(a[719]), .Z(n29582) );
  AND U30350 ( .A(n29583), .B(n29582), .Z(n29636) );
  XOR U30351 ( .A(a[716]), .B(n42197), .Z(n29625) );
  NANDN U30352 ( .A(n29625), .B(n42173), .Z(n29586) );
  NANDN U30353 ( .A(n29584), .B(n42172), .Z(n29585) );
  NAND U30354 ( .A(n29586), .B(n29585), .Z(n29634) );
  NAND U30355 ( .A(b[7]), .B(a[712]), .Z(n29635) );
  XNOR U30356 ( .A(n29634), .B(n29635), .Z(n29637) );
  XOR U30357 ( .A(n29636), .B(n29637), .Z(n29643) );
  NANDN U30358 ( .A(n29587), .B(n42093), .Z(n29589) );
  XOR U30359 ( .A(n42134), .B(a[718]), .Z(n29628) );
  NANDN U30360 ( .A(n29628), .B(n42095), .Z(n29588) );
  NAND U30361 ( .A(n29589), .B(n29588), .Z(n29641) );
  NANDN U30362 ( .A(n29590), .B(n42231), .Z(n29592) );
  XOR U30363 ( .A(n221), .B(a[714]), .Z(n29631) );
  NANDN U30364 ( .A(n29631), .B(n42234), .Z(n29591) );
  AND U30365 ( .A(n29592), .B(n29591), .Z(n29640) );
  XNOR U30366 ( .A(n29641), .B(n29640), .Z(n29642) );
  XNOR U30367 ( .A(n29643), .B(n29642), .Z(n29647) );
  NANDN U30368 ( .A(n29594), .B(n29593), .Z(n29598) );
  NAND U30369 ( .A(n29596), .B(n29595), .Z(n29597) );
  AND U30370 ( .A(n29598), .B(n29597), .Z(n29646) );
  XOR U30371 ( .A(n29647), .B(n29646), .Z(n29648) );
  NANDN U30372 ( .A(n29600), .B(n29599), .Z(n29604) );
  NANDN U30373 ( .A(n29602), .B(n29601), .Z(n29603) );
  NAND U30374 ( .A(n29604), .B(n29603), .Z(n29649) );
  XOR U30375 ( .A(n29648), .B(n29649), .Z(n29616) );
  OR U30376 ( .A(n29606), .B(n29605), .Z(n29610) );
  NANDN U30377 ( .A(n29608), .B(n29607), .Z(n29609) );
  NAND U30378 ( .A(n29610), .B(n29609), .Z(n29617) );
  XNOR U30379 ( .A(n29616), .B(n29617), .Z(n29618) );
  XNOR U30380 ( .A(n29619), .B(n29618), .Z(n29652) );
  XNOR U30381 ( .A(n29652), .B(sreg[1736]), .Z(n29654) );
  NAND U30382 ( .A(n29611), .B(sreg[1735]), .Z(n29615) );
  OR U30383 ( .A(n29613), .B(n29612), .Z(n29614) );
  AND U30384 ( .A(n29615), .B(n29614), .Z(n29653) );
  XOR U30385 ( .A(n29654), .B(n29653), .Z(c[1736]) );
  NANDN U30386 ( .A(n29617), .B(n29616), .Z(n29621) );
  NAND U30387 ( .A(n29619), .B(n29618), .Z(n29620) );
  NAND U30388 ( .A(n29621), .B(n29620), .Z(n29660) );
  NAND U30389 ( .A(b[0]), .B(a[721]), .Z(n29622) );
  XNOR U30390 ( .A(b[1]), .B(n29622), .Z(n29624) );
  NAND U30391 ( .A(n118), .B(a[720]), .Z(n29623) );
  AND U30392 ( .A(n29624), .B(n29623), .Z(n29677) );
  XOR U30393 ( .A(a[717]), .B(n42197), .Z(n29666) );
  NANDN U30394 ( .A(n29666), .B(n42173), .Z(n29627) );
  NANDN U30395 ( .A(n29625), .B(n42172), .Z(n29626) );
  NAND U30396 ( .A(n29627), .B(n29626), .Z(n29675) );
  NAND U30397 ( .A(b[7]), .B(a[713]), .Z(n29676) );
  XNOR U30398 ( .A(n29675), .B(n29676), .Z(n29678) );
  XOR U30399 ( .A(n29677), .B(n29678), .Z(n29684) );
  NANDN U30400 ( .A(n29628), .B(n42093), .Z(n29630) );
  XOR U30401 ( .A(n42134), .B(a[719]), .Z(n29669) );
  NANDN U30402 ( .A(n29669), .B(n42095), .Z(n29629) );
  NAND U30403 ( .A(n29630), .B(n29629), .Z(n29682) );
  NANDN U30404 ( .A(n29631), .B(n42231), .Z(n29633) );
  XOR U30405 ( .A(n221), .B(a[715]), .Z(n29672) );
  NANDN U30406 ( .A(n29672), .B(n42234), .Z(n29632) );
  AND U30407 ( .A(n29633), .B(n29632), .Z(n29681) );
  XNOR U30408 ( .A(n29682), .B(n29681), .Z(n29683) );
  XNOR U30409 ( .A(n29684), .B(n29683), .Z(n29688) );
  NANDN U30410 ( .A(n29635), .B(n29634), .Z(n29639) );
  NAND U30411 ( .A(n29637), .B(n29636), .Z(n29638) );
  AND U30412 ( .A(n29639), .B(n29638), .Z(n29687) );
  XOR U30413 ( .A(n29688), .B(n29687), .Z(n29689) );
  NANDN U30414 ( .A(n29641), .B(n29640), .Z(n29645) );
  NANDN U30415 ( .A(n29643), .B(n29642), .Z(n29644) );
  NAND U30416 ( .A(n29645), .B(n29644), .Z(n29690) );
  XOR U30417 ( .A(n29689), .B(n29690), .Z(n29657) );
  OR U30418 ( .A(n29647), .B(n29646), .Z(n29651) );
  NANDN U30419 ( .A(n29649), .B(n29648), .Z(n29650) );
  NAND U30420 ( .A(n29651), .B(n29650), .Z(n29658) );
  XNOR U30421 ( .A(n29657), .B(n29658), .Z(n29659) );
  XNOR U30422 ( .A(n29660), .B(n29659), .Z(n29693) );
  XNOR U30423 ( .A(n29693), .B(sreg[1737]), .Z(n29695) );
  NAND U30424 ( .A(n29652), .B(sreg[1736]), .Z(n29656) );
  OR U30425 ( .A(n29654), .B(n29653), .Z(n29655) );
  AND U30426 ( .A(n29656), .B(n29655), .Z(n29694) );
  XOR U30427 ( .A(n29695), .B(n29694), .Z(c[1737]) );
  NANDN U30428 ( .A(n29658), .B(n29657), .Z(n29662) );
  NAND U30429 ( .A(n29660), .B(n29659), .Z(n29661) );
  NAND U30430 ( .A(n29662), .B(n29661), .Z(n29701) );
  NAND U30431 ( .A(b[0]), .B(a[722]), .Z(n29663) );
  XNOR U30432 ( .A(b[1]), .B(n29663), .Z(n29665) );
  NAND U30433 ( .A(n118), .B(a[721]), .Z(n29664) );
  AND U30434 ( .A(n29665), .B(n29664), .Z(n29718) );
  XOR U30435 ( .A(a[718]), .B(n42197), .Z(n29707) );
  NANDN U30436 ( .A(n29707), .B(n42173), .Z(n29668) );
  NANDN U30437 ( .A(n29666), .B(n42172), .Z(n29667) );
  NAND U30438 ( .A(n29668), .B(n29667), .Z(n29716) );
  NAND U30439 ( .A(b[7]), .B(a[714]), .Z(n29717) );
  XNOR U30440 ( .A(n29716), .B(n29717), .Z(n29719) );
  XOR U30441 ( .A(n29718), .B(n29719), .Z(n29725) );
  NANDN U30442 ( .A(n29669), .B(n42093), .Z(n29671) );
  XOR U30443 ( .A(n42134), .B(a[720]), .Z(n29710) );
  NANDN U30444 ( .A(n29710), .B(n42095), .Z(n29670) );
  NAND U30445 ( .A(n29671), .B(n29670), .Z(n29723) );
  NANDN U30446 ( .A(n29672), .B(n42231), .Z(n29674) );
  XOR U30447 ( .A(n221), .B(a[716]), .Z(n29713) );
  NANDN U30448 ( .A(n29713), .B(n42234), .Z(n29673) );
  AND U30449 ( .A(n29674), .B(n29673), .Z(n29722) );
  XNOR U30450 ( .A(n29723), .B(n29722), .Z(n29724) );
  XNOR U30451 ( .A(n29725), .B(n29724), .Z(n29729) );
  NANDN U30452 ( .A(n29676), .B(n29675), .Z(n29680) );
  NAND U30453 ( .A(n29678), .B(n29677), .Z(n29679) );
  AND U30454 ( .A(n29680), .B(n29679), .Z(n29728) );
  XOR U30455 ( .A(n29729), .B(n29728), .Z(n29730) );
  NANDN U30456 ( .A(n29682), .B(n29681), .Z(n29686) );
  NANDN U30457 ( .A(n29684), .B(n29683), .Z(n29685) );
  NAND U30458 ( .A(n29686), .B(n29685), .Z(n29731) );
  XOR U30459 ( .A(n29730), .B(n29731), .Z(n29698) );
  OR U30460 ( .A(n29688), .B(n29687), .Z(n29692) );
  NANDN U30461 ( .A(n29690), .B(n29689), .Z(n29691) );
  NAND U30462 ( .A(n29692), .B(n29691), .Z(n29699) );
  XNOR U30463 ( .A(n29698), .B(n29699), .Z(n29700) );
  XNOR U30464 ( .A(n29701), .B(n29700), .Z(n29734) );
  XNOR U30465 ( .A(n29734), .B(sreg[1738]), .Z(n29736) );
  NAND U30466 ( .A(n29693), .B(sreg[1737]), .Z(n29697) );
  OR U30467 ( .A(n29695), .B(n29694), .Z(n29696) );
  AND U30468 ( .A(n29697), .B(n29696), .Z(n29735) );
  XOR U30469 ( .A(n29736), .B(n29735), .Z(c[1738]) );
  NANDN U30470 ( .A(n29699), .B(n29698), .Z(n29703) );
  NAND U30471 ( .A(n29701), .B(n29700), .Z(n29702) );
  NAND U30472 ( .A(n29703), .B(n29702), .Z(n29742) );
  NAND U30473 ( .A(b[0]), .B(a[723]), .Z(n29704) );
  XNOR U30474 ( .A(b[1]), .B(n29704), .Z(n29706) );
  NAND U30475 ( .A(n118), .B(a[722]), .Z(n29705) );
  AND U30476 ( .A(n29706), .B(n29705), .Z(n29759) );
  XOR U30477 ( .A(a[719]), .B(n42197), .Z(n29748) );
  NANDN U30478 ( .A(n29748), .B(n42173), .Z(n29709) );
  NANDN U30479 ( .A(n29707), .B(n42172), .Z(n29708) );
  NAND U30480 ( .A(n29709), .B(n29708), .Z(n29757) );
  NAND U30481 ( .A(b[7]), .B(a[715]), .Z(n29758) );
  XNOR U30482 ( .A(n29757), .B(n29758), .Z(n29760) );
  XOR U30483 ( .A(n29759), .B(n29760), .Z(n29766) );
  NANDN U30484 ( .A(n29710), .B(n42093), .Z(n29712) );
  XOR U30485 ( .A(n42134), .B(a[721]), .Z(n29751) );
  NANDN U30486 ( .A(n29751), .B(n42095), .Z(n29711) );
  NAND U30487 ( .A(n29712), .B(n29711), .Z(n29764) );
  NANDN U30488 ( .A(n29713), .B(n42231), .Z(n29715) );
  XOR U30489 ( .A(n221), .B(a[717]), .Z(n29754) );
  NANDN U30490 ( .A(n29754), .B(n42234), .Z(n29714) );
  AND U30491 ( .A(n29715), .B(n29714), .Z(n29763) );
  XNOR U30492 ( .A(n29764), .B(n29763), .Z(n29765) );
  XNOR U30493 ( .A(n29766), .B(n29765), .Z(n29770) );
  NANDN U30494 ( .A(n29717), .B(n29716), .Z(n29721) );
  NAND U30495 ( .A(n29719), .B(n29718), .Z(n29720) );
  AND U30496 ( .A(n29721), .B(n29720), .Z(n29769) );
  XOR U30497 ( .A(n29770), .B(n29769), .Z(n29771) );
  NANDN U30498 ( .A(n29723), .B(n29722), .Z(n29727) );
  NANDN U30499 ( .A(n29725), .B(n29724), .Z(n29726) );
  NAND U30500 ( .A(n29727), .B(n29726), .Z(n29772) );
  XOR U30501 ( .A(n29771), .B(n29772), .Z(n29739) );
  OR U30502 ( .A(n29729), .B(n29728), .Z(n29733) );
  NANDN U30503 ( .A(n29731), .B(n29730), .Z(n29732) );
  NAND U30504 ( .A(n29733), .B(n29732), .Z(n29740) );
  XNOR U30505 ( .A(n29739), .B(n29740), .Z(n29741) );
  XNOR U30506 ( .A(n29742), .B(n29741), .Z(n29775) );
  XNOR U30507 ( .A(n29775), .B(sreg[1739]), .Z(n29777) );
  NAND U30508 ( .A(n29734), .B(sreg[1738]), .Z(n29738) );
  OR U30509 ( .A(n29736), .B(n29735), .Z(n29737) );
  AND U30510 ( .A(n29738), .B(n29737), .Z(n29776) );
  XOR U30511 ( .A(n29777), .B(n29776), .Z(c[1739]) );
  NANDN U30512 ( .A(n29740), .B(n29739), .Z(n29744) );
  NAND U30513 ( .A(n29742), .B(n29741), .Z(n29743) );
  NAND U30514 ( .A(n29744), .B(n29743), .Z(n29783) );
  NAND U30515 ( .A(b[0]), .B(a[724]), .Z(n29745) );
  XNOR U30516 ( .A(b[1]), .B(n29745), .Z(n29747) );
  NAND U30517 ( .A(n118), .B(a[723]), .Z(n29746) );
  AND U30518 ( .A(n29747), .B(n29746), .Z(n29800) );
  XOR U30519 ( .A(a[720]), .B(n42197), .Z(n29789) );
  NANDN U30520 ( .A(n29789), .B(n42173), .Z(n29750) );
  NANDN U30521 ( .A(n29748), .B(n42172), .Z(n29749) );
  NAND U30522 ( .A(n29750), .B(n29749), .Z(n29798) );
  NAND U30523 ( .A(b[7]), .B(a[716]), .Z(n29799) );
  XNOR U30524 ( .A(n29798), .B(n29799), .Z(n29801) );
  XOR U30525 ( .A(n29800), .B(n29801), .Z(n29807) );
  NANDN U30526 ( .A(n29751), .B(n42093), .Z(n29753) );
  XOR U30527 ( .A(n42134), .B(a[722]), .Z(n29792) );
  NANDN U30528 ( .A(n29792), .B(n42095), .Z(n29752) );
  NAND U30529 ( .A(n29753), .B(n29752), .Z(n29805) );
  NANDN U30530 ( .A(n29754), .B(n42231), .Z(n29756) );
  XOR U30531 ( .A(n221), .B(a[718]), .Z(n29795) );
  NANDN U30532 ( .A(n29795), .B(n42234), .Z(n29755) );
  AND U30533 ( .A(n29756), .B(n29755), .Z(n29804) );
  XNOR U30534 ( .A(n29805), .B(n29804), .Z(n29806) );
  XNOR U30535 ( .A(n29807), .B(n29806), .Z(n29811) );
  NANDN U30536 ( .A(n29758), .B(n29757), .Z(n29762) );
  NAND U30537 ( .A(n29760), .B(n29759), .Z(n29761) );
  AND U30538 ( .A(n29762), .B(n29761), .Z(n29810) );
  XOR U30539 ( .A(n29811), .B(n29810), .Z(n29812) );
  NANDN U30540 ( .A(n29764), .B(n29763), .Z(n29768) );
  NANDN U30541 ( .A(n29766), .B(n29765), .Z(n29767) );
  NAND U30542 ( .A(n29768), .B(n29767), .Z(n29813) );
  XOR U30543 ( .A(n29812), .B(n29813), .Z(n29780) );
  OR U30544 ( .A(n29770), .B(n29769), .Z(n29774) );
  NANDN U30545 ( .A(n29772), .B(n29771), .Z(n29773) );
  NAND U30546 ( .A(n29774), .B(n29773), .Z(n29781) );
  XNOR U30547 ( .A(n29780), .B(n29781), .Z(n29782) );
  XNOR U30548 ( .A(n29783), .B(n29782), .Z(n29816) );
  XNOR U30549 ( .A(n29816), .B(sreg[1740]), .Z(n29818) );
  NAND U30550 ( .A(n29775), .B(sreg[1739]), .Z(n29779) );
  OR U30551 ( .A(n29777), .B(n29776), .Z(n29778) );
  AND U30552 ( .A(n29779), .B(n29778), .Z(n29817) );
  XOR U30553 ( .A(n29818), .B(n29817), .Z(c[1740]) );
  NANDN U30554 ( .A(n29781), .B(n29780), .Z(n29785) );
  NAND U30555 ( .A(n29783), .B(n29782), .Z(n29784) );
  NAND U30556 ( .A(n29785), .B(n29784), .Z(n29824) );
  NAND U30557 ( .A(b[0]), .B(a[725]), .Z(n29786) );
  XNOR U30558 ( .A(b[1]), .B(n29786), .Z(n29788) );
  NAND U30559 ( .A(n118), .B(a[724]), .Z(n29787) );
  AND U30560 ( .A(n29788), .B(n29787), .Z(n29841) );
  XOR U30561 ( .A(a[721]), .B(n42197), .Z(n29830) );
  NANDN U30562 ( .A(n29830), .B(n42173), .Z(n29791) );
  NANDN U30563 ( .A(n29789), .B(n42172), .Z(n29790) );
  NAND U30564 ( .A(n29791), .B(n29790), .Z(n29839) );
  NAND U30565 ( .A(b[7]), .B(a[717]), .Z(n29840) );
  XNOR U30566 ( .A(n29839), .B(n29840), .Z(n29842) );
  XOR U30567 ( .A(n29841), .B(n29842), .Z(n29848) );
  NANDN U30568 ( .A(n29792), .B(n42093), .Z(n29794) );
  XOR U30569 ( .A(n42134), .B(a[723]), .Z(n29833) );
  NANDN U30570 ( .A(n29833), .B(n42095), .Z(n29793) );
  NAND U30571 ( .A(n29794), .B(n29793), .Z(n29846) );
  NANDN U30572 ( .A(n29795), .B(n42231), .Z(n29797) );
  XOR U30573 ( .A(n222), .B(a[719]), .Z(n29836) );
  NANDN U30574 ( .A(n29836), .B(n42234), .Z(n29796) );
  AND U30575 ( .A(n29797), .B(n29796), .Z(n29845) );
  XNOR U30576 ( .A(n29846), .B(n29845), .Z(n29847) );
  XNOR U30577 ( .A(n29848), .B(n29847), .Z(n29852) );
  NANDN U30578 ( .A(n29799), .B(n29798), .Z(n29803) );
  NAND U30579 ( .A(n29801), .B(n29800), .Z(n29802) );
  AND U30580 ( .A(n29803), .B(n29802), .Z(n29851) );
  XOR U30581 ( .A(n29852), .B(n29851), .Z(n29853) );
  NANDN U30582 ( .A(n29805), .B(n29804), .Z(n29809) );
  NANDN U30583 ( .A(n29807), .B(n29806), .Z(n29808) );
  NAND U30584 ( .A(n29809), .B(n29808), .Z(n29854) );
  XOR U30585 ( .A(n29853), .B(n29854), .Z(n29821) );
  OR U30586 ( .A(n29811), .B(n29810), .Z(n29815) );
  NANDN U30587 ( .A(n29813), .B(n29812), .Z(n29814) );
  NAND U30588 ( .A(n29815), .B(n29814), .Z(n29822) );
  XNOR U30589 ( .A(n29821), .B(n29822), .Z(n29823) );
  XNOR U30590 ( .A(n29824), .B(n29823), .Z(n29857) );
  XNOR U30591 ( .A(n29857), .B(sreg[1741]), .Z(n29859) );
  NAND U30592 ( .A(n29816), .B(sreg[1740]), .Z(n29820) );
  OR U30593 ( .A(n29818), .B(n29817), .Z(n29819) );
  AND U30594 ( .A(n29820), .B(n29819), .Z(n29858) );
  XOR U30595 ( .A(n29859), .B(n29858), .Z(c[1741]) );
  NANDN U30596 ( .A(n29822), .B(n29821), .Z(n29826) );
  NAND U30597 ( .A(n29824), .B(n29823), .Z(n29825) );
  NAND U30598 ( .A(n29826), .B(n29825), .Z(n29865) );
  NAND U30599 ( .A(b[0]), .B(a[726]), .Z(n29827) );
  XNOR U30600 ( .A(b[1]), .B(n29827), .Z(n29829) );
  NAND U30601 ( .A(n118), .B(a[725]), .Z(n29828) );
  AND U30602 ( .A(n29829), .B(n29828), .Z(n29882) );
  XOR U30603 ( .A(a[722]), .B(n42197), .Z(n29871) );
  NANDN U30604 ( .A(n29871), .B(n42173), .Z(n29832) );
  NANDN U30605 ( .A(n29830), .B(n42172), .Z(n29831) );
  NAND U30606 ( .A(n29832), .B(n29831), .Z(n29880) );
  NAND U30607 ( .A(b[7]), .B(a[718]), .Z(n29881) );
  XNOR U30608 ( .A(n29880), .B(n29881), .Z(n29883) );
  XOR U30609 ( .A(n29882), .B(n29883), .Z(n29889) );
  NANDN U30610 ( .A(n29833), .B(n42093), .Z(n29835) );
  XOR U30611 ( .A(n42134), .B(a[724]), .Z(n29874) );
  NANDN U30612 ( .A(n29874), .B(n42095), .Z(n29834) );
  NAND U30613 ( .A(n29835), .B(n29834), .Z(n29887) );
  NANDN U30614 ( .A(n29836), .B(n42231), .Z(n29838) );
  XOR U30615 ( .A(n222), .B(a[720]), .Z(n29877) );
  NANDN U30616 ( .A(n29877), .B(n42234), .Z(n29837) );
  AND U30617 ( .A(n29838), .B(n29837), .Z(n29886) );
  XNOR U30618 ( .A(n29887), .B(n29886), .Z(n29888) );
  XNOR U30619 ( .A(n29889), .B(n29888), .Z(n29893) );
  NANDN U30620 ( .A(n29840), .B(n29839), .Z(n29844) );
  NAND U30621 ( .A(n29842), .B(n29841), .Z(n29843) );
  AND U30622 ( .A(n29844), .B(n29843), .Z(n29892) );
  XOR U30623 ( .A(n29893), .B(n29892), .Z(n29894) );
  NANDN U30624 ( .A(n29846), .B(n29845), .Z(n29850) );
  NANDN U30625 ( .A(n29848), .B(n29847), .Z(n29849) );
  NAND U30626 ( .A(n29850), .B(n29849), .Z(n29895) );
  XOR U30627 ( .A(n29894), .B(n29895), .Z(n29862) );
  OR U30628 ( .A(n29852), .B(n29851), .Z(n29856) );
  NANDN U30629 ( .A(n29854), .B(n29853), .Z(n29855) );
  NAND U30630 ( .A(n29856), .B(n29855), .Z(n29863) );
  XNOR U30631 ( .A(n29862), .B(n29863), .Z(n29864) );
  XNOR U30632 ( .A(n29865), .B(n29864), .Z(n29898) );
  XNOR U30633 ( .A(n29898), .B(sreg[1742]), .Z(n29900) );
  NAND U30634 ( .A(n29857), .B(sreg[1741]), .Z(n29861) );
  OR U30635 ( .A(n29859), .B(n29858), .Z(n29860) );
  AND U30636 ( .A(n29861), .B(n29860), .Z(n29899) );
  XOR U30637 ( .A(n29900), .B(n29899), .Z(c[1742]) );
  NANDN U30638 ( .A(n29863), .B(n29862), .Z(n29867) );
  NAND U30639 ( .A(n29865), .B(n29864), .Z(n29866) );
  NAND U30640 ( .A(n29867), .B(n29866), .Z(n29906) );
  NAND U30641 ( .A(b[0]), .B(a[727]), .Z(n29868) );
  XNOR U30642 ( .A(b[1]), .B(n29868), .Z(n29870) );
  NAND U30643 ( .A(n118), .B(a[726]), .Z(n29869) );
  AND U30644 ( .A(n29870), .B(n29869), .Z(n29923) );
  XOR U30645 ( .A(a[723]), .B(n42197), .Z(n29912) );
  NANDN U30646 ( .A(n29912), .B(n42173), .Z(n29873) );
  NANDN U30647 ( .A(n29871), .B(n42172), .Z(n29872) );
  NAND U30648 ( .A(n29873), .B(n29872), .Z(n29921) );
  NAND U30649 ( .A(b[7]), .B(a[719]), .Z(n29922) );
  XNOR U30650 ( .A(n29921), .B(n29922), .Z(n29924) );
  XOR U30651 ( .A(n29923), .B(n29924), .Z(n29930) );
  NANDN U30652 ( .A(n29874), .B(n42093), .Z(n29876) );
  XOR U30653 ( .A(n42134), .B(a[725]), .Z(n29915) );
  NANDN U30654 ( .A(n29915), .B(n42095), .Z(n29875) );
  NAND U30655 ( .A(n29876), .B(n29875), .Z(n29928) );
  NANDN U30656 ( .A(n29877), .B(n42231), .Z(n29879) );
  XOR U30657 ( .A(n222), .B(a[721]), .Z(n29918) );
  NANDN U30658 ( .A(n29918), .B(n42234), .Z(n29878) );
  AND U30659 ( .A(n29879), .B(n29878), .Z(n29927) );
  XNOR U30660 ( .A(n29928), .B(n29927), .Z(n29929) );
  XNOR U30661 ( .A(n29930), .B(n29929), .Z(n29934) );
  NANDN U30662 ( .A(n29881), .B(n29880), .Z(n29885) );
  NAND U30663 ( .A(n29883), .B(n29882), .Z(n29884) );
  AND U30664 ( .A(n29885), .B(n29884), .Z(n29933) );
  XOR U30665 ( .A(n29934), .B(n29933), .Z(n29935) );
  NANDN U30666 ( .A(n29887), .B(n29886), .Z(n29891) );
  NANDN U30667 ( .A(n29889), .B(n29888), .Z(n29890) );
  NAND U30668 ( .A(n29891), .B(n29890), .Z(n29936) );
  XOR U30669 ( .A(n29935), .B(n29936), .Z(n29903) );
  OR U30670 ( .A(n29893), .B(n29892), .Z(n29897) );
  NANDN U30671 ( .A(n29895), .B(n29894), .Z(n29896) );
  NAND U30672 ( .A(n29897), .B(n29896), .Z(n29904) );
  XNOR U30673 ( .A(n29903), .B(n29904), .Z(n29905) );
  XNOR U30674 ( .A(n29906), .B(n29905), .Z(n29939) );
  XNOR U30675 ( .A(n29939), .B(sreg[1743]), .Z(n29941) );
  NAND U30676 ( .A(n29898), .B(sreg[1742]), .Z(n29902) );
  OR U30677 ( .A(n29900), .B(n29899), .Z(n29901) );
  AND U30678 ( .A(n29902), .B(n29901), .Z(n29940) );
  XOR U30679 ( .A(n29941), .B(n29940), .Z(c[1743]) );
  NANDN U30680 ( .A(n29904), .B(n29903), .Z(n29908) );
  NAND U30681 ( .A(n29906), .B(n29905), .Z(n29907) );
  NAND U30682 ( .A(n29908), .B(n29907), .Z(n29947) );
  NAND U30683 ( .A(b[0]), .B(a[728]), .Z(n29909) );
  XNOR U30684 ( .A(b[1]), .B(n29909), .Z(n29911) );
  NAND U30685 ( .A(n119), .B(a[727]), .Z(n29910) );
  AND U30686 ( .A(n29911), .B(n29910), .Z(n29964) );
  XOR U30687 ( .A(a[724]), .B(n42197), .Z(n29953) );
  NANDN U30688 ( .A(n29953), .B(n42173), .Z(n29914) );
  NANDN U30689 ( .A(n29912), .B(n42172), .Z(n29913) );
  NAND U30690 ( .A(n29914), .B(n29913), .Z(n29962) );
  NAND U30691 ( .A(b[7]), .B(a[720]), .Z(n29963) );
  XNOR U30692 ( .A(n29962), .B(n29963), .Z(n29965) );
  XOR U30693 ( .A(n29964), .B(n29965), .Z(n29971) );
  NANDN U30694 ( .A(n29915), .B(n42093), .Z(n29917) );
  XOR U30695 ( .A(n42134), .B(a[726]), .Z(n29956) );
  NANDN U30696 ( .A(n29956), .B(n42095), .Z(n29916) );
  NAND U30697 ( .A(n29917), .B(n29916), .Z(n29969) );
  NANDN U30698 ( .A(n29918), .B(n42231), .Z(n29920) );
  XOR U30699 ( .A(n222), .B(a[722]), .Z(n29959) );
  NANDN U30700 ( .A(n29959), .B(n42234), .Z(n29919) );
  AND U30701 ( .A(n29920), .B(n29919), .Z(n29968) );
  XNOR U30702 ( .A(n29969), .B(n29968), .Z(n29970) );
  XNOR U30703 ( .A(n29971), .B(n29970), .Z(n29975) );
  NANDN U30704 ( .A(n29922), .B(n29921), .Z(n29926) );
  NAND U30705 ( .A(n29924), .B(n29923), .Z(n29925) );
  AND U30706 ( .A(n29926), .B(n29925), .Z(n29974) );
  XOR U30707 ( .A(n29975), .B(n29974), .Z(n29976) );
  NANDN U30708 ( .A(n29928), .B(n29927), .Z(n29932) );
  NANDN U30709 ( .A(n29930), .B(n29929), .Z(n29931) );
  NAND U30710 ( .A(n29932), .B(n29931), .Z(n29977) );
  XOR U30711 ( .A(n29976), .B(n29977), .Z(n29944) );
  OR U30712 ( .A(n29934), .B(n29933), .Z(n29938) );
  NANDN U30713 ( .A(n29936), .B(n29935), .Z(n29937) );
  NAND U30714 ( .A(n29938), .B(n29937), .Z(n29945) );
  XNOR U30715 ( .A(n29944), .B(n29945), .Z(n29946) );
  XNOR U30716 ( .A(n29947), .B(n29946), .Z(n29980) );
  XNOR U30717 ( .A(n29980), .B(sreg[1744]), .Z(n29982) );
  NAND U30718 ( .A(n29939), .B(sreg[1743]), .Z(n29943) );
  OR U30719 ( .A(n29941), .B(n29940), .Z(n29942) );
  AND U30720 ( .A(n29943), .B(n29942), .Z(n29981) );
  XOR U30721 ( .A(n29982), .B(n29981), .Z(c[1744]) );
  NANDN U30722 ( .A(n29945), .B(n29944), .Z(n29949) );
  NAND U30723 ( .A(n29947), .B(n29946), .Z(n29948) );
  NAND U30724 ( .A(n29949), .B(n29948), .Z(n29988) );
  NAND U30725 ( .A(b[0]), .B(a[729]), .Z(n29950) );
  XNOR U30726 ( .A(b[1]), .B(n29950), .Z(n29952) );
  NAND U30727 ( .A(n119), .B(a[728]), .Z(n29951) );
  AND U30728 ( .A(n29952), .B(n29951), .Z(n30005) );
  XOR U30729 ( .A(a[725]), .B(n42197), .Z(n29994) );
  NANDN U30730 ( .A(n29994), .B(n42173), .Z(n29955) );
  NANDN U30731 ( .A(n29953), .B(n42172), .Z(n29954) );
  NAND U30732 ( .A(n29955), .B(n29954), .Z(n30003) );
  NAND U30733 ( .A(b[7]), .B(a[721]), .Z(n30004) );
  XNOR U30734 ( .A(n30003), .B(n30004), .Z(n30006) );
  XOR U30735 ( .A(n30005), .B(n30006), .Z(n30012) );
  NANDN U30736 ( .A(n29956), .B(n42093), .Z(n29958) );
  XOR U30737 ( .A(n42134), .B(a[727]), .Z(n29997) );
  NANDN U30738 ( .A(n29997), .B(n42095), .Z(n29957) );
  NAND U30739 ( .A(n29958), .B(n29957), .Z(n30010) );
  NANDN U30740 ( .A(n29959), .B(n42231), .Z(n29961) );
  XOR U30741 ( .A(n222), .B(a[723]), .Z(n30000) );
  NANDN U30742 ( .A(n30000), .B(n42234), .Z(n29960) );
  AND U30743 ( .A(n29961), .B(n29960), .Z(n30009) );
  XNOR U30744 ( .A(n30010), .B(n30009), .Z(n30011) );
  XNOR U30745 ( .A(n30012), .B(n30011), .Z(n30016) );
  NANDN U30746 ( .A(n29963), .B(n29962), .Z(n29967) );
  NAND U30747 ( .A(n29965), .B(n29964), .Z(n29966) );
  AND U30748 ( .A(n29967), .B(n29966), .Z(n30015) );
  XOR U30749 ( .A(n30016), .B(n30015), .Z(n30017) );
  NANDN U30750 ( .A(n29969), .B(n29968), .Z(n29973) );
  NANDN U30751 ( .A(n29971), .B(n29970), .Z(n29972) );
  NAND U30752 ( .A(n29973), .B(n29972), .Z(n30018) );
  XOR U30753 ( .A(n30017), .B(n30018), .Z(n29985) );
  OR U30754 ( .A(n29975), .B(n29974), .Z(n29979) );
  NANDN U30755 ( .A(n29977), .B(n29976), .Z(n29978) );
  NAND U30756 ( .A(n29979), .B(n29978), .Z(n29986) );
  XNOR U30757 ( .A(n29985), .B(n29986), .Z(n29987) );
  XNOR U30758 ( .A(n29988), .B(n29987), .Z(n30021) );
  XNOR U30759 ( .A(n30021), .B(sreg[1745]), .Z(n30023) );
  NAND U30760 ( .A(n29980), .B(sreg[1744]), .Z(n29984) );
  OR U30761 ( .A(n29982), .B(n29981), .Z(n29983) );
  AND U30762 ( .A(n29984), .B(n29983), .Z(n30022) );
  XOR U30763 ( .A(n30023), .B(n30022), .Z(c[1745]) );
  NANDN U30764 ( .A(n29986), .B(n29985), .Z(n29990) );
  NAND U30765 ( .A(n29988), .B(n29987), .Z(n29989) );
  NAND U30766 ( .A(n29990), .B(n29989), .Z(n30029) );
  NAND U30767 ( .A(b[0]), .B(a[730]), .Z(n29991) );
  XNOR U30768 ( .A(b[1]), .B(n29991), .Z(n29993) );
  NAND U30769 ( .A(n119), .B(a[729]), .Z(n29992) );
  AND U30770 ( .A(n29993), .B(n29992), .Z(n30046) );
  XOR U30771 ( .A(a[726]), .B(n42197), .Z(n30035) );
  NANDN U30772 ( .A(n30035), .B(n42173), .Z(n29996) );
  NANDN U30773 ( .A(n29994), .B(n42172), .Z(n29995) );
  NAND U30774 ( .A(n29996), .B(n29995), .Z(n30044) );
  NAND U30775 ( .A(b[7]), .B(a[722]), .Z(n30045) );
  XNOR U30776 ( .A(n30044), .B(n30045), .Z(n30047) );
  XOR U30777 ( .A(n30046), .B(n30047), .Z(n30053) );
  NANDN U30778 ( .A(n29997), .B(n42093), .Z(n29999) );
  XOR U30779 ( .A(n42134), .B(a[728]), .Z(n30038) );
  NANDN U30780 ( .A(n30038), .B(n42095), .Z(n29998) );
  NAND U30781 ( .A(n29999), .B(n29998), .Z(n30051) );
  NANDN U30782 ( .A(n30000), .B(n42231), .Z(n30002) );
  XOR U30783 ( .A(n222), .B(a[724]), .Z(n30041) );
  NANDN U30784 ( .A(n30041), .B(n42234), .Z(n30001) );
  AND U30785 ( .A(n30002), .B(n30001), .Z(n30050) );
  XNOR U30786 ( .A(n30051), .B(n30050), .Z(n30052) );
  XNOR U30787 ( .A(n30053), .B(n30052), .Z(n30057) );
  NANDN U30788 ( .A(n30004), .B(n30003), .Z(n30008) );
  NAND U30789 ( .A(n30006), .B(n30005), .Z(n30007) );
  AND U30790 ( .A(n30008), .B(n30007), .Z(n30056) );
  XOR U30791 ( .A(n30057), .B(n30056), .Z(n30058) );
  NANDN U30792 ( .A(n30010), .B(n30009), .Z(n30014) );
  NANDN U30793 ( .A(n30012), .B(n30011), .Z(n30013) );
  NAND U30794 ( .A(n30014), .B(n30013), .Z(n30059) );
  XOR U30795 ( .A(n30058), .B(n30059), .Z(n30026) );
  OR U30796 ( .A(n30016), .B(n30015), .Z(n30020) );
  NANDN U30797 ( .A(n30018), .B(n30017), .Z(n30019) );
  NAND U30798 ( .A(n30020), .B(n30019), .Z(n30027) );
  XNOR U30799 ( .A(n30026), .B(n30027), .Z(n30028) );
  XNOR U30800 ( .A(n30029), .B(n30028), .Z(n30062) );
  XNOR U30801 ( .A(n30062), .B(sreg[1746]), .Z(n30064) );
  NAND U30802 ( .A(n30021), .B(sreg[1745]), .Z(n30025) );
  OR U30803 ( .A(n30023), .B(n30022), .Z(n30024) );
  AND U30804 ( .A(n30025), .B(n30024), .Z(n30063) );
  XOR U30805 ( .A(n30064), .B(n30063), .Z(c[1746]) );
  NANDN U30806 ( .A(n30027), .B(n30026), .Z(n30031) );
  NAND U30807 ( .A(n30029), .B(n30028), .Z(n30030) );
  NAND U30808 ( .A(n30031), .B(n30030), .Z(n30070) );
  NAND U30809 ( .A(b[0]), .B(a[731]), .Z(n30032) );
  XNOR U30810 ( .A(b[1]), .B(n30032), .Z(n30034) );
  NAND U30811 ( .A(n119), .B(a[730]), .Z(n30033) );
  AND U30812 ( .A(n30034), .B(n30033), .Z(n30087) );
  XOR U30813 ( .A(a[727]), .B(n42197), .Z(n30076) );
  NANDN U30814 ( .A(n30076), .B(n42173), .Z(n30037) );
  NANDN U30815 ( .A(n30035), .B(n42172), .Z(n30036) );
  NAND U30816 ( .A(n30037), .B(n30036), .Z(n30085) );
  NAND U30817 ( .A(b[7]), .B(a[723]), .Z(n30086) );
  XNOR U30818 ( .A(n30085), .B(n30086), .Z(n30088) );
  XOR U30819 ( .A(n30087), .B(n30088), .Z(n30094) );
  NANDN U30820 ( .A(n30038), .B(n42093), .Z(n30040) );
  XOR U30821 ( .A(n42134), .B(a[729]), .Z(n30079) );
  NANDN U30822 ( .A(n30079), .B(n42095), .Z(n30039) );
  NAND U30823 ( .A(n30040), .B(n30039), .Z(n30092) );
  NANDN U30824 ( .A(n30041), .B(n42231), .Z(n30043) );
  XOR U30825 ( .A(n222), .B(a[725]), .Z(n30082) );
  NANDN U30826 ( .A(n30082), .B(n42234), .Z(n30042) );
  AND U30827 ( .A(n30043), .B(n30042), .Z(n30091) );
  XNOR U30828 ( .A(n30092), .B(n30091), .Z(n30093) );
  XNOR U30829 ( .A(n30094), .B(n30093), .Z(n30098) );
  NANDN U30830 ( .A(n30045), .B(n30044), .Z(n30049) );
  NAND U30831 ( .A(n30047), .B(n30046), .Z(n30048) );
  AND U30832 ( .A(n30049), .B(n30048), .Z(n30097) );
  XOR U30833 ( .A(n30098), .B(n30097), .Z(n30099) );
  NANDN U30834 ( .A(n30051), .B(n30050), .Z(n30055) );
  NANDN U30835 ( .A(n30053), .B(n30052), .Z(n30054) );
  NAND U30836 ( .A(n30055), .B(n30054), .Z(n30100) );
  XOR U30837 ( .A(n30099), .B(n30100), .Z(n30067) );
  OR U30838 ( .A(n30057), .B(n30056), .Z(n30061) );
  NANDN U30839 ( .A(n30059), .B(n30058), .Z(n30060) );
  NAND U30840 ( .A(n30061), .B(n30060), .Z(n30068) );
  XNOR U30841 ( .A(n30067), .B(n30068), .Z(n30069) );
  XNOR U30842 ( .A(n30070), .B(n30069), .Z(n30103) );
  XNOR U30843 ( .A(n30103), .B(sreg[1747]), .Z(n30105) );
  NAND U30844 ( .A(n30062), .B(sreg[1746]), .Z(n30066) );
  OR U30845 ( .A(n30064), .B(n30063), .Z(n30065) );
  AND U30846 ( .A(n30066), .B(n30065), .Z(n30104) );
  XOR U30847 ( .A(n30105), .B(n30104), .Z(c[1747]) );
  NANDN U30848 ( .A(n30068), .B(n30067), .Z(n30072) );
  NAND U30849 ( .A(n30070), .B(n30069), .Z(n30071) );
  NAND U30850 ( .A(n30072), .B(n30071), .Z(n30111) );
  NAND U30851 ( .A(b[0]), .B(a[732]), .Z(n30073) );
  XNOR U30852 ( .A(b[1]), .B(n30073), .Z(n30075) );
  NAND U30853 ( .A(n119), .B(a[731]), .Z(n30074) );
  AND U30854 ( .A(n30075), .B(n30074), .Z(n30128) );
  XOR U30855 ( .A(a[728]), .B(n42197), .Z(n30117) );
  NANDN U30856 ( .A(n30117), .B(n42173), .Z(n30078) );
  NANDN U30857 ( .A(n30076), .B(n42172), .Z(n30077) );
  NAND U30858 ( .A(n30078), .B(n30077), .Z(n30126) );
  NAND U30859 ( .A(b[7]), .B(a[724]), .Z(n30127) );
  XNOR U30860 ( .A(n30126), .B(n30127), .Z(n30129) );
  XOR U30861 ( .A(n30128), .B(n30129), .Z(n30135) );
  NANDN U30862 ( .A(n30079), .B(n42093), .Z(n30081) );
  XOR U30863 ( .A(n42134), .B(a[730]), .Z(n30120) );
  NANDN U30864 ( .A(n30120), .B(n42095), .Z(n30080) );
  NAND U30865 ( .A(n30081), .B(n30080), .Z(n30133) );
  NANDN U30866 ( .A(n30082), .B(n42231), .Z(n30084) );
  XOR U30867 ( .A(n222), .B(a[726]), .Z(n30123) );
  NANDN U30868 ( .A(n30123), .B(n42234), .Z(n30083) );
  AND U30869 ( .A(n30084), .B(n30083), .Z(n30132) );
  XNOR U30870 ( .A(n30133), .B(n30132), .Z(n30134) );
  XNOR U30871 ( .A(n30135), .B(n30134), .Z(n30139) );
  NANDN U30872 ( .A(n30086), .B(n30085), .Z(n30090) );
  NAND U30873 ( .A(n30088), .B(n30087), .Z(n30089) );
  AND U30874 ( .A(n30090), .B(n30089), .Z(n30138) );
  XOR U30875 ( .A(n30139), .B(n30138), .Z(n30140) );
  NANDN U30876 ( .A(n30092), .B(n30091), .Z(n30096) );
  NANDN U30877 ( .A(n30094), .B(n30093), .Z(n30095) );
  NAND U30878 ( .A(n30096), .B(n30095), .Z(n30141) );
  XOR U30879 ( .A(n30140), .B(n30141), .Z(n30108) );
  OR U30880 ( .A(n30098), .B(n30097), .Z(n30102) );
  NANDN U30881 ( .A(n30100), .B(n30099), .Z(n30101) );
  NAND U30882 ( .A(n30102), .B(n30101), .Z(n30109) );
  XNOR U30883 ( .A(n30108), .B(n30109), .Z(n30110) );
  XNOR U30884 ( .A(n30111), .B(n30110), .Z(n30144) );
  XNOR U30885 ( .A(n30144), .B(sreg[1748]), .Z(n30146) );
  NAND U30886 ( .A(n30103), .B(sreg[1747]), .Z(n30107) );
  OR U30887 ( .A(n30105), .B(n30104), .Z(n30106) );
  AND U30888 ( .A(n30107), .B(n30106), .Z(n30145) );
  XOR U30889 ( .A(n30146), .B(n30145), .Z(c[1748]) );
  NANDN U30890 ( .A(n30109), .B(n30108), .Z(n30113) );
  NAND U30891 ( .A(n30111), .B(n30110), .Z(n30112) );
  NAND U30892 ( .A(n30113), .B(n30112), .Z(n30152) );
  NAND U30893 ( .A(b[0]), .B(a[733]), .Z(n30114) );
  XNOR U30894 ( .A(b[1]), .B(n30114), .Z(n30116) );
  NAND U30895 ( .A(n119), .B(a[732]), .Z(n30115) );
  AND U30896 ( .A(n30116), .B(n30115), .Z(n30169) );
  XOR U30897 ( .A(a[729]), .B(n42197), .Z(n30158) );
  NANDN U30898 ( .A(n30158), .B(n42173), .Z(n30119) );
  NANDN U30899 ( .A(n30117), .B(n42172), .Z(n30118) );
  NAND U30900 ( .A(n30119), .B(n30118), .Z(n30167) );
  NAND U30901 ( .A(b[7]), .B(a[725]), .Z(n30168) );
  XNOR U30902 ( .A(n30167), .B(n30168), .Z(n30170) );
  XOR U30903 ( .A(n30169), .B(n30170), .Z(n30176) );
  NANDN U30904 ( .A(n30120), .B(n42093), .Z(n30122) );
  XOR U30905 ( .A(n42134), .B(a[731]), .Z(n30161) );
  NANDN U30906 ( .A(n30161), .B(n42095), .Z(n30121) );
  NAND U30907 ( .A(n30122), .B(n30121), .Z(n30174) );
  NANDN U30908 ( .A(n30123), .B(n42231), .Z(n30125) );
  XOR U30909 ( .A(n222), .B(a[727]), .Z(n30164) );
  NANDN U30910 ( .A(n30164), .B(n42234), .Z(n30124) );
  AND U30911 ( .A(n30125), .B(n30124), .Z(n30173) );
  XNOR U30912 ( .A(n30174), .B(n30173), .Z(n30175) );
  XNOR U30913 ( .A(n30176), .B(n30175), .Z(n30180) );
  NANDN U30914 ( .A(n30127), .B(n30126), .Z(n30131) );
  NAND U30915 ( .A(n30129), .B(n30128), .Z(n30130) );
  AND U30916 ( .A(n30131), .B(n30130), .Z(n30179) );
  XOR U30917 ( .A(n30180), .B(n30179), .Z(n30181) );
  NANDN U30918 ( .A(n30133), .B(n30132), .Z(n30137) );
  NANDN U30919 ( .A(n30135), .B(n30134), .Z(n30136) );
  NAND U30920 ( .A(n30137), .B(n30136), .Z(n30182) );
  XOR U30921 ( .A(n30181), .B(n30182), .Z(n30149) );
  OR U30922 ( .A(n30139), .B(n30138), .Z(n30143) );
  NANDN U30923 ( .A(n30141), .B(n30140), .Z(n30142) );
  NAND U30924 ( .A(n30143), .B(n30142), .Z(n30150) );
  XNOR U30925 ( .A(n30149), .B(n30150), .Z(n30151) );
  XNOR U30926 ( .A(n30152), .B(n30151), .Z(n30185) );
  XNOR U30927 ( .A(n30185), .B(sreg[1749]), .Z(n30187) );
  NAND U30928 ( .A(n30144), .B(sreg[1748]), .Z(n30148) );
  OR U30929 ( .A(n30146), .B(n30145), .Z(n30147) );
  AND U30930 ( .A(n30148), .B(n30147), .Z(n30186) );
  XOR U30931 ( .A(n30187), .B(n30186), .Z(c[1749]) );
  NANDN U30932 ( .A(n30150), .B(n30149), .Z(n30154) );
  NAND U30933 ( .A(n30152), .B(n30151), .Z(n30153) );
  NAND U30934 ( .A(n30154), .B(n30153), .Z(n30193) );
  NAND U30935 ( .A(b[0]), .B(a[734]), .Z(n30155) );
  XNOR U30936 ( .A(b[1]), .B(n30155), .Z(n30157) );
  NAND U30937 ( .A(n119), .B(a[733]), .Z(n30156) );
  AND U30938 ( .A(n30157), .B(n30156), .Z(n30210) );
  XOR U30939 ( .A(a[730]), .B(n42197), .Z(n30199) );
  NANDN U30940 ( .A(n30199), .B(n42173), .Z(n30160) );
  NANDN U30941 ( .A(n30158), .B(n42172), .Z(n30159) );
  NAND U30942 ( .A(n30160), .B(n30159), .Z(n30208) );
  NAND U30943 ( .A(b[7]), .B(a[726]), .Z(n30209) );
  XNOR U30944 ( .A(n30208), .B(n30209), .Z(n30211) );
  XOR U30945 ( .A(n30210), .B(n30211), .Z(n30217) );
  NANDN U30946 ( .A(n30161), .B(n42093), .Z(n30163) );
  XOR U30947 ( .A(n42134), .B(a[732]), .Z(n30202) );
  NANDN U30948 ( .A(n30202), .B(n42095), .Z(n30162) );
  NAND U30949 ( .A(n30163), .B(n30162), .Z(n30215) );
  NANDN U30950 ( .A(n30164), .B(n42231), .Z(n30166) );
  XOR U30951 ( .A(n222), .B(a[728]), .Z(n30205) );
  NANDN U30952 ( .A(n30205), .B(n42234), .Z(n30165) );
  AND U30953 ( .A(n30166), .B(n30165), .Z(n30214) );
  XNOR U30954 ( .A(n30215), .B(n30214), .Z(n30216) );
  XNOR U30955 ( .A(n30217), .B(n30216), .Z(n30221) );
  NANDN U30956 ( .A(n30168), .B(n30167), .Z(n30172) );
  NAND U30957 ( .A(n30170), .B(n30169), .Z(n30171) );
  AND U30958 ( .A(n30172), .B(n30171), .Z(n30220) );
  XOR U30959 ( .A(n30221), .B(n30220), .Z(n30222) );
  NANDN U30960 ( .A(n30174), .B(n30173), .Z(n30178) );
  NANDN U30961 ( .A(n30176), .B(n30175), .Z(n30177) );
  NAND U30962 ( .A(n30178), .B(n30177), .Z(n30223) );
  XOR U30963 ( .A(n30222), .B(n30223), .Z(n30190) );
  OR U30964 ( .A(n30180), .B(n30179), .Z(n30184) );
  NANDN U30965 ( .A(n30182), .B(n30181), .Z(n30183) );
  NAND U30966 ( .A(n30184), .B(n30183), .Z(n30191) );
  XNOR U30967 ( .A(n30190), .B(n30191), .Z(n30192) );
  XNOR U30968 ( .A(n30193), .B(n30192), .Z(n30226) );
  XNOR U30969 ( .A(n30226), .B(sreg[1750]), .Z(n30228) );
  NAND U30970 ( .A(n30185), .B(sreg[1749]), .Z(n30189) );
  OR U30971 ( .A(n30187), .B(n30186), .Z(n30188) );
  AND U30972 ( .A(n30189), .B(n30188), .Z(n30227) );
  XOR U30973 ( .A(n30228), .B(n30227), .Z(c[1750]) );
  NANDN U30974 ( .A(n30191), .B(n30190), .Z(n30195) );
  NAND U30975 ( .A(n30193), .B(n30192), .Z(n30194) );
  NAND U30976 ( .A(n30195), .B(n30194), .Z(n30234) );
  NAND U30977 ( .A(b[0]), .B(a[735]), .Z(n30196) );
  XNOR U30978 ( .A(b[1]), .B(n30196), .Z(n30198) );
  NAND U30979 ( .A(n120), .B(a[734]), .Z(n30197) );
  AND U30980 ( .A(n30198), .B(n30197), .Z(n30251) );
  XOR U30981 ( .A(a[731]), .B(n42197), .Z(n30240) );
  NANDN U30982 ( .A(n30240), .B(n42173), .Z(n30201) );
  NANDN U30983 ( .A(n30199), .B(n42172), .Z(n30200) );
  NAND U30984 ( .A(n30201), .B(n30200), .Z(n30249) );
  NAND U30985 ( .A(b[7]), .B(a[727]), .Z(n30250) );
  XNOR U30986 ( .A(n30249), .B(n30250), .Z(n30252) );
  XOR U30987 ( .A(n30251), .B(n30252), .Z(n30258) );
  NANDN U30988 ( .A(n30202), .B(n42093), .Z(n30204) );
  XOR U30989 ( .A(n42134), .B(a[733]), .Z(n30243) );
  NANDN U30990 ( .A(n30243), .B(n42095), .Z(n30203) );
  NAND U30991 ( .A(n30204), .B(n30203), .Z(n30256) );
  NANDN U30992 ( .A(n30205), .B(n42231), .Z(n30207) );
  XOR U30993 ( .A(n222), .B(a[729]), .Z(n30246) );
  NANDN U30994 ( .A(n30246), .B(n42234), .Z(n30206) );
  AND U30995 ( .A(n30207), .B(n30206), .Z(n30255) );
  XNOR U30996 ( .A(n30256), .B(n30255), .Z(n30257) );
  XNOR U30997 ( .A(n30258), .B(n30257), .Z(n30262) );
  NANDN U30998 ( .A(n30209), .B(n30208), .Z(n30213) );
  NAND U30999 ( .A(n30211), .B(n30210), .Z(n30212) );
  AND U31000 ( .A(n30213), .B(n30212), .Z(n30261) );
  XOR U31001 ( .A(n30262), .B(n30261), .Z(n30263) );
  NANDN U31002 ( .A(n30215), .B(n30214), .Z(n30219) );
  NANDN U31003 ( .A(n30217), .B(n30216), .Z(n30218) );
  NAND U31004 ( .A(n30219), .B(n30218), .Z(n30264) );
  XOR U31005 ( .A(n30263), .B(n30264), .Z(n30231) );
  OR U31006 ( .A(n30221), .B(n30220), .Z(n30225) );
  NANDN U31007 ( .A(n30223), .B(n30222), .Z(n30224) );
  NAND U31008 ( .A(n30225), .B(n30224), .Z(n30232) );
  XNOR U31009 ( .A(n30231), .B(n30232), .Z(n30233) );
  XNOR U31010 ( .A(n30234), .B(n30233), .Z(n30267) );
  XNOR U31011 ( .A(n30267), .B(sreg[1751]), .Z(n30269) );
  NAND U31012 ( .A(n30226), .B(sreg[1750]), .Z(n30230) );
  OR U31013 ( .A(n30228), .B(n30227), .Z(n30229) );
  AND U31014 ( .A(n30230), .B(n30229), .Z(n30268) );
  XOR U31015 ( .A(n30269), .B(n30268), .Z(c[1751]) );
  NANDN U31016 ( .A(n30232), .B(n30231), .Z(n30236) );
  NAND U31017 ( .A(n30234), .B(n30233), .Z(n30235) );
  NAND U31018 ( .A(n30236), .B(n30235), .Z(n30275) );
  NAND U31019 ( .A(b[0]), .B(a[736]), .Z(n30237) );
  XNOR U31020 ( .A(b[1]), .B(n30237), .Z(n30239) );
  NAND U31021 ( .A(n120), .B(a[735]), .Z(n30238) );
  AND U31022 ( .A(n30239), .B(n30238), .Z(n30292) );
  XOR U31023 ( .A(a[732]), .B(n42197), .Z(n30281) );
  NANDN U31024 ( .A(n30281), .B(n42173), .Z(n30242) );
  NANDN U31025 ( .A(n30240), .B(n42172), .Z(n30241) );
  NAND U31026 ( .A(n30242), .B(n30241), .Z(n30290) );
  NAND U31027 ( .A(b[7]), .B(a[728]), .Z(n30291) );
  XNOR U31028 ( .A(n30290), .B(n30291), .Z(n30293) );
  XOR U31029 ( .A(n30292), .B(n30293), .Z(n30299) );
  NANDN U31030 ( .A(n30243), .B(n42093), .Z(n30245) );
  XOR U31031 ( .A(n42134), .B(a[734]), .Z(n30284) );
  NANDN U31032 ( .A(n30284), .B(n42095), .Z(n30244) );
  NAND U31033 ( .A(n30245), .B(n30244), .Z(n30297) );
  NANDN U31034 ( .A(n30246), .B(n42231), .Z(n30248) );
  XOR U31035 ( .A(n222), .B(a[730]), .Z(n30287) );
  NANDN U31036 ( .A(n30287), .B(n42234), .Z(n30247) );
  AND U31037 ( .A(n30248), .B(n30247), .Z(n30296) );
  XNOR U31038 ( .A(n30297), .B(n30296), .Z(n30298) );
  XNOR U31039 ( .A(n30299), .B(n30298), .Z(n30303) );
  NANDN U31040 ( .A(n30250), .B(n30249), .Z(n30254) );
  NAND U31041 ( .A(n30252), .B(n30251), .Z(n30253) );
  AND U31042 ( .A(n30254), .B(n30253), .Z(n30302) );
  XOR U31043 ( .A(n30303), .B(n30302), .Z(n30304) );
  NANDN U31044 ( .A(n30256), .B(n30255), .Z(n30260) );
  NANDN U31045 ( .A(n30258), .B(n30257), .Z(n30259) );
  NAND U31046 ( .A(n30260), .B(n30259), .Z(n30305) );
  XOR U31047 ( .A(n30304), .B(n30305), .Z(n30272) );
  OR U31048 ( .A(n30262), .B(n30261), .Z(n30266) );
  NANDN U31049 ( .A(n30264), .B(n30263), .Z(n30265) );
  NAND U31050 ( .A(n30266), .B(n30265), .Z(n30273) );
  XNOR U31051 ( .A(n30272), .B(n30273), .Z(n30274) );
  XNOR U31052 ( .A(n30275), .B(n30274), .Z(n30308) );
  XNOR U31053 ( .A(n30308), .B(sreg[1752]), .Z(n30310) );
  NAND U31054 ( .A(n30267), .B(sreg[1751]), .Z(n30271) );
  OR U31055 ( .A(n30269), .B(n30268), .Z(n30270) );
  AND U31056 ( .A(n30271), .B(n30270), .Z(n30309) );
  XOR U31057 ( .A(n30310), .B(n30309), .Z(c[1752]) );
  NANDN U31058 ( .A(n30273), .B(n30272), .Z(n30277) );
  NAND U31059 ( .A(n30275), .B(n30274), .Z(n30276) );
  NAND U31060 ( .A(n30277), .B(n30276), .Z(n30316) );
  NAND U31061 ( .A(b[0]), .B(a[737]), .Z(n30278) );
  XNOR U31062 ( .A(b[1]), .B(n30278), .Z(n30280) );
  NAND U31063 ( .A(n120), .B(a[736]), .Z(n30279) );
  AND U31064 ( .A(n30280), .B(n30279), .Z(n30333) );
  XOR U31065 ( .A(a[733]), .B(n42197), .Z(n30322) );
  NANDN U31066 ( .A(n30322), .B(n42173), .Z(n30283) );
  NANDN U31067 ( .A(n30281), .B(n42172), .Z(n30282) );
  NAND U31068 ( .A(n30283), .B(n30282), .Z(n30331) );
  NAND U31069 ( .A(b[7]), .B(a[729]), .Z(n30332) );
  XNOR U31070 ( .A(n30331), .B(n30332), .Z(n30334) );
  XOR U31071 ( .A(n30333), .B(n30334), .Z(n30340) );
  NANDN U31072 ( .A(n30284), .B(n42093), .Z(n30286) );
  XOR U31073 ( .A(n42134), .B(a[735]), .Z(n30325) );
  NANDN U31074 ( .A(n30325), .B(n42095), .Z(n30285) );
  NAND U31075 ( .A(n30286), .B(n30285), .Z(n30338) );
  NANDN U31076 ( .A(n30287), .B(n42231), .Z(n30289) );
  XOR U31077 ( .A(n223), .B(a[731]), .Z(n30328) );
  NANDN U31078 ( .A(n30328), .B(n42234), .Z(n30288) );
  AND U31079 ( .A(n30289), .B(n30288), .Z(n30337) );
  XNOR U31080 ( .A(n30338), .B(n30337), .Z(n30339) );
  XNOR U31081 ( .A(n30340), .B(n30339), .Z(n30344) );
  NANDN U31082 ( .A(n30291), .B(n30290), .Z(n30295) );
  NAND U31083 ( .A(n30293), .B(n30292), .Z(n30294) );
  AND U31084 ( .A(n30295), .B(n30294), .Z(n30343) );
  XOR U31085 ( .A(n30344), .B(n30343), .Z(n30345) );
  NANDN U31086 ( .A(n30297), .B(n30296), .Z(n30301) );
  NANDN U31087 ( .A(n30299), .B(n30298), .Z(n30300) );
  NAND U31088 ( .A(n30301), .B(n30300), .Z(n30346) );
  XOR U31089 ( .A(n30345), .B(n30346), .Z(n30313) );
  OR U31090 ( .A(n30303), .B(n30302), .Z(n30307) );
  NANDN U31091 ( .A(n30305), .B(n30304), .Z(n30306) );
  NAND U31092 ( .A(n30307), .B(n30306), .Z(n30314) );
  XNOR U31093 ( .A(n30313), .B(n30314), .Z(n30315) );
  XNOR U31094 ( .A(n30316), .B(n30315), .Z(n30349) );
  XNOR U31095 ( .A(n30349), .B(sreg[1753]), .Z(n30351) );
  NAND U31096 ( .A(n30308), .B(sreg[1752]), .Z(n30312) );
  OR U31097 ( .A(n30310), .B(n30309), .Z(n30311) );
  AND U31098 ( .A(n30312), .B(n30311), .Z(n30350) );
  XOR U31099 ( .A(n30351), .B(n30350), .Z(c[1753]) );
  NANDN U31100 ( .A(n30314), .B(n30313), .Z(n30318) );
  NAND U31101 ( .A(n30316), .B(n30315), .Z(n30317) );
  NAND U31102 ( .A(n30318), .B(n30317), .Z(n30357) );
  NAND U31103 ( .A(b[0]), .B(a[738]), .Z(n30319) );
  XNOR U31104 ( .A(b[1]), .B(n30319), .Z(n30321) );
  NAND U31105 ( .A(n120), .B(a[737]), .Z(n30320) );
  AND U31106 ( .A(n30321), .B(n30320), .Z(n30374) );
  XOR U31107 ( .A(a[734]), .B(n42197), .Z(n30363) );
  NANDN U31108 ( .A(n30363), .B(n42173), .Z(n30324) );
  NANDN U31109 ( .A(n30322), .B(n42172), .Z(n30323) );
  NAND U31110 ( .A(n30324), .B(n30323), .Z(n30372) );
  NAND U31111 ( .A(b[7]), .B(a[730]), .Z(n30373) );
  XNOR U31112 ( .A(n30372), .B(n30373), .Z(n30375) );
  XOR U31113 ( .A(n30374), .B(n30375), .Z(n30381) );
  NANDN U31114 ( .A(n30325), .B(n42093), .Z(n30327) );
  XOR U31115 ( .A(n42134), .B(a[736]), .Z(n30366) );
  NANDN U31116 ( .A(n30366), .B(n42095), .Z(n30326) );
  NAND U31117 ( .A(n30327), .B(n30326), .Z(n30379) );
  NANDN U31118 ( .A(n30328), .B(n42231), .Z(n30330) );
  XOR U31119 ( .A(n223), .B(a[732]), .Z(n30369) );
  NANDN U31120 ( .A(n30369), .B(n42234), .Z(n30329) );
  AND U31121 ( .A(n30330), .B(n30329), .Z(n30378) );
  XNOR U31122 ( .A(n30379), .B(n30378), .Z(n30380) );
  XNOR U31123 ( .A(n30381), .B(n30380), .Z(n30385) );
  NANDN U31124 ( .A(n30332), .B(n30331), .Z(n30336) );
  NAND U31125 ( .A(n30334), .B(n30333), .Z(n30335) );
  AND U31126 ( .A(n30336), .B(n30335), .Z(n30384) );
  XOR U31127 ( .A(n30385), .B(n30384), .Z(n30386) );
  NANDN U31128 ( .A(n30338), .B(n30337), .Z(n30342) );
  NANDN U31129 ( .A(n30340), .B(n30339), .Z(n30341) );
  NAND U31130 ( .A(n30342), .B(n30341), .Z(n30387) );
  XOR U31131 ( .A(n30386), .B(n30387), .Z(n30354) );
  OR U31132 ( .A(n30344), .B(n30343), .Z(n30348) );
  NANDN U31133 ( .A(n30346), .B(n30345), .Z(n30347) );
  NAND U31134 ( .A(n30348), .B(n30347), .Z(n30355) );
  XNOR U31135 ( .A(n30354), .B(n30355), .Z(n30356) );
  XNOR U31136 ( .A(n30357), .B(n30356), .Z(n30390) );
  XNOR U31137 ( .A(n30390), .B(sreg[1754]), .Z(n30392) );
  NAND U31138 ( .A(n30349), .B(sreg[1753]), .Z(n30353) );
  OR U31139 ( .A(n30351), .B(n30350), .Z(n30352) );
  AND U31140 ( .A(n30353), .B(n30352), .Z(n30391) );
  XOR U31141 ( .A(n30392), .B(n30391), .Z(c[1754]) );
  NANDN U31142 ( .A(n30355), .B(n30354), .Z(n30359) );
  NAND U31143 ( .A(n30357), .B(n30356), .Z(n30358) );
  NAND U31144 ( .A(n30359), .B(n30358), .Z(n30398) );
  NAND U31145 ( .A(b[0]), .B(a[739]), .Z(n30360) );
  XNOR U31146 ( .A(b[1]), .B(n30360), .Z(n30362) );
  NAND U31147 ( .A(n120), .B(a[738]), .Z(n30361) );
  AND U31148 ( .A(n30362), .B(n30361), .Z(n30415) );
  XOR U31149 ( .A(a[735]), .B(n42197), .Z(n30404) );
  NANDN U31150 ( .A(n30404), .B(n42173), .Z(n30365) );
  NANDN U31151 ( .A(n30363), .B(n42172), .Z(n30364) );
  NAND U31152 ( .A(n30365), .B(n30364), .Z(n30413) );
  NAND U31153 ( .A(b[7]), .B(a[731]), .Z(n30414) );
  XNOR U31154 ( .A(n30413), .B(n30414), .Z(n30416) );
  XOR U31155 ( .A(n30415), .B(n30416), .Z(n30422) );
  NANDN U31156 ( .A(n30366), .B(n42093), .Z(n30368) );
  XOR U31157 ( .A(n42134), .B(a[737]), .Z(n30407) );
  NANDN U31158 ( .A(n30407), .B(n42095), .Z(n30367) );
  NAND U31159 ( .A(n30368), .B(n30367), .Z(n30420) );
  NANDN U31160 ( .A(n30369), .B(n42231), .Z(n30371) );
  XOR U31161 ( .A(n223), .B(a[733]), .Z(n30410) );
  NANDN U31162 ( .A(n30410), .B(n42234), .Z(n30370) );
  AND U31163 ( .A(n30371), .B(n30370), .Z(n30419) );
  XNOR U31164 ( .A(n30420), .B(n30419), .Z(n30421) );
  XNOR U31165 ( .A(n30422), .B(n30421), .Z(n30426) );
  NANDN U31166 ( .A(n30373), .B(n30372), .Z(n30377) );
  NAND U31167 ( .A(n30375), .B(n30374), .Z(n30376) );
  AND U31168 ( .A(n30377), .B(n30376), .Z(n30425) );
  XOR U31169 ( .A(n30426), .B(n30425), .Z(n30427) );
  NANDN U31170 ( .A(n30379), .B(n30378), .Z(n30383) );
  NANDN U31171 ( .A(n30381), .B(n30380), .Z(n30382) );
  NAND U31172 ( .A(n30383), .B(n30382), .Z(n30428) );
  XOR U31173 ( .A(n30427), .B(n30428), .Z(n30395) );
  OR U31174 ( .A(n30385), .B(n30384), .Z(n30389) );
  NANDN U31175 ( .A(n30387), .B(n30386), .Z(n30388) );
  NAND U31176 ( .A(n30389), .B(n30388), .Z(n30396) );
  XNOR U31177 ( .A(n30395), .B(n30396), .Z(n30397) );
  XNOR U31178 ( .A(n30398), .B(n30397), .Z(n30431) );
  XNOR U31179 ( .A(n30431), .B(sreg[1755]), .Z(n30433) );
  NAND U31180 ( .A(n30390), .B(sreg[1754]), .Z(n30394) );
  OR U31181 ( .A(n30392), .B(n30391), .Z(n30393) );
  AND U31182 ( .A(n30394), .B(n30393), .Z(n30432) );
  XOR U31183 ( .A(n30433), .B(n30432), .Z(c[1755]) );
  NANDN U31184 ( .A(n30396), .B(n30395), .Z(n30400) );
  NAND U31185 ( .A(n30398), .B(n30397), .Z(n30399) );
  NAND U31186 ( .A(n30400), .B(n30399), .Z(n30439) );
  NAND U31187 ( .A(b[0]), .B(a[740]), .Z(n30401) );
  XNOR U31188 ( .A(b[1]), .B(n30401), .Z(n30403) );
  NAND U31189 ( .A(n120), .B(a[739]), .Z(n30402) );
  AND U31190 ( .A(n30403), .B(n30402), .Z(n30456) );
  XOR U31191 ( .A(a[736]), .B(n42197), .Z(n30445) );
  NANDN U31192 ( .A(n30445), .B(n42173), .Z(n30406) );
  NANDN U31193 ( .A(n30404), .B(n42172), .Z(n30405) );
  NAND U31194 ( .A(n30406), .B(n30405), .Z(n30454) );
  NAND U31195 ( .A(b[7]), .B(a[732]), .Z(n30455) );
  XNOR U31196 ( .A(n30454), .B(n30455), .Z(n30457) );
  XOR U31197 ( .A(n30456), .B(n30457), .Z(n30463) );
  NANDN U31198 ( .A(n30407), .B(n42093), .Z(n30409) );
  XOR U31199 ( .A(n42134), .B(a[738]), .Z(n30448) );
  NANDN U31200 ( .A(n30448), .B(n42095), .Z(n30408) );
  NAND U31201 ( .A(n30409), .B(n30408), .Z(n30461) );
  NANDN U31202 ( .A(n30410), .B(n42231), .Z(n30412) );
  XOR U31203 ( .A(n223), .B(a[734]), .Z(n30451) );
  NANDN U31204 ( .A(n30451), .B(n42234), .Z(n30411) );
  AND U31205 ( .A(n30412), .B(n30411), .Z(n30460) );
  XNOR U31206 ( .A(n30461), .B(n30460), .Z(n30462) );
  XNOR U31207 ( .A(n30463), .B(n30462), .Z(n30467) );
  NANDN U31208 ( .A(n30414), .B(n30413), .Z(n30418) );
  NAND U31209 ( .A(n30416), .B(n30415), .Z(n30417) );
  AND U31210 ( .A(n30418), .B(n30417), .Z(n30466) );
  XOR U31211 ( .A(n30467), .B(n30466), .Z(n30468) );
  NANDN U31212 ( .A(n30420), .B(n30419), .Z(n30424) );
  NANDN U31213 ( .A(n30422), .B(n30421), .Z(n30423) );
  NAND U31214 ( .A(n30424), .B(n30423), .Z(n30469) );
  XOR U31215 ( .A(n30468), .B(n30469), .Z(n30436) );
  OR U31216 ( .A(n30426), .B(n30425), .Z(n30430) );
  NANDN U31217 ( .A(n30428), .B(n30427), .Z(n30429) );
  NAND U31218 ( .A(n30430), .B(n30429), .Z(n30437) );
  XNOR U31219 ( .A(n30436), .B(n30437), .Z(n30438) );
  XNOR U31220 ( .A(n30439), .B(n30438), .Z(n30472) );
  XNOR U31221 ( .A(n30472), .B(sreg[1756]), .Z(n30474) );
  NAND U31222 ( .A(n30431), .B(sreg[1755]), .Z(n30435) );
  OR U31223 ( .A(n30433), .B(n30432), .Z(n30434) );
  AND U31224 ( .A(n30435), .B(n30434), .Z(n30473) );
  XOR U31225 ( .A(n30474), .B(n30473), .Z(c[1756]) );
  NANDN U31226 ( .A(n30437), .B(n30436), .Z(n30441) );
  NAND U31227 ( .A(n30439), .B(n30438), .Z(n30440) );
  NAND U31228 ( .A(n30441), .B(n30440), .Z(n30480) );
  NAND U31229 ( .A(b[0]), .B(a[741]), .Z(n30442) );
  XNOR U31230 ( .A(b[1]), .B(n30442), .Z(n30444) );
  NAND U31231 ( .A(n120), .B(a[740]), .Z(n30443) );
  AND U31232 ( .A(n30444), .B(n30443), .Z(n30497) );
  XOR U31233 ( .A(a[737]), .B(n42197), .Z(n30486) );
  NANDN U31234 ( .A(n30486), .B(n42173), .Z(n30447) );
  NANDN U31235 ( .A(n30445), .B(n42172), .Z(n30446) );
  NAND U31236 ( .A(n30447), .B(n30446), .Z(n30495) );
  NAND U31237 ( .A(b[7]), .B(a[733]), .Z(n30496) );
  XNOR U31238 ( .A(n30495), .B(n30496), .Z(n30498) );
  XOR U31239 ( .A(n30497), .B(n30498), .Z(n30504) );
  NANDN U31240 ( .A(n30448), .B(n42093), .Z(n30450) );
  XOR U31241 ( .A(n42134), .B(a[739]), .Z(n30489) );
  NANDN U31242 ( .A(n30489), .B(n42095), .Z(n30449) );
  NAND U31243 ( .A(n30450), .B(n30449), .Z(n30502) );
  NANDN U31244 ( .A(n30451), .B(n42231), .Z(n30453) );
  XOR U31245 ( .A(n223), .B(a[735]), .Z(n30492) );
  NANDN U31246 ( .A(n30492), .B(n42234), .Z(n30452) );
  AND U31247 ( .A(n30453), .B(n30452), .Z(n30501) );
  XNOR U31248 ( .A(n30502), .B(n30501), .Z(n30503) );
  XNOR U31249 ( .A(n30504), .B(n30503), .Z(n30508) );
  NANDN U31250 ( .A(n30455), .B(n30454), .Z(n30459) );
  NAND U31251 ( .A(n30457), .B(n30456), .Z(n30458) );
  AND U31252 ( .A(n30459), .B(n30458), .Z(n30507) );
  XOR U31253 ( .A(n30508), .B(n30507), .Z(n30509) );
  NANDN U31254 ( .A(n30461), .B(n30460), .Z(n30465) );
  NANDN U31255 ( .A(n30463), .B(n30462), .Z(n30464) );
  NAND U31256 ( .A(n30465), .B(n30464), .Z(n30510) );
  XOR U31257 ( .A(n30509), .B(n30510), .Z(n30477) );
  OR U31258 ( .A(n30467), .B(n30466), .Z(n30471) );
  NANDN U31259 ( .A(n30469), .B(n30468), .Z(n30470) );
  NAND U31260 ( .A(n30471), .B(n30470), .Z(n30478) );
  XNOR U31261 ( .A(n30477), .B(n30478), .Z(n30479) );
  XNOR U31262 ( .A(n30480), .B(n30479), .Z(n30513) );
  XNOR U31263 ( .A(n30513), .B(sreg[1757]), .Z(n30515) );
  NAND U31264 ( .A(n30472), .B(sreg[1756]), .Z(n30476) );
  OR U31265 ( .A(n30474), .B(n30473), .Z(n30475) );
  AND U31266 ( .A(n30476), .B(n30475), .Z(n30514) );
  XOR U31267 ( .A(n30515), .B(n30514), .Z(c[1757]) );
  NANDN U31268 ( .A(n30478), .B(n30477), .Z(n30482) );
  NAND U31269 ( .A(n30480), .B(n30479), .Z(n30481) );
  NAND U31270 ( .A(n30482), .B(n30481), .Z(n30521) );
  NAND U31271 ( .A(b[0]), .B(a[742]), .Z(n30483) );
  XNOR U31272 ( .A(b[1]), .B(n30483), .Z(n30485) );
  NAND U31273 ( .A(n121), .B(a[741]), .Z(n30484) );
  AND U31274 ( .A(n30485), .B(n30484), .Z(n30538) );
  XOR U31275 ( .A(a[738]), .B(n42197), .Z(n30527) );
  NANDN U31276 ( .A(n30527), .B(n42173), .Z(n30488) );
  NANDN U31277 ( .A(n30486), .B(n42172), .Z(n30487) );
  NAND U31278 ( .A(n30488), .B(n30487), .Z(n30536) );
  NAND U31279 ( .A(b[7]), .B(a[734]), .Z(n30537) );
  XNOR U31280 ( .A(n30536), .B(n30537), .Z(n30539) );
  XOR U31281 ( .A(n30538), .B(n30539), .Z(n30545) );
  NANDN U31282 ( .A(n30489), .B(n42093), .Z(n30491) );
  XOR U31283 ( .A(n42134), .B(a[740]), .Z(n30530) );
  NANDN U31284 ( .A(n30530), .B(n42095), .Z(n30490) );
  NAND U31285 ( .A(n30491), .B(n30490), .Z(n30543) );
  NANDN U31286 ( .A(n30492), .B(n42231), .Z(n30494) );
  XOR U31287 ( .A(n223), .B(a[736]), .Z(n30533) );
  NANDN U31288 ( .A(n30533), .B(n42234), .Z(n30493) );
  AND U31289 ( .A(n30494), .B(n30493), .Z(n30542) );
  XNOR U31290 ( .A(n30543), .B(n30542), .Z(n30544) );
  XNOR U31291 ( .A(n30545), .B(n30544), .Z(n30549) );
  NANDN U31292 ( .A(n30496), .B(n30495), .Z(n30500) );
  NAND U31293 ( .A(n30498), .B(n30497), .Z(n30499) );
  AND U31294 ( .A(n30500), .B(n30499), .Z(n30548) );
  XOR U31295 ( .A(n30549), .B(n30548), .Z(n30550) );
  NANDN U31296 ( .A(n30502), .B(n30501), .Z(n30506) );
  NANDN U31297 ( .A(n30504), .B(n30503), .Z(n30505) );
  NAND U31298 ( .A(n30506), .B(n30505), .Z(n30551) );
  XOR U31299 ( .A(n30550), .B(n30551), .Z(n30518) );
  OR U31300 ( .A(n30508), .B(n30507), .Z(n30512) );
  NANDN U31301 ( .A(n30510), .B(n30509), .Z(n30511) );
  NAND U31302 ( .A(n30512), .B(n30511), .Z(n30519) );
  XNOR U31303 ( .A(n30518), .B(n30519), .Z(n30520) );
  XNOR U31304 ( .A(n30521), .B(n30520), .Z(n30554) );
  XNOR U31305 ( .A(n30554), .B(sreg[1758]), .Z(n30556) );
  NAND U31306 ( .A(n30513), .B(sreg[1757]), .Z(n30517) );
  OR U31307 ( .A(n30515), .B(n30514), .Z(n30516) );
  AND U31308 ( .A(n30517), .B(n30516), .Z(n30555) );
  XOR U31309 ( .A(n30556), .B(n30555), .Z(c[1758]) );
  NANDN U31310 ( .A(n30519), .B(n30518), .Z(n30523) );
  NAND U31311 ( .A(n30521), .B(n30520), .Z(n30522) );
  NAND U31312 ( .A(n30523), .B(n30522), .Z(n30562) );
  NAND U31313 ( .A(b[0]), .B(a[743]), .Z(n30524) );
  XNOR U31314 ( .A(b[1]), .B(n30524), .Z(n30526) );
  NAND U31315 ( .A(n121), .B(a[742]), .Z(n30525) );
  AND U31316 ( .A(n30526), .B(n30525), .Z(n30579) );
  XOR U31317 ( .A(a[739]), .B(n42197), .Z(n30568) );
  NANDN U31318 ( .A(n30568), .B(n42173), .Z(n30529) );
  NANDN U31319 ( .A(n30527), .B(n42172), .Z(n30528) );
  NAND U31320 ( .A(n30529), .B(n30528), .Z(n30577) );
  NAND U31321 ( .A(b[7]), .B(a[735]), .Z(n30578) );
  XNOR U31322 ( .A(n30577), .B(n30578), .Z(n30580) );
  XOR U31323 ( .A(n30579), .B(n30580), .Z(n30586) );
  NANDN U31324 ( .A(n30530), .B(n42093), .Z(n30532) );
  XOR U31325 ( .A(n42134), .B(a[741]), .Z(n30571) );
  NANDN U31326 ( .A(n30571), .B(n42095), .Z(n30531) );
  NAND U31327 ( .A(n30532), .B(n30531), .Z(n30584) );
  NANDN U31328 ( .A(n30533), .B(n42231), .Z(n30535) );
  XOR U31329 ( .A(n223), .B(a[737]), .Z(n30574) );
  NANDN U31330 ( .A(n30574), .B(n42234), .Z(n30534) );
  AND U31331 ( .A(n30535), .B(n30534), .Z(n30583) );
  XNOR U31332 ( .A(n30584), .B(n30583), .Z(n30585) );
  XNOR U31333 ( .A(n30586), .B(n30585), .Z(n30590) );
  NANDN U31334 ( .A(n30537), .B(n30536), .Z(n30541) );
  NAND U31335 ( .A(n30539), .B(n30538), .Z(n30540) );
  AND U31336 ( .A(n30541), .B(n30540), .Z(n30589) );
  XOR U31337 ( .A(n30590), .B(n30589), .Z(n30591) );
  NANDN U31338 ( .A(n30543), .B(n30542), .Z(n30547) );
  NANDN U31339 ( .A(n30545), .B(n30544), .Z(n30546) );
  NAND U31340 ( .A(n30547), .B(n30546), .Z(n30592) );
  XOR U31341 ( .A(n30591), .B(n30592), .Z(n30559) );
  OR U31342 ( .A(n30549), .B(n30548), .Z(n30553) );
  NANDN U31343 ( .A(n30551), .B(n30550), .Z(n30552) );
  NAND U31344 ( .A(n30553), .B(n30552), .Z(n30560) );
  XNOR U31345 ( .A(n30559), .B(n30560), .Z(n30561) );
  XNOR U31346 ( .A(n30562), .B(n30561), .Z(n30595) );
  XNOR U31347 ( .A(n30595), .B(sreg[1759]), .Z(n30597) );
  NAND U31348 ( .A(n30554), .B(sreg[1758]), .Z(n30558) );
  OR U31349 ( .A(n30556), .B(n30555), .Z(n30557) );
  AND U31350 ( .A(n30558), .B(n30557), .Z(n30596) );
  XOR U31351 ( .A(n30597), .B(n30596), .Z(c[1759]) );
  NANDN U31352 ( .A(n30560), .B(n30559), .Z(n30564) );
  NAND U31353 ( .A(n30562), .B(n30561), .Z(n30563) );
  NAND U31354 ( .A(n30564), .B(n30563), .Z(n30603) );
  NAND U31355 ( .A(b[0]), .B(a[744]), .Z(n30565) );
  XNOR U31356 ( .A(b[1]), .B(n30565), .Z(n30567) );
  NAND U31357 ( .A(n121), .B(a[743]), .Z(n30566) );
  AND U31358 ( .A(n30567), .B(n30566), .Z(n30620) );
  XOR U31359 ( .A(a[740]), .B(n42197), .Z(n30609) );
  NANDN U31360 ( .A(n30609), .B(n42173), .Z(n30570) );
  NANDN U31361 ( .A(n30568), .B(n42172), .Z(n30569) );
  NAND U31362 ( .A(n30570), .B(n30569), .Z(n30618) );
  NAND U31363 ( .A(b[7]), .B(a[736]), .Z(n30619) );
  XNOR U31364 ( .A(n30618), .B(n30619), .Z(n30621) );
  XOR U31365 ( .A(n30620), .B(n30621), .Z(n30627) );
  NANDN U31366 ( .A(n30571), .B(n42093), .Z(n30573) );
  XOR U31367 ( .A(n42134), .B(a[742]), .Z(n30612) );
  NANDN U31368 ( .A(n30612), .B(n42095), .Z(n30572) );
  NAND U31369 ( .A(n30573), .B(n30572), .Z(n30625) );
  NANDN U31370 ( .A(n30574), .B(n42231), .Z(n30576) );
  XOR U31371 ( .A(n223), .B(a[738]), .Z(n30615) );
  NANDN U31372 ( .A(n30615), .B(n42234), .Z(n30575) );
  AND U31373 ( .A(n30576), .B(n30575), .Z(n30624) );
  XNOR U31374 ( .A(n30625), .B(n30624), .Z(n30626) );
  XNOR U31375 ( .A(n30627), .B(n30626), .Z(n30631) );
  NANDN U31376 ( .A(n30578), .B(n30577), .Z(n30582) );
  NAND U31377 ( .A(n30580), .B(n30579), .Z(n30581) );
  AND U31378 ( .A(n30582), .B(n30581), .Z(n30630) );
  XOR U31379 ( .A(n30631), .B(n30630), .Z(n30632) );
  NANDN U31380 ( .A(n30584), .B(n30583), .Z(n30588) );
  NANDN U31381 ( .A(n30586), .B(n30585), .Z(n30587) );
  NAND U31382 ( .A(n30588), .B(n30587), .Z(n30633) );
  XOR U31383 ( .A(n30632), .B(n30633), .Z(n30600) );
  OR U31384 ( .A(n30590), .B(n30589), .Z(n30594) );
  NANDN U31385 ( .A(n30592), .B(n30591), .Z(n30593) );
  NAND U31386 ( .A(n30594), .B(n30593), .Z(n30601) );
  XNOR U31387 ( .A(n30600), .B(n30601), .Z(n30602) );
  XNOR U31388 ( .A(n30603), .B(n30602), .Z(n30636) );
  XNOR U31389 ( .A(n30636), .B(sreg[1760]), .Z(n30638) );
  NAND U31390 ( .A(n30595), .B(sreg[1759]), .Z(n30599) );
  OR U31391 ( .A(n30597), .B(n30596), .Z(n30598) );
  AND U31392 ( .A(n30599), .B(n30598), .Z(n30637) );
  XOR U31393 ( .A(n30638), .B(n30637), .Z(c[1760]) );
  NANDN U31394 ( .A(n30601), .B(n30600), .Z(n30605) );
  NAND U31395 ( .A(n30603), .B(n30602), .Z(n30604) );
  NAND U31396 ( .A(n30605), .B(n30604), .Z(n30644) );
  NAND U31397 ( .A(b[0]), .B(a[745]), .Z(n30606) );
  XNOR U31398 ( .A(b[1]), .B(n30606), .Z(n30608) );
  NAND U31399 ( .A(n121), .B(a[744]), .Z(n30607) );
  AND U31400 ( .A(n30608), .B(n30607), .Z(n30661) );
  XOR U31401 ( .A(a[741]), .B(n42197), .Z(n30650) );
  NANDN U31402 ( .A(n30650), .B(n42173), .Z(n30611) );
  NANDN U31403 ( .A(n30609), .B(n42172), .Z(n30610) );
  NAND U31404 ( .A(n30611), .B(n30610), .Z(n30659) );
  NAND U31405 ( .A(b[7]), .B(a[737]), .Z(n30660) );
  XNOR U31406 ( .A(n30659), .B(n30660), .Z(n30662) );
  XOR U31407 ( .A(n30661), .B(n30662), .Z(n30668) );
  NANDN U31408 ( .A(n30612), .B(n42093), .Z(n30614) );
  XOR U31409 ( .A(n42134), .B(a[743]), .Z(n30653) );
  NANDN U31410 ( .A(n30653), .B(n42095), .Z(n30613) );
  NAND U31411 ( .A(n30614), .B(n30613), .Z(n30666) );
  NANDN U31412 ( .A(n30615), .B(n42231), .Z(n30617) );
  XOR U31413 ( .A(n223), .B(a[739]), .Z(n30656) );
  NANDN U31414 ( .A(n30656), .B(n42234), .Z(n30616) );
  AND U31415 ( .A(n30617), .B(n30616), .Z(n30665) );
  XNOR U31416 ( .A(n30666), .B(n30665), .Z(n30667) );
  XNOR U31417 ( .A(n30668), .B(n30667), .Z(n30672) );
  NANDN U31418 ( .A(n30619), .B(n30618), .Z(n30623) );
  NAND U31419 ( .A(n30621), .B(n30620), .Z(n30622) );
  AND U31420 ( .A(n30623), .B(n30622), .Z(n30671) );
  XOR U31421 ( .A(n30672), .B(n30671), .Z(n30673) );
  NANDN U31422 ( .A(n30625), .B(n30624), .Z(n30629) );
  NANDN U31423 ( .A(n30627), .B(n30626), .Z(n30628) );
  NAND U31424 ( .A(n30629), .B(n30628), .Z(n30674) );
  XOR U31425 ( .A(n30673), .B(n30674), .Z(n30641) );
  OR U31426 ( .A(n30631), .B(n30630), .Z(n30635) );
  NANDN U31427 ( .A(n30633), .B(n30632), .Z(n30634) );
  NAND U31428 ( .A(n30635), .B(n30634), .Z(n30642) );
  XNOR U31429 ( .A(n30641), .B(n30642), .Z(n30643) );
  XNOR U31430 ( .A(n30644), .B(n30643), .Z(n30677) );
  XNOR U31431 ( .A(n30677), .B(sreg[1761]), .Z(n30679) );
  NAND U31432 ( .A(n30636), .B(sreg[1760]), .Z(n30640) );
  OR U31433 ( .A(n30638), .B(n30637), .Z(n30639) );
  AND U31434 ( .A(n30640), .B(n30639), .Z(n30678) );
  XOR U31435 ( .A(n30679), .B(n30678), .Z(c[1761]) );
  NANDN U31436 ( .A(n30642), .B(n30641), .Z(n30646) );
  NAND U31437 ( .A(n30644), .B(n30643), .Z(n30645) );
  NAND U31438 ( .A(n30646), .B(n30645), .Z(n30685) );
  NAND U31439 ( .A(b[0]), .B(a[746]), .Z(n30647) );
  XNOR U31440 ( .A(b[1]), .B(n30647), .Z(n30649) );
  NAND U31441 ( .A(n121), .B(a[745]), .Z(n30648) );
  AND U31442 ( .A(n30649), .B(n30648), .Z(n30702) );
  XOR U31443 ( .A(a[742]), .B(n42197), .Z(n30691) );
  NANDN U31444 ( .A(n30691), .B(n42173), .Z(n30652) );
  NANDN U31445 ( .A(n30650), .B(n42172), .Z(n30651) );
  NAND U31446 ( .A(n30652), .B(n30651), .Z(n30700) );
  NAND U31447 ( .A(b[7]), .B(a[738]), .Z(n30701) );
  XNOR U31448 ( .A(n30700), .B(n30701), .Z(n30703) );
  XOR U31449 ( .A(n30702), .B(n30703), .Z(n30709) );
  NANDN U31450 ( .A(n30653), .B(n42093), .Z(n30655) );
  XOR U31451 ( .A(n42134), .B(a[744]), .Z(n30694) );
  NANDN U31452 ( .A(n30694), .B(n42095), .Z(n30654) );
  NAND U31453 ( .A(n30655), .B(n30654), .Z(n30707) );
  NANDN U31454 ( .A(n30656), .B(n42231), .Z(n30658) );
  XOR U31455 ( .A(n223), .B(a[740]), .Z(n30697) );
  NANDN U31456 ( .A(n30697), .B(n42234), .Z(n30657) );
  AND U31457 ( .A(n30658), .B(n30657), .Z(n30706) );
  XNOR U31458 ( .A(n30707), .B(n30706), .Z(n30708) );
  XNOR U31459 ( .A(n30709), .B(n30708), .Z(n30713) );
  NANDN U31460 ( .A(n30660), .B(n30659), .Z(n30664) );
  NAND U31461 ( .A(n30662), .B(n30661), .Z(n30663) );
  AND U31462 ( .A(n30664), .B(n30663), .Z(n30712) );
  XOR U31463 ( .A(n30713), .B(n30712), .Z(n30714) );
  NANDN U31464 ( .A(n30666), .B(n30665), .Z(n30670) );
  NANDN U31465 ( .A(n30668), .B(n30667), .Z(n30669) );
  NAND U31466 ( .A(n30670), .B(n30669), .Z(n30715) );
  XOR U31467 ( .A(n30714), .B(n30715), .Z(n30682) );
  OR U31468 ( .A(n30672), .B(n30671), .Z(n30676) );
  NANDN U31469 ( .A(n30674), .B(n30673), .Z(n30675) );
  NAND U31470 ( .A(n30676), .B(n30675), .Z(n30683) );
  XNOR U31471 ( .A(n30682), .B(n30683), .Z(n30684) );
  XNOR U31472 ( .A(n30685), .B(n30684), .Z(n30718) );
  XNOR U31473 ( .A(n30718), .B(sreg[1762]), .Z(n30720) );
  NAND U31474 ( .A(n30677), .B(sreg[1761]), .Z(n30681) );
  OR U31475 ( .A(n30679), .B(n30678), .Z(n30680) );
  AND U31476 ( .A(n30681), .B(n30680), .Z(n30719) );
  XOR U31477 ( .A(n30720), .B(n30719), .Z(c[1762]) );
  NANDN U31478 ( .A(n30683), .B(n30682), .Z(n30687) );
  NAND U31479 ( .A(n30685), .B(n30684), .Z(n30686) );
  NAND U31480 ( .A(n30687), .B(n30686), .Z(n30726) );
  NAND U31481 ( .A(b[0]), .B(a[747]), .Z(n30688) );
  XNOR U31482 ( .A(b[1]), .B(n30688), .Z(n30690) );
  NAND U31483 ( .A(n121), .B(a[746]), .Z(n30689) );
  AND U31484 ( .A(n30690), .B(n30689), .Z(n30743) );
  XOR U31485 ( .A(a[743]), .B(n42197), .Z(n30732) );
  NANDN U31486 ( .A(n30732), .B(n42173), .Z(n30693) );
  NANDN U31487 ( .A(n30691), .B(n42172), .Z(n30692) );
  NAND U31488 ( .A(n30693), .B(n30692), .Z(n30741) );
  NAND U31489 ( .A(b[7]), .B(a[739]), .Z(n30742) );
  XNOR U31490 ( .A(n30741), .B(n30742), .Z(n30744) );
  XOR U31491 ( .A(n30743), .B(n30744), .Z(n30750) );
  NANDN U31492 ( .A(n30694), .B(n42093), .Z(n30696) );
  XOR U31493 ( .A(n42134), .B(a[745]), .Z(n30735) );
  NANDN U31494 ( .A(n30735), .B(n42095), .Z(n30695) );
  NAND U31495 ( .A(n30696), .B(n30695), .Z(n30748) );
  NANDN U31496 ( .A(n30697), .B(n42231), .Z(n30699) );
  XOR U31497 ( .A(n223), .B(a[741]), .Z(n30738) );
  NANDN U31498 ( .A(n30738), .B(n42234), .Z(n30698) );
  AND U31499 ( .A(n30699), .B(n30698), .Z(n30747) );
  XNOR U31500 ( .A(n30748), .B(n30747), .Z(n30749) );
  XNOR U31501 ( .A(n30750), .B(n30749), .Z(n30754) );
  NANDN U31502 ( .A(n30701), .B(n30700), .Z(n30705) );
  NAND U31503 ( .A(n30703), .B(n30702), .Z(n30704) );
  AND U31504 ( .A(n30705), .B(n30704), .Z(n30753) );
  XOR U31505 ( .A(n30754), .B(n30753), .Z(n30755) );
  NANDN U31506 ( .A(n30707), .B(n30706), .Z(n30711) );
  NANDN U31507 ( .A(n30709), .B(n30708), .Z(n30710) );
  NAND U31508 ( .A(n30711), .B(n30710), .Z(n30756) );
  XOR U31509 ( .A(n30755), .B(n30756), .Z(n30723) );
  OR U31510 ( .A(n30713), .B(n30712), .Z(n30717) );
  NANDN U31511 ( .A(n30715), .B(n30714), .Z(n30716) );
  NAND U31512 ( .A(n30717), .B(n30716), .Z(n30724) );
  XNOR U31513 ( .A(n30723), .B(n30724), .Z(n30725) );
  XNOR U31514 ( .A(n30726), .B(n30725), .Z(n30759) );
  XNOR U31515 ( .A(n30759), .B(sreg[1763]), .Z(n30761) );
  NAND U31516 ( .A(n30718), .B(sreg[1762]), .Z(n30722) );
  OR U31517 ( .A(n30720), .B(n30719), .Z(n30721) );
  AND U31518 ( .A(n30722), .B(n30721), .Z(n30760) );
  XOR U31519 ( .A(n30761), .B(n30760), .Z(c[1763]) );
  NANDN U31520 ( .A(n30724), .B(n30723), .Z(n30728) );
  NAND U31521 ( .A(n30726), .B(n30725), .Z(n30727) );
  NAND U31522 ( .A(n30728), .B(n30727), .Z(n30767) );
  NAND U31523 ( .A(b[0]), .B(a[748]), .Z(n30729) );
  XNOR U31524 ( .A(b[1]), .B(n30729), .Z(n30731) );
  NAND U31525 ( .A(n121), .B(a[747]), .Z(n30730) );
  AND U31526 ( .A(n30731), .B(n30730), .Z(n30784) );
  XOR U31527 ( .A(a[744]), .B(n42197), .Z(n30773) );
  NANDN U31528 ( .A(n30773), .B(n42173), .Z(n30734) );
  NANDN U31529 ( .A(n30732), .B(n42172), .Z(n30733) );
  NAND U31530 ( .A(n30734), .B(n30733), .Z(n30782) );
  NAND U31531 ( .A(b[7]), .B(a[740]), .Z(n30783) );
  XNOR U31532 ( .A(n30782), .B(n30783), .Z(n30785) );
  XOR U31533 ( .A(n30784), .B(n30785), .Z(n30791) );
  NANDN U31534 ( .A(n30735), .B(n42093), .Z(n30737) );
  XOR U31535 ( .A(n42134), .B(a[746]), .Z(n30776) );
  NANDN U31536 ( .A(n30776), .B(n42095), .Z(n30736) );
  NAND U31537 ( .A(n30737), .B(n30736), .Z(n30789) );
  NANDN U31538 ( .A(n30738), .B(n42231), .Z(n30740) );
  XOR U31539 ( .A(n223), .B(a[742]), .Z(n30779) );
  NANDN U31540 ( .A(n30779), .B(n42234), .Z(n30739) );
  AND U31541 ( .A(n30740), .B(n30739), .Z(n30788) );
  XNOR U31542 ( .A(n30789), .B(n30788), .Z(n30790) );
  XNOR U31543 ( .A(n30791), .B(n30790), .Z(n30795) );
  NANDN U31544 ( .A(n30742), .B(n30741), .Z(n30746) );
  NAND U31545 ( .A(n30744), .B(n30743), .Z(n30745) );
  AND U31546 ( .A(n30746), .B(n30745), .Z(n30794) );
  XOR U31547 ( .A(n30795), .B(n30794), .Z(n30796) );
  NANDN U31548 ( .A(n30748), .B(n30747), .Z(n30752) );
  NANDN U31549 ( .A(n30750), .B(n30749), .Z(n30751) );
  NAND U31550 ( .A(n30752), .B(n30751), .Z(n30797) );
  XOR U31551 ( .A(n30796), .B(n30797), .Z(n30764) );
  OR U31552 ( .A(n30754), .B(n30753), .Z(n30758) );
  NANDN U31553 ( .A(n30756), .B(n30755), .Z(n30757) );
  NAND U31554 ( .A(n30758), .B(n30757), .Z(n30765) );
  XNOR U31555 ( .A(n30764), .B(n30765), .Z(n30766) );
  XNOR U31556 ( .A(n30767), .B(n30766), .Z(n30800) );
  XNOR U31557 ( .A(n30800), .B(sreg[1764]), .Z(n30802) );
  NAND U31558 ( .A(n30759), .B(sreg[1763]), .Z(n30763) );
  OR U31559 ( .A(n30761), .B(n30760), .Z(n30762) );
  AND U31560 ( .A(n30763), .B(n30762), .Z(n30801) );
  XOR U31561 ( .A(n30802), .B(n30801), .Z(c[1764]) );
  NANDN U31562 ( .A(n30765), .B(n30764), .Z(n30769) );
  NAND U31563 ( .A(n30767), .B(n30766), .Z(n30768) );
  NAND U31564 ( .A(n30769), .B(n30768), .Z(n30808) );
  NAND U31565 ( .A(b[0]), .B(a[749]), .Z(n30770) );
  XNOR U31566 ( .A(b[1]), .B(n30770), .Z(n30772) );
  NAND U31567 ( .A(n122), .B(a[748]), .Z(n30771) );
  AND U31568 ( .A(n30772), .B(n30771), .Z(n30825) );
  XOR U31569 ( .A(a[745]), .B(n42197), .Z(n30814) );
  NANDN U31570 ( .A(n30814), .B(n42173), .Z(n30775) );
  NANDN U31571 ( .A(n30773), .B(n42172), .Z(n30774) );
  NAND U31572 ( .A(n30775), .B(n30774), .Z(n30823) );
  NAND U31573 ( .A(b[7]), .B(a[741]), .Z(n30824) );
  XNOR U31574 ( .A(n30823), .B(n30824), .Z(n30826) );
  XOR U31575 ( .A(n30825), .B(n30826), .Z(n30832) );
  NANDN U31576 ( .A(n30776), .B(n42093), .Z(n30778) );
  XOR U31577 ( .A(n42134), .B(a[747]), .Z(n30817) );
  NANDN U31578 ( .A(n30817), .B(n42095), .Z(n30777) );
  NAND U31579 ( .A(n30778), .B(n30777), .Z(n30830) );
  NANDN U31580 ( .A(n30779), .B(n42231), .Z(n30781) );
  XOR U31581 ( .A(n224), .B(a[743]), .Z(n30820) );
  NANDN U31582 ( .A(n30820), .B(n42234), .Z(n30780) );
  AND U31583 ( .A(n30781), .B(n30780), .Z(n30829) );
  XNOR U31584 ( .A(n30830), .B(n30829), .Z(n30831) );
  XNOR U31585 ( .A(n30832), .B(n30831), .Z(n30836) );
  NANDN U31586 ( .A(n30783), .B(n30782), .Z(n30787) );
  NAND U31587 ( .A(n30785), .B(n30784), .Z(n30786) );
  AND U31588 ( .A(n30787), .B(n30786), .Z(n30835) );
  XOR U31589 ( .A(n30836), .B(n30835), .Z(n30837) );
  NANDN U31590 ( .A(n30789), .B(n30788), .Z(n30793) );
  NANDN U31591 ( .A(n30791), .B(n30790), .Z(n30792) );
  NAND U31592 ( .A(n30793), .B(n30792), .Z(n30838) );
  XOR U31593 ( .A(n30837), .B(n30838), .Z(n30805) );
  OR U31594 ( .A(n30795), .B(n30794), .Z(n30799) );
  NANDN U31595 ( .A(n30797), .B(n30796), .Z(n30798) );
  NAND U31596 ( .A(n30799), .B(n30798), .Z(n30806) );
  XNOR U31597 ( .A(n30805), .B(n30806), .Z(n30807) );
  XNOR U31598 ( .A(n30808), .B(n30807), .Z(n30841) );
  XNOR U31599 ( .A(n30841), .B(sreg[1765]), .Z(n30843) );
  NAND U31600 ( .A(n30800), .B(sreg[1764]), .Z(n30804) );
  OR U31601 ( .A(n30802), .B(n30801), .Z(n30803) );
  AND U31602 ( .A(n30804), .B(n30803), .Z(n30842) );
  XOR U31603 ( .A(n30843), .B(n30842), .Z(c[1765]) );
  NANDN U31604 ( .A(n30806), .B(n30805), .Z(n30810) );
  NAND U31605 ( .A(n30808), .B(n30807), .Z(n30809) );
  NAND U31606 ( .A(n30810), .B(n30809), .Z(n30849) );
  NAND U31607 ( .A(b[0]), .B(a[750]), .Z(n30811) );
  XNOR U31608 ( .A(b[1]), .B(n30811), .Z(n30813) );
  NAND U31609 ( .A(n122), .B(a[749]), .Z(n30812) );
  AND U31610 ( .A(n30813), .B(n30812), .Z(n30866) );
  XOR U31611 ( .A(a[746]), .B(n42197), .Z(n30855) );
  NANDN U31612 ( .A(n30855), .B(n42173), .Z(n30816) );
  NANDN U31613 ( .A(n30814), .B(n42172), .Z(n30815) );
  NAND U31614 ( .A(n30816), .B(n30815), .Z(n30864) );
  NAND U31615 ( .A(b[7]), .B(a[742]), .Z(n30865) );
  XNOR U31616 ( .A(n30864), .B(n30865), .Z(n30867) );
  XOR U31617 ( .A(n30866), .B(n30867), .Z(n30873) );
  NANDN U31618 ( .A(n30817), .B(n42093), .Z(n30819) );
  XOR U31619 ( .A(n42134), .B(a[748]), .Z(n30858) );
  NANDN U31620 ( .A(n30858), .B(n42095), .Z(n30818) );
  NAND U31621 ( .A(n30819), .B(n30818), .Z(n30871) );
  NANDN U31622 ( .A(n30820), .B(n42231), .Z(n30822) );
  XOR U31623 ( .A(n224), .B(a[744]), .Z(n30861) );
  NANDN U31624 ( .A(n30861), .B(n42234), .Z(n30821) );
  AND U31625 ( .A(n30822), .B(n30821), .Z(n30870) );
  XNOR U31626 ( .A(n30871), .B(n30870), .Z(n30872) );
  XNOR U31627 ( .A(n30873), .B(n30872), .Z(n30877) );
  NANDN U31628 ( .A(n30824), .B(n30823), .Z(n30828) );
  NAND U31629 ( .A(n30826), .B(n30825), .Z(n30827) );
  AND U31630 ( .A(n30828), .B(n30827), .Z(n30876) );
  XOR U31631 ( .A(n30877), .B(n30876), .Z(n30878) );
  NANDN U31632 ( .A(n30830), .B(n30829), .Z(n30834) );
  NANDN U31633 ( .A(n30832), .B(n30831), .Z(n30833) );
  NAND U31634 ( .A(n30834), .B(n30833), .Z(n30879) );
  XOR U31635 ( .A(n30878), .B(n30879), .Z(n30846) );
  OR U31636 ( .A(n30836), .B(n30835), .Z(n30840) );
  NANDN U31637 ( .A(n30838), .B(n30837), .Z(n30839) );
  NAND U31638 ( .A(n30840), .B(n30839), .Z(n30847) );
  XNOR U31639 ( .A(n30846), .B(n30847), .Z(n30848) );
  XNOR U31640 ( .A(n30849), .B(n30848), .Z(n30882) );
  XNOR U31641 ( .A(n30882), .B(sreg[1766]), .Z(n30884) );
  NAND U31642 ( .A(n30841), .B(sreg[1765]), .Z(n30845) );
  OR U31643 ( .A(n30843), .B(n30842), .Z(n30844) );
  AND U31644 ( .A(n30845), .B(n30844), .Z(n30883) );
  XOR U31645 ( .A(n30884), .B(n30883), .Z(c[1766]) );
  NANDN U31646 ( .A(n30847), .B(n30846), .Z(n30851) );
  NAND U31647 ( .A(n30849), .B(n30848), .Z(n30850) );
  NAND U31648 ( .A(n30851), .B(n30850), .Z(n30890) );
  NAND U31649 ( .A(b[0]), .B(a[751]), .Z(n30852) );
  XNOR U31650 ( .A(b[1]), .B(n30852), .Z(n30854) );
  NAND U31651 ( .A(n122), .B(a[750]), .Z(n30853) );
  AND U31652 ( .A(n30854), .B(n30853), .Z(n30907) );
  XOR U31653 ( .A(a[747]), .B(n42197), .Z(n30896) );
  NANDN U31654 ( .A(n30896), .B(n42173), .Z(n30857) );
  NANDN U31655 ( .A(n30855), .B(n42172), .Z(n30856) );
  NAND U31656 ( .A(n30857), .B(n30856), .Z(n30905) );
  NAND U31657 ( .A(b[7]), .B(a[743]), .Z(n30906) );
  XNOR U31658 ( .A(n30905), .B(n30906), .Z(n30908) );
  XOR U31659 ( .A(n30907), .B(n30908), .Z(n30914) );
  NANDN U31660 ( .A(n30858), .B(n42093), .Z(n30860) );
  XOR U31661 ( .A(n42134), .B(a[749]), .Z(n30899) );
  NANDN U31662 ( .A(n30899), .B(n42095), .Z(n30859) );
  NAND U31663 ( .A(n30860), .B(n30859), .Z(n30912) );
  NANDN U31664 ( .A(n30861), .B(n42231), .Z(n30863) );
  XOR U31665 ( .A(n224), .B(a[745]), .Z(n30902) );
  NANDN U31666 ( .A(n30902), .B(n42234), .Z(n30862) );
  AND U31667 ( .A(n30863), .B(n30862), .Z(n30911) );
  XNOR U31668 ( .A(n30912), .B(n30911), .Z(n30913) );
  XNOR U31669 ( .A(n30914), .B(n30913), .Z(n30918) );
  NANDN U31670 ( .A(n30865), .B(n30864), .Z(n30869) );
  NAND U31671 ( .A(n30867), .B(n30866), .Z(n30868) );
  AND U31672 ( .A(n30869), .B(n30868), .Z(n30917) );
  XOR U31673 ( .A(n30918), .B(n30917), .Z(n30919) );
  NANDN U31674 ( .A(n30871), .B(n30870), .Z(n30875) );
  NANDN U31675 ( .A(n30873), .B(n30872), .Z(n30874) );
  NAND U31676 ( .A(n30875), .B(n30874), .Z(n30920) );
  XOR U31677 ( .A(n30919), .B(n30920), .Z(n30887) );
  OR U31678 ( .A(n30877), .B(n30876), .Z(n30881) );
  NANDN U31679 ( .A(n30879), .B(n30878), .Z(n30880) );
  NAND U31680 ( .A(n30881), .B(n30880), .Z(n30888) );
  XNOR U31681 ( .A(n30887), .B(n30888), .Z(n30889) );
  XNOR U31682 ( .A(n30890), .B(n30889), .Z(n30923) );
  XNOR U31683 ( .A(n30923), .B(sreg[1767]), .Z(n30925) );
  NAND U31684 ( .A(n30882), .B(sreg[1766]), .Z(n30886) );
  OR U31685 ( .A(n30884), .B(n30883), .Z(n30885) );
  AND U31686 ( .A(n30886), .B(n30885), .Z(n30924) );
  XOR U31687 ( .A(n30925), .B(n30924), .Z(c[1767]) );
  NANDN U31688 ( .A(n30888), .B(n30887), .Z(n30892) );
  NAND U31689 ( .A(n30890), .B(n30889), .Z(n30891) );
  NAND U31690 ( .A(n30892), .B(n30891), .Z(n30931) );
  NAND U31691 ( .A(b[0]), .B(a[752]), .Z(n30893) );
  XNOR U31692 ( .A(b[1]), .B(n30893), .Z(n30895) );
  NAND U31693 ( .A(n122), .B(a[751]), .Z(n30894) );
  AND U31694 ( .A(n30895), .B(n30894), .Z(n30948) );
  XOR U31695 ( .A(a[748]), .B(n42197), .Z(n30937) );
  NANDN U31696 ( .A(n30937), .B(n42173), .Z(n30898) );
  NANDN U31697 ( .A(n30896), .B(n42172), .Z(n30897) );
  NAND U31698 ( .A(n30898), .B(n30897), .Z(n30946) );
  NAND U31699 ( .A(b[7]), .B(a[744]), .Z(n30947) );
  XNOR U31700 ( .A(n30946), .B(n30947), .Z(n30949) );
  XOR U31701 ( .A(n30948), .B(n30949), .Z(n30955) );
  NANDN U31702 ( .A(n30899), .B(n42093), .Z(n30901) );
  XOR U31703 ( .A(n42134), .B(a[750]), .Z(n30940) );
  NANDN U31704 ( .A(n30940), .B(n42095), .Z(n30900) );
  NAND U31705 ( .A(n30901), .B(n30900), .Z(n30953) );
  NANDN U31706 ( .A(n30902), .B(n42231), .Z(n30904) );
  XOR U31707 ( .A(n224), .B(a[746]), .Z(n30943) );
  NANDN U31708 ( .A(n30943), .B(n42234), .Z(n30903) );
  AND U31709 ( .A(n30904), .B(n30903), .Z(n30952) );
  XNOR U31710 ( .A(n30953), .B(n30952), .Z(n30954) );
  XNOR U31711 ( .A(n30955), .B(n30954), .Z(n30959) );
  NANDN U31712 ( .A(n30906), .B(n30905), .Z(n30910) );
  NAND U31713 ( .A(n30908), .B(n30907), .Z(n30909) );
  AND U31714 ( .A(n30910), .B(n30909), .Z(n30958) );
  XOR U31715 ( .A(n30959), .B(n30958), .Z(n30960) );
  NANDN U31716 ( .A(n30912), .B(n30911), .Z(n30916) );
  NANDN U31717 ( .A(n30914), .B(n30913), .Z(n30915) );
  NAND U31718 ( .A(n30916), .B(n30915), .Z(n30961) );
  XOR U31719 ( .A(n30960), .B(n30961), .Z(n30928) );
  OR U31720 ( .A(n30918), .B(n30917), .Z(n30922) );
  NANDN U31721 ( .A(n30920), .B(n30919), .Z(n30921) );
  NAND U31722 ( .A(n30922), .B(n30921), .Z(n30929) );
  XNOR U31723 ( .A(n30928), .B(n30929), .Z(n30930) );
  XNOR U31724 ( .A(n30931), .B(n30930), .Z(n30964) );
  XNOR U31725 ( .A(n30964), .B(sreg[1768]), .Z(n30966) );
  NAND U31726 ( .A(n30923), .B(sreg[1767]), .Z(n30927) );
  OR U31727 ( .A(n30925), .B(n30924), .Z(n30926) );
  AND U31728 ( .A(n30927), .B(n30926), .Z(n30965) );
  XOR U31729 ( .A(n30966), .B(n30965), .Z(c[1768]) );
  NANDN U31730 ( .A(n30929), .B(n30928), .Z(n30933) );
  NAND U31731 ( .A(n30931), .B(n30930), .Z(n30932) );
  NAND U31732 ( .A(n30933), .B(n30932), .Z(n30972) );
  NAND U31733 ( .A(b[0]), .B(a[753]), .Z(n30934) );
  XNOR U31734 ( .A(b[1]), .B(n30934), .Z(n30936) );
  NAND U31735 ( .A(n122), .B(a[752]), .Z(n30935) );
  AND U31736 ( .A(n30936), .B(n30935), .Z(n30989) );
  XOR U31737 ( .A(a[749]), .B(n42197), .Z(n30978) );
  NANDN U31738 ( .A(n30978), .B(n42173), .Z(n30939) );
  NANDN U31739 ( .A(n30937), .B(n42172), .Z(n30938) );
  NAND U31740 ( .A(n30939), .B(n30938), .Z(n30987) );
  NAND U31741 ( .A(b[7]), .B(a[745]), .Z(n30988) );
  XNOR U31742 ( .A(n30987), .B(n30988), .Z(n30990) );
  XOR U31743 ( .A(n30989), .B(n30990), .Z(n30996) );
  NANDN U31744 ( .A(n30940), .B(n42093), .Z(n30942) );
  XOR U31745 ( .A(n42134), .B(a[751]), .Z(n30981) );
  NANDN U31746 ( .A(n30981), .B(n42095), .Z(n30941) );
  NAND U31747 ( .A(n30942), .B(n30941), .Z(n30994) );
  NANDN U31748 ( .A(n30943), .B(n42231), .Z(n30945) );
  XOR U31749 ( .A(n224), .B(a[747]), .Z(n30984) );
  NANDN U31750 ( .A(n30984), .B(n42234), .Z(n30944) );
  AND U31751 ( .A(n30945), .B(n30944), .Z(n30993) );
  XNOR U31752 ( .A(n30994), .B(n30993), .Z(n30995) );
  XNOR U31753 ( .A(n30996), .B(n30995), .Z(n31000) );
  NANDN U31754 ( .A(n30947), .B(n30946), .Z(n30951) );
  NAND U31755 ( .A(n30949), .B(n30948), .Z(n30950) );
  AND U31756 ( .A(n30951), .B(n30950), .Z(n30999) );
  XOR U31757 ( .A(n31000), .B(n30999), .Z(n31001) );
  NANDN U31758 ( .A(n30953), .B(n30952), .Z(n30957) );
  NANDN U31759 ( .A(n30955), .B(n30954), .Z(n30956) );
  NAND U31760 ( .A(n30957), .B(n30956), .Z(n31002) );
  XOR U31761 ( .A(n31001), .B(n31002), .Z(n30969) );
  OR U31762 ( .A(n30959), .B(n30958), .Z(n30963) );
  NANDN U31763 ( .A(n30961), .B(n30960), .Z(n30962) );
  NAND U31764 ( .A(n30963), .B(n30962), .Z(n30970) );
  XNOR U31765 ( .A(n30969), .B(n30970), .Z(n30971) );
  XNOR U31766 ( .A(n30972), .B(n30971), .Z(n31005) );
  XNOR U31767 ( .A(n31005), .B(sreg[1769]), .Z(n31007) );
  NAND U31768 ( .A(n30964), .B(sreg[1768]), .Z(n30968) );
  OR U31769 ( .A(n30966), .B(n30965), .Z(n30967) );
  AND U31770 ( .A(n30968), .B(n30967), .Z(n31006) );
  XOR U31771 ( .A(n31007), .B(n31006), .Z(c[1769]) );
  NANDN U31772 ( .A(n30970), .B(n30969), .Z(n30974) );
  NAND U31773 ( .A(n30972), .B(n30971), .Z(n30973) );
  NAND U31774 ( .A(n30974), .B(n30973), .Z(n31013) );
  NAND U31775 ( .A(b[0]), .B(a[754]), .Z(n30975) );
  XNOR U31776 ( .A(b[1]), .B(n30975), .Z(n30977) );
  NAND U31777 ( .A(n122), .B(a[753]), .Z(n30976) );
  AND U31778 ( .A(n30977), .B(n30976), .Z(n31030) );
  XOR U31779 ( .A(a[750]), .B(n42197), .Z(n31019) );
  NANDN U31780 ( .A(n31019), .B(n42173), .Z(n30980) );
  NANDN U31781 ( .A(n30978), .B(n42172), .Z(n30979) );
  NAND U31782 ( .A(n30980), .B(n30979), .Z(n31028) );
  NAND U31783 ( .A(b[7]), .B(a[746]), .Z(n31029) );
  XNOR U31784 ( .A(n31028), .B(n31029), .Z(n31031) );
  XOR U31785 ( .A(n31030), .B(n31031), .Z(n31037) );
  NANDN U31786 ( .A(n30981), .B(n42093), .Z(n30983) );
  XOR U31787 ( .A(n42134), .B(a[752]), .Z(n31022) );
  NANDN U31788 ( .A(n31022), .B(n42095), .Z(n30982) );
  NAND U31789 ( .A(n30983), .B(n30982), .Z(n31035) );
  NANDN U31790 ( .A(n30984), .B(n42231), .Z(n30986) );
  XOR U31791 ( .A(n224), .B(a[748]), .Z(n31025) );
  NANDN U31792 ( .A(n31025), .B(n42234), .Z(n30985) );
  AND U31793 ( .A(n30986), .B(n30985), .Z(n31034) );
  XNOR U31794 ( .A(n31035), .B(n31034), .Z(n31036) );
  XNOR U31795 ( .A(n31037), .B(n31036), .Z(n31041) );
  NANDN U31796 ( .A(n30988), .B(n30987), .Z(n30992) );
  NAND U31797 ( .A(n30990), .B(n30989), .Z(n30991) );
  AND U31798 ( .A(n30992), .B(n30991), .Z(n31040) );
  XOR U31799 ( .A(n31041), .B(n31040), .Z(n31042) );
  NANDN U31800 ( .A(n30994), .B(n30993), .Z(n30998) );
  NANDN U31801 ( .A(n30996), .B(n30995), .Z(n30997) );
  NAND U31802 ( .A(n30998), .B(n30997), .Z(n31043) );
  XOR U31803 ( .A(n31042), .B(n31043), .Z(n31010) );
  OR U31804 ( .A(n31000), .B(n30999), .Z(n31004) );
  NANDN U31805 ( .A(n31002), .B(n31001), .Z(n31003) );
  NAND U31806 ( .A(n31004), .B(n31003), .Z(n31011) );
  XNOR U31807 ( .A(n31010), .B(n31011), .Z(n31012) );
  XNOR U31808 ( .A(n31013), .B(n31012), .Z(n31046) );
  XNOR U31809 ( .A(n31046), .B(sreg[1770]), .Z(n31048) );
  NAND U31810 ( .A(n31005), .B(sreg[1769]), .Z(n31009) );
  OR U31811 ( .A(n31007), .B(n31006), .Z(n31008) );
  AND U31812 ( .A(n31009), .B(n31008), .Z(n31047) );
  XOR U31813 ( .A(n31048), .B(n31047), .Z(c[1770]) );
  NANDN U31814 ( .A(n31011), .B(n31010), .Z(n31015) );
  NAND U31815 ( .A(n31013), .B(n31012), .Z(n31014) );
  NAND U31816 ( .A(n31015), .B(n31014), .Z(n31054) );
  NAND U31817 ( .A(b[0]), .B(a[755]), .Z(n31016) );
  XNOR U31818 ( .A(b[1]), .B(n31016), .Z(n31018) );
  NAND U31819 ( .A(n122), .B(a[754]), .Z(n31017) );
  AND U31820 ( .A(n31018), .B(n31017), .Z(n31071) );
  XOR U31821 ( .A(a[751]), .B(n42197), .Z(n31060) );
  NANDN U31822 ( .A(n31060), .B(n42173), .Z(n31021) );
  NANDN U31823 ( .A(n31019), .B(n42172), .Z(n31020) );
  NAND U31824 ( .A(n31021), .B(n31020), .Z(n31069) );
  NAND U31825 ( .A(b[7]), .B(a[747]), .Z(n31070) );
  XNOR U31826 ( .A(n31069), .B(n31070), .Z(n31072) );
  XOR U31827 ( .A(n31071), .B(n31072), .Z(n31078) );
  NANDN U31828 ( .A(n31022), .B(n42093), .Z(n31024) );
  XOR U31829 ( .A(n42134), .B(a[753]), .Z(n31063) );
  NANDN U31830 ( .A(n31063), .B(n42095), .Z(n31023) );
  NAND U31831 ( .A(n31024), .B(n31023), .Z(n31076) );
  NANDN U31832 ( .A(n31025), .B(n42231), .Z(n31027) );
  XOR U31833 ( .A(n224), .B(a[749]), .Z(n31066) );
  NANDN U31834 ( .A(n31066), .B(n42234), .Z(n31026) );
  AND U31835 ( .A(n31027), .B(n31026), .Z(n31075) );
  XNOR U31836 ( .A(n31076), .B(n31075), .Z(n31077) );
  XNOR U31837 ( .A(n31078), .B(n31077), .Z(n31082) );
  NANDN U31838 ( .A(n31029), .B(n31028), .Z(n31033) );
  NAND U31839 ( .A(n31031), .B(n31030), .Z(n31032) );
  AND U31840 ( .A(n31033), .B(n31032), .Z(n31081) );
  XOR U31841 ( .A(n31082), .B(n31081), .Z(n31083) );
  NANDN U31842 ( .A(n31035), .B(n31034), .Z(n31039) );
  NANDN U31843 ( .A(n31037), .B(n31036), .Z(n31038) );
  NAND U31844 ( .A(n31039), .B(n31038), .Z(n31084) );
  XOR U31845 ( .A(n31083), .B(n31084), .Z(n31051) );
  OR U31846 ( .A(n31041), .B(n31040), .Z(n31045) );
  NANDN U31847 ( .A(n31043), .B(n31042), .Z(n31044) );
  NAND U31848 ( .A(n31045), .B(n31044), .Z(n31052) );
  XNOR U31849 ( .A(n31051), .B(n31052), .Z(n31053) );
  XNOR U31850 ( .A(n31054), .B(n31053), .Z(n31087) );
  XNOR U31851 ( .A(n31087), .B(sreg[1771]), .Z(n31089) );
  NAND U31852 ( .A(n31046), .B(sreg[1770]), .Z(n31050) );
  OR U31853 ( .A(n31048), .B(n31047), .Z(n31049) );
  AND U31854 ( .A(n31050), .B(n31049), .Z(n31088) );
  XOR U31855 ( .A(n31089), .B(n31088), .Z(c[1771]) );
  NANDN U31856 ( .A(n31052), .B(n31051), .Z(n31056) );
  NAND U31857 ( .A(n31054), .B(n31053), .Z(n31055) );
  NAND U31858 ( .A(n31056), .B(n31055), .Z(n31095) );
  NAND U31859 ( .A(b[0]), .B(a[756]), .Z(n31057) );
  XNOR U31860 ( .A(b[1]), .B(n31057), .Z(n31059) );
  NAND U31861 ( .A(n123), .B(a[755]), .Z(n31058) );
  AND U31862 ( .A(n31059), .B(n31058), .Z(n31112) );
  XOR U31863 ( .A(a[752]), .B(n42197), .Z(n31101) );
  NANDN U31864 ( .A(n31101), .B(n42173), .Z(n31062) );
  NANDN U31865 ( .A(n31060), .B(n42172), .Z(n31061) );
  NAND U31866 ( .A(n31062), .B(n31061), .Z(n31110) );
  NAND U31867 ( .A(b[7]), .B(a[748]), .Z(n31111) );
  XNOR U31868 ( .A(n31110), .B(n31111), .Z(n31113) );
  XOR U31869 ( .A(n31112), .B(n31113), .Z(n31119) );
  NANDN U31870 ( .A(n31063), .B(n42093), .Z(n31065) );
  XOR U31871 ( .A(n42134), .B(a[754]), .Z(n31104) );
  NANDN U31872 ( .A(n31104), .B(n42095), .Z(n31064) );
  NAND U31873 ( .A(n31065), .B(n31064), .Z(n31117) );
  NANDN U31874 ( .A(n31066), .B(n42231), .Z(n31068) );
  XOR U31875 ( .A(n224), .B(a[750]), .Z(n31107) );
  NANDN U31876 ( .A(n31107), .B(n42234), .Z(n31067) );
  AND U31877 ( .A(n31068), .B(n31067), .Z(n31116) );
  XNOR U31878 ( .A(n31117), .B(n31116), .Z(n31118) );
  XNOR U31879 ( .A(n31119), .B(n31118), .Z(n31123) );
  NANDN U31880 ( .A(n31070), .B(n31069), .Z(n31074) );
  NAND U31881 ( .A(n31072), .B(n31071), .Z(n31073) );
  AND U31882 ( .A(n31074), .B(n31073), .Z(n31122) );
  XOR U31883 ( .A(n31123), .B(n31122), .Z(n31124) );
  NANDN U31884 ( .A(n31076), .B(n31075), .Z(n31080) );
  NANDN U31885 ( .A(n31078), .B(n31077), .Z(n31079) );
  NAND U31886 ( .A(n31080), .B(n31079), .Z(n31125) );
  XOR U31887 ( .A(n31124), .B(n31125), .Z(n31092) );
  OR U31888 ( .A(n31082), .B(n31081), .Z(n31086) );
  NANDN U31889 ( .A(n31084), .B(n31083), .Z(n31085) );
  NAND U31890 ( .A(n31086), .B(n31085), .Z(n31093) );
  XNOR U31891 ( .A(n31092), .B(n31093), .Z(n31094) );
  XNOR U31892 ( .A(n31095), .B(n31094), .Z(n31128) );
  XNOR U31893 ( .A(n31128), .B(sreg[1772]), .Z(n31130) );
  NAND U31894 ( .A(n31087), .B(sreg[1771]), .Z(n31091) );
  OR U31895 ( .A(n31089), .B(n31088), .Z(n31090) );
  AND U31896 ( .A(n31091), .B(n31090), .Z(n31129) );
  XOR U31897 ( .A(n31130), .B(n31129), .Z(c[1772]) );
  NANDN U31898 ( .A(n31093), .B(n31092), .Z(n31097) );
  NAND U31899 ( .A(n31095), .B(n31094), .Z(n31096) );
  NAND U31900 ( .A(n31097), .B(n31096), .Z(n31136) );
  NAND U31901 ( .A(b[0]), .B(a[757]), .Z(n31098) );
  XNOR U31902 ( .A(b[1]), .B(n31098), .Z(n31100) );
  NAND U31903 ( .A(n123), .B(a[756]), .Z(n31099) );
  AND U31904 ( .A(n31100), .B(n31099), .Z(n31153) );
  XOR U31905 ( .A(a[753]), .B(n42197), .Z(n31142) );
  NANDN U31906 ( .A(n31142), .B(n42173), .Z(n31103) );
  NANDN U31907 ( .A(n31101), .B(n42172), .Z(n31102) );
  NAND U31908 ( .A(n31103), .B(n31102), .Z(n31151) );
  NAND U31909 ( .A(b[7]), .B(a[749]), .Z(n31152) );
  XNOR U31910 ( .A(n31151), .B(n31152), .Z(n31154) );
  XOR U31911 ( .A(n31153), .B(n31154), .Z(n31160) );
  NANDN U31912 ( .A(n31104), .B(n42093), .Z(n31106) );
  XOR U31913 ( .A(n42134), .B(a[755]), .Z(n31145) );
  NANDN U31914 ( .A(n31145), .B(n42095), .Z(n31105) );
  NAND U31915 ( .A(n31106), .B(n31105), .Z(n31158) );
  NANDN U31916 ( .A(n31107), .B(n42231), .Z(n31109) );
  XOR U31917 ( .A(n224), .B(a[751]), .Z(n31148) );
  NANDN U31918 ( .A(n31148), .B(n42234), .Z(n31108) );
  AND U31919 ( .A(n31109), .B(n31108), .Z(n31157) );
  XNOR U31920 ( .A(n31158), .B(n31157), .Z(n31159) );
  XNOR U31921 ( .A(n31160), .B(n31159), .Z(n31164) );
  NANDN U31922 ( .A(n31111), .B(n31110), .Z(n31115) );
  NAND U31923 ( .A(n31113), .B(n31112), .Z(n31114) );
  AND U31924 ( .A(n31115), .B(n31114), .Z(n31163) );
  XOR U31925 ( .A(n31164), .B(n31163), .Z(n31165) );
  NANDN U31926 ( .A(n31117), .B(n31116), .Z(n31121) );
  NANDN U31927 ( .A(n31119), .B(n31118), .Z(n31120) );
  NAND U31928 ( .A(n31121), .B(n31120), .Z(n31166) );
  XOR U31929 ( .A(n31165), .B(n31166), .Z(n31133) );
  OR U31930 ( .A(n31123), .B(n31122), .Z(n31127) );
  NANDN U31931 ( .A(n31125), .B(n31124), .Z(n31126) );
  NAND U31932 ( .A(n31127), .B(n31126), .Z(n31134) );
  XNOR U31933 ( .A(n31133), .B(n31134), .Z(n31135) );
  XNOR U31934 ( .A(n31136), .B(n31135), .Z(n31169) );
  XNOR U31935 ( .A(n31169), .B(sreg[1773]), .Z(n31171) );
  NAND U31936 ( .A(n31128), .B(sreg[1772]), .Z(n31132) );
  OR U31937 ( .A(n31130), .B(n31129), .Z(n31131) );
  AND U31938 ( .A(n31132), .B(n31131), .Z(n31170) );
  XOR U31939 ( .A(n31171), .B(n31170), .Z(c[1773]) );
  NANDN U31940 ( .A(n31134), .B(n31133), .Z(n31138) );
  NAND U31941 ( .A(n31136), .B(n31135), .Z(n31137) );
  NAND U31942 ( .A(n31138), .B(n31137), .Z(n31177) );
  NAND U31943 ( .A(b[0]), .B(a[758]), .Z(n31139) );
  XNOR U31944 ( .A(b[1]), .B(n31139), .Z(n31141) );
  NAND U31945 ( .A(n123), .B(a[757]), .Z(n31140) );
  AND U31946 ( .A(n31141), .B(n31140), .Z(n31194) );
  XOR U31947 ( .A(a[754]), .B(n42197), .Z(n31183) );
  NANDN U31948 ( .A(n31183), .B(n42173), .Z(n31144) );
  NANDN U31949 ( .A(n31142), .B(n42172), .Z(n31143) );
  NAND U31950 ( .A(n31144), .B(n31143), .Z(n31192) );
  NAND U31951 ( .A(b[7]), .B(a[750]), .Z(n31193) );
  XNOR U31952 ( .A(n31192), .B(n31193), .Z(n31195) );
  XOR U31953 ( .A(n31194), .B(n31195), .Z(n31201) );
  NANDN U31954 ( .A(n31145), .B(n42093), .Z(n31147) );
  XOR U31955 ( .A(n42134), .B(a[756]), .Z(n31186) );
  NANDN U31956 ( .A(n31186), .B(n42095), .Z(n31146) );
  NAND U31957 ( .A(n31147), .B(n31146), .Z(n31199) );
  NANDN U31958 ( .A(n31148), .B(n42231), .Z(n31150) );
  XOR U31959 ( .A(n224), .B(a[752]), .Z(n31189) );
  NANDN U31960 ( .A(n31189), .B(n42234), .Z(n31149) );
  AND U31961 ( .A(n31150), .B(n31149), .Z(n31198) );
  XNOR U31962 ( .A(n31199), .B(n31198), .Z(n31200) );
  XNOR U31963 ( .A(n31201), .B(n31200), .Z(n31205) );
  NANDN U31964 ( .A(n31152), .B(n31151), .Z(n31156) );
  NAND U31965 ( .A(n31154), .B(n31153), .Z(n31155) );
  AND U31966 ( .A(n31156), .B(n31155), .Z(n31204) );
  XOR U31967 ( .A(n31205), .B(n31204), .Z(n31206) );
  NANDN U31968 ( .A(n31158), .B(n31157), .Z(n31162) );
  NANDN U31969 ( .A(n31160), .B(n31159), .Z(n31161) );
  NAND U31970 ( .A(n31162), .B(n31161), .Z(n31207) );
  XOR U31971 ( .A(n31206), .B(n31207), .Z(n31174) );
  OR U31972 ( .A(n31164), .B(n31163), .Z(n31168) );
  NANDN U31973 ( .A(n31166), .B(n31165), .Z(n31167) );
  NAND U31974 ( .A(n31168), .B(n31167), .Z(n31175) );
  XNOR U31975 ( .A(n31174), .B(n31175), .Z(n31176) );
  XNOR U31976 ( .A(n31177), .B(n31176), .Z(n31210) );
  XNOR U31977 ( .A(n31210), .B(sreg[1774]), .Z(n31212) );
  NAND U31978 ( .A(n31169), .B(sreg[1773]), .Z(n31173) );
  OR U31979 ( .A(n31171), .B(n31170), .Z(n31172) );
  AND U31980 ( .A(n31173), .B(n31172), .Z(n31211) );
  XOR U31981 ( .A(n31212), .B(n31211), .Z(c[1774]) );
  NANDN U31982 ( .A(n31175), .B(n31174), .Z(n31179) );
  NAND U31983 ( .A(n31177), .B(n31176), .Z(n31178) );
  NAND U31984 ( .A(n31179), .B(n31178), .Z(n31218) );
  NAND U31985 ( .A(b[0]), .B(a[759]), .Z(n31180) );
  XNOR U31986 ( .A(b[1]), .B(n31180), .Z(n31182) );
  NAND U31987 ( .A(n123), .B(a[758]), .Z(n31181) );
  AND U31988 ( .A(n31182), .B(n31181), .Z(n31235) );
  XOR U31989 ( .A(a[755]), .B(n42197), .Z(n31224) );
  NANDN U31990 ( .A(n31224), .B(n42173), .Z(n31185) );
  NANDN U31991 ( .A(n31183), .B(n42172), .Z(n31184) );
  NAND U31992 ( .A(n31185), .B(n31184), .Z(n31233) );
  NAND U31993 ( .A(b[7]), .B(a[751]), .Z(n31234) );
  XNOR U31994 ( .A(n31233), .B(n31234), .Z(n31236) );
  XOR U31995 ( .A(n31235), .B(n31236), .Z(n31242) );
  NANDN U31996 ( .A(n31186), .B(n42093), .Z(n31188) );
  XOR U31997 ( .A(n42134), .B(a[757]), .Z(n31227) );
  NANDN U31998 ( .A(n31227), .B(n42095), .Z(n31187) );
  NAND U31999 ( .A(n31188), .B(n31187), .Z(n31240) );
  NANDN U32000 ( .A(n31189), .B(n42231), .Z(n31191) );
  XOR U32001 ( .A(n224), .B(a[753]), .Z(n31230) );
  NANDN U32002 ( .A(n31230), .B(n42234), .Z(n31190) );
  AND U32003 ( .A(n31191), .B(n31190), .Z(n31239) );
  XNOR U32004 ( .A(n31240), .B(n31239), .Z(n31241) );
  XNOR U32005 ( .A(n31242), .B(n31241), .Z(n31246) );
  NANDN U32006 ( .A(n31193), .B(n31192), .Z(n31197) );
  NAND U32007 ( .A(n31195), .B(n31194), .Z(n31196) );
  AND U32008 ( .A(n31197), .B(n31196), .Z(n31245) );
  XOR U32009 ( .A(n31246), .B(n31245), .Z(n31247) );
  NANDN U32010 ( .A(n31199), .B(n31198), .Z(n31203) );
  NANDN U32011 ( .A(n31201), .B(n31200), .Z(n31202) );
  NAND U32012 ( .A(n31203), .B(n31202), .Z(n31248) );
  XOR U32013 ( .A(n31247), .B(n31248), .Z(n31215) );
  OR U32014 ( .A(n31205), .B(n31204), .Z(n31209) );
  NANDN U32015 ( .A(n31207), .B(n31206), .Z(n31208) );
  NAND U32016 ( .A(n31209), .B(n31208), .Z(n31216) );
  XNOR U32017 ( .A(n31215), .B(n31216), .Z(n31217) );
  XNOR U32018 ( .A(n31218), .B(n31217), .Z(n31251) );
  XNOR U32019 ( .A(n31251), .B(sreg[1775]), .Z(n31253) );
  NAND U32020 ( .A(n31210), .B(sreg[1774]), .Z(n31214) );
  OR U32021 ( .A(n31212), .B(n31211), .Z(n31213) );
  AND U32022 ( .A(n31214), .B(n31213), .Z(n31252) );
  XOR U32023 ( .A(n31253), .B(n31252), .Z(c[1775]) );
  NANDN U32024 ( .A(n31216), .B(n31215), .Z(n31220) );
  NAND U32025 ( .A(n31218), .B(n31217), .Z(n31219) );
  NAND U32026 ( .A(n31220), .B(n31219), .Z(n31259) );
  NAND U32027 ( .A(b[0]), .B(a[760]), .Z(n31221) );
  XNOR U32028 ( .A(b[1]), .B(n31221), .Z(n31223) );
  NAND U32029 ( .A(n123), .B(a[759]), .Z(n31222) );
  AND U32030 ( .A(n31223), .B(n31222), .Z(n31276) );
  XOR U32031 ( .A(a[756]), .B(n42197), .Z(n31265) );
  NANDN U32032 ( .A(n31265), .B(n42173), .Z(n31226) );
  NANDN U32033 ( .A(n31224), .B(n42172), .Z(n31225) );
  NAND U32034 ( .A(n31226), .B(n31225), .Z(n31274) );
  NAND U32035 ( .A(b[7]), .B(a[752]), .Z(n31275) );
  XNOR U32036 ( .A(n31274), .B(n31275), .Z(n31277) );
  XOR U32037 ( .A(n31276), .B(n31277), .Z(n31283) );
  NANDN U32038 ( .A(n31227), .B(n42093), .Z(n31229) );
  XOR U32039 ( .A(n42134), .B(a[758]), .Z(n31268) );
  NANDN U32040 ( .A(n31268), .B(n42095), .Z(n31228) );
  NAND U32041 ( .A(n31229), .B(n31228), .Z(n31281) );
  NANDN U32042 ( .A(n31230), .B(n42231), .Z(n31232) );
  XOR U32043 ( .A(n224), .B(a[754]), .Z(n31271) );
  NANDN U32044 ( .A(n31271), .B(n42234), .Z(n31231) );
  AND U32045 ( .A(n31232), .B(n31231), .Z(n31280) );
  XNOR U32046 ( .A(n31281), .B(n31280), .Z(n31282) );
  XNOR U32047 ( .A(n31283), .B(n31282), .Z(n31287) );
  NANDN U32048 ( .A(n31234), .B(n31233), .Z(n31238) );
  NAND U32049 ( .A(n31236), .B(n31235), .Z(n31237) );
  AND U32050 ( .A(n31238), .B(n31237), .Z(n31286) );
  XOR U32051 ( .A(n31287), .B(n31286), .Z(n31288) );
  NANDN U32052 ( .A(n31240), .B(n31239), .Z(n31244) );
  NANDN U32053 ( .A(n31242), .B(n31241), .Z(n31243) );
  NAND U32054 ( .A(n31244), .B(n31243), .Z(n31289) );
  XOR U32055 ( .A(n31288), .B(n31289), .Z(n31256) );
  OR U32056 ( .A(n31246), .B(n31245), .Z(n31250) );
  NANDN U32057 ( .A(n31248), .B(n31247), .Z(n31249) );
  NAND U32058 ( .A(n31250), .B(n31249), .Z(n31257) );
  XNOR U32059 ( .A(n31256), .B(n31257), .Z(n31258) );
  XNOR U32060 ( .A(n31259), .B(n31258), .Z(n31292) );
  XNOR U32061 ( .A(n31292), .B(sreg[1776]), .Z(n31294) );
  NAND U32062 ( .A(n31251), .B(sreg[1775]), .Z(n31255) );
  OR U32063 ( .A(n31253), .B(n31252), .Z(n31254) );
  AND U32064 ( .A(n31255), .B(n31254), .Z(n31293) );
  XOR U32065 ( .A(n31294), .B(n31293), .Z(c[1776]) );
  NANDN U32066 ( .A(n31257), .B(n31256), .Z(n31261) );
  NAND U32067 ( .A(n31259), .B(n31258), .Z(n31260) );
  NAND U32068 ( .A(n31261), .B(n31260), .Z(n31300) );
  NAND U32069 ( .A(b[0]), .B(a[761]), .Z(n31262) );
  XNOR U32070 ( .A(b[1]), .B(n31262), .Z(n31264) );
  NAND U32071 ( .A(n123), .B(a[760]), .Z(n31263) );
  AND U32072 ( .A(n31264), .B(n31263), .Z(n31317) );
  XOR U32073 ( .A(a[757]), .B(n42197), .Z(n31306) );
  NANDN U32074 ( .A(n31306), .B(n42173), .Z(n31267) );
  NANDN U32075 ( .A(n31265), .B(n42172), .Z(n31266) );
  NAND U32076 ( .A(n31267), .B(n31266), .Z(n31315) );
  NAND U32077 ( .A(b[7]), .B(a[753]), .Z(n31316) );
  XNOR U32078 ( .A(n31315), .B(n31316), .Z(n31318) );
  XOR U32079 ( .A(n31317), .B(n31318), .Z(n31324) );
  NANDN U32080 ( .A(n31268), .B(n42093), .Z(n31270) );
  XOR U32081 ( .A(n42134), .B(a[759]), .Z(n31309) );
  NANDN U32082 ( .A(n31309), .B(n42095), .Z(n31269) );
  NAND U32083 ( .A(n31270), .B(n31269), .Z(n31322) );
  NANDN U32084 ( .A(n31271), .B(n42231), .Z(n31273) );
  XOR U32085 ( .A(n225), .B(a[755]), .Z(n31312) );
  NANDN U32086 ( .A(n31312), .B(n42234), .Z(n31272) );
  AND U32087 ( .A(n31273), .B(n31272), .Z(n31321) );
  XNOR U32088 ( .A(n31322), .B(n31321), .Z(n31323) );
  XNOR U32089 ( .A(n31324), .B(n31323), .Z(n31328) );
  NANDN U32090 ( .A(n31275), .B(n31274), .Z(n31279) );
  NAND U32091 ( .A(n31277), .B(n31276), .Z(n31278) );
  AND U32092 ( .A(n31279), .B(n31278), .Z(n31327) );
  XOR U32093 ( .A(n31328), .B(n31327), .Z(n31329) );
  NANDN U32094 ( .A(n31281), .B(n31280), .Z(n31285) );
  NANDN U32095 ( .A(n31283), .B(n31282), .Z(n31284) );
  NAND U32096 ( .A(n31285), .B(n31284), .Z(n31330) );
  XOR U32097 ( .A(n31329), .B(n31330), .Z(n31297) );
  OR U32098 ( .A(n31287), .B(n31286), .Z(n31291) );
  NANDN U32099 ( .A(n31289), .B(n31288), .Z(n31290) );
  NAND U32100 ( .A(n31291), .B(n31290), .Z(n31298) );
  XNOR U32101 ( .A(n31297), .B(n31298), .Z(n31299) );
  XNOR U32102 ( .A(n31300), .B(n31299), .Z(n31333) );
  XNOR U32103 ( .A(n31333), .B(sreg[1777]), .Z(n31335) );
  NAND U32104 ( .A(n31292), .B(sreg[1776]), .Z(n31296) );
  OR U32105 ( .A(n31294), .B(n31293), .Z(n31295) );
  AND U32106 ( .A(n31296), .B(n31295), .Z(n31334) );
  XOR U32107 ( .A(n31335), .B(n31334), .Z(c[1777]) );
  NANDN U32108 ( .A(n31298), .B(n31297), .Z(n31302) );
  NAND U32109 ( .A(n31300), .B(n31299), .Z(n31301) );
  NAND U32110 ( .A(n31302), .B(n31301), .Z(n31341) );
  NAND U32111 ( .A(b[0]), .B(a[762]), .Z(n31303) );
  XNOR U32112 ( .A(b[1]), .B(n31303), .Z(n31305) );
  NAND U32113 ( .A(n123), .B(a[761]), .Z(n31304) );
  AND U32114 ( .A(n31305), .B(n31304), .Z(n31358) );
  XOR U32115 ( .A(a[758]), .B(n42197), .Z(n31347) );
  NANDN U32116 ( .A(n31347), .B(n42173), .Z(n31308) );
  NANDN U32117 ( .A(n31306), .B(n42172), .Z(n31307) );
  NAND U32118 ( .A(n31308), .B(n31307), .Z(n31356) );
  NAND U32119 ( .A(b[7]), .B(a[754]), .Z(n31357) );
  XNOR U32120 ( .A(n31356), .B(n31357), .Z(n31359) );
  XOR U32121 ( .A(n31358), .B(n31359), .Z(n31365) );
  NANDN U32122 ( .A(n31309), .B(n42093), .Z(n31311) );
  XOR U32123 ( .A(n42134), .B(a[760]), .Z(n31350) );
  NANDN U32124 ( .A(n31350), .B(n42095), .Z(n31310) );
  NAND U32125 ( .A(n31311), .B(n31310), .Z(n31363) );
  NANDN U32126 ( .A(n31312), .B(n42231), .Z(n31314) );
  XOR U32127 ( .A(n225), .B(a[756]), .Z(n31353) );
  NANDN U32128 ( .A(n31353), .B(n42234), .Z(n31313) );
  AND U32129 ( .A(n31314), .B(n31313), .Z(n31362) );
  XNOR U32130 ( .A(n31363), .B(n31362), .Z(n31364) );
  XNOR U32131 ( .A(n31365), .B(n31364), .Z(n31369) );
  NANDN U32132 ( .A(n31316), .B(n31315), .Z(n31320) );
  NAND U32133 ( .A(n31318), .B(n31317), .Z(n31319) );
  AND U32134 ( .A(n31320), .B(n31319), .Z(n31368) );
  XOR U32135 ( .A(n31369), .B(n31368), .Z(n31370) );
  NANDN U32136 ( .A(n31322), .B(n31321), .Z(n31326) );
  NANDN U32137 ( .A(n31324), .B(n31323), .Z(n31325) );
  NAND U32138 ( .A(n31326), .B(n31325), .Z(n31371) );
  XOR U32139 ( .A(n31370), .B(n31371), .Z(n31338) );
  OR U32140 ( .A(n31328), .B(n31327), .Z(n31332) );
  NANDN U32141 ( .A(n31330), .B(n31329), .Z(n31331) );
  NAND U32142 ( .A(n31332), .B(n31331), .Z(n31339) );
  XNOR U32143 ( .A(n31338), .B(n31339), .Z(n31340) );
  XNOR U32144 ( .A(n31341), .B(n31340), .Z(n31374) );
  XNOR U32145 ( .A(n31374), .B(sreg[1778]), .Z(n31376) );
  NAND U32146 ( .A(n31333), .B(sreg[1777]), .Z(n31337) );
  OR U32147 ( .A(n31335), .B(n31334), .Z(n31336) );
  AND U32148 ( .A(n31337), .B(n31336), .Z(n31375) );
  XOR U32149 ( .A(n31376), .B(n31375), .Z(c[1778]) );
  NANDN U32150 ( .A(n31339), .B(n31338), .Z(n31343) );
  NAND U32151 ( .A(n31341), .B(n31340), .Z(n31342) );
  NAND U32152 ( .A(n31343), .B(n31342), .Z(n31382) );
  NAND U32153 ( .A(b[0]), .B(a[763]), .Z(n31344) );
  XNOR U32154 ( .A(b[1]), .B(n31344), .Z(n31346) );
  NAND U32155 ( .A(n124), .B(a[762]), .Z(n31345) );
  AND U32156 ( .A(n31346), .B(n31345), .Z(n31399) );
  XOR U32157 ( .A(a[759]), .B(n42197), .Z(n31388) );
  NANDN U32158 ( .A(n31388), .B(n42173), .Z(n31349) );
  NANDN U32159 ( .A(n31347), .B(n42172), .Z(n31348) );
  NAND U32160 ( .A(n31349), .B(n31348), .Z(n31397) );
  NAND U32161 ( .A(b[7]), .B(a[755]), .Z(n31398) );
  XNOR U32162 ( .A(n31397), .B(n31398), .Z(n31400) );
  XOR U32163 ( .A(n31399), .B(n31400), .Z(n31406) );
  NANDN U32164 ( .A(n31350), .B(n42093), .Z(n31352) );
  XOR U32165 ( .A(n42134), .B(a[761]), .Z(n31391) );
  NANDN U32166 ( .A(n31391), .B(n42095), .Z(n31351) );
  NAND U32167 ( .A(n31352), .B(n31351), .Z(n31404) );
  NANDN U32168 ( .A(n31353), .B(n42231), .Z(n31355) );
  XOR U32169 ( .A(n225), .B(a[757]), .Z(n31394) );
  NANDN U32170 ( .A(n31394), .B(n42234), .Z(n31354) );
  AND U32171 ( .A(n31355), .B(n31354), .Z(n31403) );
  XNOR U32172 ( .A(n31404), .B(n31403), .Z(n31405) );
  XNOR U32173 ( .A(n31406), .B(n31405), .Z(n31410) );
  NANDN U32174 ( .A(n31357), .B(n31356), .Z(n31361) );
  NAND U32175 ( .A(n31359), .B(n31358), .Z(n31360) );
  AND U32176 ( .A(n31361), .B(n31360), .Z(n31409) );
  XOR U32177 ( .A(n31410), .B(n31409), .Z(n31411) );
  NANDN U32178 ( .A(n31363), .B(n31362), .Z(n31367) );
  NANDN U32179 ( .A(n31365), .B(n31364), .Z(n31366) );
  NAND U32180 ( .A(n31367), .B(n31366), .Z(n31412) );
  XOR U32181 ( .A(n31411), .B(n31412), .Z(n31379) );
  OR U32182 ( .A(n31369), .B(n31368), .Z(n31373) );
  NANDN U32183 ( .A(n31371), .B(n31370), .Z(n31372) );
  NAND U32184 ( .A(n31373), .B(n31372), .Z(n31380) );
  XNOR U32185 ( .A(n31379), .B(n31380), .Z(n31381) );
  XNOR U32186 ( .A(n31382), .B(n31381), .Z(n31415) );
  XNOR U32187 ( .A(n31415), .B(sreg[1779]), .Z(n31417) );
  NAND U32188 ( .A(n31374), .B(sreg[1778]), .Z(n31378) );
  OR U32189 ( .A(n31376), .B(n31375), .Z(n31377) );
  AND U32190 ( .A(n31378), .B(n31377), .Z(n31416) );
  XOR U32191 ( .A(n31417), .B(n31416), .Z(c[1779]) );
  NANDN U32192 ( .A(n31380), .B(n31379), .Z(n31384) );
  NAND U32193 ( .A(n31382), .B(n31381), .Z(n31383) );
  NAND U32194 ( .A(n31384), .B(n31383), .Z(n31423) );
  NAND U32195 ( .A(b[0]), .B(a[764]), .Z(n31385) );
  XNOR U32196 ( .A(b[1]), .B(n31385), .Z(n31387) );
  NAND U32197 ( .A(n124), .B(a[763]), .Z(n31386) );
  AND U32198 ( .A(n31387), .B(n31386), .Z(n31440) );
  XOR U32199 ( .A(a[760]), .B(n42197), .Z(n31429) );
  NANDN U32200 ( .A(n31429), .B(n42173), .Z(n31390) );
  NANDN U32201 ( .A(n31388), .B(n42172), .Z(n31389) );
  NAND U32202 ( .A(n31390), .B(n31389), .Z(n31438) );
  NAND U32203 ( .A(b[7]), .B(a[756]), .Z(n31439) );
  XNOR U32204 ( .A(n31438), .B(n31439), .Z(n31441) );
  XOR U32205 ( .A(n31440), .B(n31441), .Z(n31447) );
  NANDN U32206 ( .A(n31391), .B(n42093), .Z(n31393) );
  XOR U32207 ( .A(n42134), .B(a[762]), .Z(n31432) );
  NANDN U32208 ( .A(n31432), .B(n42095), .Z(n31392) );
  NAND U32209 ( .A(n31393), .B(n31392), .Z(n31445) );
  NANDN U32210 ( .A(n31394), .B(n42231), .Z(n31396) );
  XOR U32211 ( .A(n225), .B(a[758]), .Z(n31435) );
  NANDN U32212 ( .A(n31435), .B(n42234), .Z(n31395) );
  AND U32213 ( .A(n31396), .B(n31395), .Z(n31444) );
  XNOR U32214 ( .A(n31445), .B(n31444), .Z(n31446) );
  XNOR U32215 ( .A(n31447), .B(n31446), .Z(n31451) );
  NANDN U32216 ( .A(n31398), .B(n31397), .Z(n31402) );
  NAND U32217 ( .A(n31400), .B(n31399), .Z(n31401) );
  AND U32218 ( .A(n31402), .B(n31401), .Z(n31450) );
  XOR U32219 ( .A(n31451), .B(n31450), .Z(n31452) );
  NANDN U32220 ( .A(n31404), .B(n31403), .Z(n31408) );
  NANDN U32221 ( .A(n31406), .B(n31405), .Z(n31407) );
  NAND U32222 ( .A(n31408), .B(n31407), .Z(n31453) );
  XOR U32223 ( .A(n31452), .B(n31453), .Z(n31420) );
  OR U32224 ( .A(n31410), .B(n31409), .Z(n31414) );
  NANDN U32225 ( .A(n31412), .B(n31411), .Z(n31413) );
  NAND U32226 ( .A(n31414), .B(n31413), .Z(n31421) );
  XNOR U32227 ( .A(n31420), .B(n31421), .Z(n31422) );
  XNOR U32228 ( .A(n31423), .B(n31422), .Z(n31456) );
  XNOR U32229 ( .A(n31456), .B(sreg[1780]), .Z(n31458) );
  NAND U32230 ( .A(n31415), .B(sreg[1779]), .Z(n31419) );
  OR U32231 ( .A(n31417), .B(n31416), .Z(n31418) );
  AND U32232 ( .A(n31419), .B(n31418), .Z(n31457) );
  XOR U32233 ( .A(n31458), .B(n31457), .Z(c[1780]) );
  NANDN U32234 ( .A(n31421), .B(n31420), .Z(n31425) );
  NAND U32235 ( .A(n31423), .B(n31422), .Z(n31424) );
  NAND U32236 ( .A(n31425), .B(n31424), .Z(n31464) );
  NAND U32237 ( .A(b[0]), .B(a[765]), .Z(n31426) );
  XNOR U32238 ( .A(b[1]), .B(n31426), .Z(n31428) );
  NAND U32239 ( .A(n124), .B(a[764]), .Z(n31427) );
  AND U32240 ( .A(n31428), .B(n31427), .Z(n31481) );
  XOR U32241 ( .A(a[761]), .B(n42197), .Z(n31470) );
  NANDN U32242 ( .A(n31470), .B(n42173), .Z(n31431) );
  NANDN U32243 ( .A(n31429), .B(n42172), .Z(n31430) );
  NAND U32244 ( .A(n31431), .B(n31430), .Z(n31479) );
  NAND U32245 ( .A(b[7]), .B(a[757]), .Z(n31480) );
  XNOR U32246 ( .A(n31479), .B(n31480), .Z(n31482) );
  XOR U32247 ( .A(n31481), .B(n31482), .Z(n31488) );
  NANDN U32248 ( .A(n31432), .B(n42093), .Z(n31434) );
  XOR U32249 ( .A(n42134), .B(a[763]), .Z(n31473) );
  NANDN U32250 ( .A(n31473), .B(n42095), .Z(n31433) );
  NAND U32251 ( .A(n31434), .B(n31433), .Z(n31486) );
  NANDN U32252 ( .A(n31435), .B(n42231), .Z(n31437) );
  XOR U32253 ( .A(n225), .B(a[759]), .Z(n31476) );
  NANDN U32254 ( .A(n31476), .B(n42234), .Z(n31436) );
  AND U32255 ( .A(n31437), .B(n31436), .Z(n31485) );
  XNOR U32256 ( .A(n31486), .B(n31485), .Z(n31487) );
  XNOR U32257 ( .A(n31488), .B(n31487), .Z(n31492) );
  NANDN U32258 ( .A(n31439), .B(n31438), .Z(n31443) );
  NAND U32259 ( .A(n31441), .B(n31440), .Z(n31442) );
  AND U32260 ( .A(n31443), .B(n31442), .Z(n31491) );
  XOR U32261 ( .A(n31492), .B(n31491), .Z(n31493) );
  NANDN U32262 ( .A(n31445), .B(n31444), .Z(n31449) );
  NANDN U32263 ( .A(n31447), .B(n31446), .Z(n31448) );
  NAND U32264 ( .A(n31449), .B(n31448), .Z(n31494) );
  XOR U32265 ( .A(n31493), .B(n31494), .Z(n31461) );
  OR U32266 ( .A(n31451), .B(n31450), .Z(n31455) );
  NANDN U32267 ( .A(n31453), .B(n31452), .Z(n31454) );
  NAND U32268 ( .A(n31455), .B(n31454), .Z(n31462) );
  XNOR U32269 ( .A(n31461), .B(n31462), .Z(n31463) );
  XNOR U32270 ( .A(n31464), .B(n31463), .Z(n31497) );
  XNOR U32271 ( .A(n31497), .B(sreg[1781]), .Z(n31499) );
  NAND U32272 ( .A(n31456), .B(sreg[1780]), .Z(n31460) );
  OR U32273 ( .A(n31458), .B(n31457), .Z(n31459) );
  AND U32274 ( .A(n31460), .B(n31459), .Z(n31498) );
  XOR U32275 ( .A(n31499), .B(n31498), .Z(c[1781]) );
  NANDN U32276 ( .A(n31462), .B(n31461), .Z(n31466) );
  NAND U32277 ( .A(n31464), .B(n31463), .Z(n31465) );
  NAND U32278 ( .A(n31466), .B(n31465), .Z(n31505) );
  NAND U32279 ( .A(b[0]), .B(a[766]), .Z(n31467) );
  XNOR U32280 ( .A(b[1]), .B(n31467), .Z(n31469) );
  NAND U32281 ( .A(n124), .B(a[765]), .Z(n31468) );
  AND U32282 ( .A(n31469), .B(n31468), .Z(n31522) );
  XOR U32283 ( .A(a[762]), .B(n42197), .Z(n31511) );
  NANDN U32284 ( .A(n31511), .B(n42173), .Z(n31472) );
  NANDN U32285 ( .A(n31470), .B(n42172), .Z(n31471) );
  NAND U32286 ( .A(n31472), .B(n31471), .Z(n31520) );
  NAND U32287 ( .A(b[7]), .B(a[758]), .Z(n31521) );
  XNOR U32288 ( .A(n31520), .B(n31521), .Z(n31523) );
  XOR U32289 ( .A(n31522), .B(n31523), .Z(n31529) );
  NANDN U32290 ( .A(n31473), .B(n42093), .Z(n31475) );
  XOR U32291 ( .A(n42134), .B(a[764]), .Z(n31514) );
  NANDN U32292 ( .A(n31514), .B(n42095), .Z(n31474) );
  NAND U32293 ( .A(n31475), .B(n31474), .Z(n31527) );
  NANDN U32294 ( .A(n31476), .B(n42231), .Z(n31478) );
  XOR U32295 ( .A(n225), .B(a[760]), .Z(n31517) );
  NANDN U32296 ( .A(n31517), .B(n42234), .Z(n31477) );
  AND U32297 ( .A(n31478), .B(n31477), .Z(n31526) );
  XNOR U32298 ( .A(n31527), .B(n31526), .Z(n31528) );
  XNOR U32299 ( .A(n31529), .B(n31528), .Z(n31533) );
  NANDN U32300 ( .A(n31480), .B(n31479), .Z(n31484) );
  NAND U32301 ( .A(n31482), .B(n31481), .Z(n31483) );
  AND U32302 ( .A(n31484), .B(n31483), .Z(n31532) );
  XOR U32303 ( .A(n31533), .B(n31532), .Z(n31534) );
  NANDN U32304 ( .A(n31486), .B(n31485), .Z(n31490) );
  NANDN U32305 ( .A(n31488), .B(n31487), .Z(n31489) );
  NAND U32306 ( .A(n31490), .B(n31489), .Z(n31535) );
  XOR U32307 ( .A(n31534), .B(n31535), .Z(n31502) );
  OR U32308 ( .A(n31492), .B(n31491), .Z(n31496) );
  NANDN U32309 ( .A(n31494), .B(n31493), .Z(n31495) );
  NAND U32310 ( .A(n31496), .B(n31495), .Z(n31503) );
  XNOR U32311 ( .A(n31502), .B(n31503), .Z(n31504) );
  XNOR U32312 ( .A(n31505), .B(n31504), .Z(n31538) );
  XNOR U32313 ( .A(n31538), .B(sreg[1782]), .Z(n31540) );
  NAND U32314 ( .A(n31497), .B(sreg[1781]), .Z(n31501) );
  OR U32315 ( .A(n31499), .B(n31498), .Z(n31500) );
  AND U32316 ( .A(n31501), .B(n31500), .Z(n31539) );
  XOR U32317 ( .A(n31540), .B(n31539), .Z(c[1782]) );
  NANDN U32318 ( .A(n31503), .B(n31502), .Z(n31507) );
  NAND U32319 ( .A(n31505), .B(n31504), .Z(n31506) );
  NAND U32320 ( .A(n31507), .B(n31506), .Z(n31546) );
  NAND U32321 ( .A(b[0]), .B(a[767]), .Z(n31508) );
  XNOR U32322 ( .A(b[1]), .B(n31508), .Z(n31510) );
  NAND U32323 ( .A(n124), .B(a[766]), .Z(n31509) );
  AND U32324 ( .A(n31510), .B(n31509), .Z(n31563) );
  XOR U32325 ( .A(a[763]), .B(n42197), .Z(n31552) );
  NANDN U32326 ( .A(n31552), .B(n42173), .Z(n31513) );
  NANDN U32327 ( .A(n31511), .B(n42172), .Z(n31512) );
  NAND U32328 ( .A(n31513), .B(n31512), .Z(n31561) );
  NAND U32329 ( .A(b[7]), .B(a[759]), .Z(n31562) );
  XNOR U32330 ( .A(n31561), .B(n31562), .Z(n31564) );
  XOR U32331 ( .A(n31563), .B(n31564), .Z(n31570) );
  NANDN U32332 ( .A(n31514), .B(n42093), .Z(n31516) );
  XOR U32333 ( .A(n42134), .B(a[765]), .Z(n31555) );
  NANDN U32334 ( .A(n31555), .B(n42095), .Z(n31515) );
  NAND U32335 ( .A(n31516), .B(n31515), .Z(n31568) );
  NANDN U32336 ( .A(n31517), .B(n42231), .Z(n31519) );
  XOR U32337 ( .A(n225), .B(a[761]), .Z(n31558) );
  NANDN U32338 ( .A(n31558), .B(n42234), .Z(n31518) );
  AND U32339 ( .A(n31519), .B(n31518), .Z(n31567) );
  XNOR U32340 ( .A(n31568), .B(n31567), .Z(n31569) );
  XNOR U32341 ( .A(n31570), .B(n31569), .Z(n31574) );
  NANDN U32342 ( .A(n31521), .B(n31520), .Z(n31525) );
  NAND U32343 ( .A(n31523), .B(n31522), .Z(n31524) );
  AND U32344 ( .A(n31525), .B(n31524), .Z(n31573) );
  XOR U32345 ( .A(n31574), .B(n31573), .Z(n31575) );
  NANDN U32346 ( .A(n31527), .B(n31526), .Z(n31531) );
  NANDN U32347 ( .A(n31529), .B(n31528), .Z(n31530) );
  NAND U32348 ( .A(n31531), .B(n31530), .Z(n31576) );
  XOR U32349 ( .A(n31575), .B(n31576), .Z(n31543) );
  OR U32350 ( .A(n31533), .B(n31532), .Z(n31537) );
  NANDN U32351 ( .A(n31535), .B(n31534), .Z(n31536) );
  NAND U32352 ( .A(n31537), .B(n31536), .Z(n31544) );
  XNOR U32353 ( .A(n31543), .B(n31544), .Z(n31545) );
  XNOR U32354 ( .A(n31546), .B(n31545), .Z(n31579) );
  XNOR U32355 ( .A(n31579), .B(sreg[1783]), .Z(n31581) );
  NAND U32356 ( .A(n31538), .B(sreg[1782]), .Z(n31542) );
  OR U32357 ( .A(n31540), .B(n31539), .Z(n31541) );
  AND U32358 ( .A(n31542), .B(n31541), .Z(n31580) );
  XOR U32359 ( .A(n31581), .B(n31580), .Z(c[1783]) );
  NANDN U32360 ( .A(n31544), .B(n31543), .Z(n31548) );
  NAND U32361 ( .A(n31546), .B(n31545), .Z(n31547) );
  NAND U32362 ( .A(n31548), .B(n31547), .Z(n31587) );
  NAND U32363 ( .A(b[0]), .B(a[768]), .Z(n31549) );
  XNOR U32364 ( .A(b[1]), .B(n31549), .Z(n31551) );
  NAND U32365 ( .A(n124), .B(a[767]), .Z(n31550) );
  AND U32366 ( .A(n31551), .B(n31550), .Z(n31604) );
  XOR U32367 ( .A(a[764]), .B(n42197), .Z(n31593) );
  NANDN U32368 ( .A(n31593), .B(n42173), .Z(n31554) );
  NANDN U32369 ( .A(n31552), .B(n42172), .Z(n31553) );
  NAND U32370 ( .A(n31554), .B(n31553), .Z(n31602) );
  NAND U32371 ( .A(b[7]), .B(a[760]), .Z(n31603) );
  XNOR U32372 ( .A(n31602), .B(n31603), .Z(n31605) );
  XOR U32373 ( .A(n31604), .B(n31605), .Z(n31611) );
  NANDN U32374 ( .A(n31555), .B(n42093), .Z(n31557) );
  XOR U32375 ( .A(n42134), .B(a[766]), .Z(n31596) );
  NANDN U32376 ( .A(n31596), .B(n42095), .Z(n31556) );
  NAND U32377 ( .A(n31557), .B(n31556), .Z(n31609) );
  NANDN U32378 ( .A(n31558), .B(n42231), .Z(n31560) );
  XOR U32379 ( .A(n225), .B(a[762]), .Z(n31599) );
  NANDN U32380 ( .A(n31599), .B(n42234), .Z(n31559) );
  AND U32381 ( .A(n31560), .B(n31559), .Z(n31608) );
  XNOR U32382 ( .A(n31609), .B(n31608), .Z(n31610) );
  XNOR U32383 ( .A(n31611), .B(n31610), .Z(n31615) );
  NANDN U32384 ( .A(n31562), .B(n31561), .Z(n31566) );
  NAND U32385 ( .A(n31564), .B(n31563), .Z(n31565) );
  AND U32386 ( .A(n31566), .B(n31565), .Z(n31614) );
  XOR U32387 ( .A(n31615), .B(n31614), .Z(n31616) );
  NANDN U32388 ( .A(n31568), .B(n31567), .Z(n31572) );
  NANDN U32389 ( .A(n31570), .B(n31569), .Z(n31571) );
  NAND U32390 ( .A(n31572), .B(n31571), .Z(n31617) );
  XOR U32391 ( .A(n31616), .B(n31617), .Z(n31584) );
  OR U32392 ( .A(n31574), .B(n31573), .Z(n31578) );
  NANDN U32393 ( .A(n31576), .B(n31575), .Z(n31577) );
  NAND U32394 ( .A(n31578), .B(n31577), .Z(n31585) );
  XNOR U32395 ( .A(n31584), .B(n31585), .Z(n31586) );
  XNOR U32396 ( .A(n31587), .B(n31586), .Z(n31620) );
  XNOR U32397 ( .A(n31620), .B(sreg[1784]), .Z(n31622) );
  NAND U32398 ( .A(n31579), .B(sreg[1783]), .Z(n31583) );
  OR U32399 ( .A(n31581), .B(n31580), .Z(n31582) );
  AND U32400 ( .A(n31583), .B(n31582), .Z(n31621) );
  XOR U32401 ( .A(n31622), .B(n31621), .Z(c[1784]) );
  NANDN U32402 ( .A(n31585), .B(n31584), .Z(n31589) );
  NAND U32403 ( .A(n31587), .B(n31586), .Z(n31588) );
  NAND U32404 ( .A(n31589), .B(n31588), .Z(n31628) );
  NAND U32405 ( .A(b[0]), .B(a[769]), .Z(n31590) );
  XNOR U32406 ( .A(b[1]), .B(n31590), .Z(n31592) );
  NAND U32407 ( .A(n124), .B(a[768]), .Z(n31591) );
  AND U32408 ( .A(n31592), .B(n31591), .Z(n31645) );
  XOR U32409 ( .A(a[765]), .B(n42197), .Z(n31634) );
  NANDN U32410 ( .A(n31634), .B(n42173), .Z(n31595) );
  NANDN U32411 ( .A(n31593), .B(n42172), .Z(n31594) );
  NAND U32412 ( .A(n31595), .B(n31594), .Z(n31643) );
  NAND U32413 ( .A(b[7]), .B(a[761]), .Z(n31644) );
  XNOR U32414 ( .A(n31643), .B(n31644), .Z(n31646) );
  XOR U32415 ( .A(n31645), .B(n31646), .Z(n31652) );
  NANDN U32416 ( .A(n31596), .B(n42093), .Z(n31598) );
  XOR U32417 ( .A(n42134), .B(a[767]), .Z(n31637) );
  NANDN U32418 ( .A(n31637), .B(n42095), .Z(n31597) );
  NAND U32419 ( .A(n31598), .B(n31597), .Z(n31650) );
  NANDN U32420 ( .A(n31599), .B(n42231), .Z(n31601) );
  XOR U32421 ( .A(n225), .B(a[763]), .Z(n31640) );
  NANDN U32422 ( .A(n31640), .B(n42234), .Z(n31600) );
  AND U32423 ( .A(n31601), .B(n31600), .Z(n31649) );
  XNOR U32424 ( .A(n31650), .B(n31649), .Z(n31651) );
  XNOR U32425 ( .A(n31652), .B(n31651), .Z(n31656) );
  NANDN U32426 ( .A(n31603), .B(n31602), .Z(n31607) );
  NAND U32427 ( .A(n31605), .B(n31604), .Z(n31606) );
  AND U32428 ( .A(n31607), .B(n31606), .Z(n31655) );
  XOR U32429 ( .A(n31656), .B(n31655), .Z(n31657) );
  NANDN U32430 ( .A(n31609), .B(n31608), .Z(n31613) );
  NANDN U32431 ( .A(n31611), .B(n31610), .Z(n31612) );
  NAND U32432 ( .A(n31613), .B(n31612), .Z(n31658) );
  XOR U32433 ( .A(n31657), .B(n31658), .Z(n31625) );
  OR U32434 ( .A(n31615), .B(n31614), .Z(n31619) );
  NANDN U32435 ( .A(n31617), .B(n31616), .Z(n31618) );
  NAND U32436 ( .A(n31619), .B(n31618), .Z(n31626) );
  XNOR U32437 ( .A(n31625), .B(n31626), .Z(n31627) );
  XNOR U32438 ( .A(n31628), .B(n31627), .Z(n31661) );
  XNOR U32439 ( .A(n31661), .B(sreg[1785]), .Z(n31663) );
  NAND U32440 ( .A(n31620), .B(sreg[1784]), .Z(n31624) );
  OR U32441 ( .A(n31622), .B(n31621), .Z(n31623) );
  AND U32442 ( .A(n31624), .B(n31623), .Z(n31662) );
  XOR U32443 ( .A(n31663), .B(n31662), .Z(c[1785]) );
  NANDN U32444 ( .A(n31626), .B(n31625), .Z(n31630) );
  NAND U32445 ( .A(n31628), .B(n31627), .Z(n31629) );
  NAND U32446 ( .A(n31630), .B(n31629), .Z(n31669) );
  NAND U32447 ( .A(b[0]), .B(a[770]), .Z(n31631) );
  XNOR U32448 ( .A(b[1]), .B(n31631), .Z(n31633) );
  NAND U32449 ( .A(n125), .B(a[769]), .Z(n31632) );
  AND U32450 ( .A(n31633), .B(n31632), .Z(n31686) );
  XOR U32451 ( .A(a[766]), .B(n42197), .Z(n31675) );
  NANDN U32452 ( .A(n31675), .B(n42173), .Z(n31636) );
  NANDN U32453 ( .A(n31634), .B(n42172), .Z(n31635) );
  NAND U32454 ( .A(n31636), .B(n31635), .Z(n31684) );
  NAND U32455 ( .A(b[7]), .B(a[762]), .Z(n31685) );
  XNOR U32456 ( .A(n31684), .B(n31685), .Z(n31687) );
  XOR U32457 ( .A(n31686), .B(n31687), .Z(n31693) );
  NANDN U32458 ( .A(n31637), .B(n42093), .Z(n31639) );
  XOR U32459 ( .A(n42134), .B(a[768]), .Z(n31678) );
  NANDN U32460 ( .A(n31678), .B(n42095), .Z(n31638) );
  NAND U32461 ( .A(n31639), .B(n31638), .Z(n31691) );
  NANDN U32462 ( .A(n31640), .B(n42231), .Z(n31642) );
  XOR U32463 ( .A(n225), .B(a[764]), .Z(n31681) );
  NANDN U32464 ( .A(n31681), .B(n42234), .Z(n31641) );
  AND U32465 ( .A(n31642), .B(n31641), .Z(n31690) );
  XNOR U32466 ( .A(n31691), .B(n31690), .Z(n31692) );
  XNOR U32467 ( .A(n31693), .B(n31692), .Z(n31697) );
  NANDN U32468 ( .A(n31644), .B(n31643), .Z(n31648) );
  NAND U32469 ( .A(n31646), .B(n31645), .Z(n31647) );
  AND U32470 ( .A(n31648), .B(n31647), .Z(n31696) );
  XOR U32471 ( .A(n31697), .B(n31696), .Z(n31698) );
  NANDN U32472 ( .A(n31650), .B(n31649), .Z(n31654) );
  NANDN U32473 ( .A(n31652), .B(n31651), .Z(n31653) );
  NAND U32474 ( .A(n31654), .B(n31653), .Z(n31699) );
  XOR U32475 ( .A(n31698), .B(n31699), .Z(n31666) );
  OR U32476 ( .A(n31656), .B(n31655), .Z(n31660) );
  NANDN U32477 ( .A(n31658), .B(n31657), .Z(n31659) );
  NAND U32478 ( .A(n31660), .B(n31659), .Z(n31667) );
  XNOR U32479 ( .A(n31666), .B(n31667), .Z(n31668) );
  XNOR U32480 ( .A(n31669), .B(n31668), .Z(n31702) );
  XNOR U32481 ( .A(n31702), .B(sreg[1786]), .Z(n31704) );
  NAND U32482 ( .A(n31661), .B(sreg[1785]), .Z(n31665) );
  OR U32483 ( .A(n31663), .B(n31662), .Z(n31664) );
  AND U32484 ( .A(n31665), .B(n31664), .Z(n31703) );
  XOR U32485 ( .A(n31704), .B(n31703), .Z(c[1786]) );
  NANDN U32486 ( .A(n31667), .B(n31666), .Z(n31671) );
  NAND U32487 ( .A(n31669), .B(n31668), .Z(n31670) );
  NAND U32488 ( .A(n31671), .B(n31670), .Z(n31710) );
  NAND U32489 ( .A(b[0]), .B(a[771]), .Z(n31672) );
  XNOR U32490 ( .A(b[1]), .B(n31672), .Z(n31674) );
  NAND U32491 ( .A(n125), .B(a[770]), .Z(n31673) );
  AND U32492 ( .A(n31674), .B(n31673), .Z(n31727) );
  XOR U32493 ( .A(a[767]), .B(n42197), .Z(n31716) );
  NANDN U32494 ( .A(n31716), .B(n42173), .Z(n31677) );
  NANDN U32495 ( .A(n31675), .B(n42172), .Z(n31676) );
  NAND U32496 ( .A(n31677), .B(n31676), .Z(n31725) );
  NAND U32497 ( .A(b[7]), .B(a[763]), .Z(n31726) );
  XNOR U32498 ( .A(n31725), .B(n31726), .Z(n31728) );
  XOR U32499 ( .A(n31727), .B(n31728), .Z(n31734) );
  NANDN U32500 ( .A(n31678), .B(n42093), .Z(n31680) );
  XOR U32501 ( .A(n42134), .B(a[769]), .Z(n31719) );
  NANDN U32502 ( .A(n31719), .B(n42095), .Z(n31679) );
  NAND U32503 ( .A(n31680), .B(n31679), .Z(n31732) );
  NANDN U32504 ( .A(n31681), .B(n42231), .Z(n31683) );
  XOR U32505 ( .A(n225), .B(a[765]), .Z(n31722) );
  NANDN U32506 ( .A(n31722), .B(n42234), .Z(n31682) );
  AND U32507 ( .A(n31683), .B(n31682), .Z(n31731) );
  XNOR U32508 ( .A(n31732), .B(n31731), .Z(n31733) );
  XNOR U32509 ( .A(n31734), .B(n31733), .Z(n31738) );
  NANDN U32510 ( .A(n31685), .B(n31684), .Z(n31689) );
  NAND U32511 ( .A(n31687), .B(n31686), .Z(n31688) );
  AND U32512 ( .A(n31689), .B(n31688), .Z(n31737) );
  XOR U32513 ( .A(n31738), .B(n31737), .Z(n31739) );
  NANDN U32514 ( .A(n31691), .B(n31690), .Z(n31695) );
  NANDN U32515 ( .A(n31693), .B(n31692), .Z(n31694) );
  NAND U32516 ( .A(n31695), .B(n31694), .Z(n31740) );
  XOR U32517 ( .A(n31739), .B(n31740), .Z(n31707) );
  OR U32518 ( .A(n31697), .B(n31696), .Z(n31701) );
  NANDN U32519 ( .A(n31699), .B(n31698), .Z(n31700) );
  NAND U32520 ( .A(n31701), .B(n31700), .Z(n31708) );
  XNOR U32521 ( .A(n31707), .B(n31708), .Z(n31709) );
  XNOR U32522 ( .A(n31710), .B(n31709), .Z(n31743) );
  XNOR U32523 ( .A(n31743), .B(sreg[1787]), .Z(n31745) );
  NAND U32524 ( .A(n31702), .B(sreg[1786]), .Z(n31706) );
  OR U32525 ( .A(n31704), .B(n31703), .Z(n31705) );
  AND U32526 ( .A(n31706), .B(n31705), .Z(n31744) );
  XOR U32527 ( .A(n31745), .B(n31744), .Z(c[1787]) );
  NANDN U32528 ( .A(n31708), .B(n31707), .Z(n31712) );
  NAND U32529 ( .A(n31710), .B(n31709), .Z(n31711) );
  NAND U32530 ( .A(n31712), .B(n31711), .Z(n31751) );
  NAND U32531 ( .A(b[0]), .B(a[772]), .Z(n31713) );
  XNOR U32532 ( .A(b[1]), .B(n31713), .Z(n31715) );
  NAND U32533 ( .A(n125), .B(a[771]), .Z(n31714) );
  AND U32534 ( .A(n31715), .B(n31714), .Z(n31768) );
  XOR U32535 ( .A(a[768]), .B(n42197), .Z(n31757) );
  NANDN U32536 ( .A(n31757), .B(n42173), .Z(n31718) );
  NANDN U32537 ( .A(n31716), .B(n42172), .Z(n31717) );
  NAND U32538 ( .A(n31718), .B(n31717), .Z(n31766) );
  NAND U32539 ( .A(b[7]), .B(a[764]), .Z(n31767) );
  XNOR U32540 ( .A(n31766), .B(n31767), .Z(n31769) );
  XOR U32541 ( .A(n31768), .B(n31769), .Z(n31775) );
  NANDN U32542 ( .A(n31719), .B(n42093), .Z(n31721) );
  XOR U32543 ( .A(n42134), .B(a[770]), .Z(n31760) );
  NANDN U32544 ( .A(n31760), .B(n42095), .Z(n31720) );
  NAND U32545 ( .A(n31721), .B(n31720), .Z(n31773) );
  NANDN U32546 ( .A(n31722), .B(n42231), .Z(n31724) );
  XOR U32547 ( .A(n225), .B(a[766]), .Z(n31763) );
  NANDN U32548 ( .A(n31763), .B(n42234), .Z(n31723) );
  AND U32549 ( .A(n31724), .B(n31723), .Z(n31772) );
  XNOR U32550 ( .A(n31773), .B(n31772), .Z(n31774) );
  XNOR U32551 ( .A(n31775), .B(n31774), .Z(n31779) );
  NANDN U32552 ( .A(n31726), .B(n31725), .Z(n31730) );
  NAND U32553 ( .A(n31728), .B(n31727), .Z(n31729) );
  AND U32554 ( .A(n31730), .B(n31729), .Z(n31778) );
  XOR U32555 ( .A(n31779), .B(n31778), .Z(n31780) );
  NANDN U32556 ( .A(n31732), .B(n31731), .Z(n31736) );
  NANDN U32557 ( .A(n31734), .B(n31733), .Z(n31735) );
  NAND U32558 ( .A(n31736), .B(n31735), .Z(n31781) );
  XOR U32559 ( .A(n31780), .B(n31781), .Z(n31748) );
  OR U32560 ( .A(n31738), .B(n31737), .Z(n31742) );
  NANDN U32561 ( .A(n31740), .B(n31739), .Z(n31741) );
  NAND U32562 ( .A(n31742), .B(n31741), .Z(n31749) );
  XNOR U32563 ( .A(n31748), .B(n31749), .Z(n31750) );
  XNOR U32564 ( .A(n31751), .B(n31750), .Z(n31784) );
  XNOR U32565 ( .A(n31784), .B(sreg[1788]), .Z(n31786) );
  NAND U32566 ( .A(n31743), .B(sreg[1787]), .Z(n31747) );
  OR U32567 ( .A(n31745), .B(n31744), .Z(n31746) );
  AND U32568 ( .A(n31747), .B(n31746), .Z(n31785) );
  XOR U32569 ( .A(n31786), .B(n31785), .Z(c[1788]) );
  NANDN U32570 ( .A(n31749), .B(n31748), .Z(n31753) );
  NAND U32571 ( .A(n31751), .B(n31750), .Z(n31752) );
  NAND U32572 ( .A(n31753), .B(n31752), .Z(n31792) );
  NAND U32573 ( .A(b[0]), .B(a[773]), .Z(n31754) );
  XNOR U32574 ( .A(b[1]), .B(n31754), .Z(n31756) );
  NAND U32575 ( .A(n125), .B(a[772]), .Z(n31755) );
  AND U32576 ( .A(n31756), .B(n31755), .Z(n31809) );
  XOR U32577 ( .A(a[769]), .B(n42197), .Z(n31798) );
  NANDN U32578 ( .A(n31798), .B(n42173), .Z(n31759) );
  NANDN U32579 ( .A(n31757), .B(n42172), .Z(n31758) );
  NAND U32580 ( .A(n31759), .B(n31758), .Z(n31807) );
  NAND U32581 ( .A(b[7]), .B(a[765]), .Z(n31808) );
  XNOR U32582 ( .A(n31807), .B(n31808), .Z(n31810) );
  XOR U32583 ( .A(n31809), .B(n31810), .Z(n31816) );
  NANDN U32584 ( .A(n31760), .B(n42093), .Z(n31762) );
  XOR U32585 ( .A(n42134), .B(a[771]), .Z(n31801) );
  NANDN U32586 ( .A(n31801), .B(n42095), .Z(n31761) );
  NAND U32587 ( .A(n31762), .B(n31761), .Z(n31814) );
  NANDN U32588 ( .A(n31763), .B(n42231), .Z(n31765) );
  XOR U32589 ( .A(n226), .B(a[767]), .Z(n31804) );
  NANDN U32590 ( .A(n31804), .B(n42234), .Z(n31764) );
  AND U32591 ( .A(n31765), .B(n31764), .Z(n31813) );
  XNOR U32592 ( .A(n31814), .B(n31813), .Z(n31815) );
  XNOR U32593 ( .A(n31816), .B(n31815), .Z(n31820) );
  NANDN U32594 ( .A(n31767), .B(n31766), .Z(n31771) );
  NAND U32595 ( .A(n31769), .B(n31768), .Z(n31770) );
  AND U32596 ( .A(n31771), .B(n31770), .Z(n31819) );
  XOR U32597 ( .A(n31820), .B(n31819), .Z(n31821) );
  NANDN U32598 ( .A(n31773), .B(n31772), .Z(n31777) );
  NANDN U32599 ( .A(n31775), .B(n31774), .Z(n31776) );
  NAND U32600 ( .A(n31777), .B(n31776), .Z(n31822) );
  XOR U32601 ( .A(n31821), .B(n31822), .Z(n31789) );
  OR U32602 ( .A(n31779), .B(n31778), .Z(n31783) );
  NANDN U32603 ( .A(n31781), .B(n31780), .Z(n31782) );
  NAND U32604 ( .A(n31783), .B(n31782), .Z(n31790) );
  XNOR U32605 ( .A(n31789), .B(n31790), .Z(n31791) );
  XNOR U32606 ( .A(n31792), .B(n31791), .Z(n31825) );
  XNOR U32607 ( .A(n31825), .B(sreg[1789]), .Z(n31827) );
  NAND U32608 ( .A(n31784), .B(sreg[1788]), .Z(n31788) );
  OR U32609 ( .A(n31786), .B(n31785), .Z(n31787) );
  AND U32610 ( .A(n31788), .B(n31787), .Z(n31826) );
  XOR U32611 ( .A(n31827), .B(n31826), .Z(c[1789]) );
  NANDN U32612 ( .A(n31790), .B(n31789), .Z(n31794) );
  NAND U32613 ( .A(n31792), .B(n31791), .Z(n31793) );
  NAND U32614 ( .A(n31794), .B(n31793), .Z(n31833) );
  NAND U32615 ( .A(b[0]), .B(a[774]), .Z(n31795) );
  XNOR U32616 ( .A(b[1]), .B(n31795), .Z(n31797) );
  NAND U32617 ( .A(n125), .B(a[773]), .Z(n31796) );
  AND U32618 ( .A(n31797), .B(n31796), .Z(n31850) );
  XOR U32619 ( .A(a[770]), .B(n42197), .Z(n31839) );
  NANDN U32620 ( .A(n31839), .B(n42173), .Z(n31800) );
  NANDN U32621 ( .A(n31798), .B(n42172), .Z(n31799) );
  NAND U32622 ( .A(n31800), .B(n31799), .Z(n31848) );
  NAND U32623 ( .A(b[7]), .B(a[766]), .Z(n31849) );
  XNOR U32624 ( .A(n31848), .B(n31849), .Z(n31851) );
  XOR U32625 ( .A(n31850), .B(n31851), .Z(n31857) );
  NANDN U32626 ( .A(n31801), .B(n42093), .Z(n31803) );
  XOR U32627 ( .A(n42134), .B(a[772]), .Z(n31842) );
  NANDN U32628 ( .A(n31842), .B(n42095), .Z(n31802) );
  NAND U32629 ( .A(n31803), .B(n31802), .Z(n31855) );
  NANDN U32630 ( .A(n31804), .B(n42231), .Z(n31806) );
  XOR U32631 ( .A(n226), .B(a[768]), .Z(n31845) );
  NANDN U32632 ( .A(n31845), .B(n42234), .Z(n31805) );
  AND U32633 ( .A(n31806), .B(n31805), .Z(n31854) );
  XNOR U32634 ( .A(n31855), .B(n31854), .Z(n31856) );
  XNOR U32635 ( .A(n31857), .B(n31856), .Z(n31861) );
  NANDN U32636 ( .A(n31808), .B(n31807), .Z(n31812) );
  NAND U32637 ( .A(n31810), .B(n31809), .Z(n31811) );
  AND U32638 ( .A(n31812), .B(n31811), .Z(n31860) );
  XOR U32639 ( .A(n31861), .B(n31860), .Z(n31862) );
  NANDN U32640 ( .A(n31814), .B(n31813), .Z(n31818) );
  NANDN U32641 ( .A(n31816), .B(n31815), .Z(n31817) );
  NAND U32642 ( .A(n31818), .B(n31817), .Z(n31863) );
  XOR U32643 ( .A(n31862), .B(n31863), .Z(n31830) );
  OR U32644 ( .A(n31820), .B(n31819), .Z(n31824) );
  NANDN U32645 ( .A(n31822), .B(n31821), .Z(n31823) );
  NAND U32646 ( .A(n31824), .B(n31823), .Z(n31831) );
  XNOR U32647 ( .A(n31830), .B(n31831), .Z(n31832) );
  XNOR U32648 ( .A(n31833), .B(n31832), .Z(n31866) );
  XNOR U32649 ( .A(n31866), .B(sreg[1790]), .Z(n31868) );
  NAND U32650 ( .A(n31825), .B(sreg[1789]), .Z(n31829) );
  OR U32651 ( .A(n31827), .B(n31826), .Z(n31828) );
  AND U32652 ( .A(n31829), .B(n31828), .Z(n31867) );
  XOR U32653 ( .A(n31868), .B(n31867), .Z(c[1790]) );
  NANDN U32654 ( .A(n31831), .B(n31830), .Z(n31835) );
  NAND U32655 ( .A(n31833), .B(n31832), .Z(n31834) );
  NAND U32656 ( .A(n31835), .B(n31834), .Z(n31874) );
  NAND U32657 ( .A(b[0]), .B(a[775]), .Z(n31836) );
  XNOR U32658 ( .A(b[1]), .B(n31836), .Z(n31838) );
  NAND U32659 ( .A(n125), .B(a[774]), .Z(n31837) );
  AND U32660 ( .A(n31838), .B(n31837), .Z(n31891) );
  XOR U32661 ( .A(a[771]), .B(n42197), .Z(n31880) );
  NANDN U32662 ( .A(n31880), .B(n42173), .Z(n31841) );
  NANDN U32663 ( .A(n31839), .B(n42172), .Z(n31840) );
  NAND U32664 ( .A(n31841), .B(n31840), .Z(n31889) );
  NAND U32665 ( .A(b[7]), .B(a[767]), .Z(n31890) );
  XNOR U32666 ( .A(n31889), .B(n31890), .Z(n31892) );
  XOR U32667 ( .A(n31891), .B(n31892), .Z(n31898) );
  NANDN U32668 ( .A(n31842), .B(n42093), .Z(n31844) );
  XOR U32669 ( .A(n42134), .B(a[773]), .Z(n31883) );
  NANDN U32670 ( .A(n31883), .B(n42095), .Z(n31843) );
  NAND U32671 ( .A(n31844), .B(n31843), .Z(n31896) );
  NANDN U32672 ( .A(n31845), .B(n42231), .Z(n31847) );
  XOR U32673 ( .A(n226), .B(a[769]), .Z(n31886) );
  NANDN U32674 ( .A(n31886), .B(n42234), .Z(n31846) );
  AND U32675 ( .A(n31847), .B(n31846), .Z(n31895) );
  XNOR U32676 ( .A(n31896), .B(n31895), .Z(n31897) );
  XNOR U32677 ( .A(n31898), .B(n31897), .Z(n31902) );
  NANDN U32678 ( .A(n31849), .B(n31848), .Z(n31853) );
  NAND U32679 ( .A(n31851), .B(n31850), .Z(n31852) );
  AND U32680 ( .A(n31853), .B(n31852), .Z(n31901) );
  XOR U32681 ( .A(n31902), .B(n31901), .Z(n31903) );
  NANDN U32682 ( .A(n31855), .B(n31854), .Z(n31859) );
  NANDN U32683 ( .A(n31857), .B(n31856), .Z(n31858) );
  NAND U32684 ( .A(n31859), .B(n31858), .Z(n31904) );
  XOR U32685 ( .A(n31903), .B(n31904), .Z(n31871) );
  OR U32686 ( .A(n31861), .B(n31860), .Z(n31865) );
  NANDN U32687 ( .A(n31863), .B(n31862), .Z(n31864) );
  NAND U32688 ( .A(n31865), .B(n31864), .Z(n31872) );
  XNOR U32689 ( .A(n31871), .B(n31872), .Z(n31873) );
  XNOR U32690 ( .A(n31874), .B(n31873), .Z(n31907) );
  XNOR U32691 ( .A(n31907), .B(sreg[1791]), .Z(n31909) );
  NAND U32692 ( .A(n31866), .B(sreg[1790]), .Z(n31870) );
  OR U32693 ( .A(n31868), .B(n31867), .Z(n31869) );
  AND U32694 ( .A(n31870), .B(n31869), .Z(n31908) );
  XOR U32695 ( .A(n31909), .B(n31908), .Z(c[1791]) );
  NANDN U32696 ( .A(n31872), .B(n31871), .Z(n31876) );
  NAND U32697 ( .A(n31874), .B(n31873), .Z(n31875) );
  NAND U32698 ( .A(n31876), .B(n31875), .Z(n31915) );
  NAND U32699 ( .A(b[0]), .B(a[776]), .Z(n31877) );
  XNOR U32700 ( .A(b[1]), .B(n31877), .Z(n31879) );
  NAND U32701 ( .A(n125), .B(a[775]), .Z(n31878) );
  AND U32702 ( .A(n31879), .B(n31878), .Z(n31932) );
  XOR U32703 ( .A(a[772]), .B(n42197), .Z(n31921) );
  NANDN U32704 ( .A(n31921), .B(n42173), .Z(n31882) );
  NANDN U32705 ( .A(n31880), .B(n42172), .Z(n31881) );
  NAND U32706 ( .A(n31882), .B(n31881), .Z(n31930) );
  NAND U32707 ( .A(b[7]), .B(a[768]), .Z(n31931) );
  XNOR U32708 ( .A(n31930), .B(n31931), .Z(n31933) );
  XOR U32709 ( .A(n31932), .B(n31933), .Z(n31939) );
  NANDN U32710 ( .A(n31883), .B(n42093), .Z(n31885) );
  XOR U32711 ( .A(n42134), .B(a[774]), .Z(n31924) );
  NANDN U32712 ( .A(n31924), .B(n42095), .Z(n31884) );
  NAND U32713 ( .A(n31885), .B(n31884), .Z(n31937) );
  NANDN U32714 ( .A(n31886), .B(n42231), .Z(n31888) );
  XOR U32715 ( .A(n226), .B(a[770]), .Z(n31927) );
  NANDN U32716 ( .A(n31927), .B(n42234), .Z(n31887) );
  AND U32717 ( .A(n31888), .B(n31887), .Z(n31936) );
  XNOR U32718 ( .A(n31937), .B(n31936), .Z(n31938) );
  XNOR U32719 ( .A(n31939), .B(n31938), .Z(n31943) );
  NANDN U32720 ( .A(n31890), .B(n31889), .Z(n31894) );
  NAND U32721 ( .A(n31892), .B(n31891), .Z(n31893) );
  AND U32722 ( .A(n31894), .B(n31893), .Z(n31942) );
  XOR U32723 ( .A(n31943), .B(n31942), .Z(n31944) );
  NANDN U32724 ( .A(n31896), .B(n31895), .Z(n31900) );
  NANDN U32725 ( .A(n31898), .B(n31897), .Z(n31899) );
  NAND U32726 ( .A(n31900), .B(n31899), .Z(n31945) );
  XOR U32727 ( .A(n31944), .B(n31945), .Z(n31912) );
  OR U32728 ( .A(n31902), .B(n31901), .Z(n31906) );
  NANDN U32729 ( .A(n31904), .B(n31903), .Z(n31905) );
  NAND U32730 ( .A(n31906), .B(n31905), .Z(n31913) );
  XNOR U32731 ( .A(n31912), .B(n31913), .Z(n31914) );
  XNOR U32732 ( .A(n31915), .B(n31914), .Z(n31948) );
  XNOR U32733 ( .A(n31948), .B(sreg[1792]), .Z(n31950) );
  NAND U32734 ( .A(n31907), .B(sreg[1791]), .Z(n31911) );
  OR U32735 ( .A(n31909), .B(n31908), .Z(n31910) );
  AND U32736 ( .A(n31911), .B(n31910), .Z(n31949) );
  XOR U32737 ( .A(n31950), .B(n31949), .Z(c[1792]) );
  NANDN U32738 ( .A(n31913), .B(n31912), .Z(n31917) );
  NAND U32739 ( .A(n31915), .B(n31914), .Z(n31916) );
  NAND U32740 ( .A(n31917), .B(n31916), .Z(n31956) );
  NAND U32741 ( .A(b[0]), .B(a[777]), .Z(n31918) );
  XNOR U32742 ( .A(b[1]), .B(n31918), .Z(n31920) );
  NAND U32743 ( .A(n126), .B(a[776]), .Z(n31919) );
  AND U32744 ( .A(n31920), .B(n31919), .Z(n31973) );
  XOR U32745 ( .A(a[773]), .B(n42197), .Z(n31962) );
  NANDN U32746 ( .A(n31962), .B(n42173), .Z(n31923) );
  NANDN U32747 ( .A(n31921), .B(n42172), .Z(n31922) );
  NAND U32748 ( .A(n31923), .B(n31922), .Z(n31971) );
  NAND U32749 ( .A(b[7]), .B(a[769]), .Z(n31972) );
  XNOR U32750 ( .A(n31971), .B(n31972), .Z(n31974) );
  XOR U32751 ( .A(n31973), .B(n31974), .Z(n31980) );
  NANDN U32752 ( .A(n31924), .B(n42093), .Z(n31926) );
  XOR U32753 ( .A(n42134), .B(a[775]), .Z(n31965) );
  NANDN U32754 ( .A(n31965), .B(n42095), .Z(n31925) );
  NAND U32755 ( .A(n31926), .B(n31925), .Z(n31978) );
  NANDN U32756 ( .A(n31927), .B(n42231), .Z(n31929) );
  XOR U32757 ( .A(n226), .B(a[771]), .Z(n31968) );
  NANDN U32758 ( .A(n31968), .B(n42234), .Z(n31928) );
  AND U32759 ( .A(n31929), .B(n31928), .Z(n31977) );
  XNOR U32760 ( .A(n31978), .B(n31977), .Z(n31979) );
  XNOR U32761 ( .A(n31980), .B(n31979), .Z(n31984) );
  NANDN U32762 ( .A(n31931), .B(n31930), .Z(n31935) );
  NAND U32763 ( .A(n31933), .B(n31932), .Z(n31934) );
  AND U32764 ( .A(n31935), .B(n31934), .Z(n31983) );
  XOR U32765 ( .A(n31984), .B(n31983), .Z(n31985) );
  NANDN U32766 ( .A(n31937), .B(n31936), .Z(n31941) );
  NANDN U32767 ( .A(n31939), .B(n31938), .Z(n31940) );
  NAND U32768 ( .A(n31941), .B(n31940), .Z(n31986) );
  XOR U32769 ( .A(n31985), .B(n31986), .Z(n31953) );
  OR U32770 ( .A(n31943), .B(n31942), .Z(n31947) );
  NANDN U32771 ( .A(n31945), .B(n31944), .Z(n31946) );
  NAND U32772 ( .A(n31947), .B(n31946), .Z(n31954) );
  XNOR U32773 ( .A(n31953), .B(n31954), .Z(n31955) );
  XNOR U32774 ( .A(n31956), .B(n31955), .Z(n31989) );
  XNOR U32775 ( .A(n31989), .B(sreg[1793]), .Z(n31991) );
  NAND U32776 ( .A(n31948), .B(sreg[1792]), .Z(n31952) );
  OR U32777 ( .A(n31950), .B(n31949), .Z(n31951) );
  AND U32778 ( .A(n31952), .B(n31951), .Z(n31990) );
  XOR U32779 ( .A(n31991), .B(n31990), .Z(c[1793]) );
  NANDN U32780 ( .A(n31954), .B(n31953), .Z(n31958) );
  NAND U32781 ( .A(n31956), .B(n31955), .Z(n31957) );
  NAND U32782 ( .A(n31958), .B(n31957), .Z(n31997) );
  NAND U32783 ( .A(b[0]), .B(a[778]), .Z(n31959) );
  XNOR U32784 ( .A(b[1]), .B(n31959), .Z(n31961) );
  NAND U32785 ( .A(n126), .B(a[777]), .Z(n31960) );
  AND U32786 ( .A(n31961), .B(n31960), .Z(n32014) );
  XOR U32787 ( .A(a[774]), .B(n42197), .Z(n32003) );
  NANDN U32788 ( .A(n32003), .B(n42173), .Z(n31964) );
  NANDN U32789 ( .A(n31962), .B(n42172), .Z(n31963) );
  NAND U32790 ( .A(n31964), .B(n31963), .Z(n32012) );
  NAND U32791 ( .A(b[7]), .B(a[770]), .Z(n32013) );
  XNOR U32792 ( .A(n32012), .B(n32013), .Z(n32015) );
  XOR U32793 ( .A(n32014), .B(n32015), .Z(n32021) );
  NANDN U32794 ( .A(n31965), .B(n42093), .Z(n31967) );
  XOR U32795 ( .A(n42134), .B(a[776]), .Z(n32006) );
  NANDN U32796 ( .A(n32006), .B(n42095), .Z(n31966) );
  NAND U32797 ( .A(n31967), .B(n31966), .Z(n32019) );
  NANDN U32798 ( .A(n31968), .B(n42231), .Z(n31970) );
  XOR U32799 ( .A(n226), .B(a[772]), .Z(n32009) );
  NANDN U32800 ( .A(n32009), .B(n42234), .Z(n31969) );
  AND U32801 ( .A(n31970), .B(n31969), .Z(n32018) );
  XNOR U32802 ( .A(n32019), .B(n32018), .Z(n32020) );
  XNOR U32803 ( .A(n32021), .B(n32020), .Z(n32025) );
  NANDN U32804 ( .A(n31972), .B(n31971), .Z(n31976) );
  NAND U32805 ( .A(n31974), .B(n31973), .Z(n31975) );
  AND U32806 ( .A(n31976), .B(n31975), .Z(n32024) );
  XOR U32807 ( .A(n32025), .B(n32024), .Z(n32026) );
  NANDN U32808 ( .A(n31978), .B(n31977), .Z(n31982) );
  NANDN U32809 ( .A(n31980), .B(n31979), .Z(n31981) );
  NAND U32810 ( .A(n31982), .B(n31981), .Z(n32027) );
  XOR U32811 ( .A(n32026), .B(n32027), .Z(n31994) );
  OR U32812 ( .A(n31984), .B(n31983), .Z(n31988) );
  NANDN U32813 ( .A(n31986), .B(n31985), .Z(n31987) );
  NAND U32814 ( .A(n31988), .B(n31987), .Z(n31995) );
  XNOR U32815 ( .A(n31994), .B(n31995), .Z(n31996) );
  XNOR U32816 ( .A(n31997), .B(n31996), .Z(n32030) );
  XNOR U32817 ( .A(n32030), .B(sreg[1794]), .Z(n32032) );
  NAND U32818 ( .A(n31989), .B(sreg[1793]), .Z(n31993) );
  OR U32819 ( .A(n31991), .B(n31990), .Z(n31992) );
  AND U32820 ( .A(n31993), .B(n31992), .Z(n32031) );
  XOR U32821 ( .A(n32032), .B(n32031), .Z(c[1794]) );
  NANDN U32822 ( .A(n31995), .B(n31994), .Z(n31999) );
  NAND U32823 ( .A(n31997), .B(n31996), .Z(n31998) );
  NAND U32824 ( .A(n31999), .B(n31998), .Z(n32038) );
  NAND U32825 ( .A(b[0]), .B(a[779]), .Z(n32000) );
  XNOR U32826 ( .A(b[1]), .B(n32000), .Z(n32002) );
  NAND U32827 ( .A(n126), .B(a[778]), .Z(n32001) );
  AND U32828 ( .A(n32002), .B(n32001), .Z(n32055) );
  XOR U32829 ( .A(a[775]), .B(n42197), .Z(n32044) );
  NANDN U32830 ( .A(n32044), .B(n42173), .Z(n32005) );
  NANDN U32831 ( .A(n32003), .B(n42172), .Z(n32004) );
  NAND U32832 ( .A(n32005), .B(n32004), .Z(n32053) );
  NAND U32833 ( .A(b[7]), .B(a[771]), .Z(n32054) );
  XNOR U32834 ( .A(n32053), .B(n32054), .Z(n32056) );
  XOR U32835 ( .A(n32055), .B(n32056), .Z(n32062) );
  NANDN U32836 ( .A(n32006), .B(n42093), .Z(n32008) );
  XOR U32837 ( .A(n42134), .B(a[777]), .Z(n32047) );
  NANDN U32838 ( .A(n32047), .B(n42095), .Z(n32007) );
  NAND U32839 ( .A(n32008), .B(n32007), .Z(n32060) );
  NANDN U32840 ( .A(n32009), .B(n42231), .Z(n32011) );
  XOR U32841 ( .A(n226), .B(a[773]), .Z(n32050) );
  NANDN U32842 ( .A(n32050), .B(n42234), .Z(n32010) );
  AND U32843 ( .A(n32011), .B(n32010), .Z(n32059) );
  XNOR U32844 ( .A(n32060), .B(n32059), .Z(n32061) );
  XNOR U32845 ( .A(n32062), .B(n32061), .Z(n32066) );
  NANDN U32846 ( .A(n32013), .B(n32012), .Z(n32017) );
  NAND U32847 ( .A(n32015), .B(n32014), .Z(n32016) );
  AND U32848 ( .A(n32017), .B(n32016), .Z(n32065) );
  XOR U32849 ( .A(n32066), .B(n32065), .Z(n32067) );
  NANDN U32850 ( .A(n32019), .B(n32018), .Z(n32023) );
  NANDN U32851 ( .A(n32021), .B(n32020), .Z(n32022) );
  NAND U32852 ( .A(n32023), .B(n32022), .Z(n32068) );
  XOR U32853 ( .A(n32067), .B(n32068), .Z(n32035) );
  OR U32854 ( .A(n32025), .B(n32024), .Z(n32029) );
  NANDN U32855 ( .A(n32027), .B(n32026), .Z(n32028) );
  NAND U32856 ( .A(n32029), .B(n32028), .Z(n32036) );
  XNOR U32857 ( .A(n32035), .B(n32036), .Z(n32037) );
  XNOR U32858 ( .A(n32038), .B(n32037), .Z(n32071) );
  XNOR U32859 ( .A(n32071), .B(sreg[1795]), .Z(n32073) );
  NAND U32860 ( .A(n32030), .B(sreg[1794]), .Z(n32034) );
  OR U32861 ( .A(n32032), .B(n32031), .Z(n32033) );
  AND U32862 ( .A(n32034), .B(n32033), .Z(n32072) );
  XOR U32863 ( .A(n32073), .B(n32072), .Z(c[1795]) );
  NANDN U32864 ( .A(n32036), .B(n32035), .Z(n32040) );
  NAND U32865 ( .A(n32038), .B(n32037), .Z(n32039) );
  NAND U32866 ( .A(n32040), .B(n32039), .Z(n32079) );
  NAND U32867 ( .A(b[0]), .B(a[780]), .Z(n32041) );
  XNOR U32868 ( .A(b[1]), .B(n32041), .Z(n32043) );
  NAND U32869 ( .A(n126), .B(a[779]), .Z(n32042) );
  AND U32870 ( .A(n32043), .B(n32042), .Z(n32096) );
  XOR U32871 ( .A(a[776]), .B(n42197), .Z(n32085) );
  NANDN U32872 ( .A(n32085), .B(n42173), .Z(n32046) );
  NANDN U32873 ( .A(n32044), .B(n42172), .Z(n32045) );
  NAND U32874 ( .A(n32046), .B(n32045), .Z(n32094) );
  NAND U32875 ( .A(b[7]), .B(a[772]), .Z(n32095) );
  XNOR U32876 ( .A(n32094), .B(n32095), .Z(n32097) );
  XOR U32877 ( .A(n32096), .B(n32097), .Z(n32103) );
  NANDN U32878 ( .A(n32047), .B(n42093), .Z(n32049) );
  XOR U32879 ( .A(n42134), .B(a[778]), .Z(n32088) );
  NANDN U32880 ( .A(n32088), .B(n42095), .Z(n32048) );
  NAND U32881 ( .A(n32049), .B(n32048), .Z(n32101) );
  NANDN U32882 ( .A(n32050), .B(n42231), .Z(n32052) );
  XOR U32883 ( .A(n226), .B(a[774]), .Z(n32091) );
  NANDN U32884 ( .A(n32091), .B(n42234), .Z(n32051) );
  AND U32885 ( .A(n32052), .B(n32051), .Z(n32100) );
  XNOR U32886 ( .A(n32101), .B(n32100), .Z(n32102) );
  XNOR U32887 ( .A(n32103), .B(n32102), .Z(n32107) );
  NANDN U32888 ( .A(n32054), .B(n32053), .Z(n32058) );
  NAND U32889 ( .A(n32056), .B(n32055), .Z(n32057) );
  AND U32890 ( .A(n32058), .B(n32057), .Z(n32106) );
  XOR U32891 ( .A(n32107), .B(n32106), .Z(n32108) );
  NANDN U32892 ( .A(n32060), .B(n32059), .Z(n32064) );
  NANDN U32893 ( .A(n32062), .B(n32061), .Z(n32063) );
  NAND U32894 ( .A(n32064), .B(n32063), .Z(n32109) );
  XOR U32895 ( .A(n32108), .B(n32109), .Z(n32076) );
  OR U32896 ( .A(n32066), .B(n32065), .Z(n32070) );
  NANDN U32897 ( .A(n32068), .B(n32067), .Z(n32069) );
  NAND U32898 ( .A(n32070), .B(n32069), .Z(n32077) );
  XNOR U32899 ( .A(n32076), .B(n32077), .Z(n32078) );
  XNOR U32900 ( .A(n32079), .B(n32078), .Z(n32112) );
  XNOR U32901 ( .A(n32112), .B(sreg[1796]), .Z(n32114) );
  NAND U32902 ( .A(n32071), .B(sreg[1795]), .Z(n32075) );
  OR U32903 ( .A(n32073), .B(n32072), .Z(n32074) );
  AND U32904 ( .A(n32075), .B(n32074), .Z(n32113) );
  XOR U32905 ( .A(n32114), .B(n32113), .Z(c[1796]) );
  NANDN U32906 ( .A(n32077), .B(n32076), .Z(n32081) );
  NAND U32907 ( .A(n32079), .B(n32078), .Z(n32080) );
  NAND U32908 ( .A(n32081), .B(n32080), .Z(n32120) );
  NAND U32909 ( .A(b[0]), .B(a[781]), .Z(n32082) );
  XNOR U32910 ( .A(b[1]), .B(n32082), .Z(n32084) );
  NAND U32911 ( .A(n126), .B(a[780]), .Z(n32083) );
  AND U32912 ( .A(n32084), .B(n32083), .Z(n32137) );
  XOR U32913 ( .A(a[777]), .B(n42197), .Z(n32126) );
  NANDN U32914 ( .A(n32126), .B(n42173), .Z(n32087) );
  NANDN U32915 ( .A(n32085), .B(n42172), .Z(n32086) );
  NAND U32916 ( .A(n32087), .B(n32086), .Z(n32135) );
  NAND U32917 ( .A(b[7]), .B(a[773]), .Z(n32136) );
  XNOR U32918 ( .A(n32135), .B(n32136), .Z(n32138) );
  XOR U32919 ( .A(n32137), .B(n32138), .Z(n32144) );
  NANDN U32920 ( .A(n32088), .B(n42093), .Z(n32090) );
  XOR U32921 ( .A(n42134), .B(a[779]), .Z(n32129) );
  NANDN U32922 ( .A(n32129), .B(n42095), .Z(n32089) );
  NAND U32923 ( .A(n32090), .B(n32089), .Z(n32142) );
  NANDN U32924 ( .A(n32091), .B(n42231), .Z(n32093) );
  XOR U32925 ( .A(n226), .B(a[775]), .Z(n32132) );
  NANDN U32926 ( .A(n32132), .B(n42234), .Z(n32092) );
  AND U32927 ( .A(n32093), .B(n32092), .Z(n32141) );
  XNOR U32928 ( .A(n32142), .B(n32141), .Z(n32143) );
  XNOR U32929 ( .A(n32144), .B(n32143), .Z(n32148) );
  NANDN U32930 ( .A(n32095), .B(n32094), .Z(n32099) );
  NAND U32931 ( .A(n32097), .B(n32096), .Z(n32098) );
  AND U32932 ( .A(n32099), .B(n32098), .Z(n32147) );
  XOR U32933 ( .A(n32148), .B(n32147), .Z(n32149) );
  NANDN U32934 ( .A(n32101), .B(n32100), .Z(n32105) );
  NANDN U32935 ( .A(n32103), .B(n32102), .Z(n32104) );
  NAND U32936 ( .A(n32105), .B(n32104), .Z(n32150) );
  XOR U32937 ( .A(n32149), .B(n32150), .Z(n32117) );
  OR U32938 ( .A(n32107), .B(n32106), .Z(n32111) );
  NANDN U32939 ( .A(n32109), .B(n32108), .Z(n32110) );
  NAND U32940 ( .A(n32111), .B(n32110), .Z(n32118) );
  XNOR U32941 ( .A(n32117), .B(n32118), .Z(n32119) );
  XNOR U32942 ( .A(n32120), .B(n32119), .Z(n32153) );
  XNOR U32943 ( .A(n32153), .B(sreg[1797]), .Z(n32155) );
  NAND U32944 ( .A(n32112), .B(sreg[1796]), .Z(n32116) );
  OR U32945 ( .A(n32114), .B(n32113), .Z(n32115) );
  AND U32946 ( .A(n32116), .B(n32115), .Z(n32154) );
  XOR U32947 ( .A(n32155), .B(n32154), .Z(c[1797]) );
  NANDN U32948 ( .A(n32118), .B(n32117), .Z(n32122) );
  NAND U32949 ( .A(n32120), .B(n32119), .Z(n32121) );
  NAND U32950 ( .A(n32122), .B(n32121), .Z(n32161) );
  NAND U32951 ( .A(b[0]), .B(a[782]), .Z(n32123) );
  XNOR U32952 ( .A(b[1]), .B(n32123), .Z(n32125) );
  NAND U32953 ( .A(n126), .B(a[781]), .Z(n32124) );
  AND U32954 ( .A(n32125), .B(n32124), .Z(n32178) );
  XOR U32955 ( .A(a[778]), .B(n42197), .Z(n32167) );
  NANDN U32956 ( .A(n32167), .B(n42173), .Z(n32128) );
  NANDN U32957 ( .A(n32126), .B(n42172), .Z(n32127) );
  NAND U32958 ( .A(n32128), .B(n32127), .Z(n32176) );
  NAND U32959 ( .A(b[7]), .B(a[774]), .Z(n32177) );
  XNOR U32960 ( .A(n32176), .B(n32177), .Z(n32179) );
  XOR U32961 ( .A(n32178), .B(n32179), .Z(n32185) );
  NANDN U32962 ( .A(n32129), .B(n42093), .Z(n32131) );
  XOR U32963 ( .A(n42134), .B(a[780]), .Z(n32170) );
  NANDN U32964 ( .A(n32170), .B(n42095), .Z(n32130) );
  NAND U32965 ( .A(n32131), .B(n32130), .Z(n32183) );
  NANDN U32966 ( .A(n32132), .B(n42231), .Z(n32134) );
  XOR U32967 ( .A(n226), .B(a[776]), .Z(n32173) );
  NANDN U32968 ( .A(n32173), .B(n42234), .Z(n32133) );
  AND U32969 ( .A(n32134), .B(n32133), .Z(n32182) );
  XNOR U32970 ( .A(n32183), .B(n32182), .Z(n32184) );
  XNOR U32971 ( .A(n32185), .B(n32184), .Z(n32189) );
  NANDN U32972 ( .A(n32136), .B(n32135), .Z(n32140) );
  NAND U32973 ( .A(n32138), .B(n32137), .Z(n32139) );
  AND U32974 ( .A(n32140), .B(n32139), .Z(n32188) );
  XOR U32975 ( .A(n32189), .B(n32188), .Z(n32190) );
  NANDN U32976 ( .A(n32142), .B(n32141), .Z(n32146) );
  NANDN U32977 ( .A(n32144), .B(n32143), .Z(n32145) );
  NAND U32978 ( .A(n32146), .B(n32145), .Z(n32191) );
  XOR U32979 ( .A(n32190), .B(n32191), .Z(n32158) );
  OR U32980 ( .A(n32148), .B(n32147), .Z(n32152) );
  NANDN U32981 ( .A(n32150), .B(n32149), .Z(n32151) );
  NAND U32982 ( .A(n32152), .B(n32151), .Z(n32159) );
  XNOR U32983 ( .A(n32158), .B(n32159), .Z(n32160) );
  XNOR U32984 ( .A(n32161), .B(n32160), .Z(n32194) );
  XNOR U32985 ( .A(n32194), .B(sreg[1798]), .Z(n32196) );
  NAND U32986 ( .A(n32153), .B(sreg[1797]), .Z(n32157) );
  OR U32987 ( .A(n32155), .B(n32154), .Z(n32156) );
  AND U32988 ( .A(n32157), .B(n32156), .Z(n32195) );
  XOR U32989 ( .A(n32196), .B(n32195), .Z(c[1798]) );
  NANDN U32990 ( .A(n32159), .B(n32158), .Z(n32163) );
  NAND U32991 ( .A(n32161), .B(n32160), .Z(n32162) );
  NAND U32992 ( .A(n32163), .B(n32162), .Z(n32202) );
  NAND U32993 ( .A(b[0]), .B(a[783]), .Z(n32164) );
  XNOR U32994 ( .A(b[1]), .B(n32164), .Z(n32166) );
  NAND U32995 ( .A(n126), .B(a[782]), .Z(n32165) );
  AND U32996 ( .A(n32166), .B(n32165), .Z(n32219) );
  XOR U32997 ( .A(a[779]), .B(n42197), .Z(n32208) );
  NANDN U32998 ( .A(n32208), .B(n42173), .Z(n32169) );
  NANDN U32999 ( .A(n32167), .B(n42172), .Z(n32168) );
  NAND U33000 ( .A(n32169), .B(n32168), .Z(n32217) );
  NAND U33001 ( .A(b[7]), .B(a[775]), .Z(n32218) );
  XNOR U33002 ( .A(n32217), .B(n32218), .Z(n32220) );
  XOR U33003 ( .A(n32219), .B(n32220), .Z(n32226) );
  NANDN U33004 ( .A(n32170), .B(n42093), .Z(n32172) );
  XOR U33005 ( .A(n42134), .B(a[781]), .Z(n32211) );
  NANDN U33006 ( .A(n32211), .B(n42095), .Z(n32171) );
  NAND U33007 ( .A(n32172), .B(n32171), .Z(n32224) );
  NANDN U33008 ( .A(n32173), .B(n42231), .Z(n32175) );
  XOR U33009 ( .A(n226), .B(a[777]), .Z(n32214) );
  NANDN U33010 ( .A(n32214), .B(n42234), .Z(n32174) );
  AND U33011 ( .A(n32175), .B(n32174), .Z(n32223) );
  XNOR U33012 ( .A(n32224), .B(n32223), .Z(n32225) );
  XNOR U33013 ( .A(n32226), .B(n32225), .Z(n32230) );
  NANDN U33014 ( .A(n32177), .B(n32176), .Z(n32181) );
  NAND U33015 ( .A(n32179), .B(n32178), .Z(n32180) );
  AND U33016 ( .A(n32181), .B(n32180), .Z(n32229) );
  XOR U33017 ( .A(n32230), .B(n32229), .Z(n32231) );
  NANDN U33018 ( .A(n32183), .B(n32182), .Z(n32187) );
  NANDN U33019 ( .A(n32185), .B(n32184), .Z(n32186) );
  NAND U33020 ( .A(n32187), .B(n32186), .Z(n32232) );
  XOR U33021 ( .A(n32231), .B(n32232), .Z(n32199) );
  OR U33022 ( .A(n32189), .B(n32188), .Z(n32193) );
  NANDN U33023 ( .A(n32191), .B(n32190), .Z(n32192) );
  NAND U33024 ( .A(n32193), .B(n32192), .Z(n32200) );
  XNOR U33025 ( .A(n32199), .B(n32200), .Z(n32201) );
  XNOR U33026 ( .A(n32202), .B(n32201), .Z(n32235) );
  XNOR U33027 ( .A(n32235), .B(sreg[1799]), .Z(n32237) );
  NAND U33028 ( .A(n32194), .B(sreg[1798]), .Z(n32198) );
  OR U33029 ( .A(n32196), .B(n32195), .Z(n32197) );
  AND U33030 ( .A(n32198), .B(n32197), .Z(n32236) );
  XOR U33031 ( .A(n32237), .B(n32236), .Z(c[1799]) );
  NANDN U33032 ( .A(n32200), .B(n32199), .Z(n32204) );
  NAND U33033 ( .A(n32202), .B(n32201), .Z(n32203) );
  NAND U33034 ( .A(n32204), .B(n32203), .Z(n32243) );
  NAND U33035 ( .A(b[0]), .B(a[784]), .Z(n32205) );
  XNOR U33036 ( .A(b[1]), .B(n32205), .Z(n32207) );
  NAND U33037 ( .A(n127), .B(a[783]), .Z(n32206) );
  AND U33038 ( .A(n32207), .B(n32206), .Z(n32260) );
  XOR U33039 ( .A(a[780]), .B(n42197), .Z(n32249) );
  NANDN U33040 ( .A(n32249), .B(n42173), .Z(n32210) );
  NANDN U33041 ( .A(n32208), .B(n42172), .Z(n32209) );
  NAND U33042 ( .A(n32210), .B(n32209), .Z(n32258) );
  NAND U33043 ( .A(b[7]), .B(a[776]), .Z(n32259) );
  XNOR U33044 ( .A(n32258), .B(n32259), .Z(n32261) );
  XOR U33045 ( .A(n32260), .B(n32261), .Z(n32267) );
  NANDN U33046 ( .A(n32211), .B(n42093), .Z(n32213) );
  XOR U33047 ( .A(n42134), .B(a[782]), .Z(n32252) );
  NANDN U33048 ( .A(n32252), .B(n42095), .Z(n32212) );
  NAND U33049 ( .A(n32213), .B(n32212), .Z(n32265) );
  NANDN U33050 ( .A(n32214), .B(n42231), .Z(n32216) );
  XOR U33051 ( .A(n226), .B(a[778]), .Z(n32255) );
  NANDN U33052 ( .A(n32255), .B(n42234), .Z(n32215) );
  AND U33053 ( .A(n32216), .B(n32215), .Z(n32264) );
  XNOR U33054 ( .A(n32265), .B(n32264), .Z(n32266) );
  XNOR U33055 ( .A(n32267), .B(n32266), .Z(n32271) );
  NANDN U33056 ( .A(n32218), .B(n32217), .Z(n32222) );
  NAND U33057 ( .A(n32220), .B(n32219), .Z(n32221) );
  AND U33058 ( .A(n32222), .B(n32221), .Z(n32270) );
  XOR U33059 ( .A(n32271), .B(n32270), .Z(n32272) );
  NANDN U33060 ( .A(n32224), .B(n32223), .Z(n32228) );
  NANDN U33061 ( .A(n32226), .B(n32225), .Z(n32227) );
  NAND U33062 ( .A(n32228), .B(n32227), .Z(n32273) );
  XOR U33063 ( .A(n32272), .B(n32273), .Z(n32240) );
  OR U33064 ( .A(n32230), .B(n32229), .Z(n32234) );
  NANDN U33065 ( .A(n32232), .B(n32231), .Z(n32233) );
  NAND U33066 ( .A(n32234), .B(n32233), .Z(n32241) );
  XNOR U33067 ( .A(n32240), .B(n32241), .Z(n32242) );
  XNOR U33068 ( .A(n32243), .B(n32242), .Z(n32276) );
  XNOR U33069 ( .A(n32276), .B(sreg[1800]), .Z(n32278) );
  NAND U33070 ( .A(n32235), .B(sreg[1799]), .Z(n32239) );
  OR U33071 ( .A(n32237), .B(n32236), .Z(n32238) );
  AND U33072 ( .A(n32239), .B(n32238), .Z(n32277) );
  XOR U33073 ( .A(n32278), .B(n32277), .Z(c[1800]) );
  NANDN U33074 ( .A(n32241), .B(n32240), .Z(n32245) );
  NAND U33075 ( .A(n32243), .B(n32242), .Z(n32244) );
  NAND U33076 ( .A(n32245), .B(n32244), .Z(n32284) );
  NAND U33077 ( .A(b[0]), .B(a[785]), .Z(n32246) );
  XNOR U33078 ( .A(b[1]), .B(n32246), .Z(n32248) );
  NAND U33079 ( .A(n127), .B(a[784]), .Z(n32247) );
  AND U33080 ( .A(n32248), .B(n32247), .Z(n32301) );
  XOR U33081 ( .A(a[781]), .B(n42197), .Z(n32290) );
  NANDN U33082 ( .A(n32290), .B(n42173), .Z(n32251) );
  NANDN U33083 ( .A(n32249), .B(n42172), .Z(n32250) );
  NAND U33084 ( .A(n32251), .B(n32250), .Z(n32299) );
  NAND U33085 ( .A(b[7]), .B(a[777]), .Z(n32300) );
  XNOR U33086 ( .A(n32299), .B(n32300), .Z(n32302) );
  XOR U33087 ( .A(n32301), .B(n32302), .Z(n32308) );
  NANDN U33088 ( .A(n32252), .B(n42093), .Z(n32254) );
  XOR U33089 ( .A(n42134), .B(a[783]), .Z(n32293) );
  NANDN U33090 ( .A(n32293), .B(n42095), .Z(n32253) );
  NAND U33091 ( .A(n32254), .B(n32253), .Z(n32306) );
  NANDN U33092 ( .A(n32255), .B(n42231), .Z(n32257) );
  XOR U33093 ( .A(n227), .B(a[779]), .Z(n32296) );
  NANDN U33094 ( .A(n32296), .B(n42234), .Z(n32256) );
  AND U33095 ( .A(n32257), .B(n32256), .Z(n32305) );
  XNOR U33096 ( .A(n32306), .B(n32305), .Z(n32307) );
  XNOR U33097 ( .A(n32308), .B(n32307), .Z(n32312) );
  NANDN U33098 ( .A(n32259), .B(n32258), .Z(n32263) );
  NAND U33099 ( .A(n32261), .B(n32260), .Z(n32262) );
  AND U33100 ( .A(n32263), .B(n32262), .Z(n32311) );
  XOR U33101 ( .A(n32312), .B(n32311), .Z(n32313) );
  NANDN U33102 ( .A(n32265), .B(n32264), .Z(n32269) );
  NANDN U33103 ( .A(n32267), .B(n32266), .Z(n32268) );
  NAND U33104 ( .A(n32269), .B(n32268), .Z(n32314) );
  XOR U33105 ( .A(n32313), .B(n32314), .Z(n32281) );
  OR U33106 ( .A(n32271), .B(n32270), .Z(n32275) );
  NANDN U33107 ( .A(n32273), .B(n32272), .Z(n32274) );
  NAND U33108 ( .A(n32275), .B(n32274), .Z(n32282) );
  XNOR U33109 ( .A(n32281), .B(n32282), .Z(n32283) );
  XNOR U33110 ( .A(n32284), .B(n32283), .Z(n32317) );
  XNOR U33111 ( .A(n32317), .B(sreg[1801]), .Z(n32319) );
  NAND U33112 ( .A(n32276), .B(sreg[1800]), .Z(n32280) );
  OR U33113 ( .A(n32278), .B(n32277), .Z(n32279) );
  AND U33114 ( .A(n32280), .B(n32279), .Z(n32318) );
  XOR U33115 ( .A(n32319), .B(n32318), .Z(c[1801]) );
  NANDN U33116 ( .A(n32282), .B(n32281), .Z(n32286) );
  NAND U33117 ( .A(n32284), .B(n32283), .Z(n32285) );
  NAND U33118 ( .A(n32286), .B(n32285), .Z(n32325) );
  NAND U33119 ( .A(b[0]), .B(a[786]), .Z(n32287) );
  XNOR U33120 ( .A(b[1]), .B(n32287), .Z(n32289) );
  NAND U33121 ( .A(n127), .B(a[785]), .Z(n32288) );
  AND U33122 ( .A(n32289), .B(n32288), .Z(n32342) );
  XOR U33123 ( .A(a[782]), .B(n42197), .Z(n32331) );
  NANDN U33124 ( .A(n32331), .B(n42173), .Z(n32292) );
  NANDN U33125 ( .A(n32290), .B(n42172), .Z(n32291) );
  NAND U33126 ( .A(n32292), .B(n32291), .Z(n32340) );
  NAND U33127 ( .A(b[7]), .B(a[778]), .Z(n32341) );
  XNOR U33128 ( .A(n32340), .B(n32341), .Z(n32343) );
  XOR U33129 ( .A(n32342), .B(n32343), .Z(n32349) );
  NANDN U33130 ( .A(n32293), .B(n42093), .Z(n32295) );
  XOR U33131 ( .A(n42134), .B(a[784]), .Z(n32334) );
  NANDN U33132 ( .A(n32334), .B(n42095), .Z(n32294) );
  NAND U33133 ( .A(n32295), .B(n32294), .Z(n32347) );
  NANDN U33134 ( .A(n32296), .B(n42231), .Z(n32298) );
  XOR U33135 ( .A(n227), .B(a[780]), .Z(n32337) );
  NANDN U33136 ( .A(n32337), .B(n42234), .Z(n32297) );
  AND U33137 ( .A(n32298), .B(n32297), .Z(n32346) );
  XNOR U33138 ( .A(n32347), .B(n32346), .Z(n32348) );
  XNOR U33139 ( .A(n32349), .B(n32348), .Z(n32353) );
  NANDN U33140 ( .A(n32300), .B(n32299), .Z(n32304) );
  NAND U33141 ( .A(n32302), .B(n32301), .Z(n32303) );
  AND U33142 ( .A(n32304), .B(n32303), .Z(n32352) );
  XOR U33143 ( .A(n32353), .B(n32352), .Z(n32354) );
  NANDN U33144 ( .A(n32306), .B(n32305), .Z(n32310) );
  NANDN U33145 ( .A(n32308), .B(n32307), .Z(n32309) );
  NAND U33146 ( .A(n32310), .B(n32309), .Z(n32355) );
  XOR U33147 ( .A(n32354), .B(n32355), .Z(n32322) );
  OR U33148 ( .A(n32312), .B(n32311), .Z(n32316) );
  NANDN U33149 ( .A(n32314), .B(n32313), .Z(n32315) );
  NAND U33150 ( .A(n32316), .B(n32315), .Z(n32323) );
  XNOR U33151 ( .A(n32322), .B(n32323), .Z(n32324) );
  XNOR U33152 ( .A(n32325), .B(n32324), .Z(n32358) );
  XNOR U33153 ( .A(n32358), .B(sreg[1802]), .Z(n32360) );
  NAND U33154 ( .A(n32317), .B(sreg[1801]), .Z(n32321) );
  OR U33155 ( .A(n32319), .B(n32318), .Z(n32320) );
  AND U33156 ( .A(n32321), .B(n32320), .Z(n32359) );
  XOR U33157 ( .A(n32360), .B(n32359), .Z(c[1802]) );
  NANDN U33158 ( .A(n32323), .B(n32322), .Z(n32327) );
  NAND U33159 ( .A(n32325), .B(n32324), .Z(n32326) );
  NAND U33160 ( .A(n32327), .B(n32326), .Z(n32366) );
  NAND U33161 ( .A(b[0]), .B(a[787]), .Z(n32328) );
  XNOR U33162 ( .A(b[1]), .B(n32328), .Z(n32330) );
  NAND U33163 ( .A(n127), .B(a[786]), .Z(n32329) );
  AND U33164 ( .A(n32330), .B(n32329), .Z(n32383) );
  XOR U33165 ( .A(a[783]), .B(n42197), .Z(n32372) );
  NANDN U33166 ( .A(n32372), .B(n42173), .Z(n32333) );
  NANDN U33167 ( .A(n32331), .B(n42172), .Z(n32332) );
  NAND U33168 ( .A(n32333), .B(n32332), .Z(n32381) );
  NAND U33169 ( .A(b[7]), .B(a[779]), .Z(n32382) );
  XNOR U33170 ( .A(n32381), .B(n32382), .Z(n32384) );
  XOR U33171 ( .A(n32383), .B(n32384), .Z(n32390) );
  NANDN U33172 ( .A(n32334), .B(n42093), .Z(n32336) );
  XOR U33173 ( .A(n42134), .B(a[785]), .Z(n32375) );
  NANDN U33174 ( .A(n32375), .B(n42095), .Z(n32335) );
  NAND U33175 ( .A(n32336), .B(n32335), .Z(n32388) );
  NANDN U33176 ( .A(n32337), .B(n42231), .Z(n32339) );
  XOR U33177 ( .A(n227), .B(a[781]), .Z(n32378) );
  NANDN U33178 ( .A(n32378), .B(n42234), .Z(n32338) );
  AND U33179 ( .A(n32339), .B(n32338), .Z(n32387) );
  XNOR U33180 ( .A(n32388), .B(n32387), .Z(n32389) );
  XNOR U33181 ( .A(n32390), .B(n32389), .Z(n32394) );
  NANDN U33182 ( .A(n32341), .B(n32340), .Z(n32345) );
  NAND U33183 ( .A(n32343), .B(n32342), .Z(n32344) );
  AND U33184 ( .A(n32345), .B(n32344), .Z(n32393) );
  XOR U33185 ( .A(n32394), .B(n32393), .Z(n32395) );
  NANDN U33186 ( .A(n32347), .B(n32346), .Z(n32351) );
  NANDN U33187 ( .A(n32349), .B(n32348), .Z(n32350) );
  NAND U33188 ( .A(n32351), .B(n32350), .Z(n32396) );
  XOR U33189 ( .A(n32395), .B(n32396), .Z(n32363) );
  OR U33190 ( .A(n32353), .B(n32352), .Z(n32357) );
  NANDN U33191 ( .A(n32355), .B(n32354), .Z(n32356) );
  NAND U33192 ( .A(n32357), .B(n32356), .Z(n32364) );
  XNOR U33193 ( .A(n32363), .B(n32364), .Z(n32365) );
  XNOR U33194 ( .A(n32366), .B(n32365), .Z(n32399) );
  XNOR U33195 ( .A(n32399), .B(sreg[1803]), .Z(n32401) );
  NAND U33196 ( .A(n32358), .B(sreg[1802]), .Z(n32362) );
  OR U33197 ( .A(n32360), .B(n32359), .Z(n32361) );
  AND U33198 ( .A(n32362), .B(n32361), .Z(n32400) );
  XOR U33199 ( .A(n32401), .B(n32400), .Z(c[1803]) );
  NANDN U33200 ( .A(n32364), .B(n32363), .Z(n32368) );
  NAND U33201 ( .A(n32366), .B(n32365), .Z(n32367) );
  NAND U33202 ( .A(n32368), .B(n32367), .Z(n32407) );
  NAND U33203 ( .A(b[0]), .B(a[788]), .Z(n32369) );
  XNOR U33204 ( .A(b[1]), .B(n32369), .Z(n32371) );
  NAND U33205 ( .A(n127), .B(a[787]), .Z(n32370) );
  AND U33206 ( .A(n32371), .B(n32370), .Z(n32424) );
  XOR U33207 ( .A(a[784]), .B(n42197), .Z(n32413) );
  NANDN U33208 ( .A(n32413), .B(n42173), .Z(n32374) );
  NANDN U33209 ( .A(n32372), .B(n42172), .Z(n32373) );
  NAND U33210 ( .A(n32374), .B(n32373), .Z(n32422) );
  NAND U33211 ( .A(b[7]), .B(a[780]), .Z(n32423) );
  XNOR U33212 ( .A(n32422), .B(n32423), .Z(n32425) );
  XOR U33213 ( .A(n32424), .B(n32425), .Z(n32431) );
  NANDN U33214 ( .A(n32375), .B(n42093), .Z(n32377) );
  XOR U33215 ( .A(n42134), .B(a[786]), .Z(n32416) );
  NANDN U33216 ( .A(n32416), .B(n42095), .Z(n32376) );
  NAND U33217 ( .A(n32377), .B(n32376), .Z(n32429) );
  NANDN U33218 ( .A(n32378), .B(n42231), .Z(n32380) );
  XOR U33219 ( .A(n227), .B(a[782]), .Z(n32419) );
  NANDN U33220 ( .A(n32419), .B(n42234), .Z(n32379) );
  AND U33221 ( .A(n32380), .B(n32379), .Z(n32428) );
  XNOR U33222 ( .A(n32429), .B(n32428), .Z(n32430) );
  XNOR U33223 ( .A(n32431), .B(n32430), .Z(n32435) );
  NANDN U33224 ( .A(n32382), .B(n32381), .Z(n32386) );
  NAND U33225 ( .A(n32384), .B(n32383), .Z(n32385) );
  AND U33226 ( .A(n32386), .B(n32385), .Z(n32434) );
  XOR U33227 ( .A(n32435), .B(n32434), .Z(n32436) );
  NANDN U33228 ( .A(n32388), .B(n32387), .Z(n32392) );
  NANDN U33229 ( .A(n32390), .B(n32389), .Z(n32391) );
  NAND U33230 ( .A(n32392), .B(n32391), .Z(n32437) );
  XOR U33231 ( .A(n32436), .B(n32437), .Z(n32404) );
  OR U33232 ( .A(n32394), .B(n32393), .Z(n32398) );
  NANDN U33233 ( .A(n32396), .B(n32395), .Z(n32397) );
  NAND U33234 ( .A(n32398), .B(n32397), .Z(n32405) );
  XNOR U33235 ( .A(n32404), .B(n32405), .Z(n32406) );
  XNOR U33236 ( .A(n32407), .B(n32406), .Z(n32440) );
  XNOR U33237 ( .A(n32440), .B(sreg[1804]), .Z(n32442) );
  NAND U33238 ( .A(n32399), .B(sreg[1803]), .Z(n32403) );
  OR U33239 ( .A(n32401), .B(n32400), .Z(n32402) );
  AND U33240 ( .A(n32403), .B(n32402), .Z(n32441) );
  XOR U33241 ( .A(n32442), .B(n32441), .Z(c[1804]) );
  NANDN U33242 ( .A(n32405), .B(n32404), .Z(n32409) );
  NAND U33243 ( .A(n32407), .B(n32406), .Z(n32408) );
  NAND U33244 ( .A(n32409), .B(n32408), .Z(n32448) );
  NAND U33245 ( .A(b[0]), .B(a[789]), .Z(n32410) );
  XNOR U33246 ( .A(b[1]), .B(n32410), .Z(n32412) );
  NAND U33247 ( .A(n127), .B(a[788]), .Z(n32411) );
  AND U33248 ( .A(n32412), .B(n32411), .Z(n32465) );
  XOR U33249 ( .A(a[785]), .B(n42197), .Z(n32454) );
  NANDN U33250 ( .A(n32454), .B(n42173), .Z(n32415) );
  NANDN U33251 ( .A(n32413), .B(n42172), .Z(n32414) );
  NAND U33252 ( .A(n32415), .B(n32414), .Z(n32463) );
  NAND U33253 ( .A(b[7]), .B(a[781]), .Z(n32464) );
  XNOR U33254 ( .A(n32463), .B(n32464), .Z(n32466) );
  XOR U33255 ( .A(n32465), .B(n32466), .Z(n32472) );
  NANDN U33256 ( .A(n32416), .B(n42093), .Z(n32418) );
  XOR U33257 ( .A(n42134), .B(a[787]), .Z(n32457) );
  NANDN U33258 ( .A(n32457), .B(n42095), .Z(n32417) );
  NAND U33259 ( .A(n32418), .B(n32417), .Z(n32470) );
  NANDN U33260 ( .A(n32419), .B(n42231), .Z(n32421) );
  XOR U33261 ( .A(n227), .B(a[783]), .Z(n32460) );
  NANDN U33262 ( .A(n32460), .B(n42234), .Z(n32420) );
  AND U33263 ( .A(n32421), .B(n32420), .Z(n32469) );
  XNOR U33264 ( .A(n32470), .B(n32469), .Z(n32471) );
  XNOR U33265 ( .A(n32472), .B(n32471), .Z(n32476) );
  NANDN U33266 ( .A(n32423), .B(n32422), .Z(n32427) );
  NAND U33267 ( .A(n32425), .B(n32424), .Z(n32426) );
  AND U33268 ( .A(n32427), .B(n32426), .Z(n32475) );
  XOR U33269 ( .A(n32476), .B(n32475), .Z(n32477) );
  NANDN U33270 ( .A(n32429), .B(n32428), .Z(n32433) );
  NANDN U33271 ( .A(n32431), .B(n32430), .Z(n32432) );
  NAND U33272 ( .A(n32433), .B(n32432), .Z(n32478) );
  XOR U33273 ( .A(n32477), .B(n32478), .Z(n32445) );
  OR U33274 ( .A(n32435), .B(n32434), .Z(n32439) );
  NANDN U33275 ( .A(n32437), .B(n32436), .Z(n32438) );
  NAND U33276 ( .A(n32439), .B(n32438), .Z(n32446) );
  XNOR U33277 ( .A(n32445), .B(n32446), .Z(n32447) );
  XNOR U33278 ( .A(n32448), .B(n32447), .Z(n32481) );
  XNOR U33279 ( .A(n32481), .B(sreg[1805]), .Z(n32483) );
  NAND U33280 ( .A(n32440), .B(sreg[1804]), .Z(n32444) );
  OR U33281 ( .A(n32442), .B(n32441), .Z(n32443) );
  AND U33282 ( .A(n32444), .B(n32443), .Z(n32482) );
  XOR U33283 ( .A(n32483), .B(n32482), .Z(c[1805]) );
  NANDN U33284 ( .A(n32446), .B(n32445), .Z(n32450) );
  NAND U33285 ( .A(n32448), .B(n32447), .Z(n32449) );
  NAND U33286 ( .A(n32450), .B(n32449), .Z(n32489) );
  NAND U33287 ( .A(b[0]), .B(a[790]), .Z(n32451) );
  XNOR U33288 ( .A(b[1]), .B(n32451), .Z(n32453) );
  NAND U33289 ( .A(n127), .B(a[789]), .Z(n32452) );
  AND U33290 ( .A(n32453), .B(n32452), .Z(n32506) );
  XOR U33291 ( .A(a[786]), .B(n42197), .Z(n32495) );
  NANDN U33292 ( .A(n32495), .B(n42173), .Z(n32456) );
  NANDN U33293 ( .A(n32454), .B(n42172), .Z(n32455) );
  NAND U33294 ( .A(n32456), .B(n32455), .Z(n32504) );
  NAND U33295 ( .A(b[7]), .B(a[782]), .Z(n32505) );
  XNOR U33296 ( .A(n32504), .B(n32505), .Z(n32507) );
  XOR U33297 ( .A(n32506), .B(n32507), .Z(n32513) );
  NANDN U33298 ( .A(n32457), .B(n42093), .Z(n32459) );
  XOR U33299 ( .A(n42134), .B(a[788]), .Z(n32498) );
  NANDN U33300 ( .A(n32498), .B(n42095), .Z(n32458) );
  NAND U33301 ( .A(n32459), .B(n32458), .Z(n32511) );
  NANDN U33302 ( .A(n32460), .B(n42231), .Z(n32462) );
  XOR U33303 ( .A(n227), .B(a[784]), .Z(n32501) );
  NANDN U33304 ( .A(n32501), .B(n42234), .Z(n32461) );
  AND U33305 ( .A(n32462), .B(n32461), .Z(n32510) );
  XNOR U33306 ( .A(n32511), .B(n32510), .Z(n32512) );
  XNOR U33307 ( .A(n32513), .B(n32512), .Z(n32517) );
  NANDN U33308 ( .A(n32464), .B(n32463), .Z(n32468) );
  NAND U33309 ( .A(n32466), .B(n32465), .Z(n32467) );
  AND U33310 ( .A(n32468), .B(n32467), .Z(n32516) );
  XOR U33311 ( .A(n32517), .B(n32516), .Z(n32518) );
  NANDN U33312 ( .A(n32470), .B(n32469), .Z(n32474) );
  NANDN U33313 ( .A(n32472), .B(n32471), .Z(n32473) );
  NAND U33314 ( .A(n32474), .B(n32473), .Z(n32519) );
  XOR U33315 ( .A(n32518), .B(n32519), .Z(n32486) );
  OR U33316 ( .A(n32476), .B(n32475), .Z(n32480) );
  NANDN U33317 ( .A(n32478), .B(n32477), .Z(n32479) );
  NAND U33318 ( .A(n32480), .B(n32479), .Z(n32487) );
  XNOR U33319 ( .A(n32486), .B(n32487), .Z(n32488) );
  XNOR U33320 ( .A(n32489), .B(n32488), .Z(n32522) );
  XNOR U33321 ( .A(n32522), .B(sreg[1806]), .Z(n32524) );
  NAND U33322 ( .A(n32481), .B(sreg[1805]), .Z(n32485) );
  OR U33323 ( .A(n32483), .B(n32482), .Z(n32484) );
  AND U33324 ( .A(n32485), .B(n32484), .Z(n32523) );
  XOR U33325 ( .A(n32524), .B(n32523), .Z(c[1806]) );
  NANDN U33326 ( .A(n32487), .B(n32486), .Z(n32491) );
  NAND U33327 ( .A(n32489), .B(n32488), .Z(n32490) );
  NAND U33328 ( .A(n32491), .B(n32490), .Z(n32530) );
  NAND U33329 ( .A(b[0]), .B(a[791]), .Z(n32492) );
  XNOR U33330 ( .A(b[1]), .B(n32492), .Z(n32494) );
  NAND U33331 ( .A(n128), .B(a[790]), .Z(n32493) );
  AND U33332 ( .A(n32494), .B(n32493), .Z(n32547) );
  XOR U33333 ( .A(a[787]), .B(n42197), .Z(n32536) );
  NANDN U33334 ( .A(n32536), .B(n42173), .Z(n32497) );
  NANDN U33335 ( .A(n32495), .B(n42172), .Z(n32496) );
  NAND U33336 ( .A(n32497), .B(n32496), .Z(n32545) );
  NAND U33337 ( .A(b[7]), .B(a[783]), .Z(n32546) );
  XNOR U33338 ( .A(n32545), .B(n32546), .Z(n32548) );
  XOR U33339 ( .A(n32547), .B(n32548), .Z(n32554) );
  NANDN U33340 ( .A(n32498), .B(n42093), .Z(n32500) );
  XOR U33341 ( .A(n42134), .B(a[789]), .Z(n32539) );
  NANDN U33342 ( .A(n32539), .B(n42095), .Z(n32499) );
  NAND U33343 ( .A(n32500), .B(n32499), .Z(n32552) );
  NANDN U33344 ( .A(n32501), .B(n42231), .Z(n32503) );
  XOR U33345 ( .A(n227), .B(a[785]), .Z(n32542) );
  NANDN U33346 ( .A(n32542), .B(n42234), .Z(n32502) );
  AND U33347 ( .A(n32503), .B(n32502), .Z(n32551) );
  XNOR U33348 ( .A(n32552), .B(n32551), .Z(n32553) );
  XNOR U33349 ( .A(n32554), .B(n32553), .Z(n32558) );
  NANDN U33350 ( .A(n32505), .B(n32504), .Z(n32509) );
  NAND U33351 ( .A(n32507), .B(n32506), .Z(n32508) );
  AND U33352 ( .A(n32509), .B(n32508), .Z(n32557) );
  XOR U33353 ( .A(n32558), .B(n32557), .Z(n32559) );
  NANDN U33354 ( .A(n32511), .B(n32510), .Z(n32515) );
  NANDN U33355 ( .A(n32513), .B(n32512), .Z(n32514) );
  NAND U33356 ( .A(n32515), .B(n32514), .Z(n32560) );
  XOR U33357 ( .A(n32559), .B(n32560), .Z(n32527) );
  OR U33358 ( .A(n32517), .B(n32516), .Z(n32521) );
  NANDN U33359 ( .A(n32519), .B(n32518), .Z(n32520) );
  NAND U33360 ( .A(n32521), .B(n32520), .Z(n32528) );
  XNOR U33361 ( .A(n32527), .B(n32528), .Z(n32529) );
  XNOR U33362 ( .A(n32530), .B(n32529), .Z(n32563) );
  XNOR U33363 ( .A(n32563), .B(sreg[1807]), .Z(n32565) );
  NAND U33364 ( .A(n32522), .B(sreg[1806]), .Z(n32526) );
  OR U33365 ( .A(n32524), .B(n32523), .Z(n32525) );
  AND U33366 ( .A(n32526), .B(n32525), .Z(n32564) );
  XOR U33367 ( .A(n32565), .B(n32564), .Z(c[1807]) );
  NANDN U33368 ( .A(n32528), .B(n32527), .Z(n32532) );
  NAND U33369 ( .A(n32530), .B(n32529), .Z(n32531) );
  NAND U33370 ( .A(n32532), .B(n32531), .Z(n32571) );
  NAND U33371 ( .A(b[0]), .B(a[792]), .Z(n32533) );
  XNOR U33372 ( .A(b[1]), .B(n32533), .Z(n32535) );
  NAND U33373 ( .A(n128), .B(a[791]), .Z(n32534) );
  AND U33374 ( .A(n32535), .B(n32534), .Z(n32588) );
  XOR U33375 ( .A(a[788]), .B(n42197), .Z(n32577) );
  NANDN U33376 ( .A(n32577), .B(n42173), .Z(n32538) );
  NANDN U33377 ( .A(n32536), .B(n42172), .Z(n32537) );
  NAND U33378 ( .A(n32538), .B(n32537), .Z(n32586) );
  NAND U33379 ( .A(b[7]), .B(a[784]), .Z(n32587) );
  XNOR U33380 ( .A(n32586), .B(n32587), .Z(n32589) );
  XOR U33381 ( .A(n32588), .B(n32589), .Z(n32595) );
  NANDN U33382 ( .A(n32539), .B(n42093), .Z(n32541) );
  XOR U33383 ( .A(n42134), .B(a[790]), .Z(n32580) );
  NANDN U33384 ( .A(n32580), .B(n42095), .Z(n32540) );
  NAND U33385 ( .A(n32541), .B(n32540), .Z(n32593) );
  NANDN U33386 ( .A(n32542), .B(n42231), .Z(n32544) );
  XOR U33387 ( .A(n227), .B(a[786]), .Z(n32583) );
  NANDN U33388 ( .A(n32583), .B(n42234), .Z(n32543) );
  AND U33389 ( .A(n32544), .B(n32543), .Z(n32592) );
  XNOR U33390 ( .A(n32593), .B(n32592), .Z(n32594) );
  XNOR U33391 ( .A(n32595), .B(n32594), .Z(n32599) );
  NANDN U33392 ( .A(n32546), .B(n32545), .Z(n32550) );
  NAND U33393 ( .A(n32548), .B(n32547), .Z(n32549) );
  AND U33394 ( .A(n32550), .B(n32549), .Z(n32598) );
  XOR U33395 ( .A(n32599), .B(n32598), .Z(n32600) );
  NANDN U33396 ( .A(n32552), .B(n32551), .Z(n32556) );
  NANDN U33397 ( .A(n32554), .B(n32553), .Z(n32555) );
  NAND U33398 ( .A(n32556), .B(n32555), .Z(n32601) );
  XOR U33399 ( .A(n32600), .B(n32601), .Z(n32568) );
  OR U33400 ( .A(n32558), .B(n32557), .Z(n32562) );
  NANDN U33401 ( .A(n32560), .B(n32559), .Z(n32561) );
  NAND U33402 ( .A(n32562), .B(n32561), .Z(n32569) );
  XNOR U33403 ( .A(n32568), .B(n32569), .Z(n32570) );
  XNOR U33404 ( .A(n32571), .B(n32570), .Z(n32604) );
  XNOR U33405 ( .A(n32604), .B(sreg[1808]), .Z(n32606) );
  NAND U33406 ( .A(n32563), .B(sreg[1807]), .Z(n32567) );
  OR U33407 ( .A(n32565), .B(n32564), .Z(n32566) );
  AND U33408 ( .A(n32567), .B(n32566), .Z(n32605) );
  XOR U33409 ( .A(n32606), .B(n32605), .Z(c[1808]) );
  NANDN U33410 ( .A(n32569), .B(n32568), .Z(n32573) );
  NAND U33411 ( .A(n32571), .B(n32570), .Z(n32572) );
  NAND U33412 ( .A(n32573), .B(n32572), .Z(n32612) );
  NAND U33413 ( .A(b[0]), .B(a[793]), .Z(n32574) );
  XNOR U33414 ( .A(b[1]), .B(n32574), .Z(n32576) );
  NAND U33415 ( .A(n128), .B(a[792]), .Z(n32575) );
  AND U33416 ( .A(n32576), .B(n32575), .Z(n32629) );
  XOR U33417 ( .A(a[789]), .B(n42197), .Z(n32618) );
  NANDN U33418 ( .A(n32618), .B(n42173), .Z(n32579) );
  NANDN U33419 ( .A(n32577), .B(n42172), .Z(n32578) );
  NAND U33420 ( .A(n32579), .B(n32578), .Z(n32627) );
  NAND U33421 ( .A(b[7]), .B(a[785]), .Z(n32628) );
  XNOR U33422 ( .A(n32627), .B(n32628), .Z(n32630) );
  XOR U33423 ( .A(n32629), .B(n32630), .Z(n32636) );
  NANDN U33424 ( .A(n32580), .B(n42093), .Z(n32582) );
  XOR U33425 ( .A(n42134), .B(a[791]), .Z(n32621) );
  NANDN U33426 ( .A(n32621), .B(n42095), .Z(n32581) );
  NAND U33427 ( .A(n32582), .B(n32581), .Z(n32634) );
  NANDN U33428 ( .A(n32583), .B(n42231), .Z(n32585) );
  XOR U33429 ( .A(n227), .B(a[787]), .Z(n32624) );
  NANDN U33430 ( .A(n32624), .B(n42234), .Z(n32584) );
  AND U33431 ( .A(n32585), .B(n32584), .Z(n32633) );
  XNOR U33432 ( .A(n32634), .B(n32633), .Z(n32635) );
  XNOR U33433 ( .A(n32636), .B(n32635), .Z(n32640) );
  NANDN U33434 ( .A(n32587), .B(n32586), .Z(n32591) );
  NAND U33435 ( .A(n32589), .B(n32588), .Z(n32590) );
  AND U33436 ( .A(n32591), .B(n32590), .Z(n32639) );
  XOR U33437 ( .A(n32640), .B(n32639), .Z(n32641) );
  NANDN U33438 ( .A(n32593), .B(n32592), .Z(n32597) );
  NANDN U33439 ( .A(n32595), .B(n32594), .Z(n32596) );
  NAND U33440 ( .A(n32597), .B(n32596), .Z(n32642) );
  XOR U33441 ( .A(n32641), .B(n32642), .Z(n32609) );
  OR U33442 ( .A(n32599), .B(n32598), .Z(n32603) );
  NANDN U33443 ( .A(n32601), .B(n32600), .Z(n32602) );
  NAND U33444 ( .A(n32603), .B(n32602), .Z(n32610) );
  XNOR U33445 ( .A(n32609), .B(n32610), .Z(n32611) );
  XNOR U33446 ( .A(n32612), .B(n32611), .Z(n32645) );
  XNOR U33447 ( .A(n32645), .B(sreg[1809]), .Z(n32647) );
  NAND U33448 ( .A(n32604), .B(sreg[1808]), .Z(n32608) );
  OR U33449 ( .A(n32606), .B(n32605), .Z(n32607) );
  AND U33450 ( .A(n32608), .B(n32607), .Z(n32646) );
  XOR U33451 ( .A(n32647), .B(n32646), .Z(c[1809]) );
  NANDN U33452 ( .A(n32610), .B(n32609), .Z(n32614) );
  NAND U33453 ( .A(n32612), .B(n32611), .Z(n32613) );
  NAND U33454 ( .A(n32614), .B(n32613), .Z(n32653) );
  NAND U33455 ( .A(b[0]), .B(a[794]), .Z(n32615) );
  XNOR U33456 ( .A(b[1]), .B(n32615), .Z(n32617) );
  NAND U33457 ( .A(n128), .B(a[793]), .Z(n32616) );
  AND U33458 ( .A(n32617), .B(n32616), .Z(n32670) );
  XOR U33459 ( .A(a[790]), .B(n42197), .Z(n32659) );
  NANDN U33460 ( .A(n32659), .B(n42173), .Z(n32620) );
  NANDN U33461 ( .A(n32618), .B(n42172), .Z(n32619) );
  NAND U33462 ( .A(n32620), .B(n32619), .Z(n32668) );
  NAND U33463 ( .A(b[7]), .B(a[786]), .Z(n32669) );
  XNOR U33464 ( .A(n32668), .B(n32669), .Z(n32671) );
  XOR U33465 ( .A(n32670), .B(n32671), .Z(n32677) );
  NANDN U33466 ( .A(n32621), .B(n42093), .Z(n32623) );
  XOR U33467 ( .A(n42134), .B(a[792]), .Z(n32662) );
  NANDN U33468 ( .A(n32662), .B(n42095), .Z(n32622) );
  NAND U33469 ( .A(n32623), .B(n32622), .Z(n32675) );
  NANDN U33470 ( .A(n32624), .B(n42231), .Z(n32626) );
  XOR U33471 ( .A(n227), .B(a[788]), .Z(n32665) );
  NANDN U33472 ( .A(n32665), .B(n42234), .Z(n32625) );
  AND U33473 ( .A(n32626), .B(n32625), .Z(n32674) );
  XNOR U33474 ( .A(n32675), .B(n32674), .Z(n32676) );
  XNOR U33475 ( .A(n32677), .B(n32676), .Z(n32681) );
  NANDN U33476 ( .A(n32628), .B(n32627), .Z(n32632) );
  NAND U33477 ( .A(n32630), .B(n32629), .Z(n32631) );
  AND U33478 ( .A(n32632), .B(n32631), .Z(n32680) );
  XOR U33479 ( .A(n32681), .B(n32680), .Z(n32682) );
  NANDN U33480 ( .A(n32634), .B(n32633), .Z(n32638) );
  NANDN U33481 ( .A(n32636), .B(n32635), .Z(n32637) );
  NAND U33482 ( .A(n32638), .B(n32637), .Z(n32683) );
  XOR U33483 ( .A(n32682), .B(n32683), .Z(n32650) );
  OR U33484 ( .A(n32640), .B(n32639), .Z(n32644) );
  NANDN U33485 ( .A(n32642), .B(n32641), .Z(n32643) );
  NAND U33486 ( .A(n32644), .B(n32643), .Z(n32651) );
  XNOR U33487 ( .A(n32650), .B(n32651), .Z(n32652) );
  XNOR U33488 ( .A(n32653), .B(n32652), .Z(n32686) );
  XNOR U33489 ( .A(n32686), .B(sreg[1810]), .Z(n32688) );
  NAND U33490 ( .A(n32645), .B(sreg[1809]), .Z(n32649) );
  OR U33491 ( .A(n32647), .B(n32646), .Z(n32648) );
  AND U33492 ( .A(n32649), .B(n32648), .Z(n32687) );
  XOR U33493 ( .A(n32688), .B(n32687), .Z(c[1810]) );
  NANDN U33494 ( .A(n32651), .B(n32650), .Z(n32655) );
  NAND U33495 ( .A(n32653), .B(n32652), .Z(n32654) );
  NAND U33496 ( .A(n32655), .B(n32654), .Z(n32694) );
  NAND U33497 ( .A(b[0]), .B(a[795]), .Z(n32656) );
  XNOR U33498 ( .A(b[1]), .B(n32656), .Z(n32658) );
  NAND U33499 ( .A(n128), .B(a[794]), .Z(n32657) );
  AND U33500 ( .A(n32658), .B(n32657), .Z(n32711) );
  XOR U33501 ( .A(a[791]), .B(n42197), .Z(n32700) );
  NANDN U33502 ( .A(n32700), .B(n42173), .Z(n32661) );
  NANDN U33503 ( .A(n32659), .B(n42172), .Z(n32660) );
  NAND U33504 ( .A(n32661), .B(n32660), .Z(n32709) );
  NAND U33505 ( .A(b[7]), .B(a[787]), .Z(n32710) );
  XNOR U33506 ( .A(n32709), .B(n32710), .Z(n32712) );
  XOR U33507 ( .A(n32711), .B(n32712), .Z(n32718) );
  NANDN U33508 ( .A(n32662), .B(n42093), .Z(n32664) );
  XOR U33509 ( .A(n42134), .B(a[793]), .Z(n32703) );
  NANDN U33510 ( .A(n32703), .B(n42095), .Z(n32663) );
  NAND U33511 ( .A(n32664), .B(n32663), .Z(n32716) );
  NANDN U33512 ( .A(n32665), .B(n42231), .Z(n32667) );
  XOR U33513 ( .A(n227), .B(a[789]), .Z(n32706) );
  NANDN U33514 ( .A(n32706), .B(n42234), .Z(n32666) );
  AND U33515 ( .A(n32667), .B(n32666), .Z(n32715) );
  XNOR U33516 ( .A(n32716), .B(n32715), .Z(n32717) );
  XNOR U33517 ( .A(n32718), .B(n32717), .Z(n32722) );
  NANDN U33518 ( .A(n32669), .B(n32668), .Z(n32673) );
  NAND U33519 ( .A(n32671), .B(n32670), .Z(n32672) );
  AND U33520 ( .A(n32673), .B(n32672), .Z(n32721) );
  XOR U33521 ( .A(n32722), .B(n32721), .Z(n32723) );
  NANDN U33522 ( .A(n32675), .B(n32674), .Z(n32679) );
  NANDN U33523 ( .A(n32677), .B(n32676), .Z(n32678) );
  NAND U33524 ( .A(n32679), .B(n32678), .Z(n32724) );
  XOR U33525 ( .A(n32723), .B(n32724), .Z(n32691) );
  OR U33526 ( .A(n32681), .B(n32680), .Z(n32685) );
  NANDN U33527 ( .A(n32683), .B(n32682), .Z(n32684) );
  NAND U33528 ( .A(n32685), .B(n32684), .Z(n32692) );
  XNOR U33529 ( .A(n32691), .B(n32692), .Z(n32693) );
  XNOR U33530 ( .A(n32694), .B(n32693), .Z(n32727) );
  XNOR U33531 ( .A(n32727), .B(sreg[1811]), .Z(n32729) );
  NAND U33532 ( .A(n32686), .B(sreg[1810]), .Z(n32690) );
  OR U33533 ( .A(n32688), .B(n32687), .Z(n32689) );
  AND U33534 ( .A(n32690), .B(n32689), .Z(n32728) );
  XOR U33535 ( .A(n32729), .B(n32728), .Z(c[1811]) );
  NANDN U33536 ( .A(n32692), .B(n32691), .Z(n32696) );
  NAND U33537 ( .A(n32694), .B(n32693), .Z(n32695) );
  NAND U33538 ( .A(n32696), .B(n32695), .Z(n32735) );
  NAND U33539 ( .A(b[0]), .B(a[796]), .Z(n32697) );
  XNOR U33540 ( .A(b[1]), .B(n32697), .Z(n32699) );
  NAND U33541 ( .A(n128), .B(a[795]), .Z(n32698) );
  AND U33542 ( .A(n32699), .B(n32698), .Z(n32752) );
  XOR U33543 ( .A(a[792]), .B(n42197), .Z(n32741) );
  NANDN U33544 ( .A(n32741), .B(n42173), .Z(n32702) );
  NANDN U33545 ( .A(n32700), .B(n42172), .Z(n32701) );
  NAND U33546 ( .A(n32702), .B(n32701), .Z(n32750) );
  NAND U33547 ( .A(b[7]), .B(a[788]), .Z(n32751) );
  XNOR U33548 ( .A(n32750), .B(n32751), .Z(n32753) );
  XOR U33549 ( .A(n32752), .B(n32753), .Z(n32759) );
  NANDN U33550 ( .A(n32703), .B(n42093), .Z(n32705) );
  XOR U33551 ( .A(n42134), .B(a[794]), .Z(n32744) );
  NANDN U33552 ( .A(n32744), .B(n42095), .Z(n32704) );
  NAND U33553 ( .A(n32705), .B(n32704), .Z(n32757) );
  NANDN U33554 ( .A(n32706), .B(n42231), .Z(n32708) );
  XOR U33555 ( .A(n227), .B(a[790]), .Z(n32747) );
  NANDN U33556 ( .A(n32747), .B(n42234), .Z(n32707) );
  AND U33557 ( .A(n32708), .B(n32707), .Z(n32756) );
  XNOR U33558 ( .A(n32757), .B(n32756), .Z(n32758) );
  XNOR U33559 ( .A(n32759), .B(n32758), .Z(n32763) );
  NANDN U33560 ( .A(n32710), .B(n32709), .Z(n32714) );
  NAND U33561 ( .A(n32712), .B(n32711), .Z(n32713) );
  AND U33562 ( .A(n32714), .B(n32713), .Z(n32762) );
  XOR U33563 ( .A(n32763), .B(n32762), .Z(n32764) );
  NANDN U33564 ( .A(n32716), .B(n32715), .Z(n32720) );
  NANDN U33565 ( .A(n32718), .B(n32717), .Z(n32719) );
  NAND U33566 ( .A(n32720), .B(n32719), .Z(n32765) );
  XOR U33567 ( .A(n32764), .B(n32765), .Z(n32732) );
  OR U33568 ( .A(n32722), .B(n32721), .Z(n32726) );
  NANDN U33569 ( .A(n32724), .B(n32723), .Z(n32725) );
  NAND U33570 ( .A(n32726), .B(n32725), .Z(n32733) );
  XNOR U33571 ( .A(n32732), .B(n32733), .Z(n32734) );
  XNOR U33572 ( .A(n32735), .B(n32734), .Z(n32768) );
  XNOR U33573 ( .A(n32768), .B(sreg[1812]), .Z(n32770) );
  NAND U33574 ( .A(n32727), .B(sreg[1811]), .Z(n32731) );
  OR U33575 ( .A(n32729), .B(n32728), .Z(n32730) );
  AND U33576 ( .A(n32731), .B(n32730), .Z(n32769) );
  XOR U33577 ( .A(n32770), .B(n32769), .Z(c[1812]) );
  NANDN U33578 ( .A(n32733), .B(n32732), .Z(n32737) );
  NAND U33579 ( .A(n32735), .B(n32734), .Z(n32736) );
  NAND U33580 ( .A(n32737), .B(n32736), .Z(n32776) );
  NAND U33581 ( .A(b[0]), .B(a[797]), .Z(n32738) );
  XNOR U33582 ( .A(b[1]), .B(n32738), .Z(n32740) );
  NAND U33583 ( .A(n128), .B(a[796]), .Z(n32739) );
  AND U33584 ( .A(n32740), .B(n32739), .Z(n32793) );
  XOR U33585 ( .A(a[793]), .B(n42197), .Z(n32782) );
  NANDN U33586 ( .A(n32782), .B(n42173), .Z(n32743) );
  NANDN U33587 ( .A(n32741), .B(n42172), .Z(n32742) );
  NAND U33588 ( .A(n32743), .B(n32742), .Z(n32791) );
  NAND U33589 ( .A(b[7]), .B(a[789]), .Z(n32792) );
  XNOR U33590 ( .A(n32791), .B(n32792), .Z(n32794) );
  XOR U33591 ( .A(n32793), .B(n32794), .Z(n32800) );
  NANDN U33592 ( .A(n32744), .B(n42093), .Z(n32746) );
  XOR U33593 ( .A(n42134), .B(a[795]), .Z(n32785) );
  NANDN U33594 ( .A(n32785), .B(n42095), .Z(n32745) );
  NAND U33595 ( .A(n32746), .B(n32745), .Z(n32798) );
  NANDN U33596 ( .A(n32747), .B(n42231), .Z(n32749) );
  XOR U33597 ( .A(n228), .B(a[791]), .Z(n32788) );
  NANDN U33598 ( .A(n32788), .B(n42234), .Z(n32748) );
  AND U33599 ( .A(n32749), .B(n32748), .Z(n32797) );
  XNOR U33600 ( .A(n32798), .B(n32797), .Z(n32799) );
  XNOR U33601 ( .A(n32800), .B(n32799), .Z(n32804) );
  NANDN U33602 ( .A(n32751), .B(n32750), .Z(n32755) );
  NAND U33603 ( .A(n32753), .B(n32752), .Z(n32754) );
  AND U33604 ( .A(n32755), .B(n32754), .Z(n32803) );
  XOR U33605 ( .A(n32804), .B(n32803), .Z(n32805) );
  NANDN U33606 ( .A(n32757), .B(n32756), .Z(n32761) );
  NANDN U33607 ( .A(n32759), .B(n32758), .Z(n32760) );
  NAND U33608 ( .A(n32761), .B(n32760), .Z(n32806) );
  XOR U33609 ( .A(n32805), .B(n32806), .Z(n32773) );
  OR U33610 ( .A(n32763), .B(n32762), .Z(n32767) );
  NANDN U33611 ( .A(n32765), .B(n32764), .Z(n32766) );
  NAND U33612 ( .A(n32767), .B(n32766), .Z(n32774) );
  XNOR U33613 ( .A(n32773), .B(n32774), .Z(n32775) );
  XNOR U33614 ( .A(n32776), .B(n32775), .Z(n32809) );
  XNOR U33615 ( .A(n32809), .B(sreg[1813]), .Z(n32811) );
  NAND U33616 ( .A(n32768), .B(sreg[1812]), .Z(n32772) );
  OR U33617 ( .A(n32770), .B(n32769), .Z(n32771) );
  AND U33618 ( .A(n32772), .B(n32771), .Z(n32810) );
  XOR U33619 ( .A(n32811), .B(n32810), .Z(c[1813]) );
  NANDN U33620 ( .A(n32774), .B(n32773), .Z(n32778) );
  NAND U33621 ( .A(n32776), .B(n32775), .Z(n32777) );
  NAND U33622 ( .A(n32778), .B(n32777), .Z(n32817) );
  NAND U33623 ( .A(b[0]), .B(a[798]), .Z(n32779) );
  XNOR U33624 ( .A(b[1]), .B(n32779), .Z(n32781) );
  NAND U33625 ( .A(n129), .B(a[797]), .Z(n32780) );
  AND U33626 ( .A(n32781), .B(n32780), .Z(n32834) );
  XOR U33627 ( .A(a[794]), .B(n42197), .Z(n32823) );
  NANDN U33628 ( .A(n32823), .B(n42173), .Z(n32784) );
  NANDN U33629 ( .A(n32782), .B(n42172), .Z(n32783) );
  NAND U33630 ( .A(n32784), .B(n32783), .Z(n32832) );
  NAND U33631 ( .A(b[7]), .B(a[790]), .Z(n32833) );
  XNOR U33632 ( .A(n32832), .B(n32833), .Z(n32835) );
  XOR U33633 ( .A(n32834), .B(n32835), .Z(n32841) );
  NANDN U33634 ( .A(n32785), .B(n42093), .Z(n32787) );
  XOR U33635 ( .A(n42134), .B(a[796]), .Z(n32826) );
  NANDN U33636 ( .A(n32826), .B(n42095), .Z(n32786) );
  NAND U33637 ( .A(n32787), .B(n32786), .Z(n32839) );
  NANDN U33638 ( .A(n32788), .B(n42231), .Z(n32790) );
  XOR U33639 ( .A(n228), .B(a[792]), .Z(n32829) );
  NANDN U33640 ( .A(n32829), .B(n42234), .Z(n32789) );
  AND U33641 ( .A(n32790), .B(n32789), .Z(n32838) );
  XNOR U33642 ( .A(n32839), .B(n32838), .Z(n32840) );
  XNOR U33643 ( .A(n32841), .B(n32840), .Z(n32845) );
  NANDN U33644 ( .A(n32792), .B(n32791), .Z(n32796) );
  NAND U33645 ( .A(n32794), .B(n32793), .Z(n32795) );
  AND U33646 ( .A(n32796), .B(n32795), .Z(n32844) );
  XOR U33647 ( .A(n32845), .B(n32844), .Z(n32846) );
  NANDN U33648 ( .A(n32798), .B(n32797), .Z(n32802) );
  NANDN U33649 ( .A(n32800), .B(n32799), .Z(n32801) );
  NAND U33650 ( .A(n32802), .B(n32801), .Z(n32847) );
  XOR U33651 ( .A(n32846), .B(n32847), .Z(n32814) );
  OR U33652 ( .A(n32804), .B(n32803), .Z(n32808) );
  NANDN U33653 ( .A(n32806), .B(n32805), .Z(n32807) );
  NAND U33654 ( .A(n32808), .B(n32807), .Z(n32815) );
  XNOR U33655 ( .A(n32814), .B(n32815), .Z(n32816) );
  XNOR U33656 ( .A(n32817), .B(n32816), .Z(n32850) );
  XNOR U33657 ( .A(n32850), .B(sreg[1814]), .Z(n32852) );
  NAND U33658 ( .A(n32809), .B(sreg[1813]), .Z(n32813) );
  OR U33659 ( .A(n32811), .B(n32810), .Z(n32812) );
  AND U33660 ( .A(n32813), .B(n32812), .Z(n32851) );
  XOR U33661 ( .A(n32852), .B(n32851), .Z(c[1814]) );
  NANDN U33662 ( .A(n32815), .B(n32814), .Z(n32819) );
  NAND U33663 ( .A(n32817), .B(n32816), .Z(n32818) );
  NAND U33664 ( .A(n32819), .B(n32818), .Z(n32858) );
  NAND U33665 ( .A(b[0]), .B(a[799]), .Z(n32820) );
  XNOR U33666 ( .A(b[1]), .B(n32820), .Z(n32822) );
  NAND U33667 ( .A(n129), .B(a[798]), .Z(n32821) );
  AND U33668 ( .A(n32822), .B(n32821), .Z(n32875) );
  XOR U33669 ( .A(a[795]), .B(n42197), .Z(n32864) );
  NANDN U33670 ( .A(n32864), .B(n42173), .Z(n32825) );
  NANDN U33671 ( .A(n32823), .B(n42172), .Z(n32824) );
  NAND U33672 ( .A(n32825), .B(n32824), .Z(n32873) );
  NAND U33673 ( .A(b[7]), .B(a[791]), .Z(n32874) );
  XNOR U33674 ( .A(n32873), .B(n32874), .Z(n32876) );
  XOR U33675 ( .A(n32875), .B(n32876), .Z(n32882) );
  NANDN U33676 ( .A(n32826), .B(n42093), .Z(n32828) );
  XOR U33677 ( .A(n42134), .B(a[797]), .Z(n32867) );
  NANDN U33678 ( .A(n32867), .B(n42095), .Z(n32827) );
  NAND U33679 ( .A(n32828), .B(n32827), .Z(n32880) );
  NANDN U33680 ( .A(n32829), .B(n42231), .Z(n32831) );
  XOR U33681 ( .A(n228), .B(a[793]), .Z(n32870) );
  NANDN U33682 ( .A(n32870), .B(n42234), .Z(n32830) );
  AND U33683 ( .A(n32831), .B(n32830), .Z(n32879) );
  XNOR U33684 ( .A(n32880), .B(n32879), .Z(n32881) );
  XNOR U33685 ( .A(n32882), .B(n32881), .Z(n32886) );
  NANDN U33686 ( .A(n32833), .B(n32832), .Z(n32837) );
  NAND U33687 ( .A(n32835), .B(n32834), .Z(n32836) );
  AND U33688 ( .A(n32837), .B(n32836), .Z(n32885) );
  XOR U33689 ( .A(n32886), .B(n32885), .Z(n32887) );
  NANDN U33690 ( .A(n32839), .B(n32838), .Z(n32843) );
  NANDN U33691 ( .A(n32841), .B(n32840), .Z(n32842) );
  NAND U33692 ( .A(n32843), .B(n32842), .Z(n32888) );
  XOR U33693 ( .A(n32887), .B(n32888), .Z(n32855) );
  OR U33694 ( .A(n32845), .B(n32844), .Z(n32849) );
  NANDN U33695 ( .A(n32847), .B(n32846), .Z(n32848) );
  NAND U33696 ( .A(n32849), .B(n32848), .Z(n32856) );
  XNOR U33697 ( .A(n32855), .B(n32856), .Z(n32857) );
  XNOR U33698 ( .A(n32858), .B(n32857), .Z(n32891) );
  XNOR U33699 ( .A(n32891), .B(sreg[1815]), .Z(n32893) );
  NAND U33700 ( .A(n32850), .B(sreg[1814]), .Z(n32854) );
  OR U33701 ( .A(n32852), .B(n32851), .Z(n32853) );
  AND U33702 ( .A(n32854), .B(n32853), .Z(n32892) );
  XOR U33703 ( .A(n32893), .B(n32892), .Z(c[1815]) );
  NANDN U33704 ( .A(n32856), .B(n32855), .Z(n32860) );
  NAND U33705 ( .A(n32858), .B(n32857), .Z(n32859) );
  NAND U33706 ( .A(n32860), .B(n32859), .Z(n32899) );
  NAND U33707 ( .A(b[0]), .B(a[800]), .Z(n32861) );
  XNOR U33708 ( .A(b[1]), .B(n32861), .Z(n32863) );
  NAND U33709 ( .A(n129), .B(a[799]), .Z(n32862) );
  AND U33710 ( .A(n32863), .B(n32862), .Z(n32916) );
  XOR U33711 ( .A(a[796]), .B(n42197), .Z(n32905) );
  NANDN U33712 ( .A(n32905), .B(n42173), .Z(n32866) );
  NANDN U33713 ( .A(n32864), .B(n42172), .Z(n32865) );
  NAND U33714 ( .A(n32866), .B(n32865), .Z(n32914) );
  NAND U33715 ( .A(b[7]), .B(a[792]), .Z(n32915) );
  XNOR U33716 ( .A(n32914), .B(n32915), .Z(n32917) );
  XOR U33717 ( .A(n32916), .B(n32917), .Z(n32923) );
  NANDN U33718 ( .A(n32867), .B(n42093), .Z(n32869) );
  XOR U33719 ( .A(n42134), .B(a[798]), .Z(n32908) );
  NANDN U33720 ( .A(n32908), .B(n42095), .Z(n32868) );
  NAND U33721 ( .A(n32869), .B(n32868), .Z(n32921) );
  NANDN U33722 ( .A(n32870), .B(n42231), .Z(n32872) );
  XOR U33723 ( .A(n228), .B(a[794]), .Z(n32911) );
  NANDN U33724 ( .A(n32911), .B(n42234), .Z(n32871) );
  AND U33725 ( .A(n32872), .B(n32871), .Z(n32920) );
  XNOR U33726 ( .A(n32921), .B(n32920), .Z(n32922) );
  XNOR U33727 ( .A(n32923), .B(n32922), .Z(n32927) );
  NANDN U33728 ( .A(n32874), .B(n32873), .Z(n32878) );
  NAND U33729 ( .A(n32876), .B(n32875), .Z(n32877) );
  AND U33730 ( .A(n32878), .B(n32877), .Z(n32926) );
  XOR U33731 ( .A(n32927), .B(n32926), .Z(n32928) );
  NANDN U33732 ( .A(n32880), .B(n32879), .Z(n32884) );
  NANDN U33733 ( .A(n32882), .B(n32881), .Z(n32883) );
  NAND U33734 ( .A(n32884), .B(n32883), .Z(n32929) );
  XOR U33735 ( .A(n32928), .B(n32929), .Z(n32896) );
  OR U33736 ( .A(n32886), .B(n32885), .Z(n32890) );
  NANDN U33737 ( .A(n32888), .B(n32887), .Z(n32889) );
  NAND U33738 ( .A(n32890), .B(n32889), .Z(n32897) );
  XNOR U33739 ( .A(n32896), .B(n32897), .Z(n32898) );
  XNOR U33740 ( .A(n32899), .B(n32898), .Z(n32932) );
  XNOR U33741 ( .A(n32932), .B(sreg[1816]), .Z(n32934) );
  NAND U33742 ( .A(n32891), .B(sreg[1815]), .Z(n32895) );
  OR U33743 ( .A(n32893), .B(n32892), .Z(n32894) );
  AND U33744 ( .A(n32895), .B(n32894), .Z(n32933) );
  XOR U33745 ( .A(n32934), .B(n32933), .Z(c[1816]) );
  NANDN U33746 ( .A(n32897), .B(n32896), .Z(n32901) );
  NAND U33747 ( .A(n32899), .B(n32898), .Z(n32900) );
  NAND U33748 ( .A(n32901), .B(n32900), .Z(n32940) );
  NAND U33749 ( .A(b[0]), .B(a[801]), .Z(n32902) );
  XNOR U33750 ( .A(b[1]), .B(n32902), .Z(n32904) );
  NAND U33751 ( .A(n129), .B(a[800]), .Z(n32903) );
  AND U33752 ( .A(n32904), .B(n32903), .Z(n32957) );
  XOR U33753 ( .A(a[797]), .B(n42197), .Z(n32946) );
  NANDN U33754 ( .A(n32946), .B(n42173), .Z(n32907) );
  NANDN U33755 ( .A(n32905), .B(n42172), .Z(n32906) );
  NAND U33756 ( .A(n32907), .B(n32906), .Z(n32955) );
  NAND U33757 ( .A(b[7]), .B(a[793]), .Z(n32956) );
  XNOR U33758 ( .A(n32955), .B(n32956), .Z(n32958) );
  XOR U33759 ( .A(n32957), .B(n32958), .Z(n32964) );
  NANDN U33760 ( .A(n32908), .B(n42093), .Z(n32910) );
  XOR U33761 ( .A(n42134), .B(a[799]), .Z(n32949) );
  NANDN U33762 ( .A(n32949), .B(n42095), .Z(n32909) );
  NAND U33763 ( .A(n32910), .B(n32909), .Z(n32962) );
  NANDN U33764 ( .A(n32911), .B(n42231), .Z(n32913) );
  XOR U33765 ( .A(n228), .B(a[795]), .Z(n32952) );
  NANDN U33766 ( .A(n32952), .B(n42234), .Z(n32912) );
  AND U33767 ( .A(n32913), .B(n32912), .Z(n32961) );
  XNOR U33768 ( .A(n32962), .B(n32961), .Z(n32963) );
  XNOR U33769 ( .A(n32964), .B(n32963), .Z(n32968) );
  NANDN U33770 ( .A(n32915), .B(n32914), .Z(n32919) );
  NAND U33771 ( .A(n32917), .B(n32916), .Z(n32918) );
  AND U33772 ( .A(n32919), .B(n32918), .Z(n32967) );
  XOR U33773 ( .A(n32968), .B(n32967), .Z(n32969) );
  NANDN U33774 ( .A(n32921), .B(n32920), .Z(n32925) );
  NANDN U33775 ( .A(n32923), .B(n32922), .Z(n32924) );
  NAND U33776 ( .A(n32925), .B(n32924), .Z(n32970) );
  XOR U33777 ( .A(n32969), .B(n32970), .Z(n32937) );
  OR U33778 ( .A(n32927), .B(n32926), .Z(n32931) );
  NANDN U33779 ( .A(n32929), .B(n32928), .Z(n32930) );
  NAND U33780 ( .A(n32931), .B(n32930), .Z(n32938) );
  XNOR U33781 ( .A(n32937), .B(n32938), .Z(n32939) );
  XNOR U33782 ( .A(n32940), .B(n32939), .Z(n32973) );
  XNOR U33783 ( .A(n32973), .B(sreg[1817]), .Z(n32975) );
  NAND U33784 ( .A(n32932), .B(sreg[1816]), .Z(n32936) );
  OR U33785 ( .A(n32934), .B(n32933), .Z(n32935) );
  AND U33786 ( .A(n32936), .B(n32935), .Z(n32974) );
  XOR U33787 ( .A(n32975), .B(n32974), .Z(c[1817]) );
  NANDN U33788 ( .A(n32938), .B(n32937), .Z(n32942) );
  NAND U33789 ( .A(n32940), .B(n32939), .Z(n32941) );
  NAND U33790 ( .A(n32942), .B(n32941), .Z(n32981) );
  NAND U33791 ( .A(b[0]), .B(a[802]), .Z(n32943) );
  XNOR U33792 ( .A(b[1]), .B(n32943), .Z(n32945) );
  NAND U33793 ( .A(n129), .B(a[801]), .Z(n32944) );
  AND U33794 ( .A(n32945), .B(n32944), .Z(n32998) );
  XOR U33795 ( .A(a[798]), .B(n42197), .Z(n32987) );
  NANDN U33796 ( .A(n32987), .B(n42173), .Z(n32948) );
  NANDN U33797 ( .A(n32946), .B(n42172), .Z(n32947) );
  NAND U33798 ( .A(n32948), .B(n32947), .Z(n32996) );
  NAND U33799 ( .A(b[7]), .B(a[794]), .Z(n32997) );
  XNOR U33800 ( .A(n32996), .B(n32997), .Z(n32999) );
  XOR U33801 ( .A(n32998), .B(n32999), .Z(n33005) );
  NANDN U33802 ( .A(n32949), .B(n42093), .Z(n32951) );
  XOR U33803 ( .A(n42134), .B(a[800]), .Z(n32990) );
  NANDN U33804 ( .A(n32990), .B(n42095), .Z(n32950) );
  NAND U33805 ( .A(n32951), .B(n32950), .Z(n33003) );
  NANDN U33806 ( .A(n32952), .B(n42231), .Z(n32954) );
  XOR U33807 ( .A(n228), .B(a[796]), .Z(n32993) );
  NANDN U33808 ( .A(n32993), .B(n42234), .Z(n32953) );
  AND U33809 ( .A(n32954), .B(n32953), .Z(n33002) );
  XNOR U33810 ( .A(n33003), .B(n33002), .Z(n33004) );
  XNOR U33811 ( .A(n33005), .B(n33004), .Z(n33009) );
  NANDN U33812 ( .A(n32956), .B(n32955), .Z(n32960) );
  NAND U33813 ( .A(n32958), .B(n32957), .Z(n32959) );
  AND U33814 ( .A(n32960), .B(n32959), .Z(n33008) );
  XOR U33815 ( .A(n33009), .B(n33008), .Z(n33010) );
  NANDN U33816 ( .A(n32962), .B(n32961), .Z(n32966) );
  NANDN U33817 ( .A(n32964), .B(n32963), .Z(n32965) );
  NAND U33818 ( .A(n32966), .B(n32965), .Z(n33011) );
  XOR U33819 ( .A(n33010), .B(n33011), .Z(n32978) );
  OR U33820 ( .A(n32968), .B(n32967), .Z(n32972) );
  NANDN U33821 ( .A(n32970), .B(n32969), .Z(n32971) );
  NAND U33822 ( .A(n32972), .B(n32971), .Z(n32979) );
  XNOR U33823 ( .A(n32978), .B(n32979), .Z(n32980) );
  XNOR U33824 ( .A(n32981), .B(n32980), .Z(n33014) );
  XNOR U33825 ( .A(n33014), .B(sreg[1818]), .Z(n33016) );
  NAND U33826 ( .A(n32973), .B(sreg[1817]), .Z(n32977) );
  OR U33827 ( .A(n32975), .B(n32974), .Z(n32976) );
  AND U33828 ( .A(n32977), .B(n32976), .Z(n33015) );
  XOR U33829 ( .A(n33016), .B(n33015), .Z(c[1818]) );
  NANDN U33830 ( .A(n32979), .B(n32978), .Z(n32983) );
  NAND U33831 ( .A(n32981), .B(n32980), .Z(n32982) );
  NAND U33832 ( .A(n32983), .B(n32982), .Z(n33022) );
  NAND U33833 ( .A(b[0]), .B(a[803]), .Z(n32984) );
  XNOR U33834 ( .A(b[1]), .B(n32984), .Z(n32986) );
  NAND U33835 ( .A(n129), .B(a[802]), .Z(n32985) );
  AND U33836 ( .A(n32986), .B(n32985), .Z(n33039) );
  XOR U33837 ( .A(a[799]), .B(n42197), .Z(n33028) );
  NANDN U33838 ( .A(n33028), .B(n42173), .Z(n32989) );
  NANDN U33839 ( .A(n32987), .B(n42172), .Z(n32988) );
  NAND U33840 ( .A(n32989), .B(n32988), .Z(n33037) );
  NAND U33841 ( .A(b[7]), .B(a[795]), .Z(n33038) );
  XNOR U33842 ( .A(n33037), .B(n33038), .Z(n33040) );
  XOR U33843 ( .A(n33039), .B(n33040), .Z(n33046) );
  NANDN U33844 ( .A(n32990), .B(n42093), .Z(n32992) );
  XOR U33845 ( .A(n42134), .B(a[801]), .Z(n33031) );
  NANDN U33846 ( .A(n33031), .B(n42095), .Z(n32991) );
  NAND U33847 ( .A(n32992), .B(n32991), .Z(n33044) );
  NANDN U33848 ( .A(n32993), .B(n42231), .Z(n32995) );
  XOR U33849 ( .A(n228), .B(a[797]), .Z(n33034) );
  NANDN U33850 ( .A(n33034), .B(n42234), .Z(n32994) );
  AND U33851 ( .A(n32995), .B(n32994), .Z(n33043) );
  XNOR U33852 ( .A(n33044), .B(n33043), .Z(n33045) );
  XNOR U33853 ( .A(n33046), .B(n33045), .Z(n33050) );
  NANDN U33854 ( .A(n32997), .B(n32996), .Z(n33001) );
  NAND U33855 ( .A(n32999), .B(n32998), .Z(n33000) );
  AND U33856 ( .A(n33001), .B(n33000), .Z(n33049) );
  XOR U33857 ( .A(n33050), .B(n33049), .Z(n33051) );
  NANDN U33858 ( .A(n33003), .B(n33002), .Z(n33007) );
  NANDN U33859 ( .A(n33005), .B(n33004), .Z(n33006) );
  NAND U33860 ( .A(n33007), .B(n33006), .Z(n33052) );
  XOR U33861 ( .A(n33051), .B(n33052), .Z(n33019) );
  OR U33862 ( .A(n33009), .B(n33008), .Z(n33013) );
  NANDN U33863 ( .A(n33011), .B(n33010), .Z(n33012) );
  NAND U33864 ( .A(n33013), .B(n33012), .Z(n33020) );
  XNOR U33865 ( .A(n33019), .B(n33020), .Z(n33021) );
  XNOR U33866 ( .A(n33022), .B(n33021), .Z(n33055) );
  XNOR U33867 ( .A(n33055), .B(sreg[1819]), .Z(n33057) );
  NAND U33868 ( .A(n33014), .B(sreg[1818]), .Z(n33018) );
  OR U33869 ( .A(n33016), .B(n33015), .Z(n33017) );
  AND U33870 ( .A(n33018), .B(n33017), .Z(n33056) );
  XOR U33871 ( .A(n33057), .B(n33056), .Z(c[1819]) );
  NANDN U33872 ( .A(n33020), .B(n33019), .Z(n33024) );
  NAND U33873 ( .A(n33022), .B(n33021), .Z(n33023) );
  NAND U33874 ( .A(n33024), .B(n33023), .Z(n33063) );
  NAND U33875 ( .A(b[0]), .B(a[804]), .Z(n33025) );
  XNOR U33876 ( .A(b[1]), .B(n33025), .Z(n33027) );
  NAND U33877 ( .A(n129), .B(a[803]), .Z(n33026) );
  AND U33878 ( .A(n33027), .B(n33026), .Z(n33080) );
  XOR U33879 ( .A(a[800]), .B(n42197), .Z(n33069) );
  NANDN U33880 ( .A(n33069), .B(n42173), .Z(n33030) );
  NANDN U33881 ( .A(n33028), .B(n42172), .Z(n33029) );
  NAND U33882 ( .A(n33030), .B(n33029), .Z(n33078) );
  NAND U33883 ( .A(b[7]), .B(a[796]), .Z(n33079) );
  XNOR U33884 ( .A(n33078), .B(n33079), .Z(n33081) );
  XOR U33885 ( .A(n33080), .B(n33081), .Z(n33087) );
  NANDN U33886 ( .A(n33031), .B(n42093), .Z(n33033) );
  XOR U33887 ( .A(n42134), .B(a[802]), .Z(n33072) );
  NANDN U33888 ( .A(n33072), .B(n42095), .Z(n33032) );
  NAND U33889 ( .A(n33033), .B(n33032), .Z(n33085) );
  NANDN U33890 ( .A(n33034), .B(n42231), .Z(n33036) );
  XOR U33891 ( .A(n228), .B(a[798]), .Z(n33075) );
  NANDN U33892 ( .A(n33075), .B(n42234), .Z(n33035) );
  AND U33893 ( .A(n33036), .B(n33035), .Z(n33084) );
  XNOR U33894 ( .A(n33085), .B(n33084), .Z(n33086) );
  XNOR U33895 ( .A(n33087), .B(n33086), .Z(n33091) );
  NANDN U33896 ( .A(n33038), .B(n33037), .Z(n33042) );
  NAND U33897 ( .A(n33040), .B(n33039), .Z(n33041) );
  AND U33898 ( .A(n33042), .B(n33041), .Z(n33090) );
  XOR U33899 ( .A(n33091), .B(n33090), .Z(n33092) );
  NANDN U33900 ( .A(n33044), .B(n33043), .Z(n33048) );
  NANDN U33901 ( .A(n33046), .B(n33045), .Z(n33047) );
  NAND U33902 ( .A(n33048), .B(n33047), .Z(n33093) );
  XOR U33903 ( .A(n33092), .B(n33093), .Z(n33060) );
  OR U33904 ( .A(n33050), .B(n33049), .Z(n33054) );
  NANDN U33905 ( .A(n33052), .B(n33051), .Z(n33053) );
  NAND U33906 ( .A(n33054), .B(n33053), .Z(n33061) );
  XNOR U33907 ( .A(n33060), .B(n33061), .Z(n33062) );
  XNOR U33908 ( .A(n33063), .B(n33062), .Z(n33096) );
  XNOR U33909 ( .A(n33096), .B(sreg[1820]), .Z(n33098) );
  NAND U33910 ( .A(n33055), .B(sreg[1819]), .Z(n33059) );
  OR U33911 ( .A(n33057), .B(n33056), .Z(n33058) );
  AND U33912 ( .A(n33059), .B(n33058), .Z(n33097) );
  XOR U33913 ( .A(n33098), .B(n33097), .Z(c[1820]) );
  NANDN U33914 ( .A(n33061), .B(n33060), .Z(n33065) );
  NAND U33915 ( .A(n33063), .B(n33062), .Z(n33064) );
  NAND U33916 ( .A(n33065), .B(n33064), .Z(n33104) );
  NAND U33917 ( .A(b[0]), .B(a[805]), .Z(n33066) );
  XNOR U33918 ( .A(b[1]), .B(n33066), .Z(n33068) );
  NAND U33919 ( .A(n130), .B(a[804]), .Z(n33067) );
  AND U33920 ( .A(n33068), .B(n33067), .Z(n33121) );
  XOR U33921 ( .A(a[801]), .B(n42197), .Z(n33110) );
  NANDN U33922 ( .A(n33110), .B(n42173), .Z(n33071) );
  NANDN U33923 ( .A(n33069), .B(n42172), .Z(n33070) );
  NAND U33924 ( .A(n33071), .B(n33070), .Z(n33119) );
  NAND U33925 ( .A(b[7]), .B(a[797]), .Z(n33120) );
  XNOR U33926 ( .A(n33119), .B(n33120), .Z(n33122) );
  XOR U33927 ( .A(n33121), .B(n33122), .Z(n33128) );
  NANDN U33928 ( .A(n33072), .B(n42093), .Z(n33074) );
  XOR U33929 ( .A(n42134), .B(a[803]), .Z(n33113) );
  NANDN U33930 ( .A(n33113), .B(n42095), .Z(n33073) );
  NAND U33931 ( .A(n33074), .B(n33073), .Z(n33126) );
  NANDN U33932 ( .A(n33075), .B(n42231), .Z(n33077) );
  XOR U33933 ( .A(n228), .B(a[799]), .Z(n33116) );
  NANDN U33934 ( .A(n33116), .B(n42234), .Z(n33076) );
  AND U33935 ( .A(n33077), .B(n33076), .Z(n33125) );
  XNOR U33936 ( .A(n33126), .B(n33125), .Z(n33127) );
  XNOR U33937 ( .A(n33128), .B(n33127), .Z(n33132) );
  NANDN U33938 ( .A(n33079), .B(n33078), .Z(n33083) );
  NAND U33939 ( .A(n33081), .B(n33080), .Z(n33082) );
  AND U33940 ( .A(n33083), .B(n33082), .Z(n33131) );
  XOR U33941 ( .A(n33132), .B(n33131), .Z(n33133) );
  NANDN U33942 ( .A(n33085), .B(n33084), .Z(n33089) );
  NANDN U33943 ( .A(n33087), .B(n33086), .Z(n33088) );
  NAND U33944 ( .A(n33089), .B(n33088), .Z(n33134) );
  XOR U33945 ( .A(n33133), .B(n33134), .Z(n33101) );
  OR U33946 ( .A(n33091), .B(n33090), .Z(n33095) );
  NANDN U33947 ( .A(n33093), .B(n33092), .Z(n33094) );
  NAND U33948 ( .A(n33095), .B(n33094), .Z(n33102) );
  XNOR U33949 ( .A(n33101), .B(n33102), .Z(n33103) );
  XNOR U33950 ( .A(n33104), .B(n33103), .Z(n33137) );
  XNOR U33951 ( .A(n33137), .B(sreg[1821]), .Z(n33139) );
  NAND U33952 ( .A(n33096), .B(sreg[1820]), .Z(n33100) );
  OR U33953 ( .A(n33098), .B(n33097), .Z(n33099) );
  AND U33954 ( .A(n33100), .B(n33099), .Z(n33138) );
  XOR U33955 ( .A(n33139), .B(n33138), .Z(c[1821]) );
  NANDN U33956 ( .A(n33102), .B(n33101), .Z(n33106) );
  NAND U33957 ( .A(n33104), .B(n33103), .Z(n33105) );
  NAND U33958 ( .A(n33106), .B(n33105), .Z(n33145) );
  NAND U33959 ( .A(b[0]), .B(a[806]), .Z(n33107) );
  XNOR U33960 ( .A(b[1]), .B(n33107), .Z(n33109) );
  NAND U33961 ( .A(n130), .B(a[805]), .Z(n33108) );
  AND U33962 ( .A(n33109), .B(n33108), .Z(n33162) );
  XOR U33963 ( .A(a[802]), .B(n42197), .Z(n33151) );
  NANDN U33964 ( .A(n33151), .B(n42173), .Z(n33112) );
  NANDN U33965 ( .A(n33110), .B(n42172), .Z(n33111) );
  NAND U33966 ( .A(n33112), .B(n33111), .Z(n33160) );
  NAND U33967 ( .A(b[7]), .B(a[798]), .Z(n33161) );
  XNOR U33968 ( .A(n33160), .B(n33161), .Z(n33163) );
  XOR U33969 ( .A(n33162), .B(n33163), .Z(n33169) );
  NANDN U33970 ( .A(n33113), .B(n42093), .Z(n33115) );
  XOR U33971 ( .A(n42134), .B(a[804]), .Z(n33154) );
  NANDN U33972 ( .A(n33154), .B(n42095), .Z(n33114) );
  NAND U33973 ( .A(n33115), .B(n33114), .Z(n33167) );
  NANDN U33974 ( .A(n33116), .B(n42231), .Z(n33118) );
  XOR U33975 ( .A(n228), .B(a[800]), .Z(n33157) );
  NANDN U33976 ( .A(n33157), .B(n42234), .Z(n33117) );
  AND U33977 ( .A(n33118), .B(n33117), .Z(n33166) );
  XNOR U33978 ( .A(n33167), .B(n33166), .Z(n33168) );
  XNOR U33979 ( .A(n33169), .B(n33168), .Z(n33173) );
  NANDN U33980 ( .A(n33120), .B(n33119), .Z(n33124) );
  NAND U33981 ( .A(n33122), .B(n33121), .Z(n33123) );
  AND U33982 ( .A(n33124), .B(n33123), .Z(n33172) );
  XOR U33983 ( .A(n33173), .B(n33172), .Z(n33174) );
  NANDN U33984 ( .A(n33126), .B(n33125), .Z(n33130) );
  NANDN U33985 ( .A(n33128), .B(n33127), .Z(n33129) );
  NAND U33986 ( .A(n33130), .B(n33129), .Z(n33175) );
  XOR U33987 ( .A(n33174), .B(n33175), .Z(n33142) );
  OR U33988 ( .A(n33132), .B(n33131), .Z(n33136) );
  NANDN U33989 ( .A(n33134), .B(n33133), .Z(n33135) );
  NAND U33990 ( .A(n33136), .B(n33135), .Z(n33143) );
  XNOR U33991 ( .A(n33142), .B(n33143), .Z(n33144) );
  XNOR U33992 ( .A(n33145), .B(n33144), .Z(n33178) );
  XNOR U33993 ( .A(n33178), .B(sreg[1822]), .Z(n33180) );
  NAND U33994 ( .A(n33137), .B(sreg[1821]), .Z(n33141) );
  OR U33995 ( .A(n33139), .B(n33138), .Z(n33140) );
  AND U33996 ( .A(n33141), .B(n33140), .Z(n33179) );
  XOR U33997 ( .A(n33180), .B(n33179), .Z(c[1822]) );
  NANDN U33998 ( .A(n33143), .B(n33142), .Z(n33147) );
  NAND U33999 ( .A(n33145), .B(n33144), .Z(n33146) );
  NAND U34000 ( .A(n33147), .B(n33146), .Z(n33186) );
  NAND U34001 ( .A(b[0]), .B(a[807]), .Z(n33148) );
  XNOR U34002 ( .A(b[1]), .B(n33148), .Z(n33150) );
  NAND U34003 ( .A(n130), .B(a[806]), .Z(n33149) );
  AND U34004 ( .A(n33150), .B(n33149), .Z(n33203) );
  XOR U34005 ( .A(a[803]), .B(n42197), .Z(n33192) );
  NANDN U34006 ( .A(n33192), .B(n42173), .Z(n33153) );
  NANDN U34007 ( .A(n33151), .B(n42172), .Z(n33152) );
  NAND U34008 ( .A(n33153), .B(n33152), .Z(n33201) );
  NAND U34009 ( .A(b[7]), .B(a[799]), .Z(n33202) );
  XNOR U34010 ( .A(n33201), .B(n33202), .Z(n33204) );
  XOR U34011 ( .A(n33203), .B(n33204), .Z(n33210) );
  NANDN U34012 ( .A(n33154), .B(n42093), .Z(n33156) );
  XOR U34013 ( .A(n42134), .B(a[805]), .Z(n33195) );
  NANDN U34014 ( .A(n33195), .B(n42095), .Z(n33155) );
  NAND U34015 ( .A(n33156), .B(n33155), .Z(n33208) );
  NANDN U34016 ( .A(n33157), .B(n42231), .Z(n33159) );
  XOR U34017 ( .A(n228), .B(a[801]), .Z(n33198) );
  NANDN U34018 ( .A(n33198), .B(n42234), .Z(n33158) );
  AND U34019 ( .A(n33159), .B(n33158), .Z(n33207) );
  XNOR U34020 ( .A(n33208), .B(n33207), .Z(n33209) );
  XNOR U34021 ( .A(n33210), .B(n33209), .Z(n33214) );
  NANDN U34022 ( .A(n33161), .B(n33160), .Z(n33165) );
  NAND U34023 ( .A(n33163), .B(n33162), .Z(n33164) );
  AND U34024 ( .A(n33165), .B(n33164), .Z(n33213) );
  XOR U34025 ( .A(n33214), .B(n33213), .Z(n33215) );
  NANDN U34026 ( .A(n33167), .B(n33166), .Z(n33171) );
  NANDN U34027 ( .A(n33169), .B(n33168), .Z(n33170) );
  NAND U34028 ( .A(n33171), .B(n33170), .Z(n33216) );
  XOR U34029 ( .A(n33215), .B(n33216), .Z(n33183) );
  OR U34030 ( .A(n33173), .B(n33172), .Z(n33177) );
  NANDN U34031 ( .A(n33175), .B(n33174), .Z(n33176) );
  NAND U34032 ( .A(n33177), .B(n33176), .Z(n33184) );
  XNOR U34033 ( .A(n33183), .B(n33184), .Z(n33185) );
  XNOR U34034 ( .A(n33186), .B(n33185), .Z(n33219) );
  XNOR U34035 ( .A(n33219), .B(sreg[1823]), .Z(n33221) );
  NAND U34036 ( .A(n33178), .B(sreg[1822]), .Z(n33182) );
  OR U34037 ( .A(n33180), .B(n33179), .Z(n33181) );
  AND U34038 ( .A(n33182), .B(n33181), .Z(n33220) );
  XOR U34039 ( .A(n33221), .B(n33220), .Z(c[1823]) );
  NANDN U34040 ( .A(n33184), .B(n33183), .Z(n33188) );
  NAND U34041 ( .A(n33186), .B(n33185), .Z(n33187) );
  NAND U34042 ( .A(n33188), .B(n33187), .Z(n33227) );
  NAND U34043 ( .A(b[0]), .B(a[808]), .Z(n33189) );
  XNOR U34044 ( .A(b[1]), .B(n33189), .Z(n33191) );
  NAND U34045 ( .A(n130), .B(a[807]), .Z(n33190) );
  AND U34046 ( .A(n33191), .B(n33190), .Z(n33244) );
  XOR U34047 ( .A(a[804]), .B(n42197), .Z(n33233) );
  NANDN U34048 ( .A(n33233), .B(n42173), .Z(n33194) );
  NANDN U34049 ( .A(n33192), .B(n42172), .Z(n33193) );
  NAND U34050 ( .A(n33194), .B(n33193), .Z(n33242) );
  NAND U34051 ( .A(b[7]), .B(a[800]), .Z(n33243) );
  XNOR U34052 ( .A(n33242), .B(n33243), .Z(n33245) );
  XOR U34053 ( .A(n33244), .B(n33245), .Z(n33251) );
  NANDN U34054 ( .A(n33195), .B(n42093), .Z(n33197) );
  XOR U34055 ( .A(n42134), .B(a[806]), .Z(n33236) );
  NANDN U34056 ( .A(n33236), .B(n42095), .Z(n33196) );
  NAND U34057 ( .A(n33197), .B(n33196), .Z(n33249) );
  NANDN U34058 ( .A(n33198), .B(n42231), .Z(n33200) );
  XOR U34059 ( .A(n228), .B(a[802]), .Z(n33239) );
  NANDN U34060 ( .A(n33239), .B(n42234), .Z(n33199) );
  AND U34061 ( .A(n33200), .B(n33199), .Z(n33248) );
  XNOR U34062 ( .A(n33249), .B(n33248), .Z(n33250) );
  XNOR U34063 ( .A(n33251), .B(n33250), .Z(n33255) );
  NANDN U34064 ( .A(n33202), .B(n33201), .Z(n33206) );
  NAND U34065 ( .A(n33204), .B(n33203), .Z(n33205) );
  AND U34066 ( .A(n33206), .B(n33205), .Z(n33254) );
  XOR U34067 ( .A(n33255), .B(n33254), .Z(n33256) );
  NANDN U34068 ( .A(n33208), .B(n33207), .Z(n33212) );
  NANDN U34069 ( .A(n33210), .B(n33209), .Z(n33211) );
  NAND U34070 ( .A(n33212), .B(n33211), .Z(n33257) );
  XOR U34071 ( .A(n33256), .B(n33257), .Z(n33224) );
  OR U34072 ( .A(n33214), .B(n33213), .Z(n33218) );
  NANDN U34073 ( .A(n33216), .B(n33215), .Z(n33217) );
  NAND U34074 ( .A(n33218), .B(n33217), .Z(n33225) );
  XNOR U34075 ( .A(n33224), .B(n33225), .Z(n33226) );
  XNOR U34076 ( .A(n33227), .B(n33226), .Z(n33260) );
  XNOR U34077 ( .A(n33260), .B(sreg[1824]), .Z(n33262) );
  NAND U34078 ( .A(n33219), .B(sreg[1823]), .Z(n33223) );
  OR U34079 ( .A(n33221), .B(n33220), .Z(n33222) );
  AND U34080 ( .A(n33223), .B(n33222), .Z(n33261) );
  XOR U34081 ( .A(n33262), .B(n33261), .Z(c[1824]) );
  NANDN U34082 ( .A(n33225), .B(n33224), .Z(n33229) );
  NAND U34083 ( .A(n33227), .B(n33226), .Z(n33228) );
  NAND U34084 ( .A(n33229), .B(n33228), .Z(n33268) );
  NAND U34085 ( .A(b[0]), .B(a[809]), .Z(n33230) );
  XNOR U34086 ( .A(b[1]), .B(n33230), .Z(n33232) );
  NAND U34087 ( .A(n130), .B(a[808]), .Z(n33231) );
  AND U34088 ( .A(n33232), .B(n33231), .Z(n33285) );
  XOR U34089 ( .A(a[805]), .B(n42197), .Z(n33274) );
  NANDN U34090 ( .A(n33274), .B(n42173), .Z(n33235) );
  NANDN U34091 ( .A(n33233), .B(n42172), .Z(n33234) );
  NAND U34092 ( .A(n33235), .B(n33234), .Z(n33283) );
  NAND U34093 ( .A(b[7]), .B(a[801]), .Z(n33284) );
  XNOR U34094 ( .A(n33283), .B(n33284), .Z(n33286) );
  XOR U34095 ( .A(n33285), .B(n33286), .Z(n33292) );
  NANDN U34096 ( .A(n33236), .B(n42093), .Z(n33238) );
  XOR U34097 ( .A(n42134), .B(a[807]), .Z(n33277) );
  NANDN U34098 ( .A(n33277), .B(n42095), .Z(n33237) );
  NAND U34099 ( .A(n33238), .B(n33237), .Z(n33290) );
  NANDN U34100 ( .A(n33239), .B(n42231), .Z(n33241) );
  XOR U34101 ( .A(n229), .B(a[803]), .Z(n33280) );
  NANDN U34102 ( .A(n33280), .B(n42234), .Z(n33240) );
  AND U34103 ( .A(n33241), .B(n33240), .Z(n33289) );
  XNOR U34104 ( .A(n33290), .B(n33289), .Z(n33291) );
  XNOR U34105 ( .A(n33292), .B(n33291), .Z(n33296) );
  NANDN U34106 ( .A(n33243), .B(n33242), .Z(n33247) );
  NAND U34107 ( .A(n33245), .B(n33244), .Z(n33246) );
  AND U34108 ( .A(n33247), .B(n33246), .Z(n33295) );
  XOR U34109 ( .A(n33296), .B(n33295), .Z(n33297) );
  NANDN U34110 ( .A(n33249), .B(n33248), .Z(n33253) );
  NANDN U34111 ( .A(n33251), .B(n33250), .Z(n33252) );
  NAND U34112 ( .A(n33253), .B(n33252), .Z(n33298) );
  XOR U34113 ( .A(n33297), .B(n33298), .Z(n33265) );
  OR U34114 ( .A(n33255), .B(n33254), .Z(n33259) );
  NANDN U34115 ( .A(n33257), .B(n33256), .Z(n33258) );
  NAND U34116 ( .A(n33259), .B(n33258), .Z(n33266) );
  XNOR U34117 ( .A(n33265), .B(n33266), .Z(n33267) );
  XNOR U34118 ( .A(n33268), .B(n33267), .Z(n33301) );
  XNOR U34119 ( .A(n33301), .B(sreg[1825]), .Z(n33303) );
  NAND U34120 ( .A(n33260), .B(sreg[1824]), .Z(n33264) );
  OR U34121 ( .A(n33262), .B(n33261), .Z(n33263) );
  AND U34122 ( .A(n33264), .B(n33263), .Z(n33302) );
  XOR U34123 ( .A(n33303), .B(n33302), .Z(c[1825]) );
  NANDN U34124 ( .A(n33266), .B(n33265), .Z(n33270) );
  NAND U34125 ( .A(n33268), .B(n33267), .Z(n33269) );
  NAND U34126 ( .A(n33270), .B(n33269), .Z(n33309) );
  NAND U34127 ( .A(b[0]), .B(a[810]), .Z(n33271) );
  XNOR U34128 ( .A(b[1]), .B(n33271), .Z(n33273) );
  NAND U34129 ( .A(n130), .B(a[809]), .Z(n33272) );
  AND U34130 ( .A(n33273), .B(n33272), .Z(n33326) );
  XOR U34131 ( .A(a[806]), .B(n42197), .Z(n33315) );
  NANDN U34132 ( .A(n33315), .B(n42173), .Z(n33276) );
  NANDN U34133 ( .A(n33274), .B(n42172), .Z(n33275) );
  NAND U34134 ( .A(n33276), .B(n33275), .Z(n33324) );
  NAND U34135 ( .A(b[7]), .B(a[802]), .Z(n33325) );
  XNOR U34136 ( .A(n33324), .B(n33325), .Z(n33327) );
  XOR U34137 ( .A(n33326), .B(n33327), .Z(n33333) );
  NANDN U34138 ( .A(n33277), .B(n42093), .Z(n33279) );
  XOR U34139 ( .A(n42134), .B(a[808]), .Z(n33318) );
  NANDN U34140 ( .A(n33318), .B(n42095), .Z(n33278) );
  NAND U34141 ( .A(n33279), .B(n33278), .Z(n33331) );
  NANDN U34142 ( .A(n33280), .B(n42231), .Z(n33282) );
  XOR U34143 ( .A(n229), .B(a[804]), .Z(n33321) );
  NANDN U34144 ( .A(n33321), .B(n42234), .Z(n33281) );
  AND U34145 ( .A(n33282), .B(n33281), .Z(n33330) );
  XNOR U34146 ( .A(n33331), .B(n33330), .Z(n33332) );
  XNOR U34147 ( .A(n33333), .B(n33332), .Z(n33337) );
  NANDN U34148 ( .A(n33284), .B(n33283), .Z(n33288) );
  NAND U34149 ( .A(n33286), .B(n33285), .Z(n33287) );
  AND U34150 ( .A(n33288), .B(n33287), .Z(n33336) );
  XOR U34151 ( .A(n33337), .B(n33336), .Z(n33338) );
  NANDN U34152 ( .A(n33290), .B(n33289), .Z(n33294) );
  NANDN U34153 ( .A(n33292), .B(n33291), .Z(n33293) );
  NAND U34154 ( .A(n33294), .B(n33293), .Z(n33339) );
  XOR U34155 ( .A(n33338), .B(n33339), .Z(n33306) );
  OR U34156 ( .A(n33296), .B(n33295), .Z(n33300) );
  NANDN U34157 ( .A(n33298), .B(n33297), .Z(n33299) );
  NAND U34158 ( .A(n33300), .B(n33299), .Z(n33307) );
  XNOR U34159 ( .A(n33306), .B(n33307), .Z(n33308) );
  XNOR U34160 ( .A(n33309), .B(n33308), .Z(n33342) );
  XNOR U34161 ( .A(n33342), .B(sreg[1826]), .Z(n33344) );
  NAND U34162 ( .A(n33301), .B(sreg[1825]), .Z(n33305) );
  OR U34163 ( .A(n33303), .B(n33302), .Z(n33304) );
  AND U34164 ( .A(n33305), .B(n33304), .Z(n33343) );
  XOR U34165 ( .A(n33344), .B(n33343), .Z(c[1826]) );
  NANDN U34166 ( .A(n33307), .B(n33306), .Z(n33311) );
  NAND U34167 ( .A(n33309), .B(n33308), .Z(n33310) );
  NAND U34168 ( .A(n33311), .B(n33310), .Z(n33350) );
  NAND U34169 ( .A(b[0]), .B(a[811]), .Z(n33312) );
  XNOR U34170 ( .A(b[1]), .B(n33312), .Z(n33314) );
  NAND U34171 ( .A(n130), .B(a[810]), .Z(n33313) );
  AND U34172 ( .A(n33314), .B(n33313), .Z(n33367) );
  XOR U34173 ( .A(a[807]), .B(n42197), .Z(n33356) );
  NANDN U34174 ( .A(n33356), .B(n42173), .Z(n33317) );
  NANDN U34175 ( .A(n33315), .B(n42172), .Z(n33316) );
  NAND U34176 ( .A(n33317), .B(n33316), .Z(n33365) );
  NAND U34177 ( .A(b[7]), .B(a[803]), .Z(n33366) );
  XNOR U34178 ( .A(n33365), .B(n33366), .Z(n33368) );
  XOR U34179 ( .A(n33367), .B(n33368), .Z(n33374) );
  NANDN U34180 ( .A(n33318), .B(n42093), .Z(n33320) );
  XOR U34181 ( .A(n42134), .B(a[809]), .Z(n33359) );
  NANDN U34182 ( .A(n33359), .B(n42095), .Z(n33319) );
  NAND U34183 ( .A(n33320), .B(n33319), .Z(n33372) );
  NANDN U34184 ( .A(n33321), .B(n42231), .Z(n33323) );
  XOR U34185 ( .A(n229), .B(a[805]), .Z(n33362) );
  NANDN U34186 ( .A(n33362), .B(n42234), .Z(n33322) );
  AND U34187 ( .A(n33323), .B(n33322), .Z(n33371) );
  XNOR U34188 ( .A(n33372), .B(n33371), .Z(n33373) );
  XNOR U34189 ( .A(n33374), .B(n33373), .Z(n33378) );
  NANDN U34190 ( .A(n33325), .B(n33324), .Z(n33329) );
  NAND U34191 ( .A(n33327), .B(n33326), .Z(n33328) );
  AND U34192 ( .A(n33329), .B(n33328), .Z(n33377) );
  XOR U34193 ( .A(n33378), .B(n33377), .Z(n33379) );
  NANDN U34194 ( .A(n33331), .B(n33330), .Z(n33335) );
  NANDN U34195 ( .A(n33333), .B(n33332), .Z(n33334) );
  NAND U34196 ( .A(n33335), .B(n33334), .Z(n33380) );
  XOR U34197 ( .A(n33379), .B(n33380), .Z(n33347) );
  OR U34198 ( .A(n33337), .B(n33336), .Z(n33341) );
  NANDN U34199 ( .A(n33339), .B(n33338), .Z(n33340) );
  NAND U34200 ( .A(n33341), .B(n33340), .Z(n33348) );
  XNOR U34201 ( .A(n33347), .B(n33348), .Z(n33349) );
  XNOR U34202 ( .A(n33350), .B(n33349), .Z(n33383) );
  XNOR U34203 ( .A(n33383), .B(sreg[1827]), .Z(n33385) );
  NAND U34204 ( .A(n33342), .B(sreg[1826]), .Z(n33346) );
  OR U34205 ( .A(n33344), .B(n33343), .Z(n33345) );
  AND U34206 ( .A(n33346), .B(n33345), .Z(n33384) );
  XOR U34207 ( .A(n33385), .B(n33384), .Z(c[1827]) );
  NANDN U34208 ( .A(n33348), .B(n33347), .Z(n33352) );
  NAND U34209 ( .A(n33350), .B(n33349), .Z(n33351) );
  NAND U34210 ( .A(n33352), .B(n33351), .Z(n33391) );
  NAND U34211 ( .A(b[0]), .B(a[812]), .Z(n33353) );
  XNOR U34212 ( .A(b[1]), .B(n33353), .Z(n33355) );
  NAND U34213 ( .A(n131), .B(a[811]), .Z(n33354) );
  AND U34214 ( .A(n33355), .B(n33354), .Z(n33408) );
  XOR U34215 ( .A(a[808]), .B(n42197), .Z(n33397) );
  NANDN U34216 ( .A(n33397), .B(n42173), .Z(n33358) );
  NANDN U34217 ( .A(n33356), .B(n42172), .Z(n33357) );
  NAND U34218 ( .A(n33358), .B(n33357), .Z(n33406) );
  NAND U34219 ( .A(b[7]), .B(a[804]), .Z(n33407) );
  XNOR U34220 ( .A(n33406), .B(n33407), .Z(n33409) );
  XOR U34221 ( .A(n33408), .B(n33409), .Z(n33415) );
  NANDN U34222 ( .A(n33359), .B(n42093), .Z(n33361) );
  XOR U34223 ( .A(n42134), .B(a[810]), .Z(n33400) );
  NANDN U34224 ( .A(n33400), .B(n42095), .Z(n33360) );
  NAND U34225 ( .A(n33361), .B(n33360), .Z(n33413) );
  NANDN U34226 ( .A(n33362), .B(n42231), .Z(n33364) );
  XOR U34227 ( .A(n229), .B(a[806]), .Z(n33403) );
  NANDN U34228 ( .A(n33403), .B(n42234), .Z(n33363) );
  AND U34229 ( .A(n33364), .B(n33363), .Z(n33412) );
  XNOR U34230 ( .A(n33413), .B(n33412), .Z(n33414) );
  XNOR U34231 ( .A(n33415), .B(n33414), .Z(n33419) );
  NANDN U34232 ( .A(n33366), .B(n33365), .Z(n33370) );
  NAND U34233 ( .A(n33368), .B(n33367), .Z(n33369) );
  AND U34234 ( .A(n33370), .B(n33369), .Z(n33418) );
  XOR U34235 ( .A(n33419), .B(n33418), .Z(n33420) );
  NANDN U34236 ( .A(n33372), .B(n33371), .Z(n33376) );
  NANDN U34237 ( .A(n33374), .B(n33373), .Z(n33375) );
  NAND U34238 ( .A(n33376), .B(n33375), .Z(n33421) );
  XOR U34239 ( .A(n33420), .B(n33421), .Z(n33388) );
  OR U34240 ( .A(n33378), .B(n33377), .Z(n33382) );
  NANDN U34241 ( .A(n33380), .B(n33379), .Z(n33381) );
  NAND U34242 ( .A(n33382), .B(n33381), .Z(n33389) );
  XNOR U34243 ( .A(n33388), .B(n33389), .Z(n33390) );
  XNOR U34244 ( .A(n33391), .B(n33390), .Z(n33424) );
  XNOR U34245 ( .A(n33424), .B(sreg[1828]), .Z(n33426) );
  NAND U34246 ( .A(n33383), .B(sreg[1827]), .Z(n33387) );
  OR U34247 ( .A(n33385), .B(n33384), .Z(n33386) );
  AND U34248 ( .A(n33387), .B(n33386), .Z(n33425) );
  XOR U34249 ( .A(n33426), .B(n33425), .Z(c[1828]) );
  NANDN U34250 ( .A(n33389), .B(n33388), .Z(n33393) );
  NAND U34251 ( .A(n33391), .B(n33390), .Z(n33392) );
  NAND U34252 ( .A(n33393), .B(n33392), .Z(n33432) );
  NAND U34253 ( .A(b[0]), .B(a[813]), .Z(n33394) );
  XNOR U34254 ( .A(b[1]), .B(n33394), .Z(n33396) );
  NAND U34255 ( .A(n131), .B(a[812]), .Z(n33395) );
  AND U34256 ( .A(n33396), .B(n33395), .Z(n33449) );
  XOR U34257 ( .A(a[809]), .B(n42197), .Z(n33438) );
  NANDN U34258 ( .A(n33438), .B(n42173), .Z(n33399) );
  NANDN U34259 ( .A(n33397), .B(n42172), .Z(n33398) );
  NAND U34260 ( .A(n33399), .B(n33398), .Z(n33447) );
  NAND U34261 ( .A(b[7]), .B(a[805]), .Z(n33448) );
  XNOR U34262 ( .A(n33447), .B(n33448), .Z(n33450) );
  XOR U34263 ( .A(n33449), .B(n33450), .Z(n33456) );
  NANDN U34264 ( .A(n33400), .B(n42093), .Z(n33402) );
  XOR U34265 ( .A(n42134), .B(a[811]), .Z(n33441) );
  NANDN U34266 ( .A(n33441), .B(n42095), .Z(n33401) );
  NAND U34267 ( .A(n33402), .B(n33401), .Z(n33454) );
  NANDN U34268 ( .A(n33403), .B(n42231), .Z(n33405) );
  XOR U34269 ( .A(n229), .B(a[807]), .Z(n33444) );
  NANDN U34270 ( .A(n33444), .B(n42234), .Z(n33404) );
  AND U34271 ( .A(n33405), .B(n33404), .Z(n33453) );
  XNOR U34272 ( .A(n33454), .B(n33453), .Z(n33455) );
  XNOR U34273 ( .A(n33456), .B(n33455), .Z(n33460) );
  NANDN U34274 ( .A(n33407), .B(n33406), .Z(n33411) );
  NAND U34275 ( .A(n33409), .B(n33408), .Z(n33410) );
  AND U34276 ( .A(n33411), .B(n33410), .Z(n33459) );
  XOR U34277 ( .A(n33460), .B(n33459), .Z(n33461) );
  NANDN U34278 ( .A(n33413), .B(n33412), .Z(n33417) );
  NANDN U34279 ( .A(n33415), .B(n33414), .Z(n33416) );
  NAND U34280 ( .A(n33417), .B(n33416), .Z(n33462) );
  XOR U34281 ( .A(n33461), .B(n33462), .Z(n33429) );
  OR U34282 ( .A(n33419), .B(n33418), .Z(n33423) );
  NANDN U34283 ( .A(n33421), .B(n33420), .Z(n33422) );
  NAND U34284 ( .A(n33423), .B(n33422), .Z(n33430) );
  XNOR U34285 ( .A(n33429), .B(n33430), .Z(n33431) );
  XNOR U34286 ( .A(n33432), .B(n33431), .Z(n33465) );
  XNOR U34287 ( .A(n33465), .B(sreg[1829]), .Z(n33467) );
  NAND U34288 ( .A(n33424), .B(sreg[1828]), .Z(n33428) );
  OR U34289 ( .A(n33426), .B(n33425), .Z(n33427) );
  AND U34290 ( .A(n33428), .B(n33427), .Z(n33466) );
  XOR U34291 ( .A(n33467), .B(n33466), .Z(c[1829]) );
  NANDN U34292 ( .A(n33430), .B(n33429), .Z(n33434) );
  NAND U34293 ( .A(n33432), .B(n33431), .Z(n33433) );
  NAND U34294 ( .A(n33434), .B(n33433), .Z(n33473) );
  NAND U34295 ( .A(b[0]), .B(a[814]), .Z(n33435) );
  XNOR U34296 ( .A(b[1]), .B(n33435), .Z(n33437) );
  NAND U34297 ( .A(n131), .B(a[813]), .Z(n33436) );
  AND U34298 ( .A(n33437), .B(n33436), .Z(n33490) );
  XOR U34299 ( .A(a[810]), .B(n42197), .Z(n33479) );
  NANDN U34300 ( .A(n33479), .B(n42173), .Z(n33440) );
  NANDN U34301 ( .A(n33438), .B(n42172), .Z(n33439) );
  NAND U34302 ( .A(n33440), .B(n33439), .Z(n33488) );
  NAND U34303 ( .A(b[7]), .B(a[806]), .Z(n33489) );
  XNOR U34304 ( .A(n33488), .B(n33489), .Z(n33491) );
  XOR U34305 ( .A(n33490), .B(n33491), .Z(n33497) );
  NANDN U34306 ( .A(n33441), .B(n42093), .Z(n33443) );
  XOR U34307 ( .A(n42134), .B(a[812]), .Z(n33482) );
  NANDN U34308 ( .A(n33482), .B(n42095), .Z(n33442) );
  NAND U34309 ( .A(n33443), .B(n33442), .Z(n33495) );
  NANDN U34310 ( .A(n33444), .B(n42231), .Z(n33446) );
  XOR U34311 ( .A(n229), .B(a[808]), .Z(n33485) );
  NANDN U34312 ( .A(n33485), .B(n42234), .Z(n33445) );
  AND U34313 ( .A(n33446), .B(n33445), .Z(n33494) );
  XNOR U34314 ( .A(n33495), .B(n33494), .Z(n33496) );
  XNOR U34315 ( .A(n33497), .B(n33496), .Z(n33501) );
  NANDN U34316 ( .A(n33448), .B(n33447), .Z(n33452) );
  NAND U34317 ( .A(n33450), .B(n33449), .Z(n33451) );
  AND U34318 ( .A(n33452), .B(n33451), .Z(n33500) );
  XOR U34319 ( .A(n33501), .B(n33500), .Z(n33502) );
  NANDN U34320 ( .A(n33454), .B(n33453), .Z(n33458) );
  NANDN U34321 ( .A(n33456), .B(n33455), .Z(n33457) );
  NAND U34322 ( .A(n33458), .B(n33457), .Z(n33503) );
  XOR U34323 ( .A(n33502), .B(n33503), .Z(n33470) );
  OR U34324 ( .A(n33460), .B(n33459), .Z(n33464) );
  NANDN U34325 ( .A(n33462), .B(n33461), .Z(n33463) );
  NAND U34326 ( .A(n33464), .B(n33463), .Z(n33471) );
  XNOR U34327 ( .A(n33470), .B(n33471), .Z(n33472) );
  XNOR U34328 ( .A(n33473), .B(n33472), .Z(n33506) );
  XNOR U34329 ( .A(n33506), .B(sreg[1830]), .Z(n33508) );
  NAND U34330 ( .A(n33465), .B(sreg[1829]), .Z(n33469) );
  OR U34331 ( .A(n33467), .B(n33466), .Z(n33468) );
  AND U34332 ( .A(n33469), .B(n33468), .Z(n33507) );
  XOR U34333 ( .A(n33508), .B(n33507), .Z(c[1830]) );
  NANDN U34334 ( .A(n33471), .B(n33470), .Z(n33475) );
  NAND U34335 ( .A(n33473), .B(n33472), .Z(n33474) );
  NAND U34336 ( .A(n33475), .B(n33474), .Z(n33514) );
  NAND U34337 ( .A(b[0]), .B(a[815]), .Z(n33476) );
  XNOR U34338 ( .A(b[1]), .B(n33476), .Z(n33478) );
  NAND U34339 ( .A(n131), .B(a[814]), .Z(n33477) );
  AND U34340 ( .A(n33478), .B(n33477), .Z(n33531) );
  XOR U34341 ( .A(a[811]), .B(n42197), .Z(n33520) );
  NANDN U34342 ( .A(n33520), .B(n42173), .Z(n33481) );
  NANDN U34343 ( .A(n33479), .B(n42172), .Z(n33480) );
  NAND U34344 ( .A(n33481), .B(n33480), .Z(n33529) );
  NAND U34345 ( .A(b[7]), .B(a[807]), .Z(n33530) );
  XNOR U34346 ( .A(n33529), .B(n33530), .Z(n33532) );
  XOR U34347 ( .A(n33531), .B(n33532), .Z(n33538) );
  NANDN U34348 ( .A(n33482), .B(n42093), .Z(n33484) );
  XOR U34349 ( .A(n42134), .B(a[813]), .Z(n33523) );
  NANDN U34350 ( .A(n33523), .B(n42095), .Z(n33483) );
  NAND U34351 ( .A(n33484), .B(n33483), .Z(n33536) );
  NANDN U34352 ( .A(n33485), .B(n42231), .Z(n33487) );
  XOR U34353 ( .A(n229), .B(a[809]), .Z(n33526) );
  NANDN U34354 ( .A(n33526), .B(n42234), .Z(n33486) );
  AND U34355 ( .A(n33487), .B(n33486), .Z(n33535) );
  XNOR U34356 ( .A(n33536), .B(n33535), .Z(n33537) );
  XNOR U34357 ( .A(n33538), .B(n33537), .Z(n33542) );
  NANDN U34358 ( .A(n33489), .B(n33488), .Z(n33493) );
  NAND U34359 ( .A(n33491), .B(n33490), .Z(n33492) );
  AND U34360 ( .A(n33493), .B(n33492), .Z(n33541) );
  XOR U34361 ( .A(n33542), .B(n33541), .Z(n33543) );
  NANDN U34362 ( .A(n33495), .B(n33494), .Z(n33499) );
  NANDN U34363 ( .A(n33497), .B(n33496), .Z(n33498) );
  NAND U34364 ( .A(n33499), .B(n33498), .Z(n33544) );
  XOR U34365 ( .A(n33543), .B(n33544), .Z(n33511) );
  OR U34366 ( .A(n33501), .B(n33500), .Z(n33505) );
  NANDN U34367 ( .A(n33503), .B(n33502), .Z(n33504) );
  NAND U34368 ( .A(n33505), .B(n33504), .Z(n33512) );
  XNOR U34369 ( .A(n33511), .B(n33512), .Z(n33513) );
  XNOR U34370 ( .A(n33514), .B(n33513), .Z(n33547) );
  XNOR U34371 ( .A(n33547), .B(sreg[1831]), .Z(n33549) );
  NAND U34372 ( .A(n33506), .B(sreg[1830]), .Z(n33510) );
  OR U34373 ( .A(n33508), .B(n33507), .Z(n33509) );
  AND U34374 ( .A(n33510), .B(n33509), .Z(n33548) );
  XOR U34375 ( .A(n33549), .B(n33548), .Z(c[1831]) );
  NANDN U34376 ( .A(n33512), .B(n33511), .Z(n33516) );
  NAND U34377 ( .A(n33514), .B(n33513), .Z(n33515) );
  NAND U34378 ( .A(n33516), .B(n33515), .Z(n33555) );
  NAND U34379 ( .A(b[0]), .B(a[816]), .Z(n33517) );
  XNOR U34380 ( .A(b[1]), .B(n33517), .Z(n33519) );
  NAND U34381 ( .A(n131), .B(a[815]), .Z(n33518) );
  AND U34382 ( .A(n33519), .B(n33518), .Z(n33572) );
  XOR U34383 ( .A(a[812]), .B(n42197), .Z(n33561) );
  NANDN U34384 ( .A(n33561), .B(n42173), .Z(n33522) );
  NANDN U34385 ( .A(n33520), .B(n42172), .Z(n33521) );
  NAND U34386 ( .A(n33522), .B(n33521), .Z(n33570) );
  NAND U34387 ( .A(b[7]), .B(a[808]), .Z(n33571) );
  XNOR U34388 ( .A(n33570), .B(n33571), .Z(n33573) );
  XOR U34389 ( .A(n33572), .B(n33573), .Z(n33579) );
  NANDN U34390 ( .A(n33523), .B(n42093), .Z(n33525) );
  XOR U34391 ( .A(n42134), .B(a[814]), .Z(n33564) );
  NANDN U34392 ( .A(n33564), .B(n42095), .Z(n33524) );
  NAND U34393 ( .A(n33525), .B(n33524), .Z(n33577) );
  NANDN U34394 ( .A(n33526), .B(n42231), .Z(n33528) );
  XOR U34395 ( .A(n229), .B(a[810]), .Z(n33567) );
  NANDN U34396 ( .A(n33567), .B(n42234), .Z(n33527) );
  AND U34397 ( .A(n33528), .B(n33527), .Z(n33576) );
  XNOR U34398 ( .A(n33577), .B(n33576), .Z(n33578) );
  XNOR U34399 ( .A(n33579), .B(n33578), .Z(n33583) );
  NANDN U34400 ( .A(n33530), .B(n33529), .Z(n33534) );
  NAND U34401 ( .A(n33532), .B(n33531), .Z(n33533) );
  AND U34402 ( .A(n33534), .B(n33533), .Z(n33582) );
  XOR U34403 ( .A(n33583), .B(n33582), .Z(n33584) );
  NANDN U34404 ( .A(n33536), .B(n33535), .Z(n33540) );
  NANDN U34405 ( .A(n33538), .B(n33537), .Z(n33539) );
  NAND U34406 ( .A(n33540), .B(n33539), .Z(n33585) );
  XOR U34407 ( .A(n33584), .B(n33585), .Z(n33552) );
  OR U34408 ( .A(n33542), .B(n33541), .Z(n33546) );
  NANDN U34409 ( .A(n33544), .B(n33543), .Z(n33545) );
  NAND U34410 ( .A(n33546), .B(n33545), .Z(n33553) );
  XNOR U34411 ( .A(n33552), .B(n33553), .Z(n33554) );
  XNOR U34412 ( .A(n33555), .B(n33554), .Z(n33588) );
  XNOR U34413 ( .A(n33588), .B(sreg[1832]), .Z(n33590) );
  NAND U34414 ( .A(n33547), .B(sreg[1831]), .Z(n33551) );
  OR U34415 ( .A(n33549), .B(n33548), .Z(n33550) );
  AND U34416 ( .A(n33551), .B(n33550), .Z(n33589) );
  XOR U34417 ( .A(n33590), .B(n33589), .Z(c[1832]) );
  NANDN U34418 ( .A(n33553), .B(n33552), .Z(n33557) );
  NAND U34419 ( .A(n33555), .B(n33554), .Z(n33556) );
  NAND U34420 ( .A(n33557), .B(n33556), .Z(n33596) );
  NAND U34421 ( .A(b[0]), .B(a[817]), .Z(n33558) );
  XNOR U34422 ( .A(b[1]), .B(n33558), .Z(n33560) );
  NAND U34423 ( .A(n131), .B(a[816]), .Z(n33559) );
  AND U34424 ( .A(n33560), .B(n33559), .Z(n33613) );
  XOR U34425 ( .A(a[813]), .B(n42197), .Z(n33602) );
  NANDN U34426 ( .A(n33602), .B(n42173), .Z(n33563) );
  NANDN U34427 ( .A(n33561), .B(n42172), .Z(n33562) );
  NAND U34428 ( .A(n33563), .B(n33562), .Z(n33611) );
  NAND U34429 ( .A(b[7]), .B(a[809]), .Z(n33612) );
  XNOR U34430 ( .A(n33611), .B(n33612), .Z(n33614) );
  XOR U34431 ( .A(n33613), .B(n33614), .Z(n33620) );
  NANDN U34432 ( .A(n33564), .B(n42093), .Z(n33566) );
  XOR U34433 ( .A(n42134), .B(a[815]), .Z(n33605) );
  NANDN U34434 ( .A(n33605), .B(n42095), .Z(n33565) );
  NAND U34435 ( .A(n33566), .B(n33565), .Z(n33618) );
  NANDN U34436 ( .A(n33567), .B(n42231), .Z(n33569) );
  XOR U34437 ( .A(n229), .B(a[811]), .Z(n33608) );
  NANDN U34438 ( .A(n33608), .B(n42234), .Z(n33568) );
  AND U34439 ( .A(n33569), .B(n33568), .Z(n33617) );
  XNOR U34440 ( .A(n33618), .B(n33617), .Z(n33619) );
  XNOR U34441 ( .A(n33620), .B(n33619), .Z(n33624) );
  NANDN U34442 ( .A(n33571), .B(n33570), .Z(n33575) );
  NAND U34443 ( .A(n33573), .B(n33572), .Z(n33574) );
  AND U34444 ( .A(n33575), .B(n33574), .Z(n33623) );
  XOR U34445 ( .A(n33624), .B(n33623), .Z(n33625) );
  NANDN U34446 ( .A(n33577), .B(n33576), .Z(n33581) );
  NANDN U34447 ( .A(n33579), .B(n33578), .Z(n33580) );
  NAND U34448 ( .A(n33581), .B(n33580), .Z(n33626) );
  XOR U34449 ( .A(n33625), .B(n33626), .Z(n33593) );
  OR U34450 ( .A(n33583), .B(n33582), .Z(n33587) );
  NANDN U34451 ( .A(n33585), .B(n33584), .Z(n33586) );
  NAND U34452 ( .A(n33587), .B(n33586), .Z(n33594) );
  XNOR U34453 ( .A(n33593), .B(n33594), .Z(n33595) );
  XNOR U34454 ( .A(n33596), .B(n33595), .Z(n33629) );
  XNOR U34455 ( .A(n33629), .B(sreg[1833]), .Z(n33631) );
  NAND U34456 ( .A(n33588), .B(sreg[1832]), .Z(n33592) );
  OR U34457 ( .A(n33590), .B(n33589), .Z(n33591) );
  AND U34458 ( .A(n33592), .B(n33591), .Z(n33630) );
  XOR U34459 ( .A(n33631), .B(n33630), .Z(c[1833]) );
  NANDN U34460 ( .A(n33594), .B(n33593), .Z(n33598) );
  NAND U34461 ( .A(n33596), .B(n33595), .Z(n33597) );
  NAND U34462 ( .A(n33598), .B(n33597), .Z(n33637) );
  NAND U34463 ( .A(b[0]), .B(a[818]), .Z(n33599) );
  XNOR U34464 ( .A(b[1]), .B(n33599), .Z(n33601) );
  NAND U34465 ( .A(n131), .B(a[817]), .Z(n33600) );
  AND U34466 ( .A(n33601), .B(n33600), .Z(n33654) );
  XOR U34467 ( .A(a[814]), .B(n42197), .Z(n33643) );
  NANDN U34468 ( .A(n33643), .B(n42173), .Z(n33604) );
  NANDN U34469 ( .A(n33602), .B(n42172), .Z(n33603) );
  NAND U34470 ( .A(n33604), .B(n33603), .Z(n33652) );
  NAND U34471 ( .A(b[7]), .B(a[810]), .Z(n33653) );
  XNOR U34472 ( .A(n33652), .B(n33653), .Z(n33655) );
  XOR U34473 ( .A(n33654), .B(n33655), .Z(n33661) );
  NANDN U34474 ( .A(n33605), .B(n42093), .Z(n33607) );
  XOR U34475 ( .A(n42134), .B(a[816]), .Z(n33646) );
  NANDN U34476 ( .A(n33646), .B(n42095), .Z(n33606) );
  NAND U34477 ( .A(n33607), .B(n33606), .Z(n33659) );
  NANDN U34478 ( .A(n33608), .B(n42231), .Z(n33610) );
  XOR U34479 ( .A(n229), .B(a[812]), .Z(n33649) );
  NANDN U34480 ( .A(n33649), .B(n42234), .Z(n33609) );
  AND U34481 ( .A(n33610), .B(n33609), .Z(n33658) );
  XNOR U34482 ( .A(n33659), .B(n33658), .Z(n33660) );
  XNOR U34483 ( .A(n33661), .B(n33660), .Z(n33665) );
  NANDN U34484 ( .A(n33612), .B(n33611), .Z(n33616) );
  NAND U34485 ( .A(n33614), .B(n33613), .Z(n33615) );
  AND U34486 ( .A(n33616), .B(n33615), .Z(n33664) );
  XOR U34487 ( .A(n33665), .B(n33664), .Z(n33666) );
  NANDN U34488 ( .A(n33618), .B(n33617), .Z(n33622) );
  NANDN U34489 ( .A(n33620), .B(n33619), .Z(n33621) );
  NAND U34490 ( .A(n33622), .B(n33621), .Z(n33667) );
  XOR U34491 ( .A(n33666), .B(n33667), .Z(n33634) );
  OR U34492 ( .A(n33624), .B(n33623), .Z(n33628) );
  NANDN U34493 ( .A(n33626), .B(n33625), .Z(n33627) );
  NAND U34494 ( .A(n33628), .B(n33627), .Z(n33635) );
  XNOR U34495 ( .A(n33634), .B(n33635), .Z(n33636) );
  XNOR U34496 ( .A(n33637), .B(n33636), .Z(n33670) );
  XNOR U34497 ( .A(n33670), .B(sreg[1834]), .Z(n33672) );
  NAND U34498 ( .A(n33629), .B(sreg[1833]), .Z(n33633) );
  OR U34499 ( .A(n33631), .B(n33630), .Z(n33632) );
  AND U34500 ( .A(n33633), .B(n33632), .Z(n33671) );
  XOR U34501 ( .A(n33672), .B(n33671), .Z(c[1834]) );
  NANDN U34502 ( .A(n33635), .B(n33634), .Z(n33639) );
  NAND U34503 ( .A(n33637), .B(n33636), .Z(n33638) );
  NAND U34504 ( .A(n33639), .B(n33638), .Z(n33678) );
  NAND U34505 ( .A(b[0]), .B(a[819]), .Z(n33640) );
  XNOR U34506 ( .A(b[1]), .B(n33640), .Z(n33642) );
  NAND U34507 ( .A(n132), .B(a[818]), .Z(n33641) );
  AND U34508 ( .A(n33642), .B(n33641), .Z(n33695) );
  XOR U34509 ( .A(a[815]), .B(n42197), .Z(n33684) );
  NANDN U34510 ( .A(n33684), .B(n42173), .Z(n33645) );
  NANDN U34511 ( .A(n33643), .B(n42172), .Z(n33644) );
  NAND U34512 ( .A(n33645), .B(n33644), .Z(n33693) );
  NAND U34513 ( .A(b[7]), .B(a[811]), .Z(n33694) );
  XNOR U34514 ( .A(n33693), .B(n33694), .Z(n33696) );
  XOR U34515 ( .A(n33695), .B(n33696), .Z(n33702) );
  NANDN U34516 ( .A(n33646), .B(n42093), .Z(n33648) );
  XOR U34517 ( .A(n42134), .B(a[817]), .Z(n33687) );
  NANDN U34518 ( .A(n33687), .B(n42095), .Z(n33647) );
  NAND U34519 ( .A(n33648), .B(n33647), .Z(n33700) );
  NANDN U34520 ( .A(n33649), .B(n42231), .Z(n33651) );
  XOR U34521 ( .A(n229), .B(a[813]), .Z(n33690) );
  NANDN U34522 ( .A(n33690), .B(n42234), .Z(n33650) );
  AND U34523 ( .A(n33651), .B(n33650), .Z(n33699) );
  XNOR U34524 ( .A(n33700), .B(n33699), .Z(n33701) );
  XNOR U34525 ( .A(n33702), .B(n33701), .Z(n33706) );
  NANDN U34526 ( .A(n33653), .B(n33652), .Z(n33657) );
  NAND U34527 ( .A(n33655), .B(n33654), .Z(n33656) );
  AND U34528 ( .A(n33657), .B(n33656), .Z(n33705) );
  XOR U34529 ( .A(n33706), .B(n33705), .Z(n33707) );
  NANDN U34530 ( .A(n33659), .B(n33658), .Z(n33663) );
  NANDN U34531 ( .A(n33661), .B(n33660), .Z(n33662) );
  NAND U34532 ( .A(n33663), .B(n33662), .Z(n33708) );
  XOR U34533 ( .A(n33707), .B(n33708), .Z(n33675) );
  OR U34534 ( .A(n33665), .B(n33664), .Z(n33669) );
  NANDN U34535 ( .A(n33667), .B(n33666), .Z(n33668) );
  NAND U34536 ( .A(n33669), .B(n33668), .Z(n33676) );
  XNOR U34537 ( .A(n33675), .B(n33676), .Z(n33677) );
  XNOR U34538 ( .A(n33678), .B(n33677), .Z(n33711) );
  XNOR U34539 ( .A(n33711), .B(sreg[1835]), .Z(n33713) );
  NAND U34540 ( .A(n33670), .B(sreg[1834]), .Z(n33674) );
  OR U34541 ( .A(n33672), .B(n33671), .Z(n33673) );
  AND U34542 ( .A(n33674), .B(n33673), .Z(n33712) );
  XOR U34543 ( .A(n33713), .B(n33712), .Z(c[1835]) );
  NANDN U34544 ( .A(n33676), .B(n33675), .Z(n33680) );
  NAND U34545 ( .A(n33678), .B(n33677), .Z(n33679) );
  NAND U34546 ( .A(n33680), .B(n33679), .Z(n33719) );
  NAND U34547 ( .A(b[0]), .B(a[820]), .Z(n33681) );
  XNOR U34548 ( .A(b[1]), .B(n33681), .Z(n33683) );
  NAND U34549 ( .A(n132), .B(a[819]), .Z(n33682) );
  AND U34550 ( .A(n33683), .B(n33682), .Z(n33736) );
  XOR U34551 ( .A(a[816]), .B(n42197), .Z(n33725) );
  NANDN U34552 ( .A(n33725), .B(n42173), .Z(n33686) );
  NANDN U34553 ( .A(n33684), .B(n42172), .Z(n33685) );
  NAND U34554 ( .A(n33686), .B(n33685), .Z(n33734) );
  NAND U34555 ( .A(b[7]), .B(a[812]), .Z(n33735) );
  XNOR U34556 ( .A(n33734), .B(n33735), .Z(n33737) );
  XOR U34557 ( .A(n33736), .B(n33737), .Z(n33743) );
  NANDN U34558 ( .A(n33687), .B(n42093), .Z(n33689) );
  XOR U34559 ( .A(n42134), .B(a[818]), .Z(n33728) );
  NANDN U34560 ( .A(n33728), .B(n42095), .Z(n33688) );
  NAND U34561 ( .A(n33689), .B(n33688), .Z(n33741) );
  NANDN U34562 ( .A(n33690), .B(n42231), .Z(n33692) );
  XOR U34563 ( .A(n229), .B(a[814]), .Z(n33731) );
  NANDN U34564 ( .A(n33731), .B(n42234), .Z(n33691) );
  AND U34565 ( .A(n33692), .B(n33691), .Z(n33740) );
  XNOR U34566 ( .A(n33741), .B(n33740), .Z(n33742) );
  XNOR U34567 ( .A(n33743), .B(n33742), .Z(n33747) );
  NANDN U34568 ( .A(n33694), .B(n33693), .Z(n33698) );
  NAND U34569 ( .A(n33696), .B(n33695), .Z(n33697) );
  AND U34570 ( .A(n33698), .B(n33697), .Z(n33746) );
  XOR U34571 ( .A(n33747), .B(n33746), .Z(n33748) );
  NANDN U34572 ( .A(n33700), .B(n33699), .Z(n33704) );
  NANDN U34573 ( .A(n33702), .B(n33701), .Z(n33703) );
  NAND U34574 ( .A(n33704), .B(n33703), .Z(n33749) );
  XOR U34575 ( .A(n33748), .B(n33749), .Z(n33716) );
  OR U34576 ( .A(n33706), .B(n33705), .Z(n33710) );
  NANDN U34577 ( .A(n33708), .B(n33707), .Z(n33709) );
  NAND U34578 ( .A(n33710), .B(n33709), .Z(n33717) );
  XNOR U34579 ( .A(n33716), .B(n33717), .Z(n33718) );
  XNOR U34580 ( .A(n33719), .B(n33718), .Z(n33752) );
  XNOR U34581 ( .A(n33752), .B(sreg[1836]), .Z(n33754) );
  NAND U34582 ( .A(n33711), .B(sreg[1835]), .Z(n33715) );
  OR U34583 ( .A(n33713), .B(n33712), .Z(n33714) );
  AND U34584 ( .A(n33715), .B(n33714), .Z(n33753) );
  XOR U34585 ( .A(n33754), .B(n33753), .Z(c[1836]) );
  NANDN U34586 ( .A(n33717), .B(n33716), .Z(n33721) );
  NAND U34587 ( .A(n33719), .B(n33718), .Z(n33720) );
  NAND U34588 ( .A(n33721), .B(n33720), .Z(n33760) );
  NAND U34589 ( .A(b[0]), .B(a[821]), .Z(n33722) );
  XNOR U34590 ( .A(b[1]), .B(n33722), .Z(n33724) );
  NAND U34591 ( .A(n132), .B(a[820]), .Z(n33723) );
  AND U34592 ( .A(n33724), .B(n33723), .Z(n33777) );
  XOR U34593 ( .A(a[817]), .B(n42197), .Z(n33766) );
  NANDN U34594 ( .A(n33766), .B(n42173), .Z(n33727) );
  NANDN U34595 ( .A(n33725), .B(n42172), .Z(n33726) );
  NAND U34596 ( .A(n33727), .B(n33726), .Z(n33775) );
  NAND U34597 ( .A(b[7]), .B(a[813]), .Z(n33776) );
  XNOR U34598 ( .A(n33775), .B(n33776), .Z(n33778) );
  XOR U34599 ( .A(n33777), .B(n33778), .Z(n33784) );
  NANDN U34600 ( .A(n33728), .B(n42093), .Z(n33730) );
  XOR U34601 ( .A(n42134), .B(a[819]), .Z(n33769) );
  NANDN U34602 ( .A(n33769), .B(n42095), .Z(n33729) );
  NAND U34603 ( .A(n33730), .B(n33729), .Z(n33782) );
  NANDN U34604 ( .A(n33731), .B(n42231), .Z(n33733) );
  XOR U34605 ( .A(n230), .B(a[815]), .Z(n33772) );
  NANDN U34606 ( .A(n33772), .B(n42234), .Z(n33732) );
  AND U34607 ( .A(n33733), .B(n33732), .Z(n33781) );
  XNOR U34608 ( .A(n33782), .B(n33781), .Z(n33783) );
  XNOR U34609 ( .A(n33784), .B(n33783), .Z(n33788) );
  NANDN U34610 ( .A(n33735), .B(n33734), .Z(n33739) );
  NAND U34611 ( .A(n33737), .B(n33736), .Z(n33738) );
  AND U34612 ( .A(n33739), .B(n33738), .Z(n33787) );
  XOR U34613 ( .A(n33788), .B(n33787), .Z(n33789) );
  NANDN U34614 ( .A(n33741), .B(n33740), .Z(n33745) );
  NANDN U34615 ( .A(n33743), .B(n33742), .Z(n33744) );
  NAND U34616 ( .A(n33745), .B(n33744), .Z(n33790) );
  XOR U34617 ( .A(n33789), .B(n33790), .Z(n33757) );
  OR U34618 ( .A(n33747), .B(n33746), .Z(n33751) );
  NANDN U34619 ( .A(n33749), .B(n33748), .Z(n33750) );
  NAND U34620 ( .A(n33751), .B(n33750), .Z(n33758) );
  XNOR U34621 ( .A(n33757), .B(n33758), .Z(n33759) );
  XNOR U34622 ( .A(n33760), .B(n33759), .Z(n33793) );
  XNOR U34623 ( .A(n33793), .B(sreg[1837]), .Z(n33795) );
  NAND U34624 ( .A(n33752), .B(sreg[1836]), .Z(n33756) );
  OR U34625 ( .A(n33754), .B(n33753), .Z(n33755) );
  AND U34626 ( .A(n33756), .B(n33755), .Z(n33794) );
  XOR U34627 ( .A(n33795), .B(n33794), .Z(c[1837]) );
  NANDN U34628 ( .A(n33758), .B(n33757), .Z(n33762) );
  NAND U34629 ( .A(n33760), .B(n33759), .Z(n33761) );
  NAND U34630 ( .A(n33762), .B(n33761), .Z(n33801) );
  NAND U34631 ( .A(b[0]), .B(a[822]), .Z(n33763) );
  XNOR U34632 ( .A(b[1]), .B(n33763), .Z(n33765) );
  NAND U34633 ( .A(n132), .B(a[821]), .Z(n33764) );
  AND U34634 ( .A(n33765), .B(n33764), .Z(n33818) );
  XOR U34635 ( .A(a[818]), .B(n42197), .Z(n33807) );
  NANDN U34636 ( .A(n33807), .B(n42173), .Z(n33768) );
  NANDN U34637 ( .A(n33766), .B(n42172), .Z(n33767) );
  NAND U34638 ( .A(n33768), .B(n33767), .Z(n33816) );
  NAND U34639 ( .A(b[7]), .B(a[814]), .Z(n33817) );
  XNOR U34640 ( .A(n33816), .B(n33817), .Z(n33819) );
  XOR U34641 ( .A(n33818), .B(n33819), .Z(n33825) );
  NANDN U34642 ( .A(n33769), .B(n42093), .Z(n33771) );
  XOR U34643 ( .A(n42134), .B(a[820]), .Z(n33810) );
  NANDN U34644 ( .A(n33810), .B(n42095), .Z(n33770) );
  NAND U34645 ( .A(n33771), .B(n33770), .Z(n33823) );
  NANDN U34646 ( .A(n33772), .B(n42231), .Z(n33774) );
  XOR U34647 ( .A(n230), .B(a[816]), .Z(n33813) );
  NANDN U34648 ( .A(n33813), .B(n42234), .Z(n33773) );
  AND U34649 ( .A(n33774), .B(n33773), .Z(n33822) );
  XNOR U34650 ( .A(n33823), .B(n33822), .Z(n33824) );
  XNOR U34651 ( .A(n33825), .B(n33824), .Z(n33829) );
  NANDN U34652 ( .A(n33776), .B(n33775), .Z(n33780) );
  NAND U34653 ( .A(n33778), .B(n33777), .Z(n33779) );
  AND U34654 ( .A(n33780), .B(n33779), .Z(n33828) );
  XOR U34655 ( .A(n33829), .B(n33828), .Z(n33830) );
  NANDN U34656 ( .A(n33782), .B(n33781), .Z(n33786) );
  NANDN U34657 ( .A(n33784), .B(n33783), .Z(n33785) );
  NAND U34658 ( .A(n33786), .B(n33785), .Z(n33831) );
  XOR U34659 ( .A(n33830), .B(n33831), .Z(n33798) );
  OR U34660 ( .A(n33788), .B(n33787), .Z(n33792) );
  NANDN U34661 ( .A(n33790), .B(n33789), .Z(n33791) );
  NAND U34662 ( .A(n33792), .B(n33791), .Z(n33799) );
  XNOR U34663 ( .A(n33798), .B(n33799), .Z(n33800) );
  XNOR U34664 ( .A(n33801), .B(n33800), .Z(n33834) );
  XNOR U34665 ( .A(n33834), .B(sreg[1838]), .Z(n33836) );
  NAND U34666 ( .A(n33793), .B(sreg[1837]), .Z(n33797) );
  OR U34667 ( .A(n33795), .B(n33794), .Z(n33796) );
  AND U34668 ( .A(n33797), .B(n33796), .Z(n33835) );
  XOR U34669 ( .A(n33836), .B(n33835), .Z(c[1838]) );
  NANDN U34670 ( .A(n33799), .B(n33798), .Z(n33803) );
  NAND U34671 ( .A(n33801), .B(n33800), .Z(n33802) );
  NAND U34672 ( .A(n33803), .B(n33802), .Z(n33842) );
  NAND U34673 ( .A(b[0]), .B(a[823]), .Z(n33804) );
  XNOR U34674 ( .A(b[1]), .B(n33804), .Z(n33806) );
  NAND U34675 ( .A(n132), .B(a[822]), .Z(n33805) );
  AND U34676 ( .A(n33806), .B(n33805), .Z(n33859) );
  XOR U34677 ( .A(a[819]), .B(n42197), .Z(n33848) );
  NANDN U34678 ( .A(n33848), .B(n42173), .Z(n33809) );
  NANDN U34679 ( .A(n33807), .B(n42172), .Z(n33808) );
  NAND U34680 ( .A(n33809), .B(n33808), .Z(n33857) );
  NAND U34681 ( .A(b[7]), .B(a[815]), .Z(n33858) );
  XNOR U34682 ( .A(n33857), .B(n33858), .Z(n33860) );
  XOR U34683 ( .A(n33859), .B(n33860), .Z(n33866) );
  NANDN U34684 ( .A(n33810), .B(n42093), .Z(n33812) );
  XOR U34685 ( .A(n42134), .B(a[821]), .Z(n33851) );
  NANDN U34686 ( .A(n33851), .B(n42095), .Z(n33811) );
  NAND U34687 ( .A(n33812), .B(n33811), .Z(n33864) );
  NANDN U34688 ( .A(n33813), .B(n42231), .Z(n33815) );
  XOR U34689 ( .A(n230), .B(a[817]), .Z(n33854) );
  NANDN U34690 ( .A(n33854), .B(n42234), .Z(n33814) );
  AND U34691 ( .A(n33815), .B(n33814), .Z(n33863) );
  XNOR U34692 ( .A(n33864), .B(n33863), .Z(n33865) );
  XNOR U34693 ( .A(n33866), .B(n33865), .Z(n33870) );
  NANDN U34694 ( .A(n33817), .B(n33816), .Z(n33821) );
  NAND U34695 ( .A(n33819), .B(n33818), .Z(n33820) );
  AND U34696 ( .A(n33821), .B(n33820), .Z(n33869) );
  XOR U34697 ( .A(n33870), .B(n33869), .Z(n33871) );
  NANDN U34698 ( .A(n33823), .B(n33822), .Z(n33827) );
  NANDN U34699 ( .A(n33825), .B(n33824), .Z(n33826) );
  NAND U34700 ( .A(n33827), .B(n33826), .Z(n33872) );
  XOR U34701 ( .A(n33871), .B(n33872), .Z(n33839) );
  OR U34702 ( .A(n33829), .B(n33828), .Z(n33833) );
  NANDN U34703 ( .A(n33831), .B(n33830), .Z(n33832) );
  NAND U34704 ( .A(n33833), .B(n33832), .Z(n33840) );
  XNOR U34705 ( .A(n33839), .B(n33840), .Z(n33841) );
  XNOR U34706 ( .A(n33842), .B(n33841), .Z(n33875) );
  XNOR U34707 ( .A(n33875), .B(sreg[1839]), .Z(n33877) );
  NAND U34708 ( .A(n33834), .B(sreg[1838]), .Z(n33838) );
  OR U34709 ( .A(n33836), .B(n33835), .Z(n33837) );
  AND U34710 ( .A(n33838), .B(n33837), .Z(n33876) );
  XOR U34711 ( .A(n33877), .B(n33876), .Z(c[1839]) );
  NANDN U34712 ( .A(n33840), .B(n33839), .Z(n33844) );
  NAND U34713 ( .A(n33842), .B(n33841), .Z(n33843) );
  NAND U34714 ( .A(n33844), .B(n33843), .Z(n33883) );
  NAND U34715 ( .A(b[0]), .B(a[824]), .Z(n33845) );
  XNOR U34716 ( .A(b[1]), .B(n33845), .Z(n33847) );
  NAND U34717 ( .A(n132), .B(a[823]), .Z(n33846) );
  AND U34718 ( .A(n33847), .B(n33846), .Z(n33900) );
  XOR U34719 ( .A(a[820]), .B(n42197), .Z(n33889) );
  NANDN U34720 ( .A(n33889), .B(n42173), .Z(n33850) );
  NANDN U34721 ( .A(n33848), .B(n42172), .Z(n33849) );
  NAND U34722 ( .A(n33850), .B(n33849), .Z(n33898) );
  NAND U34723 ( .A(b[7]), .B(a[816]), .Z(n33899) );
  XNOR U34724 ( .A(n33898), .B(n33899), .Z(n33901) );
  XOR U34725 ( .A(n33900), .B(n33901), .Z(n33907) );
  NANDN U34726 ( .A(n33851), .B(n42093), .Z(n33853) );
  XOR U34727 ( .A(n42134), .B(a[822]), .Z(n33892) );
  NANDN U34728 ( .A(n33892), .B(n42095), .Z(n33852) );
  NAND U34729 ( .A(n33853), .B(n33852), .Z(n33905) );
  NANDN U34730 ( .A(n33854), .B(n42231), .Z(n33856) );
  XOR U34731 ( .A(n230), .B(a[818]), .Z(n33895) );
  NANDN U34732 ( .A(n33895), .B(n42234), .Z(n33855) );
  AND U34733 ( .A(n33856), .B(n33855), .Z(n33904) );
  XNOR U34734 ( .A(n33905), .B(n33904), .Z(n33906) );
  XNOR U34735 ( .A(n33907), .B(n33906), .Z(n33911) );
  NANDN U34736 ( .A(n33858), .B(n33857), .Z(n33862) );
  NAND U34737 ( .A(n33860), .B(n33859), .Z(n33861) );
  AND U34738 ( .A(n33862), .B(n33861), .Z(n33910) );
  XOR U34739 ( .A(n33911), .B(n33910), .Z(n33912) );
  NANDN U34740 ( .A(n33864), .B(n33863), .Z(n33868) );
  NANDN U34741 ( .A(n33866), .B(n33865), .Z(n33867) );
  NAND U34742 ( .A(n33868), .B(n33867), .Z(n33913) );
  XOR U34743 ( .A(n33912), .B(n33913), .Z(n33880) );
  OR U34744 ( .A(n33870), .B(n33869), .Z(n33874) );
  NANDN U34745 ( .A(n33872), .B(n33871), .Z(n33873) );
  NAND U34746 ( .A(n33874), .B(n33873), .Z(n33881) );
  XNOR U34747 ( .A(n33880), .B(n33881), .Z(n33882) );
  XNOR U34748 ( .A(n33883), .B(n33882), .Z(n33916) );
  XNOR U34749 ( .A(n33916), .B(sreg[1840]), .Z(n33918) );
  NAND U34750 ( .A(n33875), .B(sreg[1839]), .Z(n33879) );
  OR U34751 ( .A(n33877), .B(n33876), .Z(n33878) );
  AND U34752 ( .A(n33879), .B(n33878), .Z(n33917) );
  XOR U34753 ( .A(n33918), .B(n33917), .Z(c[1840]) );
  NANDN U34754 ( .A(n33881), .B(n33880), .Z(n33885) );
  NAND U34755 ( .A(n33883), .B(n33882), .Z(n33884) );
  NAND U34756 ( .A(n33885), .B(n33884), .Z(n33924) );
  NAND U34757 ( .A(b[0]), .B(a[825]), .Z(n33886) );
  XNOR U34758 ( .A(b[1]), .B(n33886), .Z(n33888) );
  NAND U34759 ( .A(n132), .B(a[824]), .Z(n33887) );
  AND U34760 ( .A(n33888), .B(n33887), .Z(n33941) );
  XOR U34761 ( .A(a[821]), .B(n42197), .Z(n33930) );
  NANDN U34762 ( .A(n33930), .B(n42173), .Z(n33891) );
  NANDN U34763 ( .A(n33889), .B(n42172), .Z(n33890) );
  NAND U34764 ( .A(n33891), .B(n33890), .Z(n33939) );
  NAND U34765 ( .A(b[7]), .B(a[817]), .Z(n33940) );
  XNOR U34766 ( .A(n33939), .B(n33940), .Z(n33942) );
  XOR U34767 ( .A(n33941), .B(n33942), .Z(n33948) );
  NANDN U34768 ( .A(n33892), .B(n42093), .Z(n33894) );
  XOR U34769 ( .A(n42134), .B(a[823]), .Z(n33933) );
  NANDN U34770 ( .A(n33933), .B(n42095), .Z(n33893) );
  NAND U34771 ( .A(n33894), .B(n33893), .Z(n33946) );
  NANDN U34772 ( .A(n33895), .B(n42231), .Z(n33897) );
  XOR U34773 ( .A(n230), .B(a[819]), .Z(n33936) );
  NANDN U34774 ( .A(n33936), .B(n42234), .Z(n33896) );
  AND U34775 ( .A(n33897), .B(n33896), .Z(n33945) );
  XNOR U34776 ( .A(n33946), .B(n33945), .Z(n33947) );
  XNOR U34777 ( .A(n33948), .B(n33947), .Z(n33952) );
  NANDN U34778 ( .A(n33899), .B(n33898), .Z(n33903) );
  NAND U34779 ( .A(n33901), .B(n33900), .Z(n33902) );
  AND U34780 ( .A(n33903), .B(n33902), .Z(n33951) );
  XOR U34781 ( .A(n33952), .B(n33951), .Z(n33953) );
  NANDN U34782 ( .A(n33905), .B(n33904), .Z(n33909) );
  NANDN U34783 ( .A(n33907), .B(n33906), .Z(n33908) );
  NAND U34784 ( .A(n33909), .B(n33908), .Z(n33954) );
  XOR U34785 ( .A(n33953), .B(n33954), .Z(n33921) );
  OR U34786 ( .A(n33911), .B(n33910), .Z(n33915) );
  NANDN U34787 ( .A(n33913), .B(n33912), .Z(n33914) );
  NAND U34788 ( .A(n33915), .B(n33914), .Z(n33922) );
  XNOR U34789 ( .A(n33921), .B(n33922), .Z(n33923) );
  XNOR U34790 ( .A(n33924), .B(n33923), .Z(n33957) );
  XNOR U34791 ( .A(n33957), .B(sreg[1841]), .Z(n33959) );
  NAND U34792 ( .A(n33916), .B(sreg[1840]), .Z(n33920) );
  OR U34793 ( .A(n33918), .B(n33917), .Z(n33919) );
  AND U34794 ( .A(n33920), .B(n33919), .Z(n33958) );
  XOR U34795 ( .A(n33959), .B(n33958), .Z(c[1841]) );
  NANDN U34796 ( .A(n33922), .B(n33921), .Z(n33926) );
  NAND U34797 ( .A(n33924), .B(n33923), .Z(n33925) );
  NAND U34798 ( .A(n33926), .B(n33925), .Z(n33965) );
  NAND U34799 ( .A(b[0]), .B(a[826]), .Z(n33927) );
  XNOR U34800 ( .A(b[1]), .B(n33927), .Z(n33929) );
  NAND U34801 ( .A(n133), .B(a[825]), .Z(n33928) );
  AND U34802 ( .A(n33929), .B(n33928), .Z(n33982) );
  XOR U34803 ( .A(a[822]), .B(n42197), .Z(n33971) );
  NANDN U34804 ( .A(n33971), .B(n42173), .Z(n33932) );
  NANDN U34805 ( .A(n33930), .B(n42172), .Z(n33931) );
  NAND U34806 ( .A(n33932), .B(n33931), .Z(n33980) );
  NAND U34807 ( .A(b[7]), .B(a[818]), .Z(n33981) );
  XNOR U34808 ( .A(n33980), .B(n33981), .Z(n33983) );
  XOR U34809 ( .A(n33982), .B(n33983), .Z(n33989) );
  NANDN U34810 ( .A(n33933), .B(n42093), .Z(n33935) );
  XOR U34811 ( .A(n42134), .B(a[824]), .Z(n33974) );
  NANDN U34812 ( .A(n33974), .B(n42095), .Z(n33934) );
  NAND U34813 ( .A(n33935), .B(n33934), .Z(n33987) );
  NANDN U34814 ( .A(n33936), .B(n42231), .Z(n33938) );
  XOR U34815 ( .A(n230), .B(a[820]), .Z(n33977) );
  NANDN U34816 ( .A(n33977), .B(n42234), .Z(n33937) );
  AND U34817 ( .A(n33938), .B(n33937), .Z(n33986) );
  XNOR U34818 ( .A(n33987), .B(n33986), .Z(n33988) );
  XNOR U34819 ( .A(n33989), .B(n33988), .Z(n33993) );
  NANDN U34820 ( .A(n33940), .B(n33939), .Z(n33944) );
  NAND U34821 ( .A(n33942), .B(n33941), .Z(n33943) );
  AND U34822 ( .A(n33944), .B(n33943), .Z(n33992) );
  XOR U34823 ( .A(n33993), .B(n33992), .Z(n33994) );
  NANDN U34824 ( .A(n33946), .B(n33945), .Z(n33950) );
  NANDN U34825 ( .A(n33948), .B(n33947), .Z(n33949) );
  NAND U34826 ( .A(n33950), .B(n33949), .Z(n33995) );
  XOR U34827 ( .A(n33994), .B(n33995), .Z(n33962) );
  OR U34828 ( .A(n33952), .B(n33951), .Z(n33956) );
  NANDN U34829 ( .A(n33954), .B(n33953), .Z(n33955) );
  NAND U34830 ( .A(n33956), .B(n33955), .Z(n33963) );
  XNOR U34831 ( .A(n33962), .B(n33963), .Z(n33964) );
  XNOR U34832 ( .A(n33965), .B(n33964), .Z(n33998) );
  XNOR U34833 ( .A(n33998), .B(sreg[1842]), .Z(n34000) );
  NAND U34834 ( .A(n33957), .B(sreg[1841]), .Z(n33961) );
  OR U34835 ( .A(n33959), .B(n33958), .Z(n33960) );
  AND U34836 ( .A(n33961), .B(n33960), .Z(n33999) );
  XOR U34837 ( .A(n34000), .B(n33999), .Z(c[1842]) );
  NANDN U34838 ( .A(n33963), .B(n33962), .Z(n33967) );
  NAND U34839 ( .A(n33965), .B(n33964), .Z(n33966) );
  NAND U34840 ( .A(n33967), .B(n33966), .Z(n34006) );
  NAND U34841 ( .A(b[0]), .B(a[827]), .Z(n33968) );
  XNOR U34842 ( .A(b[1]), .B(n33968), .Z(n33970) );
  NAND U34843 ( .A(n133), .B(a[826]), .Z(n33969) );
  AND U34844 ( .A(n33970), .B(n33969), .Z(n34023) );
  XOR U34845 ( .A(a[823]), .B(n42197), .Z(n34012) );
  NANDN U34846 ( .A(n34012), .B(n42173), .Z(n33973) );
  NANDN U34847 ( .A(n33971), .B(n42172), .Z(n33972) );
  NAND U34848 ( .A(n33973), .B(n33972), .Z(n34021) );
  NAND U34849 ( .A(b[7]), .B(a[819]), .Z(n34022) );
  XNOR U34850 ( .A(n34021), .B(n34022), .Z(n34024) );
  XOR U34851 ( .A(n34023), .B(n34024), .Z(n34030) );
  NANDN U34852 ( .A(n33974), .B(n42093), .Z(n33976) );
  XOR U34853 ( .A(n42134), .B(a[825]), .Z(n34015) );
  NANDN U34854 ( .A(n34015), .B(n42095), .Z(n33975) );
  NAND U34855 ( .A(n33976), .B(n33975), .Z(n34028) );
  NANDN U34856 ( .A(n33977), .B(n42231), .Z(n33979) );
  XOR U34857 ( .A(n230), .B(a[821]), .Z(n34018) );
  NANDN U34858 ( .A(n34018), .B(n42234), .Z(n33978) );
  AND U34859 ( .A(n33979), .B(n33978), .Z(n34027) );
  XNOR U34860 ( .A(n34028), .B(n34027), .Z(n34029) );
  XNOR U34861 ( .A(n34030), .B(n34029), .Z(n34034) );
  NANDN U34862 ( .A(n33981), .B(n33980), .Z(n33985) );
  NAND U34863 ( .A(n33983), .B(n33982), .Z(n33984) );
  AND U34864 ( .A(n33985), .B(n33984), .Z(n34033) );
  XOR U34865 ( .A(n34034), .B(n34033), .Z(n34035) );
  NANDN U34866 ( .A(n33987), .B(n33986), .Z(n33991) );
  NANDN U34867 ( .A(n33989), .B(n33988), .Z(n33990) );
  NAND U34868 ( .A(n33991), .B(n33990), .Z(n34036) );
  XOR U34869 ( .A(n34035), .B(n34036), .Z(n34003) );
  OR U34870 ( .A(n33993), .B(n33992), .Z(n33997) );
  NANDN U34871 ( .A(n33995), .B(n33994), .Z(n33996) );
  NAND U34872 ( .A(n33997), .B(n33996), .Z(n34004) );
  XNOR U34873 ( .A(n34003), .B(n34004), .Z(n34005) );
  XNOR U34874 ( .A(n34006), .B(n34005), .Z(n34039) );
  XNOR U34875 ( .A(n34039), .B(sreg[1843]), .Z(n34041) );
  NAND U34876 ( .A(n33998), .B(sreg[1842]), .Z(n34002) );
  OR U34877 ( .A(n34000), .B(n33999), .Z(n34001) );
  AND U34878 ( .A(n34002), .B(n34001), .Z(n34040) );
  XOR U34879 ( .A(n34041), .B(n34040), .Z(c[1843]) );
  NANDN U34880 ( .A(n34004), .B(n34003), .Z(n34008) );
  NAND U34881 ( .A(n34006), .B(n34005), .Z(n34007) );
  NAND U34882 ( .A(n34008), .B(n34007), .Z(n34047) );
  NAND U34883 ( .A(b[0]), .B(a[828]), .Z(n34009) );
  XNOR U34884 ( .A(b[1]), .B(n34009), .Z(n34011) );
  NAND U34885 ( .A(n133), .B(a[827]), .Z(n34010) );
  AND U34886 ( .A(n34011), .B(n34010), .Z(n34064) );
  XOR U34887 ( .A(a[824]), .B(n42197), .Z(n34053) );
  NANDN U34888 ( .A(n34053), .B(n42173), .Z(n34014) );
  NANDN U34889 ( .A(n34012), .B(n42172), .Z(n34013) );
  NAND U34890 ( .A(n34014), .B(n34013), .Z(n34062) );
  NAND U34891 ( .A(b[7]), .B(a[820]), .Z(n34063) );
  XNOR U34892 ( .A(n34062), .B(n34063), .Z(n34065) );
  XOR U34893 ( .A(n34064), .B(n34065), .Z(n34071) );
  NANDN U34894 ( .A(n34015), .B(n42093), .Z(n34017) );
  XOR U34895 ( .A(n42134), .B(a[826]), .Z(n34056) );
  NANDN U34896 ( .A(n34056), .B(n42095), .Z(n34016) );
  NAND U34897 ( .A(n34017), .B(n34016), .Z(n34069) );
  NANDN U34898 ( .A(n34018), .B(n42231), .Z(n34020) );
  XOR U34899 ( .A(n230), .B(a[822]), .Z(n34059) );
  NANDN U34900 ( .A(n34059), .B(n42234), .Z(n34019) );
  AND U34901 ( .A(n34020), .B(n34019), .Z(n34068) );
  XNOR U34902 ( .A(n34069), .B(n34068), .Z(n34070) );
  XNOR U34903 ( .A(n34071), .B(n34070), .Z(n34075) );
  NANDN U34904 ( .A(n34022), .B(n34021), .Z(n34026) );
  NAND U34905 ( .A(n34024), .B(n34023), .Z(n34025) );
  AND U34906 ( .A(n34026), .B(n34025), .Z(n34074) );
  XOR U34907 ( .A(n34075), .B(n34074), .Z(n34076) );
  NANDN U34908 ( .A(n34028), .B(n34027), .Z(n34032) );
  NANDN U34909 ( .A(n34030), .B(n34029), .Z(n34031) );
  NAND U34910 ( .A(n34032), .B(n34031), .Z(n34077) );
  XOR U34911 ( .A(n34076), .B(n34077), .Z(n34044) );
  OR U34912 ( .A(n34034), .B(n34033), .Z(n34038) );
  NANDN U34913 ( .A(n34036), .B(n34035), .Z(n34037) );
  NAND U34914 ( .A(n34038), .B(n34037), .Z(n34045) );
  XNOR U34915 ( .A(n34044), .B(n34045), .Z(n34046) );
  XNOR U34916 ( .A(n34047), .B(n34046), .Z(n34080) );
  XNOR U34917 ( .A(n34080), .B(sreg[1844]), .Z(n34082) );
  NAND U34918 ( .A(n34039), .B(sreg[1843]), .Z(n34043) );
  OR U34919 ( .A(n34041), .B(n34040), .Z(n34042) );
  AND U34920 ( .A(n34043), .B(n34042), .Z(n34081) );
  XOR U34921 ( .A(n34082), .B(n34081), .Z(c[1844]) );
  NANDN U34922 ( .A(n34045), .B(n34044), .Z(n34049) );
  NAND U34923 ( .A(n34047), .B(n34046), .Z(n34048) );
  NAND U34924 ( .A(n34049), .B(n34048), .Z(n34088) );
  NAND U34925 ( .A(b[0]), .B(a[829]), .Z(n34050) );
  XNOR U34926 ( .A(b[1]), .B(n34050), .Z(n34052) );
  NAND U34927 ( .A(n133), .B(a[828]), .Z(n34051) );
  AND U34928 ( .A(n34052), .B(n34051), .Z(n34105) );
  XOR U34929 ( .A(a[825]), .B(n42197), .Z(n34094) );
  NANDN U34930 ( .A(n34094), .B(n42173), .Z(n34055) );
  NANDN U34931 ( .A(n34053), .B(n42172), .Z(n34054) );
  NAND U34932 ( .A(n34055), .B(n34054), .Z(n34103) );
  NAND U34933 ( .A(b[7]), .B(a[821]), .Z(n34104) );
  XNOR U34934 ( .A(n34103), .B(n34104), .Z(n34106) );
  XOR U34935 ( .A(n34105), .B(n34106), .Z(n34112) );
  NANDN U34936 ( .A(n34056), .B(n42093), .Z(n34058) );
  XOR U34937 ( .A(n42134), .B(a[827]), .Z(n34097) );
  NANDN U34938 ( .A(n34097), .B(n42095), .Z(n34057) );
  NAND U34939 ( .A(n34058), .B(n34057), .Z(n34110) );
  NANDN U34940 ( .A(n34059), .B(n42231), .Z(n34061) );
  XOR U34941 ( .A(n230), .B(a[823]), .Z(n34100) );
  NANDN U34942 ( .A(n34100), .B(n42234), .Z(n34060) );
  AND U34943 ( .A(n34061), .B(n34060), .Z(n34109) );
  XNOR U34944 ( .A(n34110), .B(n34109), .Z(n34111) );
  XNOR U34945 ( .A(n34112), .B(n34111), .Z(n34116) );
  NANDN U34946 ( .A(n34063), .B(n34062), .Z(n34067) );
  NAND U34947 ( .A(n34065), .B(n34064), .Z(n34066) );
  AND U34948 ( .A(n34067), .B(n34066), .Z(n34115) );
  XOR U34949 ( .A(n34116), .B(n34115), .Z(n34117) );
  NANDN U34950 ( .A(n34069), .B(n34068), .Z(n34073) );
  NANDN U34951 ( .A(n34071), .B(n34070), .Z(n34072) );
  NAND U34952 ( .A(n34073), .B(n34072), .Z(n34118) );
  XOR U34953 ( .A(n34117), .B(n34118), .Z(n34085) );
  OR U34954 ( .A(n34075), .B(n34074), .Z(n34079) );
  NANDN U34955 ( .A(n34077), .B(n34076), .Z(n34078) );
  NAND U34956 ( .A(n34079), .B(n34078), .Z(n34086) );
  XNOR U34957 ( .A(n34085), .B(n34086), .Z(n34087) );
  XNOR U34958 ( .A(n34088), .B(n34087), .Z(n34121) );
  XNOR U34959 ( .A(n34121), .B(sreg[1845]), .Z(n34123) );
  NAND U34960 ( .A(n34080), .B(sreg[1844]), .Z(n34084) );
  OR U34961 ( .A(n34082), .B(n34081), .Z(n34083) );
  AND U34962 ( .A(n34084), .B(n34083), .Z(n34122) );
  XOR U34963 ( .A(n34123), .B(n34122), .Z(c[1845]) );
  NANDN U34964 ( .A(n34086), .B(n34085), .Z(n34090) );
  NAND U34965 ( .A(n34088), .B(n34087), .Z(n34089) );
  NAND U34966 ( .A(n34090), .B(n34089), .Z(n34129) );
  NAND U34967 ( .A(b[0]), .B(a[830]), .Z(n34091) );
  XNOR U34968 ( .A(b[1]), .B(n34091), .Z(n34093) );
  NAND U34969 ( .A(n133), .B(a[829]), .Z(n34092) );
  AND U34970 ( .A(n34093), .B(n34092), .Z(n34146) );
  XOR U34971 ( .A(a[826]), .B(n42197), .Z(n34135) );
  NANDN U34972 ( .A(n34135), .B(n42173), .Z(n34096) );
  NANDN U34973 ( .A(n34094), .B(n42172), .Z(n34095) );
  NAND U34974 ( .A(n34096), .B(n34095), .Z(n34144) );
  NAND U34975 ( .A(b[7]), .B(a[822]), .Z(n34145) );
  XNOR U34976 ( .A(n34144), .B(n34145), .Z(n34147) );
  XOR U34977 ( .A(n34146), .B(n34147), .Z(n34153) );
  NANDN U34978 ( .A(n34097), .B(n42093), .Z(n34099) );
  XOR U34979 ( .A(n42134), .B(a[828]), .Z(n34138) );
  NANDN U34980 ( .A(n34138), .B(n42095), .Z(n34098) );
  NAND U34981 ( .A(n34099), .B(n34098), .Z(n34151) );
  NANDN U34982 ( .A(n34100), .B(n42231), .Z(n34102) );
  XOR U34983 ( .A(n230), .B(a[824]), .Z(n34141) );
  NANDN U34984 ( .A(n34141), .B(n42234), .Z(n34101) );
  AND U34985 ( .A(n34102), .B(n34101), .Z(n34150) );
  XNOR U34986 ( .A(n34151), .B(n34150), .Z(n34152) );
  XNOR U34987 ( .A(n34153), .B(n34152), .Z(n34157) );
  NANDN U34988 ( .A(n34104), .B(n34103), .Z(n34108) );
  NAND U34989 ( .A(n34106), .B(n34105), .Z(n34107) );
  AND U34990 ( .A(n34108), .B(n34107), .Z(n34156) );
  XOR U34991 ( .A(n34157), .B(n34156), .Z(n34158) );
  NANDN U34992 ( .A(n34110), .B(n34109), .Z(n34114) );
  NANDN U34993 ( .A(n34112), .B(n34111), .Z(n34113) );
  NAND U34994 ( .A(n34114), .B(n34113), .Z(n34159) );
  XOR U34995 ( .A(n34158), .B(n34159), .Z(n34126) );
  OR U34996 ( .A(n34116), .B(n34115), .Z(n34120) );
  NANDN U34997 ( .A(n34118), .B(n34117), .Z(n34119) );
  NAND U34998 ( .A(n34120), .B(n34119), .Z(n34127) );
  XNOR U34999 ( .A(n34126), .B(n34127), .Z(n34128) );
  XNOR U35000 ( .A(n34129), .B(n34128), .Z(n34162) );
  XNOR U35001 ( .A(n34162), .B(sreg[1846]), .Z(n34164) );
  NAND U35002 ( .A(n34121), .B(sreg[1845]), .Z(n34125) );
  OR U35003 ( .A(n34123), .B(n34122), .Z(n34124) );
  AND U35004 ( .A(n34125), .B(n34124), .Z(n34163) );
  XOR U35005 ( .A(n34164), .B(n34163), .Z(c[1846]) );
  NANDN U35006 ( .A(n34127), .B(n34126), .Z(n34131) );
  NAND U35007 ( .A(n34129), .B(n34128), .Z(n34130) );
  NAND U35008 ( .A(n34131), .B(n34130), .Z(n34170) );
  NAND U35009 ( .A(b[0]), .B(a[831]), .Z(n34132) );
  XNOR U35010 ( .A(b[1]), .B(n34132), .Z(n34134) );
  NAND U35011 ( .A(n133), .B(a[830]), .Z(n34133) );
  AND U35012 ( .A(n34134), .B(n34133), .Z(n34187) );
  XOR U35013 ( .A(a[827]), .B(n42197), .Z(n34176) );
  NANDN U35014 ( .A(n34176), .B(n42173), .Z(n34137) );
  NANDN U35015 ( .A(n34135), .B(n42172), .Z(n34136) );
  NAND U35016 ( .A(n34137), .B(n34136), .Z(n34185) );
  NAND U35017 ( .A(b[7]), .B(a[823]), .Z(n34186) );
  XNOR U35018 ( .A(n34185), .B(n34186), .Z(n34188) );
  XOR U35019 ( .A(n34187), .B(n34188), .Z(n34194) );
  NANDN U35020 ( .A(n34138), .B(n42093), .Z(n34140) );
  XOR U35021 ( .A(n42134), .B(a[829]), .Z(n34179) );
  NANDN U35022 ( .A(n34179), .B(n42095), .Z(n34139) );
  NAND U35023 ( .A(n34140), .B(n34139), .Z(n34192) );
  NANDN U35024 ( .A(n34141), .B(n42231), .Z(n34143) );
  XOR U35025 ( .A(n230), .B(a[825]), .Z(n34182) );
  NANDN U35026 ( .A(n34182), .B(n42234), .Z(n34142) );
  AND U35027 ( .A(n34143), .B(n34142), .Z(n34191) );
  XNOR U35028 ( .A(n34192), .B(n34191), .Z(n34193) );
  XNOR U35029 ( .A(n34194), .B(n34193), .Z(n34198) );
  NANDN U35030 ( .A(n34145), .B(n34144), .Z(n34149) );
  NAND U35031 ( .A(n34147), .B(n34146), .Z(n34148) );
  AND U35032 ( .A(n34149), .B(n34148), .Z(n34197) );
  XOR U35033 ( .A(n34198), .B(n34197), .Z(n34199) );
  NANDN U35034 ( .A(n34151), .B(n34150), .Z(n34155) );
  NANDN U35035 ( .A(n34153), .B(n34152), .Z(n34154) );
  NAND U35036 ( .A(n34155), .B(n34154), .Z(n34200) );
  XOR U35037 ( .A(n34199), .B(n34200), .Z(n34167) );
  OR U35038 ( .A(n34157), .B(n34156), .Z(n34161) );
  NANDN U35039 ( .A(n34159), .B(n34158), .Z(n34160) );
  NAND U35040 ( .A(n34161), .B(n34160), .Z(n34168) );
  XNOR U35041 ( .A(n34167), .B(n34168), .Z(n34169) );
  XNOR U35042 ( .A(n34170), .B(n34169), .Z(n34203) );
  XNOR U35043 ( .A(n34203), .B(sreg[1847]), .Z(n34205) );
  NAND U35044 ( .A(n34162), .B(sreg[1846]), .Z(n34166) );
  OR U35045 ( .A(n34164), .B(n34163), .Z(n34165) );
  AND U35046 ( .A(n34166), .B(n34165), .Z(n34204) );
  XOR U35047 ( .A(n34205), .B(n34204), .Z(c[1847]) );
  NANDN U35048 ( .A(n34168), .B(n34167), .Z(n34172) );
  NAND U35049 ( .A(n34170), .B(n34169), .Z(n34171) );
  NAND U35050 ( .A(n34172), .B(n34171), .Z(n34211) );
  NAND U35051 ( .A(b[0]), .B(a[832]), .Z(n34173) );
  XNOR U35052 ( .A(b[1]), .B(n34173), .Z(n34175) );
  NAND U35053 ( .A(n133), .B(a[831]), .Z(n34174) );
  AND U35054 ( .A(n34175), .B(n34174), .Z(n34228) );
  XOR U35055 ( .A(a[828]), .B(n42197), .Z(n34217) );
  NANDN U35056 ( .A(n34217), .B(n42173), .Z(n34178) );
  NANDN U35057 ( .A(n34176), .B(n42172), .Z(n34177) );
  NAND U35058 ( .A(n34178), .B(n34177), .Z(n34226) );
  NAND U35059 ( .A(b[7]), .B(a[824]), .Z(n34227) );
  XNOR U35060 ( .A(n34226), .B(n34227), .Z(n34229) );
  XOR U35061 ( .A(n34228), .B(n34229), .Z(n34235) );
  NANDN U35062 ( .A(n34179), .B(n42093), .Z(n34181) );
  XOR U35063 ( .A(n42134), .B(a[830]), .Z(n34220) );
  NANDN U35064 ( .A(n34220), .B(n42095), .Z(n34180) );
  NAND U35065 ( .A(n34181), .B(n34180), .Z(n34233) );
  NANDN U35066 ( .A(n34182), .B(n42231), .Z(n34184) );
  XOR U35067 ( .A(n230), .B(a[826]), .Z(n34223) );
  NANDN U35068 ( .A(n34223), .B(n42234), .Z(n34183) );
  AND U35069 ( .A(n34184), .B(n34183), .Z(n34232) );
  XNOR U35070 ( .A(n34233), .B(n34232), .Z(n34234) );
  XNOR U35071 ( .A(n34235), .B(n34234), .Z(n34239) );
  NANDN U35072 ( .A(n34186), .B(n34185), .Z(n34190) );
  NAND U35073 ( .A(n34188), .B(n34187), .Z(n34189) );
  AND U35074 ( .A(n34190), .B(n34189), .Z(n34238) );
  XOR U35075 ( .A(n34239), .B(n34238), .Z(n34240) );
  NANDN U35076 ( .A(n34192), .B(n34191), .Z(n34196) );
  NANDN U35077 ( .A(n34194), .B(n34193), .Z(n34195) );
  NAND U35078 ( .A(n34196), .B(n34195), .Z(n34241) );
  XOR U35079 ( .A(n34240), .B(n34241), .Z(n34208) );
  OR U35080 ( .A(n34198), .B(n34197), .Z(n34202) );
  NANDN U35081 ( .A(n34200), .B(n34199), .Z(n34201) );
  NAND U35082 ( .A(n34202), .B(n34201), .Z(n34209) );
  XNOR U35083 ( .A(n34208), .B(n34209), .Z(n34210) );
  XNOR U35084 ( .A(n34211), .B(n34210), .Z(n34244) );
  XNOR U35085 ( .A(n34244), .B(sreg[1848]), .Z(n34246) );
  NAND U35086 ( .A(n34203), .B(sreg[1847]), .Z(n34207) );
  OR U35087 ( .A(n34205), .B(n34204), .Z(n34206) );
  AND U35088 ( .A(n34207), .B(n34206), .Z(n34245) );
  XOR U35089 ( .A(n34246), .B(n34245), .Z(c[1848]) );
  NANDN U35090 ( .A(n34209), .B(n34208), .Z(n34213) );
  NAND U35091 ( .A(n34211), .B(n34210), .Z(n34212) );
  NAND U35092 ( .A(n34213), .B(n34212), .Z(n34252) );
  NAND U35093 ( .A(b[0]), .B(a[833]), .Z(n34214) );
  XNOR U35094 ( .A(b[1]), .B(n34214), .Z(n34216) );
  NAND U35095 ( .A(n134), .B(a[832]), .Z(n34215) );
  AND U35096 ( .A(n34216), .B(n34215), .Z(n34269) );
  XOR U35097 ( .A(a[829]), .B(n42197), .Z(n34258) );
  NANDN U35098 ( .A(n34258), .B(n42173), .Z(n34219) );
  NANDN U35099 ( .A(n34217), .B(n42172), .Z(n34218) );
  NAND U35100 ( .A(n34219), .B(n34218), .Z(n34267) );
  NAND U35101 ( .A(b[7]), .B(a[825]), .Z(n34268) );
  XNOR U35102 ( .A(n34267), .B(n34268), .Z(n34270) );
  XOR U35103 ( .A(n34269), .B(n34270), .Z(n34276) );
  NANDN U35104 ( .A(n34220), .B(n42093), .Z(n34222) );
  XOR U35105 ( .A(n42134), .B(a[831]), .Z(n34261) );
  NANDN U35106 ( .A(n34261), .B(n42095), .Z(n34221) );
  NAND U35107 ( .A(n34222), .B(n34221), .Z(n34274) );
  NANDN U35108 ( .A(n34223), .B(n42231), .Z(n34225) );
  XOR U35109 ( .A(n231), .B(a[827]), .Z(n34264) );
  NANDN U35110 ( .A(n34264), .B(n42234), .Z(n34224) );
  AND U35111 ( .A(n34225), .B(n34224), .Z(n34273) );
  XNOR U35112 ( .A(n34274), .B(n34273), .Z(n34275) );
  XNOR U35113 ( .A(n34276), .B(n34275), .Z(n34280) );
  NANDN U35114 ( .A(n34227), .B(n34226), .Z(n34231) );
  NAND U35115 ( .A(n34229), .B(n34228), .Z(n34230) );
  AND U35116 ( .A(n34231), .B(n34230), .Z(n34279) );
  XOR U35117 ( .A(n34280), .B(n34279), .Z(n34281) );
  NANDN U35118 ( .A(n34233), .B(n34232), .Z(n34237) );
  NANDN U35119 ( .A(n34235), .B(n34234), .Z(n34236) );
  NAND U35120 ( .A(n34237), .B(n34236), .Z(n34282) );
  XOR U35121 ( .A(n34281), .B(n34282), .Z(n34249) );
  OR U35122 ( .A(n34239), .B(n34238), .Z(n34243) );
  NANDN U35123 ( .A(n34241), .B(n34240), .Z(n34242) );
  NAND U35124 ( .A(n34243), .B(n34242), .Z(n34250) );
  XNOR U35125 ( .A(n34249), .B(n34250), .Z(n34251) );
  XNOR U35126 ( .A(n34252), .B(n34251), .Z(n34285) );
  XNOR U35127 ( .A(n34285), .B(sreg[1849]), .Z(n34287) );
  NAND U35128 ( .A(n34244), .B(sreg[1848]), .Z(n34248) );
  OR U35129 ( .A(n34246), .B(n34245), .Z(n34247) );
  AND U35130 ( .A(n34248), .B(n34247), .Z(n34286) );
  XOR U35131 ( .A(n34287), .B(n34286), .Z(c[1849]) );
  NANDN U35132 ( .A(n34250), .B(n34249), .Z(n34254) );
  NAND U35133 ( .A(n34252), .B(n34251), .Z(n34253) );
  NAND U35134 ( .A(n34254), .B(n34253), .Z(n34293) );
  NAND U35135 ( .A(b[0]), .B(a[834]), .Z(n34255) );
  XNOR U35136 ( .A(b[1]), .B(n34255), .Z(n34257) );
  NAND U35137 ( .A(n134), .B(a[833]), .Z(n34256) );
  AND U35138 ( .A(n34257), .B(n34256), .Z(n34310) );
  XOR U35139 ( .A(a[830]), .B(n42197), .Z(n34299) );
  NANDN U35140 ( .A(n34299), .B(n42173), .Z(n34260) );
  NANDN U35141 ( .A(n34258), .B(n42172), .Z(n34259) );
  NAND U35142 ( .A(n34260), .B(n34259), .Z(n34308) );
  NAND U35143 ( .A(b[7]), .B(a[826]), .Z(n34309) );
  XNOR U35144 ( .A(n34308), .B(n34309), .Z(n34311) );
  XOR U35145 ( .A(n34310), .B(n34311), .Z(n34317) );
  NANDN U35146 ( .A(n34261), .B(n42093), .Z(n34263) );
  XOR U35147 ( .A(n42134), .B(a[832]), .Z(n34302) );
  NANDN U35148 ( .A(n34302), .B(n42095), .Z(n34262) );
  NAND U35149 ( .A(n34263), .B(n34262), .Z(n34315) );
  NANDN U35150 ( .A(n34264), .B(n42231), .Z(n34266) );
  XOR U35151 ( .A(n231), .B(a[828]), .Z(n34305) );
  NANDN U35152 ( .A(n34305), .B(n42234), .Z(n34265) );
  AND U35153 ( .A(n34266), .B(n34265), .Z(n34314) );
  XNOR U35154 ( .A(n34315), .B(n34314), .Z(n34316) );
  XNOR U35155 ( .A(n34317), .B(n34316), .Z(n34321) );
  NANDN U35156 ( .A(n34268), .B(n34267), .Z(n34272) );
  NAND U35157 ( .A(n34270), .B(n34269), .Z(n34271) );
  AND U35158 ( .A(n34272), .B(n34271), .Z(n34320) );
  XOR U35159 ( .A(n34321), .B(n34320), .Z(n34322) );
  NANDN U35160 ( .A(n34274), .B(n34273), .Z(n34278) );
  NANDN U35161 ( .A(n34276), .B(n34275), .Z(n34277) );
  NAND U35162 ( .A(n34278), .B(n34277), .Z(n34323) );
  XOR U35163 ( .A(n34322), .B(n34323), .Z(n34290) );
  OR U35164 ( .A(n34280), .B(n34279), .Z(n34284) );
  NANDN U35165 ( .A(n34282), .B(n34281), .Z(n34283) );
  NAND U35166 ( .A(n34284), .B(n34283), .Z(n34291) );
  XNOR U35167 ( .A(n34290), .B(n34291), .Z(n34292) );
  XNOR U35168 ( .A(n34293), .B(n34292), .Z(n34326) );
  XNOR U35169 ( .A(n34326), .B(sreg[1850]), .Z(n34328) );
  NAND U35170 ( .A(n34285), .B(sreg[1849]), .Z(n34289) );
  OR U35171 ( .A(n34287), .B(n34286), .Z(n34288) );
  AND U35172 ( .A(n34289), .B(n34288), .Z(n34327) );
  XOR U35173 ( .A(n34328), .B(n34327), .Z(c[1850]) );
  NANDN U35174 ( .A(n34291), .B(n34290), .Z(n34295) );
  NAND U35175 ( .A(n34293), .B(n34292), .Z(n34294) );
  NAND U35176 ( .A(n34295), .B(n34294), .Z(n34334) );
  NAND U35177 ( .A(b[0]), .B(a[835]), .Z(n34296) );
  XNOR U35178 ( .A(b[1]), .B(n34296), .Z(n34298) );
  NAND U35179 ( .A(n134), .B(a[834]), .Z(n34297) );
  AND U35180 ( .A(n34298), .B(n34297), .Z(n34351) );
  XOR U35181 ( .A(a[831]), .B(n42197), .Z(n34340) );
  NANDN U35182 ( .A(n34340), .B(n42173), .Z(n34301) );
  NANDN U35183 ( .A(n34299), .B(n42172), .Z(n34300) );
  NAND U35184 ( .A(n34301), .B(n34300), .Z(n34349) );
  NAND U35185 ( .A(b[7]), .B(a[827]), .Z(n34350) );
  XNOR U35186 ( .A(n34349), .B(n34350), .Z(n34352) );
  XOR U35187 ( .A(n34351), .B(n34352), .Z(n34358) );
  NANDN U35188 ( .A(n34302), .B(n42093), .Z(n34304) );
  XOR U35189 ( .A(n42134), .B(a[833]), .Z(n34343) );
  NANDN U35190 ( .A(n34343), .B(n42095), .Z(n34303) );
  NAND U35191 ( .A(n34304), .B(n34303), .Z(n34356) );
  NANDN U35192 ( .A(n34305), .B(n42231), .Z(n34307) );
  XOR U35193 ( .A(n231), .B(a[829]), .Z(n34346) );
  NANDN U35194 ( .A(n34346), .B(n42234), .Z(n34306) );
  AND U35195 ( .A(n34307), .B(n34306), .Z(n34355) );
  XNOR U35196 ( .A(n34356), .B(n34355), .Z(n34357) );
  XNOR U35197 ( .A(n34358), .B(n34357), .Z(n34362) );
  NANDN U35198 ( .A(n34309), .B(n34308), .Z(n34313) );
  NAND U35199 ( .A(n34311), .B(n34310), .Z(n34312) );
  AND U35200 ( .A(n34313), .B(n34312), .Z(n34361) );
  XOR U35201 ( .A(n34362), .B(n34361), .Z(n34363) );
  NANDN U35202 ( .A(n34315), .B(n34314), .Z(n34319) );
  NANDN U35203 ( .A(n34317), .B(n34316), .Z(n34318) );
  NAND U35204 ( .A(n34319), .B(n34318), .Z(n34364) );
  XOR U35205 ( .A(n34363), .B(n34364), .Z(n34331) );
  OR U35206 ( .A(n34321), .B(n34320), .Z(n34325) );
  NANDN U35207 ( .A(n34323), .B(n34322), .Z(n34324) );
  NAND U35208 ( .A(n34325), .B(n34324), .Z(n34332) );
  XNOR U35209 ( .A(n34331), .B(n34332), .Z(n34333) );
  XNOR U35210 ( .A(n34334), .B(n34333), .Z(n34367) );
  XNOR U35211 ( .A(n34367), .B(sreg[1851]), .Z(n34369) );
  NAND U35212 ( .A(n34326), .B(sreg[1850]), .Z(n34330) );
  OR U35213 ( .A(n34328), .B(n34327), .Z(n34329) );
  AND U35214 ( .A(n34330), .B(n34329), .Z(n34368) );
  XOR U35215 ( .A(n34369), .B(n34368), .Z(c[1851]) );
  NANDN U35216 ( .A(n34332), .B(n34331), .Z(n34336) );
  NAND U35217 ( .A(n34334), .B(n34333), .Z(n34335) );
  NAND U35218 ( .A(n34336), .B(n34335), .Z(n34375) );
  NAND U35219 ( .A(b[0]), .B(a[836]), .Z(n34337) );
  XNOR U35220 ( .A(b[1]), .B(n34337), .Z(n34339) );
  NAND U35221 ( .A(n134), .B(a[835]), .Z(n34338) );
  AND U35222 ( .A(n34339), .B(n34338), .Z(n34392) );
  XOR U35223 ( .A(a[832]), .B(n42197), .Z(n34381) );
  NANDN U35224 ( .A(n34381), .B(n42173), .Z(n34342) );
  NANDN U35225 ( .A(n34340), .B(n42172), .Z(n34341) );
  NAND U35226 ( .A(n34342), .B(n34341), .Z(n34390) );
  NAND U35227 ( .A(b[7]), .B(a[828]), .Z(n34391) );
  XNOR U35228 ( .A(n34390), .B(n34391), .Z(n34393) );
  XOR U35229 ( .A(n34392), .B(n34393), .Z(n34399) );
  NANDN U35230 ( .A(n34343), .B(n42093), .Z(n34345) );
  XOR U35231 ( .A(n42134), .B(a[834]), .Z(n34384) );
  NANDN U35232 ( .A(n34384), .B(n42095), .Z(n34344) );
  NAND U35233 ( .A(n34345), .B(n34344), .Z(n34397) );
  NANDN U35234 ( .A(n34346), .B(n42231), .Z(n34348) );
  XOR U35235 ( .A(n231), .B(a[830]), .Z(n34387) );
  NANDN U35236 ( .A(n34387), .B(n42234), .Z(n34347) );
  AND U35237 ( .A(n34348), .B(n34347), .Z(n34396) );
  XNOR U35238 ( .A(n34397), .B(n34396), .Z(n34398) );
  XNOR U35239 ( .A(n34399), .B(n34398), .Z(n34403) );
  NANDN U35240 ( .A(n34350), .B(n34349), .Z(n34354) );
  NAND U35241 ( .A(n34352), .B(n34351), .Z(n34353) );
  AND U35242 ( .A(n34354), .B(n34353), .Z(n34402) );
  XOR U35243 ( .A(n34403), .B(n34402), .Z(n34404) );
  NANDN U35244 ( .A(n34356), .B(n34355), .Z(n34360) );
  NANDN U35245 ( .A(n34358), .B(n34357), .Z(n34359) );
  NAND U35246 ( .A(n34360), .B(n34359), .Z(n34405) );
  XOR U35247 ( .A(n34404), .B(n34405), .Z(n34372) );
  OR U35248 ( .A(n34362), .B(n34361), .Z(n34366) );
  NANDN U35249 ( .A(n34364), .B(n34363), .Z(n34365) );
  NAND U35250 ( .A(n34366), .B(n34365), .Z(n34373) );
  XNOR U35251 ( .A(n34372), .B(n34373), .Z(n34374) );
  XNOR U35252 ( .A(n34375), .B(n34374), .Z(n34408) );
  XNOR U35253 ( .A(n34408), .B(sreg[1852]), .Z(n34410) );
  NAND U35254 ( .A(n34367), .B(sreg[1851]), .Z(n34371) );
  OR U35255 ( .A(n34369), .B(n34368), .Z(n34370) );
  AND U35256 ( .A(n34371), .B(n34370), .Z(n34409) );
  XOR U35257 ( .A(n34410), .B(n34409), .Z(c[1852]) );
  NANDN U35258 ( .A(n34373), .B(n34372), .Z(n34377) );
  NAND U35259 ( .A(n34375), .B(n34374), .Z(n34376) );
  NAND U35260 ( .A(n34377), .B(n34376), .Z(n34416) );
  NAND U35261 ( .A(b[0]), .B(a[837]), .Z(n34378) );
  XNOR U35262 ( .A(b[1]), .B(n34378), .Z(n34380) );
  NAND U35263 ( .A(n134), .B(a[836]), .Z(n34379) );
  AND U35264 ( .A(n34380), .B(n34379), .Z(n34433) );
  XOR U35265 ( .A(a[833]), .B(n42197), .Z(n34422) );
  NANDN U35266 ( .A(n34422), .B(n42173), .Z(n34383) );
  NANDN U35267 ( .A(n34381), .B(n42172), .Z(n34382) );
  NAND U35268 ( .A(n34383), .B(n34382), .Z(n34431) );
  NAND U35269 ( .A(b[7]), .B(a[829]), .Z(n34432) );
  XNOR U35270 ( .A(n34431), .B(n34432), .Z(n34434) );
  XOR U35271 ( .A(n34433), .B(n34434), .Z(n34440) );
  NANDN U35272 ( .A(n34384), .B(n42093), .Z(n34386) );
  XOR U35273 ( .A(n42134), .B(a[835]), .Z(n34425) );
  NANDN U35274 ( .A(n34425), .B(n42095), .Z(n34385) );
  NAND U35275 ( .A(n34386), .B(n34385), .Z(n34438) );
  NANDN U35276 ( .A(n34387), .B(n42231), .Z(n34389) );
  XOR U35277 ( .A(n231), .B(a[831]), .Z(n34428) );
  NANDN U35278 ( .A(n34428), .B(n42234), .Z(n34388) );
  AND U35279 ( .A(n34389), .B(n34388), .Z(n34437) );
  XNOR U35280 ( .A(n34438), .B(n34437), .Z(n34439) );
  XNOR U35281 ( .A(n34440), .B(n34439), .Z(n34444) );
  NANDN U35282 ( .A(n34391), .B(n34390), .Z(n34395) );
  NAND U35283 ( .A(n34393), .B(n34392), .Z(n34394) );
  AND U35284 ( .A(n34395), .B(n34394), .Z(n34443) );
  XOR U35285 ( .A(n34444), .B(n34443), .Z(n34445) );
  NANDN U35286 ( .A(n34397), .B(n34396), .Z(n34401) );
  NANDN U35287 ( .A(n34399), .B(n34398), .Z(n34400) );
  NAND U35288 ( .A(n34401), .B(n34400), .Z(n34446) );
  XOR U35289 ( .A(n34445), .B(n34446), .Z(n34413) );
  OR U35290 ( .A(n34403), .B(n34402), .Z(n34407) );
  NANDN U35291 ( .A(n34405), .B(n34404), .Z(n34406) );
  NAND U35292 ( .A(n34407), .B(n34406), .Z(n34414) );
  XNOR U35293 ( .A(n34413), .B(n34414), .Z(n34415) );
  XNOR U35294 ( .A(n34416), .B(n34415), .Z(n34449) );
  XNOR U35295 ( .A(n34449), .B(sreg[1853]), .Z(n34451) );
  NAND U35296 ( .A(n34408), .B(sreg[1852]), .Z(n34412) );
  OR U35297 ( .A(n34410), .B(n34409), .Z(n34411) );
  AND U35298 ( .A(n34412), .B(n34411), .Z(n34450) );
  XOR U35299 ( .A(n34451), .B(n34450), .Z(c[1853]) );
  NANDN U35300 ( .A(n34414), .B(n34413), .Z(n34418) );
  NAND U35301 ( .A(n34416), .B(n34415), .Z(n34417) );
  NAND U35302 ( .A(n34418), .B(n34417), .Z(n34457) );
  NAND U35303 ( .A(b[0]), .B(a[838]), .Z(n34419) );
  XNOR U35304 ( .A(b[1]), .B(n34419), .Z(n34421) );
  NAND U35305 ( .A(n134), .B(a[837]), .Z(n34420) );
  AND U35306 ( .A(n34421), .B(n34420), .Z(n34474) );
  XOR U35307 ( .A(a[834]), .B(n42197), .Z(n34463) );
  NANDN U35308 ( .A(n34463), .B(n42173), .Z(n34424) );
  NANDN U35309 ( .A(n34422), .B(n42172), .Z(n34423) );
  NAND U35310 ( .A(n34424), .B(n34423), .Z(n34472) );
  NAND U35311 ( .A(b[7]), .B(a[830]), .Z(n34473) );
  XNOR U35312 ( .A(n34472), .B(n34473), .Z(n34475) );
  XOR U35313 ( .A(n34474), .B(n34475), .Z(n34481) );
  NANDN U35314 ( .A(n34425), .B(n42093), .Z(n34427) );
  XOR U35315 ( .A(n42134), .B(a[836]), .Z(n34466) );
  NANDN U35316 ( .A(n34466), .B(n42095), .Z(n34426) );
  NAND U35317 ( .A(n34427), .B(n34426), .Z(n34479) );
  NANDN U35318 ( .A(n34428), .B(n42231), .Z(n34430) );
  XOR U35319 ( .A(n231), .B(a[832]), .Z(n34469) );
  NANDN U35320 ( .A(n34469), .B(n42234), .Z(n34429) );
  AND U35321 ( .A(n34430), .B(n34429), .Z(n34478) );
  XNOR U35322 ( .A(n34479), .B(n34478), .Z(n34480) );
  XNOR U35323 ( .A(n34481), .B(n34480), .Z(n34485) );
  NANDN U35324 ( .A(n34432), .B(n34431), .Z(n34436) );
  NAND U35325 ( .A(n34434), .B(n34433), .Z(n34435) );
  AND U35326 ( .A(n34436), .B(n34435), .Z(n34484) );
  XOR U35327 ( .A(n34485), .B(n34484), .Z(n34486) );
  NANDN U35328 ( .A(n34438), .B(n34437), .Z(n34442) );
  NANDN U35329 ( .A(n34440), .B(n34439), .Z(n34441) );
  NAND U35330 ( .A(n34442), .B(n34441), .Z(n34487) );
  XOR U35331 ( .A(n34486), .B(n34487), .Z(n34454) );
  OR U35332 ( .A(n34444), .B(n34443), .Z(n34448) );
  NANDN U35333 ( .A(n34446), .B(n34445), .Z(n34447) );
  NAND U35334 ( .A(n34448), .B(n34447), .Z(n34455) );
  XNOR U35335 ( .A(n34454), .B(n34455), .Z(n34456) );
  XNOR U35336 ( .A(n34457), .B(n34456), .Z(n34490) );
  XNOR U35337 ( .A(n34490), .B(sreg[1854]), .Z(n34492) );
  NAND U35338 ( .A(n34449), .B(sreg[1853]), .Z(n34453) );
  OR U35339 ( .A(n34451), .B(n34450), .Z(n34452) );
  AND U35340 ( .A(n34453), .B(n34452), .Z(n34491) );
  XOR U35341 ( .A(n34492), .B(n34491), .Z(c[1854]) );
  NANDN U35342 ( .A(n34455), .B(n34454), .Z(n34459) );
  NAND U35343 ( .A(n34457), .B(n34456), .Z(n34458) );
  NAND U35344 ( .A(n34459), .B(n34458), .Z(n34498) );
  NAND U35345 ( .A(b[0]), .B(a[839]), .Z(n34460) );
  XNOR U35346 ( .A(b[1]), .B(n34460), .Z(n34462) );
  NAND U35347 ( .A(n134), .B(a[838]), .Z(n34461) );
  AND U35348 ( .A(n34462), .B(n34461), .Z(n34515) );
  XOR U35349 ( .A(a[835]), .B(n42197), .Z(n34504) );
  NANDN U35350 ( .A(n34504), .B(n42173), .Z(n34465) );
  NANDN U35351 ( .A(n34463), .B(n42172), .Z(n34464) );
  NAND U35352 ( .A(n34465), .B(n34464), .Z(n34513) );
  NAND U35353 ( .A(b[7]), .B(a[831]), .Z(n34514) );
  XNOR U35354 ( .A(n34513), .B(n34514), .Z(n34516) );
  XOR U35355 ( .A(n34515), .B(n34516), .Z(n34522) );
  NANDN U35356 ( .A(n34466), .B(n42093), .Z(n34468) );
  XOR U35357 ( .A(n42134), .B(a[837]), .Z(n34507) );
  NANDN U35358 ( .A(n34507), .B(n42095), .Z(n34467) );
  NAND U35359 ( .A(n34468), .B(n34467), .Z(n34520) );
  NANDN U35360 ( .A(n34469), .B(n42231), .Z(n34471) );
  XOR U35361 ( .A(n231), .B(a[833]), .Z(n34510) );
  NANDN U35362 ( .A(n34510), .B(n42234), .Z(n34470) );
  AND U35363 ( .A(n34471), .B(n34470), .Z(n34519) );
  XNOR U35364 ( .A(n34520), .B(n34519), .Z(n34521) );
  XNOR U35365 ( .A(n34522), .B(n34521), .Z(n34526) );
  NANDN U35366 ( .A(n34473), .B(n34472), .Z(n34477) );
  NAND U35367 ( .A(n34475), .B(n34474), .Z(n34476) );
  AND U35368 ( .A(n34477), .B(n34476), .Z(n34525) );
  XOR U35369 ( .A(n34526), .B(n34525), .Z(n34527) );
  NANDN U35370 ( .A(n34479), .B(n34478), .Z(n34483) );
  NANDN U35371 ( .A(n34481), .B(n34480), .Z(n34482) );
  NAND U35372 ( .A(n34483), .B(n34482), .Z(n34528) );
  XOR U35373 ( .A(n34527), .B(n34528), .Z(n34495) );
  OR U35374 ( .A(n34485), .B(n34484), .Z(n34489) );
  NANDN U35375 ( .A(n34487), .B(n34486), .Z(n34488) );
  NAND U35376 ( .A(n34489), .B(n34488), .Z(n34496) );
  XNOR U35377 ( .A(n34495), .B(n34496), .Z(n34497) );
  XNOR U35378 ( .A(n34498), .B(n34497), .Z(n34531) );
  XNOR U35379 ( .A(n34531), .B(sreg[1855]), .Z(n34533) );
  NAND U35380 ( .A(n34490), .B(sreg[1854]), .Z(n34494) );
  OR U35381 ( .A(n34492), .B(n34491), .Z(n34493) );
  AND U35382 ( .A(n34494), .B(n34493), .Z(n34532) );
  XOR U35383 ( .A(n34533), .B(n34532), .Z(c[1855]) );
  NANDN U35384 ( .A(n34496), .B(n34495), .Z(n34500) );
  NAND U35385 ( .A(n34498), .B(n34497), .Z(n34499) );
  NAND U35386 ( .A(n34500), .B(n34499), .Z(n34539) );
  NAND U35387 ( .A(b[0]), .B(a[840]), .Z(n34501) );
  XNOR U35388 ( .A(b[1]), .B(n34501), .Z(n34503) );
  NAND U35389 ( .A(n135), .B(a[839]), .Z(n34502) );
  AND U35390 ( .A(n34503), .B(n34502), .Z(n34556) );
  XOR U35391 ( .A(a[836]), .B(n42197), .Z(n34545) );
  NANDN U35392 ( .A(n34545), .B(n42173), .Z(n34506) );
  NANDN U35393 ( .A(n34504), .B(n42172), .Z(n34505) );
  NAND U35394 ( .A(n34506), .B(n34505), .Z(n34554) );
  NAND U35395 ( .A(b[7]), .B(a[832]), .Z(n34555) );
  XNOR U35396 ( .A(n34554), .B(n34555), .Z(n34557) );
  XOR U35397 ( .A(n34556), .B(n34557), .Z(n34563) );
  NANDN U35398 ( .A(n34507), .B(n42093), .Z(n34509) );
  XOR U35399 ( .A(n42134), .B(a[838]), .Z(n34548) );
  NANDN U35400 ( .A(n34548), .B(n42095), .Z(n34508) );
  NAND U35401 ( .A(n34509), .B(n34508), .Z(n34561) );
  NANDN U35402 ( .A(n34510), .B(n42231), .Z(n34512) );
  XOR U35403 ( .A(n231), .B(a[834]), .Z(n34551) );
  NANDN U35404 ( .A(n34551), .B(n42234), .Z(n34511) );
  AND U35405 ( .A(n34512), .B(n34511), .Z(n34560) );
  XNOR U35406 ( .A(n34561), .B(n34560), .Z(n34562) );
  XNOR U35407 ( .A(n34563), .B(n34562), .Z(n34567) );
  NANDN U35408 ( .A(n34514), .B(n34513), .Z(n34518) );
  NAND U35409 ( .A(n34516), .B(n34515), .Z(n34517) );
  AND U35410 ( .A(n34518), .B(n34517), .Z(n34566) );
  XOR U35411 ( .A(n34567), .B(n34566), .Z(n34568) );
  NANDN U35412 ( .A(n34520), .B(n34519), .Z(n34524) );
  NANDN U35413 ( .A(n34522), .B(n34521), .Z(n34523) );
  NAND U35414 ( .A(n34524), .B(n34523), .Z(n34569) );
  XOR U35415 ( .A(n34568), .B(n34569), .Z(n34536) );
  OR U35416 ( .A(n34526), .B(n34525), .Z(n34530) );
  NANDN U35417 ( .A(n34528), .B(n34527), .Z(n34529) );
  NAND U35418 ( .A(n34530), .B(n34529), .Z(n34537) );
  XNOR U35419 ( .A(n34536), .B(n34537), .Z(n34538) );
  XNOR U35420 ( .A(n34539), .B(n34538), .Z(n34572) );
  XNOR U35421 ( .A(n34572), .B(sreg[1856]), .Z(n34574) );
  NAND U35422 ( .A(n34531), .B(sreg[1855]), .Z(n34535) );
  OR U35423 ( .A(n34533), .B(n34532), .Z(n34534) );
  AND U35424 ( .A(n34535), .B(n34534), .Z(n34573) );
  XOR U35425 ( .A(n34574), .B(n34573), .Z(c[1856]) );
  NANDN U35426 ( .A(n34537), .B(n34536), .Z(n34541) );
  NAND U35427 ( .A(n34539), .B(n34538), .Z(n34540) );
  NAND U35428 ( .A(n34541), .B(n34540), .Z(n34580) );
  NAND U35429 ( .A(b[0]), .B(a[841]), .Z(n34542) );
  XNOR U35430 ( .A(b[1]), .B(n34542), .Z(n34544) );
  NAND U35431 ( .A(n135), .B(a[840]), .Z(n34543) );
  AND U35432 ( .A(n34544), .B(n34543), .Z(n34597) );
  XOR U35433 ( .A(a[837]), .B(n42197), .Z(n34586) );
  NANDN U35434 ( .A(n34586), .B(n42173), .Z(n34547) );
  NANDN U35435 ( .A(n34545), .B(n42172), .Z(n34546) );
  NAND U35436 ( .A(n34547), .B(n34546), .Z(n34595) );
  NAND U35437 ( .A(b[7]), .B(a[833]), .Z(n34596) );
  XNOR U35438 ( .A(n34595), .B(n34596), .Z(n34598) );
  XOR U35439 ( .A(n34597), .B(n34598), .Z(n34604) );
  NANDN U35440 ( .A(n34548), .B(n42093), .Z(n34550) );
  XOR U35441 ( .A(n42134), .B(a[839]), .Z(n34589) );
  NANDN U35442 ( .A(n34589), .B(n42095), .Z(n34549) );
  NAND U35443 ( .A(n34550), .B(n34549), .Z(n34602) );
  NANDN U35444 ( .A(n34551), .B(n42231), .Z(n34553) );
  XOR U35445 ( .A(n231), .B(a[835]), .Z(n34592) );
  NANDN U35446 ( .A(n34592), .B(n42234), .Z(n34552) );
  AND U35447 ( .A(n34553), .B(n34552), .Z(n34601) );
  XNOR U35448 ( .A(n34602), .B(n34601), .Z(n34603) );
  XNOR U35449 ( .A(n34604), .B(n34603), .Z(n34608) );
  NANDN U35450 ( .A(n34555), .B(n34554), .Z(n34559) );
  NAND U35451 ( .A(n34557), .B(n34556), .Z(n34558) );
  AND U35452 ( .A(n34559), .B(n34558), .Z(n34607) );
  XOR U35453 ( .A(n34608), .B(n34607), .Z(n34609) );
  NANDN U35454 ( .A(n34561), .B(n34560), .Z(n34565) );
  NANDN U35455 ( .A(n34563), .B(n34562), .Z(n34564) );
  NAND U35456 ( .A(n34565), .B(n34564), .Z(n34610) );
  XOR U35457 ( .A(n34609), .B(n34610), .Z(n34577) );
  OR U35458 ( .A(n34567), .B(n34566), .Z(n34571) );
  NANDN U35459 ( .A(n34569), .B(n34568), .Z(n34570) );
  NAND U35460 ( .A(n34571), .B(n34570), .Z(n34578) );
  XNOR U35461 ( .A(n34577), .B(n34578), .Z(n34579) );
  XNOR U35462 ( .A(n34580), .B(n34579), .Z(n34613) );
  XNOR U35463 ( .A(n34613), .B(sreg[1857]), .Z(n34615) );
  NAND U35464 ( .A(n34572), .B(sreg[1856]), .Z(n34576) );
  OR U35465 ( .A(n34574), .B(n34573), .Z(n34575) );
  AND U35466 ( .A(n34576), .B(n34575), .Z(n34614) );
  XOR U35467 ( .A(n34615), .B(n34614), .Z(c[1857]) );
  NANDN U35468 ( .A(n34578), .B(n34577), .Z(n34582) );
  NAND U35469 ( .A(n34580), .B(n34579), .Z(n34581) );
  NAND U35470 ( .A(n34582), .B(n34581), .Z(n34621) );
  NAND U35471 ( .A(b[0]), .B(a[842]), .Z(n34583) );
  XNOR U35472 ( .A(b[1]), .B(n34583), .Z(n34585) );
  NAND U35473 ( .A(n135), .B(a[841]), .Z(n34584) );
  AND U35474 ( .A(n34585), .B(n34584), .Z(n34638) );
  XOR U35475 ( .A(a[838]), .B(n42197), .Z(n34627) );
  NANDN U35476 ( .A(n34627), .B(n42173), .Z(n34588) );
  NANDN U35477 ( .A(n34586), .B(n42172), .Z(n34587) );
  NAND U35478 ( .A(n34588), .B(n34587), .Z(n34636) );
  NAND U35479 ( .A(b[7]), .B(a[834]), .Z(n34637) );
  XNOR U35480 ( .A(n34636), .B(n34637), .Z(n34639) );
  XOR U35481 ( .A(n34638), .B(n34639), .Z(n34645) );
  NANDN U35482 ( .A(n34589), .B(n42093), .Z(n34591) );
  XOR U35483 ( .A(n42134), .B(a[840]), .Z(n34630) );
  NANDN U35484 ( .A(n34630), .B(n42095), .Z(n34590) );
  NAND U35485 ( .A(n34591), .B(n34590), .Z(n34643) );
  NANDN U35486 ( .A(n34592), .B(n42231), .Z(n34594) );
  XOR U35487 ( .A(n231), .B(a[836]), .Z(n34633) );
  NANDN U35488 ( .A(n34633), .B(n42234), .Z(n34593) );
  AND U35489 ( .A(n34594), .B(n34593), .Z(n34642) );
  XNOR U35490 ( .A(n34643), .B(n34642), .Z(n34644) );
  XNOR U35491 ( .A(n34645), .B(n34644), .Z(n34649) );
  NANDN U35492 ( .A(n34596), .B(n34595), .Z(n34600) );
  NAND U35493 ( .A(n34598), .B(n34597), .Z(n34599) );
  AND U35494 ( .A(n34600), .B(n34599), .Z(n34648) );
  XOR U35495 ( .A(n34649), .B(n34648), .Z(n34650) );
  NANDN U35496 ( .A(n34602), .B(n34601), .Z(n34606) );
  NANDN U35497 ( .A(n34604), .B(n34603), .Z(n34605) );
  NAND U35498 ( .A(n34606), .B(n34605), .Z(n34651) );
  XOR U35499 ( .A(n34650), .B(n34651), .Z(n34618) );
  OR U35500 ( .A(n34608), .B(n34607), .Z(n34612) );
  NANDN U35501 ( .A(n34610), .B(n34609), .Z(n34611) );
  NAND U35502 ( .A(n34612), .B(n34611), .Z(n34619) );
  XNOR U35503 ( .A(n34618), .B(n34619), .Z(n34620) );
  XNOR U35504 ( .A(n34621), .B(n34620), .Z(n34654) );
  XNOR U35505 ( .A(n34654), .B(sreg[1858]), .Z(n34656) );
  NAND U35506 ( .A(n34613), .B(sreg[1857]), .Z(n34617) );
  OR U35507 ( .A(n34615), .B(n34614), .Z(n34616) );
  AND U35508 ( .A(n34617), .B(n34616), .Z(n34655) );
  XOR U35509 ( .A(n34656), .B(n34655), .Z(c[1858]) );
  NANDN U35510 ( .A(n34619), .B(n34618), .Z(n34623) );
  NAND U35511 ( .A(n34621), .B(n34620), .Z(n34622) );
  NAND U35512 ( .A(n34623), .B(n34622), .Z(n34662) );
  NAND U35513 ( .A(b[0]), .B(a[843]), .Z(n34624) );
  XNOR U35514 ( .A(b[1]), .B(n34624), .Z(n34626) );
  NAND U35515 ( .A(n135), .B(a[842]), .Z(n34625) );
  AND U35516 ( .A(n34626), .B(n34625), .Z(n34679) );
  XOR U35517 ( .A(a[839]), .B(n42197), .Z(n34668) );
  NANDN U35518 ( .A(n34668), .B(n42173), .Z(n34629) );
  NANDN U35519 ( .A(n34627), .B(n42172), .Z(n34628) );
  NAND U35520 ( .A(n34629), .B(n34628), .Z(n34677) );
  NAND U35521 ( .A(b[7]), .B(a[835]), .Z(n34678) );
  XNOR U35522 ( .A(n34677), .B(n34678), .Z(n34680) );
  XOR U35523 ( .A(n34679), .B(n34680), .Z(n34686) );
  NANDN U35524 ( .A(n34630), .B(n42093), .Z(n34632) );
  XOR U35525 ( .A(n42134), .B(a[841]), .Z(n34671) );
  NANDN U35526 ( .A(n34671), .B(n42095), .Z(n34631) );
  NAND U35527 ( .A(n34632), .B(n34631), .Z(n34684) );
  NANDN U35528 ( .A(n34633), .B(n42231), .Z(n34635) );
  XOR U35529 ( .A(n231), .B(a[837]), .Z(n34674) );
  NANDN U35530 ( .A(n34674), .B(n42234), .Z(n34634) );
  AND U35531 ( .A(n34635), .B(n34634), .Z(n34683) );
  XNOR U35532 ( .A(n34684), .B(n34683), .Z(n34685) );
  XNOR U35533 ( .A(n34686), .B(n34685), .Z(n34690) );
  NANDN U35534 ( .A(n34637), .B(n34636), .Z(n34641) );
  NAND U35535 ( .A(n34639), .B(n34638), .Z(n34640) );
  AND U35536 ( .A(n34641), .B(n34640), .Z(n34689) );
  XOR U35537 ( .A(n34690), .B(n34689), .Z(n34691) );
  NANDN U35538 ( .A(n34643), .B(n34642), .Z(n34647) );
  NANDN U35539 ( .A(n34645), .B(n34644), .Z(n34646) );
  NAND U35540 ( .A(n34647), .B(n34646), .Z(n34692) );
  XOR U35541 ( .A(n34691), .B(n34692), .Z(n34659) );
  OR U35542 ( .A(n34649), .B(n34648), .Z(n34653) );
  NANDN U35543 ( .A(n34651), .B(n34650), .Z(n34652) );
  NAND U35544 ( .A(n34653), .B(n34652), .Z(n34660) );
  XNOR U35545 ( .A(n34659), .B(n34660), .Z(n34661) );
  XNOR U35546 ( .A(n34662), .B(n34661), .Z(n34695) );
  XNOR U35547 ( .A(n34695), .B(sreg[1859]), .Z(n34697) );
  NAND U35548 ( .A(n34654), .B(sreg[1858]), .Z(n34658) );
  OR U35549 ( .A(n34656), .B(n34655), .Z(n34657) );
  AND U35550 ( .A(n34658), .B(n34657), .Z(n34696) );
  XOR U35551 ( .A(n34697), .B(n34696), .Z(c[1859]) );
  NANDN U35552 ( .A(n34660), .B(n34659), .Z(n34664) );
  NAND U35553 ( .A(n34662), .B(n34661), .Z(n34663) );
  NAND U35554 ( .A(n34664), .B(n34663), .Z(n34703) );
  NAND U35555 ( .A(b[0]), .B(a[844]), .Z(n34665) );
  XNOR U35556 ( .A(b[1]), .B(n34665), .Z(n34667) );
  NAND U35557 ( .A(n135), .B(a[843]), .Z(n34666) );
  AND U35558 ( .A(n34667), .B(n34666), .Z(n34720) );
  XOR U35559 ( .A(a[840]), .B(n42197), .Z(n34709) );
  NANDN U35560 ( .A(n34709), .B(n42173), .Z(n34670) );
  NANDN U35561 ( .A(n34668), .B(n42172), .Z(n34669) );
  NAND U35562 ( .A(n34670), .B(n34669), .Z(n34718) );
  NAND U35563 ( .A(b[7]), .B(a[836]), .Z(n34719) );
  XNOR U35564 ( .A(n34718), .B(n34719), .Z(n34721) );
  XOR U35565 ( .A(n34720), .B(n34721), .Z(n34727) );
  NANDN U35566 ( .A(n34671), .B(n42093), .Z(n34673) );
  XOR U35567 ( .A(n42134), .B(a[842]), .Z(n34712) );
  NANDN U35568 ( .A(n34712), .B(n42095), .Z(n34672) );
  NAND U35569 ( .A(n34673), .B(n34672), .Z(n34725) );
  NANDN U35570 ( .A(n34674), .B(n42231), .Z(n34676) );
  XOR U35571 ( .A(n231), .B(a[838]), .Z(n34715) );
  NANDN U35572 ( .A(n34715), .B(n42234), .Z(n34675) );
  AND U35573 ( .A(n34676), .B(n34675), .Z(n34724) );
  XNOR U35574 ( .A(n34725), .B(n34724), .Z(n34726) );
  XNOR U35575 ( .A(n34727), .B(n34726), .Z(n34731) );
  NANDN U35576 ( .A(n34678), .B(n34677), .Z(n34682) );
  NAND U35577 ( .A(n34680), .B(n34679), .Z(n34681) );
  AND U35578 ( .A(n34682), .B(n34681), .Z(n34730) );
  XOR U35579 ( .A(n34731), .B(n34730), .Z(n34732) );
  NANDN U35580 ( .A(n34684), .B(n34683), .Z(n34688) );
  NANDN U35581 ( .A(n34686), .B(n34685), .Z(n34687) );
  NAND U35582 ( .A(n34688), .B(n34687), .Z(n34733) );
  XOR U35583 ( .A(n34732), .B(n34733), .Z(n34700) );
  OR U35584 ( .A(n34690), .B(n34689), .Z(n34694) );
  NANDN U35585 ( .A(n34692), .B(n34691), .Z(n34693) );
  NAND U35586 ( .A(n34694), .B(n34693), .Z(n34701) );
  XNOR U35587 ( .A(n34700), .B(n34701), .Z(n34702) );
  XNOR U35588 ( .A(n34703), .B(n34702), .Z(n34736) );
  XNOR U35589 ( .A(n34736), .B(sreg[1860]), .Z(n34738) );
  NAND U35590 ( .A(n34695), .B(sreg[1859]), .Z(n34699) );
  OR U35591 ( .A(n34697), .B(n34696), .Z(n34698) );
  AND U35592 ( .A(n34699), .B(n34698), .Z(n34737) );
  XOR U35593 ( .A(n34738), .B(n34737), .Z(c[1860]) );
  NANDN U35594 ( .A(n34701), .B(n34700), .Z(n34705) );
  NAND U35595 ( .A(n34703), .B(n34702), .Z(n34704) );
  NAND U35596 ( .A(n34705), .B(n34704), .Z(n34744) );
  NAND U35597 ( .A(b[0]), .B(a[845]), .Z(n34706) );
  XNOR U35598 ( .A(b[1]), .B(n34706), .Z(n34708) );
  NAND U35599 ( .A(n135), .B(a[844]), .Z(n34707) );
  AND U35600 ( .A(n34708), .B(n34707), .Z(n34761) );
  XOR U35601 ( .A(a[841]), .B(n42197), .Z(n34750) );
  NANDN U35602 ( .A(n34750), .B(n42173), .Z(n34711) );
  NANDN U35603 ( .A(n34709), .B(n42172), .Z(n34710) );
  NAND U35604 ( .A(n34711), .B(n34710), .Z(n34759) );
  NAND U35605 ( .A(b[7]), .B(a[837]), .Z(n34760) );
  XNOR U35606 ( .A(n34759), .B(n34760), .Z(n34762) );
  XOR U35607 ( .A(n34761), .B(n34762), .Z(n34768) );
  NANDN U35608 ( .A(n34712), .B(n42093), .Z(n34714) );
  XOR U35609 ( .A(n42134), .B(a[843]), .Z(n34753) );
  NANDN U35610 ( .A(n34753), .B(n42095), .Z(n34713) );
  NAND U35611 ( .A(n34714), .B(n34713), .Z(n34766) );
  NANDN U35612 ( .A(n34715), .B(n42231), .Z(n34717) );
  XOR U35613 ( .A(n232), .B(a[839]), .Z(n34756) );
  NANDN U35614 ( .A(n34756), .B(n42234), .Z(n34716) );
  AND U35615 ( .A(n34717), .B(n34716), .Z(n34765) );
  XNOR U35616 ( .A(n34766), .B(n34765), .Z(n34767) );
  XNOR U35617 ( .A(n34768), .B(n34767), .Z(n34772) );
  NANDN U35618 ( .A(n34719), .B(n34718), .Z(n34723) );
  NAND U35619 ( .A(n34721), .B(n34720), .Z(n34722) );
  AND U35620 ( .A(n34723), .B(n34722), .Z(n34771) );
  XOR U35621 ( .A(n34772), .B(n34771), .Z(n34773) );
  NANDN U35622 ( .A(n34725), .B(n34724), .Z(n34729) );
  NANDN U35623 ( .A(n34727), .B(n34726), .Z(n34728) );
  NAND U35624 ( .A(n34729), .B(n34728), .Z(n34774) );
  XOR U35625 ( .A(n34773), .B(n34774), .Z(n34741) );
  OR U35626 ( .A(n34731), .B(n34730), .Z(n34735) );
  NANDN U35627 ( .A(n34733), .B(n34732), .Z(n34734) );
  NAND U35628 ( .A(n34735), .B(n34734), .Z(n34742) );
  XNOR U35629 ( .A(n34741), .B(n34742), .Z(n34743) );
  XNOR U35630 ( .A(n34744), .B(n34743), .Z(n34777) );
  XNOR U35631 ( .A(n34777), .B(sreg[1861]), .Z(n34779) );
  NAND U35632 ( .A(n34736), .B(sreg[1860]), .Z(n34740) );
  OR U35633 ( .A(n34738), .B(n34737), .Z(n34739) );
  AND U35634 ( .A(n34740), .B(n34739), .Z(n34778) );
  XOR U35635 ( .A(n34779), .B(n34778), .Z(c[1861]) );
  NANDN U35636 ( .A(n34742), .B(n34741), .Z(n34746) );
  NAND U35637 ( .A(n34744), .B(n34743), .Z(n34745) );
  NAND U35638 ( .A(n34746), .B(n34745), .Z(n34785) );
  NAND U35639 ( .A(b[0]), .B(a[846]), .Z(n34747) );
  XNOR U35640 ( .A(b[1]), .B(n34747), .Z(n34749) );
  NAND U35641 ( .A(n135), .B(a[845]), .Z(n34748) );
  AND U35642 ( .A(n34749), .B(n34748), .Z(n34802) );
  XOR U35643 ( .A(a[842]), .B(n42197), .Z(n34791) );
  NANDN U35644 ( .A(n34791), .B(n42173), .Z(n34752) );
  NANDN U35645 ( .A(n34750), .B(n42172), .Z(n34751) );
  NAND U35646 ( .A(n34752), .B(n34751), .Z(n34800) );
  NAND U35647 ( .A(b[7]), .B(a[838]), .Z(n34801) );
  XNOR U35648 ( .A(n34800), .B(n34801), .Z(n34803) );
  XOR U35649 ( .A(n34802), .B(n34803), .Z(n34809) );
  NANDN U35650 ( .A(n34753), .B(n42093), .Z(n34755) );
  XOR U35651 ( .A(n42134), .B(a[844]), .Z(n34794) );
  NANDN U35652 ( .A(n34794), .B(n42095), .Z(n34754) );
  NAND U35653 ( .A(n34755), .B(n34754), .Z(n34807) );
  NANDN U35654 ( .A(n34756), .B(n42231), .Z(n34758) );
  XOR U35655 ( .A(n232), .B(a[840]), .Z(n34797) );
  NANDN U35656 ( .A(n34797), .B(n42234), .Z(n34757) );
  AND U35657 ( .A(n34758), .B(n34757), .Z(n34806) );
  XNOR U35658 ( .A(n34807), .B(n34806), .Z(n34808) );
  XNOR U35659 ( .A(n34809), .B(n34808), .Z(n34813) );
  NANDN U35660 ( .A(n34760), .B(n34759), .Z(n34764) );
  NAND U35661 ( .A(n34762), .B(n34761), .Z(n34763) );
  AND U35662 ( .A(n34764), .B(n34763), .Z(n34812) );
  XOR U35663 ( .A(n34813), .B(n34812), .Z(n34814) );
  NANDN U35664 ( .A(n34766), .B(n34765), .Z(n34770) );
  NANDN U35665 ( .A(n34768), .B(n34767), .Z(n34769) );
  NAND U35666 ( .A(n34770), .B(n34769), .Z(n34815) );
  XOR U35667 ( .A(n34814), .B(n34815), .Z(n34782) );
  OR U35668 ( .A(n34772), .B(n34771), .Z(n34776) );
  NANDN U35669 ( .A(n34774), .B(n34773), .Z(n34775) );
  NAND U35670 ( .A(n34776), .B(n34775), .Z(n34783) );
  XNOR U35671 ( .A(n34782), .B(n34783), .Z(n34784) );
  XNOR U35672 ( .A(n34785), .B(n34784), .Z(n34818) );
  XNOR U35673 ( .A(n34818), .B(sreg[1862]), .Z(n34820) );
  NAND U35674 ( .A(n34777), .B(sreg[1861]), .Z(n34781) );
  OR U35675 ( .A(n34779), .B(n34778), .Z(n34780) );
  AND U35676 ( .A(n34781), .B(n34780), .Z(n34819) );
  XOR U35677 ( .A(n34820), .B(n34819), .Z(c[1862]) );
  NANDN U35678 ( .A(n34783), .B(n34782), .Z(n34787) );
  NAND U35679 ( .A(n34785), .B(n34784), .Z(n34786) );
  NAND U35680 ( .A(n34787), .B(n34786), .Z(n34826) );
  NAND U35681 ( .A(b[0]), .B(a[847]), .Z(n34788) );
  XNOR U35682 ( .A(b[1]), .B(n34788), .Z(n34790) );
  NAND U35683 ( .A(n136), .B(a[846]), .Z(n34789) );
  AND U35684 ( .A(n34790), .B(n34789), .Z(n34843) );
  XOR U35685 ( .A(a[843]), .B(n42197), .Z(n34832) );
  NANDN U35686 ( .A(n34832), .B(n42173), .Z(n34793) );
  NANDN U35687 ( .A(n34791), .B(n42172), .Z(n34792) );
  NAND U35688 ( .A(n34793), .B(n34792), .Z(n34841) );
  NAND U35689 ( .A(b[7]), .B(a[839]), .Z(n34842) );
  XNOR U35690 ( .A(n34841), .B(n34842), .Z(n34844) );
  XOR U35691 ( .A(n34843), .B(n34844), .Z(n34850) );
  NANDN U35692 ( .A(n34794), .B(n42093), .Z(n34796) );
  XOR U35693 ( .A(n42134), .B(a[845]), .Z(n34835) );
  NANDN U35694 ( .A(n34835), .B(n42095), .Z(n34795) );
  NAND U35695 ( .A(n34796), .B(n34795), .Z(n34848) );
  NANDN U35696 ( .A(n34797), .B(n42231), .Z(n34799) );
  XOR U35697 ( .A(n232), .B(a[841]), .Z(n34838) );
  NANDN U35698 ( .A(n34838), .B(n42234), .Z(n34798) );
  AND U35699 ( .A(n34799), .B(n34798), .Z(n34847) );
  XNOR U35700 ( .A(n34848), .B(n34847), .Z(n34849) );
  XNOR U35701 ( .A(n34850), .B(n34849), .Z(n34854) );
  NANDN U35702 ( .A(n34801), .B(n34800), .Z(n34805) );
  NAND U35703 ( .A(n34803), .B(n34802), .Z(n34804) );
  AND U35704 ( .A(n34805), .B(n34804), .Z(n34853) );
  XOR U35705 ( .A(n34854), .B(n34853), .Z(n34855) );
  NANDN U35706 ( .A(n34807), .B(n34806), .Z(n34811) );
  NANDN U35707 ( .A(n34809), .B(n34808), .Z(n34810) );
  NAND U35708 ( .A(n34811), .B(n34810), .Z(n34856) );
  XOR U35709 ( .A(n34855), .B(n34856), .Z(n34823) );
  OR U35710 ( .A(n34813), .B(n34812), .Z(n34817) );
  NANDN U35711 ( .A(n34815), .B(n34814), .Z(n34816) );
  NAND U35712 ( .A(n34817), .B(n34816), .Z(n34824) );
  XNOR U35713 ( .A(n34823), .B(n34824), .Z(n34825) );
  XNOR U35714 ( .A(n34826), .B(n34825), .Z(n34859) );
  XNOR U35715 ( .A(n34859), .B(sreg[1863]), .Z(n34861) );
  NAND U35716 ( .A(n34818), .B(sreg[1862]), .Z(n34822) );
  OR U35717 ( .A(n34820), .B(n34819), .Z(n34821) );
  AND U35718 ( .A(n34822), .B(n34821), .Z(n34860) );
  XOR U35719 ( .A(n34861), .B(n34860), .Z(c[1863]) );
  NANDN U35720 ( .A(n34824), .B(n34823), .Z(n34828) );
  NAND U35721 ( .A(n34826), .B(n34825), .Z(n34827) );
  NAND U35722 ( .A(n34828), .B(n34827), .Z(n34867) );
  NAND U35723 ( .A(b[0]), .B(a[848]), .Z(n34829) );
  XNOR U35724 ( .A(b[1]), .B(n34829), .Z(n34831) );
  NAND U35725 ( .A(n136), .B(a[847]), .Z(n34830) );
  AND U35726 ( .A(n34831), .B(n34830), .Z(n34884) );
  XOR U35727 ( .A(a[844]), .B(n42197), .Z(n34873) );
  NANDN U35728 ( .A(n34873), .B(n42173), .Z(n34834) );
  NANDN U35729 ( .A(n34832), .B(n42172), .Z(n34833) );
  NAND U35730 ( .A(n34834), .B(n34833), .Z(n34882) );
  NAND U35731 ( .A(b[7]), .B(a[840]), .Z(n34883) );
  XNOR U35732 ( .A(n34882), .B(n34883), .Z(n34885) );
  XOR U35733 ( .A(n34884), .B(n34885), .Z(n34891) );
  NANDN U35734 ( .A(n34835), .B(n42093), .Z(n34837) );
  XOR U35735 ( .A(n42134), .B(a[846]), .Z(n34876) );
  NANDN U35736 ( .A(n34876), .B(n42095), .Z(n34836) );
  NAND U35737 ( .A(n34837), .B(n34836), .Z(n34889) );
  NANDN U35738 ( .A(n34838), .B(n42231), .Z(n34840) );
  XOR U35739 ( .A(n232), .B(a[842]), .Z(n34879) );
  NANDN U35740 ( .A(n34879), .B(n42234), .Z(n34839) );
  AND U35741 ( .A(n34840), .B(n34839), .Z(n34888) );
  XNOR U35742 ( .A(n34889), .B(n34888), .Z(n34890) );
  XNOR U35743 ( .A(n34891), .B(n34890), .Z(n34895) );
  NANDN U35744 ( .A(n34842), .B(n34841), .Z(n34846) );
  NAND U35745 ( .A(n34844), .B(n34843), .Z(n34845) );
  AND U35746 ( .A(n34846), .B(n34845), .Z(n34894) );
  XOR U35747 ( .A(n34895), .B(n34894), .Z(n34896) );
  NANDN U35748 ( .A(n34848), .B(n34847), .Z(n34852) );
  NANDN U35749 ( .A(n34850), .B(n34849), .Z(n34851) );
  NAND U35750 ( .A(n34852), .B(n34851), .Z(n34897) );
  XOR U35751 ( .A(n34896), .B(n34897), .Z(n34864) );
  OR U35752 ( .A(n34854), .B(n34853), .Z(n34858) );
  NANDN U35753 ( .A(n34856), .B(n34855), .Z(n34857) );
  NAND U35754 ( .A(n34858), .B(n34857), .Z(n34865) );
  XNOR U35755 ( .A(n34864), .B(n34865), .Z(n34866) );
  XNOR U35756 ( .A(n34867), .B(n34866), .Z(n34900) );
  XNOR U35757 ( .A(n34900), .B(sreg[1864]), .Z(n34902) );
  NAND U35758 ( .A(n34859), .B(sreg[1863]), .Z(n34863) );
  OR U35759 ( .A(n34861), .B(n34860), .Z(n34862) );
  AND U35760 ( .A(n34863), .B(n34862), .Z(n34901) );
  XOR U35761 ( .A(n34902), .B(n34901), .Z(c[1864]) );
  NANDN U35762 ( .A(n34865), .B(n34864), .Z(n34869) );
  NAND U35763 ( .A(n34867), .B(n34866), .Z(n34868) );
  NAND U35764 ( .A(n34869), .B(n34868), .Z(n34908) );
  NAND U35765 ( .A(b[0]), .B(a[849]), .Z(n34870) );
  XNOR U35766 ( .A(b[1]), .B(n34870), .Z(n34872) );
  NAND U35767 ( .A(n136), .B(a[848]), .Z(n34871) );
  AND U35768 ( .A(n34872), .B(n34871), .Z(n34925) );
  XOR U35769 ( .A(a[845]), .B(n42197), .Z(n34914) );
  NANDN U35770 ( .A(n34914), .B(n42173), .Z(n34875) );
  NANDN U35771 ( .A(n34873), .B(n42172), .Z(n34874) );
  NAND U35772 ( .A(n34875), .B(n34874), .Z(n34923) );
  NAND U35773 ( .A(b[7]), .B(a[841]), .Z(n34924) );
  XNOR U35774 ( .A(n34923), .B(n34924), .Z(n34926) );
  XOR U35775 ( .A(n34925), .B(n34926), .Z(n34932) );
  NANDN U35776 ( .A(n34876), .B(n42093), .Z(n34878) );
  XOR U35777 ( .A(n42134), .B(a[847]), .Z(n34917) );
  NANDN U35778 ( .A(n34917), .B(n42095), .Z(n34877) );
  NAND U35779 ( .A(n34878), .B(n34877), .Z(n34930) );
  NANDN U35780 ( .A(n34879), .B(n42231), .Z(n34881) );
  XOR U35781 ( .A(n232), .B(a[843]), .Z(n34920) );
  NANDN U35782 ( .A(n34920), .B(n42234), .Z(n34880) );
  AND U35783 ( .A(n34881), .B(n34880), .Z(n34929) );
  XNOR U35784 ( .A(n34930), .B(n34929), .Z(n34931) );
  XNOR U35785 ( .A(n34932), .B(n34931), .Z(n34936) );
  NANDN U35786 ( .A(n34883), .B(n34882), .Z(n34887) );
  NAND U35787 ( .A(n34885), .B(n34884), .Z(n34886) );
  AND U35788 ( .A(n34887), .B(n34886), .Z(n34935) );
  XOR U35789 ( .A(n34936), .B(n34935), .Z(n34937) );
  NANDN U35790 ( .A(n34889), .B(n34888), .Z(n34893) );
  NANDN U35791 ( .A(n34891), .B(n34890), .Z(n34892) );
  NAND U35792 ( .A(n34893), .B(n34892), .Z(n34938) );
  XOR U35793 ( .A(n34937), .B(n34938), .Z(n34905) );
  OR U35794 ( .A(n34895), .B(n34894), .Z(n34899) );
  NANDN U35795 ( .A(n34897), .B(n34896), .Z(n34898) );
  NAND U35796 ( .A(n34899), .B(n34898), .Z(n34906) );
  XNOR U35797 ( .A(n34905), .B(n34906), .Z(n34907) );
  XNOR U35798 ( .A(n34908), .B(n34907), .Z(n34941) );
  XNOR U35799 ( .A(n34941), .B(sreg[1865]), .Z(n34943) );
  NAND U35800 ( .A(n34900), .B(sreg[1864]), .Z(n34904) );
  OR U35801 ( .A(n34902), .B(n34901), .Z(n34903) );
  AND U35802 ( .A(n34904), .B(n34903), .Z(n34942) );
  XOR U35803 ( .A(n34943), .B(n34942), .Z(c[1865]) );
  NANDN U35804 ( .A(n34906), .B(n34905), .Z(n34910) );
  NAND U35805 ( .A(n34908), .B(n34907), .Z(n34909) );
  NAND U35806 ( .A(n34910), .B(n34909), .Z(n34949) );
  NAND U35807 ( .A(b[0]), .B(a[850]), .Z(n34911) );
  XNOR U35808 ( .A(b[1]), .B(n34911), .Z(n34913) );
  NAND U35809 ( .A(n136), .B(a[849]), .Z(n34912) );
  AND U35810 ( .A(n34913), .B(n34912), .Z(n34966) );
  XOR U35811 ( .A(a[846]), .B(n42197), .Z(n34955) );
  NANDN U35812 ( .A(n34955), .B(n42173), .Z(n34916) );
  NANDN U35813 ( .A(n34914), .B(n42172), .Z(n34915) );
  NAND U35814 ( .A(n34916), .B(n34915), .Z(n34964) );
  NAND U35815 ( .A(b[7]), .B(a[842]), .Z(n34965) );
  XNOR U35816 ( .A(n34964), .B(n34965), .Z(n34967) );
  XOR U35817 ( .A(n34966), .B(n34967), .Z(n34973) );
  NANDN U35818 ( .A(n34917), .B(n42093), .Z(n34919) );
  XOR U35819 ( .A(n42134), .B(a[848]), .Z(n34958) );
  NANDN U35820 ( .A(n34958), .B(n42095), .Z(n34918) );
  NAND U35821 ( .A(n34919), .B(n34918), .Z(n34971) );
  NANDN U35822 ( .A(n34920), .B(n42231), .Z(n34922) );
  XOR U35823 ( .A(n232), .B(a[844]), .Z(n34961) );
  NANDN U35824 ( .A(n34961), .B(n42234), .Z(n34921) );
  AND U35825 ( .A(n34922), .B(n34921), .Z(n34970) );
  XNOR U35826 ( .A(n34971), .B(n34970), .Z(n34972) );
  XNOR U35827 ( .A(n34973), .B(n34972), .Z(n34977) );
  NANDN U35828 ( .A(n34924), .B(n34923), .Z(n34928) );
  NAND U35829 ( .A(n34926), .B(n34925), .Z(n34927) );
  AND U35830 ( .A(n34928), .B(n34927), .Z(n34976) );
  XOR U35831 ( .A(n34977), .B(n34976), .Z(n34978) );
  NANDN U35832 ( .A(n34930), .B(n34929), .Z(n34934) );
  NANDN U35833 ( .A(n34932), .B(n34931), .Z(n34933) );
  NAND U35834 ( .A(n34934), .B(n34933), .Z(n34979) );
  XOR U35835 ( .A(n34978), .B(n34979), .Z(n34946) );
  OR U35836 ( .A(n34936), .B(n34935), .Z(n34940) );
  NANDN U35837 ( .A(n34938), .B(n34937), .Z(n34939) );
  NAND U35838 ( .A(n34940), .B(n34939), .Z(n34947) );
  XNOR U35839 ( .A(n34946), .B(n34947), .Z(n34948) );
  XNOR U35840 ( .A(n34949), .B(n34948), .Z(n34982) );
  XNOR U35841 ( .A(n34982), .B(sreg[1866]), .Z(n34984) );
  NAND U35842 ( .A(n34941), .B(sreg[1865]), .Z(n34945) );
  OR U35843 ( .A(n34943), .B(n34942), .Z(n34944) );
  AND U35844 ( .A(n34945), .B(n34944), .Z(n34983) );
  XOR U35845 ( .A(n34984), .B(n34983), .Z(c[1866]) );
  NANDN U35846 ( .A(n34947), .B(n34946), .Z(n34951) );
  NAND U35847 ( .A(n34949), .B(n34948), .Z(n34950) );
  NAND U35848 ( .A(n34951), .B(n34950), .Z(n34990) );
  NAND U35849 ( .A(b[0]), .B(a[851]), .Z(n34952) );
  XNOR U35850 ( .A(b[1]), .B(n34952), .Z(n34954) );
  NAND U35851 ( .A(n136), .B(a[850]), .Z(n34953) );
  AND U35852 ( .A(n34954), .B(n34953), .Z(n35007) );
  XOR U35853 ( .A(a[847]), .B(n42197), .Z(n34996) );
  NANDN U35854 ( .A(n34996), .B(n42173), .Z(n34957) );
  NANDN U35855 ( .A(n34955), .B(n42172), .Z(n34956) );
  NAND U35856 ( .A(n34957), .B(n34956), .Z(n35005) );
  NAND U35857 ( .A(b[7]), .B(a[843]), .Z(n35006) );
  XNOR U35858 ( .A(n35005), .B(n35006), .Z(n35008) );
  XOR U35859 ( .A(n35007), .B(n35008), .Z(n35014) );
  NANDN U35860 ( .A(n34958), .B(n42093), .Z(n34960) );
  XOR U35861 ( .A(n42134), .B(a[849]), .Z(n34999) );
  NANDN U35862 ( .A(n34999), .B(n42095), .Z(n34959) );
  NAND U35863 ( .A(n34960), .B(n34959), .Z(n35012) );
  NANDN U35864 ( .A(n34961), .B(n42231), .Z(n34963) );
  XOR U35865 ( .A(n232), .B(a[845]), .Z(n35002) );
  NANDN U35866 ( .A(n35002), .B(n42234), .Z(n34962) );
  AND U35867 ( .A(n34963), .B(n34962), .Z(n35011) );
  XNOR U35868 ( .A(n35012), .B(n35011), .Z(n35013) );
  XNOR U35869 ( .A(n35014), .B(n35013), .Z(n35018) );
  NANDN U35870 ( .A(n34965), .B(n34964), .Z(n34969) );
  NAND U35871 ( .A(n34967), .B(n34966), .Z(n34968) );
  AND U35872 ( .A(n34969), .B(n34968), .Z(n35017) );
  XOR U35873 ( .A(n35018), .B(n35017), .Z(n35019) );
  NANDN U35874 ( .A(n34971), .B(n34970), .Z(n34975) );
  NANDN U35875 ( .A(n34973), .B(n34972), .Z(n34974) );
  NAND U35876 ( .A(n34975), .B(n34974), .Z(n35020) );
  XOR U35877 ( .A(n35019), .B(n35020), .Z(n34987) );
  OR U35878 ( .A(n34977), .B(n34976), .Z(n34981) );
  NANDN U35879 ( .A(n34979), .B(n34978), .Z(n34980) );
  NAND U35880 ( .A(n34981), .B(n34980), .Z(n34988) );
  XNOR U35881 ( .A(n34987), .B(n34988), .Z(n34989) );
  XNOR U35882 ( .A(n34990), .B(n34989), .Z(n35023) );
  XNOR U35883 ( .A(n35023), .B(sreg[1867]), .Z(n35025) );
  NAND U35884 ( .A(n34982), .B(sreg[1866]), .Z(n34986) );
  OR U35885 ( .A(n34984), .B(n34983), .Z(n34985) );
  AND U35886 ( .A(n34986), .B(n34985), .Z(n35024) );
  XOR U35887 ( .A(n35025), .B(n35024), .Z(c[1867]) );
  NANDN U35888 ( .A(n34988), .B(n34987), .Z(n34992) );
  NAND U35889 ( .A(n34990), .B(n34989), .Z(n34991) );
  NAND U35890 ( .A(n34992), .B(n34991), .Z(n35031) );
  NAND U35891 ( .A(b[0]), .B(a[852]), .Z(n34993) );
  XNOR U35892 ( .A(b[1]), .B(n34993), .Z(n34995) );
  NAND U35893 ( .A(n136), .B(a[851]), .Z(n34994) );
  AND U35894 ( .A(n34995), .B(n34994), .Z(n35048) );
  XOR U35895 ( .A(a[848]), .B(n42197), .Z(n35037) );
  NANDN U35896 ( .A(n35037), .B(n42173), .Z(n34998) );
  NANDN U35897 ( .A(n34996), .B(n42172), .Z(n34997) );
  NAND U35898 ( .A(n34998), .B(n34997), .Z(n35046) );
  NAND U35899 ( .A(b[7]), .B(a[844]), .Z(n35047) );
  XNOR U35900 ( .A(n35046), .B(n35047), .Z(n35049) );
  XOR U35901 ( .A(n35048), .B(n35049), .Z(n35055) );
  NANDN U35902 ( .A(n34999), .B(n42093), .Z(n35001) );
  XOR U35903 ( .A(n42134), .B(a[850]), .Z(n35040) );
  NANDN U35904 ( .A(n35040), .B(n42095), .Z(n35000) );
  NAND U35905 ( .A(n35001), .B(n35000), .Z(n35053) );
  NANDN U35906 ( .A(n35002), .B(n42231), .Z(n35004) );
  XOR U35907 ( .A(n232), .B(a[846]), .Z(n35043) );
  NANDN U35908 ( .A(n35043), .B(n42234), .Z(n35003) );
  AND U35909 ( .A(n35004), .B(n35003), .Z(n35052) );
  XNOR U35910 ( .A(n35053), .B(n35052), .Z(n35054) );
  XNOR U35911 ( .A(n35055), .B(n35054), .Z(n35059) );
  NANDN U35912 ( .A(n35006), .B(n35005), .Z(n35010) );
  NAND U35913 ( .A(n35008), .B(n35007), .Z(n35009) );
  AND U35914 ( .A(n35010), .B(n35009), .Z(n35058) );
  XOR U35915 ( .A(n35059), .B(n35058), .Z(n35060) );
  NANDN U35916 ( .A(n35012), .B(n35011), .Z(n35016) );
  NANDN U35917 ( .A(n35014), .B(n35013), .Z(n35015) );
  NAND U35918 ( .A(n35016), .B(n35015), .Z(n35061) );
  XOR U35919 ( .A(n35060), .B(n35061), .Z(n35028) );
  OR U35920 ( .A(n35018), .B(n35017), .Z(n35022) );
  NANDN U35921 ( .A(n35020), .B(n35019), .Z(n35021) );
  NAND U35922 ( .A(n35022), .B(n35021), .Z(n35029) );
  XNOR U35923 ( .A(n35028), .B(n35029), .Z(n35030) );
  XNOR U35924 ( .A(n35031), .B(n35030), .Z(n35064) );
  XNOR U35925 ( .A(n35064), .B(sreg[1868]), .Z(n35066) );
  NAND U35926 ( .A(n35023), .B(sreg[1867]), .Z(n35027) );
  OR U35927 ( .A(n35025), .B(n35024), .Z(n35026) );
  AND U35928 ( .A(n35027), .B(n35026), .Z(n35065) );
  XOR U35929 ( .A(n35066), .B(n35065), .Z(c[1868]) );
  NANDN U35930 ( .A(n35029), .B(n35028), .Z(n35033) );
  NAND U35931 ( .A(n35031), .B(n35030), .Z(n35032) );
  NAND U35932 ( .A(n35033), .B(n35032), .Z(n35072) );
  NAND U35933 ( .A(b[0]), .B(a[853]), .Z(n35034) );
  XNOR U35934 ( .A(b[1]), .B(n35034), .Z(n35036) );
  NAND U35935 ( .A(n136), .B(a[852]), .Z(n35035) );
  AND U35936 ( .A(n35036), .B(n35035), .Z(n35089) );
  XOR U35937 ( .A(a[849]), .B(n42197), .Z(n35078) );
  NANDN U35938 ( .A(n35078), .B(n42173), .Z(n35039) );
  NANDN U35939 ( .A(n35037), .B(n42172), .Z(n35038) );
  NAND U35940 ( .A(n35039), .B(n35038), .Z(n35087) );
  NAND U35941 ( .A(b[7]), .B(a[845]), .Z(n35088) );
  XNOR U35942 ( .A(n35087), .B(n35088), .Z(n35090) );
  XOR U35943 ( .A(n35089), .B(n35090), .Z(n35096) );
  NANDN U35944 ( .A(n35040), .B(n42093), .Z(n35042) );
  XOR U35945 ( .A(n42134), .B(a[851]), .Z(n35081) );
  NANDN U35946 ( .A(n35081), .B(n42095), .Z(n35041) );
  NAND U35947 ( .A(n35042), .B(n35041), .Z(n35094) );
  NANDN U35948 ( .A(n35043), .B(n42231), .Z(n35045) );
  XOR U35949 ( .A(n232), .B(a[847]), .Z(n35084) );
  NANDN U35950 ( .A(n35084), .B(n42234), .Z(n35044) );
  AND U35951 ( .A(n35045), .B(n35044), .Z(n35093) );
  XNOR U35952 ( .A(n35094), .B(n35093), .Z(n35095) );
  XNOR U35953 ( .A(n35096), .B(n35095), .Z(n35100) );
  NANDN U35954 ( .A(n35047), .B(n35046), .Z(n35051) );
  NAND U35955 ( .A(n35049), .B(n35048), .Z(n35050) );
  AND U35956 ( .A(n35051), .B(n35050), .Z(n35099) );
  XOR U35957 ( .A(n35100), .B(n35099), .Z(n35101) );
  NANDN U35958 ( .A(n35053), .B(n35052), .Z(n35057) );
  NANDN U35959 ( .A(n35055), .B(n35054), .Z(n35056) );
  NAND U35960 ( .A(n35057), .B(n35056), .Z(n35102) );
  XOR U35961 ( .A(n35101), .B(n35102), .Z(n35069) );
  OR U35962 ( .A(n35059), .B(n35058), .Z(n35063) );
  NANDN U35963 ( .A(n35061), .B(n35060), .Z(n35062) );
  NAND U35964 ( .A(n35063), .B(n35062), .Z(n35070) );
  XNOR U35965 ( .A(n35069), .B(n35070), .Z(n35071) );
  XNOR U35966 ( .A(n35072), .B(n35071), .Z(n35105) );
  XNOR U35967 ( .A(n35105), .B(sreg[1869]), .Z(n35107) );
  NAND U35968 ( .A(n35064), .B(sreg[1868]), .Z(n35068) );
  OR U35969 ( .A(n35066), .B(n35065), .Z(n35067) );
  AND U35970 ( .A(n35068), .B(n35067), .Z(n35106) );
  XOR U35971 ( .A(n35107), .B(n35106), .Z(c[1869]) );
  NANDN U35972 ( .A(n35070), .B(n35069), .Z(n35074) );
  NAND U35973 ( .A(n35072), .B(n35071), .Z(n35073) );
  NAND U35974 ( .A(n35074), .B(n35073), .Z(n35113) );
  NAND U35975 ( .A(b[0]), .B(a[854]), .Z(n35075) );
  XNOR U35976 ( .A(b[1]), .B(n35075), .Z(n35077) );
  NAND U35977 ( .A(n137), .B(a[853]), .Z(n35076) );
  AND U35978 ( .A(n35077), .B(n35076), .Z(n35130) );
  XOR U35979 ( .A(a[850]), .B(n42197), .Z(n35119) );
  NANDN U35980 ( .A(n35119), .B(n42173), .Z(n35080) );
  NANDN U35981 ( .A(n35078), .B(n42172), .Z(n35079) );
  NAND U35982 ( .A(n35080), .B(n35079), .Z(n35128) );
  NAND U35983 ( .A(b[7]), .B(a[846]), .Z(n35129) );
  XNOR U35984 ( .A(n35128), .B(n35129), .Z(n35131) );
  XOR U35985 ( .A(n35130), .B(n35131), .Z(n35137) );
  NANDN U35986 ( .A(n35081), .B(n42093), .Z(n35083) );
  XOR U35987 ( .A(n42134), .B(a[852]), .Z(n35122) );
  NANDN U35988 ( .A(n35122), .B(n42095), .Z(n35082) );
  NAND U35989 ( .A(n35083), .B(n35082), .Z(n35135) );
  NANDN U35990 ( .A(n35084), .B(n42231), .Z(n35086) );
  XOR U35991 ( .A(n232), .B(a[848]), .Z(n35125) );
  NANDN U35992 ( .A(n35125), .B(n42234), .Z(n35085) );
  AND U35993 ( .A(n35086), .B(n35085), .Z(n35134) );
  XNOR U35994 ( .A(n35135), .B(n35134), .Z(n35136) );
  XNOR U35995 ( .A(n35137), .B(n35136), .Z(n35141) );
  NANDN U35996 ( .A(n35088), .B(n35087), .Z(n35092) );
  NAND U35997 ( .A(n35090), .B(n35089), .Z(n35091) );
  AND U35998 ( .A(n35092), .B(n35091), .Z(n35140) );
  XOR U35999 ( .A(n35141), .B(n35140), .Z(n35142) );
  NANDN U36000 ( .A(n35094), .B(n35093), .Z(n35098) );
  NANDN U36001 ( .A(n35096), .B(n35095), .Z(n35097) );
  NAND U36002 ( .A(n35098), .B(n35097), .Z(n35143) );
  XOR U36003 ( .A(n35142), .B(n35143), .Z(n35110) );
  OR U36004 ( .A(n35100), .B(n35099), .Z(n35104) );
  NANDN U36005 ( .A(n35102), .B(n35101), .Z(n35103) );
  NAND U36006 ( .A(n35104), .B(n35103), .Z(n35111) );
  XNOR U36007 ( .A(n35110), .B(n35111), .Z(n35112) );
  XNOR U36008 ( .A(n35113), .B(n35112), .Z(n35146) );
  XNOR U36009 ( .A(n35146), .B(sreg[1870]), .Z(n35148) );
  NAND U36010 ( .A(n35105), .B(sreg[1869]), .Z(n35109) );
  OR U36011 ( .A(n35107), .B(n35106), .Z(n35108) );
  AND U36012 ( .A(n35109), .B(n35108), .Z(n35147) );
  XOR U36013 ( .A(n35148), .B(n35147), .Z(c[1870]) );
  NANDN U36014 ( .A(n35111), .B(n35110), .Z(n35115) );
  NAND U36015 ( .A(n35113), .B(n35112), .Z(n35114) );
  NAND U36016 ( .A(n35115), .B(n35114), .Z(n35154) );
  NAND U36017 ( .A(b[0]), .B(a[855]), .Z(n35116) );
  XNOR U36018 ( .A(b[1]), .B(n35116), .Z(n35118) );
  NAND U36019 ( .A(n137), .B(a[854]), .Z(n35117) );
  AND U36020 ( .A(n35118), .B(n35117), .Z(n35171) );
  XOR U36021 ( .A(a[851]), .B(n42197), .Z(n35160) );
  NANDN U36022 ( .A(n35160), .B(n42173), .Z(n35121) );
  NANDN U36023 ( .A(n35119), .B(n42172), .Z(n35120) );
  NAND U36024 ( .A(n35121), .B(n35120), .Z(n35169) );
  NAND U36025 ( .A(b[7]), .B(a[847]), .Z(n35170) );
  XNOR U36026 ( .A(n35169), .B(n35170), .Z(n35172) );
  XOR U36027 ( .A(n35171), .B(n35172), .Z(n35178) );
  NANDN U36028 ( .A(n35122), .B(n42093), .Z(n35124) );
  XOR U36029 ( .A(n42134), .B(a[853]), .Z(n35163) );
  NANDN U36030 ( .A(n35163), .B(n42095), .Z(n35123) );
  NAND U36031 ( .A(n35124), .B(n35123), .Z(n35176) );
  NANDN U36032 ( .A(n35125), .B(n42231), .Z(n35127) );
  XOR U36033 ( .A(n232), .B(a[849]), .Z(n35166) );
  NANDN U36034 ( .A(n35166), .B(n42234), .Z(n35126) );
  AND U36035 ( .A(n35127), .B(n35126), .Z(n35175) );
  XNOR U36036 ( .A(n35176), .B(n35175), .Z(n35177) );
  XNOR U36037 ( .A(n35178), .B(n35177), .Z(n35182) );
  NANDN U36038 ( .A(n35129), .B(n35128), .Z(n35133) );
  NAND U36039 ( .A(n35131), .B(n35130), .Z(n35132) );
  AND U36040 ( .A(n35133), .B(n35132), .Z(n35181) );
  XOR U36041 ( .A(n35182), .B(n35181), .Z(n35183) );
  NANDN U36042 ( .A(n35135), .B(n35134), .Z(n35139) );
  NANDN U36043 ( .A(n35137), .B(n35136), .Z(n35138) );
  NAND U36044 ( .A(n35139), .B(n35138), .Z(n35184) );
  XOR U36045 ( .A(n35183), .B(n35184), .Z(n35151) );
  OR U36046 ( .A(n35141), .B(n35140), .Z(n35145) );
  NANDN U36047 ( .A(n35143), .B(n35142), .Z(n35144) );
  NAND U36048 ( .A(n35145), .B(n35144), .Z(n35152) );
  XNOR U36049 ( .A(n35151), .B(n35152), .Z(n35153) );
  XNOR U36050 ( .A(n35154), .B(n35153), .Z(n35187) );
  XNOR U36051 ( .A(n35187), .B(sreg[1871]), .Z(n35189) );
  NAND U36052 ( .A(n35146), .B(sreg[1870]), .Z(n35150) );
  OR U36053 ( .A(n35148), .B(n35147), .Z(n35149) );
  AND U36054 ( .A(n35150), .B(n35149), .Z(n35188) );
  XOR U36055 ( .A(n35189), .B(n35188), .Z(c[1871]) );
  NANDN U36056 ( .A(n35152), .B(n35151), .Z(n35156) );
  NAND U36057 ( .A(n35154), .B(n35153), .Z(n35155) );
  NAND U36058 ( .A(n35156), .B(n35155), .Z(n35195) );
  NAND U36059 ( .A(b[0]), .B(a[856]), .Z(n35157) );
  XNOR U36060 ( .A(b[1]), .B(n35157), .Z(n35159) );
  NAND U36061 ( .A(n137), .B(a[855]), .Z(n35158) );
  AND U36062 ( .A(n35159), .B(n35158), .Z(n35212) );
  XOR U36063 ( .A(a[852]), .B(n42197), .Z(n35201) );
  NANDN U36064 ( .A(n35201), .B(n42173), .Z(n35162) );
  NANDN U36065 ( .A(n35160), .B(n42172), .Z(n35161) );
  NAND U36066 ( .A(n35162), .B(n35161), .Z(n35210) );
  NAND U36067 ( .A(b[7]), .B(a[848]), .Z(n35211) );
  XNOR U36068 ( .A(n35210), .B(n35211), .Z(n35213) );
  XOR U36069 ( .A(n35212), .B(n35213), .Z(n35219) );
  NANDN U36070 ( .A(n35163), .B(n42093), .Z(n35165) );
  XOR U36071 ( .A(n42134), .B(a[854]), .Z(n35204) );
  NANDN U36072 ( .A(n35204), .B(n42095), .Z(n35164) );
  NAND U36073 ( .A(n35165), .B(n35164), .Z(n35217) );
  NANDN U36074 ( .A(n35166), .B(n42231), .Z(n35168) );
  XOR U36075 ( .A(n232), .B(a[850]), .Z(n35207) );
  NANDN U36076 ( .A(n35207), .B(n42234), .Z(n35167) );
  AND U36077 ( .A(n35168), .B(n35167), .Z(n35216) );
  XNOR U36078 ( .A(n35217), .B(n35216), .Z(n35218) );
  XNOR U36079 ( .A(n35219), .B(n35218), .Z(n35223) );
  NANDN U36080 ( .A(n35170), .B(n35169), .Z(n35174) );
  NAND U36081 ( .A(n35172), .B(n35171), .Z(n35173) );
  AND U36082 ( .A(n35174), .B(n35173), .Z(n35222) );
  XOR U36083 ( .A(n35223), .B(n35222), .Z(n35224) );
  NANDN U36084 ( .A(n35176), .B(n35175), .Z(n35180) );
  NANDN U36085 ( .A(n35178), .B(n35177), .Z(n35179) );
  NAND U36086 ( .A(n35180), .B(n35179), .Z(n35225) );
  XOR U36087 ( .A(n35224), .B(n35225), .Z(n35192) );
  OR U36088 ( .A(n35182), .B(n35181), .Z(n35186) );
  NANDN U36089 ( .A(n35184), .B(n35183), .Z(n35185) );
  NAND U36090 ( .A(n35186), .B(n35185), .Z(n35193) );
  XNOR U36091 ( .A(n35192), .B(n35193), .Z(n35194) );
  XNOR U36092 ( .A(n35195), .B(n35194), .Z(n35228) );
  XNOR U36093 ( .A(n35228), .B(sreg[1872]), .Z(n35230) );
  NAND U36094 ( .A(n35187), .B(sreg[1871]), .Z(n35191) );
  OR U36095 ( .A(n35189), .B(n35188), .Z(n35190) );
  AND U36096 ( .A(n35191), .B(n35190), .Z(n35229) );
  XOR U36097 ( .A(n35230), .B(n35229), .Z(c[1872]) );
  NANDN U36098 ( .A(n35193), .B(n35192), .Z(n35197) );
  NAND U36099 ( .A(n35195), .B(n35194), .Z(n35196) );
  NAND U36100 ( .A(n35197), .B(n35196), .Z(n35236) );
  NAND U36101 ( .A(b[0]), .B(a[857]), .Z(n35198) );
  XNOR U36102 ( .A(b[1]), .B(n35198), .Z(n35200) );
  NAND U36103 ( .A(n137), .B(a[856]), .Z(n35199) );
  AND U36104 ( .A(n35200), .B(n35199), .Z(n35253) );
  XOR U36105 ( .A(a[853]), .B(n42197), .Z(n35242) );
  NANDN U36106 ( .A(n35242), .B(n42173), .Z(n35203) );
  NANDN U36107 ( .A(n35201), .B(n42172), .Z(n35202) );
  NAND U36108 ( .A(n35203), .B(n35202), .Z(n35251) );
  NAND U36109 ( .A(b[7]), .B(a[849]), .Z(n35252) );
  XNOR U36110 ( .A(n35251), .B(n35252), .Z(n35254) );
  XOR U36111 ( .A(n35253), .B(n35254), .Z(n35260) );
  NANDN U36112 ( .A(n35204), .B(n42093), .Z(n35206) );
  XOR U36113 ( .A(n42134), .B(a[855]), .Z(n35245) );
  NANDN U36114 ( .A(n35245), .B(n42095), .Z(n35205) );
  NAND U36115 ( .A(n35206), .B(n35205), .Z(n35258) );
  NANDN U36116 ( .A(n35207), .B(n42231), .Z(n35209) );
  XOR U36117 ( .A(n233), .B(a[851]), .Z(n35248) );
  NANDN U36118 ( .A(n35248), .B(n42234), .Z(n35208) );
  AND U36119 ( .A(n35209), .B(n35208), .Z(n35257) );
  XNOR U36120 ( .A(n35258), .B(n35257), .Z(n35259) );
  XNOR U36121 ( .A(n35260), .B(n35259), .Z(n35264) );
  NANDN U36122 ( .A(n35211), .B(n35210), .Z(n35215) );
  NAND U36123 ( .A(n35213), .B(n35212), .Z(n35214) );
  AND U36124 ( .A(n35215), .B(n35214), .Z(n35263) );
  XOR U36125 ( .A(n35264), .B(n35263), .Z(n35265) );
  NANDN U36126 ( .A(n35217), .B(n35216), .Z(n35221) );
  NANDN U36127 ( .A(n35219), .B(n35218), .Z(n35220) );
  NAND U36128 ( .A(n35221), .B(n35220), .Z(n35266) );
  XOR U36129 ( .A(n35265), .B(n35266), .Z(n35233) );
  OR U36130 ( .A(n35223), .B(n35222), .Z(n35227) );
  NANDN U36131 ( .A(n35225), .B(n35224), .Z(n35226) );
  NAND U36132 ( .A(n35227), .B(n35226), .Z(n35234) );
  XNOR U36133 ( .A(n35233), .B(n35234), .Z(n35235) );
  XNOR U36134 ( .A(n35236), .B(n35235), .Z(n35269) );
  XNOR U36135 ( .A(n35269), .B(sreg[1873]), .Z(n35271) );
  NAND U36136 ( .A(n35228), .B(sreg[1872]), .Z(n35232) );
  OR U36137 ( .A(n35230), .B(n35229), .Z(n35231) );
  AND U36138 ( .A(n35232), .B(n35231), .Z(n35270) );
  XOR U36139 ( .A(n35271), .B(n35270), .Z(c[1873]) );
  NANDN U36140 ( .A(n35234), .B(n35233), .Z(n35238) );
  NAND U36141 ( .A(n35236), .B(n35235), .Z(n35237) );
  NAND U36142 ( .A(n35238), .B(n35237), .Z(n35277) );
  NAND U36143 ( .A(b[0]), .B(a[858]), .Z(n35239) );
  XNOR U36144 ( .A(b[1]), .B(n35239), .Z(n35241) );
  NAND U36145 ( .A(n137), .B(a[857]), .Z(n35240) );
  AND U36146 ( .A(n35241), .B(n35240), .Z(n35294) );
  XOR U36147 ( .A(a[854]), .B(n42197), .Z(n35283) );
  NANDN U36148 ( .A(n35283), .B(n42173), .Z(n35244) );
  NANDN U36149 ( .A(n35242), .B(n42172), .Z(n35243) );
  NAND U36150 ( .A(n35244), .B(n35243), .Z(n35292) );
  NAND U36151 ( .A(b[7]), .B(a[850]), .Z(n35293) );
  XNOR U36152 ( .A(n35292), .B(n35293), .Z(n35295) );
  XOR U36153 ( .A(n35294), .B(n35295), .Z(n35301) );
  NANDN U36154 ( .A(n35245), .B(n42093), .Z(n35247) );
  XOR U36155 ( .A(n42134), .B(a[856]), .Z(n35286) );
  NANDN U36156 ( .A(n35286), .B(n42095), .Z(n35246) );
  NAND U36157 ( .A(n35247), .B(n35246), .Z(n35299) );
  NANDN U36158 ( .A(n35248), .B(n42231), .Z(n35250) );
  XOR U36159 ( .A(n233), .B(a[852]), .Z(n35289) );
  NANDN U36160 ( .A(n35289), .B(n42234), .Z(n35249) );
  AND U36161 ( .A(n35250), .B(n35249), .Z(n35298) );
  XNOR U36162 ( .A(n35299), .B(n35298), .Z(n35300) );
  XNOR U36163 ( .A(n35301), .B(n35300), .Z(n35305) );
  NANDN U36164 ( .A(n35252), .B(n35251), .Z(n35256) );
  NAND U36165 ( .A(n35254), .B(n35253), .Z(n35255) );
  AND U36166 ( .A(n35256), .B(n35255), .Z(n35304) );
  XOR U36167 ( .A(n35305), .B(n35304), .Z(n35306) );
  NANDN U36168 ( .A(n35258), .B(n35257), .Z(n35262) );
  NANDN U36169 ( .A(n35260), .B(n35259), .Z(n35261) );
  NAND U36170 ( .A(n35262), .B(n35261), .Z(n35307) );
  XOR U36171 ( .A(n35306), .B(n35307), .Z(n35274) );
  OR U36172 ( .A(n35264), .B(n35263), .Z(n35268) );
  NANDN U36173 ( .A(n35266), .B(n35265), .Z(n35267) );
  NAND U36174 ( .A(n35268), .B(n35267), .Z(n35275) );
  XNOR U36175 ( .A(n35274), .B(n35275), .Z(n35276) );
  XNOR U36176 ( .A(n35277), .B(n35276), .Z(n35310) );
  XNOR U36177 ( .A(n35310), .B(sreg[1874]), .Z(n35312) );
  NAND U36178 ( .A(n35269), .B(sreg[1873]), .Z(n35273) );
  OR U36179 ( .A(n35271), .B(n35270), .Z(n35272) );
  AND U36180 ( .A(n35273), .B(n35272), .Z(n35311) );
  XOR U36181 ( .A(n35312), .B(n35311), .Z(c[1874]) );
  NANDN U36182 ( .A(n35275), .B(n35274), .Z(n35279) );
  NAND U36183 ( .A(n35277), .B(n35276), .Z(n35278) );
  NAND U36184 ( .A(n35279), .B(n35278), .Z(n35318) );
  NAND U36185 ( .A(b[0]), .B(a[859]), .Z(n35280) );
  XNOR U36186 ( .A(b[1]), .B(n35280), .Z(n35282) );
  NAND U36187 ( .A(n137), .B(a[858]), .Z(n35281) );
  AND U36188 ( .A(n35282), .B(n35281), .Z(n35335) );
  XOR U36189 ( .A(a[855]), .B(n42197), .Z(n35324) );
  NANDN U36190 ( .A(n35324), .B(n42173), .Z(n35285) );
  NANDN U36191 ( .A(n35283), .B(n42172), .Z(n35284) );
  NAND U36192 ( .A(n35285), .B(n35284), .Z(n35333) );
  NAND U36193 ( .A(b[7]), .B(a[851]), .Z(n35334) );
  XNOR U36194 ( .A(n35333), .B(n35334), .Z(n35336) );
  XOR U36195 ( .A(n35335), .B(n35336), .Z(n35342) );
  NANDN U36196 ( .A(n35286), .B(n42093), .Z(n35288) );
  XOR U36197 ( .A(n42134), .B(a[857]), .Z(n35327) );
  NANDN U36198 ( .A(n35327), .B(n42095), .Z(n35287) );
  NAND U36199 ( .A(n35288), .B(n35287), .Z(n35340) );
  NANDN U36200 ( .A(n35289), .B(n42231), .Z(n35291) );
  XOR U36201 ( .A(n233), .B(a[853]), .Z(n35330) );
  NANDN U36202 ( .A(n35330), .B(n42234), .Z(n35290) );
  AND U36203 ( .A(n35291), .B(n35290), .Z(n35339) );
  XNOR U36204 ( .A(n35340), .B(n35339), .Z(n35341) );
  XNOR U36205 ( .A(n35342), .B(n35341), .Z(n35346) );
  NANDN U36206 ( .A(n35293), .B(n35292), .Z(n35297) );
  NAND U36207 ( .A(n35295), .B(n35294), .Z(n35296) );
  AND U36208 ( .A(n35297), .B(n35296), .Z(n35345) );
  XOR U36209 ( .A(n35346), .B(n35345), .Z(n35347) );
  NANDN U36210 ( .A(n35299), .B(n35298), .Z(n35303) );
  NANDN U36211 ( .A(n35301), .B(n35300), .Z(n35302) );
  NAND U36212 ( .A(n35303), .B(n35302), .Z(n35348) );
  XOR U36213 ( .A(n35347), .B(n35348), .Z(n35315) );
  OR U36214 ( .A(n35305), .B(n35304), .Z(n35309) );
  NANDN U36215 ( .A(n35307), .B(n35306), .Z(n35308) );
  NAND U36216 ( .A(n35309), .B(n35308), .Z(n35316) );
  XNOR U36217 ( .A(n35315), .B(n35316), .Z(n35317) );
  XNOR U36218 ( .A(n35318), .B(n35317), .Z(n35351) );
  XNOR U36219 ( .A(n35351), .B(sreg[1875]), .Z(n35353) );
  NAND U36220 ( .A(n35310), .B(sreg[1874]), .Z(n35314) );
  OR U36221 ( .A(n35312), .B(n35311), .Z(n35313) );
  AND U36222 ( .A(n35314), .B(n35313), .Z(n35352) );
  XOR U36223 ( .A(n35353), .B(n35352), .Z(c[1875]) );
  NANDN U36224 ( .A(n35316), .B(n35315), .Z(n35320) );
  NAND U36225 ( .A(n35318), .B(n35317), .Z(n35319) );
  NAND U36226 ( .A(n35320), .B(n35319), .Z(n35359) );
  NAND U36227 ( .A(b[0]), .B(a[860]), .Z(n35321) );
  XNOR U36228 ( .A(b[1]), .B(n35321), .Z(n35323) );
  NAND U36229 ( .A(n137), .B(a[859]), .Z(n35322) );
  AND U36230 ( .A(n35323), .B(n35322), .Z(n35376) );
  XOR U36231 ( .A(a[856]), .B(n42197), .Z(n35365) );
  NANDN U36232 ( .A(n35365), .B(n42173), .Z(n35326) );
  NANDN U36233 ( .A(n35324), .B(n42172), .Z(n35325) );
  NAND U36234 ( .A(n35326), .B(n35325), .Z(n35374) );
  NAND U36235 ( .A(b[7]), .B(a[852]), .Z(n35375) );
  XNOR U36236 ( .A(n35374), .B(n35375), .Z(n35377) );
  XOR U36237 ( .A(n35376), .B(n35377), .Z(n35383) );
  NANDN U36238 ( .A(n35327), .B(n42093), .Z(n35329) );
  XOR U36239 ( .A(n42134), .B(a[858]), .Z(n35368) );
  NANDN U36240 ( .A(n35368), .B(n42095), .Z(n35328) );
  NAND U36241 ( .A(n35329), .B(n35328), .Z(n35381) );
  NANDN U36242 ( .A(n35330), .B(n42231), .Z(n35332) );
  XOR U36243 ( .A(n233), .B(a[854]), .Z(n35371) );
  NANDN U36244 ( .A(n35371), .B(n42234), .Z(n35331) );
  AND U36245 ( .A(n35332), .B(n35331), .Z(n35380) );
  XNOR U36246 ( .A(n35381), .B(n35380), .Z(n35382) );
  XNOR U36247 ( .A(n35383), .B(n35382), .Z(n35387) );
  NANDN U36248 ( .A(n35334), .B(n35333), .Z(n35338) );
  NAND U36249 ( .A(n35336), .B(n35335), .Z(n35337) );
  AND U36250 ( .A(n35338), .B(n35337), .Z(n35386) );
  XOR U36251 ( .A(n35387), .B(n35386), .Z(n35388) );
  NANDN U36252 ( .A(n35340), .B(n35339), .Z(n35344) );
  NANDN U36253 ( .A(n35342), .B(n35341), .Z(n35343) );
  NAND U36254 ( .A(n35344), .B(n35343), .Z(n35389) );
  XOR U36255 ( .A(n35388), .B(n35389), .Z(n35356) );
  OR U36256 ( .A(n35346), .B(n35345), .Z(n35350) );
  NANDN U36257 ( .A(n35348), .B(n35347), .Z(n35349) );
  NAND U36258 ( .A(n35350), .B(n35349), .Z(n35357) );
  XNOR U36259 ( .A(n35356), .B(n35357), .Z(n35358) );
  XNOR U36260 ( .A(n35359), .B(n35358), .Z(n35392) );
  XNOR U36261 ( .A(n35392), .B(sreg[1876]), .Z(n35394) );
  NAND U36262 ( .A(n35351), .B(sreg[1875]), .Z(n35355) );
  OR U36263 ( .A(n35353), .B(n35352), .Z(n35354) );
  AND U36264 ( .A(n35355), .B(n35354), .Z(n35393) );
  XOR U36265 ( .A(n35394), .B(n35393), .Z(c[1876]) );
  NANDN U36266 ( .A(n35357), .B(n35356), .Z(n35361) );
  NAND U36267 ( .A(n35359), .B(n35358), .Z(n35360) );
  NAND U36268 ( .A(n35361), .B(n35360), .Z(n35400) );
  NAND U36269 ( .A(b[0]), .B(a[861]), .Z(n35362) );
  XNOR U36270 ( .A(b[1]), .B(n35362), .Z(n35364) );
  NAND U36271 ( .A(n138), .B(a[860]), .Z(n35363) );
  AND U36272 ( .A(n35364), .B(n35363), .Z(n35417) );
  XOR U36273 ( .A(a[857]), .B(n42197), .Z(n35406) );
  NANDN U36274 ( .A(n35406), .B(n42173), .Z(n35367) );
  NANDN U36275 ( .A(n35365), .B(n42172), .Z(n35366) );
  NAND U36276 ( .A(n35367), .B(n35366), .Z(n35415) );
  NAND U36277 ( .A(b[7]), .B(a[853]), .Z(n35416) );
  XNOR U36278 ( .A(n35415), .B(n35416), .Z(n35418) );
  XOR U36279 ( .A(n35417), .B(n35418), .Z(n35424) );
  NANDN U36280 ( .A(n35368), .B(n42093), .Z(n35370) );
  XOR U36281 ( .A(n42134), .B(a[859]), .Z(n35409) );
  NANDN U36282 ( .A(n35409), .B(n42095), .Z(n35369) );
  NAND U36283 ( .A(n35370), .B(n35369), .Z(n35422) );
  NANDN U36284 ( .A(n35371), .B(n42231), .Z(n35373) );
  XOR U36285 ( .A(n233), .B(a[855]), .Z(n35412) );
  NANDN U36286 ( .A(n35412), .B(n42234), .Z(n35372) );
  AND U36287 ( .A(n35373), .B(n35372), .Z(n35421) );
  XNOR U36288 ( .A(n35422), .B(n35421), .Z(n35423) );
  XNOR U36289 ( .A(n35424), .B(n35423), .Z(n35428) );
  NANDN U36290 ( .A(n35375), .B(n35374), .Z(n35379) );
  NAND U36291 ( .A(n35377), .B(n35376), .Z(n35378) );
  AND U36292 ( .A(n35379), .B(n35378), .Z(n35427) );
  XOR U36293 ( .A(n35428), .B(n35427), .Z(n35429) );
  NANDN U36294 ( .A(n35381), .B(n35380), .Z(n35385) );
  NANDN U36295 ( .A(n35383), .B(n35382), .Z(n35384) );
  NAND U36296 ( .A(n35385), .B(n35384), .Z(n35430) );
  XOR U36297 ( .A(n35429), .B(n35430), .Z(n35397) );
  OR U36298 ( .A(n35387), .B(n35386), .Z(n35391) );
  NANDN U36299 ( .A(n35389), .B(n35388), .Z(n35390) );
  NAND U36300 ( .A(n35391), .B(n35390), .Z(n35398) );
  XNOR U36301 ( .A(n35397), .B(n35398), .Z(n35399) );
  XNOR U36302 ( .A(n35400), .B(n35399), .Z(n35433) );
  XNOR U36303 ( .A(n35433), .B(sreg[1877]), .Z(n35435) );
  NAND U36304 ( .A(n35392), .B(sreg[1876]), .Z(n35396) );
  OR U36305 ( .A(n35394), .B(n35393), .Z(n35395) );
  AND U36306 ( .A(n35396), .B(n35395), .Z(n35434) );
  XOR U36307 ( .A(n35435), .B(n35434), .Z(c[1877]) );
  NANDN U36308 ( .A(n35398), .B(n35397), .Z(n35402) );
  NAND U36309 ( .A(n35400), .B(n35399), .Z(n35401) );
  NAND U36310 ( .A(n35402), .B(n35401), .Z(n35441) );
  NAND U36311 ( .A(b[0]), .B(a[862]), .Z(n35403) );
  XNOR U36312 ( .A(b[1]), .B(n35403), .Z(n35405) );
  NAND U36313 ( .A(n138), .B(a[861]), .Z(n35404) );
  AND U36314 ( .A(n35405), .B(n35404), .Z(n35458) );
  XOR U36315 ( .A(a[858]), .B(n42197), .Z(n35447) );
  NANDN U36316 ( .A(n35447), .B(n42173), .Z(n35408) );
  NANDN U36317 ( .A(n35406), .B(n42172), .Z(n35407) );
  NAND U36318 ( .A(n35408), .B(n35407), .Z(n35456) );
  NAND U36319 ( .A(b[7]), .B(a[854]), .Z(n35457) );
  XNOR U36320 ( .A(n35456), .B(n35457), .Z(n35459) );
  XOR U36321 ( .A(n35458), .B(n35459), .Z(n35465) );
  NANDN U36322 ( .A(n35409), .B(n42093), .Z(n35411) );
  XOR U36323 ( .A(n42134), .B(a[860]), .Z(n35450) );
  NANDN U36324 ( .A(n35450), .B(n42095), .Z(n35410) );
  NAND U36325 ( .A(n35411), .B(n35410), .Z(n35463) );
  NANDN U36326 ( .A(n35412), .B(n42231), .Z(n35414) );
  XOR U36327 ( .A(n233), .B(a[856]), .Z(n35453) );
  NANDN U36328 ( .A(n35453), .B(n42234), .Z(n35413) );
  AND U36329 ( .A(n35414), .B(n35413), .Z(n35462) );
  XNOR U36330 ( .A(n35463), .B(n35462), .Z(n35464) );
  XNOR U36331 ( .A(n35465), .B(n35464), .Z(n35469) );
  NANDN U36332 ( .A(n35416), .B(n35415), .Z(n35420) );
  NAND U36333 ( .A(n35418), .B(n35417), .Z(n35419) );
  AND U36334 ( .A(n35420), .B(n35419), .Z(n35468) );
  XOR U36335 ( .A(n35469), .B(n35468), .Z(n35470) );
  NANDN U36336 ( .A(n35422), .B(n35421), .Z(n35426) );
  NANDN U36337 ( .A(n35424), .B(n35423), .Z(n35425) );
  NAND U36338 ( .A(n35426), .B(n35425), .Z(n35471) );
  XOR U36339 ( .A(n35470), .B(n35471), .Z(n35438) );
  OR U36340 ( .A(n35428), .B(n35427), .Z(n35432) );
  NANDN U36341 ( .A(n35430), .B(n35429), .Z(n35431) );
  NAND U36342 ( .A(n35432), .B(n35431), .Z(n35439) );
  XNOR U36343 ( .A(n35438), .B(n35439), .Z(n35440) );
  XNOR U36344 ( .A(n35441), .B(n35440), .Z(n35474) );
  XNOR U36345 ( .A(n35474), .B(sreg[1878]), .Z(n35476) );
  NAND U36346 ( .A(n35433), .B(sreg[1877]), .Z(n35437) );
  OR U36347 ( .A(n35435), .B(n35434), .Z(n35436) );
  AND U36348 ( .A(n35437), .B(n35436), .Z(n35475) );
  XOR U36349 ( .A(n35476), .B(n35475), .Z(c[1878]) );
  NANDN U36350 ( .A(n35439), .B(n35438), .Z(n35443) );
  NAND U36351 ( .A(n35441), .B(n35440), .Z(n35442) );
  NAND U36352 ( .A(n35443), .B(n35442), .Z(n35482) );
  NAND U36353 ( .A(b[0]), .B(a[863]), .Z(n35444) );
  XNOR U36354 ( .A(b[1]), .B(n35444), .Z(n35446) );
  NAND U36355 ( .A(n138), .B(a[862]), .Z(n35445) );
  AND U36356 ( .A(n35446), .B(n35445), .Z(n35499) );
  XOR U36357 ( .A(a[859]), .B(n42197), .Z(n35488) );
  NANDN U36358 ( .A(n35488), .B(n42173), .Z(n35449) );
  NANDN U36359 ( .A(n35447), .B(n42172), .Z(n35448) );
  NAND U36360 ( .A(n35449), .B(n35448), .Z(n35497) );
  NAND U36361 ( .A(b[7]), .B(a[855]), .Z(n35498) );
  XNOR U36362 ( .A(n35497), .B(n35498), .Z(n35500) );
  XOR U36363 ( .A(n35499), .B(n35500), .Z(n35506) );
  NANDN U36364 ( .A(n35450), .B(n42093), .Z(n35452) );
  XOR U36365 ( .A(n42134), .B(a[861]), .Z(n35491) );
  NANDN U36366 ( .A(n35491), .B(n42095), .Z(n35451) );
  NAND U36367 ( .A(n35452), .B(n35451), .Z(n35504) );
  NANDN U36368 ( .A(n35453), .B(n42231), .Z(n35455) );
  XOR U36369 ( .A(n233), .B(a[857]), .Z(n35494) );
  NANDN U36370 ( .A(n35494), .B(n42234), .Z(n35454) );
  AND U36371 ( .A(n35455), .B(n35454), .Z(n35503) );
  XNOR U36372 ( .A(n35504), .B(n35503), .Z(n35505) );
  XNOR U36373 ( .A(n35506), .B(n35505), .Z(n35510) );
  NANDN U36374 ( .A(n35457), .B(n35456), .Z(n35461) );
  NAND U36375 ( .A(n35459), .B(n35458), .Z(n35460) );
  AND U36376 ( .A(n35461), .B(n35460), .Z(n35509) );
  XOR U36377 ( .A(n35510), .B(n35509), .Z(n35511) );
  NANDN U36378 ( .A(n35463), .B(n35462), .Z(n35467) );
  NANDN U36379 ( .A(n35465), .B(n35464), .Z(n35466) );
  NAND U36380 ( .A(n35467), .B(n35466), .Z(n35512) );
  XOR U36381 ( .A(n35511), .B(n35512), .Z(n35479) );
  OR U36382 ( .A(n35469), .B(n35468), .Z(n35473) );
  NANDN U36383 ( .A(n35471), .B(n35470), .Z(n35472) );
  NAND U36384 ( .A(n35473), .B(n35472), .Z(n35480) );
  XNOR U36385 ( .A(n35479), .B(n35480), .Z(n35481) );
  XNOR U36386 ( .A(n35482), .B(n35481), .Z(n35515) );
  XNOR U36387 ( .A(n35515), .B(sreg[1879]), .Z(n35517) );
  NAND U36388 ( .A(n35474), .B(sreg[1878]), .Z(n35478) );
  OR U36389 ( .A(n35476), .B(n35475), .Z(n35477) );
  AND U36390 ( .A(n35478), .B(n35477), .Z(n35516) );
  XOR U36391 ( .A(n35517), .B(n35516), .Z(c[1879]) );
  NANDN U36392 ( .A(n35480), .B(n35479), .Z(n35484) );
  NAND U36393 ( .A(n35482), .B(n35481), .Z(n35483) );
  NAND U36394 ( .A(n35484), .B(n35483), .Z(n35523) );
  NAND U36395 ( .A(b[0]), .B(a[864]), .Z(n35485) );
  XNOR U36396 ( .A(b[1]), .B(n35485), .Z(n35487) );
  NAND U36397 ( .A(n138), .B(a[863]), .Z(n35486) );
  AND U36398 ( .A(n35487), .B(n35486), .Z(n35540) );
  XOR U36399 ( .A(a[860]), .B(n42197), .Z(n35529) );
  NANDN U36400 ( .A(n35529), .B(n42173), .Z(n35490) );
  NANDN U36401 ( .A(n35488), .B(n42172), .Z(n35489) );
  NAND U36402 ( .A(n35490), .B(n35489), .Z(n35538) );
  NAND U36403 ( .A(b[7]), .B(a[856]), .Z(n35539) );
  XNOR U36404 ( .A(n35538), .B(n35539), .Z(n35541) );
  XOR U36405 ( .A(n35540), .B(n35541), .Z(n35547) );
  NANDN U36406 ( .A(n35491), .B(n42093), .Z(n35493) );
  XOR U36407 ( .A(n42134), .B(a[862]), .Z(n35532) );
  NANDN U36408 ( .A(n35532), .B(n42095), .Z(n35492) );
  NAND U36409 ( .A(n35493), .B(n35492), .Z(n35545) );
  NANDN U36410 ( .A(n35494), .B(n42231), .Z(n35496) );
  XOR U36411 ( .A(n233), .B(a[858]), .Z(n35535) );
  NANDN U36412 ( .A(n35535), .B(n42234), .Z(n35495) );
  AND U36413 ( .A(n35496), .B(n35495), .Z(n35544) );
  XNOR U36414 ( .A(n35545), .B(n35544), .Z(n35546) );
  XNOR U36415 ( .A(n35547), .B(n35546), .Z(n35551) );
  NANDN U36416 ( .A(n35498), .B(n35497), .Z(n35502) );
  NAND U36417 ( .A(n35500), .B(n35499), .Z(n35501) );
  AND U36418 ( .A(n35502), .B(n35501), .Z(n35550) );
  XOR U36419 ( .A(n35551), .B(n35550), .Z(n35552) );
  NANDN U36420 ( .A(n35504), .B(n35503), .Z(n35508) );
  NANDN U36421 ( .A(n35506), .B(n35505), .Z(n35507) );
  NAND U36422 ( .A(n35508), .B(n35507), .Z(n35553) );
  XOR U36423 ( .A(n35552), .B(n35553), .Z(n35520) );
  OR U36424 ( .A(n35510), .B(n35509), .Z(n35514) );
  NANDN U36425 ( .A(n35512), .B(n35511), .Z(n35513) );
  NAND U36426 ( .A(n35514), .B(n35513), .Z(n35521) );
  XNOR U36427 ( .A(n35520), .B(n35521), .Z(n35522) );
  XNOR U36428 ( .A(n35523), .B(n35522), .Z(n35556) );
  XNOR U36429 ( .A(n35556), .B(sreg[1880]), .Z(n35558) );
  NAND U36430 ( .A(n35515), .B(sreg[1879]), .Z(n35519) );
  OR U36431 ( .A(n35517), .B(n35516), .Z(n35518) );
  AND U36432 ( .A(n35519), .B(n35518), .Z(n35557) );
  XOR U36433 ( .A(n35558), .B(n35557), .Z(c[1880]) );
  NANDN U36434 ( .A(n35521), .B(n35520), .Z(n35525) );
  NAND U36435 ( .A(n35523), .B(n35522), .Z(n35524) );
  NAND U36436 ( .A(n35525), .B(n35524), .Z(n35564) );
  NAND U36437 ( .A(b[0]), .B(a[865]), .Z(n35526) );
  XNOR U36438 ( .A(b[1]), .B(n35526), .Z(n35528) );
  NAND U36439 ( .A(n138), .B(a[864]), .Z(n35527) );
  AND U36440 ( .A(n35528), .B(n35527), .Z(n35581) );
  XOR U36441 ( .A(a[861]), .B(n42197), .Z(n35570) );
  NANDN U36442 ( .A(n35570), .B(n42173), .Z(n35531) );
  NANDN U36443 ( .A(n35529), .B(n42172), .Z(n35530) );
  NAND U36444 ( .A(n35531), .B(n35530), .Z(n35579) );
  NAND U36445 ( .A(b[7]), .B(a[857]), .Z(n35580) );
  XNOR U36446 ( .A(n35579), .B(n35580), .Z(n35582) );
  XOR U36447 ( .A(n35581), .B(n35582), .Z(n35588) );
  NANDN U36448 ( .A(n35532), .B(n42093), .Z(n35534) );
  XOR U36449 ( .A(n42134), .B(a[863]), .Z(n35573) );
  NANDN U36450 ( .A(n35573), .B(n42095), .Z(n35533) );
  NAND U36451 ( .A(n35534), .B(n35533), .Z(n35586) );
  NANDN U36452 ( .A(n35535), .B(n42231), .Z(n35537) );
  XOR U36453 ( .A(n233), .B(a[859]), .Z(n35576) );
  NANDN U36454 ( .A(n35576), .B(n42234), .Z(n35536) );
  AND U36455 ( .A(n35537), .B(n35536), .Z(n35585) );
  XNOR U36456 ( .A(n35586), .B(n35585), .Z(n35587) );
  XNOR U36457 ( .A(n35588), .B(n35587), .Z(n35592) );
  NANDN U36458 ( .A(n35539), .B(n35538), .Z(n35543) );
  NAND U36459 ( .A(n35541), .B(n35540), .Z(n35542) );
  AND U36460 ( .A(n35543), .B(n35542), .Z(n35591) );
  XOR U36461 ( .A(n35592), .B(n35591), .Z(n35593) );
  NANDN U36462 ( .A(n35545), .B(n35544), .Z(n35549) );
  NANDN U36463 ( .A(n35547), .B(n35546), .Z(n35548) );
  NAND U36464 ( .A(n35549), .B(n35548), .Z(n35594) );
  XOR U36465 ( .A(n35593), .B(n35594), .Z(n35561) );
  OR U36466 ( .A(n35551), .B(n35550), .Z(n35555) );
  NANDN U36467 ( .A(n35553), .B(n35552), .Z(n35554) );
  NAND U36468 ( .A(n35555), .B(n35554), .Z(n35562) );
  XNOR U36469 ( .A(n35561), .B(n35562), .Z(n35563) );
  XNOR U36470 ( .A(n35564), .B(n35563), .Z(n35597) );
  XNOR U36471 ( .A(n35597), .B(sreg[1881]), .Z(n35599) );
  NAND U36472 ( .A(n35556), .B(sreg[1880]), .Z(n35560) );
  OR U36473 ( .A(n35558), .B(n35557), .Z(n35559) );
  AND U36474 ( .A(n35560), .B(n35559), .Z(n35598) );
  XOR U36475 ( .A(n35599), .B(n35598), .Z(c[1881]) );
  NANDN U36476 ( .A(n35562), .B(n35561), .Z(n35566) );
  NAND U36477 ( .A(n35564), .B(n35563), .Z(n35565) );
  NAND U36478 ( .A(n35566), .B(n35565), .Z(n35605) );
  NAND U36479 ( .A(b[0]), .B(a[866]), .Z(n35567) );
  XNOR U36480 ( .A(b[1]), .B(n35567), .Z(n35569) );
  NAND U36481 ( .A(n138), .B(a[865]), .Z(n35568) );
  AND U36482 ( .A(n35569), .B(n35568), .Z(n35622) );
  XOR U36483 ( .A(a[862]), .B(n42197), .Z(n35611) );
  NANDN U36484 ( .A(n35611), .B(n42173), .Z(n35572) );
  NANDN U36485 ( .A(n35570), .B(n42172), .Z(n35571) );
  NAND U36486 ( .A(n35572), .B(n35571), .Z(n35620) );
  NAND U36487 ( .A(b[7]), .B(a[858]), .Z(n35621) );
  XNOR U36488 ( .A(n35620), .B(n35621), .Z(n35623) );
  XOR U36489 ( .A(n35622), .B(n35623), .Z(n35629) );
  NANDN U36490 ( .A(n35573), .B(n42093), .Z(n35575) );
  XOR U36491 ( .A(n42134), .B(a[864]), .Z(n35614) );
  NANDN U36492 ( .A(n35614), .B(n42095), .Z(n35574) );
  NAND U36493 ( .A(n35575), .B(n35574), .Z(n35627) );
  NANDN U36494 ( .A(n35576), .B(n42231), .Z(n35578) );
  XOR U36495 ( .A(n233), .B(a[860]), .Z(n35617) );
  NANDN U36496 ( .A(n35617), .B(n42234), .Z(n35577) );
  AND U36497 ( .A(n35578), .B(n35577), .Z(n35626) );
  XNOR U36498 ( .A(n35627), .B(n35626), .Z(n35628) );
  XNOR U36499 ( .A(n35629), .B(n35628), .Z(n35633) );
  NANDN U36500 ( .A(n35580), .B(n35579), .Z(n35584) );
  NAND U36501 ( .A(n35582), .B(n35581), .Z(n35583) );
  AND U36502 ( .A(n35584), .B(n35583), .Z(n35632) );
  XOR U36503 ( .A(n35633), .B(n35632), .Z(n35634) );
  NANDN U36504 ( .A(n35586), .B(n35585), .Z(n35590) );
  NANDN U36505 ( .A(n35588), .B(n35587), .Z(n35589) );
  NAND U36506 ( .A(n35590), .B(n35589), .Z(n35635) );
  XOR U36507 ( .A(n35634), .B(n35635), .Z(n35602) );
  OR U36508 ( .A(n35592), .B(n35591), .Z(n35596) );
  NANDN U36509 ( .A(n35594), .B(n35593), .Z(n35595) );
  NAND U36510 ( .A(n35596), .B(n35595), .Z(n35603) );
  XNOR U36511 ( .A(n35602), .B(n35603), .Z(n35604) );
  XNOR U36512 ( .A(n35605), .B(n35604), .Z(n35638) );
  XNOR U36513 ( .A(n35638), .B(sreg[1882]), .Z(n35640) );
  NAND U36514 ( .A(n35597), .B(sreg[1881]), .Z(n35601) );
  OR U36515 ( .A(n35599), .B(n35598), .Z(n35600) );
  AND U36516 ( .A(n35601), .B(n35600), .Z(n35639) );
  XOR U36517 ( .A(n35640), .B(n35639), .Z(c[1882]) );
  NANDN U36518 ( .A(n35603), .B(n35602), .Z(n35607) );
  NAND U36519 ( .A(n35605), .B(n35604), .Z(n35606) );
  NAND U36520 ( .A(n35607), .B(n35606), .Z(n35646) );
  NAND U36521 ( .A(b[0]), .B(a[867]), .Z(n35608) );
  XNOR U36522 ( .A(b[1]), .B(n35608), .Z(n35610) );
  NAND U36523 ( .A(n138), .B(a[866]), .Z(n35609) );
  AND U36524 ( .A(n35610), .B(n35609), .Z(n35663) );
  XOR U36525 ( .A(a[863]), .B(n42197), .Z(n35652) );
  NANDN U36526 ( .A(n35652), .B(n42173), .Z(n35613) );
  NANDN U36527 ( .A(n35611), .B(n42172), .Z(n35612) );
  NAND U36528 ( .A(n35613), .B(n35612), .Z(n35661) );
  NAND U36529 ( .A(b[7]), .B(a[859]), .Z(n35662) );
  XNOR U36530 ( .A(n35661), .B(n35662), .Z(n35664) );
  XOR U36531 ( .A(n35663), .B(n35664), .Z(n35670) );
  NANDN U36532 ( .A(n35614), .B(n42093), .Z(n35616) );
  XOR U36533 ( .A(n42134), .B(a[865]), .Z(n35655) );
  NANDN U36534 ( .A(n35655), .B(n42095), .Z(n35615) );
  NAND U36535 ( .A(n35616), .B(n35615), .Z(n35668) );
  NANDN U36536 ( .A(n35617), .B(n42231), .Z(n35619) );
  XOR U36537 ( .A(n233), .B(a[861]), .Z(n35658) );
  NANDN U36538 ( .A(n35658), .B(n42234), .Z(n35618) );
  AND U36539 ( .A(n35619), .B(n35618), .Z(n35667) );
  XNOR U36540 ( .A(n35668), .B(n35667), .Z(n35669) );
  XNOR U36541 ( .A(n35670), .B(n35669), .Z(n35674) );
  NANDN U36542 ( .A(n35621), .B(n35620), .Z(n35625) );
  NAND U36543 ( .A(n35623), .B(n35622), .Z(n35624) );
  AND U36544 ( .A(n35625), .B(n35624), .Z(n35673) );
  XOR U36545 ( .A(n35674), .B(n35673), .Z(n35675) );
  NANDN U36546 ( .A(n35627), .B(n35626), .Z(n35631) );
  NANDN U36547 ( .A(n35629), .B(n35628), .Z(n35630) );
  NAND U36548 ( .A(n35631), .B(n35630), .Z(n35676) );
  XOR U36549 ( .A(n35675), .B(n35676), .Z(n35643) );
  OR U36550 ( .A(n35633), .B(n35632), .Z(n35637) );
  NANDN U36551 ( .A(n35635), .B(n35634), .Z(n35636) );
  NAND U36552 ( .A(n35637), .B(n35636), .Z(n35644) );
  XNOR U36553 ( .A(n35643), .B(n35644), .Z(n35645) );
  XNOR U36554 ( .A(n35646), .B(n35645), .Z(n35679) );
  XNOR U36555 ( .A(n35679), .B(sreg[1883]), .Z(n35681) );
  NAND U36556 ( .A(n35638), .B(sreg[1882]), .Z(n35642) );
  OR U36557 ( .A(n35640), .B(n35639), .Z(n35641) );
  AND U36558 ( .A(n35642), .B(n35641), .Z(n35680) );
  XOR U36559 ( .A(n35681), .B(n35680), .Z(c[1883]) );
  NANDN U36560 ( .A(n35644), .B(n35643), .Z(n35648) );
  NAND U36561 ( .A(n35646), .B(n35645), .Z(n35647) );
  NAND U36562 ( .A(n35648), .B(n35647), .Z(n35687) );
  NAND U36563 ( .A(b[0]), .B(a[868]), .Z(n35649) );
  XNOR U36564 ( .A(b[1]), .B(n35649), .Z(n35651) );
  NAND U36565 ( .A(n139), .B(a[867]), .Z(n35650) );
  AND U36566 ( .A(n35651), .B(n35650), .Z(n35704) );
  XOR U36567 ( .A(a[864]), .B(n42197), .Z(n35693) );
  NANDN U36568 ( .A(n35693), .B(n42173), .Z(n35654) );
  NANDN U36569 ( .A(n35652), .B(n42172), .Z(n35653) );
  NAND U36570 ( .A(n35654), .B(n35653), .Z(n35702) );
  NAND U36571 ( .A(b[7]), .B(a[860]), .Z(n35703) );
  XNOR U36572 ( .A(n35702), .B(n35703), .Z(n35705) );
  XOR U36573 ( .A(n35704), .B(n35705), .Z(n35711) );
  NANDN U36574 ( .A(n35655), .B(n42093), .Z(n35657) );
  XOR U36575 ( .A(n42134), .B(a[866]), .Z(n35696) );
  NANDN U36576 ( .A(n35696), .B(n42095), .Z(n35656) );
  NAND U36577 ( .A(n35657), .B(n35656), .Z(n35709) );
  NANDN U36578 ( .A(n35658), .B(n42231), .Z(n35660) );
  XOR U36579 ( .A(n233), .B(a[862]), .Z(n35699) );
  NANDN U36580 ( .A(n35699), .B(n42234), .Z(n35659) );
  AND U36581 ( .A(n35660), .B(n35659), .Z(n35708) );
  XNOR U36582 ( .A(n35709), .B(n35708), .Z(n35710) );
  XNOR U36583 ( .A(n35711), .B(n35710), .Z(n35715) );
  NANDN U36584 ( .A(n35662), .B(n35661), .Z(n35666) );
  NAND U36585 ( .A(n35664), .B(n35663), .Z(n35665) );
  AND U36586 ( .A(n35666), .B(n35665), .Z(n35714) );
  XOR U36587 ( .A(n35715), .B(n35714), .Z(n35716) );
  NANDN U36588 ( .A(n35668), .B(n35667), .Z(n35672) );
  NANDN U36589 ( .A(n35670), .B(n35669), .Z(n35671) );
  NAND U36590 ( .A(n35672), .B(n35671), .Z(n35717) );
  XOR U36591 ( .A(n35716), .B(n35717), .Z(n35684) );
  OR U36592 ( .A(n35674), .B(n35673), .Z(n35678) );
  NANDN U36593 ( .A(n35676), .B(n35675), .Z(n35677) );
  NAND U36594 ( .A(n35678), .B(n35677), .Z(n35685) );
  XNOR U36595 ( .A(n35684), .B(n35685), .Z(n35686) );
  XNOR U36596 ( .A(n35687), .B(n35686), .Z(n35720) );
  XNOR U36597 ( .A(n35720), .B(sreg[1884]), .Z(n35722) );
  NAND U36598 ( .A(n35679), .B(sreg[1883]), .Z(n35683) );
  OR U36599 ( .A(n35681), .B(n35680), .Z(n35682) );
  AND U36600 ( .A(n35683), .B(n35682), .Z(n35721) );
  XOR U36601 ( .A(n35722), .B(n35721), .Z(c[1884]) );
  NANDN U36602 ( .A(n35685), .B(n35684), .Z(n35689) );
  NAND U36603 ( .A(n35687), .B(n35686), .Z(n35688) );
  NAND U36604 ( .A(n35689), .B(n35688), .Z(n35728) );
  NAND U36605 ( .A(b[0]), .B(a[869]), .Z(n35690) );
  XNOR U36606 ( .A(b[1]), .B(n35690), .Z(n35692) );
  NAND U36607 ( .A(n139), .B(a[868]), .Z(n35691) );
  AND U36608 ( .A(n35692), .B(n35691), .Z(n35745) );
  XOR U36609 ( .A(a[865]), .B(n42197), .Z(n35734) );
  NANDN U36610 ( .A(n35734), .B(n42173), .Z(n35695) );
  NANDN U36611 ( .A(n35693), .B(n42172), .Z(n35694) );
  NAND U36612 ( .A(n35695), .B(n35694), .Z(n35743) );
  NAND U36613 ( .A(b[7]), .B(a[861]), .Z(n35744) );
  XNOR U36614 ( .A(n35743), .B(n35744), .Z(n35746) );
  XOR U36615 ( .A(n35745), .B(n35746), .Z(n35752) );
  NANDN U36616 ( .A(n35696), .B(n42093), .Z(n35698) );
  XOR U36617 ( .A(n42134), .B(a[867]), .Z(n35737) );
  NANDN U36618 ( .A(n35737), .B(n42095), .Z(n35697) );
  NAND U36619 ( .A(n35698), .B(n35697), .Z(n35750) );
  NANDN U36620 ( .A(n35699), .B(n42231), .Z(n35701) );
  XOR U36621 ( .A(n234), .B(a[863]), .Z(n35740) );
  NANDN U36622 ( .A(n35740), .B(n42234), .Z(n35700) );
  AND U36623 ( .A(n35701), .B(n35700), .Z(n35749) );
  XNOR U36624 ( .A(n35750), .B(n35749), .Z(n35751) );
  XNOR U36625 ( .A(n35752), .B(n35751), .Z(n35756) );
  NANDN U36626 ( .A(n35703), .B(n35702), .Z(n35707) );
  NAND U36627 ( .A(n35705), .B(n35704), .Z(n35706) );
  AND U36628 ( .A(n35707), .B(n35706), .Z(n35755) );
  XOR U36629 ( .A(n35756), .B(n35755), .Z(n35757) );
  NANDN U36630 ( .A(n35709), .B(n35708), .Z(n35713) );
  NANDN U36631 ( .A(n35711), .B(n35710), .Z(n35712) );
  NAND U36632 ( .A(n35713), .B(n35712), .Z(n35758) );
  XOR U36633 ( .A(n35757), .B(n35758), .Z(n35725) );
  OR U36634 ( .A(n35715), .B(n35714), .Z(n35719) );
  NANDN U36635 ( .A(n35717), .B(n35716), .Z(n35718) );
  NAND U36636 ( .A(n35719), .B(n35718), .Z(n35726) );
  XNOR U36637 ( .A(n35725), .B(n35726), .Z(n35727) );
  XNOR U36638 ( .A(n35728), .B(n35727), .Z(n35761) );
  XNOR U36639 ( .A(n35761), .B(sreg[1885]), .Z(n35763) );
  NAND U36640 ( .A(n35720), .B(sreg[1884]), .Z(n35724) );
  OR U36641 ( .A(n35722), .B(n35721), .Z(n35723) );
  AND U36642 ( .A(n35724), .B(n35723), .Z(n35762) );
  XOR U36643 ( .A(n35763), .B(n35762), .Z(c[1885]) );
  NANDN U36644 ( .A(n35726), .B(n35725), .Z(n35730) );
  NAND U36645 ( .A(n35728), .B(n35727), .Z(n35729) );
  NAND U36646 ( .A(n35730), .B(n35729), .Z(n35769) );
  NAND U36647 ( .A(b[0]), .B(a[870]), .Z(n35731) );
  XNOR U36648 ( .A(b[1]), .B(n35731), .Z(n35733) );
  NAND U36649 ( .A(n139), .B(a[869]), .Z(n35732) );
  AND U36650 ( .A(n35733), .B(n35732), .Z(n35786) );
  XOR U36651 ( .A(a[866]), .B(n42197), .Z(n35775) );
  NANDN U36652 ( .A(n35775), .B(n42173), .Z(n35736) );
  NANDN U36653 ( .A(n35734), .B(n42172), .Z(n35735) );
  NAND U36654 ( .A(n35736), .B(n35735), .Z(n35784) );
  NAND U36655 ( .A(b[7]), .B(a[862]), .Z(n35785) );
  XNOR U36656 ( .A(n35784), .B(n35785), .Z(n35787) );
  XOR U36657 ( .A(n35786), .B(n35787), .Z(n35793) );
  NANDN U36658 ( .A(n35737), .B(n42093), .Z(n35739) );
  XOR U36659 ( .A(n42134), .B(a[868]), .Z(n35778) );
  NANDN U36660 ( .A(n35778), .B(n42095), .Z(n35738) );
  NAND U36661 ( .A(n35739), .B(n35738), .Z(n35791) );
  NANDN U36662 ( .A(n35740), .B(n42231), .Z(n35742) );
  XOR U36663 ( .A(n234), .B(a[864]), .Z(n35781) );
  NANDN U36664 ( .A(n35781), .B(n42234), .Z(n35741) );
  AND U36665 ( .A(n35742), .B(n35741), .Z(n35790) );
  XNOR U36666 ( .A(n35791), .B(n35790), .Z(n35792) );
  XNOR U36667 ( .A(n35793), .B(n35792), .Z(n35797) );
  NANDN U36668 ( .A(n35744), .B(n35743), .Z(n35748) );
  NAND U36669 ( .A(n35746), .B(n35745), .Z(n35747) );
  AND U36670 ( .A(n35748), .B(n35747), .Z(n35796) );
  XOR U36671 ( .A(n35797), .B(n35796), .Z(n35798) );
  NANDN U36672 ( .A(n35750), .B(n35749), .Z(n35754) );
  NANDN U36673 ( .A(n35752), .B(n35751), .Z(n35753) );
  NAND U36674 ( .A(n35754), .B(n35753), .Z(n35799) );
  XOR U36675 ( .A(n35798), .B(n35799), .Z(n35766) );
  OR U36676 ( .A(n35756), .B(n35755), .Z(n35760) );
  NANDN U36677 ( .A(n35758), .B(n35757), .Z(n35759) );
  NAND U36678 ( .A(n35760), .B(n35759), .Z(n35767) );
  XNOR U36679 ( .A(n35766), .B(n35767), .Z(n35768) );
  XNOR U36680 ( .A(n35769), .B(n35768), .Z(n35802) );
  XNOR U36681 ( .A(n35802), .B(sreg[1886]), .Z(n35804) );
  NAND U36682 ( .A(n35761), .B(sreg[1885]), .Z(n35765) );
  OR U36683 ( .A(n35763), .B(n35762), .Z(n35764) );
  AND U36684 ( .A(n35765), .B(n35764), .Z(n35803) );
  XOR U36685 ( .A(n35804), .B(n35803), .Z(c[1886]) );
  NANDN U36686 ( .A(n35767), .B(n35766), .Z(n35771) );
  NAND U36687 ( .A(n35769), .B(n35768), .Z(n35770) );
  NAND U36688 ( .A(n35771), .B(n35770), .Z(n35810) );
  NAND U36689 ( .A(b[0]), .B(a[871]), .Z(n35772) );
  XNOR U36690 ( .A(b[1]), .B(n35772), .Z(n35774) );
  NAND U36691 ( .A(n139), .B(a[870]), .Z(n35773) );
  AND U36692 ( .A(n35774), .B(n35773), .Z(n35827) );
  XOR U36693 ( .A(a[867]), .B(n42197), .Z(n35816) );
  NANDN U36694 ( .A(n35816), .B(n42173), .Z(n35777) );
  NANDN U36695 ( .A(n35775), .B(n42172), .Z(n35776) );
  NAND U36696 ( .A(n35777), .B(n35776), .Z(n35825) );
  NAND U36697 ( .A(b[7]), .B(a[863]), .Z(n35826) );
  XNOR U36698 ( .A(n35825), .B(n35826), .Z(n35828) );
  XOR U36699 ( .A(n35827), .B(n35828), .Z(n35834) );
  NANDN U36700 ( .A(n35778), .B(n42093), .Z(n35780) );
  XOR U36701 ( .A(n42134), .B(a[869]), .Z(n35819) );
  NANDN U36702 ( .A(n35819), .B(n42095), .Z(n35779) );
  NAND U36703 ( .A(n35780), .B(n35779), .Z(n35832) );
  NANDN U36704 ( .A(n35781), .B(n42231), .Z(n35783) );
  XOR U36705 ( .A(n234), .B(a[865]), .Z(n35822) );
  NANDN U36706 ( .A(n35822), .B(n42234), .Z(n35782) );
  AND U36707 ( .A(n35783), .B(n35782), .Z(n35831) );
  XNOR U36708 ( .A(n35832), .B(n35831), .Z(n35833) );
  XNOR U36709 ( .A(n35834), .B(n35833), .Z(n35838) );
  NANDN U36710 ( .A(n35785), .B(n35784), .Z(n35789) );
  NAND U36711 ( .A(n35787), .B(n35786), .Z(n35788) );
  AND U36712 ( .A(n35789), .B(n35788), .Z(n35837) );
  XOR U36713 ( .A(n35838), .B(n35837), .Z(n35839) );
  NANDN U36714 ( .A(n35791), .B(n35790), .Z(n35795) );
  NANDN U36715 ( .A(n35793), .B(n35792), .Z(n35794) );
  NAND U36716 ( .A(n35795), .B(n35794), .Z(n35840) );
  XOR U36717 ( .A(n35839), .B(n35840), .Z(n35807) );
  OR U36718 ( .A(n35797), .B(n35796), .Z(n35801) );
  NANDN U36719 ( .A(n35799), .B(n35798), .Z(n35800) );
  NAND U36720 ( .A(n35801), .B(n35800), .Z(n35808) );
  XNOR U36721 ( .A(n35807), .B(n35808), .Z(n35809) );
  XNOR U36722 ( .A(n35810), .B(n35809), .Z(n35843) );
  XNOR U36723 ( .A(n35843), .B(sreg[1887]), .Z(n35845) );
  NAND U36724 ( .A(n35802), .B(sreg[1886]), .Z(n35806) );
  OR U36725 ( .A(n35804), .B(n35803), .Z(n35805) );
  AND U36726 ( .A(n35806), .B(n35805), .Z(n35844) );
  XOR U36727 ( .A(n35845), .B(n35844), .Z(c[1887]) );
  NANDN U36728 ( .A(n35808), .B(n35807), .Z(n35812) );
  NAND U36729 ( .A(n35810), .B(n35809), .Z(n35811) );
  NAND U36730 ( .A(n35812), .B(n35811), .Z(n35851) );
  NAND U36731 ( .A(b[0]), .B(a[872]), .Z(n35813) );
  XNOR U36732 ( .A(b[1]), .B(n35813), .Z(n35815) );
  NAND U36733 ( .A(n139), .B(a[871]), .Z(n35814) );
  AND U36734 ( .A(n35815), .B(n35814), .Z(n35868) );
  XOR U36735 ( .A(a[868]), .B(n42197), .Z(n35857) );
  NANDN U36736 ( .A(n35857), .B(n42173), .Z(n35818) );
  NANDN U36737 ( .A(n35816), .B(n42172), .Z(n35817) );
  NAND U36738 ( .A(n35818), .B(n35817), .Z(n35866) );
  NAND U36739 ( .A(b[7]), .B(a[864]), .Z(n35867) );
  XNOR U36740 ( .A(n35866), .B(n35867), .Z(n35869) );
  XOR U36741 ( .A(n35868), .B(n35869), .Z(n35875) );
  NANDN U36742 ( .A(n35819), .B(n42093), .Z(n35821) );
  XOR U36743 ( .A(n42134), .B(a[870]), .Z(n35860) );
  NANDN U36744 ( .A(n35860), .B(n42095), .Z(n35820) );
  NAND U36745 ( .A(n35821), .B(n35820), .Z(n35873) );
  NANDN U36746 ( .A(n35822), .B(n42231), .Z(n35824) );
  XOR U36747 ( .A(n234), .B(a[866]), .Z(n35863) );
  NANDN U36748 ( .A(n35863), .B(n42234), .Z(n35823) );
  AND U36749 ( .A(n35824), .B(n35823), .Z(n35872) );
  XNOR U36750 ( .A(n35873), .B(n35872), .Z(n35874) );
  XNOR U36751 ( .A(n35875), .B(n35874), .Z(n35879) );
  NANDN U36752 ( .A(n35826), .B(n35825), .Z(n35830) );
  NAND U36753 ( .A(n35828), .B(n35827), .Z(n35829) );
  AND U36754 ( .A(n35830), .B(n35829), .Z(n35878) );
  XOR U36755 ( .A(n35879), .B(n35878), .Z(n35880) );
  NANDN U36756 ( .A(n35832), .B(n35831), .Z(n35836) );
  NANDN U36757 ( .A(n35834), .B(n35833), .Z(n35835) );
  NAND U36758 ( .A(n35836), .B(n35835), .Z(n35881) );
  XOR U36759 ( .A(n35880), .B(n35881), .Z(n35848) );
  OR U36760 ( .A(n35838), .B(n35837), .Z(n35842) );
  NANDN U36761 ( .A(n35840), .B(n35839), .Z(n35841) );
  NAND U36762 ( .A(n35842), .B(n35841), .Z(n35849) );
  XNOR U36763 ( .A(n35848), .B(n35849), .Z(n35850) );
  XNOR U36764 ( .A(n35851), .B(n35850), .Z(n35884) );
  XNOR U36765 ( .A(n35884), .B(sreg[1888]), .Z(n35886) );
  NAND U36766 ( .A(n35843), .B(sreg[1887]), .Z(n35847) );
  OR U36767 ( .A(n35845), .B(n35844), .Z(n35846) );
  AND U36768 ( .A(n35847), .B(n35846), .Z(n35885) );
  XOR U36769 ( .A(n35886), .B(n35885), .Z(c[1888]) );
  NANDN U36770 ( .A(n35849), .B(n35848), .Z(n35853) );
  NAND U36771 ( .A(n35851), .B(n35850), .Z(n35852) );
  NAND U36772 ( .A(n35853), .B(n35852), .Z(n35892) );
  NAND U36773 ( .A(b[0]), .B(a[873]), .Z(n35854) );
  XNOR U36774 ( .A(b[1]), .B(n35854), .Z(n35856) );
  NAND U36775 ( .A(n139), .B(a[872]), .Z(n35855) );
  AND U36776 ( .A(n35856), .B(n35855), .Z(n35909) );
  XOR U36777 ( .A(a[869]), .B(n42197), .Z(n35898) );
  NANDN U36778 ( .A(n35898), .B(n42173), .Z(n35859) );
  NANDN U36779 ( .A(n35857), .B(n42172), .Z(n35858) );
  NAND U36780 ( .A(n35859), .B(n35858), .Z(n35907) );
  NAND U36781 ( .A(b[7]), .B(a[865]), .Z(n35908) );
  XNOR U36782 ( .A(n35907), .B(n35908), .Z(n35910) );
  XOR U36783 ( .A(n35909), .B(n35910), .Z(n35916) );
  NANDN U36784 ( .A(n35860), .B(n42093), .Z(n35862) );
  XOR U36785 ( .A(n42134), .B(a[871]), .Z(n35901) );
  NANDN U36786 ( .A(n35901), .B(n42095), .Z(n35861) );
  NAND U36787 ( .A(n35862), .B(n35861), .Z(n35914) );
  NANDN U36788 ( .A(n35863), .B(n42231), .Z(n35865) );
  XOR U36789 ( .A(n234), .B(a[867]), .Z(n35904) );
  NANDN U36790 ( .A(n35904), .B(n42234), .Z(n35864) );
  AND U36791 ( .A(n35865), .B(n35864), .Z(n35913) );
  XNOR U36792 ( .A(n35914), .B(n35913), .Z(n35915) );
  XNOR U36793 ( .A(n35916), .B(n35915), .Z(n35920) );
  NANDN U36794 ( .A(n35867), .B(n35866), .Z(n35871) );
  NAND U36795 ( .A(n35869), .B(n35868), .Z(n35870) );
  AND U36796 ( .A(n35871), .B(n35870), .Z(n35919) );
  XOR U36797 ( .A(n35920), .B(n35919), .Z(n35921) );
  NANDN U36798 ( .A(n35873), .B(n35872), .Z(n35877) );
  NANDN U36799 ( .A(n35875), .B(n35874), .Z(n35876) );
  NAND U36800 ( .A(n35877), .B(n35876), .Z(n35922) );
  XOR U36801 ( .A(n35921), .B(n35922), .Z(n35889) );
  OR U36802 ( .A(n35879), .B(n35878), .Z(n35883) );
  NANDN U36803 ( .A(n35881), .B(n35880), .Z(n35882) );
  NAND U36804 ( .A(n35883), .B(n35882), .Z(n35890) );
  XNOR U36805 ( .A(n35889), .B(n35890), .Z(n35891) );
  XNOR U36806 ( .A(n35892), .B(n35891), .Z(n35925) );
  XNOR U36807 ( .A(n35925), .B(sreg[1889]), .Z(n35927) );
  NAND U36808 ( .A(n35884), .B(sreg[1888]), .Z(n35888) );
  OR U36809 ( .A(n35886), .B(n35885), .Z(n35887) );
  AND U36810 ( .A(n35888), .B(n35887), .Z(n35926) );
  XOR U36811 ( .A(n35927), .B(n35926), .Z(c[1889]) );
  NANDN U36812 ( .A(n35890), .B(n35889), .Z(n35894) );
  NAND U36813 ( .A(n35892), .B(n35891), .Z(n35893) );
  NAND U36814 ( .A(n35894), .B(n35893), .Z(n35933) );
  NAND U36815 ( .A(b[0]), .B(a[874]), .Z(n35895) );
  XNOR U36816 ( .A(b[1]), .B(n35895), .Z(n35897) );
  NAND U36817 ( .A(n139), .B(a[873]), .Z(n35896) );
  AND U36818 ( .A(n35897), .B(n35896), .Z(n35950) );
  XOR U36819 ( .A(a[870]), .B(n42197), .Z(n35939) );
  NANDN U36820 ( .A(n35939), .B(n42173), .Z(n35900) );
  NANDN U36821 ( .A(n35898), .B(n42172), .Z(n35899) );
  NAND U36822 ( .A(n35900), .B(n35899), .Z(n35948) );
  NAND U36823 ( .A(b[7]), .B(a[866]), .Z(n35949) );
  XNOR U36824 ( .A(n35948), .B(n35949), .Z(n35951) );
  XOR U36825 ( .A(n35950), .B(n35951), .Z(n35957) );
  NANDN U36826 ( .A(n35901), .B(n42093), .Z(n35903) );
  XOR U36827 ( .A(n42134), .B(a[872]), .Z(n35942) );
  NANDN U36828 ( .A(n35942), .B(n42095), .Z(n35902) );
  NAND U36829 ( .A(n35903), .B(n35902), .Z(n35955) );
  NANDN U36830 ( .A(n35904), .B(n42231), .Z(n35906) );
  XOR U36831 ( .A(n234), .B(a[868]), .Z(n35945) );
  NANDN U36832 ( .A(n35945), .B(n42234), .Z(n35905) );
  AND U36833 ( .A(n35906), .B(n35905), .Z(n35954) );
  XNOR U36834 ( .A(n35955), .B(n35954), .Z(n35956) );
  XNOR U36835 ( .A(n35957), .B(n35956), .Z(n35961) );
  NANDN U36836 ( .A(n35908), .B(n35907), .Z(n35912) );
  NAND U36837 ( .A(n35910), .B(n35909), .Z(n35911) );
  AND U36838 ( .A(n35912), .B(n35911), .Z(n35960) );
  XOR U36839 ( .A(n35961), .B(n35960), .Z(n35962) );
  NANDN U36840 ( .A(n35914), .B(n35913), .Z(n35918) );
  NANDN U36841 ( .A(n35916), .B(n35915), .Z(n35917) );
  NAND U36842 ( .A(n35918), .B(n35917), .Z(n35963) );
  XOR U36843 ( .A(n35962), .B(n35963), .Z(n35930) );
  OR U36844 ( .A(n35920), .B(n35919), .Z(n35924) );
  NANDN U36845 ( .A(n35922), .B(n35921), .Z(n35923) );
  NAND U36846 ( .A(n35924), .B(n35923), .Z(n35931) );
  XNOR U36847 ( .A(n35930), .B(n35931), .Z(n35932) );
  XNOR U36848 ( .A(n35933), .B(n35932), .Z(n35966) );
  XNOR U36849 ( .A(n35966), .B(sreg[1890]), .Z(n35968) );
  NAND U36850 ( .A(n35925), .B(sreg[1889]), .Z(n35929) );
  OR U36851 ( .A(n35927), .B(n35926), .Z(n35928) );
  AND U36852 ( .A(n35929), .B(n35928), .Z(n35967) );
  XOR U36853 ( .A(n35968), .B(n35967), .Z(c[1890]) );
  NANDN U36854 ( .A(n35931), .B(n35930), .Z(n35935) );
  NAND U36855 ( .A(n35933), .B(n35932), .Z(n35934) );
  NAND U36856 ( .A(n35935), .B(n35934), .Z(n35974) );
  NAND U36857 ( .A(b[0]), .B(a[875]), .Z(n35936) );
  XNOR U36858 ( .A(b[1]), .B(n35936), .Z(n35938) );
  NAND U36859 ( .A(n140), .B(a[874]), .Z(n35937) );
  AND U36860 ( .A(n35938), .B(n35937), .Z(n35991) );
  XOR U36861 ( .A(a[871]), .B(n42197), .Z(n35980) );
  NANDN U36862 ( .A(n35980), .B(n42173), .Z(n35941) );
  NANDN U36863 ( .A(n35939), .B(n42172), .Z(n35940) );
  NAND U36864 ( .A(n35941), .B(n35940), .Z(n35989) );
  NAND U36865 ( .A(b[7]), .B(a[867]), .Z(n35990) );
  XNOR U36866 ( .A(n35989), .B(n35990), .Z(n35992) );
  XOR U36867 ( .A(n35991), .B(n35992), .Z(n35998) );
  NANDN U36868 ( .A(n35942), .B(n42093), .Z(n35944) );
  XOR U36869 ( .A(n42134), .B(a[873]), .Z(n35983) );
  NANDN U36870 ( .A(n35983), .B(n42095), .Z(n35943) );
  NAND U36871 ( .A(n35944), .B(n35943), .Z(n35996) );
  NANDN U36872 ( .A(n35945), .B(n42231), .Z(n35947) );
  XOR U36873 ( .A(n234), .B(a[869]), .Z(n35986) );
  NANDN U36874 ( .A(n35986), .B(n42234), .Z(n35946) );
  AND U36875 ( .A(n35947), .B(n35946), .Z(n35995) );
  XNOR U36876 ( .A(n35996), .B(n35995), .Z(n35997) );
  XNOR U36877 ( .A(n35998), .B(n35997), .Z(n36002) );
  NANDN U36878 ( .A(n35949), .B(n35948), .Z(n35953) );
  NAND U36879 ( .A(n35951), .B(n35950), .Z(n35952) );
  AND U36880 ( .A(n35953), .B(n35952), .Z(n36001) );
  XOR U36881 ( .A(n36002), .B(n36001), .Z(n36003) );
  NANDN U36882 ( .A(n35955), .B(n35954), .Z(n35959) );
  NANDN U36883 ( .A(n35957), .B(n35956), .Z(n35958) );
  NAND U36884 ( .A(n35959), .B(n35958), .Z(n36004) );
  XOR U36885 ( .A(n36003), .B(n36004), .Z(n35971) );
  OR U36886 ( .A(n35961), .B(n35960), .Z(n35965) );
  NANDN U36887 ( .A(n35963), .B(n35962), .Z(n35964) );
  NAND U36888 ( .A(n35965), .B(n35964), .Z(n35972) );
  XNOR U36889 ( .A(n35971), .B(n35972), .Z(n35973) );
  XNOR U36890 ( .A(n35974), .B(n35973), .Z(n36007) );
  XNOR U36891 ( .A(n36007), .B(sreg[1891]), .Z(n36009) );
  NAND U36892 ( .A(n35966), .B(sreg[1890]), .Z(n35970) );
  OR U36893 ( .A(n35968), .B(n35967), .Z(n35969) );
  AND U36894 ( .A(n35970), .B(n35969), .Z(n36008) );
  XOR U36895 ( .A(n36009), .B(n36008), .Z(c[1891]) );
  NANDN U36896 ( .A(n35972), .B(n35971), .Z(n35976) );
  NAND U36897 ( .A(n35974), .B(n35973), .Z(n35975) );
  NAND U36898 ( .A(n35976), .B(n35975), .Z(n36015) );
  NAND U36899 ( .A(b[0]), .B(a[876]), .Z(n35977) );
  XNOR U36900 ( .A(b[1]), .B(n35977), .Z(n35979) );
  NAND U36901 ( .A(n140), .B(a[875]), .Z(n35978) );
  AND U36902 ( .A(n35979), .B(n35978), .Z(n36032) );
  XOR U36903 ( .A(a[872]), .B(n42197), .Z(n36021) );
  NANDN U36904 ( .A(n36021), .B(n42173), .Z(n35982) );
  NANDN U36905 ( .A(n35980), .B(n42172), .Z(n35981) );
  NAND U36906 ( .A(n35982), .B(n35981), .Z(n36030) );
  NAND U36907 ( .A(b[7]), .B(a[868]), .Z(n36031) );
  XNOR U36908 ( .A(n36030), .B(n36031), .Z(n36033) );
  XOR U36909 ( .A(n36032), .B(n36033), .Z(n36039) );
  NANDN U36910 ( .A(n35983), .B(n42093), .Z(n35985) );
  XOR U36911 ( .A(n42134), .B(a[874]), .Z(n36024) );
  NANDN U36912 ( .A(n36024), .B(n42095), .Z(n35984) );
  NAND U36913 ( .A(n35985), .B(n35984), .Z(n36037) );
  NANDN U36914 ( .A(n35986), .B(n42231), .Z(n35988) );
  XOR U36915 ( .A(n234), .B(a[870]), .Z(n36027) );
  NANDN U36916 ( .A(n36027), .B(n42234), .Z(n35987) );
  AND U36917 ( .A(n35988), .B(n35987), .Z(n36036) );
  XNOR U36918 ( .A(n36037), .B(n36036), .Z(n36038) );
  XNOR U36919 ( .A(n36039), .B(n36038), .Z(n36043) );
  NANDN U36920 ( .A(n35990), .B(n35989), .Z(n35994) );
  NAND U36921 ( .A(n35992), .B(n35991), .Z(n35993) );
  AND U36922 ( .A(n35994), .B(n35993), .Z(n36042) );
  XOR U36923 ( .A(n36043), .B(n36042), .Z(n36044) );
  NANDN U36924 ( .A(n35996), .B(n35995), .Z(n36000) );
  NANDN U36925 ( .A(n35998), .B(n35997), .Z(n35999) );
  NAND U36926 ( .A(n36000), .B(n35999), .Z(n36045) );
  XOR U36927 ( .A(n36044), .B(n36045), .Z(n36012) );
  OR U36928 ( .A(n36002), .B(n36001), .Z(n36006) );
  NANDN U36929 ( .A(n36004), .B(n36003), .Z(n36005) );
  NAND U36930 ( .A(n36006), .B(n36005), .Z(n36013) );
  XNOR U36931 ( .A(n36012), .B(n36013), .Z(n36014) );
  XNOR U36932 ( .A(n36015), .B(n36014), .Z(n36048) );
  XNOR U36933 ( .A(n36048), .B(sreg[1892]), .Z(n36050) );
  NAND U36934 ( .A(n36007), .B(sreg[1891]), .Z(n36011) );
  OR U36935 ( .A(n36009), .B(n36008), .Z(n36010) );
  AND U36936 ( .A(n36011), .B(n36010), .Z(n36049) );
  XOR U36937 ( .A(n36050), .B(n36049), .Z(c[1892]) );
  NANDN U36938 ( .A(n36013), .B(n36012), .Z(n36017) );
  NAND U36939 ( .A(n36015), .B(n36014), .Z(n36016) );
  NAND U36940 ( .A(n36017), .B(n36016), .Z(n36056) );
  NAND U36941 ( .A(b[0]), .B(a[877]), .Z(n36018) );
  XNOR U36942 ( .A(b[1]), .B(n36018), .Z(n36020) );
  NAND U36943 ( .A(n140), .B(a[876]), .Z(n36019) );
  AND U36944 ( .A(n36020), .B(n36019), .Z(n36073) );
  XOR U36945 ( .A(a[873]), .B(n42197), .Z(n36062) );
  NANDN U36946 ( .A(n36062), .B(n42173), .Z(n36023) );
  NANDN U36947 ( .A(n36021), .B(n42172), .Z(n36022) );
  NAND U36948 ( .A(n36023), .B(n36022), .Z(n36071) );
  NAND U36949 ( .A(b[7]), .B(a[869]), .Z(n36072) );
  XNOR U36950 ( .A(n36071), .B(n36072), .Z(n36074) );
  XOR U36951 ( .A(n36073), .B(n36074), .Z(n36080) );
  NANDN U36952 ( .A(n36024), .B(n42093), .Z(n36026) );
  XOR U36953 ( .A(n42134), .B(a[875]), .Z(n36065) );
  NANDN U36954 ( .A(n36065), .B(n42095), .Z(n36025) );
  NAND U36955 ( .A(n36026), .B(n36025), .Z(n36078) );
  NANDN U36956 ( .A(n36027), .B(n42231), .Z(n36029) );
  XOR U36957 ( .A(n234), .B(a[871]), .Z(n36068) );
  NANDN U36958 ( .A(n36068), .B(n42234), .Z(n36028) );
  AND U36959 ( .A(n36029), .B(n36028), .Z(n36077) );
  XNOR U36960 ( .A(n36078), .B(n36077), .Z(n36079) );
  XNOR U36961 ( .A(n36080), .B(n36079), .Z(n36084) );
  NANDN U36962 ( .A(n36031), .B(n36030), .Z(n36035) );
  NAND U36963 ( .A(n36033), .B(n36032), .Z(n36034) );
  AND U36964 ( .A(n36035), .B(n36034), .Z(n36083) );
  XOR U36965 ( .A(n36084), .B(n36083), .Z(n36085) );
  NANDN U36966 ( .A(n36037), .B(n36036), .Z(n36041) );
  NANDN U36967 ( .A(n36039), .B(n36038), .Z(n36040) );
  NAND U36968 ( .A(n36041), .B(n36040), .Z(n36086) );
  XOR U36969 ( .A(n36085), .B(n36086), .Z(n36053) );
  OR U36970 ( .A(n36043), .B(n36042), .Z(n36047) );
  NANDN U36971 ( .A(n36045), .B(n36044), .Z(n36046) );
  NAND U36972 ( .A(n36047), .B(n36046), .Z(n36054) );
  XNOR U36973 ( .A(n36053), .B(n36054), .Z(n36055) );
  XNOR U36974 ( .A(n36056), .B(n36055), .Z(n36089) );
  XNOR U36975 ( .A(n36089), .B(sreg[1893]), .Z(n36091) );
  NAND U36976 ( .A(n36048), .B(sreg[1892]), .Z(n36052) );
  OR U36977 ( .A(n36050), .B(n36049), .Z(n36051) );
  AND U36978 ( .A(n36052), .B(n36051), .Z(n36090) );
  XOR U36979 ( .A(n36091), .B(n36090), .Z(c[1893]) );
  NANDN U36980 ( .A(n36054), .B(n36053), .Z(n36058) );
  NAND U36981 ( .A(n36056), .B(n36055), .Z(n36057) );
  NAND U36982 ( .A(n36058), .B(n36057), .Z(n36097) );
  NAND U36983 ( .A(b[0]), .B(a[878]), .Z(n36059) );
  XNOR U36984 ( .A(b[1]), .B(n36059), .Z(n36061) );
  NAND U36985 ( .A(n140), .B(a[877]), .Z(n36060) );
  AND U36986 ( .A(n36061), .B(n36060), .Z(n36114) );
  XOR U36987 ( .A(a[874]), .B(n42197), .Z(n36103) );
  NANDN U36988 ( .A(n36103), .B(n42173), .Z(n36064) );
  NANDN U36989 ( .A(n36062), .B(n42172), .Z(n36063) );
  NAND U36990 ( .A(n36064), .B(n36063), .Z(n36112) );
  NAND U36991 ( .A(b[7]), .B(a[870]), .Z(n36113) );
  XNOR U36992 ( .A(n36112), .B(n36113), .Z(n36115) );
  XOR U36993 ( .A(n36114), .B(n36115), .Z(n36121) );
  NANDN U36994 ( .A(n36065), .B(n42093), .Z(n36067) );
  XOR U36995 ( .A(n42134), .B(a[876]), .Z(n36106) );
  NANDN U36996 ( .A(n36106), .B(n42095), .Z(n36066) );
  NAND U36997 ( .A(n36067), .B(n36066), .Z(n36119) );
  NANDN U36998 ( .A(n36068), .B(n42231), .Z(n36070) );
  XOR U36999 ( .A(n234), .B(a[872]), .Z(n36109) );
  NANDN U37000 ( .A(n36109), .B(n42234), .Z(n36069) );
  AND U37001 ( .A(n36070), .B(n36069), .Z(n36118) );
  XNOR U37002 ( .A(n36119), .B(n36118), .Z(n36120) );
  XNOR U37003 ( .A(n36121), .B(n36120), .Z(n36125) );
  NANDN U37004 ( .A(n36072), .B(n36071), .Z(n36076) );
  NAND U37005 ( .A(n36074), .B(n36073), .Z(n36075) );
  AND U37006 ( .A(n36076), .B(n36075), .Z(n36124) );
  XOR U37007 ( .A(n36125), .B(n36124), .Z(n36126) );
  NANDN U37008 ( .A(n36078), .B(n36077), .Z(n36082) );
  NANDN U37009 ( .A(n36080), .B(n36079), .Z(n36081) );
  NAND U37010 ( .A(n36082), .B(n36081), .Z(n36127) );
  XOR U37011 ( .A(n36126), .B(n36127), .Z(n36094) );
  OR U37012 ( .A(n36084), .B(n36083), .Z(n36088) );
  NANDN U37013 ( .A(n36086), .B(n36085), .Z(n36087) );
  NAND U37014 ( .A(n36088), .B(n36087), .Z(n36095) );
  XNOR U37015 ( .A(n36094), .B(n36095), .Z(n36096) );
  XNOR U37016 ( .A(n36097), .B(n36096), .Z(n36130) );
  XNOR U37017 ( .A(n36130), .B(sreg[1894]), .Z(n36132) );
  NAND U37018 ( .A(n36089), .B(sreg[1893]), .Z(n36093) );
  OR U37019 ( .A(n36091), .B(n36090), .Z(n36092) );
  AND U37020 ( .A(n36093), .B(n36092), .Z(n36131) );
  XOR U37021 ( .A(n36132), .B(n36131), .Z(c[1894]) );
  NANDN U37022 ( .A(n36095), .B(n36094), .Z(n36099) );
  NAND U37023 ( .A(n36097), .B(n36096), .Z(n36098) );
  NAND U37024 ( .A(n36099), .B(n36098), .Z(n36138) );
  NAND U37025 ( .A(b[0]), .B(a[879]), .Z(n36100) );
  XNOR U37026 ( .A(b[1]), .B(n36100), .Z(n36102) );
  NAND U37027 ( .A(n140), .B(a[878]), .Z(n36101) );
  AND U37028 ( .A(n36102), .B(n36101), .Z(n36155) );
  XOR U37029 ( .A(a[875]), .B(n42197), .Z(n36144) );
  NANDN U37030 ( .A(n36144), .B(n42173), .Z(n36105) );
  NANDN U37031 ( .A(n36103), .B(n42172), .Z(n36104) );
  NAND U37032 ( .A(n36105), .B(n36104), .Z(n36153) );
  NAND U37033 ( .A(b[7]), .B(a[871]), .Z(n36154) );
  XNOR U37034 ( .A(n36153), .B(n36154), .Z(n36156) );
  XOR U37035 ( .A(n36155), .B(n36156), .Z(n36162) );
  NANDN U37036 ( .A(n36106), .B(n42093), .Z(n36108) );
  XOR U37037 ( .A(n42134), .B(a[877]), .Z(n36147) );
  NANDN U37038 ( .A(n36147), .B(n42095), .Z(n36107) );
  NAND U37039 ( .A(n36108), .B(n36107), .Z(n36160) );
  NANDN U37040 ( .A(n36109), .B(n42231), .Z(n36111) );
  XOR U37041 ( .A(n234), .B(a[873]), .Z(n36150) );
  NANDN U37042 ( .A(n36150), .B(n42234), .Z(n36110) );
  AND U37043 ( .A(n36111), .B(n36110), .Z(n36159) );
  XNOR U37044 ( .A(n36160), .B(n36159), .Z(n36161) );
  XNOR U37045 ( .A(n36162), .B(n36161), .Z(n36166) );
  NANDN U37046 ( .A(n36113), .B(n36112), .Z(n36117) );
  NAND U37047 ( .A(n36115), .B(n36114), .Z(n36116) );
  AND U37048 ( .A(n36117), .B(n36116), .Z(n36165) );
  XOR U37049 ( .A(n36166), .B(n36165), .Z(n36167) );
  NANDN U37050 ( .A(n36119), .B(n36118), .Z(n36123) );
  NANDN U37051 ( .A(n36121), .B(n36120), .Z(n36122) );
  NAND U37052 ( .A(n36123), .B(n36122), .Z(n36168) );
  XOR U37053 ( .A(n36167), .B(n36168), .Z(n36135) );
  OR U37054 ( .A(n36125), .B(n36124), .Z(n36129) );
  NANDN U37055 ( .A(n36127), .B(n36126), .Z(n36128) );
  NAND U37056 ( .A(n36129), .B(n36128), .Z(n36136) );
  XNOR U37057 ( .A(n36135), .B(n36136), .Z(n36137) );
  XNOR U37058 ( .A(n36138), .B(n36137), .Z(n36171) );
  XNOR U37059 ( .A(n36171), .B(sreg[1895]), .Z(n36173) );
  NAND U37060 ( .A(n36130), .B(sreg[1894]), .Z(n36134) );
  OR U37061 ( .A(n36132), .B(n36131), .Z(n36133) );
  AND U37062 ( .A(n36134), .B(n36133), .Z(n36172) );
  XOR U37063 ( .A(n36173), .B(n36172), .Z(c[1895]) );
  NANDN U37064 ( .A(n36136), .B(n36135), .Z(n36140) );
  NAND U37065 ( .A(n36138), .B(n36137), .Z(n36139) );
  NAND U37066 ( .A(n36140), .B(n36139), .Z(n36179) );
  NAND U37067 ( .A(b[0]), .B(a[880]), .Z(n36141) );
  XNOR U37068 ( .A(b[1]), .B(n36141), .Z(n36143) );
  NAND U37069 ( .A(n140), .B(a[879]), .Z(n36142) );
  AND U37070 ( .A(n36143), .B(n36142), .Z(n36196) );
  XOR U37071 ( .A(a[876]), .B(n42197), .Z(n36185) );
  NANDN U37072 ( .A(n36185), .B(n42173), .Z(n36146) );
  NANDN U37073 ( .A(n36144), .B(n42172), .Z(n36145) );
  NAND U37074 ( .A(n36146), .B(n36145), .Z(n36194) );
  NAND U37075 ( .A(b[7]), .B(a[872]), .Z(n36195) );
  XNOR U37076 ( .A(n36194), .B(n36195), .Z(n36197) );
  XOR U37077 ( .A(n36196), .B(n36197), .Z(n36203) );
  NANDN U37078 ( .A(n36147), .B(n42093), .Z(n36149) );
  XOR U37079 ( .A(n42134), .B(a[878]), .Z(n36188) );
  NANDN U37080 ( .A(n36188), .B(n42095), .Z(n36148) );
  NAND U37081 ( .A(n36149), .B(n36148), .Z(n36201) );
  NANDN U37082 ( .A(n36150), .B(n42231), .Z(n36152) );
  XOR U37083 ( .A(n234), .B(a[874]), .Z(n36191) );
  NANDN U37084 ( .A(n36191), .B(n42234), .Z(n36151) );
  AND U37085 ( .A(n36152), .B(n36151), .Z(n36200) );
  XNOR U37086 ( .A(n36201), .B(n36200), .Z(n36202) );
  XNOR U37087 ( .A(n36203), .B(n36202), .Z(n36207) );
  NANDN U37088 ( .A(n36154), .B(n36153), .Z(n36158) );
  NAND U37089 ( .A(n36156), .B(n36155), .Z(n36157) );
  AND U37090 ( .A(n36158), .B(n36157), .Z(n36206) );
  XOR U37091 ( .A(n36207), .B(n36206), .Z(n36208) );
  NANDN U37092 ( .A(n36160), .B(n36159), .Z(n36164) );
  NANDN U37093 ( .A(n36162), .B(n36161), .Z(n36163) );
  NAND U37094 ( .A(n36164), .B(n36163), .Z(n36209) );
  XOR U37095 ( .A(n36208), .B(n36209), .Z(n36176) );
  OR U37096 ( .A(n36166), .B(n36165), .Z(n36170) );
  NANDN U37097 ( .A(n36168), .B(n36167), .Z(n36169) );
  NAND U37098 ( .A(n36170), .B(n36169), .Z(n36177) );
  XNOR U37099 ( .A(n36176), .B(n36177), .Z(n36178) );
  XNOR U37100 ( .A(n36179), .B(n36178), .Z(n36212) );
  XNOR U37101 ( .A(n36212), .B(sreg[1896]), .Z(n36214) );
  NAND U37102 ( .A(n36171), .B(sreg[1895]), .Z(n36175) );
  OR U37103 ( .A(n36173), .B(n36172), .Z(n36174) );
  AND U37104 ( .A(n36175), .B(n36174), .Z(n36213) );
  XOR U37105 ( .A(n36214), .B(n36213), .Z(c[1896]) );
  NANDN U37106 ( .A(n36177), .B(n36176), .Z(n36181) );
  NAND U37107 ( .A(n36179), .B(n36178), .Z(n36180) );
  NAND U37108 ( .A(n36181), .B(n36180), .Z(n36220) );
  NAND U37109 ( .A(b[0]), .B(a[881]), .Z(n36182) );
  XNOR U37110 ( .A(b[1]), .B(n36182), .Z(n36184) );
  NAND U37111 ( .A(n140), .B(a[880]), .Z(n36183) );
  AND U37112 ( .A(n36184), .B(n36183), .Z(n36237) );
  XOR U37113 ( .A(a[877]), .B(n42197), .Z(n36226) );
  NANDN U37114 ( .A(n36226), .B(n42173), .Z(n36187) );
  NANDN U37115 ( .A(n36185), .B(n42172), .Z(n36186) );
  NAND U37116 ( .A(n36187), .B(n36186), .Z(n36235) );
  NAND U37117 ( .A(b[7]), .B(a[873]), .Z(n36236) );
  XNOR U37118 ( .A(n36235), .B(n36236), .Z(n36238) );
  XOR U37119 ( .A(n36237), .B(n36238), .Z(n36244) );
  NANDN U37120 ( .A(n36188), .B(n42093), .Z(n36190) );
  XOR U37121 ( .A(n42134), .B(a[879]), .Z(n36229) );
  NANDN U37122 ( .A(n36229), .B(n42095), .Z(n36189) );
  NAND U37123 ( .A(n36190), .B(n36189), .Z(n36242) );
  NANDN U37124 ( .A(n36191), .B(n42231), .Z(n36193) );
  XOR U37125 ( .A(n235), .B(a[875]), .Z(n36232) );
  NANDN U37126 ( .A(n36232), .B(n42234), .Z(n36192) );
  AND U37127 ( .A(n36193), .B(n36192), .Z(n36241) );
  XNOR U37128 ( .A(n36242), .B(n36241), .Z(n36243) );
  XNOR U37129 ( .A(n36244), .B(n36243), .Z(n36248) );
  NANDN U37130 ( .A(n36195), .B(n36194), .Z(n36199) );
  NAND U37131 ( .A(n36197), .B(n36196), .Z(n36198) );
  AND U37132 ( .A(n36199), .B(n36198), .Z(n36247) );
  XOR U37133 ( .A(n36248), .B(n36247), .Z(n36249) );
  NANDN U37134 ( .A(n36201), .B(n36200), .Z(n36205) );
  NANDN U37135 ( .A(n36203), .B(n36202), .Z(n36204) );
  NAND U37136 ( .A(n36205), .B(n36204), .Z(n36250) );
  XOR U37137 ( .A(n36249), .B(n36250), .Z(n36217) );
  OR U37138 ( .A(n36207), .B(n36206), .Z(n36211) );
  NANDN U37139 ( .A(n36209), .B(n36208), .Z(n36210) );
  NAND U37140 ( .A(n36211), .B(n36210), .Z(n36218) );
  XNOR U37141 ( .A(n36217), .B(n36218), .Z(n36219) );
  XNOR U37142 ( .A(n36220), .B(n36219), .Z(n36253) );
  XNOR U37143 ( .A(n36253), .B(sreg[1897]), .Z(n36255) );
  NAND U37144 ( .A(n36212), .B(sreg[1896]), .Z(n36216) );
  OR U37145 ( .A(n36214), .B(n36213), .Z(n36215) );
  AND U37146 ( .A(n36216), .B(n36215), .Z(n36254) );
  XOR U37147 ( .A(n36255), .B(n36254), .Z(c[1897]) );
  NANDN U37148 ( .A(n36218), .B(n36217), .Z(n36222) );
  NAND U37149 ( .A(n36220), .B(n36219), .Z(n36221) );
  NAND U37150 ( .A(n36222), .B(n36221), .Z(n36261) );
  NAND U37151 ( .A(b[0]), .B(a[882]), .Z(n36223) );
  XNOR U37152 ( .A(b[1]), .B(n36223), .Z(n36225) );
  NAND U37153 ( .A(n141), .B(a[881]), .Z(n36224) );
  AND U37154 ( .A(n36225), .B(n36224), .Z(n36278) );
  XOR U37155 ( .A(a[878]), .B(n42197), .Z(n36267) );
  NANDN U37156 ( .A(n36267), .B(n42173), .Z(n36228) );
  NANDN U37157 ( .A(n36226), .B(n42172), .Z(n36227) );
  NAND U37158 ( .A(n36228), .B(n36227), .Z(n36276) );
  NAND U37159 ( .A(b[7]), .B(a[874]), .Z(n36277) );
  XNOR U37160 ( .A(n36276), .B(n36277), .Z(n36279) );
  XOR U37161 ( .A(n36278), .B(n36279), .Z(n36285) );
  NANDN U37162 ( .A(n36229), .B(n42093), .Z(n36231) );
  XOR U37163 ( .A(n42134), .B(a[880]), .Z(n36270) );
  NANDN U37164 ( .A(n36270), .B(n42095), .Z(n36230) );
  NAND U37165 ( .A(n36231), .B(n36230), .Z(n36283) );
  NANDN U37166 ( .A(n36232), .B(n42231), .Z(n36234) );
  XOR U37167 ( .A(n235), .B(a[876]), .Z(n36273) );
  NANDN U37168 ( .A(n36273), .B(n42234), .Z(n36233) );
  AND U37169 ( .A(n36234), .B(n36233), .Z(n36282) );
  XNOR U37170 ( .A(n36283), .B(n36282), .Z(n36284) );
  XNOR U37171 ( .A(n36285), .B(n36284), .Z(n36289) );
  NANDN U37172 ( .A(n36236), .B(n36235), .Z(n36240) );
  NAND U37173 ( .A(n36238), .B(n36237), .Z(n36239) );
  AND U37174 ( .A(n36240), .B(n36239), .Z(n36288) );
  XOR U37175 ( .A(n36289), .B(n36288), .Z(n36290) );
  NANDN U37176 ( .A(n36242), .B(n36241), .Z(n36246) );
  NANDN U37177 ( .A(n36244), .B(n36243), .Z(n36245) );
  NAND U37178 ( .A(n36246), .B(n36245), .Z(n36291) );
  XOR U37179 ( .A(n36290), .B(n36291), .Z(n36258) );
  OR U37180 ( .A(n36248), .B(n36247), .Z(n36252) );
  NANDN U37181 ( .A(n36250), .B(n36249), .Z(n36251) );
  NAND U37182 ( .A(n36252), .B(n36251), .Z(n36259) );
  XNOR U37183 ( .A(n36258), .B(n36259), .Z(n36260) );
  XNOR U37184 ( .A(n36261), .B(n36260), .Z(n36294) );
  XNOR U37185 ( .A(n36294), .B(sreg[1898]), .Z(n36296) );
  NAND U37186 ( .A(n36253), .B(sreg[1897]), .Z(n36257) );
  OR U37187 ( .A(n36255), .B(n36254), .Z(n36256) );
  AND U37188 ( .A(n36257), .B(n36256), .Z(n36295) );
  XOR U37189 ( .A(n36296), .B(n36295), .Z(c[1898]) );
  NANDN U37190 ( .A(n36259), .B(n36258), .Z(n36263) );
  NAND U37191 ( .A(n36261), .B(n36260), .Z(n36262) );
  NAND U37192 ( .A(n36263), .B(n36262), .Z(n36302) );
  NAND U37193 ( .A(b[0]), .B(a[883]), .Z(n36264) );
  XNOR U37194 ( .A(b[1]), .B(n36264), .Z(n36266) );
  NAND U37195 ( .A(n141), .B(a[882]), .Z(n36265) );
  AND U37196 ( .A(n36266), .B(n36265), .Z(n36319) );
  XOR U37197 ( .A(a[879]), .B(n42197), .Z(n36308) );
  NANDN U37198 ( .A(n36308), .B(n42173), .Z(n36269) );
  NANDN U37199 ( .A(n36267), .B(n42172), .Z(n36268) );
  NAND U37200 ( .A(n36269), .B(n36268), .Z(n36317) );
  NAND U37201 ( .A(b[7]), .B(a[875]), .Z(n36318) );
  XNOR U37202 ( .A(n36317), .B(n36318), .Z(n36320) );
  XOR U37203 ( .A(n36319), .B(n36320), .Z(n36326) );
  NANDN U37204 ( .A(n36270), .B(n42093), .Z(n36272) );
  XOR U37205 ( .A(n42134), .B(a[881]), .Z(n36311) );
  NANDN U37206 ( .A(n36311), .B(n42095), .Z(n36271) );
  NAND U37207 ( .A(n36272), .B(n36271), .Z(n36324) );
  NANDN U37208 ( .A(n36273), .B(n42231), .Z(n36275) );
  XOR U37209 ( .A(n235), .B(a[877]), .Z(n36314) );
  NANDN U37210 ( .A(n36314), .B(n42234), .Z(n36274) );
  AND U37211 ( .A(n36275), .B(n36274), .Z(n36323) );
  XNOR U37212 ( .A(n36324), .B(n36323), .Z(n36325) );
  XNOR U37213 ( .A(n36326), .B(n36325), .Z(n36330) );
  NANDN U37214 ( .A(n36277), .B(n36276), .Z(n36281) );
  NAND U37215 ( .A(n36279), .B(n36278), .Z(n36280) );
  AND U37216 ( .A(n36281), .B(n36280), .Z(n36329) );
  XOR U37217 ( .A(n36330), .B(n36329), .Z(n36331) );
  NANDN U37218 ( .A(n36283), .B(n36282), .Z(n36287) );
  NANDN U37219 ( .A(n36285), .B(n36284), .Z(n36286) );
  NAND U37220 ( .A(n36287), .B(n36286), .Z(n36332) );
  XOR U37221 ( .A(n36331), .B(n36332), .Z(n36299) );
  OR U37222 ( .A(n36289), .B(n36288), .Z(n36293) );
  NANDN U37223 ( .A(n36291), .B(n36290), .Z(n36292) );
  NAND U37224 ( .A(n36293), .B(n36292), .Z(n36300) );
  XNOR U37225 ( .A(n36299), .B(n36300), .Z(n36301) );
  XNOR U37226 ( .A(n36302), .B(n36301), .Z(n36335) );
  XNOR U37227 ( .A(n36335), .B(sreg[1899]), .Z(n36337) );
  NAND U37228 ( .A(n36294), .B(sreg[1898]), .Z(n36298) );
  OR U37229 ( .A(n36296), .B(n36295), .Z(n36297) );
  AND U37230 ( .A(n36298), .B(n36297), .Z(n36336) );
  XOR U37231 ( .A(n36337), .B(n36336), .Z(c[1899]) );
  NANDN U37232 ( .A(n36300), .B(n36299), .Z(n36304) );
  NAND U37233 ( .A(n36302), .B(n36301), .Z(n36303) );
  NAND U37234 ( .A(n36304), .B(n36303), .Z(n36343) );
  NAND U37235 ( .A(b[0]), .B(a[884]), .Z(n36305) );
  XNOR U37236 ( .A(b[1]), .B(n36305), .Z(n36307) );
  NAND U37237 ( .A(n141), .B(a[883]), .Z(n36306) );
  AND U37238 ( .A(n36307), .B(n36306), .Z(n36360) );
  XOR U37239 ( .A(a[880]), .B(n42197), .Z(n36349) );
  NANDN U37240 ( .A(n36349), .B(n42173), .Z(n36310) );
  NANDN U37241 ( .A(n36308), .B(n42172), .Z(n36309) );
  NAND U37242 ( .A(n36310), .B(n36309), .Z(n36358) );
  NAND U37243 ( .A(b[7]), .B(a[876]), .Z(n36359) );
  XNOR U37244 ( .A(n36358), .B(n36359), .Z(n36361) );
  XOR U37245 ( .A(n36360), .B(n36361), .Z(n36367) );
  NANDN U37246 ( .A(n36311), .B(n42093), .Z(n36313) );
  XOR U37247 ( .A(n42134), .B(a[882]), .Z(n36352) );
  NANDN U37248 ( .A(n36352), .B(n42095), .Z(n36312) );
  NAND U37249 ( .A(n36313), .B(n36312), .Z(n36365) );
  NANDN U37250 ( .A(n36314), .B(n42231), .Z(n36316) );
  XOR U37251 ( .A(n235), .B(a[878]), .Z(n36355) );
  NANDN U37252 ( .A(n36355), .B(n42234), .Z(n36315) );
  AND U37253 ( .A(n36316), .B(n36315), .Z(n36364) );
  XNOR U37254 ( .A(n36365), .B(n36364), .Z(n36366) );
  XNOR U37255 ( .A(n36367), .B(n36366), .Z(n36371) );
  NANDN U37256 ( .A(n36318), .B(n36317), .Z(n36322) );
  NAND U37257 ( .A(n36320), .B(n36319), .Z(n36321) );
  AND U37258 ( .A(n36322), .B(n36321), .Z(n36370) );
  XOR U37259 ( .A(n36371), .B(n36370), .Z(n36372) );
  NANDN U37260 ( .A(n36324), .B(n36323), .Z(n36328) );
  NANDN U37261 ( .A(n36326), .B(n36325), .Z(n36327) );
  NAND U37262 ( .A(n36328), .B(n36327), .Z(n36373) );
  XOR U37263 ( .A(n36372), .B(n36373), .Z(n36340) );
  OR U37264 ( .A(n36330), .B(n36329), .Z(n36334) );
  NANDN U37265 ( .A(n36332), .B(n36331), .Z(n36333) );
  NAND U37266 ( .A(n36334), .B(n36333), .Z(n36341) );
  XNOR U37267 ( .A(n36340), .B(n36341), .Z(n36342) );
  XNOR U37268 ( .A(n36343), .B(n36342), .Z(n36376) );
  XNOR U37269 ( .A(n36376), .B(sreg[1900]), .Z(n36378) );
  NAND U37270 ( .A(n36335), .B(sreg[1899]), .Z(n36339) );
  OR U37271 ( .A(n36337), .B(n36336), .Z(n36338) );
  AND U37272 ( .A(n36339), .B(n36338), .Z(n36377) );
  XOR U37273 ( .A(n36378), .B(n36377), .Z(c[1900]) );
  NANDN U37274 ( .A(n36341), .B(n36340), .Z(n36345) );
  NAND U37275 ( .A(n36343), .B(n36342), .Z(n36344) );
  NAND U37276 ( .A(n36345), .B(n36344), .Z(n36384) );
  NAND U37277 ( .A(b[0]), .B(a[885]), .Z(n36346) );
  XNOR U37278 ( .A(b[1]), .B(n36346), .Z(n36348) );
  NAND U37279 ( .A(n141), .B(a[884]), .Z(n36347) );
  AND U37280 ( .A(n36348), .B(n36347), .Z(n36401) );
  XOR U37281 ( .A(a[881]), .B(n42197), .Z(n36390) );
  NANDN U37282 ( .A(n36390), .B(n42173), .Z(n36351) );
  NANDN U37283 ( .A(n36349), .B(n42172), .Z(n36350) );
  NAND U37284 ( .A(n36351), .B(n36350), .Z(n36399) );
  NAND U37285 ( .A(b[7]), .B(a[877]), .Z(n36400) );
  XNOR U37286 ( .A(n36399), .B(n36400), .Z(n36402) );
  XOR U37287 ( .A(n36401), .B(n36402), .Z(n36408) );
  NANDN U37288 ( .A(n36352), .B(n42093), .Z(n36354) );
  XOR U37289 ( .A(n42134), .B(a[883]), .Z(n36393) );
  NANDN U37290 ( .A(n36393), .B(n42095), .Z(n36353) );
  NAND U37291 ( .A(n36354), .B(n36353), .Z(n36406) );
  NANDN U37292 ( .A(n36355), .B(n42231), .Z(n36357) );
  XOR U37293 ( .A(n235), .B(a[879]), .Z(n36396) );
  NANDN U37294 ( .A(n36396), .B(n42234), .Z(n36356) );
  AND U37295 ( .A(n36357), .B(n36356), .Z(n36405) );
  XNOR U37296 ( .A(n36406), .B(n36405), .Z(n36407) );
  XNOR U37297 ( .A(n36408), .B(n36407), .Z(n36412) );
  NANDN U37298 ( .A(n36359), .B(n36358), .Z(n36363) );
  NAND U37299 ( .A(n36361), .B(n36360), .Z(n36362) );
  AND U37300 ( .A(n36363), .B(n36362), .Z(n36411) );
  XOR U37301 ( .A(n36412), .B(n36411), .Z(n36413) );
  NANDN U37302 ( .A(n36365), .B(n36364), .Z(n36369) );
  NANDN U37303 ( .A(n36367), .B(n36366), .Z(n36368) );
  NAND U37304 ( .A(n36369), .B(n36368), .Z(n36414) );
  XOR U37305 ( .A(n36413), .B(n36414), .Z(n36381) );
  OR U37306 ( .A(n36371), .B(n36370), .Z(n36375) );
  NANDN U37307 ( .A(n36373), .B(n36372), .Z(n36374) );
  NAND U37308 ( .A(n36375), .B(n36374), .Z(n36382) );
  XNOR U37309 ( .A(n36381), .B(n36382), .Z(n36383) );
  XNOR U37310 ( .A(n36384), .B(n36383), .Z(n36417) );
  XNOR U37311 ( .A(n36417), .B(sreg[1901]), .Z(n36419) );
  NAND U37312 ( .A(n36376), .B(sreg[1900]), .Z(n36380) );
  OR U37313 ( .A(n36378), .B(n36377), .Z(n36379) );
  AND U37314 ( .A(n36380), .B(n36379), .Z(n36418) );
  XOR U37315 ( .A(n36419), .B(n36418), .Z(c[1901]) );
  NANDN U37316 ( .A(n36382), .B(n36381), .Z(n36386) );
  NAND U37317 ( .A(n36384), .B(n36383), .Z(n36385) );
  NAND U37318 ( .A(n36386), .B(n36385), .Z(n36425) );
  NAND U37319 ( .A(b[0]), .B(a[886]), .Z(n36387) );
  XNOR U37320 ( .A(b[1]), .B(n36387), .Z(n36389) );
  NAND U37321 ( .A(n141), .B(a[885]), .Z(n36388) );
  AND U37322 ( .A(n36389), .B(n36388), .Z(n36442) );
  XOR U37323 ( .A(a[882]), .B(n42197), .Z(n36431) );
  NANDN U37324 ( .A(n36431), .B(n42173), .Z(n36392) );
  NANDN U37325 ( .A(n36390), .B(n42172), .Z(n36391) );
  NAND U37326 ( .A(n36392), .B(n36391), .Z(n36440) );
  NAND U37327 ( .A(b[7]), .B(a[878]), .Z(n36441) );
  XNOR U37328 ( .A(n36440), .B(n36441), .Z(n36443) );
  XOR U37329 ( .A(n36442), .B(n36443), .Z(n36449) );
  NANDN U37330 ( .A(n36393), .B(n42093), .Z(n36395) );
  XOR U37331 ( .A(n42134), .B(a[884]), .Z(n36434) );
  NANDN U37332 ( .A(n36434), .B(n42095), .Z(n36394) );
  NAND U37333 ( .A(n36395), .B(n36394), .Z(n36447) );
  NANDN U37334 ( .A(n36396), .B(n42231), .Z(n36398) );
  XOR U37335 ( .A(n235), .B(a[880]), .Z(n36437) );
  NANDN U37336 ( .A(n36437), .B(n42234), .Z(n36397) );
  AND U37337 ( .A(n36398), .B(n36397), .Z(n36446) );
  XNOR U37338 ( .A(n36447), .B(n36446), .Z(n36448) );
  XNOR U37339 ( .A(n36449), .B(n36448), .Z(n36453) );
  NANDN U37340 ( .A(n36400), .B(n36399), .Z(n36404) );
  NAND U37341 ( .A(n36402), .B(n36401), .Z(n36403) );
  AND U37342 ( .A(n36404), .B(n36403), .Z(n36452) );
  XOR U37343 ( .A(n36453), .B(n36452), .Z(n36454) );
  NANDN U37344 ( .A(n36406), .B(n36405), .Z(n36410) );
  NANDN U37345 ( .A(n36408), .B(n36407), .Z(n36409) );
  NAND U37346 ( .A(n36410), .B(n36409), .Z(n36455) );
  XOR U37347 ( .A(n36454), .B(n36455), .Z(n36422) );
  OR U37348 ( .A(n36412), .B(n36411), .Z(n36416) );
  NANDN U37349 ( .A(n36414), .B(n36413), .Z(n36415) );
  NAND U37350 ( .A(n36416), .B(n36415), .Z(n36423) );
  XNOR U37351 ( .A(n36422), .B(n36423), .Z(n36424) );
  XNOR U37352 ( .A(n36425), .B(n36424), .Z(n36458) );
  XNOR U37353 ( .A(n36458), .B(sreg[1902]), .Z(n36460) );
  NAND U37354 ( .A(n36417), .B(sreg[1901]), .Z(n36421) );
  OR U37355 ( .A(n36419), .B(n36418), .Z(n36420) );
  AND U37356 ( .A(n36421), .B(n36420), .Z(n36459) );
  XOR U37357 ( .A(n36460), .B(n36459), .Z(c[1902]) );
  NANDN U37358 ( .A(n36423), .B(n36422), .Z(n36427) );
  NAND U37359 ( .A(n36425), .B(n36424), .Z(n36426) );
  NAND U37360 ( .A(n36427), .B(n36426), .Z(n36466) );
  NAND U37361 ( .A(b[0]), .B(a[887]), .Z(n36428) );
  XNOR U37362 ( .A(b[1]), .B(n36428), .Z(n36430) );
  NAND U37363 ( .A(n141), .B(a[886]), .Z(n36429) );
  AND U37364 ( .A(n36430), .B(n36429), .Z(n36483) );
  XOR U37365 ( .A(a[883]), .B(n42197), .Z(n36472) );
  NANDN U37366 ( .A(n36472), .B(n42173), .Z(n36433) );
  NANDN U37367 ( .A(n36431), .B(n42172), .Z(n36432) );
  NAND U37368 ( .A(n36433), .B(n36432), .Z(n36481) );
  NAND U37369 ( .A(b[7]), .B(a[879]), .Z(n36482) );
  XNOR U37370 ( .A(n36481), .B(n36482), .Z(n36484) );
  XOR U37371 ( .A(n36483), .B(n36484), .Z(n36490) );
  NANDN U37372 ( .A(n36434), .B(n42093), .Z(n36436) );
  XOR U37373 ( .A(n42134), .B(a[885]), .Z(n36475) );
  NANDN U37374 ( .A(n36475), .B(n42095), .Z(n36435) );
  NAND U37375 ( .A(n36436), .B(n36435), .Z(n36488) );
  NANDN U37376 ( .A(n36437), .B(n42231), .Z(n36439) );
  XOR U37377 ( .A(n235), .B(a[881]), .Z(n36478) );
  NANDN U37378 ( .A(n36478), .B(n42234), .Z(n36438) );
  AND U37379 ( .A(n36439), .B(n36438), .Z(n36487) );
  XNOR U37380 ( .A(n36488), .B(n36487), .Z(n36489) );
  XNOR U37381 ( .A(n36490), .B(n36489), .Z(n36494) );
  NANDN U37382 ( .A(n36441), .B(n36440), .Z(n36445) );
  NAND U37383 ( .A(n36443), .B(n36442), .Z(n36444) );
  AND U37384 ( .A(n36445), .B(n36444), .Z(n36493) );
  XOR U37385 ( .A(n36494), .B(n36493), .Z(n36495) );
  NANDN U37386 ( .A(n36447), .B(n36446), .Z(n36451) );
  NANDN U37387 ( .A(n36449), .B(n36448), .Z(n36450) );
  NAND U37388 ( .A(n36451), .B(n36450), .Z(n36496) );
  XOR U37389 ( .A(n36495), .B(n36496), .Z(n36463) );
  OR U37390 ( .A(n36453), .B(n36452), .Z(n36457) );
  NANDN U37391 ( .A(n36455), .B(n36454), .Z(n36456) );
  NAND U37392 ( .A(n36457), .B(n36456), .Z(n36464) );
  XNOR U37393 ( .A(n36463), .B(n36464), .Z(n36465) );
  XNOR U37394 ( .A(n36466), .B(n36465), .Z(n36499) );
  XNOR U37395 ( .A(n36499), .B(sreg[1903]), .Z(n36501) );
  NAND U37396 ( .A(n36458), .B(sreg[1902]), .Z(n36462) );
  OR U37397 ( .A(n36460), .B(n36459), .Z(n36461) );
  AND U37398 ( .A(n36462), .B(n36461), .Z(n36500) );
  XOR U37399 ( .A(n36501), .B(n36500), .Z(c[1903]) );
  NANDN U37400 ( .A(n36464), .B(n36463), .Z(n36468) );
  NAND U37401 ( .A(n36466), .B(n36465), .Z(n36467) );
  NAND U37402 ( .A(n36468), .B(n36467), .Z(n36507) );
  NAND U37403 ( .A(b[0]), .B(a[888]), .Z(n36469) );
  XNOR U37404 ( .A(b[1]), .B(n36469), .Z(n36471) );
  NAND U37405 ( .A(n141), .B(a[887]), .Z(n36470) );
  AND U37406 ( .A(n36471), .B(n36470), .Z(n36524) );
  XOR U37407 ( .A(a[884]), .B(n42197), .Z(n36513) );
  NANDN U37408 ( .A(n36513), .B(n42173), .Z(n36474) );
  NANDN U37409 ( .A(n36472), .B(n42172), .Z(n36473) );
  NAND U37410 ( .A(n36474), .B(n36473), .Z(n36522) );
  NAND U37411 ( .A(b[7]), .B(a[880]), .Z(n36523) );
  XNOR U37412 ( .A(n36522), .B(n36523), .Z(n36525) );
  XOR U37413 ( .A(n36524), .B(n36525), .Z(n36531) );
  NANDN U37414 ( .A(n36475), .B(n42093), .Z(n36477) );
  XOR U37415 ( .A(n42134), .B(a[886]), .Z(n36516) );
  NANDN U37416 ( .A(n36516), .B(n42095), .Z(n36476) );
  NAND U37417 ( .A(n36477), .B(n36476), .Z(n36529) );
  NANDN U37418 ( .A(n36478), .B(n42231), .Z(n36480) );
  XOR U37419 ( .A(n235), .B(a[882]), .Z(n36519) );
  NANDN U37420 ( .A(n36519), .B(n42234), .Z(n36479) );
  AND U37421 ( .A(n36480), .B(n36479), .Z(n36528) );
  XNOR U37422 ( .A(n36529), .B(n36528), .Z(n36530) );
  XNOR U37423 ( .A(n36531), .B(n36530), .Z(n36535) );
  NANDN U37424 ( .A(n36482), .B(n36481), .Z(n36486) );
  NAND U37425 ( .A(n36484), .B(n36483), .Z(n36485) );
  AND U37426 ( .A(n36486), .B(n36485), .Z(n36534) );
  XOR U37427 ( .A(n36535), .B(n36534), .Z(n36536) );
  NANDN U37428 ( .A(n36488), .B(n36487), .Z(n36492) );
  NANDN U37429 ( .A(n36490), .B(n36489), .Z(n36491) );
  NAND U37430 ( .A(n36492), .B(n36491), .Z(n36537) );
  XOR U37431 ( .A(n36536), .B(n36537), .Z(n36504) );
  OR U37432 ( .A(n36494), .B(n36493), .Z(n36498) );
  NANDN U37433 ( .A(n36496), .B(n36495), .Z(n36497) );
  NAND U37434 ( .A(n36498), .B(n36497), .Z(n36505) );
  XNOR U37435 ( .A(n36504), .B(n36505), .Z(n36506) );
  XNOR U37436 ( .A(n36507), .B(n36506), .Z(n36540) );
  XNOR U37437 ( .A(n36540), .B(sreg[1904]), .Z(n36542) );
  NAND U37438 ( .A(n36499), .B(sreg[1903]), .Z(n36503) );
  OR U37439 ( .A(n36501), .B(n36500), .Z(n36502) );
  AND U37440 ( .A(n36503), .B(n36502), .Z(n36541) );
  XOR U37441 ( .A(n36542), .B(n36541), .Z(c[1904]) );
  NANDN U37442 ( .A(n36505), .B(n36504), .Z(n36509) );
  NAND U37443 ( .A(n36507), .B(n36506), .Z(n36508) );
  NAND U37444 ( .A(n36509), .B(n36508), .Z(n36548) );
  NAND U37445 ( .A(b[0]), .B(a[889]), .Z(n36510) );
  XNOR U37446 ( .A(b[1]), .B(n36510), .Z(n36512) );
  NAND U37447 ( .A(n142), .B(a[888]), .Z(n36511) );
  AND U37448 ( .A(n36512), .B(n36511), .Z(n36565) );
  XOR U37449 ( .A(a[885]), .B(n42197), .Z(n36554) );
  NANDN U37450 ( .A(n36554), .B(n42173), .Z(n36515) );
  NANDN U37451 ( .A(n36513), .B(n42172), .Z(n36514) );
  NAND U37452 ( .A(n36515), .B(n36514), .Z(n36563) );
  NAND U37453 ( .A(b[7]), .B(a[881]), .Z(n36564) );
  XNOR U37454 ( .A(n36563), .B(n36564), .Z(n36566) );
  XOR U37455 ( .A(n36565), .B(n36566), .Z(n36572) );
  NANDN U37456 ( .A(n36516), .B(n42093), .Z(n36518) );
  XOR U37457 ( .A(n42134), .B(a[887]), .Z(n36557) );
  NANDN U37458 ( .A(n36557), .B(n42095), .Z(n36517) );
  NAND U37459 ( .A(n36518), .B(n36517), .Z(n36570) );
  NANDN U37460 ( .A(n36519), .B(n42231), .Z(n36521) );
  XOR U37461 ( .A(n235), .B(a[883]), .Z(n36560) );
  NANDN U37462 ( .A(n36560), .B(n42234), .Z(n36520) );
  AND U37463 ( .A(n36521), .B(n36520), .Z(n36569) );
  XNOR U37464 ( .A(n36570), .B(n36569), .Z(n36571) );
  XNOR U37465 ( .A(n36572), .B(n36571), .Z(n36576) );
  NANDN U37466 ( .A(n36523), .B(n36522), .Z(n36527) );
  NAND U37467 ( .A(n36525), .B(n36524), .Z(n36526) );
  AND U37468 ( .A(n36527), .B(n36526), .Z(n36575) );
  XOR U37469 ( .A(n36576), .B(n36575), .Z(n36577) );
  NANDN U37470 ( .A(n36529), .B(n36528), .Z(n36533) );
  NANDN U37471 ( .A(n36531), .B(n36530), .Z(n36532) );
  NAND U37472 ( .A(n36533), .B(n36532), .Z(n36578) );
  XOR U37473 ( .A(n36577), .B(n36578), .Z(n36545) );
  OR U37474 ( .A(n36535), .B(n36534), .Z(n36539) );
  NANDN U37475 ( .A(n36537), .B(n36536), .Z(n36538) );
  NAND U37476 ( .A(n36539), .B(n36538), .Z(n36546) );
  XNOR U37477 ( .A(n36545), .B(n36546), .Z(n36547) );
  XNOR U37478 ( .A(n36548), .B(n36547), .Z(n36581) );
  XNOR U37479 ( .A(n36581), .B(sreg[1905]), .Z(n36583) );
  NAND U37480 ( .A(n36540), .B(sreg[1904]), .Z(n36544) );
  OR U37481 ( .A(n36542), .B(n36541), .Z(n36543) );
  AND U37482 ( .A(n36544), .B(n36543), .Z(n36582) );
  XOR U37483 ( .A(n36583), .B(n36582), .Z(c[1905]) );
  NANDN U37484 ( .A(n36546), .B(n36545), .Z(n36550) );
  NAND U37485 ( .A(n36548), .B(n36547), .Z(n36549) );
  NAND U37486 ( .A(n36550), .B(n36549), .Z(n36589) );
  NAND U37487 ( .A(b[0]), .B(a[890]), .Z(n36551) );
  XNOR U37488 ( .A(b[1]), .B(n36551), .Z(n36553) );
  NAND U37489 ( .A(n142), .B(a[889]), .Z(n36552) );
  AND U37490 ( .A(n36553), .B(n36552), .Z(n36606) );
  XOR U37491 ( .A(a[886]), .B(n42197), .Z(n36595) );
  NANDN U37492 ( .A(n36595), .B(n42173), .Z(n36556) );
  NANDN U37493 ( .A(n36554), .B(n42172), .Z(n36555) );
  NAND U37494 ( .A(n36556), .B(n36555), .Z(n36604) );
  NAND U37495 ( .A(b[7]), .B(a[882]), .Z(n36605) );
  XNOR U37496 ( .A(n36604), .B(n36605), .Z(n36607) );
  XOR U37497 ( .A(n36606), .B(n36607), .Z(n36613) );
  NANDN U37498 ( .A(n36557), .B(n42093), .Z(n36559) );
  XOR U37499 ( .A(n42134), .B(a[888]), .Z(n36598) );
  NANDN U37500 ( .A(n36598), .B(n42095), .Z(n36558) );
  NAND U37501 ( .A(n36559), .B(n36558), .Z(n36611) );
  NANDN U37502 ( .A(n36560), .B(n42231), .Z(n36562) );
  XOR U37503 ( .A(n235), .B(a[884]), .Z(n36601) );
  NANDN U37504 ( .A(n36601), .B(n42234), .Z(n36561) );
  AND U37505 ( .A(n36562), .B(n36561), .Z(n36610) );
  XNOR U37506 ( .A(n36611), .B(n36610), .Z(n36612) );
  XNOR U37507 ( .A(n36613), .B(n36612), .Z(n36617) );
  NANDN U37508 ( .A(n36564), .B(n36563), .Z(n36568) );
  NAND U37509 ( .A(n36566), .B(n36565), .Z(n36567) );
  AND U37510 ( .A(n36568), .B(n36567), .Z(n36616) );
  XOR U37511 ( .A(n36617), .B(n36616), .Z(n36618) );
  NANDN U37512 ( .A(n36570), .B(n36569), .Z(n36574) );
  NANDN U37513 ( .A(n36572), .B(n36571), .Z(n36573) );
  NAND U37514 ( .A(n36574), .B(n36573), .Z(n36619) );
  XOR U37515 ( .A(n36618), .B(n36619), .Z(n36586) );
  OR U37516 ( .A(n36576), .B(n36575), .Z(n36580) );
  NANDN U37517 ( .A(n36578), .B(n36577), .Z(n36579) );
  NAND U37518 ( .A(n36580), .B(n36579), .Z(n36587) );
  XNOR U37519 ( .A(n36586), .B(n36587), .Z(n36588) );
  XNOR U37520 ( .A(n36589), .B(n36588), .Z(n36622) );
  XNOR U37521 ( .A(n36622), .B(sreg[1906]), .Z(n36624) );
  NAND U37522 ( .A(n36581), .B(sreg[1905]), .Z(n36585) );
  OR U37523 ( .A(n36583), .B(n36582), .Z(n36584) );
  AND U37524 ( .A(n36585), .B(n36584), .Z(n36623) );
  XOR U37525 ( .A(n36624), .B(n36623), .Z(c[1906]) );
  NANDN U37526 ( .A(n36587), .B(n36586), .Z(n36591) );
  NAND U37527 ( .A(n36589), .B(n36588), .Z(n36590) );
  NAND U37528 ( .A(n36591), .B(n36590), .Z(n36630) );
  NAND U37529 ( .A(b[0]), .B(a[891]), .Z(n36592) );
  XNOR U37530 ( .A(b[1]), .B(n36592), .Z(n36594) );
  NAND U37531 ( .A(n142), .B(a[890]), .Z(n36593) );
  AND U37532 ( .A(n36594), .B(n36593), .Z(n36647) );
  XOR U37533 ( .A(a[887]), .B(n42197), .Z(n36636) );
  NANDN U37534 ( .A(n36636), .B(n42173), .Z(n36597) );
  NANDN U37535 ( .A(n36595), .B(n42172), .Z(n36596) );
  NAND U37536 ( .A(n36597), .B(n36596), .Z(n36645) );
  NAND U37537 ( .A(b[7]), .B(a[883]), .Z(n36646) );
  XNOR U37538 ( .A(n36645), .B(n36646), .Z(n36648) );
  XOR U37539 ( .A(n36647), .B(n36648), .Z(n36654) );
  NANDN U37540 ( .A(n36598), .B(n42093), .Z(n36600) );
  XOR U37541 ( .A(n42134), .B(a[889]), .Z(n36639) );
  NANDN U37542 ( .A(n36639), .B(n42095), .Z(n36599) );
  NAND U37543 ( .A(n36600), .B(n36599), .Z(n36652) );
  NANDN U37544 ( .A(n36601), .B(n42231), .Z(n36603) );
  XOR U37545 ( .A(n235), .B(a[885]), .Z(n36642) );
  NANDN U37546 ( .A(n36642), .B(n42234), .Z(n36602) );
  AND U37547 ( .A(n36603), .B(n36602), .Z(n36651) );
  XNOR U37548 ( .A(n36652), .B(n36651), .Z(n36653) );
  XNOR U37549 ( .A(n36654), .B(n36653), .Z(n36658) );
  NANDN U37550 ( .A(n36605), .B(n36604), .Z(n36609) );
  NAND U37551 ( .A(n36607), .B(n36606), .Z(n36608) );
  AND U37552 ( .A(n36609), .B(n36608), .Z(n36657) );
  XOR U37553 ( .A(n36658), .B(n36657), .Z(n36659) );
  NANDN U37554 ( .A(n36611), .B(n36610), .Z(n36615) );
  NANDN U37555 ( .A(n36613), .B(n36612), .Z(n36614) );
  NAND U37556 ( .A(n36615), .B(n36614), .Z(n36660) );
  XOR U37557 ( .A(n36659), .B(n36660), .Z(n36627) );
  OR U37558 ( .A(n36617), .B(n36616), .Z(n36621) );
  NANDN U37559 ( .A(n36619), .B(n36618), .Z(n36620) );
  NAND U37560 ( .A(n36621), .B(n36620), .Z(n36628) );
  XNOR U37561 ( .A(n36627), .B(n36628), .Z(n36629) );
  XNOR U37562 ( .A(n36630), .B(n36629), .Z(n36663) );
  XNOR U37563 ( .A(n36663), .B(sreg[1907]), .Z(n36665) );
  NAND U37564 ( .A(n36622), .B(sreg[1906]), .Z(n36626) );
  OR U37565 ( .A(n36624), .B(n36623), .Z(n36625) );
  AND U37566 ( .A(n36626), .B(n36625), .Z(n36664) );
  XOR U37567 ( .A(n36665), .B(n36664), .Z(c[1907]) );
  NANDN U37568 ( .A(n36628), .B(n36627), .Z(n36632) );
  NAND U37569 ( .A(n36630), .B(n36629), .Z(n36631) );
  NAND U37570 ( .A(n36632), .B(n36631), .Z(n36671) );
  NAND U37571 ( .A(b[0]), .B(a[892]), .Z(n36633) );
  XNOR U37572 ( .A(b[1]), .B(n36633), .Z(n36635) );
  NAND U37573 ( .A(n142), .B(a[891]), .Z(n36634) );
  AND U37574 ( .A(n36635), .B(n36634), .Z(n36688) );
  XOR U37575 ( .A(a[888]), .B(n42197), .Z(n36677) );
  NANDN U37576 ( .A(n36677), .B(n42173), .Z(n36638) );
  NANDN U37577 ( .A(n36636), .B(n42172), .Z(n36637) );
  NAND U37578 ( .A(n36638), .B(n36637), .Z(n36686) );
  NAND U37579 ( .A(b[7]), .B(a[884]), .Z(n36687) );
  XNOR U37580 ( .A(n36686), .B(n36687), .Z(n36689) );
  XOR U37581 ( .A(n36688), .B(n36689), .Z(n36695) );
  NANDN U37582 ( .A(n36639), .B(n42093), .Z(n36641) );
  XOR U37583 ( .A(n42134), .B(a[890]), .Z(n36680) );
  NANDN U37584 ( .A(n36680), .B(n42095), .Z(n36640) );
  NAND U37585 ( .A(n36641), .B(n36640), .Z(n36693) );
  NANDN U37586 ( .A(n36642), .B(n42231), .Z(n36644) );
  XOR U37587 ( .A(n235), .B(a[886]), .Z(n36683) );
  NANDN U37588 ( .A(n36683), .B(n42234), .Z(n36643) );
  AND U37589 ( .A(n36644), .B(n36643), .Z(n36692) );
  XNOR U37590 ( .A(n36693), .B(n36692), .Z(n36694) );
  XNOR U37591 ( .A(n36695), .B(n36694), .Z(n36699) );
  NANDN U37592 ( .A(n36646), .B(n36645), .Z(n36650) );
  NAND U37593 ( .A(n36648), .B(n36647), .Z(n36649) );
  AND U37594 ( .A(n36650), .B(n36649), .Z(n36698) );
  XOR U37595 ( .A(n36699), .B(n36698), .Z(n36700) );
  NANDN U37596 ( .A(n36652), .B(n36651), .Z(n36656) );
  NANDN U37597 ( .A(n36654), .B(n36653), .Z(n36655) );
  NAND U37598 ( .A(n36656), .B(n36655), .Z(n36701) );
  XOR U37599 ( .A(n36700), .B(n36701), .Z(n36668) );
  OR U37600 ( .A(n36658), .B(n36657), .Z(n36662) );
  NANDN U37601 ( .A(n36660), .B(n36659), .Z(n36661) );
  NAND U37602 ( .A(n36662), .B(n36661), .Z(n36669) );
  XNOR U37603 ( .A(n36668), .B(n36669), .Z(n36670) );
  XNOR U37604 ( .A(n36671), .B(n36670), .Z(n36704) );
  XNOR U37605 ( .A(n36704), .B(sreg[1908]), .Z(n36706) );
  NAND U37606 ( .A(n36663), .B(sreg[1907]), .Z(n36667) );
  OR U37607 ( .A(n36665), .B(n36664), .Z(n36666) );
  AND U37608 ( .A(n36667), .B(n36666), .Z(n36705) );
  XOR U37609 ( .A(n36706), .B(n36705), .Z(c[1908]) );
  NANDN U37610 ( .A(n36669), .B(n36668), .Z(n36673) );
  NAND U37611 ( .A(n36671), .B(n36670), .Z(n36672) );
  NAND U37612 ( .A(n36673), .B(n36672), .Z(n36712) );
  NAND U37613 ( .A(b[0]), .B(a[893]), .Z(n36674) );
  XNOR U37614 ( .A(b[1]), .B(n36674), .Z(n36676) );
  NAND U37615 ( .A(n142), .B(a[892]), .Z(n36675) );
  AND U37616 ( .A(n36676), .B(n36675), .Z(n36729) );
  XOR U37617 ( .A(a[889]), .B(n42197), .Z(n36718) );
  NANDN U37618 ( .A(n36718), .B(n42173), .Z(n36679) );
  NANDN U37619 ( .A(n36677), .B(n42172), .Z(n36678) );
  NAND U37620 ( .A(n36679), .B(n36678), .Z(n36727) );
  NAND U37621 ( .A(b[7]), .B(a[885]), .Z(n36728) );
  XNOR U37622 ( .A(n36727), .B(n36728), .Z(n36730) );
  XOR U37623 ( .A(n36729), .B(n36730), .Z(n36736) );
  NANDN U37624 ( .A(n36680), .B(n42093), .Z(n36682) );
  XOR U37625 ( .A(n42134), .B(a[891]), .Z(n36721) );
  NANDN U37626 ( .A(n36721), .B(n42095), .Z(n36681) );
  NAND U37627 ( .A(n36682), .B(n36681), .Z(n36734) );
  NANDN U37628 ( .A(n36683), .B(n42231), .Z(n36685) );
  XOR U37629 ( .A(n236), .B(a[887]), .Z(n36724) );
  NANDN U37630 ( .A(n36724), .B(n42234), .Z(n36684) );
  AND U37631 ( .A(n36685), .B(n36684), .Z(n36733) );
  XNOR U37632 ( .A(n36734), .B(n36733), .Z(n36735) );
  XNOR U37633 ( .A(n36736), .B(n36735), .Z(n36740) );
  NANDN U37634 ( .A(n36687), .B(n36686), .Z(n36691) );
  NAND U37635 ( .A(n36689), .B(n36688), .Z(n36690) );
  AND U37636 ( .A(n36691), .B(n36690), .Z(n36739) );
  XOR U37637 ( .A(n36740), .B(n36739), .Z(n36741) );
  NANDN U37638 ( .A(n36693), .B(n36692), .Z(n36697) );
  NANDN U37639 ( .A(n36695), .B(n36694), .Z(n36696) );
  NAND U37640 ( .A(n36697), .B(n36696), .Z(n36742) );
  XOR U37641 ( .A(n36741), .B(n36742), .Z(n36709) );
  OR U37642 ( .A(n36699), .B(n36698), .Z(n36703) );
  NANDN U37643 ( .A(n36701), .B(n36700), .Z(n36702) );
  NAND U37644 ( .A(n36703), .B(n36702), .Z(n36710) );
  XNOR U37645 ( .A(n36709), .B(n36710), .Z(n36711) );
  XNOR U37646 ( .A(n36712), .B(n36711), .Z(n36745) );
  XNOR U37647 ( .A(n36745), .B(sreg[1909]), .Z(n36747) );
  NAND U37648 ( .A(n36704), .B(sreg[1908]), .Z(n36708) );
  OR U37649 ( .A(n36706), .B(n36705), .Z(n36707) );
  AND U37650 ( .A(n36708), .B(n36707), .Z(n36746) );
  XOR U37651 ( .A(n36747), .B(n36746), .Z(c[1909]) );
  NANDN U37652 ( .A(n36710), .B(n36709), .Z(n36714) );
  NAND U37653 ( .A(n36712), .B(n36711), .Z(n36713) );
  NAND U37654 ( .A(n36714), .B(n36713), .Z(n36753) );
  NAND U37655 ( .A(b[0]), .B(a[894]), .Z(n36715) );
  XNOR U37656 ( .A(b[1]), .B(n36715), .Z(n36717) );
  NAND U37657 ( .A(n142), .B(a[893]), .Z(n36716) );
  AND U37658 ( .A(n36717), .B(n36716), .Z(n36770) );
  XOR U37659 ( .A(a[890]), .B(n42197), .Z(n36759) );
  NANDN U37660 ( .A(n36759), .B(n42173), .Z(n36720) );
  NANDN U37661 ( .A(n36718), .B(n42172), .Z(n36719) );
  NAND U37662 ( .A(n36720), .B(n36719), .Z(n36768) );
  NAND U37663 ( .A(b[7]), .B(a[886]), .Z(n36769) );
  XNOR U37664 ( .A(n36768), .B(n36769), .Z(n36771) );
  XOR U37665 ( .A(n36770), .B(n36771), .Z(n36777) );
  NANDN U37666 ( .A(n36721), .B(n42093), .Z(n36723) );
  XOR U37667 ( .A(n42134), .B(a[892]), .Z(n36762) );
  NANDN U37668 ( .A(n36762), .B(n42095), .Z(n36722) );
  NAND U37669 ( .A(n36723), .B(n36722), .Z(n36775) );
  NANDN U37670 ( .A(n36724), .B(n42231), .Z(n36726) );
  XOR U37671 ( .A(n236), .B(a[888]), .Z(n36765) );
  NANDN U37672 ( .A(n36765), .B(n42234), .Z(n36725) );
  AND U37673 ( .A(n36726), .B(n36725), .Z(n36774) );
  XNOR U37674 ( .A(n36775), .B(n36774), .Z(n36776) );
  XNOR U37675 ( .A(n36777), .B(n36776), .Z(n36781) );
  NANDN U37676 ( .A(n36728), .B(n36727), .Z(n36732) );
  NAND U37677 ( .A(n36730), .B(n36729), .Z(n36731) );
  AND U37678 ( .A(n36732), .B(n36731), .Z(n36780) );
  XOR U37679 ( .A(n36781), .B(n36780), .Z(n36782) );
  NANDN U37680 ( .A(n36734), .B(n36733), .Z(n36738) );
  NANDN U37681 ( .A(n36736), .B(n36735), .Z(n36737) );
  NAND U37682 ( .A(n36738), .B(n36737), .Z(n36783) );
  XOR U37683 ( .A(n36782), .B(n36783), .Z(n36750) );
  OR U37684 ( .A(n36740), .B(n36739), .Z(n36744) );
  NANDN U37685 ( .A(n36742), .B(n36741), .Z(n36743) );
  NAND U37686 ( .A(n36744), .B(n36743), .Z(n36751) );
  XNOR U37687 ( .A(n36750), .B(n36751), .Z(n36752) );
  XNOR U37688 ( .A(n36753), .B(n36752), .Z(n36786) );
  XNOR U37689 ( .A(n36786), .B(sreg[1910]), .Z(n36788) );
  NAND U37690 ( .A(n36745), .B(sreg[1909]), .Z(n36749) );
  OR U37691 ( .A(n36747), .B(n36746), .Z(n36748) );
  AND U37692 ( .A(n36749), .B(n36748), .Z(n36787) );
  XOR U37693 ( .A(n36788), .B(n36787), .Z(c[1910]) );
  NANDN U37694 ( .A(n36751), .B(n36750), .Z(n36755) );
  NAND U37695 ( .A(n36753), .B(n36752), .Z(n36754) );
  NAND U37696 ( .A(n36755), .B(n36754), .Z(n36794) );
  NAND U37697 ( .A(b[0]), .B(a[895]), .Z(n36756) );
  XNOR U37698 ( .A(b[1]), .B(n36756), .Z(n36758) );
  NAND U37699 ( .A(n142), .B(a[894]), .Z(n36757) );
  AND U37700 ( .A(n36758), .B(n36757), .Z(n36811) );
  XOR U37701 ( .A(a[891]), .B(n42197), .Z(n36800) );
  NANDN U37702 ( .A(n36800), .B(n42173), .Z(n36761) );
  NANDN U37703 ( .A(n36759), .B(n42172), .Z(n36760) );
  NAND U37704 ( .A(n36761), .B(n36760), .Z(n36809) );
  NAND U37705 ( .A(b[7]), .B(a[887]), .Z(n36810) );
  XNOR U37706 ( .A(n36809), .B(n36810), .Z(n36812) );
  XOR U37707 ( .A(n36811), .B(n36812), .Z(n36818) );
  NANDN U37708 ( .A(n36762), .B(n42093), .Z(n36764) );
  XOR U37709 ( .A(n42134), .B(a[893]), .Z(n36803) );
  NANDN U37710 ( .A(n36803), .B(n42095), .Z(n36763) );
  NAND U37711 ( .A(n36764), .B(n36763), .Z(n36816) );
  NANDN U37712 ( .A(n36765), .B(n42231), .Z(n36767) );
  XOR U37713 ( .A(n236), .B(a[889]), .Z(n36806) );
  NANDN U37714 ( .A(n36806), .B(n42234), .Z(n36766) );
  AND U37715 ( .A(n36767), .B(n36766), .Z(n36815) );
  XNOR U37716 ( .A(n36816), .B(n36815), .Z(n36817) );
  XNOR U37717 ( .A(n36818), .B(n36817), .Z(n36822) );
  NANDN U37718 ( .A(n36769), .B(n36768), .Z(n36773) );
  NAND U37719 ( .A(n36771), .B(n36770), .Z(n36772) );
  AND U37720 ( .A(n36773), .B(n36772), .Z(n36821) );
  XOR U37721 ( .A(n36822), .B(n36821), .Z(n36823) );
  NANDN U37722 ( .A(n36775), .B(n36774), .Z(n36779) );
  NANDN U37723 ( .A(n36777), .B(n36776), .Z(n36778) );
  NAND U37724 ( .A(n36779), .B(n36778), .Z(n36824) );
  XOR U37725 ( .A(n36823), .B(n36824), .Z(n36791) );
  OR U37726 ( .A(n36781), .B(n36780), .Z(n36785) );
  NANDN U37727 ( .A(n36783), .B(n36782), .Z(n36784) );
  NAND U37728 ( .A(n36785), .B(n36784), .Z(n36792) );
  XNOR U37729 ( .A(n36791), .B(n36792), .Z(n36793) );
  XNOR U37730 ( .A(n36794), .B(n36793), .Z(n36827) );
  XNOR U37731 ( .A(n36827), .B(sreg[1911]), .Z(n36829) );
  NAND U37732 ( .A(n36786), .B(sreg[1910]), .Z(n36790) );
  OR U37733 ( .A(n36788), .B(n36787), .Z(n36789) );
  AND U37734 ( .A(n36790), .B(n36789), .Z(n36828) );
  XOR U37735 ( .A(n36829), .B(n36828), .Z(c[1911]) );
  NANDN U37736 ( .A(n36792), .B(n36791), .Z(n36796) );
  NAND U37737 ( .A(n36794), .B(n36793), .Z(n36795) );
  NAND U37738 ( .A(n36796), .B(n36795), .Z(n36835) );
  NAND U37739 ( .A(b[0]), .B(a[896]), .Z(n36797) );
  XNOR U37740 ( .A(b[1]), .B(n36797), .Z(n36799) );
  NAND U37741 ( .A(n143), .B(a[895]), .Z(n36798) );
  AND U37742 ( .A(n36799), .B(n36798), .Z(n36852) );
  XOR U37743 ( .A(a[892]), .B(n42197), .Z(n36841) );
  NANDN U37744 ( .A(n36841), .B(n42173), .Z(n36802) );
  NANDN U37745 ( .A(n36800), .B(n42172), .Z(n36801) );
  NAND U37746 ( .A(n36802), .B(n36801), .Z(n36850) );
  NAND U37747 ( .A(b[7]), .B(a[888]), .Z(n36851) );
  XNOR U37748 ( .A(n36850), .B(n36851), .Z(n36853) );
  XOR U37749 ( .A(n36852), .B(n36853), .Z(n36859) );
  NANDN U37750 ( .A(n36803), .B(n42093), .Z(n36805) );
  XOR U37751 ( .A(n42134), .B(a[894]), .Z(n36844) );
  NANDN U37752 ( .A(n36844), .B(n42095), .Z(n36804) );
  NAND U37753 ( .A(n36805), .B(n36804), .Z(n36857) );
  NANDN U37754 ( .A(n36806), .B(n42231), .Z(n36808) );
  XOR U37755 ( .A(n236), .B(a[890]), .Z(n36847) );
  NANDN U37756 ( .A(n36847), .B(n42234), .Z(n36807) );
  AND U37757 ( .A(n36808), .B(n36807), .Z(n36856) );
  XNOR U37758 ( .A(n36857), .B(n36856), .Z(n36858) );
  XNOR U37759 ( .A(n36859), .B(n36858), .Z(n36863) );
  NANDN U37760 ( .A(n36810), .B(n36809), .Z(n36814) );
  NAND U37761 ( .A(n36812), .B(n36811), .Z(n36813) );
  AND U37762 ( .A(n36814), .B(n36813), .Z(n36862) );
  XOR U37763 ( .A(n36863), .B(n36862), .Z(n36864) );
  NANDN U37764 ( .A(n36816), .B(n36815), .Z(n36820) );
  NANDN U37765 ( .A(n36818), .B(n36817), .Z(n36819) );
  NAND U37766 ( .A(n36820), .B(n36819), .Z(n36865) );
  XOR U37767 ( .A(n36864), .B(n36865), .Z(n36832) );
  OR U37768 ( .A(n36822), .B(n36821), .Z(n36826) );
  NANDN U37769 ( .A(n36824), .B(n36823), .Z(n36825) );
  NAND U37770 ( .A(n36826), .B(n36825), .Z(n36833) );
  XNOR U37771 ( .A(n36832), .B(n36833), .Z(n36834) );
  XNOR U37772 ( .A(n36835), .B(n36834), .Z(n36868) );
  XNOR U37773 ( .A(n36868), .B(sreg[1912]), .Z(n36870) );
  NAND U37774 ( .A(n36827), .B(sreg[1911]), .Z(n36831) );
  OR U37775 ( .A(n36829), .B(n36828), .Z(n36830) );
  AND U37776 ( .A(n36831), .B(n36830), .Z(n36869) );
  XOR U37777 ( .A(n36870), .B(n36869), .Z(c[1912]) );
  NANDN U37778 ( .A(n36833), .B(n36832), .Z(n36837) );
  NAND U37779 ( .A(n36835), .B(n36834), .Z(n36836) );
  NAND U37780 ( .A(n36837), .B(n36836), .Z(n36876) );
  NAND U37781 ( .A(b[0]), .B(a[897]), .Z(n36838) );
  XNOR U37782 ( .A(b[1]), .B(n36838), .Z(n36840) );
  NAND U37783 ( .A(n143), .B(a[896]), .Z(n36839) );
  AND U37784 ( .A(n36840), .B(n36839), .Z(n36893) );
  XOR U37785 ( .A(a[893]), .B(n42197), .Z(n36882) );
  NANDN U37786 ( .A(n36882), .B(n42173), .Z(n36843) );
  NANDN U37787 ( .A(n36841), .B(n42172), .Z(n36842) );
  NAND U37788 ( .A(n36843), .B(n36842), .Z(n36891) );
  NAND U37789 ( .A(b[7]), .B(a[889]), .Z(n36892) );
  XNOR U37790 ( .A(n36891), .B(n36892), .Z(n36894) );
  XOR U37791 ( .A(n36893), .B(n36894), .Z(n36900) );
  NANDN U37792 ( .A(n36844), .B(n42093), .Z(n36846) );
  XOR U37793 ( .A(n42134), .B(a[895]), .Z(n36885) );
  NANDN U37794 ( .A(n36885), .B(n42095), .Z(n36845) );
  NAND U37795 ( .A(n36846), .B(n36845), .Z(n36898) );
  NANDN U37796 ( .A(n36847), .B(n42231), .Z(n36849) );
  XOR U37797 ( .A(n236), .B(a[891]), .Z(n36888) );
  NANDN U37798 ( .A(n36888), .B(n42234), .Z(n36848) );
  AND U37799 ( .A(n36849), .B(n36848), .Z(n36897) );
  XNOR U37800 ( .A(n36898), .B(n36897), .Z(n36899) );
  XNOR U37801 ( .A(n36900), .B(n36899), .Z(n36904) );
  NANDN U37802 ( .A(n36851), .B(n36850), .Z(n36855) );
  NAND U37803 ( .A(n36853), .B(n36852), .Z(n36854) );
  AND U37804 ( .A(n36855), .B(n36854), .Z(n36903) );
  XOR U37805 ( .A(n36904), .B(n36903), .Z(n36905) );
  NANDN U37806 ( .A(n36857), .B(n36856), .Z(n36861) );
  NANDN U37807 ( .A(n36859), .B(n36858), .Z(n36860) );
  NAND U37808 ( .A(n36861), .B(n36860), .Z(n36906) );
  XOR U37809 ( .A(n36905), .B(n36906), .Z(n36873) );
  OR U37810 ( .A(n36863), .B(n36862), .Z(n36867) );
  NANDN U37811 ( .A(n36865), .B(n36864), .Z(n36866) );
  NAND U37812 ( .A(n36867), .B(n36866), .Z(n36874) );
  XNOR U37813 ( .A(n36873), .B(n36874), .Z(n36875) );
  XNOR U37814 ( .A(n36876), .B(n36875), .Z(n36909) );
  XNOR U37815 ( .A(n36909), .B(sreg[1913]), .Z(n36911) );
  NAND U37816 ( .A(n36868), .B(sreg[1912]), .Z(n36872) );
  OR U37817 ( .A(n36870), .B(n36869), .Z(n36871) );
  AND U37818 ( .A(n36872), .B(n36871), .Z(n36910) );
  XOR U37819 ( .A(n36911), .B(n36910), .Z(c[1913]) );
  NANDN U37820 ( .A(n36874), .B(n36873), .Z(n36878) );
  NAND U37821 ( .A(n36876), .B(n36875), .Z(n36877) );
  NAND U37822 ( .A(n36878), .B(n36877), .Z(n36917) );
  NAND U37823 ( .A(b[0]), .B(a[898]), .Z(n36879) );
  XNOR U37824 ( .A(b[1]), .B(n36879), .Z(n36881) );
  NAND U37825 ( .A(n143), .B(a[897]), .Z(n36880) );
  AND U37826 ( .A(n36881), .B(n36880), .Z(n36934) );
  XOR U37827 ( .A(a[894]), .B(n42197), .Z(n36923) );
  NANDN U37828 ( .A(n36923), .B(n42173), .Z(n36884) );
  NANDN U37829 ( .A(n36882), .B(n42172), .Z(n36883) );
  NAND U37830 ( .A(n36884), .B(n36883), .Z(n36932) );
  NAND U37831 ( .A(b[7]), .B(a[890]), .Z(n36933) );
  XNOR U37832 ( .A(n36932), .B(n36933), .Z(n36935) );
  XOR U37833 ( .A(n36934), .B(n36935), .Z(n36941) );
  NANDN U37834 ( .A(n36885), .B(n42093), .Z(n36887) );
  XOR U37835 ( .A(n42134), .B(a[896]), .Z(n36926) );
  NANDN U37836 ( .A(n36926), .B(n42095), .Z(n36886) );
  NAND U37837 ( .A(n36887), .B(n36886), .Z(n36939) );
  NANDN U37838 ( .A(n36888), .B(n42231), .Z(n36890) );
  XOR U37839 ( .A(n236), .B(a[892]), .Z(n36929) );
  NANDN U37840 ( .A(n36929), .B(n42234), .Z(n36889) );
  AND U37841 ( .A(n36890), .B(n36889), .Z(n36938) );
  XNOR U37842 ( .A(n36939), .B(n36938), .Z(n36940) );
  XNOR U37843 ( .A(n36941), .B(n36940), .Z(n36945) );
  NANDN U37844 ( .A(n36892), .B(n36891), .Z(n36896) );
  NAND U37845 ( .A(n36894), .B(n36893), .Z(n36895) );
  AND U37846 ( .A(n36896), .B(n36895), .Z(n36944) );
  XOR U37847 ( .A(n36945), .B(n36944), .Z(n36946) );
  NANDN U37848 ( .A(n36898), .B(n36897), .Z(n36902) );
  NANDN U37849 ( .A(n36900), .B(n36899), .Z(n36901) );
  NAND U37850 ( .A(n36902), .B(n36901), .Z(n36947) );
  XOR U37851 ( .A(n36946), .B(n36947), .Z(n36914) );
  OR U37852 ( .A(n36904), .B(n36903), .Z(n36908) );
  NANDN U37853 ( .A(n36906), .B(n36905), .Z(n36907) );
  NAND U37854 ( .A(n36908), .B(n36907), .Z(n36915) );
  XNOR U37855 ( .A(n36914), .B(n36915), .Z(n36916) );
  XNOR U37856 ( .A(n36917), .B(n36916), .Z(n36950) );
  XNOR U37857 ( .A(n36950), .B(sreg[1914]), .Z(n36952) );
  NAND U37858 ( .A(n36909), .B(sreg[1913]), .Z(n36913) );
  OR U37859 ( .A(n36911), .B(n36910), .Z(n36912) );
  AND U37860 ( .A(n36913), .B(n36912), .Z(n36951) );
  XOR U37861 ( .A(n36952), .B(n36951), .Z(c[1914]) );
  NANDN U37862 ( .A(n36915), .B(n36914), .Z(n36919) );
  NAND U37863 ( .A(n36917), .B(n36916), .Z(n36918) );
  NAND U37864 ( .A(n36919), .B(n36918), .Z(n36958) );
  NAND U37865 ( .A(b[0]), .B(a[899]), .Z(n36920) );
  XNOR U37866 ( .A(b[1]), .B(n36920), .Z(n36922) );
  NAND U37867 ( .A(n143), .B(a[898]), .Z(n36921) );
  AND U37868 ( .A(n36922), .B(n36921), .Z(n36975) );
  XOR U37869 ( .A(a[895]), .B(n42197), .Z(n36964) );
  NANDN U37870 ( .A(n36964), .B(n42173), .Z(n36925) );
  NANDN U37871 ( .A(n36923), .B(n42172), .Z(n36924) );
  NAND U37872 ( .A(n36925), .B(n36924), .Z(n36973) );
  NAND U37873 ( .A(b[7]), .B(a[891]), .Z(n36974) );
  XNOR U37874 ( .A(n36973), .B(n36974), .Z(n36976) );
  XOR U37875 ( .A(n36975), .B(n36976), .Z(n36982) );
  NANDN U37876 ( .A(n36926), .B(n42093), .Z(n36928) );
  XOR U37877 ( .A(n42134), .B(a[897]), .Z(n36967) );
  NANDN U37878 ( .A(n36967), .B(n42095), .Z(n36927) );
  NAND U37879 ( .A(n36928), .B(n36927), .Z(n36980) );
  NANDN U37880 ( .A(n36929), .B(n42231), .Z(n36931) );
  XOR U37881 ( .A(n236), .B(a[893]), .Z(n36970) );
  NANDN U37882 ( .A(n36970), .B(n42234), .Z(n36930) );
  AND U37883 ( .A(n36931), .B(n36930), .Z(n36979) );
  XNOR U37884 ( .A(n36980), .B(n36979), .Z(n36981) );
  XNOR U37885 ( .A(n36982), .B(n36981), .Z(n36986) );
  NANDN U37886 ( .A(n36933), .B(n36932), .Z(n36937) );
  NAND U37887 ( .A(n36935), .B(n36934), .Z(n36936) );
  AND U37888 ( .A(n36937), .B(n36936), .Z(n36985) );
  XOR U37889 ( .A(n36986), .B(n36985), .Z(n36987) );
  NANDN U37890 ( .A(n36939), .B(n36938), .Z(n36943) );
  NANDN U37891 ( .A(n36941), .B(n36940), .Z(n36942) );
  NAND U37892 ( .A(n36943), .B(n36942), .Z(n36988) );
  XOR U37893 ( .A(n36987), .B(n36988), .Z(n36955) );
  OR U37894 ( .A(n36945), .B(n36944), .Z(n36949) );
  NANDN U37895 ( .A(n36947), .B(n36946), .Z(n36948) );
  NAND U37896 ( .A(n36949), .B(n36948), .Z(n36956) );
  XNOR U37897 ( .A(n36955), .B(n36956), .Z(n36957) );
  XNOR U37898 ( .A(n36958), .B(n36957), .Z(n36991) );
  XNOR U37899 ( .A(n36991), .B(sreg[1915]), .Z(n36993) );
  NAND U37900 ( .A(n36950), .B(sreg[1914]), .Z(n36954) );
  OR U37901 ( .A(n36952), .B(n36951), .Z(n36953) );
  AND U37902 ( .A(n36954), .B(n36953), .Z(n36992) );
  XOR U37903 ( .A(n36993), .B(n36992), .Z(c[1915]) );
  NANDN U37904 ( .A(n36956), .B(n36955), .Z(n36960) );
  NAND U37905 ( .A(n36958), .B(n36957), .Z(n36959) );
  NAND U37906 ( .A(n36960), .B(n36959), .Z(n36999) );
  NAND U37907 ( .A(b[0]), .B(a[900]), .Z(n36961) );
  XNOR U37908 ( .A(b[1]), .B(n36961), .Z(n36963) );
  NAND U37909 ( .A(n143), .B(a[899]), .Z(n36962) );
  AND U37910 ( .A(n36963), .B(n36962), .Z(n37016) );
  XOR U37911 ( .A(a[896]), .B(n42197), .Z(n37005) );
  NANDN U37912 ( .A(n37005), .B(n42173), .Z(n36966) );
  NANDN U37913 ( .A(n36964), .B(n42172), .Z(n36965) );
  NAND U37914 ( .A(n36966), .B(n36965), .Z(n37014) );
  NAND U37915 ( .A(b[7]), .B(a[892]), .Z(n37015) );
  XNOR U37916 ( .A(n37014), .B(n37015), .Z(n37017) );
  XOR U37917 ( .A(n37016), .B(n37017), .Z(n37023) );
  NANDN U37918 ( .A(n36967), .B(n42093), .Z(n36969) );
  XOR U37919 ( .A(n42134), .B(a[898]), .Z(n37008) );
  NANDN U37920 ( .A(n37008), .B(n42095), .Z(n36968) );
  NAND U37921 ( .A(n36969), .B(n36968), .Z(n37021) );
  NANDN U37922 ( .A(n36970), .B(n42231), .Z(n36972) );
  XOR U37923 ( .A(n236), .B(a[894]), .Z(n37011) );
  NANDN U37924 ( .A(n37011), .B(n42234), .Z(n36971) );
  AND U37925 ( .A(n36972), .B(n36971), .Z(n37020) );
  XNOR U37926 ( .A(n37021), .B(n37020), .Z(n37022) );
  XNOR U37927 ( .A(n37023), .B(n37022), .Z(n37027) );
  NANDN U37928 ( .A(n36974), .B(n36973), .Z(n36978) );
  NAND U37929 ( .A(n36976), .B(n36975), .Z(n36977) );
  AND U37930 ( .A(n36978), .B(n36977), .Z(n37026) );
  XOR U37931 ( .A(n37027), .B(n37026), .Z(n37028) );
  NANDN U37932 ( .A(n36980), .B(n36979), .Z(n36984) );
  NANDN U37933 ( .A(n36982), .B(n36981), .Z(n36983) );
  NAND U37934 ( .A(n36984), .B(n36983), .Z(n37029) );
  XOR U37935 ( .A(n37028), .B(n37029), .Z(n36996) );
  OR U37936 ( .A(n36986), .B(n36985), .Z(n36990) );
  NANDN U37937 ( .A(n36988), .B(n36987), .Z(n36989) );
  NAND U37938 ( .A(n36990), .B(n36989), .Z(n36997) );
  XNOR U37939 ( .A(n36996), .B(n36997), .Z(n36998) );
  XNOR U37940 ( .A(n36999), .B(n36998), .Z(n37032) );
  XNOR U37941 ( .A(n37032), .B(sreg[1916]), .Z(n37034) );
  NAND U37942 ( .A(n36991), .B(sreg[1915]), .Z(n36995) );
  OR U37943 ( .A(n36993), .B(n36992), .Z(n36994) );
  AND U37944 ( .A(n36995), .B(n36994), .Z(n37033) );
  XOR U37945 ( .A(n37034), .B(n37033), .Z(c[1916]) );
  NANDN U37946 ( .A(n36997), .B(n36996), .Z(n37001) );
  NAND U37947 ( .A(n36999), .B(n36998), .Z(n37000) );
  NAND U37948 ( .A(n37001), .B(n37000), .Z(n37040) );
  NAND U37949 ( .A(b[0]), .B(a[901]), .Z(n37002) );
  XNOR U37950 ( .A(b[1]), .B(n37002), .Z(n37004) );
  NAND U37951 ( .A(n143), .B(a[900]), .Z(n37003) );
  AND U37952 ( .A(n37004), .B(n37003), .Z(n37057) );
  XOR U37953 ( .A(a[897]), .B(n42197), .Z(n37046) );
  NANDN U37954 ( .A(n37046), .B(n42173), .Z(n37007) );
  NANDN U37955 ( .A(n37005), .B(n42172), .Z(n37006) );
  NAND U37956 ( .A(n37007), .B(n37006), .Z(n37055) );
  NAND U37957 ( .A(b[7]), .B(a[893]), .Z(n37056) );
  XNOR U37958 ( .A(n37055), .B(n37056), .Z(n37058) );
  XOR U37959 ( .A(n37057), .B(n37058), .Z(n37064) );
  NANDN U37960 ( .A(n37008), .B(n42093), .Z(n37010) );
  XOR U37961 ( .A(n42134), .B(a[899]), .Z(n37049) );
  NANDN U37962 ( .A(n37049), .B(n42095), .Z(n37009) );
  NAND U37963 ( .A(n37010), .B(n37009), .Z(n37062) );
  NANDN U37964 ( .A(n37011), .B(n42231), .Z(n37013) );
  XOR U37965 ( .A(n236), .B(a[895]), .Z(n37052) );
  NANDN U37966 ( .A(n37052), .B(n42234), .Z(n37012) );
  AND U37967 ( .A(n37013), .B(n37012), .Z(n37061) );
  XNOR U37968 ( .A(n37062), .B(n37061), .Z(n37063) );
  XNOR U37969 ( .A(n37064), .B(n37063), .Z(n37068) );
  NANDN U37970 ( .A(n37015), .B(n37014), .Z(n37019) );
  NAND U37971 ( .A(n37017), .B(n37016), .Z(n37018) );
  AND U37972 ( .A(n37019), .B(n37018), .Z(n37067) );
  XOR U37973 ( .A(n37068), .B(n37067), .Z(n37069) );
  NANDN U37974 ( .A(n37021), .B(n37020), .Z(n37025) );
  NANDN U37975 ( .A(n37023), .B(n37022), .Z(n37024) );
  NAND U37976 ( .A(n37025), .B(n37024), .Z(n37070) );
  XOR U37977 ( .A(n37069), .B(n37070), .Z(n37037) );
  OR U37978 ( .A(n37027), .B(n37026), .Z(n37031) );
  NANDN U37979 ( .A(n37029), .B(n37028), .Z(n37030) );
  NAND U37980 ( .A(n37031), .B(n37030), .Z(n37038) );
  XNOR U37981 ( .A(n37037), .B(n37038), .Z(n37039) );
  XNOR U37982 ( .A(n37040), .B(n37039), .Z(n37073) );
  XNOR U37983 ( .A(n37073), .B(sreg[1917]), .Z(n37075) );
  NAND U37984 ( .A(n37032), .B(sreg[1916]), .Z(n37036) );
  OR U37985 ( .A(n37034), .B(n37033), .Z(n37035) );
  AND U37986 ( .A(n37036), .B(n37035), .Z(n37074) );
  XOR U37987 ( .A(n37075), .B(n37074), .Z(c[1917]) );
  NANDN U37988 ( .A(n37038), .B(n37037), .Z(n37042) );
  NAND U37989 ( .A(n37040), .B(n37039), .Z(n37041) );
  NAND U37990 ( .A(n37042), .B(n37041), .Z(n37081) );
  NAND U37991 ( .A(b[0]), .B(a[902]), .Z(n37043) );
  XNOR U37992 ( .A(b[1]), .B(n37043), .Z(n37045) );
  NAND U37993 ( .A(n143), .B(a[901]), .Z(n37044) );
  AND U37994 ( .A(n37045), .B(n37044), .Z(n37098) );
  XOR U37995 ( .A(a[898]), .B(n42197), .Z(n37087) );
  NANDN U37996 ( .A(n37087), .B(n42173), .Z(n37048) );
  NANDN U37997 ( .A(n37046), .B(n42172), .Z(n37047) );
  NAND U37998 ( .A(n37048), .B(n37047), .Z(n37096) );
  NAND U37999 ( .A(b[7]), .B(a[894]), .Z(n37097) );
  XNOR U38000 ( .A(n37096), .B(n37097), .Z(n37099) );
  XOR U38001 ( .A(n37098), .B(n37099), .Z(n37105) );
  NANDN U38002 ( .A(n37049), .B(n42093), .Z(n37051) );
  XOR U38003 ( .A(n42134), .B(a[900]), .Z(n37090) );
  NANDN U38004 ( .A(n37090), .B(n42095), .Z(n37050) );
  NAND U38005 ( .A(n37051), .B(n37050), .Z(n37103) );
  NANDN U38006 ( .A(n37052), .B(n42231), .Z(n37054) );
  XOR U38007 ( .A(n236), .B(a[896]), .Z(n37093) );
  NANDN U38008 ( .A(n37093), .B(n42234), .Z(n37053) );
  AND U38009 ( .A(n37054), .B(n37053), .Z(n37102) );
  XNOR U38010 ( .A(n37103), .B(n37102), .Z(n37104) );
  XNOR U38011 ( .A(n37105), .B(n37104), .Z(n37109) );
  NANDN U38012 ( .A(n37056), .B(n37055), .Z(n37060) );
  NAND U38013 ( .A(n37058), .B(n37057), .Z(n37059) );
  AND U38014 ( .A(n37060), .B(n37059), .Z(n37108) );
  XOR U38015 ( .A(n37109), .B(n37108), .Z(n37110) );
  NANDN U38016 ( .A(n37062), .B(n37061), .Z(n37066) );
  NANDN U38017 ( .A(n37064), .B(n37063), .Z(n37065) );
  NAND U38018 ( .A(n37066), .B(n37065), .Z(n37111) );
  XOR U38019 ( .A(n37110), .B(n37111), .Z(n37078) );
  OR U38020 ( .A(n37068), .B(n37067), .Z(n37072) );
  NANDN U38021 ( .A(n37070), .B(n37069), .Z(n37071) );
  NAND U38022 ( .A(n37072), .B(n37071), .Z(n37079) );
  XNOR U38023 ( .A(n37078), .B(n37079), .Z(n37080) );
  XNOR U38024 ( .A(n37081), .B(n37080), .Z(n37114) );
  XNOR U38025 ( .A(n37114), .B(sreg[1918]), .Z(n37116) );
  NAND U38026 ( .A(n37073), .B(sreg[1917]), .Z(n37077) );
  OR U38027 ( .A(n37075), .B(n37074), .Z(n37076) );
  AND U38028 ( .A(n37077), .B(n37076), .Z(n37115) );
  XOR U38029 ( .A(n37116), .B(n37115), .Z(c[1918]) );
  NANDN U38030 ( .A(n37079), .B(n37078), .Z(n37083) );
  NAND U38031 ( .A(n37081), .B(n37080), .Z(n37082) );
  NAND U38032 ( .A(n37083), .B(n37082), .Z(n37122) );
  NAND U38033 ( .A(b[0]), .B(a[903]), .Z(n37084) );
  XNOR U38034 ( .A(b[1]), .B(n37084), .Z(n37086) );
  NAND U38035 ( .A(n144), .B(a[902]), .Z(n37085) );
  AND U38036 ( .A(n37086), .B(n37085), .Z(n37139) );
  XOR U38037 ( .A(a[899]), .B(n42197), .Z(n37128) );
  NANDN U38038 ( .A(n37128), .B(n42173), .Z(n37089) );
  NANDN U38039 ( .A(n37087), .B(n42172), .Z(n37088) );
  NAND U38040 ( .A(n37089), .B(n37088), .Z(n37137) );
  NAND U38041 ( .A(b[7]), .B(a[895]), .Z(n37138) );
  XNOR U38042 ( .A(n37137), .B(n37138), .Z(n37140) );
  XOR U38043 ( .A(n37139), .B(n37140), .Z(n37146) );
  NANDN U38044 ( .A(n37090), .B(n42093), .Z(n37092) );
  XOR U38045 ( .A(n42134), .B(a[901]), .Z(n37131) );
  NANDN U38046 ( .A(n37131), .B(n42095), .Z(n37091) );
  NAND U38047 ( .A(n37092), .B(n37091), .Z(n37144) );
  NANDN U38048 ( .A(n37093), .B(n42231), .Z(n37095) );
  XOR U38049 ( .A(n236), .B(a[897]), .Z(n37134) );
  NANDN U38050 ( .A(n37134), .B(n42234), .Z(n37094) );
  AND U38051 ( .A(n37095), .B(n37094), .Z(n37143) );
  XNOR U38052 ( .A(n37144), .B(n37143), .Z(n37145) );
  XNOR U38053 ( .A(n37146), .B(n37145), .Z(n37150) );
  NANDN U38054 ( .A(n37097), .B(n37096), .Z(n37101) );
  NAND U38055 ( .A(n37099), .B(n37098), .Z(n37100) );
  AND U38056 ( .A(n37101), .B(n37100), .Z(n37149) );
  XOR U38057 ( .A(n37150), .B(n37149), .Z(n37151) );
  NANDN U38058 ( .A(n37103), .B(n37102), .Z(n37107) );
  NANDN U38059 ( .A(n37105), .B(n37104), .Z(n37106) );
  NAND U38060 ( .A(n37107), .B(n37106), .Z(n37152) );
  XOR U38061 ( .A(n37151), .B(n37152), .Z(n37119) );
  OR U38062 ( .A(n37109), .B(n37108), .Z(n37113) );
  NANDN U38063 ( .A(n37111), .B(n37110), .Z(n37112) );
  NAND U38064 ( .A(n37113), .B(n37112), .Z(n37120) );
  XNOR U38065 ( .A(n37119), .B(n37120), .Z(n37121) );
  XNOR U38066 ( .A(n37122), .B(n37121), .Z(n37155) );
  XNOR U38067 ( .A(n37155), .B(sreg[1919]), .Z(n37157) );
  NAND U38068 ( .A(n37114), .B(sreg[1918]), .Z(n37118) );
  OR U38069 ( .A(n37116), .B(n37115), .Z(n37117) );
  AND U38070 ( .A(n37118), .B(n37117), .Z(n37156) );
  XOR U38071 ( .A(n37157), .B(n37156), .Z(c[1919]) );
  NANDN U38072 ( .A(n37120), .B(n37119), .Z(n37124) );
  NAND U38073 ( .A(n37122), .B(n37121), .Z(n37123) );
  NAND U38074 ( .A(n37124), .B(n37123), .Z(n37163) );
  NAND U38075 ( .A(b[0]), .B(a[904]), .Z(n37125) );
  XNOR U38076 ( .A(b[1]), .B(n37125), .Z(n37127) );
  NAND U38077 ( .A(n144), .B(a[903]), .Z(n37126) );
  AND U38078 ( .A(n37127), .B(n37126), .Z(n37180) );
  XOR U38079 ( .A(a[900]), .B(n42197), .Z(n37169) );
  NANDN U38080 ( .A(n37169), .B(n42173), .Z(n37130) );
  NANDN U38081 ( .A(n37128), .B(n42172), .Z(n37129) );
  NAND U38082 ( .A(n37130), .B(n37129), .Z(n37178) );
  NAND U38083 ( .A(b[7]), .B(a[896]), .Z(n37179) );
  XNOR U38084 ( .A(n37178), .B(n37179), .Z(n37181) );
  XOR U38085 ( .A(n37180), .B(n37181), .Z(n37187) );
  NANDN U38086 ( .A(n37131), .B(n42093), .Z(n37133) );
  XOR U38087 ( .A(n42134), .B(a[902]), .Z(n37172) );
  NANDN U38088 ( .A(n37172), .B(n42095), .Z(n37132) );
  NAND U38089 ( .A(n37133), .B(n37132), .Z(n37185) );
  NANDN U38090 ( .A(n37134), .B(n42231), .Z(n37136) );
  XOR U38091 ( .A(n236), .B(a[898]), .Z(n37175) );
  NANDN U38092 ( .A(n37175), .B(n42234), .Z(n37135) );
  AND U38093 ( .A(n37136), .B(n37135), .Z(n37184) );
  XNOR U38094 ( .A(n37185), .B(n37184), .Z(n37186) );
  XNOR U38095 ( .A(n37187), .B(n37186), .Z(n37191) );
  NANDN U38096 ( .A(n37138), .B(n37137), .Z(n37142) );
  NAND U38097 ( .A(n37140), .B(n37139), .Z(n37141) );
  AND U38098 ( .A(n37142), .B(n37141), .Z(n37190) );
  XOR U38099 ( .A(n37191), .B(n37190), .Z(n37192) );
  NANDN U38100 ( .A(n37144), .B(n37143), .Z(n37148) );
  NANDN U38101 ( .A(n37146), .B(n37145), .Z(n37147) );
  NAND U38102 ( .A(n37148), .B(n37147), .Z(n37193) );
  XOR U38103 ( .A(n37192), .B(n37193), .Z(n37160) );
  OR U38104 ( .A(n37150), .B(n37149), .Z(n37154) );
  NANDN U38105 ( .A(n37152), .B(n37151), .Z(n37153) );
  NAND U38106 ( .A(n37154), .B(n37153), .Z(n37161) );
  XNOR U38107 ( .A(n37160), .B(n37161), .Z(n37162) );
  XNOR U38108 ( .A(n37163), .B(n37162), .Z(n37196) );
  XNOR U38109 ( .A(n37196), .B(sreg[1920]), .Z(n37198) );
  NAND U38110 ( .A(n37155), .B(sreg[1919]), .Z(n37159) );
  OR U38111 ( .A(n37157), .B(n37156), .Z(n37158) );
  AND U38112 ( .A(n37159), .B(n37158), .Z(n37197) );
  XOR U38113 ( .A(n37198), .B(n37197), .Z(c[1920]) );
  NANDN U38114 ( .A(n37161), .B(n37160), .Z(n37165) );
  NAND U38115 ( .A(n37163), .B(n37162), .Z(n37164) );
  NAND U38116 ( .A(n37165), .B(n37164), .Z(n37204) );
  NAND U38117 ( .A(b[0]), .B(a[905]), .Z(n37166) );
  XNOR U38118 ( .A(b[1]), .B(n37166), .Z(n37168) );
  NAND U38119 ( .A(n144), .B(a[904]), .Z(n37167) );
  AND U38120 ( .A(n37168), .B(n37167), .Z(n37221) );
  XOR U38121 ( .A(a[901]), .B(n42197), .Z(n37210) );
  NANDN U38122 ( .A(n37210), .B(n42173), .Z(n37171) );
  NANDN U38123 ( .A(n37169), .B(n42172), .Z(n37170) );
  NAND U38124 ( .A(n37171), .B(n37170), .Z(n37219) );
  NAND U38125 ( .A(b[7]), .B(a[897]), .Z(n37220) );
  XNOR U38126 ( .A(n37219), .B(n37220), .Z(n37222) );
  XOR U38127 ( .A(n37221), .B(n37222), .Z(n37228) );
  NANDN U38128 ( .A(n37172), .B(n42093), .Z(n37174) );
  XOR U38129 ( .A(n42134), .B(a[903]), .Z(n37213) );
  NANDN U38130 ( .A(n37213), .B(n42095), .Z(n37173) );
  NAND U38131 ( .A(n37174), .B(n37173), .Z(n37226) );
  NANDN U38132 ( .A(n37175), .B(n42231), .Z(n37177) );
  XOR U38133 ( .A(n237), .B(a[899]), .Z(n37216) );
  NANDN U38134 ( .A(n37216), .B(n42234), .Z(n37176) );
  AND U38135 ( .A(n37177), .B(n37176), .Z(n37225) );
  XNOR U38136 ( .A(n37226), .B(n37225), .Z(n37227) );
  XNOR U38137 ( .A(n37228), .B(n37227), .Z(n37232) );
  NANDN U38138 ( .A(n37179), .B(n37178), .Z(n37183) );
  NAND U38139 ( .A(n37181), .B(n37180), .Z(n37182) );
  AND U38140 ( .A(n37183), .B(n37182), .Z(n37231) );
  XOR U38141 ( .A(n37232), .B(n37231), .Z(n37233) );
  NANDN U38142 ( .A(n37185), .B(n37184), .Z(n37189) );
  NANDN U38143 ( .A(n37187), .B(n37186), .Z(n37188) );
  NAND U38144 ( .A(n37189), .B(n37188), .Z(n37234) );
  XOR U38145 ( .A(n37233), .B(n37234), .Z(n37201) );
  OR U38146 ( .A(n37191), .B(n37190), .Z(n37195) );
  NANDN U38147 ( .A(n37193), .B(n37192), .Z(n37194) );
  NAND U38148 ( .A(n37195), .B(n37194), .Z(n37202) );
  XNOR U38149 ( .A(n37201), .B(n37202), .Z(n37203) );
  XNOR U38150 ( .A(n37204), .B(n37203), .Z(n37237) );
  XNOR U38151 ( .A(n37237), .B(sreg[1921]), .Z(n37239) );
  NAND U38152 ( .A(n37196), .B(sreg[1920]), .Z(n37200) );
  OR U38153 ( .A(n37198), .B(n37197), .Z(n37199) );
  AND U38154 ( .A(n37200), .B(n37199), .Z(n37238) );
  XOR U38155 ( .A(n37239), .B(n37238), .Z(c[1921]) );
  NANDN U38156 ( .A(n37202), .B(n37201), .Z(n37206) );
  NAND U38157 ( .A(n37204), .B(n37203), .Z(n37205) );
  NAND U38158 ( .A(n37206), .B(n37205), .Z(n37245) );
  NAND U38159 ( .A(b[0]), .B(a[906]), .Z(n37207) );
  XNOR U38160 ( .A(b[1]), .B(n37207), .Z(n37209) );
  NAND U38161 ( .A(n144), .B(a[905]), .Z(n37208) );
  AND U38162 ( .A(n37209), .B(n37208), .Z(n37262) );
  XOR U38163 ( .A(a[902]), .B(n42197), .Z(n37251) );
  NANDN U38164 ( .A(n37251), .B(n42173), .Z(n37212) );
  NANDN U38165 ( .A(n37210), .B(n42172), .Z(n37211) );
  NAND U38166 ( .A(n37212), .B(n37211), .Z(n37260) );
  NAND U38167 ( .A(b[7]), .B(a[898]), .Z(n37261) );
  XNOR U38168 ( .A(n37260), .B(n37261), .Z(n37263) );
  XOR U38169 ( .A(n37262), .B(n37263), .Z(n37269) );
  NANDN U38170 ( .A(n37213), .B(n42093), .Z(n37215) );
  XOR U38171 ( .A(n42134), .B(a[904]), .Z(n37254) );
  NANDN U38172 ( .A(n37254), .B(n42095), .Z(n37214) );
  NAND U38173 ( .A(n37215), .B(n37214), .Z(n37267) );
  NANDN U38174 ( .A(n37216), .B(n42231), .Z(n37218) );
  XOR U38175 ( .A(n237), .B(a[900]), .Z(n37257) );
  NANDN U38176 ( .A(n37257), .B(n42234), .Z(n37217) );
  AND U38177 ( .A(n37218), .B(n37217), .Z(n37266) );
  XNOR U38178 ( .A(n37267), .B(n37266), .Z(n37268) );
  XNOR U38179 ( .A(n37269), .B(n37268), .Z(n37273) );
  NANDN U38180 ( .A(n37220), .B(n37219), .Z(n37224) );
  NAND U38181 ( .A(n37222), .B(n37221), .Z(n37223) );
  AND U38182 ( .A(n37224), .B(n37223), .Z(n37272) );
  XOR U38183 ( .A(n37273), .B(n37272), .Z(n37274) );
  NANDN U38184 ( .A(n37226), .B(n37225), .Z(n37230) );
  NANDN U38185 ( .A(n37228), .B(n37227), .Z(n37229) );
  NAND U38186 ( .A(n37230), .B(n37229), .Z(n37275) );
  XOR U38187 ( .A(n37274), .B(n37275), .Z(n37242) );
  OR U38188 ( .A(n37232), .B(n37231), .Z(n37236) );
  NANDN U38189 ( .A(n37234), .B(n37233), .Z(n37235) );
  NAND U38190 ( .A(n37236), .B(n37235), .Z(n37243) );
  XNOR U38191 ( .A(n37242), .B(n37243), .Z(n37244) );
  XNOR U38192 ( .A(n37245), .B(n37244), .Z(n37278) );
  XNOR U38193 ( .A(n37278), .B(sreg[1922]), .Z(n37280) );
  NAND U38194 ( .A(n37237), .B(sreg[1921]), .Z(n37241) );
  OR U38195 ( .A(n37239), .B(n37238), .Z(n37240) );
  AND U38196 ( .A(n37241), .B(n37240), .Z(n37279) );
  XOR U38197 ( .A(n37280), .B(n37279), .Z(c[1922]) );
  NANDN U38198 ( .A(n37243), .B(n37242), .Z(n37247) );
  NAND U38199 ( .A(n37245), .B(n37244), .Z(n37246) );
  NAND U38200 ( .A(n37247), .B(n37246), .Z(n37286) );
  NAND U38201 ( .A(b[0]), .B(a[907]), .Z(n37248) );
  XNOR U38202 ( .A(b[1]), .B(n37248), .Z(n37250) );
  NAND U38203 ( .A(n144), .B(a[906]), .Z(n37249) );
  AND U38204 ( .A(n37250), .B(n37249), .Z(n37303) );
  XOR U38205 ( .A(a[903]), .B(n42197), .Z(n37292) );
  NANDN U38206 ( .A(n37292), .B(n42173), .Z(n37253) );
  NANDN U38207 ( .A(n37251), .B(n42172), .Z(n37252) );
  NAND U38208 ( .A(n37253), .B(n37252), .Z(n37301) );
  NAND U38209 ( .A(b[7]), .B(a[899]), .Z(n37302) );
  XNOR U38210 ( .A(n37301), .B(n37302), .Z(n37304) );
  XOR U38211 ( .A(n37303), .B(n37304), .Z(n37310) );
  NANDN U38212 ( .A(n37254), .B(n42093), .Z(n37256) );
  XOR U38213 ( .A(n42134), .B(a[905]), .Z(n37295) );
  NANDN U38214 ( .A(n37295), .B(n42095), .Z(n37255) );
  NAND U38215 ( .A(n37256), .B(n37255), .Z(n37308) );
  NANDN U38216 ( .A(n37257), .B(n42231), .Z(n37259) );
  XOR U38217 ( .A(n237), .B(a[901]), .Z(n37298) );
  NANDN U38218 ( .A(n37298), .B(n42234), .Z(n37258) );
  AND U38219 ( .A(n37259), .B(n37258), .Z(n37307) );
  XNOR U38220 ( .A(n37308), .B(n37307), .Z(n37309) );
  XNOR U38221 ( .A(n37310), .B(n37309), .Z(n37314) );
  NANDN U38222 ( .A(n37261), .B(n37260), .Z(n37265) );
  NAND U38223 ( .A(n37263), .B(n37262), .Z(n37264) );
  AND U38224 ( .A(n37265), .B(n37264), .Z(n37313) );
  XOR U38225 ( .A(n37314), .B(n37313), .Z(n37315) );
  NANDN U38226 ( .A(n37267), .B(n37266), .Z(n37271) );
  NANDN U38227 ( .A(n37269), .B(n37268), .Z(n37270) );
  NAND U38228 ( .A(n37271), .B(n37270), .Z(n37316) );
  XOR U38229 ( .A(n37315), .B(n37316), .Z(n37283) );
  OR U38230 ( .A(n37273), .B(n37272), .Z(n37277) );
  NANDN U38231 ( .A(n37275), .B(n37274), .Z(n37276) );
  NAND U38232 ( .A(n37277), .B(n37276), .Z(n37284) );
  XNOR U38233 ( .A(n37283), .B(n37284), .Z(n37285) );
  XNOR U38234 ( .A(n37286), .B(n37285), .Z(n37319) );
  XNOR U38235 ( .A(n37319), .B(sreg[1923]), .Z(n37321) );
  NAND U38236 ( .A(n37278), .B(sreg[1922]), .Z(n37282) );
  OR U38237 ( .A(n37280), .B(n37279), .Z(n37281) );
  AND U38238 ( .A(n37282), .B(n37281), .Z(n37320) );
  XOR U38239 ( .A(n37321), .B(n37320), .Z(c[1923]) );
  NANDN U38240 ( .A(n37284), .B(n37283), .Z(n37288) );
  NAND U38241 ( .A(n37286), .B(n37285), .Z(n37287) );
  NAND U38242 ( .A(n37288), .B(n37287), .Z(n37327) );
  NAND U38243 ( .A(b[0]), .B(a[908]), .Z(n37289) );
  XNOR U38244 ( .A(b[1]), .B(n37289), .Z(n37291) );
  NAND U38245 ( .A(n144), .B(a[907]), .Z(n37290) );
  AND U38246 ( .A(n37291), .B(n37290), .Z(n37344) );
  XOR U38247 ( .A(a[904]), .B(n42197), .Z(n37333) );
  NANDN U38248 ( .A(n37333), .B(n42173), .Z(n37294) );
  NANDN U38249 ( .A(n37292), .B(n42172), .Z(n37293) );
  NAND U38250 ( .A(n37294), .B(n37293), .Z(n37342) );
  NAND U38251 ( .A(b[7]), .B(a[900]), .Z(n37343) );
  XNOR U38252 ( .A(n37342), .B(n37343), .Z(n37345) );
  XOR U38253 ( .A(n37344), .B(n37345), .Z(n37351) );
  NANDN U38254 ( .A(n37295), .B(n42093), .Z(n37297) );
  XOR U38255 ( .A(n42134), .B(a[906]), .Z(n37336) );
  NANDN U38256 ( .A(n37336), .B(n42095), .Z(n37296) );
  NAND U38257 ( .A(n37297), .B(n37296), .Z(n37349) );
  NANDN U38258 ( .A(n37298), .B(n42231), .Z(n37300) );
  XOR U38259 ( .A(n237), .B(a[902]), .Z(n37339) );
  NANDN U38260 ( .A(n37339), .B(n42234), .Z(n37299) );
  AND U38261 ( .A(n37300), .B(n37299), .Z(n37348) );
  XNOR U38262 ( .A(n37349), .B(n37348), .Z(n37350) );
  XNOR U38263 ( .A(n37351), .B(n37350), .Z(n37355) );
  NANDN U38264 ( .A(n37302), .B(n37301), .Z(n37306) );
  NAND U38265 ( .A(n37304), .B(n37303), .Z(n37305) );
  AND U38266 ( .A(n37306), .B(n37305), .Z(n37354) );
  XOR U38267 ( .A(n37355), .B(n37354), .Z(n37356) );
  NANDN U38268 ( .A(n37308), .B(n37307), .Z(n37312) );
  NANDN U38269 ( .A(n37310), .B(n37309), .Z(n37311) );
  NAND U38270 ( .A(n37312), .B(n37311), .Z(n37357) );
  XOR U38271 ( .A(n37356), .B(n37357), .Z(n37324) );
  OR U38272 ( .A(n37314), .B(n37313), .Z(n37318) );
  NANDN U38273 ( .A(n37316), .B(n37315), .Z(n37317) );
  NAND U38274 ( .A(n37318), .B(n37317), .Z(n37325) );
  XNOR U38275 ( .A(n37324), .B(n37325), .Z(n37326) );
  XNOR U38276 ( .A(n37327), .B(n37326), .Z(n37360) );
  XNOR U38277 ( .A(n37360), .B(sreg[1924]), .Z(n37362) );
  NAND U38278 ( .A(n37319), .B(sreg[1923]), .Z(n37323) );
  OR U38279 ( .A(n37321), .B(n37320), .Z(n37322) );
  AND U38280 ( .A(n37323), .B(n37322), .Z(n37361) );
  XOR U38281 ( .A(n37362), .B(n37361), .Z(c[1924]) );
  NANDN U38282 ( .A(n37325), .B(n37324), .Z(n37329) );
  NAND U38283 ( .A(n37327), .B(n37326), .Z(n37328) );
  NAND U38284 ( .A(n37329), .B(n37328), .Z(n37368) );
  NAND U38285 ( .A(b[0]), .B(a[909]), .Z(n37330) );
  XNOR U38286 ( .A(b[1]), .B(n37330), .Z(n37332) );
  NAND U38287 ( .A(n144), .B(a[908]), .Z(n37331) );
  AND U38288 ( .A(n37332), .B(n37331), .Z(n37385) );
  XOR U38289 ( .A(a[905]), .B(n42197), .Z(n37374) );
  NANDN U38290 ( .A(n37374), .B(n42173), .Z(n37335) );
  NANDN U38291 ( .A(n37333), .B(n42172), .Z(n37334) );
  NAND U38292 ( .A(n37335), .B(n37334), .Z(n37383) );
  NAND U38293 ( .A(b[7]), .B(a[901]), .Z(n37384) );
  XNOR U38294 ( .A(n37383), .B(n37384), .Z(n37386) );
  XOR U38295 ( .A(n37385), .B(n37386), .Z(n37392) );
  NANDN U38296 ( .A(n37336), .B(n42093), .Z(n37338) );
  XOR U38297 ( .A(n42134), .B(a[907]), .Z(n37377) );
  NANDN U38298 ( .A(n37377), .B(n42095), .Z(n37337) );
  NAND U38299 ( .A(n37338), .B(n37337), .Z(n37390) );
  NANDN U38300 ( .A(n37339), .B(n42231), .Z(n37341) );
  XOR U38301 ( .A(n237), .B(a[903]), .Z(n37380) );
  NANDN U38302 ( .A(n37380), .B(n42234), .Z(n37340) );
  AND U38303 ( .A(n37341), .B(n37340), .Z(n37389) );
  XNOR U38304 ( .A(n37390), .B(n37389), .Z(n37391) );
  XNOR U38305 ( .A(n37392), .B(n37391), .Z(n37396) );
  NANDN U38306 ( .A(n37343), .B(n37342), .Z(n37347) );
  NAND U38307 ( .A(n37345), .B(n37344), .Z(n37346) );
  AND U38308 ( .A(n37347), .B(n37346), .Z(n37395) );
  XOR U38309 ( .A(n37396), .B(n37395), .Z(n37397) );
  NANDN U38310 ( .A(n37349), .B(n37348), .Z(n37353) );
  NANDN U38311 ( .A(n37351), .B(n37350), .Z(n37352) );
  NAND U38312 ( .A(n37353), .B(n37352), .Z(n37398) );
  XOR U38313 ( .A(n37397), .B(n37398), .Z(n37365) );
  OR U38314 ( .A(n37355), .B(n37354), .Z(n37359) );
  NANDN U38315 ( .A(n37357), .B(n37356), .Z(n37358) );
  NAND U38316 ( .A(n37359), .B(n37358), .Z(n37366) );
  XNOR U38317 ( .A(n37365), .B(n37366), .Z(n37367) );
  XNOR U38318 ( .A(n37368), .B(n37367), .Z(n37401) );
  XNOR U38319 ( .A(n37401), .B(sreg[1925]), .Z(n37403) );
  NAND U38320 ( .A(n37360), .B(sreg[1924]), .Z(n37364) );
  OR U38321 ( .A(n37362), .B(n37361), .Z(n37363) );
  AND U38322 ( .A(n37364), .B(n37363), .Z(n37402) );
  XOR U38323 ( .A(n37403), .B(n37402), .Z(c[1925]) );
  NANDN U38324 ( .A(n37366), .B(n37365), .Z(n37370) );
  NAND U38325 ( .A(n37368), .B(n37367), .Z(n37369) );
  NAND U38326 ( .A(n37370), .B(n37369), .Z(n37409) );
  NAND U38327 ( .A(b[0]), .B(a[910]), .Z(n37371) );
  XNOR U38328 ( .A(b[1]), .B(n37371), .Z(n37373) );
  NAND U38329 ( .A(n145), .B(a[909]), .Z(n37372) );
  AND U38330 ( .A(n37373), .B(n37372), .Z(n37426) );
  XOR U38331 ( .A(a[906]), .B(n42197), .Z(n37415) );
  NANDN U38332 ( .A(n37415), .B(n42173), .Z(n37376) );
  NANDN U38333 ( .A(n37374), .B(n42172), .Z(n37375) );
  NAND U38334 ( .A(n37376), .B(n37375), .Z(n37424) );
  NAND U38335 ( .A(b[7]), .B(a[902]), .Z(n37425) );
  XNOR U38336 ( .A(n37424), .B(n37425), .Z(n37427) );
  XOR U38337 ( .A(n37426), .B(n37427), .Z(n37433) );
  NANDN U38338 ( .A(n37377), .B(n42093), .Z(n37379) );
  XOR U38339 ( .A(n42134), .B(a[908]), .Z(n37418) );
  NANDN U38340 ( .A(n37418), .B(n42095), .Z(n37378) );
  NAND U38341 ( .A(n37379), .B(n37378), .Z(n37431) );
  NANDN U38342 ( .A(n37380), .B(n42231), .Z(n37382) );
  XOR U38343 ( .A(n237), .B(a[904]), .Z(n37421) );
  NANDN U38344 ( .A(n37421), .B(n42234), .Z(n37381) );
  AND U38345 ( .A(n37382), .B(n37381), .Z(n37430) );
  XNOR U38346 ( .A(n37431), .B(n37430), .Z(n37432) );
  XNOR U38347 ( .A(n37433), .B(n37432), .Z(n37437) );
  NANDN U38348 ( .A(n37384), .B(n37383), .Z(n37388) );
  NAND U38349 ( .A(n37386), .B(n37385), .Z(n37387) );
  AND U38350 ( .A(n37388), .B(n37387), .Z(n37436) );
  XOR U38351 ( .A(n37437), .B(n37436), .Z(n37438) );
  NANDN U38352 ( .A(n37390), .B(n37389), .Z(n37394) );
  NANDN U38353 ( .A(n37392), .B(n37391), .Z(n37393) );
  NAND U38354 ( .A(n37394), .B(n37393), .Z(n37439) );
  XOR U38355 ( .A(n37438), .B(n37439), .Z(n37406) );
  OR U38356 ( .A(n37396), .B(n37395), .Z(n37400) );
  NANDN U38357 ( .A(n37398), .B(n37397), .Z(n37399) );
  NAND U38358 ( .A(n37400), .B(n37399), .Z(n37407) );
  XNOR U38359 ( .A(n37406), .B(n37407), .Z(n37408) );
  XNOR U38360 ( .A(n37409), .B(n37408), .Z(n37442) );
  XNOR U38361 ( .A(n37442), .B(sreg[1926]), .Z(n37444) );
  NAND U38362 ( .A(n37401), .B(sreg[1925]), .Z(n37405) );
  OR U38363 ( .A(n37403), .B(n37402), .Z(n37404) );
  AND U38364 ( .A(n37405), .B(n37404), .Z(n37443) );
  XOR U38365 ( .A(n37444), .B(n37443), .Z(c[1926]) );
  NANDN U38366 ( .A(n37407), .B(n37406), .Z(n37411) );
  NAND U38367 ( .A(n37409), .B(n37408), .Z(n37410) );
  NAND U38368 ( .A(n37411), .B(n37410), .Z(n37450) );
  NAND U38369 ( .A(b[0]), .B(a[911]), .Z(n37412) );
  XNOR U38370 ( .A(b[1]), .B(n37412), .Z(n37414) );
  NAND U38371 ( .A(n145), .B(a[910]), .Z(n37413) );
  AND U38372 ( .A(n37414), .B(n37413), .Z(n37467) );
  XOR U38373 ( .A(a[907]), .B(n42197), .Z(n37456) );
  NANDN U38374 ( .A(n37456), .B(n42173), .Z(n37417) );
  NANDN U38375 ( .A(n37415), .B(n42172), .Z(n37416) );
  NAND U38376 ( .A(n37417), .B(n37416), .Z(n37465) );
  NAND U38377 ( .A(b[7]), .B(a[903]), .Z(n37466) );
  XNOR U38378 ( .A(n37465), .B(n37466), .Z(n37468) );
  XOR U38379 ( .A(n37467), .B(n37468), .Z(n37474) );
  NANDN U38380 ( .A(n37418), .B(n42093), .Z(n37420) );
  XOR U38381 ( .A(n42134), .B(a[909]), .Z(n37459) );
  NANDN U38382 ( .A(n37459), .B(n42095), .Z(n37419) );
  NAND U38383 ( .A(n37420), .B(n37419), .Z(n37472) );
  NANDN U38384 ( .A(n37421), .B(n42231), .Z(n37423) );
  XOR U38385 ( .A(n237), .B(a[905]), .Z(n37462) );
  NANDN U38386 ( .A(n37462), .B(n42234), .Z(n37422) );
  AND U38387 ( .A(n37423), .B(n37422), .Z(n37471) );
  XNOR U38388 ( .A(n37472), .B(n37471), .Z(n37473) );
  XNOR U38389 ( .A(n37474), .B(n37473), .Z(n37478) );
  NANDN U38390 ( .A(n37425), .B(n37424), .Z(n37429) );
  NAND U38391 ( .A(n37427), .B(n37426), .Z(n37428) );
  AND U38392 ( .A(n37429), .B(n37428), .Z(n37477) );
  XOR U38393 ( .A(n37478), .B(n37477), .Z(n37479) );
  NANDN U38394 ( .A(n37431), .B(n37430), .Z(n37435) );
  NANDN U38395 ( .A(n37433), .B(n37432), .Z(n37434) );
  NAND U38396 ( .A(n37435), .B(n37434), .Z(n37480) );
  XOR U38397 ( .A(n37479), .B(n37480), .Z(n37447) );
  OR U38398 ( .A(n37437), .B(n37436), .Z(n37441) );
  NANDN U38399 ( .A(n37439), .B(n37438), .Z(n37440) );
  NAND U38400 ( .A(n37441), .B(n37440), .Z(n37448) );
  XNOR U38401 ( .A(n37447), .B(n37448), .Z(n37449) );
  XNOR U38402 ( .A(n37450), .B(n37449), .Z(n37483) );
  XNOR U38403 ( .A(n37483), .B(sreg[1927]), .Z(n37485) );
  NAND U38404 ( .A(n37442), .B(sreg[1926]), .Z(n37446) );
  OR U38405 ( .A(n37444), .B(n37443), .Z(n37445) );
  AND U38406 ( .A(n37446), .B(n37445), .Z(n37484) );
  XOR U38407 ( .A(n37485), .B(n37484), .Z(c[1927]) );
  NANDN U38408 ( .A(n37448), .B(n37447), .Z(n37452) );
  NAND U38409 ( .A(n37450), .B(n37449), .Z(n37451) );
  NAND U38410 ( .A(n37452), .B(n37451), .Z(n37491) );
  NAND U38411 ( .A(b[0]), .B(a[912]), .Z(n37453) );
  XNOR U38412 ( .A(b[1]), .B(n37453), .Z(n37455) );
  NAND U38413 ( .A(n145), .B(a[911]), .Z(n37454) );
  AND U38414 ( .A(n37455), .B(n37454), .Z(n37508) );
  XOR U38415 ( .A(a[908]), .B(n42197), .Z(n37497) );
  NANDN U38416 ( .A(n37497), .B(n42173), .Z(n37458) );
  NANDN U38417 ( .A(n37456), .B(n42172), .Z(n37457) );
  NAND U38418 ( .A(n37458), .B(n37457), .Z(n37506) );
  NAND U38419 ( .A(b[7]), .B(a[904]), .Z(n37507) );
  XNOR U38420 ( .A(n37506), .B(n37507), .Z(n37509) );
  XOR U38421 ( .A(n37508), .B(n37509), .Z(n37515) );
  NANDN U38422 ( .A(n37459), .B(n42093), .Z(n37461) );
  XOR U38423 ( .A(n42134), .B(a[910]), .Z(n37500) );
  NANDN U38424 ( .A(n37500), .B(n42095), .Z(n37460) );
  NAND U38425 ( .A(n37461), .B(n37460), .Z(n37513) );
  NANDN U38426 ( .A(n37462), .B(n42231), .Z(n37464) );
  XOR U38427 ( .A(n237), .B(a[906]), .Z(n37503) );
  NANDN U38428 ( .A(n37503), .B(n42234), .Z(n37463) );
  AND U38429 ( .A(n37464), .B(n37463), .Z(n37512) );
  XNOR U38430 ( .A(n37513), .B(n37512), .Z(n37514) );
  XNOR U38431 ( .A(n37515), .B(n37514), .Z(n37519) );
  NANDN U38432 ( .A(n37466), .B(n37465), .Z(n37470) );
  NAND U38433 ( .A(n37468), .B(n37467), .Z(n37469) );
  AND U38434 ( .A(n37470), .B(n37469), .Z(n37518) );
  XOR U38435 ( .A(n37519), .B(n37518), .Z(n37520) );
  NANDN U38436 ( .A(n37472), .B(n37471), .Z(n37476) );
  NANDN U38437 ( .A(n37474), .B(n37473), .Z(n37475) );
  NAND U38438 ( .A(n37476), .B(n37475), .Z(n37521) );
  XOR U38439 ( .A(n37520), .B(n37521), .Z(n37488) );
  OR U38440 ( .A(n37478), .B(n37477), .Z(n37482) );
  NANDN U38441 ( .A(n37480), .B(n37479), .Z(n37481) );
  NAND U38442 ( .A(n37482), .B(n37481), .Z(n37489) );
  XNOR U38443 ( .A(n37488), .B(n37489), .Z(n37490) );
  XNOR U38444 ( .A(n37491), .B(n37490), .Z(n37524) );
  XNOR U38445 ( .A(n37524), .B(sreg[1928]), .Z(n37526) );
  NAND U38446 ( .A(n37483), .B(sreg[1927]), .Z(n37487) );
  OR U38447 ( .A(n37485), .B(n37484), .Z(n37486) );
  AND U38448 ( .A(n37487), .B(n37486), .Z(n37525) );
  XOR U38449 ( .A(n37526), .B(n37525), .Z(c[1928]) );
  NANDN U38450 ( .A(n37489), .B(n37488), .Z(n37493) );
  NAND U38451 ( .A(n37491), .B(n37490), .Z(n37492) );
  NAND U38452 ( .A(n37493), .B(n37492), .Z(n37532) );
  NAND U38453 ( .A(b[0]), .B(a[913]), .Z(n37494) );
  XNOR U38454 ( .A(b[1]), .B(n37494), .Z(n37496) );
  NAND U38455 ( .A(n145), .B(a[912]), .Z(n37495) );
  AND U38456 ( .A(n37496), .B(n37495), .Z(n37549) );
  XOR U38457 ( .A(a[909]), .B(n42197), .Z(n37538) );
  NANDN U38458 ( .A(n37538), .B(n42173), .Z(n37499) );
  NANDN U38459 ( .A(n37497), .B(n42172), .Z(n37498) );
  NAND U38460 ( .A(n37499), .B(n37498), .Z(n37547) );
  NAND U38461 ( .A(b[7]), .B(a[905]), .Z(n37548) );
  XNOR U38462 ( .A(n37547), .B(n37548), .Z(n37550) );
  XOR U38463 ( .A(n37549), .B(n37550), .Z(n37556) );
  NANDN U38464 ( .A(n37500), .B(n42093), .Z(n37502) );
  XOR U38465 ( .A(n42134), .B(a[911]), .Z(n37541) );
  NANDN U38466 ( .A(n37541), .B(n42095), .Z(n37501) );
  NAND U38467 ( .A(n37502), .B(n37501), .Z(n37554) );
  NANDN U38468 ( .A(n37503), .B(n42231), .Z(n37505) );
  XOR U38469 ( .A(n237), .B(a[907]), .Z(n37544) );
  NANDN U38470 ( .A(n37544), .B(n42234), .Z(n37504) );
  AND U38471 ( .A(n37505), .B(n37504), .Z(n37553) );
  XNOR U38472 ( .A(n37554), .B(n37553), .Z(n37555) );
  XNOR U38473 ( .A(n37556), .B(n37555), .Z(n37560) );
  NANDN U38474 ( .A(n37507), .B(n37506), .Z(n37511) );
  NAND U38475 ( .A(n37509), .B(n37508), .Z(n37510) );
  AND U38476 ( .A(n37511), .B(n37510), .Z(n37559) );
  XOR U38477 ( .A(n37560), .B(n37559), .Z(n37561) );
  NANDN U38478 ( .A(n37513), .B(n37512), .Z(n37517) );
  NANDN U38479 ( .A(n37515), .B(n37514), .Z(n37516) );
  NAND U38480 ( .A(n37517), .B(n37516), .Z(n37562) );
  XOR U38481 ( .A(n37561), .B(n37562), .Z(n37529) );
  OR U38482 ( .A(n37519), .B(n37518), .Z(n37523) );
  NANDN U38483 ( .A(n37521), .B(n37520), .Z(n37522) );
  NAND U38484 ( .A(n37523), .B(n37522), .Z(n37530) );
  XNOR U38485 ( .A(n37529), .B(n37530), .Z(n37531) );
  XNOR U38486 ( .A(n37532), .B(n37531), .Z(n37565) );
  XNOR U38487 ( .A(n37565), .B(sreg[1929]), .Z(n37567) );
  NAND U38488 ( .A(n37524), .B(sreg[1928]), .Z(n37528) );
  OR U38489 ( .A(n37526), .B(n37525), .Z(n37527) );
  AND U38490 ( .A(n37528), .B(n37527), .Z(n37566) );
  XOR U38491 ( .A(n37567), .B(n37566), .Z(c[1929]) );
  NANDN U38492 ( .A(n37530), .B(n37529), .Z(n37534) );
  NAND U38493 ( .A(n37532), .B(n37531), .Z(n37533) );
  NAND U38494 ( .A(n37534), .B(n37533), .Z(n37573) );
  NAND U38495 ( .A(b[0]), .B(a[914]), .Z(n37535) );
  XNOR U38496 ( .A(b[1]), .B(n37535), .Z(n37537) );
  NAND U38497 ( .A(n145), .B(a[913]), .Z(n37536) );
  AND U38498 ( .A(n37537), .B(n37536), .Z(n37590) );
  XOR U38499 ( .A(a[910]), .B(n42197), .Z(n37579) );
  NANDN U38500 ( .A(n37579), .B(n42173), .Z(n37540) );
  NANDN U38501 ( .A(n37538), .B(n42172), .Z(n37539) );
  NAND U38502 ( .A(n37540), .B(n37539), .Z(n37588) );
  NAND U38503 ( .A(b[7]), .B(a[906]), .Z(n37589) );
  XNOR U38504 ( .A(n37588), .B(n37589), .Z(n37591) );
  XOR U38505 ( .A(n37590), .B(n37591), .Z(n37597) );
  NANDN U38506 ( .A(n37541), .B(n42093), .Z(n37543) );
  XOR U38507 ( .A(n42134), .B(a[912]), .Z(n37582) );
  NANDN U38508 ( .A(n37582), .B(n42095), .Z(n37542) );
  NAND U38509 ( .A(n37543), .B(n37542), .Z(n37595) );
  NANDN U38510 ( .A(n37544), .B(n42231), .Z(n37546) );
  XOR U38511 ( .A(n237), .B(a[908]), .Z(n37585) );
  NANDN U38512 ( .A(n37585), .B(n42234), .Z(n37545) );
  AND U38513 ( .A(n37546), .B(n37545), .Z(n37594) );
  XNOR U38514 ( .A(n37595), .B(n37594), .Z(n37596) );
  XNOR U38515 ( .A(n37597), .B(n37596), .Z(n37601) );
  NANDN U38516 ( .A(n37548), .B(n37547), .Z(n37552) );
  NAND U38517 ( .A(n37550), .B(n37549), .Z(n37551) );
  AND U38518 ( .A(n37552), .B(n37551), .Z(n37600) );
  XOR U38519 ( .A(n37601), .B(n37600), .Z(n37602) );
  NANDN U38520 ( .A(n37554), .B(n37553), .Z(n37558) );
  NANDN U38521 ( .A(n37556), .B(n37555), .Z(n37557) );
  NAND U38522 ( .A(n37558), .B(n37557), .Z(n37603) );
  XOR U38523 ( .A(n37602), .B(n37603), .Z(n37570) );
  OR U38524 ( .A(n37560), .B(n37559), .Z(n37564) );
  NANDN U38525 ( .A(n37562), .B(n37561), .Z(n37563) );
  NAND U38526 ( .A(n37564), .B(n37563), .Z(n37571) );
  XNOR U38527 ( .A(n37570), .B(n37571), .Z(n37572) );
  XNOR U38528 ( .A(n37573), .B(n37572), .Z(n37606) );
  XNOR U38529 ( .A(n37606), .B(sreg[1930]), .Z(n37608) );
  NAND U38530 ( .A(n37565), .B(sreg[1929]), .Z(n37569) );
  OR U38531 ( .A(n37567), .B(n37566), .Z(n37568) );
  AND U38532 ( .A(n37569), .B(n37568), .Z(n37607) );
  XOR U38533 ( .A(n37608), .B(n37607), .Z(c[1930]) );
  NANDN U38534 ( .A(n37571), .B(n37570), .Z(n37575) );
  NAND U38535 ( .A(n37573), .B(n37572), .Z(n37574) );
  NAND U38536 ( .A(n37575), .B(n37574), .Z(n37614) );
  NAND U38537 ( .A(b[0]), .B(a[915]), .Z(n37576) );
  XNOR U38538 ( .A(b[1]), .B(n37576), .Z(n37578) );
  NAND U38539 ( .A(n145), .B(a[914]), .Z(n37577) );
  AND U38540 ( .A(n37578), .B(n37577), .Z(n37631) );
  XOR U38541 ( .A(a[911]), .B(n42197), .Z(n37620) );
  NANDN U38542 ( .A(n37620), .B(n42173), .Z(n37581) );
  NANDN U38543 ( .A(n37579), .B(n42172), .Z(n37580) );
  NAND U38544 ( .A(n37581), .B(n37580), .Z(n37629) );
  NAND U38545 ( .A(b[7]), .B(a[907]), .Z(n37630) );
  XNOR U38546 ( .A(n37629), .B(n37630), .Z(n37632) );
  XOR U38547 ( .A(n37631), .B(n37632), .Z(n37638) );
  NANDN U38548 ( .A(n37582), .B(n42093), .Z(n37584) );
  XOR U38549 ( .A(n42134), .B(a[913]), .Z(n37623) );
  NANDN U38550 ( .A(n37623), .B(n42095), .Z(n37583) );
  NAND U38551 ( .A(n37584), .B(n37583), .Z(n37636) );
  NANDN U38552 ( .A(n37585), .B(n42231), .Z(n37587) );
  XOR U38553 ( .A(n237), .B(a[909]), .Z(n37626) );
  NANDN U38554 ( .A(n37626), .B(n42234), .Z(n37586) );
  AND U38555 ( .A(n37587), .B(n37586), .Z(n37635) );
  XNOR U38556 ( .A(n37636), .B(n37635), .Z(n37637) );
  XNOR U38557 ( .A(n37638), .B(n37637), .Z(n37642) );
  NANDN U38558 ( .A(n37589), .B(n37588), .Z(n37593) );
  NAND U38559 ( .A(n37591), .B(n37590), .Z(n37592) );
  AND U38560 ( .A(n37593), .B(n37592), .Z(n37641) );
  XOR U38561 ( .A(n37642), .B(n37641), .Z(n37643) );
  NANDN U38562 ( .A(n37595), .B(n37594), .Z(n37599) );
  NANDN U38563 ( .A(n37597), .B(n37596), .Z(n37598) );
  NAND U38564 ( .A(n37599), .B(n37598), .Z(n37644) );
  XOR U38565 ( .A(n37643), .B(n37644), .Z(n37611) );
  OR U38566 ( .A(n37601), .B(n37600), .Z(n37605) );
  NANDN U38567 ( .A(n37603), .B(n37602), .Z(n37604) );
  NAND U38568 ( .A(n37605), .B(n37604), .Z(n37612) );
  XNOR U38569 ( .A(n37611), .B(n37612), .Z(n37613) );
  XNOR U38570 ( .A(n37614), .B(n37613), .Z(n37647) );
  XNOR U38571 ( .A(n37647), .B(sreg[1931]), .Z(n37649) );
  NAND U38572 ( .A(n37606), .B(sreg[1930]), .Z(n37610) );
  OR U38573 ( .A(n37608), .B(n37607), .Z(n37609) );
  AND U38574 ( .A(n37610), .B(n37609), .Z(n37648) );
  XOR U38575 ( .A(n37649), .B(n37648), .Z(c[1931]) );
  NANDN U38576 ( .A(n37612), .B(n37611), .Z(n37616) );
  NAND U38577 ( .A(n37614), .B(n37613), .Z(n37615) );
  NAND U38578 ( .A(n37616), .B(n37615), .Z(n37655) );
  NAND U38579 ( .A(b[0]), .B(a[916]), .Z(n37617) );
  XNOR U38580 ( .A(b[1]), .B(n37617), .Z(n37619) );
  NAND U38581 ( .A(n145), .B(a[915]), .Z(n37618) );
  AND U38582 ( .A(n37619), .B(n37618), .Z(n37672) );
  XOR U38583 ( .A(a[912]), .B(n42197), .Z(n37661) );
  NANDN U38584 ( .A(n37661), .B(n42173), .Z(n37622) );
  NANDN U38585 ( .A(n37620), .B(n42172), .Z(n37621) );
  NAND U38586 ( .A(n37622), .B(n37621), .Z(n37670) );
  NAND U38587 ( .A(b[7]), .B(a[908]), .Z(n37671) );
  XNOR U38588 ( .A(n37670), .B(n37671), .Z(n37673) );
  XOR U38589 ( .A(n37672), .B(n37673), .Z(n37679) );
  NANDN U38590 ( .A(n37623), .B(n42093), .Z(n37625) );
  XOR U38591 ( .A(n42134), .B(a[914]), .Z(n37664) );
  NANDN U38592 ( .A(n37664), .B(n42095), .Z(n37624) );
  NAND U38593 ( .A(n37625), .B(n37624), .Z(n37677) );
  NANDN U38594 ( .A(n37626), .B(n42231), .Z(n37628) );
  XOR U38595 ( .A(n237), .B(a[910]), .Z(n37667) );
  NANDN U38596 ( .A(n37667), .B(n42234), .Z(n37627) );
  AND U38597 ( .A(n37628), .B(n37627), .Z(n37676) );
  XNOR U38598 ( .A(n37677), .B(n37676), .Z(n37678) );
  XNOR U38599 ( .A(n37679), .B(n37678), .Z(n37683) );
  NANDN U38600 ( .A(n37630), .B(n37629), .Z(n37634) );
  NAND U38601 ( .A(n37632), .B(n37631), .Z(n37633) );
  AND U38602 ( .A(n37634), .B(n37633), .Z(n37682) );
  XOR U38603 ( .A(n37683), .B(n37682), .Z(n37684) );
  NANDN U38604 ( .A(n37636), .B(n37635), .Z(n37640) );
  NANDN U38605 ( .A(n37638), .B(n37637), .Z(n37639) );
  NAND U38606 ( .A(n37640), .B(n37639), .Z(n37685) );
  XOR U38607 ( .A(n37684), .B(n37685), .Z(n37652) );
  OR U38608 ( .A(n37642), .B(n37641), .Z(n37646) );
  NANDN U38609 ( .A(n37644), .B(n37643), .Z(n37645) );
  NAND U38610 ( .A(n37646), .B(n37645), .Z(n37653) );
  XNOR U38611 ( .A(n37652), .B(n37653), .Z(n37654) );
  XNOR U38612 ( .A(n37655), .B(n37654), .Z(n37688) );
  XNOR U38613 ( .A(n37688), .B(sreg[1932]), .Z(n37690) );
  NAND U38614 ( .A(n37647), .B(sreg[1931]), .Z(n37651) );
  OR U38615 ( .A(n37649), .B(n37648), .Z(n37650) );
  AND U38616 ( .A(n37651), .B(n37650), .Z(n37689) );
  XOR U38617 ( .A(n37690), .B(n37689), .Z(c[1932]) );
  NANDN U38618 ( .A(n37653), .B(n37652), .Z(n37657) );
  NAND U38619 ( .A(n37655), .B(n37654), .Z(n37656) );
  NAND U38620 ( .A(n37657), .B(n37656), .Z(n37696) );
  NAND U38621 ( .A(b[0]), .B(a[917]), .Z(n37658) );
  XNOR U38622 ( .A(b[1]), .B(n37658), .Z(n37660) );
  NAND U38623 ( .A(n146), .B(a[916]), .Z(n37659) );
  AND U38624 ( .A(n37660), .B(n37659), .Z(n37713) );
  XOR U38625 ( .A(a[913]), .B(n42197), .Z(n37702) );
  NANDN U38626 ( .A(n37702), .B(n42173), .Z(n37663) );
  NANDN U38627 ( .A(n37661), .B(n42172), .Z(n37662) );
  NAND U38628 ( .A(n37663), .B(n37662), .Z(n37711) );
  NAND U38629 ( .A(b[7]), .B(a[909]), .Z(n37712) );
  XNOR U38630 ( .A(n37711), .B(n37712), .Z(n37714) );
  XOR U38631 ( .A(n37713), .B(n37714), .Z(n37720) );
  NANDN U38632 ( .A(n37664), .B(n42093), .Z(n37666) );
  XOR U38633 ( .A(n42134), .B(a[915]), .Z(n37705) );
  NANDN U38634 ( .A(n37705), .B(n42095), .Z(n37665) );
  NAND U38635 ( .A(n37666), .B(n37665), .Z(n37718) );
  NANDN U38636 ( .A(n37667), .B(n42231), .Z(n37669) );
  XOR U38637 ( .A(n238), .B(a[911]), .Z(n37708) );
  NANDN U38638 ( .A(n37708), .B(n42234), .Z(n37668) );
  AND U38639 ( .A(n37669), .B(n37668), .Z(n37717) );
  XNOR U38640 ( .A(n37718), .B(n37717), .Z(n37719) );
  XNOR U38641 ( .A(n37720), .B(n37719), .Z(n37724) );
  NANDN U38642 ( .A(n37671), .B(n37670), .Z(n37675) );
  NAND U38643 ( .A(n37673), .B(n37672), .Z(n37674) );
  AND U38644 ( .A(n37675), .B(n37674), .Z(n37723) );
  XOR U38645 ( .A(n37724), .B(n37723), .Z(n37725) );
  NANDN U38646 ( .A(n37677), .B(n37676), .Z(n37681) );
  NANDN U38647 ( .A(n37679), .B(n37678), .Z(n37680) );
  NAND U38648 ( .A(n37681), .B(n37680), .Z(n37726) );
  XOR U38649 ( .A(n37725), .B(n37726), .Z(n37693) );
  OR U38650 ( .A(n37683), .B(n37682), .Z(n37687) );
  NANDN U38651 ( .A(n37685), .B(n37684), .Z(n37686) );
  NAND U38652 ( .A(n37687), .B(n37686), .Z(n37694) );
  XNOR U38653 ( .A(n37693), .B(n37694), .Z(n37695) );
  XNOR U38654 ( .A(n37696), .B(n37695), .Z(n37729) );
  XNOR U38655 ( .A(n37729), .B(sreg[1933]), .Z(n37731) );
  NAND U38656 ( .A(n37688), .B(sreg[1932]), .Z(n37692) );
  OR U38657 ( .A(n37690), .B(n37689), .Z(n37691) );
  AND U38658 ( .A(n37692), .B(n37691), .Z(n37730) );
  XOR U38659 ( .A(n37731), .B(n37730), .Z(c[1933]) );
  NANDN U38660 ( .A(n37694), .B(n37693), .Z(n37698) );
  NAND U38661 ( .A(n37696), .B(n37695), .Z(n37697) );
  NAND U38662 ( .A(n37698), .B(n37697), .Z(n37737) );
  NAND U38663 ( .A(b[0]), .B(a[918]), .Z(n37699) );
  XNOR U38664 ( .A(b[1]), .B(n37699), .Z(n37701) );
  NAND U38665 ( .A(n146), .B(a[917]), .Z(n37700) );
  AND U38666 ( .A(n37701), .B(n37700), .Z(n37754) );
  XOR U38667 ( .A(a[914]), .B(n42197), .Z(n37743) );
  NANDN U38668 ( .A(n37743), .B(n42173), .Z(n37704) );
  NANDN U38669 ( .A(n37702), .B(n42172), .Z(n37703) );
  NAND U38670 ( .A(n37704), .B(n37703), .Z(n37752) );
  NAND U38671 ( .A(b[7]), .B(a[910]), .Z(n37753) );
  XNOR U38672 ( .A(n37752), .B(n37753), .Z(n37755) );
  XOR U38673 ( .A(n37754), .B(n37755), .Z(n37761) );
  NANDN U38674 ( .A(n37705), .B(n42093), .Z(n37707) );
  XOR U38675 ( .A(n42134), .B(a[916]), .Z(n37746) );
  NANDN U38676 ( .A(n37746), .B(n42095), .Z(n37706) );
  NAND U38677 ( .A(n37707), .B(n37706), .Z(n37759) );
  NANDN U38678 ( .A(n37708), .B(n42231), .Z(n37710) );
  XOR U38679 ( .A(n238), .B(a[912]), .Z(n37749) );
  NANDN U38680 ( .A(n37749), .B(n42234), .Z(n37709) );
  AND U38681 ( .A(n37710), .B(n37709), .Z(n37758) );
  XNOR U38682 ( .A(n37759), .B(n37758), .Z(n37760) );
  XNOR U38683 ( .A(n37761), .B(n37760), .Z(n37765) );
  NANDN U38684 ( .A(n37712), .B(n37711), .Z(n37716) );
  NAND U38685 ( .A(n37714), .B(n37713), .Z(n37715) );
  AND U38686 ( .A(n37716), .B(n37715), .Z(n37764) );
  XOR U38687 ( .A(n37765), .B(n37764), .Z(n37766) );
  NANDN U38688 ( .A(n37718), .B(n37717), .Z(n37722) );
  NANDN U38689 ( .A(n37720), .B(n37719), .Z(n37721) );
  NAND U38690 ( .A(n37722), .B(n37721), .Z(n37767) );
  XOR U38691 ( .A(n37766), .B(n37767), .Z(n37734) );
  OR U38692 ( .A(n37724), .B(n37723), .Z(n37728) );
  NANDN U38693 ( .A(n37726), .B(n37725), .Z(n37727) );
  NAND U38694 ( .A(n37728), .B(n37727), .Z(n37735) );
  XNOR U38695 ( .A(n37734), .B(n37735), .Z(n37736) );
  XNOR U38696 ( .A(n37737), .B(n37736), .Z(n37770) );
  XNOR U38697 ( .A(n37770), .B(sreg[1934]), .Z(n37772) );
  NAND U38698 ( .A(n37729), .B(sreg[1933]), .Z(n37733) );
  OR U38699 ( .A(n37731), .B(n37730), .Z(n37732) );
  AND U38700 ( .A(n37733), .B(n37732), .Z(n37771) );
  XOR U38701 ( .A(n37772), .B(n37771), .Z(c[1934]) );
  NANDN U38702 ( .A(n37735), .B(n37734), .Z(n37739) );
  NAND U38703 ( .A(n37737), .B(n37736), .Z(n37738) );
  NAND U38704 ( .A(n37739), .B(n37738), .Z(n37778) );
  NAND U38705 ( .A(b[0]), .B(a[919]), .Z(n37740) );
  XNOR U38706 ( .A(b[1]), .B(n37740), .Z(n37742) );
  NAND U38707 ( .A(n146), .B(a[918]), .Z(n37741) );
  AND U38708 ( .A(n37742), .B(n37741), .Z(n37795) );
  XOR U38709 ( .A(a[915]), .B(n42197), .Z(n37784) );
  NANDN U38710 ( .A(n37784), .B(n42173), .Z(n37745) );
  NANDN U38711 ( .A(n37743), .B(n42172), .Z(n37744) );
  NAND U38712 ( .A(n37745), .B(n37744), .Z(n37793) );
  NAND U38713 ( .A(b[7]), .B(a[911]), .Z(n37794) );
  XNOR U38714 ( .A(n37793), .B(n37794), .Z(n37796) );
  XOR U38715 ( .A(n37795), .B(n37796), .Z(n37802) );
  NANDN U38716 ( .A(n37746), .B(n42093), .Z(n37748) );
  XOR U38717 ( .A(n42134), .B(a[917]), .Z(n37787) );
  NANDN U38718 ( .A(n37787), .B(n42095), .Z(n37747) );
  NAND U38719 ( .A(n37748), .B(n37747), .Z(n37800) );
  NANDN U38720 ( .A(n37749), .B(n42231), .Z(n37751) );
  XOR U38721 ( .A(n238), .B(a[913]), .Z(n37790) );
  NANDN U38722 ( .A(n37790), .B(n42234), .Z(n37750) );
  AND U38723 ( .A(n37751), .B(n37750), .Z(n37799) );
  XNOR U38724 ( .A(n37800), .B(n37799), .Z(n37801) );
  XNOR U38725 ( .A(n37802), .B(n37801), .Z(n37806) );
  NANDN U38726 ( .A(n37753), .B(n37752), .Z(n37757) );
  NAND U38727 ( .A(n37755), .B(n37754), .Z(n37756) );
  AND U38728 ( .A(n37757), .B(n37756), .Z(n37805) );
  XOR U38729 ( .A(n37806), .B(n37805), .Z(n37807) );
  NANDN U38730 ( .A(n37759), .B(n37758), .Z(n37763) );
  NANDN U38731 ( .A(n37761), .B(n37760), .Z(n37762) );
  NAND U38732 ( .A(n37763), .B(n37762), .Z(n37808) );
  XOR U38733 ( .A(n37807), .B(n37808), .Z(n37775) );
  OR U38734 ( .A(n37765), .B(n37764), .Z(n37769) );
  NANDN U38735 ( .A(n37767), .B(n37766), .Z(n37768) );
  NAND U38736 ( .A(n37769), .B(n37768), .Z(n37776) );
  XNOR U38737 ( .A(n37775), .B(n37776), .Z(n37777) );
  XNOR U38738 ( .A(n37778), .B(n37777), .Z(n37811) );
  XNOR U38739 ( .A(n37811), .B(sreg[1935]), .Z(n37813) );
  NAND U38740 ( .A(n37770), .B(sreg[1934]), .Z(n37774) );
  OR U38741 ( .A(n37772), .B(n37771), .Z(n37773) );
  AND U38742 ( .A(n37774), .B(n37773), .Z(n37812) );
  XOR U38743 ( .A(n37813), .B(n37812), .Z(c[1935]) );
  NANDN U38744 ( .A(n37776), .B(n37775), .Z(n37780) );
  NAND U38745 ( .A(n37778), .B(n37777), .Z(n37779) );
  NAND U38746 ( .A(n37780), .B(n37779), .Z(n37819) );
  NAND U38747 ( .A(b[0]), .B(a[920]), .Z(n37781) );
  XNOR U38748 ( .A(b[1]), .B(n37781), .Z(n37783) );
  NAND U38749 ( .A(n146), .B(a[919]), .Z(n37782) );
  AND U38750 ( .A(n37783), .B(n37782), .Z(n37836) );
  XOR U38751 ( .A(a[916]), .B(n42197), .Z(n37825) );
  NANDN U38752 ( .A(n37825), .B(n42173), .Z(n37786) );
  NANDN U38753 ( .A(n37784), .B(n42172), .Z(n37785) );
  NAND U38754 ( .A(n37786), .B(n37785), .Z(n37834) );
  NAND U38755 ( .A(b[7]), .B(a[912]), .Z(n37835) );
  XNOR U38756 ( .A(n37834), .B(n37835), .Z(n37837) );
  XOR U38757 ( .A(n37836), .B(n37837), .Z(n37843) );
  NANDN U38758 ( .A(n37787), .B(n42093), .Z(n37789) );
  XOR U38759 ( .A(n42134), .B(a[918]), .Z(n37828) );
  NANDN U38760 ( .A(n37828), .B(n42095), .Z(n37788) );
  NAND U38761 ( .A(n37789), .B(n37788), .Z(n37841) );
  NANDN U38762 ( .A(n37790), .B(n42231), .Z(n37792) );
  XOR U38763 ( .A(n238), .B(a[914]), .Z(n37831) );
  NANDN U38764 ( .A(n37831), .B(n42234), .Z(n37791) );
  AND U38765 ( .A(n37792), .B(n37791), .Z(n37840) );
  XNOR U38766 ( .A(n37841), .B(n37840), .Z(n37842) );
  XNOR U38767 ( .A(n37843), .B(n37842), .Z(n37847) );
  NANDN U38768 ( .A(n37794), .B(n37793), .Z(n37798) );
  NAND U38769 ( .A(n37796), .B(n37795), .Z(n37797) );
  AND U38770 ( .A(n37798), .B(n37797), .Z(n37846) );
  XOR U38771 ( .A(n37847), .B(n37846), .Z(n37848) );
  NANDN U38772 ( .A(n37800), .B(n37799), .Z(n37804) );
  NANDN U38773 ( .A(n37802), .B(n37801), .Z(n37803) );
  NAND U38774 ( .A(n37804), .B(n37803), .Z(n37849) );
  XOR U38775 ( .A(n37848), .B(n37849), .Z(n37816) );
  OR U38776 ( .A(n37806), .B(n37805), .Z(n37810) );
  NANDN U38777 ( .A(n37808), .B(n37807), .Z(n37809) );
  NAND U38778 ( .A(n37810), .B(n37809), .Z(n37817) );
  XNOR U38779 ( .A(n37816), .B(n37817), .Z(n37818) );
  XNOR U38780 ( .A(n37819), .B(n37818), .Z(n37852) );
  XNOR U38781 ( .A(n37852), .B(sreg[1936]), .Z(n37854) );
  NAND U38782 ( .A(n37811), .B(sreg[1935]), .Z(n37815) );
  OR U38783 ( .A(n37813), .B(n37812), .Z(n37814) );
  AND U38784 ( .A(n37815), .B(n37814), .Z(n37853) );
  XOR U38785 ( .A(n37854), .B(n37853), .Z(c[1936]) );
  NANDN U38786 ( .A(n37817), .B(n37816), .Z(n37821) );
  NAND U38787 ( .A(n37819), .B(n37818), .Z(n37820) );
  NAND U38788 ( .A(n37821), .B(n37820), .Z(n37860) );
  NAND U38789 ( .A(b[0]), .B(a[921]), .Z(n37822) );
  XNOR U38790 ( .A(b[1]), .B(n37822), .Z(n37824) );
  NAND U38791 ( .A(n146), .B(a[920]), .Z(n37823) );
  AND U38792 ( .A(n37824), .B(n37823), .Z(n37877) );
  XOR U38793 ( .A(a[917]), .B(n42197), .Z(n37866) );
  NANDN U38794 ( .A(n37866), .B(n42173), .Z(n37827) );
  NANDN U38795 ( .A(n37825), .B(n42172), .Z(n37826) );
  NAND U38796 ( .A(n37827), .B(n37826), .Z(n37875) );
  NAND U38797 ( .A(b[7]), .B(a[913]), .Z(n37876) );
  XNOR U38798 ( .A(n37875), .B(n37876), .Z(n37878) );
  XOR U38799 ( .A(n37877), .B(n37878), .Z(n37884) );
  NANDN U38800 ( .A(n37828), .B(n42093), .Z(n37830) );
  XOR U38801 ( .A(n42134), .B(a[919]), .Z(n37869) );
  NANDN U38802 ( .A(n37869), .B(n42095), .Z(n37829) );
  NAND U38803 ( .A(n37830), .B(n37829), .Z(n37882) );
  NANDN U38804 ( .A(n37831), .B(n42231), .Z(n37833) );
  XOR U38805 ( .A(n238), .B(a[915]), .Z(n37872) );
  NANDN U38806 ( .A(n37872), .B(n42234), .Z(n37832) );
  AND U38807 ( .A(n37833), .B(n37832), .Z(n37881) );
  XNOR U38808 ( .A(n37882), .B(n37881), .Z(n37883) );
  XNOR U38809 ( .A(n37884), .B(n37883), .Z(n37888) );
  NANDN U38810 ( .A(n37835), .B(n37834), .Z(n37839) );
  NAND U38811 ( .A(n37837), .B(n37836), .Z(n37838) );
  AND U38812 ( .A(n37839), .B(n37838), .Z(n37887) );
  XOR U38813 ( .A(n37888), .B(n37887), .Z(n37889) );
  NANDN U38814 ( .A(n37841), .B(n37840), .Z(n37845) );
  NANDN U38815 ( .A(n37843), .B(n37842), .Z(n37844) );
  NAND U38816 ( .A(n37845), .B(n37844), .Z(n37890) );
  XOR U38817 ( .A(n37889), .B(n37890), .Z(n37857) );
  OR U38818 ( .A(n37847), .B(n37846), .Z(n37851) );
  NANDN U38819 ( .A(n37849), .B(n37848), .Z(n37850) );
  NAND U38820 ( .A(n37851), .B(n37850), .Z(n37858) );
  XNOR U38821 ( .A(n37857), .B(n37858), .Z(n37859) );
  XNOR U38822 ( .A(n37860), .B(n37859), .Z(n37893) );
  XNOR U38823 ( .A(n37893), .B(sreg[1937]), .Z(n37895) );
  NAND U38824 ( .A(n37852), .B(sreg[1936]), .Z(n37856) );
  OR U38825 ( .A(n37854), .B(n37853), .Z(n37855) );
  AND U38826 ( .A(n37856), .B(n37855), .Z(n37894) );
  XOR U38827 ( .A(n37895), .B(n37894), .Z(c[1937]) );
  NANDN U38828 ( .A(n37858), .B(n37857), .Z(n37862) );
  NAND U38829 ( .A(n37860), .B(n37859), .Z(n37861) );
  NAND U38830 ( .A(n37862), .B(n37861), .Z(n37901) );
  NAND U38831 ( .A(b[0]), .B(a[922]), .Z(n37863) );
  XNOR U38832 ( .A(b[1]), .B(n37863), .Z(n37865) );
  NAND U38833 ( .A(n146), .B(a[921]), .Z(n37864) );
  AND U38834 ( .A(n37865), .B(n37864), .Z(n37918) );
  XOR U38835 ( .A(a[918]), .B(n42197), .Z(n37907) );
  NANDN U38836 ( .A(n37907), .B(n42173), .Z(n37868) );
  NANDN U38837 ( .A(n37866), .B(n42172), .Z(n37867) );
  NAND U38838 ( .A(n37868), .B(n37867), .Z(n37916) );
  NAND U38839 ( .A(b[7]), .B(a[914]), .Z(n37917) );
  XNOR U38840 ( .A(n37916), .B(n37917), .Z(n37919) );
  XOR U38841 ( .A(n37918), .B(n37919), .Z(n37925) );
  NANDN U38842 ( .A(n37869), .B(n42093), .Z(n37871) );
  XOR U38843 ( .A(n42134), .B(a[920]), .Z(n37910) );
  NANDN U38844 ( .A(n37910), .B(n42095), .Z(n37870) );
  NAND U38845 ( .A(n37871), .B(n37870), .Z(n37923) );
  NANDN U38846 ( .A(n37872), .B(n42231), .Z(n37874) );
  XOR U38847 ( .A(n238), .B(a[916]), .Z(n37913) );
  NANDN U38848 ( .A(n37913), .B(n42234), .Z(n37873) );
  AND U38849 ( .A(n37874), .B(n37873), .Z(n37922) );
  XNOR U38850 ( .A(n37923), .B(n37922), .Z(n37924) );
  XNOR U38851 ( .A(n37925), .B(n37924), .Z(n37929) );
  NANDN U38852 ( .A(n37876), .B(n37875), .Z(n37880) );
  NAND U38853 ( .A(n37878), .B(n37877), .Z(n37879) );
  AND U38854 ( .A(n37880), .B(n37879), .Z(n37928) );
  XOR U38855 ( .A(n37929), .B(n37928), .Z(n37930) );
  NANDN U38856 ( .A(n37882), .B(n37881), .Z(n37886) );
  NANDN U38857 ( .A(n37884), .B(n37883), .Z(n37885) );
  NAND U38858 ( .A(n37886), .B(n37885), .Z(n37931) );
  XOR U38859 ( .A(n37930), .B(n37931), .Z(n37898) );
  OR U38860 ( .A(n37888), .B(n37887), .Z(n37892) );
  NANDN U38861 ( .A(n37890), .B(n37889), .Z(n37891) );
  NAND U38862 ( .A(n37892), .B(n37891), .Z(n37899) );
  XNOR U38863 ( .A(n37898), .B(n37899), .Z(n37900) );
  XNOR U38864 ( .A(n37901), .B(n37900), .Z(n37934) );
  XNOR U38865 ( .A(n37934), .B(sreg[1938]), .Z(n37936) );
  NAND U38866 ( .A(n37893), .B(sreg[1937]), .Z(n37897) );
  OR U38867 ( .A(n37895), .B(n37894), .Z(n37896) );
  AND U38868 ( .A(n37897), .B(n37896), .Z(n37935) );
  XOR U38869 ( .A(n37936), .B(n37935), .Z(c[1938]) );
  NANDN U38870 ( .A(n37899), .B(n37898), .Z(n37903) );
  NAND U38871 ( .A(n37901), .B(n37900), .Z(n37902) );
  NAND U38872 ( .A(n37903), .B(n37902), .Z(n37942) );
  NAND U38873 ( .A(b[0]), .B(a[923]), .Z(n37904) );
  XNOR U38874 ( .A(b[1]), .B(n37904), .Z(n37906) );
  NAND U38875 ( .A(n146), .B(a[922]), .Z(n37905) );
  AND U38876 ( .A(n37906), .B(n37905), .Z(n37959) );
  XOR U38877 ( .A(a[919]), .B(n42197), .Z(n37948) );
  NANDN U38878 ( .A(n37948), .B(n42173), .Z(n37909) );
  NANDN U38879 ( .A(n37907), .B(n42172), .Z(n37908) );
  NAND U38880 ( .A(n37909), .B(n37908), .Z(n37957) );
  NAND U38881 ( .A(b[7]), .B(a[915]), .Z(n37958) );
  XNOR U38882 ( .A(n37957), .B(n37958), .Z(n37960) );
  XOR U38883 ( .A(n37959), .B(n37960), .Z(n37966) );
  NANDN U38884 ( .A(n37910), .B(n42093), .Z(n37912) );
  XOR U38885 ( .A(n42134), .B(a[921]), .Z(n37951) );
  NANDN U38886 ( .A(n37951), .B(n42095), .Z(n37911) );
  NAND U38887 ( .A(n37912), .B(n37911), .Z(n37964) );
  NANDN U38888 ( .A(n37913), .B(n42231), .Z(n37915) );
  XOR U38889 ( .A(n238), .B(a[917]), .Z(n37954) );
  NANDN U38890 ( .A(n37954), .B(n42234), .Z(n37914) );
  AND U38891 ( .A(n37915), .B(n37914), .Z(n37963) );
  XNOR U38892 ( .A(n37964), .B(n37963), .Z(n37965) );
  XNOR U38893 ( .A(n37966), .B(n37965), .Z(n37970) );
  NANDN U38894 ( .A(n37917), .B(n37916), .Z(n37921) );
  NAND U38895 ( .A(n37919), .B(n37918), .Z(n37920) );
  AND U38896 ( .A(n37921), .B(n37920), .Z(n37969) );
  XOR U38897 ( .A(n37970), .B(n37969), .Z(n37971) );
  NANDN U38898 ( .A(n37923), .B(n37922), .Z(n37927) );
  NANDN U38899 ( .A(n37925), .B(n37924), .Z(n37926) );
  NAND U38900 ( .A(n37927), .B(n37926), .Z(n37972) );
  XOR U38901 ( .A(n37971), .B(n37972), .Z(n37939) );
  OR U38902 ( .A(n37929), .B(n37928), .Z(n37933) );
  NANDN U38903 ( .A(n37931), .B(n37930), .Z(n37932) );
  NAND U38904 ( .A(n37933), .B(n37932), .Z(n37940) );
  XNOR U38905 ( .A(n37939), .B(n37940), .Z(n37941) );
  XNOR U38906 ( .A(n37942), .B(n37941), .Z(n37975) );
  XNOR U38907 ( .A(n37975), .B(sreg[1939]), .Z(n37977) );
  NAND U38908 ( .A(n37934), .B(sreg[1938]), .Z(n37938) );
  OR U38909 ( .A(n37936), .B(n37935), .Z(n37937) );
  AND U38910 ( .A(n37938), .B(n37937), .Z(n37976) );
  XOR U38911 ( .A(n37977), .B(n37976), .Z(c[1939]) );
  NANDN U38912 ( .A(n37940), .B(n37939), .Z(n37944) );
  NAND U38913 ( .A(n37942), .B(n37941), .Z(n37943) );
  NAND U38914 ( .A(n37944), .B(n37943), .Z(n37983) );
  NAND U38915 ( .A(b[0]), .B(a[924]), .Z(n37945) );
  XNOR U38916 ( .A(b[1]), .B(n37945), .Z(n37947) );
  NAND U38917 ( .A(n147), .B(a[923]), .Z(n37946) );
  AND U38918 ( .A(n37947), .B(n37946), .Z(n38000) );
  XOR U38919 ( .A(a[920]), .B(n42197), .Z(n37989) );
  NANDN U38920 ( .A(n37989), .B(n42173), .Z(n37950) );
  NANDN U38921 ( .A(n37948), .B(n42172), .Z(n37949) );
  NAND U38922 ( .A(n37950), .B(n37949), .Z(n37998) );
  NAND U38923 ( .A(b[7]), .B(a[916]), .Z(n37999) );
  XNOR U38924 ( .A(n37998), .B(n37999), .Z(n38001) );
  XOR U38925 ( .A(n38000), .B(n38001), .Z(n38007) );
  NANDN U38926 ( .A(n37951), .B(n42093), .Z(n37953) );
  XOR U38927 ( .A(n42134), .B(a[922]), .Z(n37992) );
  NANDN U38928 ( .A(n37992), .B(n42095), .Z(n37952) );
  NAND U38929 ( .A(n37953), .B(n37952), .Z(n38005) );
  NANDN U38930 ( .A(n37954), .B(n42231), .Z(n37956) );
  XOR U38931 ( .A(n238), .B(a[918]), .Z(n37995) );
  NANDN U38932 ( .A(n37995), .B(n42234), .Z(n37955) );
  AND U38933 ( .A(n37956), .B(n37955), .Z(n38004) );
  XNOR U38934 ( .A(n38005), .B(n38004), .Z(n38006) );
  XNOR U38935 ( .A(n38007), .B(n38006), .Z(n38011) );
  NANDN U38936 ( .A(n37958), .B(n37957), .Z(n37962) );
  NAND U38937 ( .A(n37960), .B(n37959), .Z(n37961) );
  AND U38938 ( .A(n37962), .B(n37961), .Z(n38010) );
  XOR U38939 ( .A(n38011), .B(n38010), .Z(n38012) );
  NANDN U38940 ( .A(n37964), .B(n37963), .Z(n37968) );
  NANDN U38941 ( .A(n37966), .B(n37965), .Z(n37967) );
  NAND U38942 ( .A(n37968), .B(n37967), .Z(n38013) );
  XOR U38943 ( .A(n38012), .B(n38013), .Z(n37980) );
  OR U38944 ( .A(n37970), .B(n37969), .Z(n37974) );
  NANDN U38945 ( .A(n37972), .B(n37971), .Z(n37973) );
  NAND U38946 ( .A(n37974), .B(n37973), .Z(n37981) );
  XNOR U38947 ( .A(n37980), .B(n37981), .Z(n37982) );
  XNOR U38948 ( .A(n37983), .B(n37982), .Z(n38016) );
  XNOR U38949 ( .A(n38016), .B(sreg[1940]), .Z(n38018) );
  NAND U38950 ( .A(n37975), .B(sreg[1939]), .Z(n37979) );
  OR U38951 ( .A(n37977), .B(n37976), .Z(n37978) );
  AND U38952 ( .A(n37979), .B(n37978), .Z(n38017) );
  XOR U38953 ( .A(n38018), .B(n38017), .Z(c[1940]) );
  NANDN U38954 ( .A(n37981), .B(n37980), .Z(n37985) );
  NAND U38955 ( .A(n37983), .B(n37982), .Z(n37984) );
  NAND U38956 ( .A(n37985), .B(n37984), .Z(n38024) );
  NAND U38957 ( .A(b[0]), .B(a[925]), .Z(n37986) );
  XNOR U38958 ( .A(b[1]), .B(n37986), .Z(n37988) );
  NAND U38959 ( .A(n147), .B(a[924]), .Z(n37987) );
  AND U38960 ( .A(n37988), .B(n37987), .Z(n38041) );
  XOR U38961 ( .A(a[921]), .B(n42197), .Z(n38030) );
  NANDN U38962 ( .A(n38030), .B(n42173), .Z(n37991) );
  NANDN U38963 ( .A(n37989), .B(n42172), .Z(n37990) );
  NAND U38964 ( .A(n37991), .B(n37990), .Z(n38039) );
  NAND U38965 ( .A(b[7]), .B(a[917]), .Z(n38040) );
  XNOR U38966 ( .A(n38039), .B(n38040), .Z(n38042) );
  XOR U38967 ( .A(n38041), .B(n38042), .Z(n38048) );
  NANDN U38968 ( .A(n37992), .B(n42093), .Z(n37994) );
  XOR U38969 ( .A(n42134), .B(a[923]), .Z(n38033) );
  NANDN U38970 ( .A(n38033), .B(n42095), .Z(n37993) );
  NAND U38971 ( .A(n37994), .B(n37993), .Z(n38046) );
  NANDN U38972 ( .A(n37995), .B(n42231), .Z(n37997) );
  XOR U38973 ( .A(n238), .B(a[919]), .Z(n38036) );
  NANDN U38974 ( .A(n38036), .B(n42234), .Z(n37996) );
  AND U38975 ( .A(n37997), .B(n37996), .Z(n38045) );
  XNOR U38976 ( .A(n38046), .B(n38045), .Z(n38047) );
  XNOR U38977 ( .A(n38048), .B(n38047), .Z(n38052) );
  NANDN U38978 ( .A(n37999), .B(n37998), .Z(n38003) );
  NAND U38979 ( .A(n38001), .B(n38000), .Z(n38002) );
  AND U38980 ( .A(n38003), .B(n38002), .Z(n38051) );
  XOR U38981 ( .A(n38052), .B(n38051), .Z(n38053) );
  NANDN U38982 ( .A(n38005), .B(n38004), .Z(n38009) );
  NANDN U38983 ( .A(n38007), .B(n38006), .Z(n38008) );
  NAND U38984 ( .A(n38009), .B(n38008), .Z(n38054) );
  XOR U38985 ( .A(n38053), .B(n38054), .Z(n38021) );
  OR U38986 ( .A(n38011), .B(n38010), .Z(n38015) );
  NANDN U38987 ( .A(n38013), .B(n38012), .Z(n38014) );
  NAND U38988 ( .A(n38015), .B(n38014), .Z(n38022) );
  XNOR U38989 ( .A(n38021), .B(n38022), .Z(n38023) );
  XNOR U38990 ( .A(n38024), .B(n38023), .Z(n38057) );
  XNOR U38991 ( .A(n38057), .B(sreg[1941]), .Z(n38059) );
  NAND U38992 ( .A(n38016), .B(sreg[1940]), .Z(n38020) );
  OR U38993 ( .A(n38018), .B(n38017), .Z(n38019) );
  AND U38994 ( .A(n38020), .B(n38019), .Z(n38058) );
  XOR U38995 ( .A(n38059), .B(n38058), .Z(c[1941]) );
  NANDN U38996 ( .A(n38022), .B(n38021), .Z(n38026) );
  NAND U38997 ( .A(n38024), .B(n38023), .Z(n38025) );
  NAND U38998 ( .A(n38026), .B(n38025), .Z(n38065) );
  NAND U38999 ( .A(b[0]), .B(a[926]), .Z(n38027) );
  XNOR U39000 ( .A(b[1]), .B(n38027), .Z(n38029) );
  NAND U39001 ( .A(n147), .B(a[925]), .Z(n38028) );
  AND U39002 ( .A(n38029), .B(n38028), .Z(n38082) );
  XOR U39003 ( .A(a[922]), .B(n42197), .Z(n38071) );
  NANDN U39004 ( .A(n38071), .B(n42173), .Z(n38032) );
  NANDN U39005 ( .A(n38030), .B(n42172), .Z(n38031) );
  NAND U39006 ( .A(n38032), .B(n38031), .Z(n38080) );
  NAND U39007 ( .A(b[7]), .B(a[918]), .Z(n38081) );
  XNOR U39008 ( .A(n38080), .B(n38081), .Z(n38083) );
  XOR U39009 ( .A(n38082), .B(n38083), .Z(n38089) );
  NANDN U39010 ( .A(n38033), .B(n42093), .Z(n38035) );
  XOR U39011 ( .A(n42134), .B(a[924]), .Z(n38074) );
  NANDN U39012 ( .A(n38074), .B(n42095), .Z(n38034) );
  NAND U39013 ( .A(n38035), .B(n38034), .Z(n38087) );
  NANDN U39014 ( .A(n38036), .B(n42231), .Z(n38038) );
  XOR U39015 ( .A(n238), .B(a[920]), .Z(n38077) );
  NANDN U39016 ( .A(n38077), .B(n42234), .Z(n38037) );
  AND U39017 ( .A(n38038), .B(n38037), .Z(n38086) );
  XNOR U39018 ( .A(n38087), .B(n38086), .Z(n38088) );
  XNOR U39019 ( .A(n38089), .B(n38088), .Z(n38093) );
  NANDN U39020 ( .A(n38040), .B(n38039), .Z(n38044) );
  NAND U39021 ( .A(n38042), .B(n38041), .Z(n38043) );
  AND U39022 ( .A(n38044), .B(n38043), .Z(n38092) );
  XOR U39023 ( .A(n38093), .B(n38092), .Z(n38094) );
  NANDN U39024 ( .A(n38046), .B(n38045), .Z(n38050) );
  NANDN U39025 ( .A(n38048), .B(n38047), .Z(n38049) );
  NAND U39026 ( .A(n38050), .B(n38049), .Z(n38095) );
  XOR U39027 ( .A(n38094), .B(n38095), .Z(n38062) );
  OR U39028 ( .A(n38052), .B(n38051), .Z(n38056) );
  NANDN U39029 ( .A(n38054), .B(n38053), .Z(n38055) );
  NAND U39030 ( .A(n38056), .B(n38055), .Z(n38063) );
  XNOR U39031 ( .A(n38062), .B(n38063), .Z(n38064) );
  XNOR U39032 ( .A(n38065), .B(n38064), .Z(n38098) );
  XNOR U39033 ( .A(n38098), .B(sreg[1942]), .Z(n38100) );
  NAND U39034 ( .A(n38057), .B(sreg[1941]), .Z(n38061) );
  OR U39035 ( .A(n38059), .B(n38058), .Z(n38060) );
  AND U39036 ( .A(n38061), .B(n38060), .Z(n38099) );
  XOR U39037 ( .A(n38100), .B(n38099), .Z(c[1942]) );
  NANDN U39038 ( .A(n38063), .B(n38062), .Z(n38067) );
  NAND U39039 ( .A(n38065), .B(n38064), .Z(n38066) );
  NAND U39040 ( .A(n38067), .B(n38066), .Z(n38106) );
  NAND U39041 ( .A(b[0]), .B(a[927]), .Z(n38068) );
  XNOR U39042 ( .A(b[1]), .B(n38068), .Z(n38070) );
  NAND U39043 ( .A(n147), .B(a[926]), .Z(n38069) );
  AND U39044 ( .A(n38070), .B(n38069), .Z(n38123) );
  XOR U39045 ( .A(a[923]), .B(n42197), .Z(n38112) );
  NANDN U39046 ( .A(n38112), .B(n42173), .Z(n38073) );
  NANDN U39047 ( .A(n38071), .B(n42172), .Z(n38072) );
  NAND U39048 ( .A(n38073), .B(n38072), .Z(n38121) );
  NAND U39049 ( .A(b[7]), .B(a[919]), .Z(n38122) );
  XNOR U39050 ( .A(n38121), .B(n38122), .Z(n38124) );
  XOR U39051 ( .A(n38123), .B(n38124), .Z(n38130) );
  NANDN U39052 ( .A(n38074), .B(n42093), .Z(n38076) );
  XOR U39053 ( .A(n42134), .B(a[925]), .Z(n38115) );
  NANDN U39054 ( .A(n38115), .B(n42095), .Z(n38075) );
  NAND U39055 ( .A(n38076), .B(n38075), .Z(n38128) );
  NANDN U39056 ( .A(n38077), .B(n42231), .Z(n38079) );
  XOR U39057 ( .A(n238), .B(a[921]), .Z(n38118) );
  NANDN U39058 ( .A(n38118), .B(n42234), .Z(n38078) );
  AND U39059 ( .A(n38079), .B(n38078), .Z(n38127) );
  XNOR U39060 ( .A(n38128), .B(n38127), .Z(n38129) );
  XNOR U39061 ( .A(n38130), .B(n38129), .Z(n38134) );
  NANDN U39062 ( .A(n38081), .B(n38080), .Z(n38085) );
  NAND U39063 ( .A(n38083), .B(n38082), .Z(n38084) );
  AND U39064 ( .A(n38085), .B(n38084), .Z(n38133) );
  XOR U39065 ( .A(n38134), .B(n38133), .Z(n38135) );
  NANDN U39066 ( .A(n38087), .B(n38086), .Z(n38091) );
  NANDN U39067 ( .A(n38089), .B(n38088), .Z(n38090) );
  NAND U39068 ( .A(n38091), .B(n38090), .Z(n38136) );
  XOR U39069 ( .A(n38135), .B(n38136), .Z(n38103) );
  OR U39070 ( .A(n38093), .B(n38092), .Z(n38097) );
  NANDN U39071 ( .A(n38095), .B(n38094), .Z(n38096) );
  NAND U39072 ( .A(n38097), .B(n38096), .Z(n38104) );
  XNOR U39073 ( .A(n38103), .B(n38104), .Z(n38105) );
  XNOR U39074 ( .A(n38106), .B(n38105), .Z(n38139) );
  XNOR U39075 ( .A(n38139), .B(sreg[1943]), .Z(n38141) );
  NAND U39076 ( .A(n38098), .B(sreg[1942]), .Z(n38102) );
  OR U39077 ( .A(n38100), .B(n38099), .Z(n38101) );
  AND U39078 ( .A(n38102), .B(n38101), .Z(n38140) );
  XOR U39079 ( .A(n38141), .B(n38140), .Z(c[1943]) );
  NANDN U39080 ( .A(n38104), .B(n38103), .Z(n38108) );
  NAND U39081 ( .A(n38106), .B(n38105), .Z(n38107) );
  NAND U39082 ( .A(n38108), .B(n38107), .Z(n38147) );
  NAND U39083 ( .A(b[0]), .B(a[928]), .Z(n38109) );
  XNOR U39084 ( .A(b[1]), .B(n38109), .Z(n38111) );
  NAND U39085 ( .A(n147), .B(a[927]), .Z(n38110) );
  AND U39086 ( .A(n38111), .B(n38110), .Z(n38164) );
  XOR U39087 ( .A(a[924]), .B(n42197), .Z(n38153) );
  NANDN U39088 ( .A(n38153), .B(n42173), .Z(n38114) );
  NANDN U39089 ( .A(n38112), .B(n42172), .Z(n38113) );
  NAND U39090 ( .A(n38114), .B(n38113), .Z(n38162) );
  NAND U39091 ( .A(b[7]), .B(a[920]), .Z(n38163) );
  XNOR U39092 ( .A(n38162), .B(n38163), .Z(n38165) );
  XOR U39093 ( .A(n38164), .B(n38165), .Z(n38171) );
  NANDN U39094 ( .A(n38115), .B(n42093), .Z(n38117) );
  XOR U39095 ( .A(n42134), .B(a[926]), .Z(n38156) );
  NANDN U39096 ( .A(n38156), .B(n42095), .Z(n38116) );
  NAND U39097 ( .A(n38117), .B(n38116), .Z(n38169) );
  NANDN U39098 ( .A(n38118), .B(n42231), .Z(n38120) );
  XOR U39099 ( .A(n238), .B(a[922]), .Z(n38159) );
  NANDN U39100 ( .A(n38159), .B(n42234), .Z(n38119) );
  AND U39101 ( .A(n38120), .B(n38119), .Z(n38168) );
  XNOR U39102 ( .A(n38169), .B(n38168), .Z(n38170) );
  XNOR U39103 ( .A(n38171), .B(n38170), .Z(n38175) );
  NANDN U39104 ( .A(n38122), .B(n38121), .Z(n38126) );
  NAND U39105 ( .A(n38124), .B(n38123), .Z(n38125) );
  AND U39106 ( .A(n38126), .B(n38125), .Z(n38174) );
  XOR U39107 ( .A(n38175), .B(n38174), .Z(n38176) );
  NANDN U39108 ( .A(n38128), .B(n38127), .Z(n38132) );
  NANDN U39109 ( .A(n38130), .B(n38129), .Z(n38131) );
  NAND U39110 ( .A(n38132), .B(n38131), .Z(n38177) );
  XOR U39111 ( .A(n38176), .B(n38177), .Z(n38144) );
  OR U39112 ( .A(n38134), .B(n38133), .Z(n38138) );
  NANDN U39113 ( .A(n38136), .B(n38135), .Z(n38137) );
  NAND U39114 ( .A(n38138), .B(n38137), .Z(n38145) );
  XNOR U39115 ( .A(n38144), .B(n38145), .Z(n38146) );
  XNOR U39116 ( .A(n38147), .B(n38146), .Z(n38180) );
  XNOR U39117 ( .A(n38180), .B(sreg[1944]), .Z(n38182) );
  NAND U39118 ( .A(n38139), .B(sreg[1943]), .Z(n38143) );
  OR U39119 ( .A(n38141), .B(n38140), .Z(n38142) );
  AND U39120 ( .A(n38143), .B(n38142), .Z(n38181) );
  XOR U39121 ( .A(n38182), .B(n38181), .Z(c[1944]) );
  NANDN U39122 ( .A(n38145), .B(n38144), .Z(n38149) );
  NAND U39123 ( .A(n38147), .B(n38146), .Z(n38148) );
  NAND U39124 ( .A(n38149), .B(n38148), .Z(n38188) );
  NAND U39125 ( .A(b[0]), .B(a[929]), .Z(n38150) );
  XNOR U39126 ( .A(b[1]), .B(n38150), .Z(n38152) );
  NAND U39127 ( .A(n147), .B(a[928]), .Z(n38151) );
  AND U39128 ( .A(n38152), .B(n38151), .Z(n38205) );
  XOR U39129 ( .A(a[925]), .B(n42197), .Z(n38194) );
  NANDN U39130 ( .A(n38194), .B(n42173), .Z(n38155) );
  NANDN U39131 ( .A(n38153), .B(n42172), .Z(n38154) );
  NAND U39132 ( .A(n38155), .B(n38154), .Z(n38203) );
  NAND U39133 ( .A(b[7]), .B(a[921]), .Z(n38204) );
  XNOR U39134 ( .A(n38203), .B(n38204), .Z(n38206) );
  XOR U39135 ( .A(n38205), .B(n38206), .Z(n38212) );
  NANDN U39136 ( .A(n38156), .B(n42093), .Z(n38158) );
  XOR U39137 ( .A(n42134), .B(a[927]), .Z(n38197) );
  NANDN U39138 ( .A(n38197), .B(n42095), .Z(n38157) );
  NAND U39139 ( .A(n38158), .B(n38157), .Z(n38210) );
  NANDN U39140 ( .A(n38159), .B(n42231), .Z(n38161) );
  XOR U39141 ( .A(n239), .B(a[923]), .Z(n38200) );
  NANDN U39142 ( .A(n38200), .B(n42234), .Z(n38160) );
  AND U39143 ( .A(n38161), .B(n38160), .Z(n38209) );
  XNOR U39144 ( .A(n38210), .B(n38209), .Z(n38211) );
  XNOR U39145 ( .A(n38212), .B(n38211), .Z(n38216) );
  NANDN U39146 ( .A(n38163), .B(n38162), .Z(n38167) );
  NAND U39147 ( .A(n38165), .B(n38164), .Z(n38166) );
  AND U39148 ( .A(n38167), .B(n38166), .Z(n38215) );
  XOR U39149 ( .A(n38216), .B(n38215), .Z(n38217) );
  NANDN U39150 ( .A(n38169), .B(n38168), .Z(n38173) );
  NANDN U39151 ( .A(n38171), .B(n38170), .Z(n38172) );
  NAND U39152 ( .A(n38173), .B(n38172), .Z(n38218) );
  XOR U39153 ( .A(n38217), .B(n38218), .Z(n38185) );
  OR U39154 ( .A(n38175), .B(n38174), .Z(n38179) );
  NANDN U39155 ( .A(n38177), .B(n38176), .Z(n38178) );
  NAND U39156 ( .A(n38179), .B(n38178), .Z(n38186) );
  XNOR U39157 ( .A(n38185), .B(n38186), .Z(n38187) );
  XNOR U39158 ( .A(n38188), .B(n38187), .Z(n38221) );
  XNOR U39159 ( .A(n38221), .B(sreg[1945]), .Z(n38223) );
  NAND U39160 ( .A(n38180), .B(sreg[1944]), .Z(n38184) );
  OR U39161 ( .A(n38182), .B(n38181), .Z(n38183) );
  AND U39162 ( .A(n38184), .B(n38183), .Z(n38222) );
  XOR U39163 ( .A(n38223), .B(n38222), .Z(c[1945]) );
  NANDN U39164 ( .A(n38186), .B(n38185), .Z(n38190) );
  NAND U39165 ( .A(n38188), .B(n38187), .Z(n38189) );
  NAND U39166 ( .A(n38190), .B(n38189), .Z(n38229) );
  NAND U39167 ( .A(b[0]), .B(a[930]), .Z(n38191) );
  XNOR U39168 ( .A(b[1]), .B(n38191), .Z(n38193) );
  NAND U39169 ( .A(n147), .B(a[929]), .Z(n38192) );
  AND U39170 ( .A(n38193), .B(n38192), .Z(n38246) );
  XOR U39171 ( .A(a[926]), .B(n42197), .Z(n38235) );
  NANDN U39172 ( .A(n38235), .B(n42173), .Z(n38196) );
  NANDN U39173 ( .A(n38194), .B(n42172), .Z(n38195) );
  NAND U39174 ( .A(n38196), .B(n38195), .Z(n38244) );
  NAND U39175 ( .A(b[7]), .B(a[922]), .Z(n38245) );
  XNOR U39176 ( .A(n38244), .B(n38245), .Z(n38247) );
  XOR U39177 ( .A(n38246), .B(n38247), .Z(n38253) );
  NANDN U39178 ( .A(n38197), .B(n42093), .Z(n38199) );
  XOR U39179 ( .A(n42134), .B(a[928]), .Z(n38238) );
  NANDN U39180 ( .A(n38238), .B(n42095), .Z(n38198) );
  NAND U39181 ( .A(n38199), .B(n38198), .Z(n38251) );
  NANDN U39182 ( .A(n38200), .B(n42231), .Z(n38202) );
  XOR U39183 ( .A(n239), .B(a[924]), .Z(n38241) );
  NANDN U39184 ( .A(n38241), .B(n42234), .Z(n38201) );
  AND U39185 ( .A(n38202), .B(n38201), .Z(n38250) );
  XNOR U39186 ( .A(n38251), .B(n38250), .Z(n38252) );
  XNOR U39187 ( .A(n38253), .B(n38252), .Z(n38257) );
  NANDN U39188 ( .A(n38204), .B(n38203), .Z(n38208) );
  NAND U39189 ( .A(n38206), .B(n38205), .Z(n38207) );
  AND U39190 ( .A(n38208), .B(n38207), .Z(n38256) );
  XOR U39191 ( .A(n38257), .B(n38256), .Z(n38258) );
  NANDN U39192 ( .A(n38210), .B(n38209), .Z(n38214) );
  NANDN U39193 ( .A(n38212), .B(n38211), .Z(n38213) );
  NAND U39194 ( .A(n38214), .B(n38213), .Z(n38259) );
  XOR U39195 ( .A(n38258), .B(n38259), .Z(n38226) );
  OR U39196 ( .A(n38216), .B(n38215), .Z(n38220) );
  NANDN U39197 ( .A(n38218), .B(n38217), .Z(n38219) );
  NAND U39198 ( .A(n38220), .B(n38219), .Z(n38227) );
  XNOR U39199 ( .A(n38226), .B(n38227), .Z(n38228) );
  XNOR U39200 ( .A(n38229), .B(n38228), .Z(n38262) );
  XNOR U39201 ( .A(n38262), .B(sreg[1946]), .Z(n38264) );
  NAND U39202 ( .A(n38221), .B(sreg[1945]), .Z(n38225) );
  OR U39203 ( .A(n38223), .B(n38222), .Z(n38224) );
  AND U39204 ( .A(n38225), .B(n38224), .Z(n38263) );
  XOR U39205 ( .A(n38264), .B(n38263), .Z(c[1946]) );
  NANDN U39206 ( .A(n38227), .B(n38226), .Z(n38231) );
  NAND U39207 ( .A(n38229), .B(n38228), .Z(n38230) );
  NAND U39208 ( .A(n38231), .B(n38230), .Z(n38270) );
  NAND U39209 ( .A(b[0]), .B(a[931]), .Z(n38232) );
  XNOR U39210 ( .A(b[1]), .B(n38232), .Z(n38234) );
  NAND U39211 ( .A(n148), .B(a[930]), .Z(n38233) );
  AND U39212 ( .A(n38234), .B(n38233), .Z(n38287) );
  XOR U39213 ( .A(a[927]), .B(n42197), .Z(n38276) );
  NANDN U39214 ( .A(n38276), .B(n42173), .Z(n38237) );
  NANDN U39215 ( .A(n38235), .B(n42172), .Z(n38236) );
  NAND U39216 ( .A(n38237), .B(n38236), .Z(n38285) );
  NAND U39217 ( .A(b[7]), .B(a[923]), .Z(n38286) );
  XNOR U39218 ( .A(n38285), .B(n38286), .Z(n38288) );
  XOR U39219 ( .A(n38287), .B(n38288), .Z(n38294) );
  NANDN U39220 ( .A(n38238), .B(n42093), .Z(n38240) );
  XOR U39221 ( .A(n42134), .B(a[929]), .Z(n38279) );
  NANDN U39222 ( .A(n38279), .B(n42095), .Z(n38239) );
  NAND U39223 ( .A(n38240), .B(n38239), .Z(n38292) );
  NANDN U39224 ( .A(n38241), .B(n42231), .Z(n38243) );
  XOR U39225 ( .A(n239), .B(a[925]), .Z(n38282) );
  NANDN U39226 ( .A(n38282), .B(n42234), .Z(n38242) );
  AND U39227 ( .A(n38243), .B(n38242), .Z(n38291) );
  XNOR U39228 ( .A(n38292), .B(n38291), .Z(n38293) );
  XNOR U39229 ( .A(n38294), .B(n38293), .Z(n38298) );
  NANDN U39230 ( .A(n38245), .B(n38244), .Z(n38249) );
  NAND U39231 ( .A(n38247), .B(n38246), .Z(n38248) );
  AND U39232 ( .A(n38249), .B(n38248), .Z(n38297) );
  XOR U39233 ( .A(n38298), .B(n38297), .Z(n38299) );
  NANDN U39234 ( .A(n38251), .B(n38250), .Z(n38255) );
  NANDN U39235 ( .A(n38253), .B(n38252), .Z(n38254) );
  NAND U39236 ( .A(n38255), .B(n38254), .Z(n38300) );
  XOR U39237 ( .A(n38299), .B(n38300), .Z(n38267) );
  OR U39238 ( .A(n38257), .B(n38256), .Z(n38261) );
  NANDN U39239 ( .A(n38259), .B(n38258), .Z(n38260) );
  NAND U39240 ( .A(n38261), .B(n38260), .Z(n38268) );
  XNOR U39241 ( .A(n38267), .B(n38268), .Z(n38269) );
  XNOR U39242 ( .A(n38270), .B(n38269), .Z(n38303) );
  XNOR U39243 ( .A(n38303), .B(sreg[1947]), .Z(n38305) );
  NAND U39244 ( .A(n38262), .B(sreg[1946]), .Z(n38266) );
  OR U39245 ( .A(n38264), .B(n38263), .Z(n38265) );
  AND U39246 ( .A(n38266), .B(n38265), .Z(n38304) );
  XOR U39247 ( .A(n38305), .B(n38304), .Z(c[1947]) );
  NANDN U39248 ( .A(n38268), .B(n38267), .Z(n38272) );
  NAND U39249 ( .A(n38270), .B(n38269), .Z(n38271) );
  NAND U39250 ( .A(n38272), .B(n38271), .Z(n38311) );
  NAND U39251 ( .A(b[0]), .B(a[932]), .Z(n38273) );
  XNOR U39252 ( .A(b[1]), .B(n38273), .Z(n38275) );
  NAND U39253 ( .A(n148), .B(a[931]), .Z(n38274) );
  AND U39254 ( .A(n38275), .B(n38274), .Z(n38328) );
  XOR U39255 ( .A(a[928]), .B(n42197), .Z(n38317) );
  NANDN U39256 ( .A(n38317), .B(n42173), .Z(n38278) );
  NANDN U39257 ( .A(n38276), .B(n42172), .Z(n38277) );
  NAND U39258 ( .A(n38278), .B(n38277), .Z(n38326) );
  NAND U39259 ( .A(b[7]), .B(a[924]), .Z(n38327) );
  XNOR U39260 ( .A(n38326), .B(n38327), .Z(n38329) );
  XOR U39261 ( .A(n38328), .B(n38329), .Z(n38335) );
  NANDN U39262 ( .A(n38279), .B(n42093), .Z(n38281) );
  XOR U39263 ( .A(n42134), .B(a[930]), .Z(n38320) );
  NANDN U39264 ( .A(n38320), .B(n42095), .Z(n38280) );
  NAND U39265 ( .A(n38281), .B(n38280), .Z(n38333) );
  NANDN U39266 ( .A(n38282), .B(n42231), .Z(n38284) );
  XOR U39267 ( .A(n239), .B(a[926]), .Z(n38323) );
  NANDN U39268 ( .A(n38323), .B(n42234), .Z(n38283) );
  AND U39269 ( .A(n38284), .B(n38283), .Z(n38332) );
  XNOR U39270 ( .A(n38333), .B(n38332), .Z(n38334) );
  XNOR U39271 ( .A(n38335), .B(n38334), .Z(n38339) );
  NANDN U39272 ( .A(n38286), .B(n38285), .Z(n38290) );
  NAND U39273 ( .A(n38288), .B(n38287), .Z(n38289) );
  AND U39274 ( .A(n38290), .B(n38289), .Z(n38338) );
  XOR U39275 ( .A(n38339), .B(n38338), .Z(n38340) );
  NANDN U39276 ( .A(n38292), .B(n38291), .Z(n38296) );
  NANDN U39277 ( .A(n38294), .B(n38293), .Z(n38295) );
  NAND U39278 ( .A(n38296), .B(n38295), .Z(n38341) );
  XOR U39279 ( .A(n38340), .B(n38341), .Z(n38308) );
  OR U39280 ( .A(n38298), .B(n38297), .Z(n38302) );
  NANDN U39281 ( .A(n38300), .B(n38299), .Z(n38301) );
  NAND U39282 ( .A(n38302), .B(n38301), .Z(n38309) );
  XNOR U39283 ( .A(n38308), .B(n38309), .Z(n38310) );
  XNOR U39284 ( .A(n38311), .B(n38310), .Z(n38344) );
  XNOR U39285 ( .A(n38344), .B(sreg[1948]), .Z(n38346) );
  NAND U39286 ( .A(n38303), .B(sreg[1947]), .Z(n38307) );
  OR U39287 ( .A(n38305), .B(n38304), .Z(n38306) );
  AND U39288 ( .A(n38307), .B(n38306), .Z(n38345) );
  XOR U39289 ( .A(n38346), .B(n38345), .Z(c[1948]) );
  NANDN U39290 ( .A(n38309), .B(n38308), .Z(n38313) );
  NAND U39291 ( .A(n38311), .B(n38310), .Z(n38312) );
  NAND U39292 ( .A(n38313), .B(n38312), .Z(n38352) );
  NAND U39293 ( .A(b[0]), .B(a[933]), .Z(n38314) );
  XNOR U39294 ( .A(b[1]), .B(n38314), .Z(n38316) );
  NAND U39295 ( .A(n148), .B(a[932]), .Z(n38315) );
  AND U39296 ( .A(n38316), .B(n38315), .Z(n38369) );
  XOR U39297 ( .A(a[929]), .B(n42197), .Z(n38358) );
  NANDN U39298 ( .A(n38358), .B(n42173), .Z(n38319) );
  NANDN U39299 ( .A(n38317), .B(n42172), .Z(n38318) );
  NAND U39300 ( .A(n38319), .B(n38318), .Z(n38367) );
  NAND U39301 ( .A(b[7]), .B(a[925]), .Z(n38368) );
  XNOR U39302 ( .A(n38367), .B(n38368), .Z(n38370) );
  XOR U39303 ( .A(n38369), .B(n38370), .Z(n38376) );
  NANDN U39304 ( .A(n38320), .B(n42093), .Z(n38322) );
  XOR U39305 ( .A(n42134), .B(a[931]), .Z(n38361) );
  NANDN U39306 ( .A(n38361), .B(n42095), .Z(n38321) );
  NAND U39307 ( .A(n38322), .B(n38321), .Z(n38374) );
  NANDN U39308 ( .A(n38323), .B(n42231), .Z(n38325) );
  XOR U39309 ( .A(n239), .B(a[927]), .Z(n38364) );
  NANDN U39310 ( .A(n38364), .B(n42234), .Z(n38324) );
  AND U39311 ( .A(n38325), .B(n38324), .Z(n38373) );
  XNOR U39312 ( .A(n38374), .B(n38373), .Z(n38375) );
  XNOR U39313 ( .A(n38376), .B(n38375), .Z(n38380) );
  NANDN U39314 ( .A(n38327), .B(n38326), .Z(n38331) );
  NAND U39315 ( .A(n38329), .B(n38328), .Z(n38330) );
  AND U39316 ( .A(n38331), .B(n38330), .Z(n38379) );
  XOR U39317 ( .A(n38380), .B(n38379), .Z(n38381) );
  NANDN U39318 ( .A(n38333), .B(n38332), .Z(n38337) );
  NANDN U39319 ( .A(n38335), .B(n38334), .Z(n38336) );
  NAND U39320 ( .A(n38337), .B(n38336), .Z(n38382) );
  XOR U39321 ( .A(n38381), .B(n38382), .Z(n38349) );
  OR U39322 ( .A(n38339), .B(n38338), .Z(n38343) );
  NANDN U39323 ( .A(n38341), .B(n38340), .Z(n38342) );
  NAND U39324 ( .A(n38343), .B(n38342), .Z(n38350) );
  XNOR U39325 ( .A(n38349), .B(n38350), .Z(n38351) );
  XNOR U39326 ( .A(n38352), .B(n38351), .Z(n38385) );
  XNOR U39327 ( .A(n38385), .B(sreg[1949]), .Z(n38387) );
  NAND U39328 ( .A(n38344), .B(sreg[1948]), .Z(n38348) );
  OR U39329 ( .A(n38346), .B(n38345), .Z(n38347) );
  AND U39330 ( .A(n38348), .B(n38347), .Z(n38386) );
  XOR U39331 ( .A(n38387), .B(n38386), .Z(c[1949]) );
  NANDN U39332 ( .A(n38350), .B(n38349), .Z(n38354) );
  NAND U39333 ( .A(n38352), .B(n38351), .Z(n38353) );
  NAND U39334 ( .A(n38354), .B(n38353), .Z(n38393) );
  NAND U39335 ( .A(b[0]), .B(a[934]), .Z(n38355) );
  XNOR U39336 ( .A(b[1]), .B(n38355), .Z(n38357) );
  NAND U39337 ( .A(n148), .B(a[933]), .Z(n38356) );
  AND U39338 ( .A(n38357), .B(n38356), .Z(n38410) );
  XOR U39339 ( .A(a[930]), .B(n42197), .Z(n38399) );
  NANDN U39340 ( .A(n38399), .B(n42173), .Z(n38360) );
  NANDN U39341 ( .A(n38358), .B(n42172), .Z(n38359) );
  NAND U39342 ( .A(n38360), .B(n38359), .Z(n38408) );
  NAND U39343 ( .A(b[7]), .B(a[926]), .Z(n38409) );
  XNOR U39344 ( .A(n38408), .B(n38409), .Z(n38411) );
  XOR U39345 ( .A(n38410), .B(n38411), .Z(n38417) );
  NANDN U39346 ( .A(n38361), .B(n42093), .Z(n38363) );
  XOR U39347 ( .A(n42134), .B(a[932]), .Z(n38402) );
  NANDN U39348 ( .A(n38402), .B(n42095), .Z(n38362) );
  NAND U39349 ( .A(n38363), .B(n38362), .Z(n38415) );
  NANDN U39350 ( .A(n38364), .B(n42231), .Z(n38366) );
  XOR U39351 ( .A(n239), .B(a[928]), .Z(n38405) );
  NANDN U39352 ( .A(n38405), .B(n42234), .Z(n38365) );
  AND U39353 ( .A(n38366), .B(n38365), .Z(n38414) );
  XNOR U39354 ( .A(n38415), .B(n38414), .Z(n38416) );
  XNOR U39355 ( .A(n38417), .B(n38416), .Z(n38421) );
  NANDN U39356 ( .A(n38368), .B(n38367), .Z(n38372) );
  NAND U39357 ( .A(n38370), .B(n38369), .Z(n38371) );
  AND U39358 ( .A(n38372), .B(n38371), .Z(n38420) );
  XOR U39359 ( .A(n38421), .B(n38420), .Z(n38422) );
  NANDN U39360 ( .A(n38374), .B(n38373), .Z(n38378) );
  NANDN U39361 ( .A(n38376), .B(n38375), .Z(n38377) );
  NAND U39362 ( .A(n38378), .B(n38377), .Z(n38423) );
  XOR U39363 ( .A(n38422), .B(n38423), .Z(n38390) );
  OR U39364 ( .A(n38380), .B(n38379), .Z(n38384) );
  NANDN U39365 ( .A(n38382), .B(n38381), .Z(n38383) );
  NAND U39366 ( .A(n38384), .B(n38383), .Z(n38391) );
  XNOR U39367 ( .A(n38390), .B(n38391), .Z(n38392) );
  XNOR U39368 ( .A(n38393), .B(n38392), .Z(n38426) );
  XNOR U39369 ( .A(n38426), .B(sreg[1950]), .Z(n38428) );
  NAND U39370 ( .A(n38385), .B(sreg[1949]), .Z(n38389) );
  OR U39371 ( .A(n38387), .B(n38386), .Z(n38388) );
  AND U39372 ( .A(n38389), .B(n38388), .Z(n38427) );
  XOR U39373 ( .A(n38428), .B(n38427), .Z(c[1950]) );
  NANDN U39374 ( .A(n38391), .B(n38390), .Z(n38395) );
  NAND U39375 ( .A(n38393), .B(n38392), .Z(n38394) );
  NAND U39376 ( .A(n38395), .B(n38394), .Z(n38434) );
  NAND U39377 ( .A(b[0]), .B(a[935]), .Z(n38396) );
  XNOR U39378 ( .A(b[1]), .B(n38396), .Z(n38398) );
  NAND U39379 ( .A(n148), .B(a[934]), .Z(n38397) );
  AND U39380 ( .A(n38398), .B(n38397), .Z(n38451) );
  XOR U39381 ( .A(a[931]), .B(n42197), .Z(n38440) );
  NANDN U39382 ( .A(n38440), .B(n42173), .Z(n38401) );
  NANDN U39383 ( .A(n38399), .B(n42172), .Z(n38400) );
  NAND U39384 ( .A(n38401), .B(n38400), .Z(n38449) );
  NAND U39385 ( .A(b[7]), .B(a[927]), .Z(n38450) );
  XNOR U39386 ( .A(n38449), .B(n38450), .Z(n38452) );
  XOR U39387 ( .A(n38451), .B(n38452), .Z(n38458) );
  NANDN U39388 ( .A(n38402), .B(n42093), .Z(n38404) );
  XOR U39389 ( .A(n42134), .B(a[933]), .Z(n38443) );
  NANDN U39390 ( .A(n38443), .B(n42095), .Z(n38403) );
  NAND U39391 ( .A(n38404), .B(n38403), .Z(n38456) );
  NANDN U39392 ( .A(n38405), .B(n42231), .Z(n38407) );
  XOR U39393 ( .A(n239), .B(a[929]), .Z(n38446) );
  NANDN U39394 ( .A(n38446), .B(n42234), .Z(n38406) );
  AND U39395 ( .A(n38407), .B(n38406), .Z(n38455) );
  XNOR U39396 ( .A(n38456), .B(n38455), .Z(n38457) );
  XNOR U39397 ( .A(n38458), .B(n38457), .Z(n38462) );
  NANDN U39398 ( .A(n38409), .B(n38408), .Z(n38413) );
  NAND U39399 ( .A(n38411), .B(n38410), .Z(n38412) );
  AND U39400 ( .A(n38413), .B(n38412), .Z(n38461) );
  XOR U39401 ( .A(n38462), .B(n38461), .Z(n38463) );
  NANDN U39402 ( .A(n38415), .B(n38414), .Z(n38419) );
  NANDN U39403 ( .A(n38417), .B(n38416), .Z(n38418) );
  NAND U39404 ( .A(n38419), .B(n38418), .Z(n38464) );
  XOR U39405 ( .A(n38463), .B(n38464), .Z(n38431) );
  OR U39406 ( .A(n38421), .B(n38420), .Z(n38425) );
  NANDN U39407 ( .A(n38423), .B(n38422), .Z(n38424) );
  NAND U39408 ( .A(n38425), .B(n38424), .Z(n38432) );
  XNOR U39409 ( .A(n38431), .B(n38432), .Z(n38433) );
  XNOR U39410 ( .A(n38434), .B(n38433), .Z(n38467) );
  XNOR U39411 ( .A(n38467), .B(sreg[1951]), .Z(n38469) );
  NAND U39412 ( .A(n38426), .B(sreg[1950]), .Z(n38430) );
  OR U39413 ( .A(n38428), .B(n38427), .Z(n38429) );
  AND U39414 ( .A(n38430), .B(n38429), .Z(n38468) );
  XOR U39415 ( .A(n38469), .B(n38468), .Z(c[1951]) );
  NANDN U39416 ( .A(n38432), .B(n38431), .Z(n38436) );
  NAND U39417 ( .A(n38434), .B(n38433), .Z(n38435) );
  NAND U39418 ( .A(n38436), .B(n38435), .Z(n38475) );
  NAND U39419 ( .A(b[0]), .B(a[936]), .Z(n38437) );
  XNOR U39420 ( .A(b[1]), .B(n38437), .Z(n38439) );
  NAND U39421 ( .A(n148), .B(a[935]), .Z(n38438) );
  AND U39422 ( .A(n38439), .B(n38438), .Z(n38492) );
  XOR U39423 ( .A(a[932]), .B(n42197), .Z(n38481) );
  NANDN U39424 ( .A(n38481), .B(n42173), .Z(n38442) );
  NANDN U39425 ( .A(n38440), .B(n42172), .Z(n38441) );
  NAND U39426 ( .A(n38442), .B(n38441), .Z(n38490) );
  NAND U39427 ( .A(b[7]), .B(a[928]), .Z(n38491) );
  XNOR U39428 ( .A(n38490), .B(n38491), .Z(n38493) );
  XOR U39429 ( .A(n38492), .B(n38493), .Z(n38499) );
  NANDN U39430 ( .A(n38443), .B(n42093), .Z(n38445) );
  XOR U39431 ( .A(n42134), .B(a[934]), .Z(n38484) );
  NANDN U39432 ( .A(n38484), .B(n42095), .Z(n38444) );
  NAND U39433 ( .A(n38445), .B(n38444), .Z(n38497) );
  NANDN U39434 ( .A(n38446), .B(n42231), .Z(n38448) );
  XOR U39435 ( .A(n239), .B(a[930]), .Z(n38487) );
  NANDN U39436 ( .A(n38487), .B(n42234), .Z(n38447) );
  AND U39437 ( .A(n38448), .B(n38447), .Z(n38496) );
  XNOR U39438 ( .A(n38497), .B(n38496), .Z(n38498) );
  XNOR U39439 ( .A(n38499), .B(n38498), .Z(n38503) );
  NANDN U39440 ( .A(n38450), .B(n38449), .Z(n38454) );
  NAND U39441 ( .A(n38452), .B(n38451), .Z(n38453) );
  AND U39442 ( .A(n38454), .B(n38453), .Z(n38502) );
  XOR U39443 ( .A(n38503), .B(n38502), .Z(n38504) );
  NANDN U39444 ( .A(n38456), .B(n38455), .Z(n38460) );
  NANDN U39445 ( .A(n38458), .B(n38457), .Z(n38459) );
  NAND U39446 ( .A(n38460), .B(n38459), .Z(n38505) );
  XOR U39447 ( .A(n38504), .B(n38505), .Z(n38472) );
  OR U39448 ( .A(n38462), .B(n38461), .Z(n38466) );
  NANDN U39449 ( .A(n38464), .B(n38463), .Z(n38465) );
  NAND U39450 ( .A(n38466), .B(n38465), .Z(n38473) );
  XNOR U39451 ( .A(n38472), .B(n38473), .Z(n38474) );
  XNOR U39452 ( .A(n38475), .B(n38474), .Z(n38508) );
  XNOR U39453 ( .A(n38508), .B(sreg[1952]), .Z(n38510) );
  NAND U39454 ( .A(n38467), .B(sreg[1951]), .Z(n38471) );
  OR U39455 ( .A(n38469), .B(n38468), .Z(n38470) );
  AND U39456 ( .A(n38471), .B(n38470), .Z(n38509) );
  XOR U39457 ( .A(n38510), .B(n38509), .Z(c[1952]) );
  NANDN U39458 ( .A(n38473), .B(n38472), .Z(n38477) );
  NAND U39459 ( .A(n38475), .B(n38474), .Z(n38476) );
  NAND U39460 ( .A(n38477), .B(n38476), .Z(n38516) );
  NAND U39461 ( .A(b[0]), .B(a[937]), .Z(n38478) );
  XNOR U39462 ( .A(b[1]), .B(n38478), .Z(n38480) );
  NAND U39463 ( .A(n148), .B(a[936]), .Z(n38479) );
  AND U39464 ( .A(n38480), .B(n38479), .Z(n38533) );
  XOR U39465 ( .A(a[933]), .B(n42197), .Z(n38522) );
  NANDN U39466 ( .A(n38522), .B(n42173), .Z(n38483) );
  NANDN U39467 ( .A(n38481), .B(n42172), .Z(n38482) );
  NAND U39468 ( .A(n38483), .B(n38482), .Z(n38531) );
  NAND U39469 ( .A(b[7]), .B(a[929]), .Z(n38532) );
  XNOR U39470 ( .A(n38531), .B(n38532), .Z(n38534) );
  XOR U39471 ( .A(n38533), .B(n38534), .Z(n38540) );
  NANDN U39472 ( .A(n38484), .B(n42093), .Z(n38486) );
  XOR U39473 ( .A(n42134), .B(a[935]), .Z(n38525) );
  NANDN U39474 ( .A(n38525), .B(n42095), .Z(n38485) );
  NAND U39475 ( .A(n38486), .B(n38485), .Z(n38538) );
  NANDN U39476 ( .A(n38487), .B(n42231), .Z(n38489) );
  XOR U39477 ( .A(n239), .B(a[931]), .Z(n38528) );
  NANDN U39478 ( .A(n38528), .B(n42234), .Z(n38488) );
  AND U39479 ( .A(n38489), .B(n38488), .Z(n38537) );
  XNOR U39480 ( .A(n38538), .B(n38537), .Z(n38539) );
  XNOR U39481 ( .A(n38540), .B(n38539), .Z(n38544) );
  NANDN U39482 ( .A(n38491), .B(n38490), .Z(n38495) );
  NAND U39483 ( .A(n38493), .B(n38492), .Z(n38494) );
  AND U39484 ( .A(n38495), .B(n38494), .Z(n38543) );
  XOR U39485 ( .A(n38544), .B(n38543), .Z(n38545) );
  NANDN U39486 ( .A(n38497), .B(n38496), .Z(n38501) );
  NANDN U39487 ( .A(n38499), .B(n38498), .Z(n38500) );
  NAND U39488 ( .A(n38501), .B(n38500), .Z(n38546) );
  XOR U39489 ( .A(n38545), .B(n38546), .Z(n38513) );
  OR U39490 ( .A(n38503), .B(n38502), .Z(n38507) );
  NANDN U39491 ( .A(n38505), .B(n38504), .Z(n38506) );
  NAND U39492 ( .A(n38507), .B(n38506), .Z(n38514) );
  XNOR U39493 ( .A(n38513), .B(n38514), .Z(n38515) );
  XNOR U39494 ( .A(n38516), .B(n38515), .Z(n38549) );
  XNOR U39495 ( .A(n38549), .B(sreg[1953]), .Z(n38551) );
  NAND U39496 ( .A(n38508), .B(sreg[1952]), .Z(n38512) );
  OR U39497 ( .A(n38510), .B(n38509), .Z(n38511) );
  AND U39498 ( .A(n38512), .B(n38511), .Z(n38550) );
  XOR U39499 ( .A(n38551), .B(n38550), .Z(c[1953]) );
  NANDN U39500 ( .A(n38514), .B(n38513), .Z(n38518) );
  NAND U39501 ( .A(n38516), .B(n38515), .Z(n38517) );
  NAND U39502 ( .A(n38518), .B(n38517), .Z(n38557) );
  NAND U39503 ( .A(b[0]), .B(a[938]), .Z(n38519) );
  XNOR U39504 ( .A(b[1]), .B(n38519), .Z(n38521) );
  NAND U39505 ( .A(n149), .B(a[937]), .Z(n38520) );
  AND U39506 ( .A(n38521), .B(n38520), .Z(n38574) );
  XOR U39507 ( .A(a[934]), .B(n42197), .Z(n38563) );
  NANDN U39508 ( .A(n38563), .B(n42173), .Z(n38524) );
  NANDN U39509 ( .A(n38522), .B(n42172), .Z(n38523) );
  NAND U39510 ( .A(n38524), .B(n38523), .Z(n38572) );
  NAND U39511 ( .A(b[7]), .B(a[930]), .Z(n38573) );
  XNOR U39512 ( .A(n38572), .B(n38573), .Z(n38575) );
  XOR U39513 ( .A(n38574), .B(n38575), .Z(n38581) );
  NANDN U39514 ( .A(n38525), .B(n42093), .Z(n38527) );
  XOR U39515 ( .A(n42134), .B(a[936]), .Z(n38566) );
  NANDN U39516 ( .A(n38566), .B(n42095), .Z(n38526) );
  NAND U39517 ( .A(n38527), .B(n38526), .Z(n38579) );
  NANDN U39518 ( .A(n38528), .B(n42231), .Z(n38530) );
  XOR U39519 ( .A(n239), .B(a[932]), .Z(n38569) );
  NANDN U39520 ( .A(n38569), .B(n42234), .Z(n38529) );
  AND U39521 ( .A(n38530), .B(n38529), .Z(n38578) );
  XNOR U39522 ( .A(n38579), .B(n38578), .Z(n38580) );
  XNOR U39523 ( .A(n38581), .B(n38580), .Z(n38585) );
  NANDN U39524 ( .A(n38532), .B(n38531), .Z(n38536) );
  NAND U39525 ( .A(n38534), .B(n38533), .Z(n38535) );
  AND U39526 ( .A(n38536), .B(n38535), .Z(n38584) );
  XOR U39527 ( .A(n38585), .B(n38584), .Z(n38586) );
  NANDN U39528 ( .A(n38538), .B(n38537), .Z(n38542) );
  NANDN U39529 ( .A(n38540), .B(n38539), .Z(n38541) );
  NAND U39530 ( .A(n38542), .B(n38541), .Z(n38587) );
  XOR U39531 ( .A(n38586), .B(n38587), .Z(n38554) );
  OR U39532 ( .A(n38544), .B(n38543), .Z(n38548) );
  NANDN U39533 ( .A(n38546), .B(n38545), .Z(n38547) );
  NAND U39534 ( .A(n38548), .B(n38547), .Z(n38555) );
  XNOR U39535 ( .A(n38554), .B(n38555), .Z(n38556) );
  XNOR U39536 ( .A(n38557), .B(n38556), .Z(n38590) );
  XNOR U39537 ( .A(n38590), .B(sreg[1954]), .Z(n38592) );
  NAND U39538 ( .A(n38549), .B(sreg[1953]), .Z(n38553) );
  OR U39539 ( .A(n38551), .B(n38550), .Z(n38552) );
  AND U39540 ( .A(n38553), .B(n38552), .Z(n38591) );
  XOR U39541 ( .A(n38592), .B(n38591), .Z(c[1954]) );
  NANDN U39542 ( .A(n38555), .B(n38554), .Z(n38559) );
  NAND U39543 ( .A(n38557), .B(n38556), .Z(n38558) );
  NAND U39544 ( .A(n38559), .B(n38558), .Z(n38598) );
  NAND U39545 ( .A(b[0]), .B(a[939]), .Z(n38560) );
  XNOR U39546 ( .A(b[1]), .B(n38560), .Z(n38562) );
  NAND U39547 ( .A(n149), .B(a[938]), .Z(n38561) );
  AND U39548 ( .A(n38562), .B(n38561), .Z(n38615) );
  XOR U39549 ( .A(a[935]), .B(n42197), .Z(n38604) );
  NANDN U39550 ( .A(n38604), .B(n42173), .Z(n38565) );
  NANDN U39551 ( .A(n38563), .B(n42172), .Z(n38564) );
  NAND U39552 ( .A(n38565), .B(n38564), .Z(n38613) );
  NAND U39553 ( .A(b[7]), .B(a[931]), .Z(n38614) );
  XNOR U39554 ( .A(n38613), .B(n38614), .Z(n38616) );
  XOR U39555 ( .A(n38615), .B(n38616), .Z(n38622) );
  NANDN U39556 ( .A(n38566), .B(n42093), .Z(n38568) );
  XOR U39557 ( .A(n42134), .B(a[937]), .Z(n38607) );
  NANDN U39558 ( .A(n38607), .B(n42095), .Z(n38567) );
  NAND U39559 ( .A(n38568), .B(n38567), .Z(n38620) );
  NANDN U39560 ( .A(n38569), .B(n42231), .Z(n38571) );
  XOR U39561 ( .A(n239), .B(a[933]), .Z(n38610) );
  NANDN U39562 ( .A(n38610), .B(n42234), .Z(n38570) );
  AND U39563 ( .A(n38571), .B(n38570), .Z(n38619) );
  XNOR U39564 ( .A(n38620), .B(n38619), .Z(n38621) );
  XNOR U39565 ( .A(n38622), .B(n38621), .Z(n38626) );
  NANDN U39566 ( .A(n38573), .B(n38572), .Z(n38577) );
  NAND U39567 ( .A(n38575), .B(n38574), .Z(n38576) );
  AND U39568 ( .A(n38577), .B(n38576), .Z(n38625) );
  XOR U39569 ( .A(n38626), .B(n38625), .Z(n38627) );
  NANDN U39570 ( .A(n38579), .B(n38578), .Z(n38583) );
  NANDN U39571 ( .A(n38581), .B(n38580), .Z(n38582) );
  NAND U39572 ( .A(n38583), .B(n38582), .Z(n38628) );
  XOR U39573 ( .A(n38627), .B(n38628), .Z(n38595) );
  OR U39574 ( .A(n38585), .B(n38584), .Z(n38589) );
  NANDN U39575 ( .A(n38587), .B(n38586), .Z(n38588) );
  NAND U39576 ( .A(n38589), .B(n38588), .Z(n38596) );
  XNOR U39577 ( .A(n38595), .B(n38596), .Z(n38597) );
  XNOR U39578 ( .A(n38598), .B(n38597), .Z(n38631) );
  XNOR U39579 ( .A(n38631), .B(sreg[1955]), .Z(n38633) );
  NAND U39580 ( .A(n38590), .B(sreg[1954]), .Z(n38594) );
  OR U39581 ( .A(n38592), .B(n38591), .Z(n38593) );
  AND U39582 ( .A(n38594), .B(n38593), .Z(n38632) );
  XOR U39583 ( .A(n38633), .B(n38632), .Z(c[1955]) );
  NANDN U39584 ( .A(n38596), .B(n38595), .Z(n38600) );
  NAND U39585 ( .A(n38598), .B(n38597), .Z(n38599) );
  NAND U39586 ( .A(n38600), .B(n38599), .Z(n38639) );
  NAND U39587 ( .A(b[0]), .B(a[940]), .Z(n38601) );
  XNOR U39588 ( .A(b[1]), .B(n38601), .Z(n38603) );
  NAND U39589 ( .A(n149), .B(a[939]), .Z(n38602) );
  AND U39590 ( .A(n38603), .B(n38602), .Z(n38656) );
  XOR U39591 ( .A(a[936]), .B(n42197), .Z(n38645) );
  NANDN U39592 ( .A(n38645), .B(n42173), .Z(n38606) );
  NANDN U39593 ( .A(n38604), .B(n42172), .Z(n38605) );
  NAND U39594 ( .A(n38606), .B(n38605), .Z(n38654) );
  NAND U39595 ( .A(b[7]), .B(a[932]), .Z(n38655) );
  XNOR U39596 ( .A(n38654), .B(n38655), .Z(n38657) );
  XOR U39597 ( .A(n38656), .B(n38657), .Z(n38663) );
  NANDN U39598 ( .A(n38607), .B(n42093), .Z(n38609) );
  XOR U39599 ( .A(n42134), .B(a[938]), .Z(n38648) );
  NANDN U39600 ( .A(n38648), .B(n42095), .Z(n38608) );
  NAND U39601 ( .A(n38609), .B(n38608), .Z(n38661) );
  NANDN U39602 ( .A(n38610), .B(n42231), .Z(n38612) );
  XOR U39603 ( .A(n239), .B(a[934]), .Z(n38651) );
  NANDN U39604 ( .A(n38651), .B(n42234), .Z(n38611) );
  AND U39605 ( .A(n38612), .B(n38611), .Z(n38660) );
  XNOR U39606 ( .A(n38661), .B(n38660), .Z(n38662) );
  XNOR U39607 ( .A(n38663), .B(n38662), .Z(n38667) );
  NANDN U39608 ( .A(n38614), .B(n38613), .Z(n38618) );
  NAND U39609 ( .A(n38616), .B(n38615), .Z(n38617) );
  AND U39610 ( .A(n38618), .B(n38617), .Z(n38666) );
  XOR U39611 ( .A(n38667), .B(n38666), .Z(n38668) );
  NANDN U39612 ( .A(n38620), .B(n38619), .Z(n38624) );
  NANDN U39613 ( .A(n38622), .B(n38621), .Z(n38623) );
  NAND U39614 ( .A(n38624), .B(n38623), .Z(n38669) );
  XOR U39615 ( .A(n38668), .B(n38669), .Z(n38636) );
  OR U39616 ( .A(n38626), .B(n38625), .Z(n38630) );
  NANDN U39617 ( .A(n38628), .B(n38627), .Z(n38629) );
  NAND U39618 ( .A(n38630), .B(n38629), .Z(n38637) );
  XNOR U39619 ( .A(n38636), .B(n38637), .Z(n38638) );
  XNOR U39620 ( .A(n38639), .B(n38638), .Z(n38672) );
  XNOR U39621 ( .A(n38672), .B(sreg[1956]), .Z(n38674) );
  NAND U39622 ( .A(n38631), .B(sreg[1955]), .Z(n38635) );
  OR U39623 ( .A(n38633), .B(n38632), .Z(n38634) );
  AND U39624 ( .A(n38635), .B(n38634), .Z(n38673) );
  XOR U39625 ( .A(n38674), .B(n38673), .Z(c[1956]) );
  NANDN U39626 ( .A(n38637), .B(n38636), .Z(n38641) );
  NAND U39627 ( .A(n38639), .B(n38638), .Z(n38640) );
  NAND U39628 ( .A(n38641), .B(n38640), .Z(n38680) );
  NAND U39629 ( .A(b[0]), .B(a[941]), .Z(n38642) );
  XNOR U39630 ( .A(b[1]), .B(n38642), .Z(n38644) );
  NAND U39631 ( .A(n149), .B(a[940]), .Z(n38643) );
  AND U39632 ( .A(n38644), .B(n38643), .Z(n38697) );
  XOR U39633 ( .A(a[937]), .B(n42197), .Z(n38686) );
  NANDN U39634 ( .A(n38686), .B(n42173), .Z(n38647) );
  NANDN U39635 ( .A(n38645), .B(n42172), .Z(n38646) );
  NAND U39636 ( .A(n38647), .B(n38646), .Z(n38695) );
  NAND U39637 ( .A(b[7]), .B(a[933]), .Z(n38696) );
  XNOR U39638 ( .A(n38695), .B(n38696), .Z(n38698) );
  XOR U39639 ( .A(n38697), .B(n38698), .Z(n38704) );
  NANDN U39640 ( .A(n38648), .B(n42093), .Z(n38650) );
  XOR U39641 ( .A(n42134), .B(a[939]), .Z(n38689) );
  NANDN U39642 ( .A(n38689), .B(n42095), .Z(n38649) );
  NAND U39643 ( .A(n38650), .B(n38649), .Z(n38702) );
  NANDN U39644 ( .A(n38651), .B(n42231), .Z(n38653) );
  XOR U39645 ( .A(n240), .B(a[935]), .Z(n38692) );
  NANDN U39646 ( .A(n38692), .B(n42234), .Z(n38652) );
  AND U39647 ( .A(n38653), .B(n38652), .Z(n38701) );
  XNOR U39648 ( .A(n38702), .B(n38701), .Z(n38703) );
  XNOR U39649 ( .A(n38704), .B(n38703), .Z(n38708) );
  NANDN U39650 ( .A(n38655), .B(n38654), .Z(n38659) );
  NAND U39651 ( .A(n38657), .B(n38656), .Z(n38658) );
  AND U39652 ( .A(n38659), .B(n38658), .Z(n38707) );
  XOR U39653 ( .A(n38708), .B(n38707), .Z(n38709) );
  NANDN U39654 ( .A(n38661), .B(n38660), .Z(n38665) );
  NANDN U39655 ( .A(n38663), .B(n38662), .Z(n38664) );
  NAND U39656 ( .A(n38665), .B(n38664), .Z(n38710) );
  XOR U39657 ( .A(n38709), .B(n38710), .Z(n38677) );
  OR U39658 ( .A(n38667), .B(n38666), .Z(n38671) );
  NANDN U39659 ( .A(n38669), .B(n38668), .Z(n38670) );
  NAND U39660 ( .A(n38671), .B(n38670), .Z(n38678) );
  XNOR U39661 ( .A(n38677), .B(n38678), .Z(n38679) );
  XNOR U39662 ( .A(n38680), .B(n38679), .Z(n38713) );
  XNOR U39663 ( .A(n38713), .B(sreg[1957]), .Z(n38715) );
  NAND U39664 ( .A(n38672), .B(sreg[1956]), .Z(n38676) );
  OR U39665 ( .A(n38674), .B(n38673), .Z(n38675) );
  AND U39666 ( .A(n38676), .B(n38675), .Z(n38714) );
  XOR U39667 ( .A(n38715), .B(n38714), .Z(c[1957]) );
  NANDN U39668 ( .A(n38678), .B(n38677), .Z(n38682) );
  NAND U39669 ( .A(n38680), .B(n38679), .Z(n38681) );
  NAND U39670 ( .A(n38682), .B(n38681), .Z(n38721) );
  NAND U39671 ( .A(b[0]), .B(a[942]), .Z(n38683) );
  XNOR U39672 ( .A(b[1]), .B(n38683), .Z(n38685) );
  NAND U39673 ( .A(n149), .B(a[941]), .Z(n38684) );
  AND U39674 ( .A(n38685), .B(n38684), .Z(n38738) );
  XOR U39675 ( .A(a[938]), .B(n42197), .Z(n38727) );
  NANDN U39676 ( .A(n38727), .B(n42173), .Z(n38688) );
  NANDN U39677 ( .A(n38686), .B(n42172), .Z(n38687) );
  NAND U39678 ( .A(n38688), .B(n38687), .Z(n38736) );
  NAND U39679 ( .A(b[7]), .B(a[934]), .Z(n38737) );
  XNOR U39680 ( .A(n38736), .B(n38737), .Z(n38739) );
  XOR U39681 ( .A(n38738), .B(n38739), .Z(n38745) );
  NANDN U39682 ( .A(n38689), .B(n42093), .Z(n38691) );
  XOR U39683 ( .A(n42134), .B(a[940]), .Z(n38730) );
  NANDN U39684 ( .A(n38730), .B(n42095), .Z(n38690) );
  NAND U39685 ( .A(n38691), .B(n38690), .Z(n38743) );
  NANDN U39686 ( .A(n38692), .B(n42231), .Z(n38694) );
  XOR U39687 ( .A(n240), .B(a[936]), .Z(n38733) );
  NANDN U39688 ( .A(n38733), .B(n42234), .Z(n38693) );
  AND U39689 ( .A(n38694), .B(n38693), .Z(n38742) );
  XNOR U39690 ( .A(n38743), .B(n38742), .Z(n38744) );
  XNOR U39691 ( .A(n38745), .B(n38744), .Z(n38749) );
  NANDN U39692 ( .A(n38696), .B(n38695), .Z(n38700) );
  NAND U39693 ( .A(n38698), .B(n38697), .Z(n38699) );
  AND U39694 ( .A(n38700), .B(n38699), .Z(n38748) );
  XOR U39695 ( .A(n38749), .B(n38748), .Z(n38750) );
  NANDN U39696 ( .A(n38702), .B(n38701), .Z(n38706) );
  NANDN U39697 ( .A(n38704), .B(n38703), .Z(n38705) );
  NAND U39698 ( .A(n38706), .B(n38705), .Z(n38751) );
  XOR U39699 ( .A(n38750), .B(n38751), .Z(n38718) );
  OR U39700 ( .A(n38708), .B(n38707), .Z(n38712) );
  NANDN U39701 ( .A(n38710), .B(n38709), .Z(n38711) );
  NAND U39702 ( .A(n38712), .B(n38711), .Z(n38719) );
  XNOR U39703 ( .A(n38718), .B(n38719), .Z(n38720) );
  XNOR U39704 ( .A(n38721), .B(n38720), .Z(n38754) );
  XNOR U39705 ( .A(n38754), .B(sreg[1958]), .Z(n38756) );
  NAND U39706 ( .A(n38713), .B(sreg[1957]), .Z(n38717) );
  OR U39707 ( .A(n38715), .B(n38714), .Z(n38716) );
  AND U39708 ( .A(n38717), .B(n38716), .Z(n38755) );
  XOR U39709 ( .A(n38756), .B(n38755), .Z(c[1958]) );
  NANDN U39710 ( .A(n38719), .B(n38718), .Z(n38723) );
  NAND U39711 ( .A(n38721), .B(n38720), .Z(n38722) );
  NAND U39712 ( .A(n38723), .B(n38722), .Z(n38762) );
  NAND U39713 ( .A(b[0]), .B(a[943]), .Z(n38724) );
  XNOR U39714 ( .A(b[1]), .B(n38724), .Z(n38726) );
  NAND U39715 ( .A(n149), .B(a[942]), .Z(n38725) );
  AND U39716 ( .A(n38726), .B(n38725), .Z(n38779) );
  XOR U39717 ( .A(a[939]), .B(n42197), .Z(n38768) );
  NANDN U39718 ( .A(n38768), .B(n42173), .Z(n38729) );
  NANDN U39719 ( .A(n38727), .B(n42172), .Z(n38728) );
  NAND U39720 ( .A(n38729), .B(n38728), .Z(n38777) );
  NAND U39721 ( .A(b[7]), .B(a[935]), .Z(n38778) );
  XNOR U39722 ( .A(n38777), .B(n38778), .Z(n38780) );
  XOR U39723 ( .A(n38779), .B(n38780), .Z(n38786) );
  NANDN U39724 ( .A(n38730), .B(n42093), .Z(n38732) );
  XOR U39725 ( .A(n42134), .B(a[941]), .Z(n38771) );
  NANDN U39726 ( .A(n38771), .B(n42095), .Z(n38731) );
  NAND U39727 ( .A(n38732), .B(n38731), .Z(n38784) );
  NANDN U39728 ( .A(n38733), .B(n42231), .Z(n38735) );
  XOR U39729 ( .A(n240), .B(a[937]), .Z(n38774) );
  NANDN U39730 ( .A(n38774), .B(n42234), .Z(n38734) );
  AND U39731 ( .A(n38735), .B(n38734), .Z(n38783) );
  XNOR U39732 ( .A(n38784), .B(n38783), .Z(n38785) );
  XNOR U39733 ( .A(n38786), .B(n38785), .Z(n38790) );
  NANDN U39734 ( .A(n38737), .B(n38736), .Z(n38741) );
  NAND U39735 ( .A(n38739), .B(n38738), .Z(n38740) );
  AND U39736 ( .A(n38741), .B(n38740), .Z(n38789) );
  XOR U39737 ( .A(n38790), .B(n38789), .Z(n38791) );
  NANDN U39738 ( .A(n38743), .B(n38742), .Z(n38747) );
  NANDN U39739 ( .A(n38745), .B(n38744), .Z(n38746) );
  NAND U39740 ( .A(n38747), .B(n38746), .Z(n38792) );
  XOR U39741 ( .A(n38791), .B(n38792), .Z(n38759) );
  OR U39742 ( .A(n38749), .B(n38748), .Z(n38753) );
  NANDN U39743 ( .A(n38751), .B(n38750), .Z(n38752) );
  NAND U39744 ( .A(n38753), .B(n38752), .Z(n38760) );
  XNOR U39745 ( .A(n38759), .B(n38760), .Z(n38761) );
  XNOR U39746 ( .A(n38762), .B(n38761), .Z(n38795) );
  XNOR U39747 ( .A(n38795), .B(sreg[1959]), .Z(n38797) );
  NAND U39748 ( .A(n38754), .B(sreg[1958]), .Z(n38758) );
  OR U39749 ( .A(n38756), .B(n38755), .Z(n38757) );
  AND U39750 ( .A(n38758), .B(n38757), .Z(n38796) );
  XOR U39751 ( .A(n38797), .B(n38796), .Z(c[1959]) );
  NANDN U39752 ( .A(n38760), .B(n38759), .Z(n38764) );
  NAND U39753 ( .A(n38762), .B(n38761), .Z(n38763) );
  NAND U39754 ( .A(n38764), .B(n38763), .Z(n38803) );
  NAND U39755 ( .A(b[0]), .B(a[944]), .Z(n38765) );
  XNOR U39756 ( .A(b[1]), .B(n38765), .Z(n38767) );
  NAND U39757 ( .A(n149), .B(a[943]), .Z(n38766) );
  AND U39758 ( .A(n38767), .B(n38766), .Z(n38820) );
  XOR U39759 ( .A(a[940]), .B(n42197), .Z(n38809) );
  NANDN U39760 ( .A(n38809), .B(n42173), .Z(n38770) );
  NANDN U39761 ( .A(n38768), .B(n42172), .Z(n38769) );
  NAND U39762 ( .A(n38770), .B(n38769), .Z(n38818) );
  NAND U39763 ( .A(b[7]), .B(a[936]), .Z(n38819) );
  XNOR U39764 ( .A(n38818), .B(n38819), .Z(n38821) );
  XOR U39765 ( .A(n38820), .B(n38821), .Z(n38827) );
  NANDN U39766 ( .A(n38771), .B(n42093), .Z(n38773) );
  XOR U39767 ( .A(n42134), .B(a[942]), .Z(n38812) );
  NANDN U39768 ( .A(n38812), .B(n42095), .Z(n38772) );
  NAND U39769 ( .A(n38773), .B(n38772), .Z(n38825) );
  NANDN U39770 ( .A(n38774), .B(n42231), .Z(n38776) );
  XOR U39771 ( .A(n240), .B(a[938]), .Z(n38815) );
  NANDN U39772 ( .A(n38815), .B(n42234), .Z(n38775) );
  AND U39773 ( .A(n38776), .B(n38775), .Z(n38824) );
  XNOR U39774 ( .A(n38825), .B(n38824), .Z(n38826) );
  XNOR U39775 ( .A(n38827), .B(n38826), .Z(n38831) );
  NANDN U39776 ( .A(n38778), .B(n38777), .Z(n38782) );
  NAND U39777 ( .A(n38780), .B(n38779), .Z(n38781) );
  AND U39778 ( .A(n38782), .B(n38781), .Z(n38830) );
  XOR U39779 ( .A(n38831), .B(n38830), .Z(n38832) );
  NANDN U39780 ( .A(n38784), .B(n38783), .Z(n38788) );
  NANDN U39781 ( .A(n38786), .B(n38785), .Z(n38787) );
  NAND U39782 ( .A(n38788), .B(n38787), .Z(n38833) );
  XOR U39783 ( .A(n38832), .B(n38833), .Z(n38800) );
  OR U39784 ( .A(n38790), .B(n38789), .Z(n38794) );
  NANDN U39785 ( .A(n38792), .B(n38791), .Z(n38793) );
  NAND U39786 ( .A(n38794), .B(n38793), .Z(n38801) );
  XNOR U39787 ( .A(n38800), .B(n38801), .Z(n38802) );
  XNOR U39788 ( .A(n38803), .B(n38802), .Z(n38836) );
  XNOR U39789 ( .A(n38836), .B(sreg[1960]), .Z(n38838) );
  NAND U39790 ( .A(n38795), .B(sreg[1959]), .Z(n38799) );
  OR U39791 ( .A(n38797), .B(n38796), .Z(n38798) );
  AND U39792 ( .A(n38799), .B(n38798), .Z(n38837) );
  XOR U39793 ( .A(n38838), .B(n38837), .Z(c[1960]) );
  NANDN U39794 ( .A(n38801), .B(n38800), .Z(n38805) );
  NAND U39795 ( .A(n38803), .B(n38802), .Z(n38804) );
  NAND U39796 ( .A(n38805), .B(n38804), .Z(n38844) );
  NAND U39797 ( .A(b[0]), .B(a[945]), .Z(n38806) );
  XNOR U39798 ( .A(b[1]), .B(n38806), .Z(n38808) );
  NAND U39799 ( .A(n150), .B(a[944]), .Z(n38807) );
  AND U39800 ( .A(n38808), .B(n38807), .Z(n38861) );
  XOR U39801 ( .A(a[941]), .B(n42197), .Z(n38850) );
  NANDN U39802 ( .A(n38850), .B(n42173), .Z(n38811) );
  NANDN U39803 ( .A(n38809), .B(n42172), .Z(n38810) );
  NAND U39804 ( .A(n38811), .B(n38810), .Z(n38859) );
  NAND U39805 ( .A(b[7]), .B(a[937]), .Z(n38860) );
  XNOR U39806 ( .A(n38859), .B(n38860), .Z(n38862) );
  XOR U39807 ( .A(n38861), .B(n38862), .Z(n38868) );
  NANDN U39808 ( .A(n38812), .B(n42093), .Z(n38814) );
  XOR U39809 ( .A(n42134), .B(a[943]), .Z(n38853) );
  NANDN U39810 ( .A(n38853), .B(n42095), .Z(n38813) );
  NAND U39811 ( .A(n38814), .B(n38813), .Z(n38866) );
  NANDN U39812 ( .A(n38815), .B(n42231), .Z(n38817) );
  XOR U39813 ( .A(n240), .B(a[939]), .Z(n38856) );
  NANDN U39814 ( .A(n38856), .B(n42234), .Z(n38816) );
  AND U39815 ( .A(n38817), .B(n38816), .Z(n38865) );
  XNOR U39816 ( .A(n38866), .B(n38865), .Z(n38867) );
  XNOR U39817 ( .A(n38868), .B(n38867), .Z(n38872) );
  NANDN U39818 ( .A(n38819), .B(n38818), .Z(n38823) );
  NAND U39819 ( .A(n38821), .B(n38820), .Z(n38822) );
  AND U39820 ( .A(n38823), .B(n38822), .Z(n38871) );
  XOR U39821 ( .A(n38872), .B(n38871), .Z(n38873) );
  NANDN U39822 ( .A(n38825), .B(n38824), .Z(n38829) );
  NANDN U39823 ( .A(n38827), .B(n38826), .Z(n38828) );
  NAND U39824 ( .A(n38829), .B(n38828), .Z(n38874) );
  XOR U39825 ( .A(n38873), .B(n38874), .Z(n38841) );
  OR U39826 ( .A(n38831), .B(n38830), .Z(n38835) );
  NANDN U39827 ( .A(n38833), .B(n38832), .Z(n38834) );
  NAND U39828 ( .A(n38835), .B(n38834), .Z(n38842) );
  XNOR U39829 ( .A(n38841), .B(n38842), .Z(n38843) );
  XNOR U39830 ( .A(n38844), .B(n38843), .Z(n38877) );
  XNOR U39831 ( .A(n38877), .B(sreg[1961]), .Z(n38879) );
  NAND U39832 ( .A(n38836), .B(sreg[1960]), .Z(n38840) );
  OR U39833 ( .A(n38838), .B(n38837), .Z(n38839) );
  AND U39834 ( .A(n38840), .B(n38839), .Z(n38878) );
  XOR U39835 ( .A(n38879), .B(n38878), .Z(c[1961]) );
  NANDN U39836 ( .A(n38842), .B(n38841), .Z(n38846) );
  NAND U39837 ( .A(n38844), .B(n38843), .Z(n38845) );
  NAND U39838 ( .A(n38846), .B(n38845), .Z(n38885) );
  NAND U39839 ( .A(b[0]), .B(a[946]), .Z(n38847) );
  XNOR U39840 ( .A(b[1]), .B(n38847), .Z(n38849) );
  NAND U39841 ( .A(n150), .B(a[945]), .Z(n38848) );
  AND U39842 ( .A(n38849), .B(n38848), .Z(n38902) );
  XOR U39843 ( .A(a[942]), .B(n42197), .Z(n38891) );
  NANDN U39844 ( .A(n38891), .B(n42173), .Z(n38852) );
  NANDN U39845 ( .A(n38850), .B(n42172), .Z(n38851) );
  NAND U39846 ( .A(n38852), .B(n38851), .Z(n38900) );
  NAND U39847 ( .A(b[7]), .B(a[938]), .Z(n38901) );
  XNOR U39848 ( .A(n38900), .B(n38901), .Z(n38903) );
  XOR U39849 ( .A(n38902), .B(n38903), .Z(n38909) );
  NANDN U39850 ( .A(n38853), .B(n42093), .Z(n38855) );
  XOR U39851 ( .A(n42134), .B(a[944]), .Z(n38894) );
  NANDN U39852 ( .A(n38894), .B(n42095), .Z(n38854) );
  NAND U39853 ( .A(n38855), .B(n38854), .Z(n38907) );
  NANDN U39854 ( .A(n38856), .B(n42231), .Z(n38858) );
  XOR U39855 ( .A(n240), .B(a[940]), .Z(n38897) );
  NANDN U39856 ( .A(n38897), .B(n42234), .Z(n38857) );
  AND U39857 ( .A(n38858), .B(n38857), .Z(n38906) );
  XNOR U39858 ( .A(n38907), .B(n38906), .Z(n38908) );
  XNOR U39859 ( .A(n38909), .B(n38908), .Z(n38913) );
  NANDN U39860 ( .A(n38860), .B(n38859), .Z(n38864) );
  NAND U39861 ( .A(n38862), .B(n38861), .Z(n38863) );
  AND U39862 ( .A(n38864), .B(n38863), .Z(n38912) );
  XOR U39863 ( .A(n38913), .B(n38912), .Z(n38914) );
  NANDN U39864 ( .A(n38866), .B(n38865), .Z(n38870) );
  NANDN U39865 ( .A(n38868), .B(n38867), .Z(n38869) );
  NAND U39866 ( .A(n38870), .B(n38869), .Z(n38915) );
  XOR U39867 ( .A(n38914), .B(n38915), .Z(n38882) );
  OR U39868 ( .A(n38872), .B(n38871), .Z(n38876) );
  NANDN U39869 ( .A(n38874), .B(n38873), .Z(n38875) );
  NAND U39870 ( .A(n38876), .B(n38875), .Z(n38883) );
  XNOR U39871 ( .A(n38882), .B(n38883), .Z(n38884) );
  XNOR U39872 ( .A(n38885), .B(n38884), .Z(n38918) );
  XNOR U39873 ( .A(n38918), .B(sreg[1962]), .Z(n38920) );
  NAND U39874 ( .A(n38877), .B(sreg[1961]), .Z(n38881) );
  OR U39875 ( .A(n38879), .B(n38878), .Z(n38880) );
  AND U39876 ( .A(n38881), .B(n38880), .Z(n38919) );
  XOR U39877 ( .A(n38920), .B(n38919), .Z(c[1962]) );
  NANDN U39878 ( .A(n38883), .B(n38882), .Z(n38887) );
  NAND U39879 ( .A(n38885), .B(n38884), .Z(n38886) );
  NAND U39880 ( .A(n38887), .B(n38886), .Z(n38926) );
  NAND U39881 ( .A(b[0]), .B(a[947]), .Z(n38888) );
  XNOR U39882 ( .A(b[1]), .B(n38888), .Z(n38890) );
  NAND U39883 ( .A(n150), .B(a[946]), .Z(n38889) );
  AND U39884 ( .A(n38890), .B(n38889), .Z(n38943) );
  XOR U39885 ( .A(a[943]), .B(n42197), .Z(n38932) );
  NANDN U39886 ( .A(n38932), .B(n42173), .Z(n38893) );
  NANDN U39887 ( .A(n38891), .B(n42172), .Z(n38892) );
  NAND U39888 ( .A(n38893), .B(n38892), .Z(n38941) );
  NAND U39889 ( .A(b[7]), .B(a[939]), .Z(n38942) );
  XNOR U39890 ( .A(n38941), .B(n38942), .Z(n38944) );
  XOR U39891 ( .A(n38943), .B(n38944), .Z(n38950) );
  NANDN U39892 ( .A(n38894), .B(n42093), .Z(n38896) );
  XOR U39893 ( .A(n42134), .B(a[945]), .Z(n38935) );
  NANDN U39894 ( .A(n38935), .B(n42095), .Z(n38895) );
  NAND U39895 ( .A(n38896), .B(n38895), .Z(n38948) );
  NANDN U39896 ( .A(n38897), .B(n42231), .Z(n38899) );
  XOR U39897 ( .A(n240), .B(a[941]), .Z(n38938) );
  NANDN U39898 ( .A(n38938), .B(n42234), .Z(n38898) );
  AND U39899 ( .A(n38899), .B(n38898), .Z(n38947) );
  XNOR U39900 ( .A(n38948), .B(n38947), .Z(n38949) );
  XNOR U39901 ( .A(n38950), .B(n38949), .Z(n38954) );
  NANDN U39902 ( .A(n38901), .B(n38900), .Z(n38905) );
  NAND U39903 ( .A(n38903), .B(n38902), .Z(n38904) );
  AND U39904 ( .A(n38905), .B(n38904), .Z(n38953) );
  XOR U39905 ( .A(n38954), .B(n38953), .Z(n38955) );
  NANDN U39906 ( .A(n38907), .B(n38906), .Z(n38911) );
  NANDN U39907 ( .A(n38909), .B(n38908), .Z(n38910) );
  NAND U39908 ( .A(n38911), .B(n38910), .Z(n38956) );
  XOR U39909 ( .A(n38955), .B(n38956), .Z(n38923) );
  OR U39910 ( .A(n38913), .B(n38912), .Z(n38917) );
  NANDN U39911 ( .A(n38915), .B(n38914), .Z(n38916) );
  NAND U39912 ( .A(n38917), .B(n38916), .Z(n38924) );
  XNOR U39913 ( .A(n38923), .B(n38924), .Z(n38925) );
  XNOR U39914 ( .A(n38926), .B(n38925), .Z(n38959) );
  XNOR U39915 ( .A(n38959), .B(sreg[1963]), .Z(n38961) );
  NAND U39916 ( .A(n38918), .B(sreg[1962]), .Z(n38922) );
  OR U39917 ( .A(n38920), .B(n38919), .Z(n38921) );
  AND U39918 ( .A(n38922), .B(n38921), .Z(n38960) );
  XOR U39919 ( .A(n38961), .B(n38960), .Z(c[1963]) );
  NANDN U39920 ( .A(n38924), .B(n38923), .Z(n38928) );
  NAND U39921 ( .A(n38926), .B(n38925), .Z(n38927) );
  NAND U39922 ( .A(n38928), .B(n38927), .Z(n38967) );
  NAND U39923 ( .A(b[0]), .B(a[948]), .Z(n38929) );
  XNOR U39924 ( .A(b[1]), .B(n38929), .Z(n38931) );
  NAND U39925 ( .A(n150), .B(a[947]), .Z(n38930) );
  AND U39926 ( .A(n38931), .B(n38930), .Z(n38984) );
  XOR U39927 ( .A(a[944]), .B(n42197), .Z(n38973) );
  NANDN U39928 ( .A(n38973), .B(n42173), .Z(n38934) );
  NANDN U39929 ( .A(n38932), .B(n42172), .Z(n38933) );
  NAND U39930 ( .A(n38934), .B(n38933), .Z(n38982) );
  NAND U39931 ( .A(b[7]), .B(a[940]), .Z(n38983) );
  XNOR U39932 ( .A(n38982), .B(n38983), .Z(n38985) );
  XOR U39933 ( .A(n38984), .B(n38985), .Z(n38991) );
  NANDN U39934 ( .A(n38935), .B(n42093), .Z(n38937) );
  XOR U39935 ( .A(n42134), .B(a[946]), .Z(n38976) );
  NANDN U39936 ( .A(n38976), .B(n42095), .Z(n38936) );
  NAND U39937 ( .A(n38937), .B(n38936), .Z(n38989) );
  NANDN U39938 ( .A(n38938), .B(n42231), .Z(n38940) );
  XOR U39939 ( .A(n240), .B(a[942]), .Z(n38979) );
  NANDN U39940 ( .A(n38979), .B(n42234), .Z(n38939) );
  AND U39941 ( .A(n38940), .B(n38939), .Z(n38988) );
  XNOR U39942 ( .A(n38989), .B(n38988), .Z(n38990) );
  XNOR U39943 ( .A(n38991), .B(n38990), .Z(n38995) );
  NANDN U39944 ( .A(n38942), .B(n38941), .Z(n38946) );
  NAND U39945 ( .A(n38944), .B(n38943), .Z(n38945) );
  AND U39946 ( .A(n38946), .B(n38945), .Z(n38994) );
  XOR U39947 ( .A(n38995), .B(n38994), .Z(n38996) );
  NANDN U39948 ( .A(n38948), .B(n38947), .Z(n38952) );
  NANDN U39949 ( .A(n38950), .B(n38949), .Z(n38951) );
  NAND U39950 ( .A(n38952), .B(n38951), .Z(n38997) );
  XOR U39951 ( .A(n38996), .B(n38997), .Z(n38964) );
  OR U39952 ( .A(n38954), .B(n38953), .Z(n38958) );
  NANDN U39953 ( .A(n38956), .B(n38955), .Z(n38957) );
  NAND U39954 ( .A(n38958), .B(n38957), .Z(n38965) );
  XNOR U39955 ( .A(n38964), .B(n38965), .Z(n38966) );
  XNOR U39956 ( .A(n38967), .B(n38966), .Z(n39000) );
  XNOR U39957 ( .A(n39000), .B(sreg[1964]), .Z(n39002) );
  NAND U39958 ( .A(n38959), .B(sreg[1963]), .Z(n38963) );
  OR U39959 ( .A(n38961), .B(n38960), .Z(n38962) );
  AND U39960 ( .A(n38963), .B(n38962), .Z(n39001) );
  XOR U39961 ( .A(n39002), .B(n39001), .Z(c[1964]) );
  NANDN U39962 ( .A(n38965), .B(n38964), .Z(n38969) );
  NAND U39963 ( .A(n38967), .B(n38966), .Z(n38968) );
  NAND U39964 ( .A(n38969), .B(n38968), .Z(n39008) );
  NAND U39965 ( .A(b[0]), .B(a[949]), .Z(n38970) );
  XNOR U39966 ( .A(b[1]), .B(n38970), .Z(n38972) );
  NAND U39967 ( .A(n150), .B(a[948]), .Z(n38971) );
  AND U39968 ( .A(n38972), .B(n38971), .Z(n39025) );
  XOR U39969 ( .A(a[945]), .B(n42197), .Z(n39014) );
  NANDN U39970 ( .A(n39014), .B(n42173), .Z(n38975) );
  NANDN U39971 ( .A(n38973), .B(n42172), .Z(n38974) );
  NAND U39972 ( .A(n38975), .B(n38974), .Z(n39023) );
  NAND U39973 ( .A(b[7]), .B(a[941]), .Z(n39024) );
  XNOR U39974 ( .A(n39023), .B(n39024), .Z(n39026) );
  XOR U39975 ( .A(n39025), .B(n39026), .Z(n39032) );
  NANDN U39976 ( .A(n38976), .B(n42093), .Z(n38978) );
  XOR U39977 ( .A(n42134), .B(a[947]), .Z(n39017) );
  NANDN U39978 ( .A(n39017), .B(n42095), .Z(n38977) );
  NAND U39979 ( .A(n38978), .B(n38977), .Z(n39030) );
  NANDN U39980 ( .A(n38979), .B(n42231), .Z(n38981) );
  XOR U39981 ( .A(n240), .B(a[943]), .Z(n39020) );
  NANDN U39982 ( .A(n39020), .B(n42234), .Z(n38980) );
  AND U39983 ( .A(n38981), .B(n38980), .Z(n39029) );
  XNOR U39984 ( .A(n39030), .B(n39029), .Z(n39031) );
  XNOR U39985 ( .A(n39032), .B(n39031), .Z(n39036) );
  NANDN U39986 ( .A(n38983), .B(n38982), .Z(n38987) );
  NAND U39987 ( .A(n38985), .B(n38984), .Z(n38986) );
  AND U39988 ( .A(n38987), .B(n38986), .Z(n39035) );
  XOR U39989 ( .A(n39036), .B(n39035), .Z(n39037) );
  NANDN U39990 ( .A(n38989), .B(n38988), .Z(n38993) );
  NANDN U39991 ( .A(n38991), .B(n38990), .Z(n38992) );
  NAND U39992 ( .A(n38993), .B(n38992), .Z(n39038) );
  XOR U39993 ( .A(n39037), .B(n39038), .Z(n39005) );
  OR U39994 ( .A(n38995), .B(n38994), .Z(n38999) );
  NANDN U39995 ( .A(n38997), .B(n38996), .Z(n38998) );
  NAND U39996 ( .A(n38999), .B(n38998), .Z(n39006) );
  XNOR U39997 ( .A(n39005), .B(n39006), .Z(n39007) );
  XNOR U39998 ( .A(n39008), .B(n39007), .Z(n39041) );
  XNOR U39999 ( .A(n39041), .B(sreg[1965]), .Z(n39043) );
  NAND U40000 ( .A(n39000), .B(sreg[1964]), .Z(n39004) );
  OR U40001 ( .A(n39002), .B(n39001), .Z(n39003) );
  AND U40002 ( .A(n39004), .B(n39003), .Z(n39042) );
  XOR U40003 ( .A(n39043), .B(n39042), .Z(c[1965]) );
  NANDN U40004 ( .A(n39006), .B(n39005), .Z(n39010) );
  NAND U40005 ( .A(n39008), .B(n39007), .Z(n39009) );
  NAND U40006 ( .A(n39010), .B(n39009), .Z(n39049) );
  NAND U40007 ( .A(b[0]), .B(a[950]), .Z(n39011) );
  XNOR U40008 ( .A(b[1]), .B(n39011), .Z(n39013) );
  NAND U40009 ( .A(n150), .B(a[949]), .Z(n39012) );
  AND U40010 ( .A(n39013), .B(n39012), .Z(n39066) );
  XOR U40011 ( .A(a[946]), .B(n42197), .Z(n39055) );
  NANDN U40012 ( .A(n39055), .B(n42173), .Z(n39016) );
  NANDN U40013 ( .A(n39014), .B(n42172), .Z(n39015) );
  NAND U40014 ( .A(n39016), .B(n39015), .Z(n39064) );
  NAND U40015 ( .A(b[7]), .B(a[942]), .Z(n39065) );
  XNOR U40016 ( .A(n39064), .B(n39065), .Z(n39067) );
  XOR U40017 ( .A(n39066), .B(n39067), .Z(n39073) );
  NANDN U40018 ( .A(n39017), .B(n42093), .Z(n39019) );
  XOR U40019 ( .A(n42134), .B(a[948]), .Z(n39058) );
  NANDN U40020 ( .A(n39058), .B(n42095), .Z(n39018) );
  NAND U40021 ( .A(n39019), .B(n39018), .Z(n39071) );
  NANDN U40022 ( .A(n39020), .B(n42231), .Z(n39022) );
  XOR U40023 ( .A(n240), .B(a[944]), .Z(n39061) );
  NANDN U40024 ( .A(n39061), .B(n42234), .Z(n39021) );
  AND U40025 ( .A(n39022), .B(n39021), .Z(n39070) );
  XNOR U40026 ( .A(n39071), .B(n39070), .Z(n39072) );
  XNOR U40027 ( .A(n39073), .B(n39072), .Z(n39077) );
  NANDN U40028 ( .A(n39024), .B(n39023), .Z(n39028) );
  NAND U40029 ( .A(n39026), .B(n39025), .Z(n39027) );
  AND U40030 ( .A(n39028), .B(n39027), .Z(n39076) );
  XOR U40031 ( .A(n39077), .B(n39076), .Z(n39078) );
  NANDN U40032 ( .A(n39030), .B(n39029), .Z(n39034) );
  NANDN U40033 ( .A(n39032), .B(n39031), .Z(n39033) );
  NAND U40034 ( .A(n39034), .B(n39033), .Z(n39079) );
  XOR U40035 ( .A(n39078), .B(n39079), .Z(n39046) );
  OR U40036 ( .A(n39036), .B(n39035), .Z(n39040) );
  NANDN U40037 ( .A(n39038), .B(n39037), .Z(n39039) );
  NAND U40038 ( .A(n39040), .B(n39039), .Z(n39047) );
  XNOR U40039 ( .A(n39046), .B(n39047), .Z(n39048) );
  XNOR U40040 ( .A(n39049), .B(n39048), .Z(n39082) );
  XNOR U40041 ( .A(n39082), .B(sreg[1966]), .Z(n39084) );
  NAND U40042 ( .A(n39041), .B(sreg[1965]), .Z(n39045) );
  OR U40043 ( .A(n39043), .B(n39042), .Z(n39044) );
  AND U40044 ( .A(n39045), .B(n39044), .Z(n39083) );
  XOR U40045 ( .A(n39084), .B(n39083), .Z(c[1966]) );
  NANDN U40046 ( .A(n39047), .B(n39046), .Z(n39051) );
  NAND U40047 ( .A(n39049), .B(n39048), .Z(n39050) );
  NAND U40048 ( .A(n39051), .B(n39050), .Z(n39090) );
  NAND U40049 ( .A(b[0]), .B(a[951]), .Z(n39052) );
  XNOR U40050 ( .A(b[1]), .B(n39052), .Z(n39054) );
  NAND U40051 ( .A(n150), .B(a[950]), .Z(n39053) );
  AND U40052 ( .A(n39054), .B(n39053), .Z(n39107) );
  XOR U40053 ( .A(a[947]), .B(n42197), .Z(n39096) );
  NANDN U40054 ( .A(n39096), .B(n42173), .Z(n39057) );
  NANDN U40055 ( .A(n39055), .B(n42172), .Z(n39056) );
  NAND U40056 ( .A(n39057), .B(n39056), .Z(n39105) );
  NAND U40057 ( .A(b[7]), .B(a[943]), .Z(n39106) );
  XNOR U40058 ( .A(n39105), .B(n39106), .Z(n39108) );
  XOR U40059 ( .A(n39107), .B(n39108), .Z(n39114) );
  NANDN U40060 ( .A(n39058), .B(n42093), .Z(n39060) );
  XOR U40061 ( .A(n42134), .B(a[949]), .Z(n39099) );
  NANDN U40062 ( .A(n39099), .B(n42095), .Z(n39059) );
  NAND U40063 ( .A(n39060), .B(n39059), .Z(n39112) );
  NANDN U40064 ( .A(n39061), .B(n42231), .Z(n39063) );
  XOR U40065 ( .A(n240), .B(a[945]), .Z(n39102) );
  NANDN U40066 ( .A(n39102), .B(n42234), .Z(n39062) );
  AND U40067 ( .A(n39063), .B(n39062), .Z(n39111) );
  XNOR U40068 ( .A(n39112), .B(n39111), .Z(n39113) );
  XNOR U40069 ( .A(n39114), .B(n39113), .Z(n39118) );
  NANDN U40070 ( .A(n39065), .B(n39064), .Z(n39069) );
  NAND U40071 ( .A(n39067), .B(n39066), .Z(n39068) );
  AND U40072 ( .A(n39069), .B(n39068), .Z(n39117) );
  XOR U40073 ( .A(n39118), .B(n39117), .Z(n39119) );
  NANDN U40074 ( .A(n39071), .B(n39070), .Z(n39075) );
  NANDN U40075 ( .A(n39073), .B(n39072), .Z(n39074) );
  NAND U40076 ( .A(n39075), .B(n39074), .Z(n39120) );
  XOR U40077 ( .A(n39119), .B(n39120), .Z(n39087) );
  OR U40078 ( .A(n39077), .B(n39076), .Z(n39081) );
  NANDN U40079 ( .A(n39079), .B(n39078), .Z(n39080) );
  NAND U40080 ( .A(n39081), .B(n39080), .Z(n39088) );
  XNOR U40081 ( .A(n39087), .B(n39088), .Z(n39089) );
  XNOR U40082 ( .A(n39090), .B(n39089), .Z(n39123) );
  XNOR U40083 ( .A(n39123), .B(sreg[1967]), .Z(n39125) );
  NAND U40084 ( .A(n39082), .B(sreg[1966]), .Z(n39086) );
  OR U40085 ( .A(n39084), .B(n39083), .Z(n39085) );
  AND U40086 ( .A(n39086), .B(n39085), .Z(n39124) );
  XOR U40087 ( .A(n39125), .B(n39124), .Z(c[1967]) );
  NANDN U40088 ( .A(n39088), .B(n39087), .Z(n39092) );
  NAND U40089 ( .A(n39090), .B(n39089), .Z(n39091) );
  NAND U40090 ( .A(n39092), .B(n39091), .Z(n39131) );
  NAND U40091 ( .A(b[0]), .B(a[952]), .Z(n39093) );
  XNOR U40092 ( .A(b[1]), .B(n39093), .Z(n39095) );
  NAND U40093 ( .A(n151), .B(a[951]), .Z(n39094) );
  AND U40094 ( .A(n39095), .B(n39094), .Z(n39148) );
  XOR U40095 ( .A(a[948]), .B(n42197), .Z(n39137) );
  NANDN U40096 ( .A(n39137), .B(n42173), .Z(n39098) );
  NANDN U40097 ( .A(n39096), .B(n42172), .Z(n39097) );
  NAND U40098 ( .A(n39098), .B(n39097), .Z(n39146) );
  NAND U40099 ( .A(b[7]), .B(a[944]), .Z(n39147) );
  XNOR U40100 ( .A(n39146), .B(n39147), .Z(n39149) );
  XOR U40101 ( .A(n39148), .B(n39149), .Z(n39155) );
  NANDN U40102 ( .A(n39099), .B(n42093), .Z(n39101) );
  XOR U40103 ( .A(n42134), .B(a[950]), .Z(n39140) );
  NANDN U40104 ( .A(n39140), .B(n42095), .Z(n39100) );
  NAND U40105 ( .A(n39101), .B(n39100), .Z(n39153) );
  NANDN U40106 ( .A(n39102), .B(n42231), .Z(n39104) );
  XOR U40107 ( .A(n240), .B(a[946]), .Z(n39143) );
  NANDN U40108 ( .A(n39143), .B(n42234), .Z(n39103) );
  AND U40109 ( .A(n39104), .B(n39103), .Z(n39152) );
  XNOR U40110 ( .A(n39153), .B(n39152), .Z(n39154) );
  XNOR U40111 ( .A(n39155), .B(n39154), .Z(n39159) );
  NANDN U40112 ( .A(n39106), .B(n39105), .Z(n39110) );
  NAND U40113 ( .A(n39108), .B(n39107), .Z(n39109) );
  AND U40114 ( .A(n39110), .B(n39109), .Z(n39158) );
  XOR U40115 ( .A(n39159), .B(n39158), .Z(n39160) );
  NANDN U40116 ( .A(n39112), .B(n39111), .Z(n39116) );
  NANDN U40117 ( .A(n39114), .B(n39113), .Z(n39115) );
  NAND U40118 ( .A(n39116), .B(n39115), .Z(n39161) );
  XOR U40119 ( .A(n39160), .B(n39161), .Z(n39128) );
  OR U40120 ( .A(n39118), .B(n39117), .Z(n39122) );
  NANDN U40121 ( .A(n39120), .B(n39119), .Z(n39121) );
  NAND U40122 ( .A(n39122), .B(n39121), .Z(n39129) );
  XNOR U40123 ( .A(n39128), .B(n39129), .Z(n39130) );
  XNOR U40124 ( .A(n39131), .B(n39130), .Z(n39164) );
  XNOR U40125 ( .A(n39164), .B(sreg[1968]), .Z(n39166) );
  NAND U40126 ( .A(n39123), .B(sreg[1967]), .Z(n39127) );
  OR U40127 ( .A(n39125), .B(n39124), .Z(n39126) );
  AND U40128 ( .A(n39127), .B(n39126), .Z(n39165) );
  XOR U40129 ( .A(n39166), .B(n39165), .Z(c[1968]) );
  NANDN U40130 ( .A(n39129), .B(n39128), .Z(n39133) );
  NAND U40131 ( .A(n39131), .B(n39130), .Z(n39132) );
  NAND U40132 ( .A(n39133), .B(n39132), .Z(n39172) );
  NAND U40133 ( .A(b[0]), .B(a[953]), .Z(n39134) );
  XNOR U40134 ( .A(b[1]), .B(n39134), .Z(n39136) );
  NAND U40135 ( .A(n151), .B(a[952]), .Z(n39135) );
  AND U40136 ( .A(n39136), .B(n39135), .Z(n39189) );
  XOR U40137 ( .A(a[949]), .B(n42197), .Z(n39178) );
  NANDN U40138 ( .A(n39178), .B(n42173), .Z(n39139) );
  NANDN U40139 ( .A(n39137), .B(n42172), .Z(n39138) );
  NAND U40140 ( .A(n39139), .B(n39138), .Z(n39187) );
  NAND U40141 ( .A(b[7]), .B(a[945]), .Z(n39188) );
  XNOR U40142 ( .A(n39187), .B(n39188), .Z(n39190) );
  XOR U40143 ( .A(n39189), .B(n39190), .Z(n39196) );
  NANDN U40144 ( .A(n39140), .B(n42093), .Z(n39142) );
  XOR U40145 ( .A(n42134), .B(a[951]), .Z(n39181) );
  NANDN U40146 ( .A(n39181), .B(n42095), .Z(n39141) );
  NAND U40147 ( .A(n39142), .B(n39141), .Z(n39194) );
  NANDN U40148 ( .A(n39143), .B(n42231), .Z(n39145) );
  XOR U40149 ( .A(n241), .B(a[947]), .Z(n39184) );
  NANDN U40150 ( .A(n39184), .B(n42234), .Z(n39144) );
  AND U40151 ( .A(n39145), .B(n39144), .Z(n39193) );
  XNOR U40152 ( .A(n39194), .B(n39193), .Z(n39195) );
  XNOR U40153 ( .A(n39196), .B(n39195), .Z(n39200) );
  NANDN U40154 ( .A(n39147), .B(n39146), .Z(n39151) );
  NAND U40155 ( .A(n39149), .B(n39148), .Z(n39150) );
  AND U40156 ( .A(n39151), .B(n39150), .Z(n39199) );
  XOR U40157 ( .A(n39200), .B(n39199), .Z(n39201) );
  NANDN U40158 ( .A(n39153), .B(n39152), .Z(n39157) );
  NANDN U40159 ( .A(n39155), .B(n39154), .Z(n39156) );
  NAND U40160 ( .A(n39157), .B(n39156), .Z(n39202) );
  XOR U40161 ( .A(n39201), .B(n39202), .Z(n39169) );
  OR U40162 ( .A(n39159), .B(n39158), .Z(n39163) );
  NANDN U40163 ( .A(n39161), .B(n39160), .Z(n39162) );
  NAND U40164 ( .A(n39163), .B(n39162), .Z(n39170) );
  XNOR U40165 ( .A(n39169), .B(n39170), .Z(n39171) );
  XNOR U40166 ( .A(n39172), .B(n39171), .Z(n39205) );
  XNOR U40167 ( .A(n39205), .B(sreg[1969]), .Z(n39207) );
  NAND U40168 ( .A(n39164), .B(sreg[1968]), .Z(n39168) );
  OR U40169 ( .A(n39166), .B(n39165), .Z(n39167) );
  AND U40170 ( .A(n39168), .B(n39167), .Z(n39206) );
  XOR U40171 ( .A(n39207), .B(n39206), .Z(c[1969]) );
  NANDN U40172 ( .A(n39170), .B(n39169), .Z(n39174) );
  NAND U40173 ( .A(n39172), .B(n39171), .Z(n39173) );
  NAND U40174 ( .A(n39174), .B(n39173), .Z(n39213) );
  NAND U40175 ( .A(b[0]), .B(a[954]), .Z(n39175) );
  XNOR U40176 ( .A(b[1]), .B(n39175), .Z(n39177) );
  NAND U40177 ( .A(n151), .B(a[953]), .Z(n39176) );
  AND U40178 ( .A(n39177), .B(n39176), .Z(n39230) );
  XOR U40179 ( .A(a[950]), .B(n42197), .Z(n39219) );
  NANDN U40180 ( .A(n39219), .B(n42173), .Z(n39180) );
  NANDN U40181 ( .A(n39178), .B(n42172), .Z(n39179) );
  NAND U40182 ( .A(n39180), .B(n39179), .Z(n39228) );
  NAND U40183 ( .A(b[7]), .B(a[946]), .Z(n39229) );
  XNOR U40184 ( .A(n39228), .B(n39229), .Z(n39231) );
  XOR U40185 ( .A(n39230), .B(n39231), .Z(n39237) );
  NANDN U40186 ( .A(n39181), .B(n42093), .Z(n39183) );
  XOR U40187 ( .A(n42134), .B(a[952]), .Z(n39222) );
  NANDN U40188 ( .A(n39222), .B(n42095), .Z(n39182) );
  NAND U40189 ( .A(n39183), .B(n39182), .Z(n39235) );
  NANDN U40190 ( .A(n39184), .B(n42231), .Z(n39186) );
  XOR U40191 ( .A(n241), .B(a[948]), .Z(n39225) );
  NANDN U40192 ( .A(n39225), .B(n42234), .Z(n39185) );
  AND U40193 ( .A(n39186), .B(n39185), .Z(n39234) );
  XNOR U40194 ( .A(n39235), .B(n39234), .Z(n39236) );
  XNOR U40195 ( .A(n39237), .B(n39236), .Z(n39241) );
  NANDN U40196 ( .A(n39188), .B(n39187), .Z(n39192) );
  NAND U40197 ( .A(n39190), .B(n39189), .Z(n39191) );
  AND U40198 ( .A(n39192), .B(n39191), .Z(n39240) );
  XOR U40199 ( .A(n39241), .B(n39240), .Z(n39242) );
  NANDN U40200 ( .A(n39194), .B(n39193), .Z(n39198) );
  NANDN U40201 ( .A(n39196), .B(n39195), .Z(n39197) );
  NAND U40202 ( .A(n39198), .B(n39197), .Z(n39243) );
  XOR U40203 ( .A(n39242), .B(n39243), .Z(n39210) );
  OR U40204 ( .A(n39200), .B(n39199), .Z(n39204) );
  NANDN U40205 ( .A(n39202), .B(n39201), .Z(n39203) );
  NAND U40206 ( .A(n39204), .B(n39203), .Z(n39211) );
  XNOR U40207 ( .A(n39210), .B(n39211), .Z(n39212) );
  XNOR U40208 ( .A(n39213), .B(n39212), .Z(n39246) );
  XNOR U40209 ( .A(n39246), .B(sreg[1970]), .Z(n39248) );
  NAND U40210 ( .A(n39205), .B(sreg[1969]), .Z(n39209) );
  OR U40211 ( .A(n39207), .B(n39206), .Z(n39208) );
  AND U40212 ( .A(n39209), .B(n39208), .Z(n39247) );
  XOR U40213 ( .A(n39248), .B(n39247), .Z(c[1970]) );
  NANDN U40214 ( .A(n39211), .B(n39210), .Z(n39215) );
  NAND U40215 ( .A(n39213), .B(n39212), .Z(n39214) );
  NAND U40216 ( .A(n39215), .B(n39214), .Z(n39254) );
  NAND U40217 ( .A(b[0]), .B(a[955]), .Z(n39216) );
  XNOR U40218 ( .A(b[1]), .B(n39216), .Z(n39218) );
  NAND U40219 ( .A(n151), .B(a[954]), .Z(n39217) );
  AND U40220 ( .A(n39218), .B(n39217), .Z(n39271) );
  XOR U40221 ( .A(a[951]), .B(n42197), .Z(n39260) );
  NANDN U40222 ( .A(n39260), .B(n42173), .Z(n39221) );
  NANDN U40223 ( .A(n39219), .B(n42172), .Z(n39220) );
  NAND U40224 ( .A(n39221), .B(n39220), .Z(n39269) );
  NAND U40225 ( .A(b[7]), .B(a[947]), .Z(n39270) );
  XNOR U40226 ( .A(n39269), .B(n39270), .Z(n39272) );
  XOR U40227 ( .A(n39271), .B(n39272), .Z(n39278) );
  NANDN U40228 ( .A(n39222), .B(n42093), .Z(n39224) );
  XOR U40229 ( .A(n42134), .B(a[953]), .Z(n39263) );
  NANDN U40230 ( .A(n39263), .B(n42095), .Z(n39223) );
  NAND U40231 ( .A(n39224), .B(n39223), .Z(n39276) );
  NANDN U40232 ( .A(n39225), .B(n42231), .Z(n39227) );
  XOR U40233 ( .A(n241), .B(a[949]), .Z(n39266) );
  NANDN U40234 ( .A(n39266), .B(n42234), .Z(n39226) );
  AND U40235 ( .A(n39227), .B(n39226), .Z(n39275) );
  XNOR U40236 ( .A(n39276), .B(n39275), .Z(n39277) );
  XNOR U40237 ( .A(n39278), .B(n39277), .Z(n39282) );
  NANDN U40238 ( .A(n39229), .B(n39228), .Z(n39233) );
  NAND U40239 ( .A(n39231), .B(n39230), .Z(n39232) );
  AND U40240 ( .A(n39233), .B(n39232), .Z(n39281) );
  XOR U40241 ( .A(n39282), .B(n39281), .Z(n39283) );
  NANDN U40242 ( .A(n39235), .B(n39234), .Z(n39239) );
  NANDN U40243 ( .A(n39237), .B(n39236), .Z(n39238) );
  NAND U40244 ( .A(n39239), .B(n39238), .Z(n39284) );
  XOR U40245 ( .A(n39283), .B(n39284), .Z(n39251) );
  OR U40246 ( .A(n39241), .B(n39240), .Z(n39245) );
  NANDN U40247 ( .A(n39243), .B(n39242), .Z(n39244) );
  NAND U40248 ( .A(n39245), .B(n39244), .Z(n39252) );
  XNOR U40249 ( .A(n39251), .B(n39252), .Z(n39253) );
  XNOR U40250 ( .A(n39254), .B(n39253), .Z(n39287) );
  XNOR U40251 ( .A(n39287), .B(sreg[1971]), .Z(n39289) );
  NAND U40252 ( .A(n39246), .B(sreg[1970]), .Z(n39250) );
  OR U40253 ( .A(n39248), .B(n39247), .Z(n39249) );
  AND U40254 ( .A(n39250), .B(n39249), .Z(n39288) );
  XOR U40255 ( .A(n39289), .B(n39288), .Z(c[1971]) );
  NANDN U40256 ( .A(n39252), .B(n39251), .Z(n39256) );
  NAND U40257 ( .A(n39254), .B(n39253), .Z(n39255) );
  NAND U40258 ( .A(n39256), .B(n39255), .Z(n39295) );
  NAND U40259 ( .A(b[0]), .B(a[956]), .Z(n39257) );
  XNOR U40260 ( .A(b[1]), .B(n39257), .Z(n39259) );
  NAND U40261 ( .A(n151), .B(a[955]), .Z(n39258) );
  AND U40262 ( .A(n39259), .B(n39258), .Z(n39312) );
  XOR U40263 ( .A(a[952]), .B(n42197), .Z(n39301) );
  NANDN U40264 ( .A(n39301), .B(n42173), .Z(n39262) );
  NANDN U40265 ( .A(n39260), .B(n42172), .Z(n39261) );
  NAND U40266 ( .A(n39262), .B(n39261), .Z(n39310) );
  NAND U40267 ( .A(b[7]), .B(a[948]), .Z(n39311) );
  XNOR U40268 ( .A(n39310), .B(n39311), .Z(n39313) );
  XOR U40269 ( .A(n39312), .B(n39313), .Z(n39319) );
  NANDN U40270 ( .A(n39263), .B(n42093), .Z(n39265) );
  XOR U40271 ( .A(n42134), .B(a[954]), .Z(n39304) );
  NANDN U40272 ( .A(n39304), .B(n42095), .Z(n39264) );
  NAND U40273 ( .A(n39265), .B(n39264), .Z(n39317) );
  NANDN U40274 ( .A(n39266), .B(n42231), .Z(n39268) );
  XOR U40275 ( .A(n241), .B(a[950]), .Z(n39307) );
  NANDN U40276 ( .A(n39307), .B(n42234), .Z(n39267) );
  AND U40277 ( .A(n39268), .B(n39267), .Z(n39316) );
  XNOR U40278 ( .A(n39317), .B(n39316), .Z(n39318) );
  XNOR U40279 ( .A(n39319), .B(n39318), .Z(n39323) );
  NANDN U40280 ( .A(n39270), .B(n39269), .Z(n39274) );
  NAND U40281 ( .A(n39272), .B(n39271), .Z(n39273) );
  AND U40282 ( .A(n39274), .B(n39273), .Z(n39322) );
  XOR U40283 ( .A(n39323), .B(n39322), .Z(n39324) );
  NANDN U40284 ( .A(n39276), .B(n39275), .Z(n39280) );
  NANDN U40285 ( .A(n39278), .B(n39277), .Z(n39279) );
  NAND U40286 ( .A(n39280), .B(n39279), .Z(n39325) );
  XOR U40287 ( .A(n39324), .B(n39325), .Z(n39292) );
  OR U40288 ( .A(n39282), .B(n39281), .Z(n39286) );
  NANDN U40289 ( .A(n39284), .B(n39283), .Z(n39285) );
  NAND U40290 ( .A(n39286), .B(n39285), .Z(n39293) );
  XNOR U40291 ( .A(n39292), .B(n39293), .Z(n39294) );
  XNOR U40292 ( .A(n39295), .B(n39294), .Z(n39328) );
  XNOR U40293 ( .A(n39328), .B(sreg[1972]), .Z(n39330) );
  NAND U40294 ( .A(n39287), .B(sreg[1971]), .Z(n39291) );
  OR U40295 ( .A(n39289), .B(n39288), .Z(n39290) );
  AND U40296 ( .A(n39291), .B(n39290), .Z(n39329) );
  XOR U40297 ( .A(n39330), .B(n39329), .Z(c[1972]) );
  NANDN U40298 ( .A(n39293), .B(n39292), .Z(n39297) );
  NAND U40299 ( .A(n39295), .B(n39294), .Z(n39296) );
  NAND U40300 ( .A(n39297), .B(n39296), .Z(n39336) );
  NAND U40301 ( .A(b[0]), .B(a[957]), .Z(n39298) );
  XNOR U40302 ( .A(b[1]), .B(n39298), .Z(n39300) );
  NAND U40303 ( .A(n151), .B(a[956]), .Z(n39299) );
  AND U40304 ( .A(n39300), .B(n39299), .Z(n39353) );
  XOR U40305 ( .A(a[953]), .B(n42197), .Z(n39342) );
  NANDN U40306 ( .A(n39342), .B(n42173), .Z(n39303) );
  NANDN U40307 ( .A(n39301), .B(n42172), .Z(n39302) );
  NAND U40308 ( .A(n39303), .B(n39302), .Z(n39351) );
  NAND U40309 ( .A(b[7]), .B(a[949]), .Z(n39352) );
  XNOR U40310 ( .A(n39351), .B(n39352), .Z(n39354) );
  XOR U40311 ( .A(n39353), .B(n39354), .Z(n39360) );
  NANDN U40312 ( .A(n39304), .B(n42093), .Z(n39306) );
  XOR U40313 ( .A(n42134), .B(a[955]), .Z(n39345) );
  NANDN U40314 ( .A(n39345), .B(n42095), .Z(n39305) );
  NAND U40315 ( .A(n39306), .B(n39305), .Z(n39358) );
  NANDN U40316 ( .A(n39307), .B(n42231), .Z(n39309) );
  XOR U40317 ( .A(n241), .B(a[951]), .Z(n39348) );
  NANDN U40318 ( .A(n39348), .B(n42234), .Z(n39308) );
  AND U40319 ( .A(n39309), .B(n39308), .Z(n39357) );
  XNOR U40320 ( .A(n39358), .B(n39357), .Z(n39359) );
  XNOR U40321 ( .A(n39360), .B(n39359), .Z(n39364) );
  NANDN U40322 ( .A(n39311), .B(n39310), .Z(n39315) );
  NAND U40323 ( .A(n39313), .B(n39312), .Z(n39314) );
  AND U40324 ( .A(n39315), .B(n39314), .Z(n39363) );
  XOR U40325 ( .A(n39364), .B(n39363), .Z(n39365) );
  NANDN U40326 ( .A(n39317), .B(n39316), .Z(n39321) );
  NANDN U40327 ( .A(n39319), .B(n39318), .Z(n39320) );
  NAND U40328 ( .A(n39321), .B(n39320), .Z(n39366) );
  XOR U40329 ( .A(n39365), .B(n39366), .Z(n39333) );
  OR U40330 ( .A(n39323), .B(n39322), .Z(n39327) );
  NANDN U40331 ( .A(n39325), .B(n39324), .Z(n39326) );
  NAND U40332 ( .A(n39327), .B(n39326), .Z(n39334) );
  XNOR U40333 ( .A(n39333), .B(n39334), .Z(n39335) );
  XNOR U40334 ( .A(n39336), .B(n39335), .Z(n39369) );
  XNOR U40335 ( .A(n39369), .B(sreg[1973]), .Z(n39371) );
  NAND U40336 ( .A(n39328), .B(sreg[1972]), .Z(n39332) );
  OR U40337 ( .A(n39330), .B(n39329), .Z(n39331) );
  AND U40338 ( .A(n39332), .B(n39331), .Z(n39370) );
  XOR U40339 ( .A(n39371), .B(n39370), .Z(c[1973]) );
  NANDN U40340 ( .A(n39334), .B(n39333), .Z(n39338) );
  NAND U40341 ( .A(n39336), .B(n39335), .Z(n39337) );
  NAND U40342 ( .A(n39338), .B(n39337), .Z(n39377) );
  NAND U40343 ( .A(b[0]), .B(a[958]), .Z(n39339) );
  XNOR U40344 ( .A(b[1]), .B(n39339), .Z(n39341) );
  NAND U40345 ( .A(n151), .B(a[957]), .Z(n39340) );
  AND U40346 ( .A(n39341), .B(n39340), .Z(n39394) );
  XOR U40347 ( .A(a[954]), .B(n42197), .Z(n39383) );
  NANDN U40348 ( .A(n39383), .B(n42173), .Z(n39344) );
  NANDN U40349 ( .A(n39342), .B(n42172), .Z(n39343) );
  NAND U40350 ( .A(n39344), .B(n39343), .Z(n39392) );
  NAND U40351 ( .A(b[7]), .B(a[950]), .Z(n39393) );
  XNOR U40352 ( .A(n39392), .B(n39393), .Z(n39395) );
  XOR U40353 ( .A(n39394), .B(n39395), .Z(n39401) );
  NANDN U40354 ( .A(n39345), .B(n42093), .Z(n39347) );
  XOR U40355 ( .A(n42134), .B(a[956]), .Z(n39386) );
  NANDN U40356 ( .A(n39386), .B(n42095), .Z(n39346) );
  NAND U40357 ( .A(n39347), .B(n39346), .Z(n39399) );
  NANDN U40358 ( .A(n39348), .B(n42231), .Z(n39350) );
  XOR U40359 ( .A(n241), .B(a[952]), .Z(n39389) );
  NANDN U40360 ( .A(n39389), .B(n42234), .Z(n39349) );
  AND U40361 ( .A(n39350), .B(n39349), .Z(n39398) );
  XNOR U40362 ( .A(n39399), .B(n39398), .Z(n39400) );
  XNOR U40363 ( .A(n39401), .B(n39400), .Z(n39405) );
  NANDN U40364 ( .A(n39352), .B(n39351), .Z(n39356) );
  NAND U40365 ( .A(n39354), .B(n39353), .Z(n39355) );
  AND U40366 ( .A(n39356), .B(n39355), .Z(n39404) );
  XOR U40367 ( .A(n39405), .B(n39404), .Z(n39406) );
  NANDN U40368 ( .A(n39358), .B(n39357), .Z(n39362) );
  NANDN U40369 ( .A(n39360), .B(n39359), .Z(n39361) );
  NAND U40370 ( .A(n39362), .B(n39361), .Z(n39407) );
  XOR U40371 ( .A(n39406), .B(n39407), .Z(n39374) );
  OR U40372 ( .A(n39364), .B(n39363), .Z(n39368) );
  NANDN U40373 ( .A(n39366), .B(n39365), .Z(n39367) );
  NAND U40374 ( .A(n39368), .B(n39367), .Z(n39375) );
  XNOR U40375 ( .A(n39374), .B(n39375), .Z(n39376) );
  XNOR U40376 ( .A(n39377), .B(n39376), .Z(n39410) );
  XNOR U40377 ( .A(n39410), .B(sreg[1974]), .Z(n39412) );
  NAND U40378 ( .A(n39369), .B(sreg[1973]), .Z(n39373) );
  OR U40379 ( .A(n39371), .B(n39370), .Z(n39372) );
  AND U40380 ( .A(n39373), .B(n39372), .Z(n39411) );
  XOR U40381 ( .A(n39412), .B(n39411), .Z(c[1974]) );
  NANDN U40382 ( .A(n39375), .B(n39374), .Z(n39379) );
  NAND U40383 ( .A(n39377), .B(n39376), .Z(n39378) );
  NAND U40384 ( .A(n39379), .B(n39378), .Z(n39418) );
  NAND U40385 ( .A(b[0]), .B(a[959]), .Z(n39380) );
  XNOR U40386 ( .A(b[1]), .B(n39380), .Z(n39382) );
  NAND U40387 ( .A(n152), .B(a[958]), .Z(n39381) );
  AND U40388 ( .A(n39382), .B(n39381), .Z(n39435) );
  XOR U40389 ( .A(a[955]), .B(n42197), .Z(n39424) );
  NANDN U40390 ( .A(n39424), .B(n42173), .Z(n39385) );
  NANDN U40391 ( .A(n39383), .B(n42172), .Z(n39384) );
  NAND U40392 ( .A(n39385), .B(n39384), .Z(n39433) );
  NAND U40393 ( .A(b[7]), .B(a[951]), .Z(n39434) );
  XNOR U40394 ( .A(n39433), .B(n39434), .Z(n39436) );
  XOR U40395 ( .A(n39435), .B(n39436), .Z(n39442) );
  NANDN U40396 ( .A(n39386), .B(n42093), .Z(n39388) );
  XOR U40397 ( .A(n42134), .B(a[957]), .Z(n39427) );
  NANDN U40398 ( .A(n39427), .B(n42095), .Z(n39387) );
  NAND U40399 ( .A(n39388), .B(n39387), .Z(n39440) );
  NANDN U40400 ( .A(n39389), .B(n42231), .Z(n39391) );
  XOR U40401 ( .A(n241), .B(a[953]), .Z(n39430) );
  NANDN U40402 ( .A(n39430), .B(n42234), .Z(n39390) );
  AND U40403 ( .A(n39391), .B(n39390), .Z(n39439) );
  XNOR U40404 ( .A(n39440), .B(n39439), .Z(n39441) );
  XNOR U40405 ( .A(n39442), .B(n39441), .Z(n39446) );
  NANDN U40406 ( .A(n39393), .B(n39392), .Z(n39397) );
  NAND U40407 ( .A(n39395), .B(n39394), .Z(n39396) );
  AND U40408 ( .A(n39397), .B(n39396), .Z(n39445) );
  XOR U40409 ( .A(n39446), .B(n39445), .Z(n39447) );
  NANDN U40410 ( .A(n39399), .B(n39398), .Z(n39403) );
  NANDN U40411 ( .A(n39401), .B(n39400), .Z(n39402) );
  NAND U40412 ( .A(n39403), .B(n39402), .Z(n39448) );
  XOR U40413 ( .A(n39447), .B(n39448), .Z(n39415) );
  OR U40414 ( .A(n39405), .B(n39404), .Z(n39409) );
  NANDN U40415 ( .A(n39407), .B(n39406), .Z(n39408) );
  NAND U40416 ( .A(n39409), .B(n39408), .Z(n39416) );
  XNOR U40417 ( .A(n39415), .B(n39416), .Z(n39417) );
  XNOR U40418 ( .A(n39418), .B(n39417), .Z(n39451) );
  XNOR U40419 ( .A(n39451), .B(sreg[1975]), .Z(n39453) );
  NAND U40420 ( .A(n39410), .B(sreg[1974]), .Z(n39414) );
  OR U40421 ( .A(n39412), .B(n39411), .Z(n39413) );
  AND U40422 ( .A(n39414), .B(n39413), .Z(n39452) );
  XOR U40423 ( .A(n39453), .B(n39452), .Z(c[1975]) );
  NANDN U40424 ( .A(n39416), .B(n39415), .Z(n39420) );
  NAND U40425 ( .A(n39418), .B(n39417), .Z(n39419) );
  NAND U40426 ( .A(n39420), .B(n39419), .Z(n39459) );
  NAND U40427 ( .A(b[0]), .B(a[960]), .Z(n39421) );
  XNOR U40428 ( .A(b[1]), .B(n39421), .Z(n39423) );
  NAND U40429 ( .A(n152), .B(a[959]), .Z(n39422) );
  AND U40430 ( .A(n39423), .B(n39422), .Z(n39476) );
  XOR U40431 ( .A(a[956]), .B(n42197), .Z(n39465) );
  NANDN U40432 ( .A(n39465), .B(n42173), .Z(n39426) );
  NANDN U40433 ( .A(n39424), .B(n42172), .Z(n39425) );
  NAND U40434 ( .A(n39426), .B(n39425), .Z(n39474) );
  NAND U40435 ( .A(b[7]), .B(a[952]), .Z(n39475) );
  XNOR U40436 ( .A(n39474), .B(n39475), .Z(n39477) );
  XOR U40437 ( .A(n39476), .B(n39477), .Z(n39483) );
  NANDN U40438 ( .A(n39427), .B(n42093), .Z(n39429) );
  XOR U40439 ( .A(n42134), .B(a[958]), .Z(n39468) );
  NANDN U40440 ( .A(n39468), .B(n42095), .Z(n39428) );
  NAND U40441 ( .A(n39429), .B(n39428), .Z(n39481) );
  NANDN U40442 ( .A(n39430), .B(n42231), .Z(n39432) );
  XOR U40443 ( .A(n241), .B(a[954]), .Z(n39471) );
  NANDN U40444 ( .A(n39471), .B(n42234), .Z(n39431) );
  AND U40445 ( .A(n39432), .B(n39431), .Z(n39480) );
  XNOR U40446 ( .A(n39481), .B(n39480), .Z(n39482) );
  XNOR U40447 ( .A(n39483), .B(n39482), .Z(n39487) );
  NANDN U40448 ( .A(n39434), .B(n39433), .Z(n39438) );
  NAND U40449 ( .A(n39436), .B(n39435), .Z(n39437) );
  AND U40450 ( .A(n39438), .B(n39437), .Z(n39486) );
  XOR U40451 ( .A(n39487), .B(n39486), .Z(n39488) );
  NANDN U40452 ( .A(n39440), .B(n39439), .Z(n39444) );
  NANDN U40453 ( .A(n39442), .B(n39441), .Z(n39443) );
  NAND U40454 ( .A(n39444), .B(n39443), .Z(n39489) );
  XOR U40455 ( .A(n39488), .B(n39489), .Z(n39456) );
  OR U40456 ( .A(n39446), .B(n39445), .Z(n39450) );
  NANDN U40457 ( .A(n39448), .B(n39447), .Z(n39449) );
  NAND U40458 ( .A(n39450), .B(n39449), .Z(n39457) );
  XNOR U40459 ( .A(n39456), .B(n39457), .Z(n39458) );
  XNOR U40460 ( .A(n39459), .B(n39458), .Z(n39492) );
  XNOR U40461 ( .A(n39492), .B(sreg[1976]), .Z(n39494) );
  NAND U40462 ( .A(n39451), .B(sreg[1975]), .Z(n39455) );
  OR U40463 ( .A(n39453), .B(n39452), .Z(n39454) );
  AND U40464 ( .A(n39455), .B(n39454), .Z(n39493) );
  XOR U40465 ( .A(n39494), .B(n39493), .Z(c[1976]) );
  NANDN U40466 ( .A(n39457), .B(n39456), .Z(n39461) );
  NAND U40467 ( .A(n39459), .B(n39458), .Z(n39460) );
  NAND U40468 ( .A(n39461), .B(n39460), .Z(n39500) );
  NAND U40469 ( .A(b[0]), .B(a[961]), .Z(n39462) );
  XNOR U40470 ( .A(b[1]), .B(n39462), .Z(n39464) );
  NAND U40471 ( .A(n152), .B(a[960]), .Z(n39463) );
  AND U40472 ( .A(n39464), .B(n39463), .Z(n39517) );
  XOR U40473 ( .A(a[957]), .B(n42197), .Z(n39506) );
  NANDN U40474 ( .A(n39506), .B(n42173), .Z(n39467) );
  NANDN U40475 ( .A(n39465), .B(n42172), .Z(n39466) );
  NAND U40476 ( .A(n39467), .B(n39466), .Z(n39515) );
  NAND U40477 ( .A(b[7]), .B(a[953]), .Z(n39516) );
  XNOR U40478 ( .A(n39515), .B(n39516), .Z(n39518) );
  XOR U40479 ( .A(n39517), .B(n39518), .Z(n39524) );
  NANDN U40480 ( .A(n39468), .B(n42093), .Z(n39470) );
  XOR U40481 ( .A(n42134), .B(a[959]), .Z(n39509) );
  NANDN U40482 ( .A(n39509), .B(n42095), .Z(n39469) );
  NAND U40483 ( .A(n39470), .B(n39469), .Z(n39522) );
  NANDN U40484 ( .A(n39471), .B(n42231), .Z(n39473) );
  XOR U40485 ( .A(n241), .B(a[955]), .Z(n39512) );
  NANDN U40486 ( .A(n39512), .B(n42234), .Z(n39472) );
  AND U40487 ( .A(n39473), .B(n39472), .Z(n39521) );
  XNOR U40488 ( .A(n39522), .B(n39521), .Z(n39523) );
  XNOR U40489 ( .A(n39524), .B(n39523), .Z(n39528) );
  NANDN U40490 ( .A(n39475), .B(n39474), .Z(n39479) );
  NAND U40491 ( .A(n39477), .B(n39476), .Z(n39478) );
  AND U40492 ( .A(n39479), .B(n39478), .Z(n39527) );
  XOR U40493 ( .A(n39528), .B(n39527), .Z(n39529) );
  NANDN U40494 ( .A(n39481), .B(n39480), .Z(n39485) );
  NANDN U40495 ( .A(n39483), .B(n39482), .Z(n39484) );
  NAND U40496 ( .A(n39485), .B(n39484), .Z(n39530) );
  XOR U40497 ( .A(n39529), .B(n39530), .Z(n39497) );
  OR U40498 ( .A(n39487), .B(n39486), .Z(n39491) );
  NANDN U40499 ( .A(n39489), .B(n39488), .Z(n39490) );
  NAND U40500 ( .A(n39491), .B(n39490), .Z(n39498) );
  XNOR U40501 ( .A(n39497), .B(n39498), .Z(n39499) );
  XNOR U40502 ( .A(n39500), .B(n39499), .Z(n39533) );
  XNOR U40503 ( .A(n39533), .B(sreg[1977]), .Z(n39535) );
  NAND U40504 ( .A(n39492), .B(sreg[1976]), .Z(n39496) );
  OR U40505 ( .A(n39494), .B(n39493), .Z(n39495) );
  AND U40506 ( .A(n39496), .B(n39495), .Z(n39534) );
  XOR U40507 ( .A(n39535), .B(n39534), .Z(c[1977]) );
  NANDN U40508 ( .A(n39498), .B(n39497), .Z(n39502) );
  NAND U40509 ( .A(n39500), .B(n39499), .Z(n39501) );
  NAND U40510 ( .A(n39502), .B(n39501), .Z(n39541) );
  NAND U40511 ( .A(b[0]), .B(a[962]), .Z(n39503) );
  XNOR U40512 ( .A(b[1]), .B(n39503), .Z(n39505) );
  NAND U40513 ( .A(n152), .B(a[961]), .Z(n39504) );
  AND U40514 ( .A(n39505), .B(n39504), .Z(n39558) );
  XOR U40515 ( .A(a[958]), .B(n42197), .Z(n39547) );
  NANDN U40516 ( .A(n39547), .B(n42173), .Z(n39508) );
  NANDN U40517 ( .A(n39506), .B(n42172), .Z(n39507) );
  NAND U40518 ( .A(n39508), .B(n39507), .Z(n39556) );
  NAND U40519 ( .A(b[7]), .B(a[954]), .Z(n39557) );
  XNOR U40520 ( .A(n39556), .B(n39557), .Z(n39559) );
  XOR U40521 ( .A(n39558), .B(n39559), .Z(n39565) );
  NANDN U40522 ( .A(n39509), .B(n42093), .Z(n39511) );
  XOR U40523 ( .A(n42134), .B(a[960]), .Z(n39550) );
  NANDN U40524 ( .A(n39550), .B(n42095), .Z(n39510) );
  NAND U40525 ( .A(n39511), .B(n39510), .Z(n39563) );
  NANDN U40526 ( .A(n39512), .B(n42231), .Z(n39514) );
  XOR U40527 ( .A(n241), .B(a[956]), .Z(n39553) );
  NANDN U40528 ( .A(n39553), .B(n42234), .Z(n39513) );
  AND U40529 ( .A(n39514), .B(n39513), .Z(n39562) );
  XNOR U40530 ( .A(n39563), .B(n39562), .Z(n39564) );
  XNOR U40531 ( .A(n39565), .B(n39564), .Z(n39569) );
  NANDN U40532 ( .A(n39516), .B(n39515), .Z(n39520) );
  NAND U40533 ( .A(n39518), .B(n39517), .Z(n39519) );
  AND U40534 ( .A(n39520), .B(n39519), .Z(n39568) );
  XOR U40535 ( .A(n39569), .B(n39568), .Z(n39570) );
  NANDN U40536 ( .A(n39522), .B(n39521), .Z(n39526) );
  NANDN U40537 ( .A(n39524), .B(n39523), .Z(n39525) );
  NAND U40538 ( .A(n39526), .B(n39525), .Z(n39571) );
  XOR U40539 ( .A(n39570), .B(n39571), .Z(n39538) );
  OR U40540 ( .A(n39528), .B(n39527), .Z(n39532) );
  NANDN U40541 ( .A(n39530), .B(n39529), .Z(n39531) );
  NAND U40542 ( .A(n39532), .B(n39531), .Z(n39539) );
  XNOR U40543 ( .A(n39538), .B(n39539), .Z(n39540) );
  XNOR U40544 ( .A(n39541), .B(n39540), .Z(n39574) );
  XNOR U40545 ( .A(n39574), .B(sreg[1978]), .Z(n39576) );
  NAND U40546 ( .A(n39533), .B(sreg[1977]), .Z(n39537) );
  OR U40547 ( .A(n39535), .B(n39534), .Z(n39536) );
  AND U40548 ( .A(n39537), .B(n39536), .Z(n39575) );
  XOR U40549 ( .A(n39576), .B(n39575), .Z(c[1978]) );
  NANDN U40550 ( .A(n39539), .B(n39538), .Z(n39543) );
  NAND U40551 ( .A(n39541), .B(n39540), .Z(n39542) );
  NAND U40552 ( .A(n39543), .B(n39542), .Z(n39582) );
  NAND U40553 ( .A(b[0]), .B(a[963]), .Z(n39544) );
  XNOR U40554 ( .A(b[1]), .B(n39544), .Z(n39546) );
  NAND U40555 ( .A(n152), .B(a[962]), .Z(n39545) );
  AND U40556 ( .A(n39546), .B(n39545), .Z(n39599) );
  XOR U40557 ( .A(a[959]), .B(n42197), .Z(n39588) );
  NANDN U40558 ( .A(n39588), .B(n42173), .Z(n39549) );
  NANDN U40559 ( .A(n39547), .B(n42172), .Z(n39548) );
  NAND U40560 ( .A(n39549), .B(n39548), .Z(n39597) );
  NAND U40561 ( .A(b[7]), .B(a[955]), .Z(n39598) );
  XNOR U40562 ( .A(n39597), .B(n39598), .Z(n39600) );
  XOR U40563 ( .A(n39599), .B(n39600), .Z(n39606) );
  NANDN U40564 ( .A(n39550), .B(n42093), .Z(n39552) );
  XOR U40565 ( .A(n42134), .B(a[961]), .Z(n39591) );
  NANDN U40566 ( .A(n39591), .B(n42095), .Z(n39551) );
  NAND U40567 ( .A(n39552), .B(n39551), .Z(n39604) );
  NANDN U40568 ( .A(n39553), .B(n42231), .Z(n39555) );
  XOR U40569 ( .A(n241), .B(a[957]), .Z(n39594) );
  NANDN U40570 ( .A(n39594), .B(n42234), .Z(n39554) );
  AND U40571 ( .A(n39555), .B(n39554), .Z(n39603) );
  XNOR U40572 ( .A(n39604), .B(n39603), .Z(n39605) );
  XNOR U40573 ( .A(n39606), .B(n39605), .Z(n39610) );
  NANDN U40574 ( .A(n39557), .B(n39556), .Z(n39561) );
  NAND U40575 ( .A(n39559), .B(n39558), .Z(n39560) );
  AND U40576 ( .A(n39561), .B(n39560), .Z(n39609) );
  XOR U40577 ( .A(n39610), .B(n39609), .Z(n39611) );
  NANDN U40578 ( .A(n39563), .B(n39562), .Z(n39567) );
  NANDN U40579 ( .A(n39565), .B(n39564), .Z(n39566) );
  NAND U40580 ( .A(n39567), .B(n39566), .Z(n39612) );
  XOR U40581 ( .A(n39611), .B(n39612), .Z(n39579) );
  OR U40582 ( .A(n39569), .B(n39568), .Z(n39573) );
  NANDN U40583 ( .A(n39571), .B(n39570), .Z(n39572) );
  NAND U40584 ( .A(n39573), .B(n39572), .Z(n39580) );
  XNOR U40585 ( .A(n39579), .B(n39580), .Z(n39581) );
  XNOR U40586 ( .A(n39582), .B(n39581), .Z(n39615) );
  XNOR U40587 ( .A(n39615), .B(sreg[1979]), .Z(n39617) );
  NAND U40588 ( .A(n39574), .B(sreg[1978]), .Z(n39578) );
  OR U40589 ( .A(n39576), .B(n39575), .Z(n39577) );
  AND U40590 ( .A(n39578), .B(n39577), .Z(n39616) );
  XOR U40591 ( .A(n39617), .B(n39616), .Z(c[1979]) );
  NANDN U40592 ( .A(n39580), .B(n39579), .Z(n39584) );
  NAND U40593 ( .A(n39582), .B(n39581), .Z(n39583) );
  NAND U40594 ( .A(n39584), .B(n39583), .Z(n39623) );
  NAND U40595 ( .A(b[0]), .B(a[964]), .Z(n39585) );
  XNOR U40596 ( .A(b[1]), .B(n39585), .Z(n39587) );
  NAND U40597 ( .A(n152), .B(a[963]), .Z(n39586) );
  AND U40598 ( .A(n39587), .B(n39586), .Z(n39640) );
  XOR U40599 ( .A(a[960]), .B(n42197), .Z(n39629) );
  NANDN U40600 ( .A(n39629), .B(n42173), .Z(n39590) );
  NANDN U40601 ( .A(n39588), .B(n42172), .Z(n39589) );
  NAND U40602 ( .A(n39590), .B(n39589), .Z(n39638) );
  NAND U40603 ( .A(b[7]), .B(a[956]), .Z(n39639) );
  XNOR U40604 ( .A(n39638), .B(n39639), .Z(n39641) );
  XOR U40605 ( .A(n39640), .B(n39641), .Z(n39647) );
  NANDN U40606 ( .A(n39591), .B(n42093), .Z(n39593) );
  XOR U40607 ( .A(n42134), .B(a[962]), .Z(n39632) );
  NANDN U40608 ( .A(n39632), .B(n42095), .Z(n39592) );
  NAND U40609 ( .A(n39593), .B(n39592), .Z(n39645) );
  NANDN U40610 ( .A(n39594), .B(n42231), .Z(n39596) );
  XOR U40611 ( .A(n241), .B(a[958]), .Z(n39635) );
  NANDN U40612 ( .A(n39635), .B(n42234), .Z(n39595) );
  AND U40613 ( .A(n39596), .B(n39595), .Z(n39644) );
  XNOR U40614 ( .A(n39645), .B(n39644), .Z(n39646) );
  XNOR U40615 ( .A(n39647), .B(n39646), .Z(n39651) );
  NANDN U40616 ( .A(n39598), .B(n39597), .Z(n39602) );
  NAND U40617 ( .A(n39600), .B(n39599), .Z(n39601) );
  AND U40618 ( .A(n39602), .B(n39601), .Z(n39650) );
  XOR U40619 ( .A(n39651), .B(n39650), .Z(n39652) );
  NANDN U40620 ( .A(n39604), .B(n39603), .Z(n39608) );
  NANDN U40621 ( .A(n39606), .B(n39605), .Z(n39607) );
  NAND U40622 ( .A(n39608), .B(n39607), .Z(n39653) );
  XOR U40623 ( .A(n39652), .B(n39653), .Z(n39620) );
  OR U40624 ( .A(n39610), .B(n39609), .Z(n39614) );
  NANDN U40625 ( .A(n39612), .B(n39611), .Z(n39613) );
  NAND U40626 ( .A(n39614), .B(n39613), .Z(n39621) );
  XNOR U40627 ( .A(n39620), .B(n39621), .Z(n39622) );
  XNOR U40628 ( .A(n39623), .B(n39622), .Z(n39656) );
  XNOR U40629 ( .A(n39656), .B(sreg[1980]), .Z(n39658) );
  NAND U40630 ( .A(n39615), .B(sreg[1979]), .Z(n39619) );
  OR U40631 ( .A(n39617), .B(n39616), .Z(n39618) );
  AND U40632 ( .A(n39619), .B(n39618), .Z(n39657) );
  XOR U40633 ( .A(n39658), .B(n39657), .Z(c[1980]) );
  NANDN U40634 ( .A(n39621), .B(n39620), .Z(n39625) );
  NAND U40635 ( .A(n39623), .B(n39622), .Z(n39624) );
  NAND U40636 ( .A(n39625), .B(n39624), .Z(n39664) );
  NAND U40637 ( .A(b[0]), .B(a[965]), .Z(n39626) );
  XNOR U40638 ( .A(b[1]), .B(n39626), .Z(n39628) );
  NAND U40639 ( .A(n152), .B(a[964]), .Z(n39627) );
  AND U40640 ( .A(n39628), .B(n39627), .Z(n39681) );
  XOR U40641 ( .A(a[961]), .B(n42197), .Z(n39670) );
  NANDN U40642 ( .A(n39670), .B(n42173), .Z(n39631) );
  NANDN U40643 ( .A(n39629), .B(n42172), .Z(n39630) );
  NAND U40644 ( .A(n39631), .B(n39630), .Z(n39679) );
  NAND U40645 ( .A(b[7]), .B(a[957]), .Z(n39680) );
  XNOR U40646 ( .A(n39679), .B(n39680), .Z(n39682) );
  XOR U40647 ( .A(n39681), .B(n39682), .Z(n39688) );
  NANDN U40648 ( .A(n39632), .B(n42093), .Z(n39634) );
  XOR U40649 ( .A(n42134), .B(a[963]), .Z(n39673) );
  NANDN U40650 ( .A(n39673), .B(n42095), .Z(n39633) );
  NAND U40651 ( .A(n39634), .B(n39633), .Z(n39686) );
  NANDN U40652 ( .A(n39635), .B(n42231), .Z(n39637) );
  XOR U40653 ( .A(n242), .B(a[959]), .Z(n39676) );
  NANDN U40654 ( .A(n39676), .B(n42234), .Z(n39636) );
  AND U40655 ( .A(n39637), .B(n39636), .Z(n39685) );
  XNOR U40656 ( .A(n39686), .B(n39685), .Z(n39687) );
  XNOR U40657 ( .A(n39688), .B(n39687), .Z(n39692) );
  NANDN U40658 ( .A(n39639), .B(n39638), .Z(n39643) );
  NAND U40659 ( .A(n39641), .B(n39640), .Z(n39642) );
  AND U40660 ( .A(n39643), .B(n39642), .Z(n39691) );
  XOR U40661 ( .A(n39692), .B(n39691), .Z(n39693) );
  NANDN U40662 ( .A(n39645), .B(n39644), .Z(n39649) );
  NANDN U40663 ( .A(n39647), .B(n39646), .Z(n39648) );
  NAND U40664 ( .A(n39649), .B(n39648), .Z(n39694) );
  XOR U40665 ( .A(n39693), .B(n39694), .Z(n39661) );
  OR U40666 ( .A(n39651), .B(n39650), .Z(n39655) );
  NANDN U40667 ( .A(n39653), .B(n39652), .Z(n39654) );
  NAND U40668 ( .A(n39655), .B(n39654), .Z(n39662) );
  XNOR U40669 ( .A(n39661), .B(n39662), .Z(n39663) );
  XNOR U40670 ( .A(n39664), .B(n39663), .Z(n39697) );
  XNOR U40671 ( .A(n39697), .B(sreg[1981]), .Z(n39699) );
  NAND U40672 ( .A(n39656), .B(sreg[1980]), .Z(n39660) );
  OR U40673 ( .A(n39658), .B(n39657), .Z(n39659) );
  AND U40674 ( .A(n39660), .B(n39659), .Z(n39698) );
  XOR U40675 ( .A(n39699), .B(n39698), .Z(c[1981]) );
  NANDN U40676 ( .A(n39662), .B(n39661), .Z(n39666) );
  NAND U40677 ( .A(n39664), .B(n39663), .Z(n39665) );
  NAND U40678 ( .A(n39666), .B(n39665), .Z(n39705) );
  NAND U40679 ( .A(b[0]), .B(a[966]), .Z(n39667) );
  XNOR U40680 ( .A(b[1]), .B(n39667), .Z(n39669) );
  NAND U40681 ( .A(n153), .B(a[965]), .Z(n39668) );
  AND U40682 ( .A(n39669), .B(n39668), .Z(n39722) );
  XOR U40683 ( .A(a[962]), .B(n42197), .Z(n39711) );
  NANDN U40684 ( .A(n39711), .B(n42173), .Z(n39672) );
  NANDN U40685 ( .A(n39670), .B(n42172), .Z(n39671) );
  NAND U40686 ( .A(n39672), .B(n39671), .Z(n39720) );
  NAND U40687 ( .A(b[7]), .B(a[958]), .Z(n39721) );
  XNOR U40688 ( .A(n39720), .B(n39721), .Z(n39723) );
  XOR U40689 ( .A(n39722), .B(n39723), .Z(n39729) );
  NANDN U40690 ( .A(n39673), .B(n42093), .Z(n39675) );
  XOR U40691 ( .A(n42134), .B(a[964]), .Z(n39714) );
  NANDN U40692 ( .A(n39714), .B(n42095), .Z(n39674) );
  NAND U40693 ( .A(n39675), .B(n39674), .Z(n39727) );
  NANDN U40694 ( .A(n39676), .B(n42231), .Z(n39678) );
  XOR U40695 ( .A(n242), .B(a[960]), .Z(n39717) );
  NANDN U40696 ( .A(n39717), .B(n42234), .Z(n39677) );
  AND U40697 ( .A(n39678), .B(n39677), .Z(n39726) );
  XNOR U40698 ( .A(n39727), .B(n39726), .Z(n39728) );
  XNOR U40699 ( .A(n39729), .B(n39728), .Z(n39733) );
  NANDN U40700 ( .A(n39680), .B(n39679), .Z(n39684) );
  NAND U40701 ( .A(n39682), .B(n39681), .Z(n39683) );
  AND U40702 ( .A(n39684), .B(n39683), .Z(n39732) );
  XOR U40703 ( .A(n39733), .B(n39732), .Z(n39734) );
  NANDN U40704 ( .A(n39686), .B(n39685), .Z(n39690) );
  NANDN U40705 ( .A(n39688), .B(n39687), .Z(n39689) );
  NAND U40706 ( .A(n39690), .B(n39689), .Z(n39735) );
  XOR U40707 ( .A(n39734), .B(n39735), .Z(n39702) );
  OR U40708 ( .A(n39692), .B(n39691), .Z(n39696) );
  NANDN U40709 ( .A(n39694), .B(n39693), .Z(n39695) );
  NAND U40710 ( .A(n39696), .B(n39695), .Z(n39703) );
  XNOR U40711 ( .A(n39702), .B(n39703), .Z(n39704) );
  XNOR U40712 ( .A(n39705), .B(n39704), .Z(n39738) );
  XNOR U40713 ( .A(n39738), .B(sreg[1982]), .Z(n39740) );
  NAND U40714 ( .A(n39697), .B(sreg[1981]), .Z(n39701) );
  OR U40715 ( .A(n39699), .B(n39698), .Z(n39700) );
  AND U40716 ( .A(n39701), .B(n39700), .Z(n39739) );
  XOR U40717 ( .A(n39740), .B(n39739), .Z(c[1982]) );
  NANDN U40718 ( .A(n39703), .B(n39702), .Z(n39707) );
  NAND U40719 ( .A(n39705), .B(n39704), .Z(n39706) );
  NAND U40720 ( .A(n39707), .B(n39706), .Z(n39746) );
  NAND U40721 ( .A(b[0]), .B(a[967]), .Z(n39708) );
  XNOR U40722 ( .A(b[1]), .B(n39708), .Z(n39710) );
  NAND U40723 ( .A(n153), .B(a[966]), .Z(n39709) );
  AND U40724 ( .A(n39710), .B(n39709), .Z(n39763) );
  XOR U40725 ( .A(a[963]), .B(n42197), .Z(n39752) );
  NANDN U40726 ( .A(n39752), .B(n42173), .Z(n39713) );
  NANDN U40727 ( .A(n39711), .B(n42172), .Z(n39712) );
  NAND U40728 ( .A(n39713), .B(n39712), .Z(n39761) );
  NAND U40729 ( .A(b[7]), .B(a[959]), .Z(n39762) );
  XNOR U40730 ( .A(n39761), .B(n39762), .Z(n39764) );
  XOR U40731 ( .A(n39763), .B(n39764), .Z(n39770) );
  NANDN U40732 ( .A(n39714), .B(n42093), .Z(n39716) );
  XOR U40733 ( .A(n42134), .B(a[965]), .Z(n39755) );
  NANDN U40734 ( .A(n39755), .B(n42095), .Z(n39715) );
  NAND U40735 ( .A(n39716), .B(n39715), .Z(n39768) );
  NANDN U40736 ( .A(n39717), .B(n42231), .Z(n39719) );
  XOR U40737 ( .A(n242), .B(a[961]), .Z(n39758) );
  NANDN U40738 ( .A(n39758), .B(n42234), .Z(n39718) );
  AND U40739 ( .A(n39719), .B(n39718), .Z(n39767) );
  XNOR U40740 ( .A(n39768), .B(n39767), .Z(n39769) );
  XNOR U40741 ( .A(n39770), .B(n39769), .Z(n39774) );
  NANDN U40742 ( .A(n39721), .B(n39720), .Z(n39725) );
  NAND U40743 ( .A(n39723), .B(n39722), .Z(n39724) );
  AND U40744 ( .A(n39725), .B(n39724), .Z(n39773) );
  XOR U40745 ( .A(n39774), .B(n39773), .Z(n39775) );
  NANDN U40746 ( .A(n39727), .B(n39726), .Z(n39731) );
  NANDN U40747 ( .A(n39729), .B(n39728), .Z(n39730) );
  NAND U40748 ( .A(n39731), .B(n39730), .Z(n39776) );
  XOR U40749 ( .A(n39775), .B(n39776), .Z(n39743) );
  OR U40750 ( .A(n39733), .B(n39732), .Z(n39737) );
  NANDN U40751 ( .A(n39735), .B(n39734), .Z(n39736) );
  NAND U40752 ( .A(n39737), .B(n39736), .Z(n39744) );
  XNOR U40753 ( .A(n39743), .B(n39744), .Z(n39745) );
  XNOR U40754 ( .A(n39746), .B(n39745), .Z(n39779) );
  XNOR U40755 ( .A(n39779), .B(sreg[1983]), .Z(n39781) );
  NAND U40756 ( .A(n39738), .B(sreg[1982]), .Z(n39742) );
  OR U40757 ( .A(n39740), .B(n39739), .Z(n39741) );
  AND U40758 ( .A(n39742), .B(n39741), .Z(n39780) );
  XOR U40759 ( .A(n39781), .B(n39780), .Z(c[1983]) );
  NANDN U40760 ( .A(n39744), .B(n39743), .Z(n39748) );
  NAND U40761 ( .A(n39746), .B(n39745), .Z(n39747) );
  NAND U40762 ( .A(n39748), .B(n39747), .Z(n39787) );
  NAND U40763 ( .A(b[0]), .B(a[968]), .Z(n39749) );
  XNOR U40764 ( .A(b[1]), .B(n39749), .Z(n39751) );
  NAND U40765 ( .A(n153), .B(a[967]), .Z(n39750) );
  AND U40766 ( .A(n39751), .B(n39750), .Z(n39804) );
  XOR U40767 ( .A(a[964]), .B(n42197), .Z(n39793) );
  NANDN U40768 ( .A(n39793), .B(n42173), .Z(n39754) );
  NANDN U40769 ( .A(n39752), .B(n42172), .Z(n39753) );
  NAND U40770 ( .A(n39754), .B(n39753), .Z(n39802) );
  NAND U40771 ( .A(b[7]), .B(a[960]), .Z(n39803) );
  XNOR U40772 ( .A(n39802), .B(n39803), .Z(n39805) );
  XOR U40773 ( .A(n39804), .B(n39805), .Z(n39811) );
  NANDN U40774 ( .A(n39755), .B(n42093), .Z(n39757) );
  XOR U40775 ( .A(n42134), .B(a[966]), .Z(n39796) );
  NANDN U40776 ( .A(n39796), .B(n42095), .Z(n39756) );
  NAND U40777 ( .A(n39757), .B(n39756), .Z(n39809) );
  NANDN U40778 ( .A(n39758), .B(n42231), .Z(n39760) );
  XOR U40779 ( .A(n242), .B(a[962]), .Z(n39799) );
  NANDN U40780 ( .A(n39799), .B(n42234), .Z(n39759) );
  AND U40781 ( .A(n39760), .B(n39759), .Z(n39808) );
  XNOR U40782 ( .A(n39809), .B(n39808), .Z(n39810) );
  XNOR U40783 ( .A(n39811), .B(n39810), .Z(n39815) );
  NANDN U40784 ( .A(n39762), .B(n39761), .Z(n39766) );
  NAND U40785 ( .A(n39764), .B(n39763), .Z(n39765) );
  AND U40786 ( .A(n39766), .B(n39765), .Z(n39814) );
  XOR U40787 ( .A(n39815), .B(n39814), .Z(n39816) );
  NANDN U40788 ( .A(n39768), .B(n39767), .Z(n39772) );
  NANDN U40789 ( .A(n39770), .B(n39769), .Z(n39771) );
  NAND U40790 ( .A(n39772), .B(n39771), .Z(n39817) );
  XOR U40791 ( .A(n39816), .B(n39817), .Z(n39784) );
  OR U40792 ( .A(n39774), .B(n39773), .Z(n39778) );
  NANDN U40793 ( .A(n39776), .B(n39775), .Z(n39777) );
  NAND U40794 ( .A(n39778), .B(n39777), .Z(n39785) );
  XNOR U40795 ( .A(n39784), .B(n39785), .Z(n39786) );
  XNOR U40796 ( .A(n39787), .B(n39786), .Z(n39820) );
  XNOR U40797 ( .A(n39820), .B(sreg[1984]), .Z(n39822) );
  NAND U40798 ( .A(n39779), .B(sreg[1983]), .Z(n39783) );
  OR U40799 ( .A(n39781), .B(n39780), .Z(n39782) );
  AND U40800 ( .A(n39783), .B(n39782), .Z(n39821) );
  XOR U40801 ( .A(n39822), .B(n39821), .Z(c[1984]) );
  NANDN U40802 ( .A(n39785), .B(n39784), .Z(n39789) );
  NAND U40803 ( .A(n39787), .B(n39786), .Z(n39788) );
  NAND U40804 ( .A(n39789), .B(n39788), .Z(n39828) );
  NAND U40805 ( .A(b[0]), .B(a[969]), .Z(n39790) );
  XNOR U40806 ( .A(b[1]), .B(n39790), .Z(n39792) );
  NAND U40807 ( .A(n153), .B(a[968]), .Z(n39791) );
  AND U40808 ( .A(n39792), .B(n39791), .Z(n39845) );
  XOR U40809 ( .A(a[965]), .B(n42197), .Z(n39834) );
  NANDN U40810 ( .A(n39834), .B(n42173), .Z(n39795) );
  NANDN U40811 ( .A(n39793), .B(n42172), .Z(n39794) );
  NAND U40812 ( .A(n39795), .B(n39794), .Z(n39843) );
  NAND U40813 ( .A(b[7]), .B(a[961]), .Z(n39844) );
  XNOR U40814 ( .A(n39843), .B(n39844), .Z(n39846) );
  XOR U40815 ( .A(n39845), .B(n39846), .Z(n39852) );
  NANDN U40816 ( .A(n39796), .B(n42093), .Z(n39798) );
  XOR U40817 ( .A(n42134), .B(a[967]), .Z(n39837) );
  NANDN U40818 ( .A(n39837), .B(n42095), .Z(n39797) );
  NAND U40819 ( .A(n39798), .B(n39797), .Z(n39850) );
  NANDN U40820 ( .A(n39799), .B(n42231), .Z(n39801) );
  XOR U40821 ( .A(n242), .B(a[963]), .Z(n39840) );
  NANDN U40822 ( .A(n39840), .B(n42234), .Z(n39800) );
  AND U40823 ( .A(n39801), .B(n39800), .Z(n39849) );
  XNOR U40824 ( .A(n39850), .B(n39849), .Z(n39851) );
  XNOR U40825 ( .A(n39852), .B(n39851), .Z(n39856) );
  NANDN U40826 ( .A(n39803), .B(n39802), .Z(n39807) );
  NAND U40827 ( .A(n39805), .B(n39804), .Z(n39806) );
  AND U40828 ( .A(n39807), .B(n39806), .Z(n39855) );
  XOR U40829 ( .A(n39856), .B(n39855), .Z(n39857) );
  NANDN U40830 ( .A(n39809), .B(n39808), .Z(n39813) );
  NANDN U40831 ( .A(n39811), .B(n39810), .Z(n39812) );
  NAND U40832 ( .A(n39813), .B(n39812), .Z(n39858) );
  XOR U40833 ( .A(n39857), .B(n39858), .Z(n39825) );
  OR U40834 ( .A(n39815), .B(n39814), .Z(n39819) );
  NANDN U40835 ( .A(n39817), .B(n39816), .Z(n39818) );
  NAND U40836 ( .A(n39819), .B(n39818), .Z(n39826) );
  XNOR U40837 ( .A(n39825), .B(n39826), .Z(n39827) );
  XNOR U40838 ( .A(n39828), .B(n39827), .Z(n39861) );
  XNOR U40839 ( .A(n39861), .B(sreg[1985]), .Z(n39863) );
  NAND U40840 ( .A(n39820), .B(sreg[1984]), .Z(n39824) );
  OR U40841 ( .A(n39822), .B(n39821), .Z(n39823) );
  AND U40842 ( .A(n39824), .B(n39823), .Z(n39862) );
  XOR U40843 ( .A(n39863), .B(n39862), .Z(c[1985]) );
  NANDN U40844 ( .A(n39826), .B(n39825), .Z(n39830) );
  NAND U40845 ( .A(n39828), .B(n39827), .Z(n39829) );
  NAND U40846 ( .A(n39830), .B(n39829), .Z(n39869) );
  NAND U40847 ( .A(b[0]), .B(a[970]), .Z(n39831) );
  XNOR U40848 ( .A(b[1]), .B(n39831), .Z(n39833) );
  NAND U40849 ( .A(n153), .B(a[969]), .Z(n39832) );
  AND U40850 ( .A(n39833), .B(n39832), .Z(n39886) );
  XOR U40851 ( .A(a[966]), .B(n42197), .Z(n39875) );
  NANDN U40852 ( .A(n39875), .B(n42173), .Z(n39836) );
  NANDN U40853 ( .A(n39834), .B(n42172), .Z(n39835) );
  NAND U40854 ( .A(n39836), .B(n39835), .Z(n39884) );
  NAND U40855 ( .A(b[7]), .B(a[962]), .Z(n39885) );
  XNOR U40856 ( .A(n39884), .B(n39885), .Z(n39887) );
  XOR U40857 ( .A(n39886), .B(n39887), .Z(n39893) );
  NANDN U40858 ( .A(n39837), .B(n42093), .Z(n39839) );
  XOR U40859 ( .A(n42134), .B(a[968]), .Z(n39878) );
  NANDN U40860 ( .A(n39878), .B(n42095), .Z(n39838) );
  NAND U40861 ( .A(n39839), .B(n39838), .Z(n39891) );
  NANDN U40862 ( .A(n39840), .B(n42231), .Z(n39842) );
  XOR U40863 ( .A(n242), .B(a[964]), .Z(n39881) );
  NANDN U40864 ( .A(n39881), .B(n42234), .Z(n39841) );
  AND U40865 ( .A(n39842), .B(n39841), .Z(n39890) );
  XNOR U40866 ( .A(n39891), .B(n39890), .Z(n39892) );
  XNOR U40867 ( .A(n39893), .B(n39892), .Z(n39897) );
  NANDN U40868 ( .A(n39844), .B(n39843), .Z(n39848) );
  NAND U40869 ( .A(n39846), .B(n39845), .Z(n39847) );
  AND U40870 ( .A(n39848), .B(n39847), .Z(n39896) );
  XOR U40871 ( .A(n39897), .B(n39896), .Z(n39898) );
  NANDN U40872 ( .A(n39850), .B(n39849), .Z(n39854) );
  NANDN U40873 ( .A(n39852), .B(n39851), .Z(n39853) );
  NAND U40874 ( .A(n39854), .B(n39853), .Z(n39899) );
  XOR U40875 ( .A(n39898), .B(n39899), .Z(n39866) );
  OR U40876 ( .A(n39856), .B(n39855), .Z(n39860) );
  NANDN U40877 ( .A(n39858), .B(n39857), .Z(n39859) );
  NAND U40878 ( .A(n39860), .B(n39859), .Z(n39867) );
  XNOR U40879 ( .A(n39866), .B(n39867), .Z(n39868) );
  XNOR U40880 ( .A(n39869), .B(n39868), .Z(n39902) );
  XNOR U40881 ( .A(n39902), .B(sreg[1986]), .Z(n39904) );
  NAND U40882 ( .A(n39861), .B(sreg[1985]), .Z(n39865) );
  OR U40883 ( .A(n39863), .B(n39862), .Z(n39864) );
  AND U40884 ( .A(n39865), .B(n39864), .Z(n39903) );
  XOR U40885 ( .A(n39904), .B(n39903), .Z(c[1986]) );
  NANDN U40886 ( .A(n39867), .B(n39866), .Z(n39871) );
  NAND U40887 ( .A(n39869), .B(n39868), .Z(n39870) );
  NAND U40888 ( .A(n39871), .B(n39870), .Z(n39910) );
  NAND U40889 ( .A(b[0]), .B(a[971]), .Z(n39872) );
  XNOR U40890 ( .A(b[1]), .B(n39872), .Z(n39874) );
  NAND U40891 ( .A(n153), .B(a[970]), .Z(n39873) );
  AND U40892 ( .A(n39874), .B(n39873), .Z(n39927) );
  XOR U40893 ( .A(a[967]), .B(n42197), .Z(n39916) );
  NANDN U40894 ( .A(n39916), .B(n42173), .Z(n39877) );
  NANDN U40895 ( .A(n39875), .B(n42172), .Z(n39876) );
  NAND U40896 ( .A(n39877), .B(n39876), .Z(n39925) );
  NAND U40897 ( .A(b[7]), .B(a[963]), .Z(n39926) );
  XNOR U40898 ( .A(n39925), .B(n39926), .Z(n39928) );
  XOR U40899 ( .A(n39927), .B(n39928), .Z(n39934) );
  NANDN U40900 ( .A(n39878), .B(n42093), .Z(n39880) );
  XOR U40901 ( .A(n42134), .B(a[969]), .Z(n39919) );
  NANDN U40902 ( .A(n39919), .B(n42095), .Z(n39879) );
  NAND U40903 ( .A(n39880), .B(n39879), .Z(n39932) );
  NANDN U40904 ( .A(n39881), .B(n42231), .Z(n39883) );
  XOR U40905 ( .A(n242), .B(a[965]), .Z(n39922) );
  NANDN U40906 ( .A(n39922), .B(n42234), .Z(n39882) );
  AND U40907 ( .A(n39883), .B(n39882), .Z(n39931) );
  XNOR U40908 ( .A(n39932), .B(n39931), .Z(n39933) );
  XNOR U40909 ( .A(n39934), .B(n39933), .Z(n39938) );
  NANDN U40910 ( .A(n39885), .B(n39884), .Z(n39889) );
  NAND U40911 ( .A(n39887), .B(n39886), .Z(n39888) );
  AND U40912 ( .A(n39889), .B(n39888), .Z(n39937) );
  XOR U40913 ( .A(n39938), .B(n39937), .Z(n39939) );
  NANDN U40914 ( .A(n39891), .B(n39890), .Z(n39895) );
  NANDN U40915 ( .A(n39893), .B(n39892), .Z(n39894) );
  NAND U40916 ( .A(n39895), .B(n39894), .Z(n39940) );
  XOR U40917 ( .A(n39939), .B(n39940), .Z(n39907) );
  OR U40918 ( .A(n39897), .B(n39896), .Z(n39901) );
  NANDN U40919 ( .A(n39899), .B(n39898), .Z(n39900) );
  NAND U40920 ( .A(n39901), .B(n39900), .Z(n39908) );
  XNOR U40921 ( .A(n39907), .B(n39908), .Z(n39909) );
  XNOR U40922 ( .A(n39910), .B(n39909), .Z(n39943) );
  XNOR U40923 ( .A(n39943), .B(sreg[1987]), .Z(n39945) );
  NAND U40924 ( .A(n39902), .B(sreg[1986]), .Z(n39906) );
  OR U40925 ( .A(n39904), .B(n39903), .Z(n39905) );
  AND U40926 ( .A(n39906), .B(n39905), .Z(n39944) );
  XOR U40927 ( .A(n39945), .B(n39944), .Z(c[1987]) );
  NANDN U40928 ( .A(n39908), .B(n39907), .Z(n39912) );
  NAND U40929 ( .A(n39910), .B(n39909), .Z(n39911) );
  NAND U40930 ( .A(n39912), .B(n39911), .Z(n39951) );
  NAND U40931 ( .A(b[0]), .B(a[972]), .Z(n39913) );
  XNOR U40932 ( .A(b[1]), .B(n39913), .Z(n39915) );
  NAND U40933 ( .A(n153), .B(a[971]), .Z(n39914) );
  AND U40934 ( .A(n39915), .B(n39914), .Z(n39968) );
  XOR U40935 ( .A(a[968]), .B(n42197), .Z(n39957) );
  NANDN U40936 ( .A(n39957), .B(n42173), .Z(n39918) );
  NANDN U40937 ( .A(n39916), .B(n42172), .Z(n39917) );
  NAND U40938 ( .A(n39918), .B(n39917), .Z(n39966) );
  NAND U40939 ( .A(b[7]), .B(a[964]), .Z(n39967) );
  XNOR U40940 ( .A(n39966), .B(n39967), .Z(n39969) );
  XOR U40941 ( .A(n39968), .B(n39969), .Z(n39975) );
  NANDN U40942 ( .A(n39919), .B(n42093), .Z(n39921) );
  XOR U40943 ( .A(n42134), .B(a[970]), .Z(n39960) );
  NANDN U40944 ( .A(n39960), .B(n42095), .Z(n39920) );
  NAND U40945 ( .A(n39921), .B(n39920), .Z(n39973) );
  NANDN U40946 ( .A(n39922), .B(n42231), .Z(n39924) );
  XOR U40947 ( .A(n242), .B(a[966]), .Z(n39963) );
  NANDN U40948 ( .A(n39963), .B(n42234), .Z(n39923) );
  AND U40949 ( .A(n39924), .B(n39923), .Z(n39972) );
  XNOR U40950 ( .A(n39973), .B(n39972), .Z(n39974) );
  XNOR U40951 ( .A(n39975), .B(n39974), .Z(n39979) );
  NANDN U40952 ( .A(n39926), .B(n39925), .Z(n39930) );
  NAND U40953 ( .A(n39928), .B(n39927), .Z(n39929) );
  AND U40954 ( .A(n39930), .B(n39929), .Z(n39978) );
  XOR U40955 ( .A(n39979), .B(n39978), .Z(n39980) );
  NANDN U40956 ( .A(n39932), .B(n39931), .Z(n39936) );
  NANDN U40957 ( .A(n39934), .B(n39933), .Z(n39935) );
  NAND U40958 ( .A(n39936), .B(n39935), .Z(n39981) );
  XOR U40959 ( .A(n39980), .B(n39981), .Z(n39948) );
  OR U40960 ( .A(n39938), .B(n39937), .Z(n39942) );
  NANDN U40961 ( .A(n39940), .B(n39939), .Z(n39941) );
  NAND U40962 ( .A(n39942), .B(n39941), .Z(n39949) );
  XNOR U40963 ( .A(n39948), .B(n39949), .Z(n39950) );
  XNOR U40964 ( .A(n39951), .B(n39950), .Z(n39984) );
  XNOR U40965 ( .A(n39984), .B(sreg[1988]), .Z(n39986) );
  NAND U40966 ( .A(n39943), .B(sreg[1987]), .Z(n39947) );
  OR U40967 ( .A(n39945), .B(n39944), .Z(n39946) );
  AND U40968 ( .A(n39947), .B(n39946), .Z(n39985) );
  XOR U40969 ( .A(n39986), .B(n39985), .Z(c[1988]) );
  NANDN U40970 ( .A(n39949), .B(n39948), .Z(n39953) );
  NAND U40971 ( .A(n39951), .B(n39950), .Z(n39952) );
  NAND U40972 ( .A(n39953), .B(n39952), .Z(n39992) );
  NAND U40973 ( .A(b[0]), .B(a[973]), .Z(n39954) );
  XNOR U40974 ( .A(b[1]), .B(n39954), .Z(n39956) );
  NAND U40975 ( .A(n154), .B(a[972]), .Z(n39955) );
  AND U40976 ( .A(n39956), .B(n39955), .Z(n40009) );
  XOR U40977 ( .A(a[969]), .B(n42197), .Z(n39998) );
  NANDN U40978 ( .A(n39998), .B(n42173), .Z(n39959) );
  NANDN U40979 ( .A(n39957), .B(n42172), .Z(n39958) );
  NAND U40980 ( .A(n39959), .B(n39958), .Z(n40007) );
  NAND U40981 ( .A(b[7]), .B(a[965]), .Z(n40008) );
  XNOR U40982 ( .A(n40007), .B(n40008), .Z(n40010) );
  XOR U40983 ( .A(n40009), .B(n40010), .Z(n40016) );
  NANDN U40984 ( .A(n39960), .B(n42093), .Z(n39962) );
  XOR U40985 ( .A(n42134), .B(a[971]), .Z(n40001) );
  NANDN U40986 ( .A(n40001), .B(n42095), .Z(n39961) );
  NAND U40987 ( .A(n39962), .B(n39961), .Z(n40014) );
  NANDN U40988 ( .A(n39963), .B(n42231), .Z(n39965) );
  XOR U40989 ( .A(n242), .B(a[967]), .Z(n40004) );
  NANDN U40990 ( .A(n40004), .B(n42234), .Z(n39964) );
  AND U40991 ( .A(n39965), .B(n39964), .Z(n40013) );
  XNOR U40992 ( .A(n40014), .B(n40013), .Z(n40015) );
  XNOR U40993 ( .A(n40016), .B(n40015), .Z(n40020) );
  NANDN U40994 ( .A(n39967), .B(n39966), .Z(n39971) );
  NAND U40995 ( .A(n39969), .B(n39968), .Z(n39970) );
  AND U40996 ( .A(n39971), .B(n39970), .Z(n40019) );
  XOR U40997 ( .A(n40020), .B(n40019), .Z(n40021) );
  NANDN U40998 ( .A(n39973), .B(n39972), .Z(n39977) );
  NANDN U40999 ( .A(n39975), .B(n39974), .Z(n39976) );
  NAND U41000 ( .A(n39977), .B(n39976), .Z(n40022) );
  XOR U41001 ( .A(n40021), .B(n40022), .Z(n39989) );
  OR U41002 ( .A(n39979), .B(n39978), .Z(n39983) );
  NANDN U41003 ( .A(n39981), .B(n39980), .Z(n39982) );
  NAND U41004 ( .A(n39983), .B(n39982), .Z(n39990) );
  XNOR U41005 ( .A(n39989), .B(n39990), .Z(n39991) );
  XNOR U41006 ( .A(n39992), .B(n39991), .Z(n40025) );
  XNOR U41007 ( .A(n40025), .B(sreg[1989]), .Z(n40027) );
  NAND U41008 ( .A(n39984), .B(sreg[1988]), .Z(n39988) );
  OR U41009 ( .A(n39986), .B(n39985), .Z(n39987) );
  AND U41010 ( .A(n39988), .B(n39987), .Z(n40026) );
  XOR U41011 ( .A(n40027), .B(n40026), .Z(c[1989]) );
  NANDN U41012 ( .A(n39990), .B(n39989), .Z(n39994) );
  NAND U41013 ( .A(n39992), .B(n39991), .Z(n39993) );
  NAND U41014 ( .A(n39994), .B(n39993), .Z(n40033) );
  NAND U41015 ( .A(b[0]), .B(a[974]), .Z(n39995) );
  XNOR U41016 ( .A(b[1]), .B(n39995), .Z(n39997) );
  NAND U41017 ( .A(n154), .B(a[973]), .Z(n39996) );
  AND U41018 ( .A(n39997), .B(n39996), .Z(n40050) );
  XOR U41019 ( .A(a[970]), .B(n42197), .Z(n40039) );
  NANDN U41020 ( .A(n40039), .B(n42173), .Z(n40000) );
  NANDN U41021 ( .A(n39998), .B(n42172), .Z(n39999) );
  NAND U41022 ( .A(n40000), .B(n39999), .Z(n40048) );
  NAND U41023 ( .A(b[7]), .B(a[966]), .Z(n40049) );
  XNOR U41024 ( .A(n40048), .B(n40049), .Z(n40051) );
  XOR U41025 ( .A(n40050), .B(n40051), .Z(n40057) );
  NANDN U41026 ( .A(n40001), .B(n42093), .Z(n40003) );
  XOR U41027 ( .A(n42134), .B(a[972]), .Z(n40042) );
  NANDN U41028 ( .A(n40042), .B(n42095), .Z(n40002) );
  NAND U41029 ( .A(n40003), .B(n40002), .Z(n40055) );
  NANDN U41030 ( .A(n40004), .B(n42231), .Z(n40006) );
  XOR U41031 ( .A(n242), .B(a[968]), .Z(n40045) );
  NANDN U41032 ( .A(n40045), .B(n42234), .Z(n40005) );
  AND U41033 ( .A(n40006), .B(n40005), .Z(n40054) );
  XNOR U41034 ( .A(n40055), .B(n40054), .Z(n40056) );
  XNOR U41035 ( .A(n40057), .B(n40056), .Z(n40061) );
  NANDN U41036 ( .A(n40008), .B(n40007), .Z(n40012) );
  NAND U41037 ( .A(n40010), .B(n40009), .Z(n40011) );
  AND U41038 ( .A(n40012), .B(n40011), .Z(n40060) );
  XOR U41039 ( .A(n40061), .B(n40060), .Z(n40062) );
  NANDN U41040 ( .A(n40014), .B(n40013), .Z(n40018) );
  NANDN U41041 ( .A(n40016), .B(n40015), .Z(n40017) );
  NAND U41042 ( .A(n40018), .B(n40017), .Z(n40063) );
  XOR U41043 ( .A(n40062), .B(n40063), .Z(n40030) );
  OR U41044 ( .A(n40020), .B(n40019), .Z(n40024) );
  NANDN U41045 ( .A(n40022), .B(n40021), .Z(n40023) );
  NAND U41046 ( .A(n40024), .B(n40023), .Z(n40031) );
  XNOR U41047 ( .A(n40030), .B(n40031), .Z(n40032) );
  XNOR U41048 ( .A(n40033), .B(n40032), .Z(n40066) );
  XNOR U41049 ( .A(n40066), .B(sreg[1990]), .Z(n40068) );
  NAND U41050 ( .A(n40025), .B(sreg[1989]), .Z(n40029) );
  OR U41051 ( .A(n40027), .B(n40026), .Z(n40028) );
  AND U41052 ( .A(n40029), .B(n40028), .Z(n40067) );
  XOR U41053 ( .A(n40068), .B(n40067), .Z(c[1990]) );
  NANDN U41054 ( .A(n40031), .B(n40030), .Z(n40035) );
  NAND U41055 ( .A(n40033), .B(n40032), .Z(n40034) );
  NAND U41056 ( .A(n40035), .B(n40034), .Z(n40074) );
  NAND U41057 ( .A(b[0]), .B(a[975]), .Z(n40036) );
  XNOR U41058 ( .A(b[1]), .B(n40036), .Z(n40038) );
  NAND U41059 ( .A(n154), .B(a[974]), .Z(n40037) );
  AND U41060 ( .A(n40038), .B(n40037), .Z(n40091) );
  XOR U41061 ( .A(a[971]), .B(n42197), .Z(n40080) );
  NANDN U41062 ( .A(n40080), .B(n42173), .Z(n40041) );
  NANDN U41063 ( .A(n40039), .B(n42172), .Z(n40040) );
  NAND U41064 ( .A(n40041), .B(n40040), .Z(n40089) );
  NAND U41065 ( .A(b[7]), .B(a[967]), .Z(n40090) );
  XNOR U41066 ( .A(n40089), .B(n40090), .Z(n40092) );
  XOR U41067 ( .A(n40091), .B(n40092), .Z(n40098) );
  NANDN U41068 ( .A(n40042), .B(n42093), .Z(n40044) );
  XOR U41069 ( .A(n42134), .B(a[973]), .Z(n40083) );
  NANDN U41070 ( .A(n40083), .B(n42095), .Z(n40043) );
  NAND U41071 ( .A(n40044), .B(n40043), .Z(n40096) );
  NANDN U41072 ( .A(n40045), .B(n42231), .Z(n40047) );
  XOR U41073 ( .A(n242), .B(a[969]), .Z(n40086) );
  NANDN U41074 ( .A(n40086), .B(n42234), .Z(n40046) );
  AND U41075 ( .A(n40047), .B(n40046), .Z(n40095) );
  XNOR U41076 ( .A(n40096), .B(n40095), .Z(n40097) );
  XNOR U41077 ( .A(n40098), .B(n40097), .Z(n40102) );
  NANDN U41078 ( .A(n40049), .B(n40048), .Z(n40053) );
  NAND U41079 ( .A(n40051), .B(n40050), .Z(n40052) );
  AND U41080 ( .A(n40053), .B(n40052), .Z(n40101) );
  XOR U41081 ( .A(n40102), .B(n40101), .Z(n40103) );
  NANDN U41082 ( .A(n40055), .B(n40054), .Z(n40059) );
  NANDN U41083 ( .A(n40057), .B(n40056), .Z(n40058) );
  NAND U41084 ( .A(n40059), .B(n40058), .Z(n40104) );
  XOR U41085 ( .A(n40103), .B(n40104), .Z(n40071) );
  OR U41086 ( .A(n40061), .B(n40060), .Z(n40065) );
  NANDN U41087 ( .A(n40063), .B(n40062), .Z(n40064) );
  NAND U41088 ( .A(n40065), .B(n40064), .Z(n40072) );
  XNOR U41089 ( .A(n40071), .B(n40072), .Z(n40073) );
  XNOR U41090 ( .A(n40074), .B(n40073), .Z(n40107) );
  XNOR U41091 ( .A(n40107), .B(sreg[1991]), .Z(n40109) );
  NAND U41092 ( .A(n40066), .B(sreg[1990]), .Z(n40070) );
  OR U41093 ( .A(n40068), .B(n40067), .Z(n40069) );
  AND U41094 ( .A(n40070), .B(n40069), .Z(n40108) );
  XOR U41095 ( .A(n40109), .B(n40108), .Z(c[1991]) );
  NANDN U41096 ( .A(n40072), .B(n40071), .Z(n40076) );
  NAND U41097 ( .A(n40074), .B(n40073), .Z(n40075) );
  NAND U41098 ( .A(n40076), .B(n40075), .Z(n40115) );
  NAND U41099 ( .A(b[0]), .B(a[976]), .Z(n40077) );
  XNOR U41100 ( .A(b[1]), .B(n40077), .Z(n40079) );
  NAND U41101 ( .A(n154), .B(a[975]), .Z(n40078) );
  AND U41102 ( .A(n40079), .B(n40078), .Z(n40132) );
  XOR U41103 ( .A(a[972]), .B(n42197), .Z(n40121) );
  NANDN U41104 ( .A(n40121), .B(n42173), .Z(n40082) );
  NANDN U41105 ( .A(n40080), .B(n42172), .Z(n40081) );
  NAND U41106 ( .A(n40082), .B(n40081), .Z(n40130) );
  NAND U41107 ( .A(b[7]), .B(a[968]), .Z(n40131) );
  XNOR U41108 ( .A(n40130), .B(n40131), .Z(n40133) );
  XOR U41109 ( .A(n40132), .B(n40133), .Z(n40139) );
  NANDN U41110 ( .A(n40083), .B(n42093), .Z(n40085) );
  XOR U41111 ( .A(n42134), .B(a[974]), .Z(n40124) );
  NANDN U41112 ( .A(n40124), .B(n42095), .Z(n40084) );
  NAND U41113 ( .A(n40085), .B(n40084), .Z(n40137) );
  NANDN U41114 ( .A(n40086), .B(n42231), .Z(n40088) );
  XOR U41115 ( .A(n242), .B(a[970]), .Z(n40127) );
  NANDN U41116 ( .A(n40127), .B(n42234), .Z(n40087) );
  AND U41117 ( .A(n40088), .B(n40087), .Z(n40136) );
  XNOR U41118 ( .A(n40137), .B(n40136), .Z(n40138) );
  XNOR U41119 ( .A(n40139), .B(n40138), .Z(n40143) );
  NANDN U41120 ( .A(n40090), .B(n40089), .Z(n40094) );
  NAND U41121 ( .A(n40092), .B(n40091), .Z(n40093) );
  AND U41122 ( .A(n40094), .B(n40093), .Z(n40142) );
  XOR U41123 ( .A(n40143), .B(n40142), .Z(n40144) );
  NANDN U41124 ( .A(n40096), .B(n40095), .Z(n40100) );
  NANDN U41125 ( .A(n40098), .B(n40097), .Z(n40099) );
  NAND U41126 ( .A(n40100), .B(n40099), .Z(n40145) );
  XOR U41127 ( .A(n40144), .B(n40145), .Z(n40112) );
  OR U41128 ( .A(n40102), .B(n40101), .Z(n40106) );
  NANDN U41129 ( .A(n40104), .B(n40103), .Z(n40105) );
  NAND U41130 ( .A(n40106), .B(n40105), .Z(n40113) );
  XNOR U41131 ( .A(n40112), .B(n40113), .Z(n40114) );
  XNOR U41132 ( .A(n40115), .B(n40114), .Z(n40148) );
  XNOR U41133 ( .A(n40148), .B(sreg[1992]), .Z(n40150) );
  NAND U41134 ( .A(n40107), .B(sreg[1991]), .Z(n40111) );
  OR U41135 ( .A(n40109), .B(n40108), .Z(n40110) );
  AND U41136 ( .A(n40111), .B(n40110), .Z(n40149) );
  XOR U41137 ( .A(n40150), .B(n40149), .Z(c[1992]) );
  NANDN U41138 ( .A(n40113), .B(n40112), .Z(n40117) );
  NAND U41139 ( .A(n40115), .B(n40114), .Z(n40116) );
  NAND U41140 ( .A(n40117), .B(n40116), .Z(n40156) );
  NAND U41141 ( .A(b[0]), .B(a[977]), .Z(n40118) );
  XNOR U41142 ( .A(b[1]), .B(n40118), .Z(n40120) );
  NAND U41143 ( .A(n154), .B(a[976]), .Z(n40119) );
  AND U41144 ( .A(n40120), .B(n40119), .Z(n40173) );
  XOR U41145 ( .A(a[973]), .B(n42197), .Z(n40162) );
  NANDN U41146 ( .A(n40162), .B(n42173), .Z(n40123) );
  NANDN U41147 ( .A(n40121), .B(n42172), .Z(n40122) );
  NAND U41148 ( .A(n40123), .B(n40122), .Z(n40171) );
  NAND U41149 ( .A(b[7]), .B(a[969]), .Z(n40172) );
  XNOR U41150 ( .A(n40171), .B(n40172), .Z(n40174) );
  XOR U41151 ( .A(n40173), .B(n40174), .Z(n40180) );
  NANDN U41152 ( .A(n40124), .B(n42093), .Z(n40126) );
  XOR U41153 ( .A(n42134), .B(a[975]), .Z(n40165) );
  NANDN U41154 ( .A(n40165), .B(n42095), .Z(n40125) );
  NAND U41155 ( .A(n40126), .B(n40125), .Z(n40178) );
  NANDN U41156 ( .A(n40127), .B(n42231), .Z(n40129) );
  XOR U41157 ( .A(n243), .B(a[971]), .Z(n40168) );
  NANDN U41158 ( .A(n40168), .B(n42234), .Z(n40128) );
  AND U41159 ( .A(n40129), .B(n40128), .Z(n40177) );
  XNOR U41160 ( .A(n40178), .B(n40177), .Z(n40179) );
  XNOR U41161 ( .A(n40180), .B(n40179), .Z(n40184) );
  NANDN U41162 ( .A(n40131), .B(n40130), .Z(n40135) );
  NAND U41163 ( .A(n40133), .B(n40132), .Z(n40134) );
  AND U41164 ( .A(n40135), .B(n40134), .Z(n40183) );
  XOR U41165 ( .A(n40184), .B(n40183), .Z(n40185) );
  NANDN U41166 ( .A(n40137), .B(n40136), .Z(n40141) );
  NANDN U41167 ( .A(n40139), .B(n40138), .Z(n40140) );
  NAND U41168 ( .A(n40141), .B(n40140), .Z(n40186) );
  XOR U41169 ( .A(n40185), .B(n40186), .Z(n40153) );
  OR U41170 ( .A(n40143), .B(n40142), .Z(n40147) );
  NANDN U41171 ( .A(n40145), .B(n40144), .Z(n40146) );
  NAND U41172 ( .A(n40147), .B(n40146), .Z(n40154) );
  XNOR U41173 ( .A(n40153), .B(n40154), .Z(n40155) );
  XNOR U41174 ( .A(n40156), .B(n40155), .Z(n40189) );
  XNOR U41175 ( .A(n40189), .B(sreg[1993]), .Z(n40191) );
  NAND U41176 ( .A(n40148), .B(sreg[1992]), .Z(n40152) );
  OR U41177 ( .A(n40150), .B(n40149), .Z(n40151) );
  AND U41178 ( .A(n40152), .B(n40151), .Z(n40190) );
  XOR U41179 ( .A(n40191), .B(n40190), .Z(c[1993]) );
  NANDN U41180 ( .A(n40154), .B(n40153), .Z(n40158) );
  NAND U41181 ( .A(n40156), .B(n40155), .Z(n40157) );
  NAND U41182 ( .A(n40158), .B(n40157), .Z(n40197) );
  NAND U41183 ( .A(b[0]), .B(a[978]), .Z(n40159) );
  XNOR U41184 ( .A(b[1]), .B(n40159), .Z(n40161) );
  NAND U41185 ( .A(n154), .B(a[977]), .Z(n40160) );
  AND U41186 ( .A(n40161), .B(n40160), .Z(n40214) );
  XOR U41187 ( .A(a[974]), .B(n42197), .Z(n40203) );
  NANDN U41188 ( .A(n40203), .B(n42173), .Z(n40164) );
  NANDN U41189 ( .A(n40162), .B(n42172), .Z(n40163) );
  NAND U41190 ( .A(n40164), .B(n40163), .Z(n40212) );
  NAND U41191 ( .A(b[7]), .B(a[970]), .Z(n40213) );
  XNOR U41192 ( .A(n40212), .B(n40213), .Z(n40215) );
  XOR U41193 ( .A(n40214), .B(n40215), .Z(n40221) );
  NANDN U41194 ( .A(n40165), .B(n42093), .Z(n40167) );
  XOR U41195 ( .A(n42134), .B(a[976]), .Z(n40206) );
  NANDN U41196 ( .A(n40206), .B(n42095), .Z(n40166) );
  NAND U41197 ( .A(n40167), .B(n40166), .Z(n40219) );
  NANDN U41198 ( .A(n40168), .B(n42231), .Z(n40170) );
  XOR U41199 ( .A(n243), .B(a[972]), .Z(n40209) );
  NANDN U41200 ( .A(n40209), .B(n42234), .Z(n40169) );
  AND U41201 ( .A(n40170), .B(n40169), .Z(n40218) );
  XNOR U41202 ( .A(n40219), .B(n40218), .Z(n40220) );
  XNOR U41203 ( .A(n40221), .B(n40220), .Z(n40225) );
  NANDN U41204 ( .A(n40172), .B(n40171), .Z(n40176) );
  NAND U41205 ( .A(n40174), .B(n40173), .Z(n40175) );
  AND U41206 ( .A(n40176), .B(n40175), .Z(n40224) );
  XOR U41207 ( .A(n40225), .B(n40224), .Z(n40226) );
  NANDN U41208 ( .A(n40178), .B(n40177), .Z(n40182) );
  NANDN U41209 ( .A(n40180), .B(n40179), .Z(n40181) );
  NAND U41210 ( .A(n40182), .B(n40181), .Z(n40227) );
  XOR U41211 ( .A(n40226), .B(n40227), .Z(n40194) );
  OR U41212 ( .A(n40184), .B(n40183), .Z(n40188) );
  NANDN U41213 ( .A(n40186), .B(n40185), .Z(n40187) );
  NAND U41214 ( .A(n40188), .B(n40187), .Z(n40195) );
  XNOR U41215 ( .A(n40194), .B(n40195), .Z(n40196) );
  XNOR U41216 ( .A(n40197), .B(n40196), .Z(n40230) );
  XNOR U41217 ( .A(n40230), .B(sreg[1994]), .Z(n40232) );
  NAND U41218 ( .A(n40189), .B(sreg[1993]), .Z(n40193) );
  OR U41219 ( .A(n40191), .B(n40190), .Z(n40192) );
  AND U41220 ( .A(n40193), .B(n40192), .Z(n40231) );
  XOR U41221 ( .A(n40232), .B(n40231), .Z(c[1994]) );
  NANDN U41222 ( .A(n40195), .B(n40194), .Z(n40199) );
  NAND U41223 ( .A(n40197), .B(n40196), .Z(n40198) );
  NAND U41224 ( .A(n40199), .B(n40198), .Z(n40238) );
  NAND U41225 ( .A(b[0]), .B(a[979]), .Z(n40200) );
  XNOR U41226 ( .A(b[1]), .B(n40200), .Z(n40202) );
  NAND U41227 ( .A(n154), .B(a[978]), .Z(n40201) );
  AND U41228 ( .A(n40202), .B(n40201), .Z(n40255) );
  XOR U41229 ( .A(a[975]), .B(n42197), .Z(n40244) );
  NANDN U41230 ( .A(n40244), .B(n42173), .Z(n40205) );
  NANDN U41231 ( .A(n40203), .B(n42172), .Z(n40204) );
  NAND U41232 ( .A(n40205), .B(n40204), .Z(n40253) );
  NAND U41233 ( .A(b[7]), .B(a[971]), .Z(n40254) );
  XNOR U41234 ( .A(n40253), .B(n40254), .Z(n40256) );
  XOR U41235 ( .A(n40255), .B(n40256), .Z(n40262) );
  NANDN U41236 ( .A(n40206), .B(n42093), .Z(n40208) );
  XOR U41237 ( .A(n42134), .B(a[977]), .Z(n40247) );
  NANDN U41238 ( .A(n40247), .B(n42095), .Z(n40207) );
  NAND U41239 ( .A(n40208), .B(n40207), .Z(n40260) );
  NANDN U41240 ( .A(n40209), .B(n42231), .Z(n40211) );
  XOR U41241 ( .A(n243), .B(a[973]), .Z(n40250) );
  NANDN U41242 ( .A(n40250), .B(n42234), .Z(n40210) );
  AND U41243 ( .A(n40211), .B(n40210), .Z(n40259) );
  XNOR U41244 ( .A(n40260), .B(n40259), .Z(n40261) );
  XNOR U41245 ( .A(n40262), .B(n40261), .Z(n40266) );
  NANDN U41246 ( .A(n40213), .B(n40212), .Z(n40217) );
  NAND U41247 ( .A(n40215), .B(n40214), .Z(n40216) );
  AND U41248 ( .A(n40217), .B(n40216), .Z(n40265) );
  XOR U41249 ( .A(n40266), .B(n40265), .Z(n40267) );
  NANDN U41250 ( .A(n40219), .B(n40218), .Z(n40223) );
  NANDN U41251 ( .A(n40221), .B(n40220), .Z(n40222) );
  NAND U41252 ( .A(n40223), .B(n40222), .Z(n40268) );
  XOR U41253 ( .A(n40267), .B(n40268), .Z(n40235) );
  OR U41254 ( .A(n40225), .B(n40224), .Z(n40229) );
  NANDN U41255 ( .A(n40227), .B(n40226), .Z(n40228) );
  NAND U41256 ( .A(n40229), .B(n40228), .Z(n40236) );
  XNOR U41257 ( .A(n40235), .B(n40236), .Z(n40237) );
  XNOR U41258 ( .A(n40238), .B(n40237), .Z(n40271) );
  XNOR U41259 ( .A(n40271), .B(sreg[1995]), .Z(n40273) );
  NAND U41260 ( .A(n40230), .B(sreg[1994]), .Z(n40234) );
  OR U41261 ( .A(n40232), .B(n40231), .Z(n40233) );
  AND U41262 ( .A(n40234), .B(n40233), .Z(n40272) );
  XOR U41263 ( .A(n40273), .B(n40272), .Z(c[1995]) );
  NANDN U41264 ( .A(n40236), .B(n40235), .Z(n40240) );
  NAND U41265 ( .A(n40238), .B(n40237), .Z(n40239) );
  NAND U41266 ( .A(n40240), .B(n40239), .Z(n40279) );
  NAND U41267 ( .A(b[0]), .B(a[980]), .Z(n40241) );
  XNOR U41268 ( .A(b[1]), .B(n40241), .Z(n40243) );
  NAND U41269 ( .A(n155), .B(a[979]), .Z(n40242) );
  AND U41270 ( .A(n40243), .B(n40242), .Z(n40296) );
  XOR U41271 ( .A(a[976]), .B(n42197), .Z(n40285) );
  NANDN U41272 ( .A(n40285), .B(n42173), .Z(n40246) );
  NANDN U41273 ( .A(n40244), .B(n42172), .Z(n40245) );
  NAND U41274 ( .A(n40246), .B(n40245), .Z(n40294) );
  NAND U41275 ( .A(b[7]), .B(a[972]), .Z(n40295) );
  XNOR U41276 ( .A(n40294), .B(n40295), .Z(n40297) );
  XOR U41277 ( .A(n40296), .B(n40297), .Z(n40303) );
  NANDN U41278 ( .A(n40247), .B(n42093), .Z(n40249) );
  XOR U41279 ( .A(n42134), .B(a[978]), .Z(n40288) );
  NANDN U41280 ( .A(n40288), .B(n42095), .Z(n40248) );
  NAND U41281 ( .A(n40249), .B(n40248), .Z(n40301) );
  NANDN U41282 ( .A(n40250), .B(n42231), .Z(n40252) );
  XOR U41283 ( .A(n243), .B(a[974]), .Z(n40291) );
  NANDN U41284 ( .A(n40291), .B(n42234), .Z(n40251) );
  AND U41285 ( .A(n40252), .B(n40251), .Z(n40300) );
  XNOR U41286 ( .A(n40301), .B(n40300), .Z(n40302) );
  XNOR U41287 ( .A(n40303), .B(n40302), .Z(n40307) );
  NANDN U41288 ( .A(n40254), .B(n40253), .Z(n40258) );
  NAND U41289 ( .A(n40256), .B(n40255), .Z(n40257) );
  AND U41290 ( .A(n40258), .B(n40257), .Z(n40306) );
  XOR U41291 ( .A(n40307), .B(n40306), .Z(n40308) );
  NANDN U41292 ( .A(n40260), .B(n40259), .Z(n40264) );
  NANDN U41293 ( .A(n40262), .B(n40261), .Z(n40263) );
  NAND U41294 ( .A(n40264), .B(n40263), .Z(n40309) );
  XOR U41295 ( .A(n40308), .B(n40309), .Z(n40276) );
  OR U41296 ( .A(n40266), .B(n40265), .Z(n40270) );
  NANDN U41297 ( .A(n40268), .B(n40267), .Z(n40269) );
  NAND U41298 ( .A(n40270), .B(n40269), .Z(n40277) );
  XNOR U41299 ( .A(n40276), .B(n40277), .Z(n40278) );
  XNOR U41300 ( .A(n40279), .B(n40278), .Z(n40312) );
  XNOR U41301 ( .A(n40312), .B(sreg[1996]), .Z(n40314) );
  NAND U41302 ( .A(n40271), .B(sreg[1995]), .Z(n40275) );
  OR U41303 ( .A(n40273), .B(n40272), .Z(n40274) );
  AND U41304 ( .A(n40275), .B(n40274), .Z(n40313) );
  XOR U41305 ( .A(n40314), .B(n40313), .Z(c[1996]) );
  NANDN U41306 ( .A(n40277), .B(n40276), .Z(n40281) );
  NAND U41307 ( .A(n40279), .B(n40278), .Z(n40280) );
  NAND U41308 ( .A(n40281), .B(n40280), .Z(n40320) );
  NAND U41309 ( .A(b[0]), .B(a[981]), .Z(n40282) );
  XNOR U41310 ( .A(b[1]), .B(n40282), .Z(n40284) );
  NAND U41311 ( .A(n155), .B(a[980]), .Z(n40283) );
  AND U41312 ( .A(n40284), .B(n40283), .Z(n40337) );
  XOR U41313 ( .A(a[977]), .B(n42197), .Z(n40326) );
  NANDN U41314 ( .A(n40326), .B(n42173), .Z(n40287) );
  NANDN U41315 ( .A(n40285), .B(n42172), .Z(n40286) );
  NAND U41316 ( .A(n40287), .B(n40286), .Z(n40335) );
  NAND U41317 ( .A(b[7]), .B(a[973]), .Z(n40336) );
  XNOR U41318 ( .A(n40335), .B(n40336), .Z(n40338) );
  XOR U41319 ( .A(n40337), .B(n40338), .Z(n40344) );
  NANDN U41320 ( .A(n40288), .B(n42093), .Z(n40290) );
  XOR U41321 ( .A(n42134), .B(a[979]), .Z(n40329) );
  NANDN U41322 ( .A(n40329), .B(n42095), .Z(n40289) );
  NAND U41323 ( .A(n40290), .B(n40289), .Z(n40342) );
  NANDN U41324 ( .A(n40291), .B(n42231), .Z(n40293) );
  XOR U41325 ( .A(n243), .B(a[975]), .Z(n40332) );
  NANDN U41326 ( .A(n40332), .B(n42234), .Z(n40292) );
  AND U41327 ( .A(n40293), .B(n40292), .Z(n40341) );
  XNOR U41328 ( .A(n40342), .B(n40341), .Z(n40343) );
  XNOR U41329 ( .A(n40344), .B(n40343), .Z(n40348) );
  NANDN U41330 ( .A(n40295), .B(n40294), .Z(n40299) );
  NAND U41331 ( .A(n40297), .B(n40296), .Z(n40298) );
  AND U41332 ( .A(n40299), .B(n40298), .Z(n40347) );
  XOR U41333 ( .A(n40348), .B(n40347), .Z(n40349) );
  NANDN U41334 ( .A(n40301), .B(n40300), .Z(n40305) );
  NANDN U41335 ( .A(n40303), .B(n40302), .Z(n40304) );
  NAND U41336 ( .A(n40305), .B(n40304), .Z(n40350) );
  XOR U41337 ( .A(n40349), .B(n40350), .Z(n40317) );
  OR U41338 ( .A(n40307), .B(n40306), .Z(n40311) );
  NANDN U41339 ( .A(n40309), .B(n40308), .Z(n40310) );
  NAND U41340 ( .A(n40311), .B(n40310), .Z(n40318) );
  XNOR U41341 ( .A(n40317), .B(n40318), .Z(n40319) );
  XNOR U41342 ( .A(n40320), .B(n40319), .Z(n40353) );
  XNOR U41343 ( .A(n40353), .B(sreg[1997]), .Z(n40355) );
  NAND U41344 ( .A(n40312), .B(sreg[1996]), .Z(n40316) );
  OR U41345 ( .A(n40314), .B(n40313), .Z(n40315) );
  AND U41346 ( .A(n40316), .B(n40315), .Z(n40354) );
  XOR U41347 ( .A(n40355), .B(n40354), .Z(c[1997]) );
  NANDN U41348 ( .A(n40318), .B(n40317), .Z(n40322) );
  NAND U41349 ( .A(n40320), .B(n40319), .Z(n40321) );
  NAND U41350 ( .A(n40322), .B(n40321), .Z(n40361) );
  NAND U41351 ( .A(b[0]), .B(a[982]), .Z(n40323) );
  XNOR U41352 ( .A(b[1]), .B(n40323), .Z(n40325) );
  NAND U41353 ( .A(n155), .B(a[981]), .Z(n40324) );
  AND U41354 ( .A(n40325), .B(n40324), .Z(n40378) );
  XOR U41355 ( .A(a[978]), .B(n42197), .Z(n40367) );
  NANDN U41356 ( .A(n40367), .B(n42173), .Z(n40328) );
  NANDN U41357 ( .A(n40326), .B(n42172), .Z(n40327) );
  NAND U41358 ( .A(n40328), .B(n40327), .Z(n40376) );
  NAND U41359 ( .A(b[7]), .B(a[974]), .Z(n40377) );
  XNOR U41360 ( .A(n40376), .B(n40377), .Z(n40379) );
  XOR U41361 ( .A(n40378), .B(n40379), .Z(n40385) );
  NANDN U41362 ( .A(n40329), .B(n42093), .Z(n40331) );
  XOR U41363 ( .A(n42134), .B(a[980]), .Z(n40370) );
  NANDN U41364 ( .A(n40370), .B(n42095), .Z(n40330) );
  NAND U41365 ( .A(n40331), .B(n40330), .Z(n40383) );
  NANDN U41366 ( .A(n40332), .B(n42231), .Z(n40334) );
  XOR U41367 ( .A(n243), .B(a[976]), .Z(n40373) );
  NANDN U41368 ( .A(n40373), .B(n42234), .Z(n40333) );
  AND U41369 ( .A(n40334), .B(n40333), .Z(n40382) );
  XNOR U41370 ( .A(n40383), .B(n40382), .Z(n40384) );
  XNOR U41371 ( .A(n40385), .B(n40384), .Z(n40389) );
  NANDN U41372 ( .A(n40336), .B(n40335), .Z(n40340) );
  NAND U41373 ( .A(n40338), .B(n40337), .Z(n40339) );
  AND U41374 ( .A(n40340), .B(n40339), .Z(n40388) );
  XOR U41375 ( .A(n40389), .B(n40388), .Z(n40390) );
  NANDN U41376 ( .A(n40342), .B(n40341), .Z(n40346) );
  NANDN U41377 ( .A(n40344), .B(n40343), .Z(n40345) );
  NAND U41378 ( .A(n40346), .B(n40345), .Z(n40391) );
  XOR U41379 ( .A(n40390), .B(n40391), .Z(n40358) );
  OR U41380 ( .A(n40348), .B(n40347), .Z(n40352) );
  NANDN U41381 ( .A(n40350), .B(n40349), .Z(n40351) );
  NAND U41382 ( .A(n40352), .B(n40351), .Z(n40359) );
  XNOR U41383 ( .A(n40358), .B(n40359), .Z(n40360) );
  XNOR U41384 ( .A(n40361), .B(n40360), .Z(n40394) );
  XNOR U41385 ( .A(n40394), .B(sreg[1998]), .Z(n40396) );
  NAND U41386 ( .A(n40353), .B(sreg[1997]), .Z(n40357) );
  OR U41387 ( .A(n40355), .B(n40354), .Z(n40356) );
  AND U41388 ( .A(n40357), .B(n40356), .Z(n40395) );
  XOR U41389 ( .A(n40396), .B(n40395), .Z(c[1998]) );
  NANDN U41390 ( .A(n40359), .B(n40358), .Z(n40363) );
  NAND U41391 ( .A(n40361), .B(n40360), .Z(n40362) );
  NAND U41392 ( .A(n40363), .B(n40362), .Z(n40402) );
  NAND U41393 ( .A(b[0]), .B(a[983]), .Z(n40364) );
  XNOR U41394 ( .A(b[1]), .B(n40364), .Z(n40366) );
  NAND U41395 ( .A(n155), .B(a[982]), .Z(n40365) );
  AND U41396 ( .A(n40366), .B(n40365), .Z(n40419) );
  XOR U41397 ( .A(a[979]), .B(n42197), .Z(n40408) );
  NANDN U41398 ( .A(n40408), .B(n42173), .Z(n40369) );
  NANDN U41399 ( .A(n40367), .B(n42172), .Z(n40368) );
  NAND U41400 ( .A(n40369), .B(n40368), .Z(n40417) );
  NAND U41401 ( .A(b[7]), .B(a[975]), .Z(n40418) );
  XNOR U41402 ( .A(n40417), .B(n40418), .Z(n40420) );
  XOR U41403 ( .A(n40419), .B(n40420), .Z(n40426) );
  NANDN U41404 ( .A(n40370), .B(n42093), .Z(n40372) );
  XOR U41405 ( .A(n42134), .B(a[981]), .Z(n40411) );
  NANDN U41406 ( .A(n40411), .B(n42095), .Z(n40371) );
  NAND U41407 ( .A(n40372), .B(n40371), .Z(n40424) );
  NANDN U41408 ( .A(n40373), .B(n42231), .Z(n40375) );
  XOR U41409 ( .A(n243), .B(a[977]), .Z(n40414) );
  NANDN U41410 ( .A(n40414), .B(n42234), .Z(n40374) );
  AND U41411 ( .A(n40375), .B(n40374), .Z(n40423) );
  XNOR U41412 ( .A(n40424), .B(n40423), .Z(n40425) );
  XNOR U41413 ( .A(n40426), .B(n40425), .Z(n40430) );
  NANDN U41414 ( .A(n40377), .B(n40376), .Z(n40381) );
  NAND U41415 ( .A(n40379), .B(n40378), .Z(n40380) );
  AND U41416 ( .A(n40381), .B(n40380), .Z(n40429) );
  XOR U41417 ( .A(n40430), .B(n40429), .Z(n40431) );
  NANDN U41418 ( .A(n40383), .B(n40382), .Z(n40387) );
  NANDN U41419 ( .A(n40385), .B(n40384), .Z(n40386) );
  NAND U41420 ( .A(n40387), .B(n40386), .Z(n40432) );
  XOR U41421 ( .A(n40431), .B(n40432), .Z(n40399) );
  OR U41422 ( .A(n40389), .B(n40388), .Z(n40393) );
  NANDN U41423 ( .A(n40391), .B(n40390), .Z(n40392) );
  NAND U41424 ( .A(n40393), .B(n40392), .Z(n40400) );
  XNOR U41425 ( .A(n40399), .B(n40400), .Z(n40401) );
  XNOR U41426 ( .A(n40402), .B(n40401), .Z(n40435) );
  XNOR U41427 ( .A(n40435), .B(sreg[1999]), .Z(n40437) );
  NAND U41428 ( .A(n40394), .B(sreg[1998]), .Z(n40398) );
  OR U41429 ( .A(n40396), .B(n40395), .Z(n40397) );
  AND U41430 ( .A(n40398), .B(n40397), .Z(n40436) );
  XOR U41431 ( .A(n40437), .B(n40436), .Z(c[1999]) );
  NANDN U41432 ( .A(n40400), .B(n40399), .Z(n40404) );
  NAND U41433 ( .A(n40402), .B(n40401), .Z(n40403) );
  NAND U41434 ( .A(n40404), .B(n40403), .Z(n40443) );
  NAND U41435 ( .A(b[0]), .B(a[984]), .Z(n40405) );
  XNOR U41436 ( .A(b[1]), .B(n40405), .Z(n40407) );
  NAND U41437 ( .A(n155), .B(a[983]), .Z(n40406) );
  AND U41438 ( .A(n40407), .B(n40406), .Z(n40460) );
  XOR U41439 ( .A(a[980]), .B(n42197), .Z(n40449) );
  NANDN U41440 ( .A(n40449), .B(n42173), .Z(n40410) );
  NANDN U41441 ( .A(n40408), .B(n42172), .Z(n40409) );
  NAND U41442 ( .A(n40410), .B(n40409), .Z(n40458) );
  NAND U41443 ( .A(b[7]), .B(a[976]), .Z(n40459) );
  XNOR U41444 ( .A(n40458), .B(n40459), .Z(n40461) );
  XOR U41445 ( .A(n40460), .B(n40461), .Z(n40467) );
  NANDN U41446 ( .A(n40411), .B(n42093), .Z(n40413) );
  XOR U41447 ( .A(n42134), .B(a[982]), .Z(n40452) );
  NANDN U41448 ( .A(n40452), .B(n42095), .Z(n40412) );
  NAND U41449 ( .A(n40413), .B(n40412), .Z(n40465) );
  NANDN U41450 ( .A(n40414), .B(n42231), .Z(n40416) );
  XOR U41451 ( .A(n243), .B(a[978]), .Z(n40455) );
  NANDN U41452 ( .A(n40455), .B(n42234), .Z(n40415) );
  AND U41453 ( .A(n40416), .B(n40415), .Z(n40464) );
  XNOR U41454 ( .A(n40465), .B(n40464), .Z(n40466) );
  XNOR U41455 ( .A(n40467), .B(n40466), .Z(n40471) );
  NANDN U41456 ( .A(n40418), .B(n40417), .Z(n40422) );
  NAND U41457 ( .A(n40420), .B(n40419), .Z(n40421) );
  AND U41458 ( .A(n40422), .B(n40421), .Z(n40470) );
  XOR U41459 ( .A(n40471), .B(n40470), .Z(n40472) );
  NANDN U41460 ( .A(n40424), .B(n40423), .Z(n40428) );
  NANDN U41461 ( .A(n40426), .B(n40425), .Z(n40427) );
  NAND U41462 ( .A(n40428), .B(n40427), .Z(n40473) );
  XOR U41463 ( .A(n40472), .B(n40473), .Z(n40440) );
  OR U41464 ( .A(n40430), .B(n40429), .Z(n40434) );
  NANDN U41465 ( .A(n40432), .B(n40431), .Z(n40433) );
  NAND U41466 ( .A(n40434), .B(n40433), .Z(n40441) );
  XNOR U41467 ( .A(n40440), .B(n40441), .Z(n40442) );
  XNOR U41468 ( .A(n40443), .B(n40442), .Z(n40476) );
  XNOR U41469 ( .A(n40476), .B(sreg[2000]), .Z(n40478) );
  NAND U41470 ( .A(n40435), .B(sreg[1999]), .Z(n40439) );
  OR U41471 ( .A(n40437), .B(n40436), .Z(n40438) );
  AND U41472 ( .A(n40439), .B(n40438), .Z(n40477) );
  XOR U41473 ( .A(n40478), .B(n40477), .Z(c[2000]) );
  NANDN U41474 ( .A(n40441), .B(n40440), .Z(n40445) );
  NAND U41475 ( .A(n40443), .B(n40442), .Z(n40444) );
  NAND U41476 ( .A(n40445), .B(n40444), .Z(n40484) );
  NAND U41477 ( .A(b[0]), .B(a[985]), .Z(n40446) );
  XNOR U41478 ( .A(b[1]), .B(n40446), .Z(n40448) );
  NAND U41479 ( .A(n155), .B(a[984]), .Z(n40447) );
  AND U41480 ( .A(n40448), .B(n40447), .Z(n40501) );
  XOR U41481 ( .A(a[981]), .B(n42197), .Z(n40490) );
  NANDN U41482 ( .A(n40490), .B(n42173), .Z(n40451) );
  NANDN U41483 ( .A(n40449), .B(n42172), .Z(n40450) );
  NAND U41484 ( .A(n40451), .B(n40450), .Z(n40499) );
  NAND U41485 ( .A(b[7]), .B(a[977]), .Z(n40500) );
  XNOR U41486 ( .A(n40499), .B(n40500), .Z(n40502) );
  XOR U41487 ( .A(n40501), .B(n40502), .Z(n40508) );
  NANDN U41488 ( .A(n40452), .B(n42093), .Z(n40454) );
  XOR U41489 ( .A(n42134), .B(a[983]), .Z(n40493) );
  NANDN U41490 ( .A(n40493), .B(n42095), .Z(n40453) );
  NAND U41491 ( .A(n40454), .B(n40453), .Z(n40506) );
  NANDN U41492 ( .A(n40455), .B(n42231), .Z(n40457) );
  XOR U41493 ( .A(n243), .B(a[979]), .Z(n40496) );
  NANDN U41494 ( .A(n40496), .B(n42234), .Z(n40456) );
  AND U41495 ( .A(n40457), .B(n40456), .Z(n40505) );
  XNOR U41496 ( .A(n40506), .B(n40505), .Z(n40507) );
  XNOR U41497 ( .A(n40508), .B(n40507), .Z(n40512) );
  NANDN U41498 ( .A(n40459), .B(n40458), .Z(n40463) );
  NAND U41499 ( .A(n40461), .B(n40460), .Z(n40462) );
  AND U41500 ( .A(n40463), .B(n40462), .Z(n40511) );
  XOR U41501 ( .A(n40512), .B(n40511), .Z(n40513) );
  NANDN U41502 ( .A(n40465), .B(n40464), .Z(n40469) );
  NANDN U41503 ( .A(n40467), .B(n40466), .Z(n40468) );
  NAND U41504 ( .A(n40469), .B(n40468), .Z(n40514) );
  XOR U41505 ( .A(n40513), .B(n40514), .Z(n40481) );
  OR U41506 ( .A(n40471), .B(n40470), .Z(n40475) );
  NANDN U41507 ( .A(n40473), .B(n40472), .Z(n40474) );
  NAND U41508 ( .A(n40475), .B(n40474), .Z(n40482) );
  XNOR U41509 ( .A(n40481), .B(n40482), .Z(n40483) );
  XNOR U41510 ( .A(n40484), .B(n40483), .Z(n40517) );
  XNOR U41511 ( .A(n40517), .B(sreg[2001]), .Z(n40519) );
  NAND U41512 ( .A(n40476), .B(sreg[2000]), .Z(n40480) );
  OR U41513 ( .A(n40478), .B(n40477), .Z(n40479) );
  AND U41514 ( .A(n40480), .B(n40479), .Z(n40518) );
  XOR U41515 ( .A(n40519), .B(n40518), .Z(c[2001]) );
  NANDN U41516 ( .A(n40482), .B(n40481), .Z(n40486) );
  NAND U41517 ( .A(n40484), .B(n40483), .Z(n40485) );
  NAND U41518 ( .A(n40486), .B(n40485), .Z(n40525) );
  NAND U41519 ( .A(b[0]), .B(a[986]), .Z(n40487) );
  XNOR U41520 ( .A(b[1]), .B(n40487), .Z(n40489) );
  NAND U41521 ( .A(n155), .B(a[985]), .Z(n40488) );
  AND U41522 ( .A(n40489), .B(n40488), .Z(n40542) );
  XOR U41523 ( .A(a[982]), .B(n42197), .Z(n40531) );
  NANDN U41524 ( .A(n40531), .B(n42173), .Z(n40492) );
  NANDN U41525 ( .A(n40490), .B(n42172), .Z(n40491) );
  NAND U41526 ( .A(n40492), .B(n40491), .Z(n40540) );
  NAND U41527 ( .A(b[7]), .B(a[978]), .Z(n40541) );
  XNOR U41528 ( .A(n40540), .B(n40541), .Z(n40543) );
  XOR U41529 ( .A(n40542), .B(n40543), .Z(n40549) );
  NANDN U41530 ( .A(n40493), .B(n42093), .Z(n40495) );
  XOR U41531 ( .A(n42134), .B(a[984]), .Z(n40534) );
  NANDN U41532 ( .A(n40534), .B(n42095), .Z(n40494) );
  NAND U41533 ( .A(n40495), .B(n40494), .Z(n40547) );
  NANDN U41534 ( .A(n40496), .B(n42231), .Z(n40498) );
  XOR U41535 ( .A(n243), .B(a[980]), .Z(n40537) );
  NANDN U41536 ( .A(n40537), .B(n42234), .Z(n40497) );
  AND U41537 ( .A(n40498), .B(n40497), .Z(n40546) );
  XNOR U41538 ( .A(n40547), .B(n40546), .Z(n40548) );
  XNOR U41539 ( .A(n40549), .B(n40548), .Z(n40553) );
  NANDN U41540 ( .A(n40500), .B(n40499), .Z(n40504) );
  NAND U41541 ( .A(n40502), .B(n40501), .Z(n40503) );
  AND U41542 ( .A(n40504), .B(n40503), .Z(n40552) );
  XOR U41543 ( .A(n40553), .B(n40552), .Z(n40554) );
  NANDN U41544 ( .A(n40506), .B(n40505), .Z(n40510) );
  NANDN U41545 ( .A(n40508), .B(n40507), .Z(n40509) );
  NAND U41546 ( .A(n40510), .B(n40509), .Z(n40555) );
  XOR U41547 ( .A(n40554), .B(n40555), .Z(n40522) );
  OR U41548 ( .A(n40512), .B(n40511), .Z(n40516) );
  NANDN U41549 ( .A(n40514), .B(n40513), .Z(n40515) );
  NAND U41550 ( .A(n40516), .B(n40515), .Z(n40523) );
  XNOR U41551 ( .A(n40522), .B(n40523), .Z(n40524) );
  XNOR U41552 ( .A(n40525), .B(n40524), .Z(n40558) );
  XNOR U41553 ( .A(n40558), .B(sreg[2002]), .Z(n40560) );
  NAND U41554 ( .A(n40517), .B(sreg[2001]), .Z(n40521) );
  OR U41555 ( .A(n40519), .B(n40518), .Z(n40520) );
  AND U41556 ( .A(n40521), .B(n40520), .Z(n40559) );
  XOR U41557 ( .A(n40560), .B(n40559), .Z(c[2002]) );
  NANDN U41558 ( .A(n40523), .B(n40522), .Z(n40527) );
  NAND U41559 ( .A(n40525), .B(n40524), .Z(n40526) );
  NAND U41560 ( .A(n40527), .B(n40526), .Z(n40566) );
  NAND U41561 ( .A(b[0]), .B(a[987]), .Z(n40528) );
  XNOR U41562 ( .A(b[1]), .B(n40528), .Z(n40530) );
  NAND U41563 ( .A(n156), .B(a[986]), .Z(n40529) );
  AND U41564 ( .A(n40530), .B(n40529), .Z(n40583) );
  XOR U41565 ( .A(a[983]), .B(n42197), .Z(n40572) );
  NANDN U41566 ( .A(n40572), .B(n42173), .Z(n40533) );
  NANDN U41567 ( .A(n40531), .B(n42172), .Z(n40532) );
  NAND U41568 ( .A(n40533), .B(n40532), .Z(n40581) );
  NAND U41569 ( .A(b[7]), .B(a[979]), .Z(n40582) );
  XNOR U41570 ( .A(n40581), .B(n40582), .Z(n40584) );
  XOR U41571 ( .A(n40583), .B(n40584), .Z(n40590) );
  NANDN U41572 ( .A(n40534), .B(n42093), .Z(n40536) );
  XOR U41573 ( .A(n42134), .B(a[985]), .Z(n40575) );
  NANDN U41574 ( .A(n40575), .B(n42095), .Z(n40535) );
  NAND U41575 ( .A(n40536), .B(n40535), .Z(n40588) );
  NANDN U41576 ( .A(n40537), .B(n42231), .Z(n40539) );
  XOR U41577 ( .A(n243), .B(a[981]), .Z(n40578) );
  NANDN U41578 ( .A(n40578), .B(n42234), .Z(n40538) );
  AND U41579 ( .A(n40539), .B(n40538), .Z(n40587) );
  XNOR U41580 ( .A(n40588), .B(n40587), .Z(n40589) );
  XNOR U41581 ( .A(n40590), .B(n40589), .Z(n40594) );
  NANDN U41582 ( .A(n40541), .B(n40540), .Z(n40545) );
  NAND U41583 ( .A(n40543), .B(n40542), .Z(n40544) );
  AND U41584 ( .A(n40545), .B(n40544), .Z(n40593) );
  XOR U41585 ( .A(n40594), .B(n40593), .Z(n40595) );
  NANDN U41586 ( .A(n40547), .B(n40546), .Z(n40551) );
  NANDN U41587 ( .A(n40549), .B(n40548), .Z(n40550) );
  NAND U41588 ( .A(n40551), .B(n40550), .Z(n40596) );
  XOR U41589 ( .A(n40595), .B(n40596), .Z(n40563) );
  OR U41590 ( .A(n40553), .B(n40552), .Z(n40557) );
  NANDN U41591 ( .A(n40555), .B(n40554), .Z(n40556) );
  NAND U41592 ( .A(n40557), .B(n40556), .Z(n40564) );
  XNOR U41593 ( .A(n40563), .B(n40564), .Z(n40565) );
  XNOR U41594 ( .A(n40566), .B(n40565), .Z(n40599) );
  XNOR U41595 ( .A(n40599), .B(sreg[2003]), .Z(n40601) );
  NAND U41596 ( .A(n40558), .B(sreg[2002]), .Z(n40562) );
  OR U41597 ( .A(n40560), .B(n40559), .Z(n40561) );
  AND U41598 ( .A(n40562), .B(n40561), .Z(n40600) );
  XOR U41599 ( .A(n40601), .B(n40600), .Z(c[2003]) );
  NANDN U41600 ( .A(n40564), .B(n40563), .Z(n40568) );
  NAND U41601 ( .A(n40566), .B(n40565), .Z(n40567) );
  NAND U41602 ( .A(n40568), .B(n40567), .Z(n40607) );
  NAND U41603 ( .A(b[0]), .B(a[988]), .Z(n40569) );
  XNOR U41604 ( .A(b[1]), .B(n40569), .Z(n40571) );
  NAND U41605 ( .A(n156), .B(a[987]), .Z(n40570) );
  AND U41606 ( .A(n40571), .B(n40570), .Z(n40624) );
  XOR U41607 ( .A(a[984]), .B(n42197), .Z(n40613) );
  NANDN U41608 ( .A(n40613), .B(n42173), .Z(n40574) );
  NANDN U41609 ( .A(n40572), .B(n42172), .Z(n40573) );
  NAND U41610 ( .A(n40574), .B(n40573), .Z(n40622) );
  NAND U41611 ( .A(b[7]), .B(a[980]), .Z(n40623) );
  XNOR U41612 ( .A(n40622), .B(n40623), .Z(n40625) );
  XOR U41613 ( .A(n40624), .B(n40625), .Z(n40631) );
  NANDN U41614 ( .A(n40575), .B(n42093), .Z(n40577) );
  XOR U41615 ( .A(n42134), .B(a[986]), .Z(n40616) );
  NANDN U41616 ( .A(n40616), .B(n42095), .Z(n40576) );
  NAND U41617 ( .A(n40577), .B(n40576), .Z(n40629) );
  NANDN U41618 ( .A(n40578), .B(n42231), .Z(n40580) );
  XOR U41619 ( .A(n243), .B(a[982]), .Z(n40619) );
  NANDN U41620 ( .A(n40619), .B(n42234), .Z(n40579) );
  AND U41621 ( .A(n40580), .B(n40579), .Z(n40628) );
  XNOR U41622 ( .A(n40629), .B(n40628), .Z(n40630) );
  XNOR U41623 ( .A(n40631), .B(n40630), .Z(n40635) );
  NANDN U41624 ( .A(n40582), .B(n40581), .Z(n40586) );
  NAND U41625 ( .A(n40584), .B(n40583), .Z(n40585) );
  AND U41626 ( .A(n40586), .B(n40585), .Z(n40634) );
  XOR U41627 ( .A(n40635), .B(n40634), .Z(n40636) );
  NANDN U41628 ( .A(n40588), .B(n40587), .Z(n40592) );
  NANDN U41629 ( .A(n40590), .B(n40589), .Z(n40591) );
  NAND U41630 ( .A(n40592), .B(n40591), .Z(n40637) );
  XOR U41631 ( .A(n40636), .B(n40637), .Z(n40604) );
  OR U41632 ( .A(n40594), .B(n40593), .Z(n40598) );
  NANDN U41633 ( .A(n40596), .B(n40595), .Z(n40597) );
  NAND U41634 ( .A(n40598), .B(n40597), .Z(n40605) );
  XNOR U41635 ( .A(n40604), .B(n40605), .Z(n40606) );
  XNOR U41636 ( .A(n40607), .B(n40606), .Z(n40640) );
  XNOR U41637 ( .A(n40640), .B(sreg[2004]), .Z(n40642) );
  NAND U41638 ( .A(n40599), .B(sreg[2003]), .Z(n40603) );
  OR U41639 ( .A(n40601), .B(n40600), .Z(n40602) );
  AND U41640 ( .A(n40603), .B(n40602), .Z(n40641) );
  XOR U41641 ( .A(n40642), .B(n40641), .Z(c[2004]) );
  NANDN U41642 ( .A(n40605), .B(n40604), .Z(n40609) );
  NAND U41643 ( .A(n40607), .B(n40606), .Z(n40608) );
  NAND U41644 ( .A(n40609), .B(n40608), .Z(n40648) );
  NAND U41645 ( .A(b[0]), .B(a[989]), .Z(n40610) );
  XNOR U41646 ( .A(b[1]), .B(n40610), .Z(n40612) );
  NAND U41647 ( .A(n156), .B(a[988]), .Z(n40611) );
  AND U41648 ( .A(n40612), .B(n40611), .Z(n40665) );
  XOR U41649 ( .A(a[985]), .B(n42197), .Z(n40654) );
  NANDN U41650 ( .A(n40654), .B(n42173), .Z(n40615) );
  NANDN U41651 ( .A(n40613), .B(n42172), .Z(n40614) );
  NAND U41652 ( .A(n40615), .B(n40614), .Z(n40663) );
  NAND U41653 ( .A(b[7]), .B(a[981]), .Z(n40664) );
  XNOR U41654 ( .A(n40663), .B(n40664), .Z(n40666) );
  XOR U41655 ( .A(n40665), .B(n40666), .Z(n40672) );
  NANDN U41656 ( .A(n40616), .B(n42093), .Z(n40618) );
  XOR U41657 ( .A(n42134), .B(a[987]), .Z(n40657) );
  NANDN U41658 ( .A(n40657), .B(n42095), .Z(n40617) );
  NAND U41659 ( .A(n40618), .B(n40617), .Z(n40670) );
  NANDN U41660 ( .A(n40619), .B(n42231), .Z(n40621) );
  XOR U41661 ( .A(n244), .B(a[983]), .Z(n40660) );
  NANDN U41662 ( .A(n40660), .B(n42234), .Z(n40620) );
  AND U41663 ( .A(n40621), .B(n40620), .Z(n40669) );
  XNOR U41664 ( .A(n40670), .B(n40669), .Z(n40671) );
  XNOR U41665 ( .A(n40672), .B(n40671), .Z(n40676) );
  NANDN U41666 ( .A(n40623), .B(n40622), .Z(n40627) );
  NAND U41667 ( .A(n40625), .B(n40624), .Z(n40626) );
  AND U41668 ( .A(n40627), .B(n40626), .Z(n40675) );
  XOR U41669 ( .A(n40676), .B(n40675), .Z(n40677) );
  NANDN U41670 ( .A(n40629), .B(n40628), .Z(n40633) );
  NANDN U41671 ( .A(n40631), .B(n40630), .Z(n40632) );
  NAND U41672 ( .A(n40633), .B(n40632), .Z(n40678) );
  XOR U41673 ( .A(n40677), .B(n40678), .Z(n40645) );
  OR U41674 ( .A(n40635), .B(n40634), .Z(n40639) );
  NANDN U41675 ( .A(n40637), .B(n40636), .Z(n40638) );
  NAND U41676 ( .A(n40639), .B(n40638), .Z(n40646) );
  XNOR U41677 ( .A(n40645), .B(n40646), .Z(n40647) );
  XNOR U41678 ( .A(n40648), .B(n40647), .Z(n40681) );
  XNOR U41679 ( .A(n40681), .B(sreg[2005]), .Z(n40683) );
  NAND U41680 ( .A(n40640), .B(sreg[2004]), .Z(n40644) );
  OR U41681 ( .A(n40642), .B(n40641), .Z(n40643) );
  AND U41682 ( .A(n40644), .B(n40643), .Z(n40682) );
  XOR U41683 ( .A(n40683), .B(n40682), .Z(c[2005]) );
  NANDN U41684 ( .A(n40646), .B(n40645), .Z(n40650) );
  NAND U41685 ( .A(n40648), .B(n40647), .Z(n40649) );
  NAND U41686 ( .A(n40650), .B(n40649), .Z(n40689) );
  NAND U41687 ( .A(b[0]), .B(a[990]), .Z(n40651) );
  XNOR U41688 ( .A(b[1]), .B(n40651), .Z(n40653) );
  NAND U41689 ( .A(n156), .B(a[989]), .Z(n40652) );
  AND U41690 ( .A(n40653), .B(n40652), .Z(n40706) );
  XOR U41691 ( .A(a[986]), .B(n42197), .Z(n40695) );
  NANDN U41692 ( .A(n40695), .B(n42173), .Z(n40656) );
  NANDN U41693 ( .A(n40654), .B(n42172), .Z(n40655) );
  NAND U41694 ( .A(n40656), .B(n40655), .Z(n40704) );
  NAND U41695 ( .A(b[7]), .B(a[982]), .Z(n40705) );
  XNOR U41696 ( .A(n40704), .B(n40705), .Z(n40707) );
  XOR U41697 ( .A(n40706), .B(n40707), .Z(n40713) );
  NANDN U41698 ( .A(n40657), .B(n42093), .Z(n40659) );
  XOR U41699 ( .A(n42134), .B(a[988]), .Z(n40698) );
  NANDN U41700 ( .A(n40698), .B(n42095), .Z(n40658) );
  NAND U41701 ( .A(n40659), .B(n40658), .Z(n40711) );
  NANDN U41702 ( .A(n40660), .B(n42231), .Z(n40662) );
  XOR U41703 ( .A(n244), .B(a[984]), .Z(n40701) );
  NANDN U41704 ( .A(n40701), .B(n42234), .Z(n40661) );
  AND U41705 ( .A(n40662), .B(n40661), .Z(n40710) );
  XNOR U41706 ( .A(n40711), .B(n40710), .Z(n40712) );
  XNOR U41707 ( .A(n40713), .B(n40712), .Z(n40717) );
  NANDN U41708 ( .A(n40664), .B(n40663), .Z(n40668) );
  NAND U41709 ( .A(n40666), .B(n40665), .Z(n40667) );
  AND U41710 ( .A(n40668), .B(n40667), .Z(n40716) );
  XOR U41711 ( .A(n40717), .B(n40716), .Z(n40718) );
  NANDN U41712 ( .A(n40670), .B(n40669), .Z(n40674) );
  NANDN U41713 ( .A(n40672), .B(n40671), .Z(n40673) );
  NAND U41714 ( .A(n40674), .B(n40673), .Z(n40719) );
  XOR U41715 ( .A(n40718), .B(n40719), .Z(n40686) );
  OR U41716 ( .A(n40676), .B(n40675), .Z(n40680) );
  NANDN U41717 ( .A(n40678), .B(n40677), .Z(n40679) );
  NAND U41718 ( .A(n40680), .B(n40679), .Z(n40687) );
  XNOR U41719 ( .A(n40686), .B(n40687), .Z(n40688) );
  XNOR U41720 ( .A(n40689), .B(n40688), .Z(n40722) );
  XNOR U41721 ( .A(n40722), .B(sreg[2006]), .Z(n40724) );
  NAND U41722 ( .A(n40681), .B(sreg[2005]), .Z(n40685) );
  OR U41723 ( .A(n40683), .B(n40682), .Z(n40684) );
  AND U41724 ( .A(n40685), .B(n40684), .Z(n40723) );
  XOR U41725 ( .A(n40724), .B(n40723), .Z(c[2006]) );
  NANDN U41726 ( .A(n40687), .B(n40686), .Z(n40691) );
  NAND U41727 ( .A(n40689), .B(n40688), .Z(n40690) );
  NAND U41728 ( .A(n40691), .B(n40690), .Z(n40730) );
  NAND U41729 ( .A(b[0]), .B(a[991]), .Z(n40692) );
  XNOR U41730 ( .A(b[1]), .B(n40692), .Z(n40694) );
  NAND U41731 ( .A(n156), .B(a[990]), .Z(n40693) );
  AND U41732 ( .A(n40694), .B(n40693), .Z(n40747) );
  XOR U41733 ( .A(a[987]), .B(n42197), .Z(n40736) );
  NANDN U41734 ( .A(n40736), .B(n42173), .Z(n40697) );
  NANDN U41735 ( .A(n40695), .B(n42172), .Z(n40696) );
  NAND U41736 ( .A(n40697), .B(n40696), .Z(n40745) );
  NAND U41737 ( .A(b[7]), .B(a[983]), .Z(n40746) );
  XNOR U41738 ( .A(n40745), .B(n40746), .Z(n40748) );
  XOR U41739 ( .A(n40747), .B(n40748), .Z(n40754) );
  NANDN U41740 ( .A(n40698), .B(n42093), .Z(n40700) );
  XOR U41741 ( .A(n42134), .B(a[989]), .Z(n40739) );
  NANDN U41742 ( .A(n40739), .B(n42095), .Z(n40699) );
  NAND U41743 ( .A(n40700), .B(n40699), .Z(n40752) );
  NANDN U41744 ( .A(n40701), .B(n42231), .Z(n40703) );
  XOR U41745 ( .A(n244), .B(a[985]), .Z(n40742) );
  NANDN U41746 ( .A(n40742), .B(n42234), .Z(n40702) );
  AND U41747 ( .A(n40703), .B(n40702), .Z(n40751) );
  XNOR U41748 ( .A(n40752), .B(n40751), .Z(n40753) );
  XNOR U41749 ( .A(n40754), .B(n40753), .Z(n40758) );
  NANDN U41750 ( .A(n40705), .B(n40704), .Z(n40709) );
  NAND U41751 ( .A(n40707), .B(n40706), .Z(n40708) );
  AND U41752 ( .A(n40709), .B(n40708), .Z(n40757) );
  XOR U41753 ( .A(n40758), .B(n40757), .Z(n40759) );
  NANDN U41754 ( .A(n40711), .B(n40710), .Z(n40715) );
  NANDN U41755 ( .A(n40713), .B(n40712), .Z(n40714) );
  NAND U41756 ( .A(n40715), .B(n40714), .Z(n40760) );
  XOR U41757 ( .A(n40759), .B(n40760), .Z(n40727) );
  OR U41758 ( .A(n40717), .B(n40716), .Z(n40721) );
  NANDN U41759 ( .A(n40719), .B(n40718), .Z(n40720) );
  NAND U41760 ( .A(n40721), .B(n40720), .Z(n40728) );
  XNOR U41761 ( .A(n40727), .B(n40728), .Z(n40729) );
  XNOR U41762 ( .A(n40730), .B(n40729), .Z(n40763) );
  XNOR U41763 ( .A(n40763), .B(sreg[2007]), .Z(n40765) );
  NAND U41764 ( .A(n40722), .B(sreg[2006]), .Z(n40726) );
  OR U41765 ( .A(n40724), .B(n40723), .Z(n40725) );
  AND U41766 ( .A(n40726), .B(n40725), .Z(n40764) );
  XOR U41767 ( .A(n40765), .B(n40764), .Z(c[2007]) );
  NANDN U41768 ( .A(n40728), .B(n40727), .Z(n40732) );
  NAND U41769 ( .A(n40730), .B(n40729), .Z(n40731) );
  NAND U41770 ( .A(n40732), .B(n40731), .Z(n40771) );
  NAND U41771 ( .A(b[0]), .B(a[992]), .Z(n40733) );
  XNOR U41772 ( .A(b[1]), .B(n40733), .Z(n40735) );
  NAND U41773 ( .A(n156), .B(a[991]), .Z(n40734) );
  AND U41774 ( .A(n40735), .B(n40734), .Z(n40788) );
  XOR U41775 ( .A(a[988]), .B(n42197), .Z(n40777) );
  NANDN U41776 ( .A(n40777), .B(n42173), .Z(n40738) );
  NANDN U41777 ( .A(n40736), .B(n42172), .Z(n40737) );
  NAND U41778 ( .A(n40738), .B(n40737), .Z(n40786) );
  NAND U41779 ( .A(b[7]), .B(a[984]), .Z(n40787) );
  XNOR U41780 ( .A(n40786), .B(n40787), .Z(n40789) );
  XOR U41781 ( .A(n40788), .B(n40789), .Z(n40795) );
  NANDN U41782 ( .A(n40739), .B(n42093), .Z(n40741) );
  XOR U41783 ( .A(n42134), .B(a[990]), .Z(n40780) );
  NANDN U41784 ( .A(n40780), .B(n42095), .Z(n40740) );
  NAND U41785 ( .A(n40741), .B(n40740), .Z(n40793) );
  NANDN U41786 ( .A(n40742), .B(n42231), .Z(n40744) );
  XOR U41787 ( .A(n244), .B(a[986]), .Z(n40783) );
  NANDN U41788 ( .A(n40783), .B(n42234), .Z(n40743) );
  AND U41789 ( .A(n40744), .B(n40743), .Z(n40792) );
  XNOR U41790 ( .A(n40793), .B(n40792), .Z(n40794) );
  XNOR U41791 ( .A(n40795), .B(n40794), .Z(n40799) );
  NANDN U41792 ( .A(n40746), .B(n40745), .Z(n40750) );
  NAND U41793 ( .A(n40748), .B(n40747), .Z(n40749) );
  AND U41794 ( .A(n40750), .B(n40749), .Z(n40798) );
  XOR U41795 ( .A(n40799), .B(n40798), .Z(n40800) );
  NANDN U41796 ( .A(n40752), .B(n40751), .Z(n40756) );
  NANDN U41797 ( .A(n40754), .B(n40753), .Z(n40755) );
  NAND U41798 ( .A(n40756), .B(n40755), .Z(n40801) );
  XOR U41799 ( .A(n40800), .B(n40801), .Z(n40768) );
  OR U41800 ( .A(n40758), .B(n40757), .Z(n40762) );
  NANDN U41801 ( .A(n40760), .B(n40759), .Z(n40761) );
  NAND U41802 ( .A(n40762), .B(n40761), .Z(n40769) );
  XNOR U41803 ( .A(n40768), .B(n40769), .Z(n40770) );
  XNOR U41804 ( .A(n40771), .B(n40770), .Z(n40804) );
  XNOR U41805 ( .A(n40804), .B(sreg[2008]), .Z(n40806) );
  NAND U41806 ( .A(n40763), .B(sreg[2007]), .Z(n40767) );
  OR U41807 ( .A(n40765), .B(n40764), .Z(n40766) );
  AND U41808 ( .A(n40767), .B(n40766), .Z(n40805) );
  XOR U41809 ( .A(n40806), .B(n40805), .Z(c[2008]) );
  NANDN U41810 ( .A(n40769), .B(n40768), .Z(n40773) );
  NAND U41811 ( .A(n40771), .B(n40770), .Z(n40772) );
  NAND U41812 ( .A(n40773), .B(n40772), .Z(n40812) );
  NAND U41813 ( .A(b[0]), .B(a[993]), .Z(n40774) );
  XNOR U41814 ( .A(b[1]), .B(n40774), .Z(n40776) );
  NAND U41815 ( .A(n156), .B(a[992]), .Z(n40775) );
  AND U41816 ( .A(n40776), .B(n40775), .Z(n40829) );
  XOR U41817 ( .A(a[989]), .B(n42197), .Z(n40818) );
  NANDN U41818 ( .A(n40818), .B(n42173), .Z(n40779) );
  NANDN U41819 ( .A(n40777), .B(n42172), .Z(n40778) );
  NAND U41820 ( .A(n40779), .B(n40778), .Z(n40827) );
  NAND U41821 ( .A(b[7]), .B(a[985]), .Z(n40828) );
  XNOR U41822 ( .A(n40827), .B(n40828), .Z(n40830) );
  XOR U41823 ( .A(n40829), .B(n40830), .Z(n40836) );
  NANDN U41824 ( .A(n40780), .B(n42093), .Z(n40782) );
  XOR U41825 ( .A(n42134), .B(a[991]), .Z(n40821) );
  NANDN U41826 ( .A(n40821), .B(n42095), .Z(n40781) );
  NAND U41827 ( .A(n40782), .B(n40781), .Z(n40834) );
  NANDN U41828 ( .A(n40783), .B(n42231), .Z(n40785) );
  XOR U41829 ( .A(n244), .B(a[987]), .Z(n40824) );
  NANDN U41830 ( .A(n40824), .B(n42234), .Z(n40784) );
  AND U41831 ( .A(n40785), .B(n40784), .Z(n40833) );
  XNOR U41832 ( .A(n40834), .B(n40833), .Z(n40835) );
  XNOR U41833 ( .A(n40836), .B(n40835), .Z(n40840) );
  NANDN U41834 ( .A(n40787), .B(n40786), .Z(n40791) );
  NAND U41835 ( .A(n40789), .B(n40788), .Z(n40790) );
  AND U41836 ( .A(n40791), .B(n40790), .Z(n40839) );
  XOR U41837 ( .A(n40840), .B(n40839), .Z(n40841) );
  NANDN U41838 ( .A(n40793), .B(n40792), .Z(n40797) );
  NANDN U41839 ( .A(n40795), .B(n40794), .Z(n40796) );
  NAND U41840 ( .A(n40797), .B(n40796), .Z(n40842) );
  XOR U41841 ( .A(n40841), .B(n40842), .Z(n40809) );
  OR U41842 ( .A(n40799), .B(n40798), .Z(n40803) );
  NANDN U41843 ( .A(n40801), .B(n40800), .Z(n40802) );
  NAND U41844 ( .A(n40803), .B(n40802), .Z(n40810) );
  XNOR U41845 ( .A(n40809), .B(n40810), .Z(n40811) );
  XNOR U41846 ( .A(n40812), .B(n40811), .Z(n40845) );
  XNOR U41847 ( .A(n40845), .B(sreg[2009]), .Z(n40847) );
  NAND U41848 ( .A(n40804), .B(sreg[2008]), .Z(n40808) );
  OR U41849 ( .A(n40806), .B(n40805), .Z(n40807) );
  AND U41850 ( .A(n40808), .B(n40807), .Z(n40846) );
  XOR U41851 ( .A(n40847), .B(n40846), .Z(c[2009]) );
  NANDN U41852 ( .A(n40810), .B(n40809), .Z(n40814) );
  NAND U41853 ( .A(n40812), .B(n40811), .Z(n40813) );
  NAND U41854 ( .A(n40814), .B(n40813), .Z(n40853) );
  NAND U41855 ( .A(b[0]), .B(a[994]), .Z(n40815) );
  XNOR U41856 ( .A(b[1]), .B(n40815), .Z(n40817) );
  NAND U41857 ( .A(n157), .B(a[993]), .Z(n40816) );
  AND U41858 ( .A(n40817), .B(n40816), .Z(n40870) );
  XOR U41859 ( .A(a[990]), .B(n42197), .Z(n40859) );
  NANDN U41860 ( .A(n40859), .B(n42173), .Z(n40820) );
  NANDN U41861 ( .A(n40818), .B(n42172), .Z(n40819) );
  NAND U41862 ( .A(n40820), .B(n40819), .Z(n40868) );
  NAND U41863 ( .A(b[7]), .B(a[986]), .Z(n40869) );
  XNOR U41864 ( .A(n40868), .B(n40869), .Z(n40871) );
  XOR U41865 ( .A(n40870), .B(n40871), .Z(n40877) );
  NANDN U41866 ( .A(n40821), .B(n42093), .Z(n40823) );
  XOR U41867 ( .A(n42134), .B(a[992]), .Z(n40862) );
  NANDN U41868 ( .A(n40862), .B(n42095), .Z(n40822) );
  NAND U41869 ( .A(n40823), .B(n40822), .Z(n40875) );
  NANDN U41870 ( .A(n40824), .B(n42231), .Z(n40826) );
  XOR U41871 ( .A(n244), .B(a[988]), .Z(n40865) );
  NANDN U41872 ( .A(n40865), .B(n42234), .Z(n40825) );
  AND U41873 ( .A(n40826), .B(n40825), .Z(n40874) );
  XNOR U41874 ( .A(n40875), .B(n40874), .Z(n40876) );
  XNOR U41875 ( .A(n40877), .B(n40876), .Z(n40881) );
  NANDN U41876 ( .A(n40828), .B(n40827), .Z(n40832) );
  NAND U41877 ( .A(n40830), .B(n40829), .Z(n40831) );
  AND U41878 ( .A(n40832), .B(n40831), .Z(n40880) );
  XOR U41879 ( .A(n40881), .B(n40880), .Z(n40882) );
  NANDN U41880 ( .A(n40834), .B(n40833), .Z(n40838) );
  NANDN U41881 ( .A(n40836), .B(n40835), .Z(n40837) );
  NAND U41882 ( .A(n40838), .B(n40837), .Z(n40883) );
  XOR U41883 ( .A(n40882), .B(n40883), .Z(n40850) );
  OR U41884 ( .A(n40840), .B(n40839), .Z(n40844) );
  NANDN U41885 ( .A(n40842), .B(n40841), .Z(n40843) );
  NAND U41886 ( .A(n40844), .B(n40843), .Z(n40851) );
  XNOR U41887 ( .A(n40850), .B(n40851), .Z(n40852) );
  XNOR U41888 ( .A(n40853), .B(n40852), .Z(n40886) );
  XNOR U41889 ( .A(n40886), .B(sreg[2010]), .Z(n40888) );
  NAND U41890 ( .A(n40845), .B(sreg[2009]), .Z(n40849) );
  OR U41891 ( .A(n40847), .B(n40846), .Z(n40848) );
  AND U41892 ( .A(n40849), .B(n40848), .Z(n40887) );
  XOR U41893 ( .A(n40888), .B(n40887), .Z(c[2010]) );
  NANDN U41894 ( .A(n40851), .B(n40850), .Z(n40855) );
  NAND U41895 ( .A(n40853), .B(n40852), .Z(n40854) );
  NAND U41896 ( .A(n40855), .B(n40854), .Z(n40894) );
  NAND U41897 ( .A(b[0]), .B(a[995]), .Z(n40856) );
  XNOR U41898 ( .A(b[1]), .B(n40856), .Z(n40858) );
  NAND U41899 ( .A(n157), .B(a[994]), .Z(n40857) );
  AND U41900 ( .A(n40858), .B(n40857), .Z(n40911) );
  XOR U41901 ( .A(a[991]), .B(n42197), .Z(n40900) );
  NANDN U41902 ( .A(n40900), .B(n42173), .Z(n40861) );
  NANDN U41903 ( .A(n40859), .B(n42172), .Z(n40860) );
  NAND U41904 ( .A(n40861), .B(n40860), .Z(n40909) );
  NAND U41905 ( .A(b[7]), .B(a[987]), .Z(n40910) );
  XNOR U41906 ( .A(n40909), .B(n40910), .Z(n40912) );
  XOR U41907 ( .A(n40911), .B(n40912), .Z(n40918) );
  NANDN U41908 ( .A(n40862), .B(n42093), .Z(n40864) );
  XOR U41909 ( .A(n42134), .B(a[993]), .Z(n40903) );
  NANDN U41910 ( .A(n40903), .B(n42095), .Z(n40863) );
  NAND U41911 ( .A(n40864), .B(n40863), .Z(n40916) );
  NANDN U41912 ( .A(n40865), .B(n42231), .Z(n40867) );
  XOR U41913 ( .A(n244), .B(a[989]), .Z(n40906) );
  NANDN U41914 ( .A(n40906), .B(n42234), .Z(n40866) );
  AND U41915 ( .A(n40867), .B(n40866), .Z(n40915) );
  XNOR U41916 ( .A(n40916), .B(n40915), .Z(n40917) );
  XNOR U41917 ( .A(n40918), .B(n40917), .Z(n40922) );
  NANDN U41918 ( .A(n40869), .B(n40868), .Z(n40873) );
  NAND U41919 ( .A(n40871), .B(n40870), .Z(n40872) );
  AND U41920 ( .A(n40873), .B(n40872), .Z(n40921) );
  XOR U41921 ( .A(n40922), .B(n40921), .Z(n40923) );
  NANDN U41922 ( .A(n40875), .B(n40874), .Z(n40879) );
  NANDN U41923 ( .A(n40877), .B(n40876), .Z(n40878) );
  NAND U41924 ( .A(n40879), .B(n40878), .Z(n40924) );
  XOR U41925 ( .A(n40923), .B(n40924), .Z(n40891) );
  OR U41926 ( .A(n40881), .B(n40880), .Z(n40885) );
  NANDN U41927 ( .A(n40883), .B(n40882), .Z(n40884) );
  NAND U41928 ( .A(n40885), .B(n40884), .Z(n40892) );
  XNOR U41929 ( .A(n40891), .B(n40892), .Z(n40893) );
  XNOR U41930 ( .A(n40894), .B(n40893), .Z(n40927) );
  XNOR U41931 ( .A(n40927), .B(sreg[2011]), .Z(n40929) );
  NAND U41932 ( .A(n40886), .B(sreg[2010]), .Z(n40890) );
  OR U41933 ( .A(n40888), .B(n40887), .Z(n40889) );
  AND U41934 ( .A(n40890), .B(n40889), .Z(n40928) );
  XOR U41935 ( .A(n40929), .B(n40928), .Z(c[2011]) );
  NANDN U41936 ( .A(n40892), .B(n40891), .Z(n40896) );
  NAND U41937 ( .A(n40894), .B(n40893), .Z(n40895) );
  NAND U41938 ( .A(n40896), .B(n40895), .Z(n40935) );
  NAND U41939 ( .A(b[0]), .B(a[996]), .Z(n40897) );
  XNOR U41940 ( .A(b[1]), .B(n40897), .Z(n40899) );
  NAND U41941 ( .A(n157), .B(a[995]), .Z(n40898) );
  AND U41942 ( .A(n40899), .B(n40898), .Z(n40952) );
  XOR U41943 ( .A(a[992]), .B(n42197), .Z(n40941) );
  NANDN U41944 ( .A(n40941), .B(n42173), .Z(n40902) );
  NANDN U41945 ( .A(n40900), .B(n42172), .Z(n40901) );
  NAND U41946 ( .A(n40902), .B(n40901), .Z(n40950) );
  NAND U41947 ( .A(b[7]), .B(a[988]), .Z(n40951) );
  XNOR U41948 ( .A(n40950), .B(n40951), .Z(n40953) );
  XOR U41949 ( .A(n40952), .B(n40953), .Z(n40959) );
  NANDN U41950 ( .A(n40903), .B(n42093), .Z(n40905) );
  XOR U41951 ( .A(n42134), .B(a[994]), .Z(n40944) );
  NANDN U41952 ( .A(n40944), .B(n42095), .Z(n40904) );
  NAND U41953 ( .A(n40905), .B(n40904), .Z(n40957) );
  NANDN U41954 ( .A(n40906), .B(n42231), .Z(n40908) );
  XOR U41955 ( .A(n244), .B(a[990]), .Z(n40947) );
  NANDN U41956 ( .A(n40947), .B(n42234), .Z(n40907) );
  AND U41957 ( .A(n40908), .B(n40907), .Z(n40956) );
  XNOR U41958 ( .A(n40957), .B(n40956), .Z(n40958) );
  XNOR U41959 ( .A(n40959), .B(n40958), .Z(n40963) );
  NANDN U41960 ( .A(n40910), .B(n40909), .Z(n40914) );
  NAND U41961 ( .A(n40912), .B(n40911), .Z(n40913) );
  AND U41962 ( .A(n40914), .B(n40913), .Z(n40962) );
  XOR U41963 ( .A(n40963), .B(n40962), .Z(n40964) );
  NANDN U41964 ( .A(n40916), .B(n40915), .Z(n40920) );
  NANDN U41965 ( .A(n40918), .B(n40917), .Z(n40919) );
  NAND U41966 ( .A(n40920), .B(n40919), .Z(n40965) );
  XOR U41967 ( .A(n40964), .B(n40965), .Z(n40932) );
  OR U41968 ( .A(n40922), .B(n40921), .Z(n40926) );
  NANDN U41969 ( .A(n40924), .B(n40923), .Z(n40925) );
  NAND U41970 ( .A(n40926), .B(n40925), .Z(n40933) );
  XNOR U41971 ( .A(n40932), .B(n40933), .Z(n40934) );
  XNOR U41972 ( .A(n40935), .B(n40934), .Z(n40968) );
  XNOR U41973 ( .A(n40968), .B(sreg[2012]), .Z(n40970) );
  NAND U41974 ( .A(n40927), .B(sreg[2011]), .Z(n40931) );
  OR U41975 ( .A(n40929), .B(n40928), .Z(n40930) );
  AND U41976 ( .A(n40931), .B(n40930), .Z(n40969) );
  XOR U41977 ( .A(n40970), .B(n40969), .Z(c[2012]) );
  NANDN U41978 ( .A(n40933), .B(n40932), .Z(n40937) );
  NAND U41979 ( .A(n40935), .B(n40934), .Z(n40936) );
  NAND U41980 ( .A(n40937), .B(n40936), .Z(n40976) );
  NAND U41981 ( .A(b[0]), .B(a[997]), .Z(n40938) );
  XNOR U41982 ( .A(b[1]), .B(n40938), .Z(n40940) );
  NAND U41983 ( .A(n157), .B(a[996]), .Z(n40939) );
  AND U41984 ( .A(n40940), .B(n40939), .Z(n40993) );
  XOR U41985 ( .A(a[993]), .B(n42197), .Z(n40982) );
  NANDN U41986 ( .A(n40982), .B(n42173), .Z(n40943) );
  NANDN U41987 ( .A(n40941), .B(n42172), .Z(n40942) );
  NAND U41988 ( .A(n40943), .B(n40942), .Z(n40991) );
  NAND U41989 ( .A(b[7]), .B(a[989]), .Z(n40992) );
  XNOR U41990 ( .A(n40991), .B(n40992), .Z(n40994) );
  XOR U41991 ( .A(n40993), .B(n40994), .Z(n41000) );
  NANDN U41992 ( .A(n40944), .B(n42093), .Z(n40946) );
  XOR U41993 ( .A(n42134), .B(a[995]), .Z(n40985) );
  NANDN U41994 ( .A(n40985), .B(n42095), .Z(n40945) );
  NAND U41995 ( .A(n40946), .B(n40945), .Z(n40998) );
  NANDN U41996 ( .A(n40947), .B(n42231), .Z(n40949) );
  XOR U41997 ( .A(n244), .B(a[991]), .Z(n40988) );
  NANDN U41998 ( .A(n40988), .B(n42234), .Z(n40948) );
  AND U41999 ( .A(n40949), .B(n40948), .Z(n40997) );
  XNOR U42000 ( .A(n40998), .B(n40997), .Z(n40999) );
  XNOR U42001 ( .A(n41000), .B(n40999), .Z(n41004) );
  NANDN U42002 ( .A(n40951), .B(n40950), .Z(n40955) );
  NAND U42003 ( .A(n40953), .B(n40952), .Z(n40954) );
  AND U42004 ( .A(n40955), .B(n40954), .Z(n41003) );
  XOR U42005 ( .A(n41004), .B(n41003), .Z(n41005) );
  NANDN U42006 ( .A(n40957), .B(n40956), .Z(n40961) );
  NANDN U42007 ( .A(n40959), .B(n40958), .Z(n40960) );
  NAND U42008 ( .A(n40961), .B(n40960), .Z(n41006) );
  XOR U42009 ( .A(n41005), .B(n41006), .Z(n40973) );
  OR U42010 ( .A(n40963), .B(n40962), .Z(n40967) );
  NANDN U42011 ( .A(n40965), .B(n40964), .Z(n40966) );
  NAND U42012 ( .A(n40967), .B(n40966), .Z(n40974) );
  XNOR U42013 ( .A(n40973), .B(n40974), .Z(n40975) );
  XNOR U42014 ( .A(n40976), .B(n40975), .Z(n41009) );
  XNOR U42015 ( .A(n41009), .B(sreg[2013]), .Z(n41011) );
  NAND U42016 ( .A(n40968), .B(sreg[2012]), .Z(n40972) );
  OR U42017 ( .A(n40970), .B(n40969), .Z(n40971) );
  AND U42018 ( .A(n40972), .B(n40971), .Z(n41010) );
  XOR U42019 ( .A(n41011), .B(n41010), .Z(c[2013]) );
  NANDN U42020 ( .A(n40974), .B(n40973), .Z(n40978) );
  NAND U42021 ( .A(n40976), .B(n40975), .Z(n40977) );
  NAND U42022 ( .A(n40978), .B(n40977), .Z(n41017) );
  NAND U42023 ( .A(b[0]), .B(a[998]), .Z(n40979) );
  XNOR U42024 ( .A(b[1]), .B(n40979), .Z(n40981) );
  NAND U42025 ( .A(n157), .B(a[997]), .Z(n40980) );
  AND U42026 ( .A(n40981), .B(n40980), .Z(n41034) );
  XOR U42027 ( .A(a[994]), .B(n42197), .Z(n41023) );
  NANDN U42028 ( .A(n41023), .B(n42173), .Z(n40984) );
  NANDN U42029 ( .A(n40982), .B(n42172), .Z(n40983) );
  NAND U42030 ( .A(n40984), .B(n40983), .Z(n41032) );
  NAND U42031 ( .A(b[7]), .B(a[990]), .Z(n41033) );
  XNOR U42032 ( .A(n41032), .B(n41033), .Z(n41035) );
  XOR U42033 ( .A(n41034), .B(n41035), .Z(n41041) );
  NANDN U42034 ( .A(n40985), .B(n42093), .Z(n40987) );
  XOR U42035 ( .A(n42134), .B(a[996]), .Z(n41026) );
  NANDN U42036 ( .A(n41026), .B(n42095), .Z(n40986) );
  NAND U42037 ( .A(n40987), .B(n40986), .Z(n41039) );
  NANDN U42038 ( .A(n40988), .B(n42231), .Z(n40990) );
  XOR U42039 ( .A(n244), .B(a[992]), .Z(n41029) );
  NANDN U42040 ( .A(n41029), .B(n42234), .Z(n40989) );
  AND U42041 ( .A(n40990), .B(n40989), .Z(n41038) );
  XNOR U42042 ( .A(n41039), .B(n41038), .Z(n41040) );
  XNOR U42043 ( .A(n41041), .B(n41040), .Z(n41045) );
  NANDN U42044 ( .A(n40992), .B(n40991), .Z(n40996) );
  NAND U42045 ( .A(n40994), .B(n40993), .Z(n40995) );
  AND U42046 ( .A(n40996), .B(n40995), .Z(n41044) );
  XOR U42047 ( .A(n41045), .B(n41044), .Z(n41046) );
  NANDN U42048 ( .A(n40998), .B(n40997), .Z(n41002) );
  NANDN U42049 ( .A(n41000), .B(n40999), .Z(n41001) );
  NAND U42050 ( .A(n41002), .B(n41001), .Z(n41047) );
  XOR U42051 ( .A(n41046), .B(n41047), .Z(n41014) );
  OR U42052 ( .A(n41004), .B(n41003), .Z(n41008) );
  NANDN U42053 ( .A(n41006), .B(n41005), .Z(n41007) );
  NAND U42054 ( .A(n41008), .B(n41007), .Z(n41015) );
  XNOR U42055 ( .A(n41014), .B(n41015), .Z(n41016) );
  XNOR U42056 ( .A(n41017), .B(n41016), .Z(n41050) );
  XNOR U42057 ( .A(n41050), .B(sreg[2014]), .Z(n41052) );
  NAND U42058 ( .A(n41009), .B(sreg[2013]), .Z(n41013) );
  OR U42059 ( .A(n41011), .B(n41010), .Z(n41012) );
  AND U42060 ( .A(n41013), .B(n41012), .Z(n41051) );
  XOR U42061 ( .A(n41052), .B(n41051), .Z(c[2014]) );
  NANDN U42062 ( .A(n41015), .B(n41014), .Z(n41019) );
  NAND U42063 ( .A(n41017), .B(n41016), .Z(n41018) );
  NAND U42064 ( .A(n41019), .B(n41018), .Z(n41058) );
  NAND U42065 ( .A(b[0]), .B(a[999]), .Z(n41020) );
  XNOR U42066 ( .A(b[1]), .B(n41020), .Z(n41022) );
  NAND U42067 ( .A(n157), .B(a[998]), .Z(n41021) );
  AND U42068 ( .A(n41022), .B(n41021), .Z(n41075) );
  XOR U42069 ( .A(a[995]), .B(n42197), .Z(n41064) );
  NANDN U42070 ( .A(n41064), .B(n42173), .Z(n41025) );
  NANDN U42071 ( .A(n41023), .B(n42172), .Z(n41024) );
  NAND U42072 ( .A(n41025), .B(n41024), .Z(n41073) );
  NAND U42073 ( .A(b[7]), .B(a[991]), .Z(n41074) );
  XNOR U42074 ( .A(n41073), .B(n41074), .Z(n41076) );
  XOR U42075 ( .A(n41075), .B(n41076), .Z(n41082) );
  NANDN U42076 ( .A(n41026), .B(n42093), .Z(n41028) );
  XOR U42077 ( .A(n42134), .B(a[997]), .Z(n41067) );
  NANDN U42078 ( .A(n41067), .B(n42095), .Z(n41027) );
  NAND U42079 ( .A(n41028), .B(n41027), .Z(n41080) );
  NANDN U42080 ( .A(n41029), .B(n42231), .Z(n41031) );
  XOR U42081 ( .A(n244), .B(a[993]), .Z(n41070) );
  NANDN U42082 ( .A(n41070), .B(n42234), .Z(n41030) );
  AND U42083 ( .A(n41031), .B(n41030), .Z(n41079) );
  XNOR U42084 ( .A(n41080), .B(n41079), .Z(n41081) );
  XNOR U42085 ( .A(n41082), .B(n41081), .Z(n41086) );
  NANDN U42086 ( .A(n41033), .B(n41032), .Z(n41037) );
  NAND U42087 ( .A(n41035), .B(n41034), .Z(n41036) );
  AND U42088 ( .A(n41037), .B(n41036), .Z(n41085) );
  XOR U42089 ( .A(n41086), .B(n41085), .Z(n41087) );
  NANDN U42090 ( .A(n41039), .B(n41038), .Z(n41043) );
  NANDN U42091 ( .A(n41041), .B(n41040), .Z(n41042) );
  NAND U42092 ( .A(n41043), .B(n41042), .Z(n41088) );
  XOR U42093 ( .A(n41087), .B(n41088), .Z(n41055) );
  OR U42094 ( .A(n41045), .B(n41044), .Z(n41049) );
  NANDN U42095 ( .A(n41047), .B(n41046), .Z(n41048) );
  NAND U42096 ( .A(n41049), .B(n41048), .Z(n41056) );
  XNOR U42097 ( .A(n41055), .B(n41056), .Z(n41057) );
  XNOR U42098 ( .A(n41058), .B(n41057), .Z(n41091) );
  XNOR U42099 ( .A(n41091), .B(sreg[2015]), .Z(n41093) );
  NAND U42100 ( .A(n41050), .B(sreg[2014]), .Z(n41054) );
  OR U42101 ( .A(n41052), .B(n41051), .Z(n41053) );
  AND U42102 ( .A(n41054), .B(n41053), .Z(n41092) );
  XOR U42103 ( .A(n41093), .B(n41092), .Z(c[2015]) );
  NANDN U42104 ( .A(n41056), .B(n41055), .Z(n41060) );
  NAND U42105 ( .A(n41058), .B(n41057), .Z(n41059) );
  NAND U42106 ( .A(n41060), .B(n41059), .Z(n41099) );
  NAND U42107 ( .A(b[0]), .B(a[1000]), .Z(n41061) );
  XNOR U42108 ( .A(b[1]), .B(n41061), .Z(n41063) );
  NAND U42109 ( .A(n157), .B(a[999]), .Z(n41062) );
  AND U42110 ( .A(n41063), .B(n41062), .Z(n41116) );
  XOR U42111 ( .A(a[996]), .B(n42197), .Z(n41105) );
  NANDN U42112 ( .A(n41105), .B(n42173), .Z(n41066) );
  NANDN U42113 ( .A(n41064), .B(n42172), .Z(n41065) );
  NAND U42114 ( .A(n41066), .B(n41065), .Z(n41114) );
  NAND U42115 ( .A(b[7]), .B(a[992]), .Z(n41115) );
  XNOR U42116 ( .A(n41114), .B(n41115), .Z(n41117) );
  XOR U42117 ( .A(n41116), .B(n41117), .Z(n41123) );
  NANDN U42118 ( .A(n41067), .B(n42093), .Z(n41069) );
  XOR U42119 ( .A(n42134), .B(a[998]), .Z(n41108) );
  NANDN U42120 ( .A(n41108), .B(n42095), .Z(n41068) );
  NAND U42121 ( .A(n41069), .B(n41068), .Z(n41121) );
  NANDN U42122 ( .A(n41070), .B(n42231), .Z(n41072) );
  XOR U42123 ( .A(n244), .B(a[994]), .Z(n41111) );
  NANDN U42124 ( .A(n41111), .B(n42234), .Z(n41071) );
  AND U42125 ( .A(n41072), .B(n41071), .Z(n41120) );
  XNOR U42126 ( .A(n41121), .B(n41120), .Z(n41122) );
  XNOR U42127 ( .A(n41123), .B(n41122), .Z(n41127) );
  NANDN U42128 ( .A(n41074), .B(n41073), .Z(n41078) );
  NAND U42129 ( .A(n41076), .B(n41075), .Z(n41077) );
  AND U42130 ( .A(n41078), .B(n41077), .Z(n41126) );
  XOR U42131 ( .A(n41127), .B(n41126), .Z(n41128) );
  NANDN U42132 ( .A(n41080), .B(n41079), .Z(n41084) );
  NANDN U42133 ( .A(n41082), .B(n41081), .Z(n41083) );
  NAND U42134 ( .A(n41084), .B(n41083), .Z(n41129) );
  XOR U42135 ( .A(n41128), .B(n41129), .Z(n41096) );
  OR U42136 ( .A(n41086), .B(n41085), .Z(n41090) );
  NANDN U42137 ( .A(n41088), .B(n41087), .Z(n41089) );
  NAND U42138 ( .A(n41090), .B(n41089), .Z(n41097) );
  XNOR U42139 ( .A(n41096), .B(n41097), .Z(n41098) );
  XNOR U42140 ( .A(n41099), .B(n41098), .Z(n41132) );
  XNOR U42141 ( .A(n41132), .B(sreg[2016]), .Z(n41134) );
  NAND U42142 ( .A(n41091), .B(sreg[2015]), .Z(n41095) );
  OR U42143 ( .A(n41093), .B(n41092), .Z(n41094) );
  AND U42144 ( .A(n41095), .B(n41094), .Z(n41133) );
  XOR U42145 ( .A(n41134), .B(n41133), .Z(c[2016]) );
  NANDN U42146 ( .A(n41097), .B(n41096), .Z(n41101) );
  NAND U42147 ( .A(n41099), .B(n41098), .Z(n41100) );
  NAND U42148 ( .A(n41101), .B(n41100), .Z(n41140) );
  NAND U42149 ( .A(b[0]), .B(a[1001]), .Z(n41102) );
  XNOR U42150 ( .A(b[1]), .B(n41102), .Z(n41104) );
  NAND U42151 ( .A(n158), .B(a[1000]), .Z(n41103) );
  AND U42152 ( .A(n41104), .B(n41103), .Z(n41157) );
  XOR U42153 ( .A(a[997]), .B(n42197), .Z(n41146) );
  NANDN U42154 ( .A(n41146), .B(n42173), .Z(n41107) );
  NANDN U42155 ( .A(n41105), .B(n42172), .Z(n41106) );
  NAND U42156 ( .A(n41107), .B(n41106), .Z(n41155) );
  NAND U42157 ( .A(b[7]), .B(a[993]), .Z(n41156) );
  XNOR U42158 ( .A(n41155), .B(n41156), .Z(n41158) );
  XOR U42159 ( .A(n41157), .B(n41158), .Z(n41164) );
  NANDN U42160 ( .A(n41108), .B(n42093), .Z(n41110) );
  XOR U42161 ( .A(n42134), .B(a[999]), .Z(n41149) );
  NANDN U42162 ( .A(n41149), .B(n42095), .Z(n41109) );
  NAND U42163 ( .A(n41110), .B(n41109), .Z(n41162) );
  NANDN U42164 ( .A(n41111), .B(n42231), .Z(n41113) );
  XOR U42165 ( .A(n245), .B(a[995]), .Z(n41152) );
  NANDN U42166 ( .A(n41152), .B(n42234), .Z(n41112) );
  AND U42167 ( .A(n41113), .B(n41112), .Z(n41161) );
  XNOR U42168 ( .A(n41162), .B(n41161), .Z(n41163) );
  XNOR U42169 ( .A(n41164), .B(n41163), .Z(n41168) );
  NANDN U42170 ( .A(n41115), .B(n41114), .Z(n41119) );
  NAND U42171 ( .A(n41117), .B(n41116), .Z(n41118) );
  AND U42172 ( .A(n41119), .B(n41118), .Z(n41167) );
  XOR U42173 ( .A(n41168), .B(n41167), .Z(n41169) );
  NANDN U42174 ( .A(n41121), .B(n41120), .Z(n41125) );
  NANDN U42175 ( .A(n41123), .B(n41122), .Z(n41124) );
  NAND U42176 ( .A(n41125), .B(n41124), .Z(n41170) );
  XOR U42177 ( .A(n41169), .B(n41170), .Z(n41137) );
  OR U42178 ( .A(n41127), .B(n41126), .Z(n41131) );
  NANDN U42179 ( .A(n41129), .B(n41128), .Z(n41130) );
  NAND U42180 ( .A(n41131), .B(n41130), .Z(n41138) );
  XNOR U42181 ( .A(n41137), .B(n41138), .Z(n41139) );
  XNOR U42182 ( .A(n41140), .B(n41139), .Z(n41173) );
  XNOR U42183 ( .A(n41173), .B(sreg[2017]), .Z(n41175) );
  NAND U42184 ( .A(n41132), .B(sreg[2016]), .Z(n41136) );
  OR U42185 ( .A(n41134), .B(n41133), .Z(n41135) );
  AND U42186 ( .A(n41136), .B(n41135), .Z(n41174) );
  XOR U42187 ( .A(n41175), .B(n41174), .Z(c[2017]) );
  NANDN U42188 ( .A(n41138), .B(n41137), .Z(n41142) );
  NAND U42189 ( .A(n41140), .B(n41139), .Z(n41141) );
  NAND U42190 ( .A(n41142), .B(n41141), .Z(n41181) );
  NAND U42191 ( .A(b[0]), .B(a[1002]), .Z(n41143) );
  XNOR U42192 ( .A(b[1]), .B(n41143), .Z(n41145) );
  NAND U42193 ( .A(n158), .B(a[1001]), .Z(n41144) );
  AND U42194 ( .A(n41145), .B(n41144), .Z(n41198) );
  XOR U42195 ( .A(a[998]), .B(n42197), .Z(n41187) );
  NANDN U42196 ( .A(n41187), .B(n42173), .Z(n41148) );
  NANDN U42197 ( .A(n41146), .B(n42172), .Z(n41147) );
  NAND U42198 ( .A(n41148), .B(n41147), .Z(n41196) );
  NAND U42199 ( .A(b[7]), .B(a[994]), .Z(n41197) );
  XNOR U42200 ( .A(n41196), .B(n41197), .Z(n41199) );
  XOR U42201 ( .A(n41198), .B(n41199), .Z(n41205) );
  NANDN U42202 ( .A(n41149), .B(n42093), .Z(n41151) );
  XOR U42203 ( .A(n42134), .B(a[1000]), .Z(n41190) );
  NANDN U42204 ( .A(n41190), .B(n42095), .Z(n41150) );
  NAND U42205 ( .A(n41151), .B(n41150), .Z(n41203) );
  NANDN U42206 ( .A(n41152), .B(n42231), .Z(n41154) );
  XOR U42207 ( .A(n245), .B(a[996]), .Z(n41193) );
  NANDN U42208 ( .A(n41193), .B(n42234), .Z(n41153) );
  AND U42209 ( .A(n41154), .B(n41153), .Z(n41202) );
  XNOR U42210 ( .A(n41203), .B(n41202), .Z(n41204) );
  XNOR U42211 ( .A(n41205), .B(n41204), .Z(n41209) );
  NANDN U42212 ( .A(n41156), .B(n41155), .Z(n41160) );
  NAND U42213 ( .A(n41158), .B(n41157), .Z(n41159) );
  AND U42214 ( .A(n41160), .B(n41159), .Z(n41208) );
  XOR U42215 ( .A(n41209), .B(n41208), .Z(n41210) );
  NANDN U42216 ( .A(n41162), .B(n41161), .Z(n41166) );
  NANDN U42217 ( .A(n41164), .B(n41163), .Z(n41165) );
  NAND U42218 ( .A(n41166), .B(n41165), .Z(n41211) );
  XOR U42219 ( .A(n41210), .B(n41211), .Z(n41178) );
  OR U42220 ( .A(n41168), .B(n41167), .Z(n41172) );
  NANDN U42221 ( .A(n41170), .B(n41169), .Z(n41171) );
  NAND U42222 ( .A(n41172), .B(n41171), .Z(n41179) );
  XNOR U42223 ( .A(n41178), .B(n41179), .Z(n41180) );
  XNOR U42224 ( .A(n41181), .B(n41180), .Z(n41214) );
  XNOR U42225 ( .A(n41214), .B(sreg[2018]), .Z(n41216) );
  NAND U42226 ( .A(n41173), .B(sreg[2017]), .Z(n41177) );
  OR U42227 ( .A(n41175), .B(n41174), .Z(n41176) );
  AND U42228 ( .A(n41177), .B(n41176), .Z(n41215) );
  XOR U42229 ( .A(n41216), .B(n41215), .Z(c[2018]) );
  NANDN U42230 ( .A(n41179), .B(n41178), .Z(n41183) );
  NAND U42231 ( .A(n41181), .B(n41180), .Z(n41182) );
  NAND U42232 ( .A(n41183), .B(n41182), .Z(n41222) );
  NAND U42233 ( .A(b[0]), .B(a[1003]), .Z(n41184) );
  XNOR U42234 ( .A(b[1]), .B(n41184), .Z(n41186) );
  NAND U42235 ( .A(n158), .B(a[1002]), .Z(n41185) );
  AND U42236 ( .A(n41186), .B(n41185), .Z(n41239) );
  XOR U42237 ( .A(a[999]), .B(n42197), .Z(n41228) );
  NANDN U42238 ( .A(n41228), .B(n42173), .Z(n41189) );
  NANDN U42239 ( .A(n41187), .B(n42172), .Z(n41188) );
  NAND U42240 ( .A(n41189), .B(n41188), .Z(n41237) );
  NAND U42241 ( .A(b[7]), .B(a[995]), .Z(n41238) );
  XNOR U42242 ( .A(n41237), .B(n41238), .Z(n41240) );
  XOR U42243 ( .A(n41239), .B(n41240), .Z(n41246) );
  NANDN U42244 ( .A(n41190), .B(n42093), .Z(n41192) );
  XOR U42245 ( .A(n42134), .B(a[1001]), .Z(n41231) );
  NANDN U42246 ( .A(n41231), .B(n42095), .Z(n41191) );
  NAND U42247 ( .A(n41192), .B(n41191), .Z(n41244) );
  NANDN U42248 ( .A(n41193), .B(n42231), .Z(n41195) );
  XOR U42249 ( .A(n245), .B(a[997]), .Z(n41234) );
  NANDN U42250 ( .A(n41234), .B(n42234), .Z(n41194) );
  AND U42251 ( .A(n41195), .B(n41194), .Z(n41243) );
  XNOR U42252 ( .A(n41244), .B(n41243), .Z(n41245) );
  XNOR U42253 ( .A(n41246), .B(n41245), .Z(n41250) );
  NANDN U42254 ( .A(n41197), .B(n41196), .Z(n41201) );
  NAND U42255 ( .A(n41199), .B(n41198), .Z(n41200) );
  AND U42256 ( .A(n41201), .B(n41200), .Z(n41249) );
  XOR U42257 ( .A(n41250), .B(n41249), .Z(n41251) );
  NANDN U42258 ( .A(n41203), .B(n41202), .Z(n41207) );
  NANDN U42259 ( .A(n41205), .B(n41204), .Z(n41206) );
  NAND U42260 ( .A(n41207), .B(n41206), .Z(n41252) );
  XOR U42261 ( .A(n41251), .B(n41252), .Z(n41219) );
  OR U42262 ( .A(n41209), .B(n41208), .Z(n41213) );
  NANDN U42263 ( .A(n41211), .B(n41210), .Z(n41212) );
  NAND U42264 ( .A(n41213), .B(n41212), .Z(n41220) );
  XNOR U42265 ( .A(n41219), .B(n41220), .Z(n41221) );
  XNOR U42266 ( .A(n41222), .B(n41221), .Z(n41255) );
  XNOR U42267 ( .A(n41255), .B(sreg[2019]), .Z(n41257) );
  NAND U42268 ( .A(n41214), .B(sreg[2018]), .Z(n41218) );
  OR U42269 ( .A(n41216), .B(n41215), .Z(n41217) );
  AND U42270 ( .A(n41218), .B(n41217), .Z(n41256) );
  XOR U42271 ( .A(n41257), .B(n41256), .Z(c[2019]) );
  NANDN U42272 ( .A(n41220), .B(n41219), .Z(n41224) );
  NAND U42273 ( .A(n41222), .B(n41221), .Z(n41223) );
  NAND U42274 ( .A(n41224), .B(n41223), .Z(n41263) );
  NAND U42275 ( .A(b[0]), .B(a[1004]), .Z(n41225) );
  XNOR U42276 ( .A(b[1]), .B(n41225), .Z(n41227) );
  NAND U42277 ( .A(n158), .B(a[1003]), .Z(n41226) );
  AND U42278 ( .A(n41227), .B(n41226), .Z(n41280) );
  XOR U42279 ( .A(a[1000]), .B(n42197), .Z(n41269) );
  NANDN U42280 ( .A(n41269), .B(n42173), .Z(n41230) );
  NANDN U42281 ( .A(n41228), .B(n42172), .Z(n41229) );
  NAND U42282 ( .A(n41230), .B(n41229), .Z(n41278) );
  NAND U42283 ( .A(b[7]), .B(a[996]), .Z(n41279) );
  XNOR U42284 ( .A(n41278), .B(n41279), .Z(n41281) );
  XOR U42285 ( .A(n41280), .B(n41281), .Z(n41287) );
  NANDN U42286 ( .A(n41231), .B(n42093), .Z(n41233) );
  XOR U42287 ( .A(n42134), .B(a[1002]), .Z(n41272) );
  NANDN U42288 ( .A(n41272), .B(n42095), .Z(n41232) );
  NAND U42289 ( .A(n41233), .B(n41232), .Z(n41285) );
  NANDN U42290 ( .A(n41234), .B(n42231), .Z(n41236) );
  XOR U42291 ( .A(n245), .B(a[998]), .Z(n41275) );
  NANDN U42292 ( .A(n41275), .B(n42234), .Z(n41235) );
  AND U42293 ( .A(n41236), .B(n41235), .Z(n41284) );
  XNOR U42294 ( .A(n41285), .B(n41284), .Z(n41286) );
  XNOR U42295 ( .A(n41287), .B(n41286), .Z(n41291) );
  NANDN U42296 ( .A(n41238), .B(n41237), .Z(n41242) );
  NAND U42297 ( .A(n41240), .B(n41239), .Z(n41241) );
  AND U42298 ( .A(n41242), .B(n41241), .Z(n41290) );
  XOR U42299 ( .A(n41291), .B(n41290), .Z(n41292) );
  NANDN U42300 ( .A(n41244), .B(n41243), .Z(n41248) );
  NANDN U42301 ( .A(n41246), .B(n41245), .Z(n41247) );
  NAND U42302 ( .A(n41248), .B(n41247), .Z(n41293) );
  XOR U42303 ( .A(n41292), .B(n41293), .Z(n41260) );
  OR U42304 ( .A(n41250), .B(n41249), .Z(n41254) );
  NANDN U42305 ( .A(n41252), .B(n41251), .Z(n41253) );
  NAND U42306 ( .A(n41254), .B(n41253), .Z(n41261) );
  XNOR U42307 ( .A(n41260), .B(n41261), .Z(n41262) );
  XNOR U42308 ( .A(n41263), .B(n41262), .Z(n41296) );
  XNOR U42309 ( .A(n41296), .B(sreg[2020]), .Z(n41298) );
  NAND U42310 ( .A(n41255), .B(sreg[2019]), .Z(n41259) );
  OR U42311 ( .A(n41257), .B(n41256), .Z(n41258) );
  AND U42312 ( .A(n41259), .B(n41258), .Z(n41297) );
  XOR U42313 ( .A(n41298), .B(n41297), .Z(c[2020]) );
  NANDN U42314 ( .A(n41261), .B(n41260), .Z(n41265) );
  NAND U42315 ( .A(n41263), .B(n41262), .Z(n41264) );
  NAND U42316 ( .A(n41265), .B(n41264), .Z(n41304) );
  NAND U42317 ( .A(b[0]), .B(a[1005]), .Z(n41266) );
  XNOR U42318 ( .A(b[1]), .B(n41266), .Z(n41268) );
  NAND U42319 ( .A(n158), .B(a[1004]), .Z(n41267) );
  AND U42320 ( .A(n41268), .B(n41267), .Z(n41321) );
  XOR U42321 ( .A(a[1001]), .B(n42197), .Z(n41310) );
  NANDN U42322 ( .A(n41310), .B(n42173), .Z(n41271) );
  NANDN U42323 ( .A(n41269), .B(n42172), .Z(n41270) );
  NAND U42324 ( .A(n41271), .B(n41270), .Z(n41319) );
  NAND U42325 ( .A(b[7]), .B(a[997]), .Z(n41320) );
  XNOR U42326 ( .A(n41319), .B(n41320), .Z(n41322) );
  XOR U42327 ( .A(n41321), .B(n41322), .Z(n41328) );
  NANDN U42328 ( .A(n41272), .B(n42093), .Z(n41274) );
  XOR U42329 ( .A(n42134), .B(a[1003]), .Z(n41313) );
  NANDN U42330 ( .A(n41313), .B(n42095), .Z(n41273) );
  NAND U42331 ( .A(n41274), .B(n41273), .Z(n41326) );
  NANDN U42332 ( .A(n41275), .B(n42231), .Z(n41277) );
  XOR U42333 ( .A(n245), .B(a[999]), .Z(n41316) );
  NANDN U42334 ( .A(n41316), .B(n42234), .Z(n41276) );
  AND U42335 ( .A(n41277), .B(n41276), .Z(n41325) );
  XNOR U42336 ( .A(n41326), .B(n41325), .Z(n41327) );
  XNOR U42337 ( .A(n41328), .B(n41327), .Z(n41332) );
  NANDN U42338 ( .A(n41279), .B(n41278), .Z(n41283) );
  NAND U42339 ( .A(n41281), .B(n41280), .Z(n41282) );
  AND U42340 ( .A(n41283), .B(n41282), .Z(n41331) );
  XOR U42341 ( .A(n41332), .B(n41331), .Z(n41333) );
  NANDN U42342 ( .A(n41285), .B(n41284), .Z(n41289) );
  NANDN U42343 ( .A(n41287), .B(n41286), .Z(n41288) );
  NAND U42344 ( .A(n41289), .B(n41288), .Z(n41334) );
  XOR U42345 ( .A(n41333), .B(n41334), .Z(n41301) );
  OR U42346 ( .A(n41291), .B(n41290), .Z(n41295) );
  NANDN U42347 ( .A(n41293), .B(n41292), .Z(n41294) );
  NAND U42348 ( .A(n41295), .B(n41294), .Z(n41302) );
  XNOR U42349 ( .A(n41301), .B(n41302), .Z(n41303) );
  XNOR U42350 ( .A(n41304), .B(n41303), .Z(n41337) );
  XNOR U42351 ( .A(n41337), .B(sreg[2021]), .Z(n41339) );
  NAND U42352 ( .A(n41296), .B(sreg[2020]), .Z(n41300) );
  OR U42353 ( .A(n41298), .B(n41297), .Z(n41299) );
  AND U42354 ( .A(n41300), .B(n41299), .Z(n41338) );
  XOR U42355 ( .A(n41339), .B(n41338), .Z(c[2021]) );
  NANDN U42356 ( .A(n41302), .B(n41301), .Z(n41306) );
  NAND U42357 ( .A(n41304), .B(n41303), .Z(n41305) );
  NAND U42358 ( .A(n41306), .B(n41305), .Z(n41345) );
  NAND U42359 ( .A(b[0]), .B(a[1006]), .Z(n41307) );
  XNOR U42360 ( .A(b[1]), .B(n41307), .Z(n41309) );
  NAND U42361 ( .A(n158), .B(a[1005]), .Z(n41308) );
  AND U42362 ( .A(n41309), .B(n41308), .Z(n41362) );
  XOR U42363 ( .A(a[1002]), .B(n42197), .Z(n41351) );
  NANDN U42364 ( .A(n41351), .B(n42173), .Z(n41312) );
  NANDN U42365 ( .A(n41310), .B(n42172), .Z(n41311) );
  NAND U42366 ( .A(n41312), .B(n41311), .Z(n41360) );
  NAND U42367 ( .A(b[7]), .B(a[998]), .Z(n41361) );
  XNOR U42368 ( .A(n41360), .B(n41361), .Z(n41363) );
  XOR U42369 ( .A(n41362), .B(n41363), .Z(n41369) );
  NANDN U42370 ( .A(n41313), .B(n42093), .Z(n41315) );
  XOR U42371 ( .A(n42134), .B(a[1004]), .Z(n41354) );
  NANDN U42372 ( .A(n41354), .B(n42095), .Z(n41314) );
  NAND U42373 ( .A(n41315), .B(n41314), .Z(n41367) );
  NANDN U42374 ( .A(n41316), .B(n42231), .Z(n41318) );
  XOR U42375 ( .A(n245), .B(a[1000]), .Z(n41357) );
  NANDN U42376 ( .A(n41357), .B(n42234), .Z(n41317) );
  AND U42377 ( .A(n41318), .B(n41317), .Z(n41366) );
  XNOR U42378 ( .A(n41367), .B(n41366), .Z(n41368) );
  XNOR U42379 ( .A(n41369), .B(n41368), .Z(n41373) );
  NANDN U42380 ( .A(n41320), .B(n41319), .Z(n41324) );
  NAND U42381 ( .A(n41322), .B(n41321), .Z(n41323) );
  AND U42382 ( .A(n41324), .B(n41323), .Z(n41372) );
  XOR U42383 ( .A(n41373), .B(n41372), .Z(n41374) );
  NANDN U42384 ( .A(n41326), .B(n41325), .Z(n41330) );
  NANDN U42385 ( .A(n41328), .B(n41327), .Z(n41329) );
  NAND U42386 ( .A(n41330), .B(n41329), .Z(n41375) );
  XOR U42387 ( .A(n41374), .B(n41375), .Z(n41342) );
  OR U42388 ( .A(n41332), .B(n41331), .Z(n41336) );
  NANDN U42389 ( .A(n41334), .B(n41333), .Z(n41335) );
  NAND U42390 ( .A(n41336), .B(n41335), .Z(n41343) );
  XNOR U42391 ( .A(n41342), .B(n41343), .Z(n41344) );
  XNOR U42392 ( .A(n41345), .B(n41344), .Z(n41378) );
  XNOR U42393 ( .A(n41378), .B(sreg[2022]), .Z(n41380) );
  NAND U42394 ( .A(n41337), .B(sreg[2021]), .Z(n41341) );
  OR U42395 ( .A(n41339), .B(n41338), .Z(n41340) );
  AND U42396 ( .A(n41341), .B(n41340), .Z(n41379) );
  XOR U42397 ( .A(n41380), .B(n41379), .Z(c[2022]) );
  NANDN U42398 ( .A(n41343), .B(n41342), .Z(n41347) );
  NAND U42399 ( .A(n41345), .B(n41344), .Z(n41346) );
  NAND U42400 ( .A(n41347), .B(n41346), .Z(n41386) );
  NAND U42401 ( .A(b[0]), .B(a[1007]), .Z(n41348) );
  XNOR U42402 ( .A(b[1]), .B(n41348), .Z(n41350) );
  NAND U42403 ( .A(n158), .B(a[1006]), .Z(n41349) );
  AND U42404 ( .A(n41350), .B(n41349), .Z(n41403) );
  XOR U42405 ( .A(a[1003]), .B(n42197), .Z(n41392) );
  NANDN U42406 ( .A(n41392), .B(n42173), .Z(n41353) );
  NANDN U42407 ( .A(n41351), .B(n42172), .Z(n41352) );
  NAND U42408 ( .A(n41353), .B(n41352), .Z(n41401) );
  NAND U42409 ( .A(b[7]), .B(a[999]), .Z(n41402) );
  XNOR U42410 ( .A(n41401), .B(n41402), .Z(n41404) );
  XOR U42411 ( .A(n41403), .B(n41404), .Z(n41410) );
  NANDN U42412 ( .A(n41354), .B(n42093), .Z(n41356) );
  XOR U42413 ( .A(n42134), .B(a[1005]), .Z(n41395) );
  NANDN U42414 ( .A(n41395), .B(n42095), .Z(n41355) );
  NAND U42415 ( .A(n41356), .B(n41355), .Z(n41408) );
  NANDN U42416 ( .A(n41357), .B(n42231), .Z(n41359) );
  XOR U42417 ( .A(n245), .B(a[1001]), .Z(n41398) );
  NANDN U42418 ( .A(n41398), .B(n42234), .Z(n41358) );
  AND U42419 ( .A(n41359), .B(n41358), .Z(n41407) );
  XNOR U42420 ( .A(n41408), .B(n41407), .Z(n41409) );
  XNOR U42421 ( .A(n41410), .B(n41409), .Z(n41414) );
  NANDN U42422 ( .A(n41361), .B(n41360), .Z(n41365) );
  NAND U42423 ( .A(n41363), .B(n41362), .Z(n41364) );
  AND U42424 ( .A(n41365), .B(n41364), .Z(n41413) );
  XOR U42425 ( .A(n41414), .B(n41413), .Z(n41415) );
  NANDN U42426 ( .A(n41367), .B(n41366), .Z(n41371) );
  NANDN U42427 ( .A(n41369), .B(n41368), .Z(n41370) );
  NAND U42428 ( .A(n41371), .B(n41370), .Z(n41416) );
  XOR U42429 ( .A(n41415), .B(n41416), .Z(n41383) );
  OR U42430 ( .A(n41373), .B(n41372), .Z(n41377) );
  NANDN U42431 ( .A(n41375), .B(n41374), .Z(n41376) );
  NAND U42432 ( .A(n41377), .B(n41376), .Z(n41384) );
  XNOR U42433 ( .A(n41383), .B(n41384), .Z(n41385) );
  XNOR U42434 ( .A(n41386), .B(n41385), .Z(n41419) );
  XNOR U42435 ( .A(n41419), .B(sreg[2023]), .Z(n41421) );
  NAND U42436 ( .A(n41378), .B(sreg[2022]), .Z(n41382) );
  OR U42437 ( .A(n41380), .B(n41379), .Z(n41381) );
  AND U42438 ( .A(n41382), .B(n41381), .Z(n41420) );
  XOR U42439 ( .A(n41421), .B(n41420), .Z(c[2023]) );
  NANDN U42440 ( .A(n41384), .B(n41383), .Z(n41388) );
  NAND U42441 ( .A(n41386), .B(n41385), .Z(n41387) );
  NAND U42442 ( .A(n41388), .B(n41387), .Z(n41427) );
  NAND U42443 ( .A(b[0]), .B(a[1008]), .Z(n41389) );
  XNOR U42444 ( .A(b[1]), .B(n41389), .Z(n41391) );
  NAND U42445 ( .A(n159), .B(a[1007]), .Z(n41390) );
  AND U42446 ( .A(n41391), .B(n41390), .Z(n41444) );
  XOR U42447 ( .A(a[1004]), .B(n42197), .Z(n41433) );
  NANDN U42448 ( .A(n41433), .B(n42173), .Z(n41394) );
  NANDN U42449 ( .A(n41392), .B(n42172), .Z(n41393) );
  NAND U42450 ( .A(n41394), .B(n41393), .Z(n41442) );
  NAND U42451 ( .A(b[7]), .B(a[1000]), .Z(n41443) );
  XNOR U42452 ( .A(n41442), .B(n41443), .Z(n41445) );
  XOR U42453 ( .A(n41444), .B(n41445), .Z(n41451) );
  NANDN U42454 ( .A(n41395), .B(n42093), .Z(n41397) );
  XOR U42455 ( .A(n42134), .B(a[1006]), .Z(n41436) );
  NANDN U42456 ( .A(n41436), .B(n42095), .Z(n41396) );
  NAND U42457 ( .A(n41397), .B(n41396), .Z(n41449) );
  NANDN U42458 ( .A(n41398), .B(n42231), .Z(n41400) );
  XOR U42459 ( .A(n245), .B(a[1002]), .Z(n41439) );
  NANDN U42460 ( .A(n41439), .B(n42234), .Z(n41399) );
  AND U42461 ( .A(n41400), .B(n41399), .Z(n41448) );
  XNOR U42462 ( .A(n41449), .B(n41448), .Z(n41450) );
  XNOR U42463 ( .A(n41451), .B(n41450), .Z(n41455) );
  NANDN U42464 ( .A(n41402), .B(n41401), .Z(n41406) );
  NAND U42465 ( .A(n41404), .B(n41403), .Z(n41405) );
  AND U42466 ( .A(n41406), .B(n41405), .Z(n41454) );
  XOR U42467 ( .A(n41455), .B(n41454), .Z(n41456) );
  NANDN U42468 ( .A(n41408), .B(n41407), .Z(n41412) );
  NANDN U42469 ( .A(n41410), .B(n41409), .Z(n41411) );
  NAND U42470 ( .A(n41412), .B(n41411), .Z(n41457) );
  XOR U42471 ( .A(n41456), .B(n41457), .Z(n41424) );
  OR U42472 ( .A(n41414), .B(n41413), .Z(n41418) );
  NANDN U42473 ( .A(n41416), .B(n41415), .Z(n41417) );
  NAND U42474 ( .A(n41418), .B(n41417), .Z(n41425) );
  XNOR U42475 ( .A(n41424), .B(n41425), .Z(n41426) );
  XNOR U42476 ( .A(n41427), .B(n41426), .Z(n41460) );
  XNOR U42477 ( .A(n41460), .B(sreg[2024]), .Z(n41462) );
  NAND U42478 ( .A(n41419), .B(sreg[2023]), .Z(n41423) );
  OR U42479 ( .A(n41421), .B(n41420), .Z(n41422) );
  AND U42480 ( .A(n41423), .B(n41422), .Z(n41461) );
  XOR U42481 ( .A(n41462), .B(n41461), .Z(c[2024]) );
  NANDN U42482 ( .A(n41425), .B(n41424), .Z(n41429) );
  NAND U42483 ( .A(n41427), .B(n41426), .Z(n41428) );
  NAND U42484 ( .A(n41429), .B(n41428), .Z(n41468) );
  NAND U42485 ( .A(b[0]), .B(a[1009]), .Z(n41430) );
  XNOR U42486 ( .A(b[1]), .B(n41430), .Z(n41432) );
  NAND U42487 ( .A(n159), .B(a[1008]), .Z(n41431) );
  AND U42488 ( .A(n41432), .B(n41431), .Z(n41485) );
  XOR U42489 ( .A(a[1005]), .B(n42197), .Z(n41474) );
  NANDN U42490 ( .A(n41474), .B(n42173), .Z(n41435) );
  NANDN U42491 ( .A(n41433), .B(n42172), .Z(n41434) );
  NAND U42492 ( .A(n41435), .B(n41434), .Z(n41483) );
  NAND U42493 ( .A(b[7]), .B(a[1001]), .Z(n41484) );
  XNOR U42494 ( .A(n41483), .B(n41484), .Z(n41486) );
  XOR U42495 ( .A(n41485), .B(n41486), .Z(n41492) );
  NANDN U42496 ( .A(n41436), .B(n42093), .Z(n41438) );
  XOR U42497 ( .A(n42134), .B(a[1007]), .Z(n41477) );
  NANDN U42498 ( .A(n41477), .B(n42095), .Z(n41437) );
  NAND U42499 ( .A(n41438), .B(n41437), .Z(n41490) );
  NANDN U42500 ( .A(n41439), .B(n42231), .Z(n41441) );
  XOR U42501 ( .A(n245), .B(a[1003]), .Z(n41480) );
  NANDN U42502 ( .A(n41480), .B(n42234), .Z(n41440) );
  AND U42503 ( .A(n41441), .B(n41440), .Z(n41489) );
  XNOR U42504 ( .A(n41490), .B(n41489), .Z(n41491) );
  XNOR U42505 ( .A(n41492), .B(n41491), .Z(n41496) );
  NANDN U42506 ( .A(n41443), .B(n41442), .Z(n41447) );
  NAND U42507 ( .A(n41445), .B(n41444), .Z(n41446) );
  AND U42508 ( .A(n41447), .B(n41446), .Z(n41495) );
  XOR U42509 ( .A(n41496), .B(n41495), .Z(n41497) );
  NANDN U42510 ( .A(n41449), .B(n41448), .Z(n41453) );
  NANDN U42511 ( .A(n41451), .B(n41450), .Z(n41452) );
  NAND U42512 ( .A(n41453), .B(n41452), .Z(n41498) );
  XOR U42513 ( .A(n41497), .B(n41498), .Z(n41465) );
  OR U42514 ( .A(n41455), .B(n41454), .Z(n41459) );
  NANDN U42515 ( .A(n41457), .B(n41456), .Z(n41458) );
  NAND U42516 ( .A(n41459), .B(n41458), .Z(n41466) );
  XNOR U42517 ( .A(n41465), .B(n41466), .Z(n41467) );
  XNOR U42518 ( .A(n41468), .B(n41467), .Z(n41501) );
  XNOR U42519 ( .A(n41501), .B(sreg[2025]), .Z(n41503) );
  NAND U42520 ( .A(n41460), .B(sreg[2024]), .Z(n41464) );
  OR U42521 ( .A(n41462), .B(n41461), .Z(n41463) );
  AND U42522 ( .A(n41464), .B(n41463), .Z(n41502) );
  XOR U42523 ( .A(n41503), .B(n41502), .Z(c[2025]) );
  NANDN U42524 ( .A(n41466), .B(n41465), .Z(n41470) );
  NAND U42525 ( .A(n41468), .B(n41467), .Z(n41469) );
  NAND U42526 ( .A(n41470), .B(n41469), .Z(n41509) );
  NAND U42527 ( .A(b[0]), .B(a[1010]), .Z(n41471) );
  XNOR U42528 ( .A(b[1]), .B(n41471), .Z(n41473) );
  NAND U42529 ( .A(n159), .B(a[1009]), .Z(n41472) );
  AND U42530 ( .A(n41473), .B(n41472), .Z(n41526) );
  XOR U42531 ( .A(a[1006]), .B(n42197), .Z(n41515) );
  NANDN U42532 ( .A(n41515), .B(n42173), .Z(n41476) );
  NANDN U42533 ( .A(n41474), .B(n42172), .Z(n41475) );
  NAND U42534 ( .A(n41476), .B(n41475), .Z(n41524) );
  NAND U42535 ( .A(b[7]), .B(a[1002]), .Z(n41525) );
  XNOR U42536 ( .A(n41524), .B(n41525), .Z(n41527) );
  XOR U42537 ( .A(n41526), .B(n41527), .Z(n41533) );
  NANDN U42538 ( .A(n41477), .B(n42093), .Z(n41479) );
  XOR U42539 ( .A(n42134), .B(a[1008]), .Z(n41518) );
  NANDN U42540 ( .A(n41518), .B(n42095), .Z(n41478) );
  NAND U42541 ( .A(n41479), .B(n41478), .Z(n41531) );
  NANDN U42542 ( .A(n41480), .B(n42231), .Z(n41482) );
  XOR U42543 ( .A(n245), .B(a[1004]), .Z(n41521) );
  NANDN U42544 ( .A(n41521), .B(n42234), .Z(n41481) );
  AND U42545 ( .A(n41482), .B(n41481), .Z(n41530) );
  XNOR U42546 ( .A(n41531), .B(n41530), .Z(n41532) );
  XNOR U42547 ( .A(n41533), .B(n41532), .Z(n41537) );
  NANDN U42548 ( .A(n41484), .B(n41483), .Z(n41488) );
  NAND U42549 ( .A(n41486), .B(n41485), .Z(n41487) );
  AND U42550 ( .A(n41488), .B(n41487), .Z(n41536) );
  XOR U42551 ( .A(n41537), .B(n41536), .Z(n41538) );
  NANDN U42552 ( .A(n41490), .B(n41489), .Z(n41494) );
  NANDN U42553 ( .A(n41492), .B(n41491), .Z(n41493) );
  NAND U42554 ( .A(n41494), .B(n41493), .Z(n41539) );
  XOR U42555 ( .A(n41538), .B(n41539), .Z(n41506) );
  OR U42556 ( .A(n41496), .B(n41495), .Z(n41500) );
  NANDN U42557 ( .A(n41498), .B(n41497), .Z(n41499) );
  NAND U42558 ( .A(n41500), .B(n41499), .Z(n41507) );
  XNOR U42559 ( .A(n41506), .B(n41507), .Z(n41508) );
  XNOR U42560 ( .A(n41509), .B(n41508), .Z(n41542) );
  XNOR U42561 ( .A(n41542), .B(sreg[2026]), .Z(n41544) );
  NAND U42562 ( .A(n41501), .B(sreg[2025]), .Z(n41505) );
  OR U42563 ( .A(n41503), .B(n41502), .Z(n41504) );
  AND U42564 ( .A(n41505), .B(n41504), .Z(n41543) );
  XOR U42565 ( .A(n41544), .B(n41543), .Z(c[2026]) );
  NANDN U42566 ( .A(n41507), .B(n41506), .Z(n41511) );
  NAND U42567 ( .A(n41509), .B(n41508), .Z(n41510) );
  NAND U42568 ( .A(n41511), .B(n41510), .Z(n41550) );
  NAND U42569 ( .A(b[0]), .B(a[1011]), .Z(n41512) );
  XNOR U42570 ( .A(b[1]), .B(n41512), .Z(n41514) );
  NAND U42571 ( .A(n159), .B(a[1010]), .Z(n41513) );
  AND U42572 ( .A(n41514), .B(n41513), .Z(n41567) );
  XOR U42573 ( .A(a[1007]), .B(n42197), .Z(n41556) );
  NANDN U42574 ( .A(n41556), .B(n42173), .Z(n41517) );
  NANDN U42575 ( .A(n41515), .B(n42172), .Z(n41516) );
  NAND U42576 ( .A(n41517), .B(n41516), .Z(n41565) );
  NAND U42577 ( .A(b[7]), .B(a[1003]), .Z(n41566) );
  XNOR U42578 ( .A(n41565), .B(n41566), .Z(n41568) );
  XOR U42579 ( .A(n41567), .B(n41568), .Z(n41574) );
  NANDN U42580 ( .A(n41518), .B(n42093), .Z(n41520) );
  XOR U42581 ( .A(n42134), .B(a[1009]), .Z(n41559) );
  NANDN U42582 ( .A(n41559), .B(n42095), .Z(n41519) );
  NAND U42583 ( .A(n41520), .B(n41519), .Z(n41572) );
  NANDN U42584 ( .A(n41521), .B(n42231), .Z(n41523) );
  XOR U42585 ( .A(n245), .B(a[1005]), .Z(n41562) );
  NANDN U42586 ( .A(n41562), .B(n42234), .Z(n41522) );
  AND U42587 ( .A(n41523), .B(n41522), .Z(n41571) );
  XNOR U42588 ( .A(n41572), .B(n41571), .Z(n41573) );
  XNOR U42589 ( .A(n41574), .B(n41573), .Z(n41578) );
  NANDN U42590 ( .A(n41525), .B(n41524), .Z(n41529) );
  NAND U42591 ( .A(n41527), .B(n41526), .Z(n41528) );
  AND U42592 ( .A(n41529), .B(n41528), .Z(n41577) );
  XOR U42593 ( .A(n41578), .B(n41577), .Z(n41579) );
  NANDN U42594 ( .A(n41531), .B(n41530), .Z(n41535) );
  NANDN U42595 ( .A(n41533), .B(n41532), .Z(n41534) );
  NAND U42596 ( .A(n41535), .B(n41534), .Z(n41580) );
  XOR U42597 ( .A(n41579), .B(n41580), .Z(n41547) );
  OR U42598 ( .A(n41537), .B(n41536), .Z(n41541) );
  NANDN U42599 ( .A(n41539), .B(n41538), .Z(n41540) );
  NAND U42600 ( .A(n41541), .B(n41540), .Z(n41548) );
  XNOR U42601 ( .A(n41547), .B(n41548), .Z(n41549) );
  XNOR U42602 ( .A(n41550), .B(n41549), .Z(n41583) );
  XNOR U42603 ( .A(n41583), .B(sreg[2027]), .Z(n41585) );
  NAND U42604 ( .A(n41542), .B(sreg[2026]), .Z(n41546) );
  OR U42605 ( .A(n41544), .B(n41543), .Z(n41545) );
  AND U42606 ( .A(n41546), .B(n41545), .Z(n41584) );
  XOR U42607 ( .A(n41585), .B(n41584), .Z(c[2027]) );
  NANDN U42608 ( .A(n41548), .B(n41547), .Z(n41552) );
  NAND U42609 ( .A(n41550), .B(n41549), .Z(n41551) );
  NAND U42610 ( .A(n41552), .B(n41551), .Z(n41591) );
  NAND U42611 ( .A(b[0]), .B(a[1012]), .Z(n41553) );
  XNOR U42612 ( .A(b[1]), .B(n41553), .Z(n41555) );
  NAND U42613 ( .A(n159), .B(a[1011]), .Z(n41554) );
  AND U42614 ( .A(n41555), .B(n41554), .Z(n41608) );
  XOR U42615 ( .A(a[1008]), .B(n42197), .Z(n41597) );
  NANDN U42616 ( .A(n41597), .B(n42173), .Z(n41558) );
  NANDN U42617 ( .A(n41556), .B(n42172), .Z(n41557) );
  NAND U42618 ( .A(n41558), .B(n41557), .Z(n41606) );
  NAND U42619 ( .A(b[7]), .B(a[1004]), .Z(n41607) );
  XNOR U42620 ( .A(n41606), .B(n41607), .Z(n41609) );
  XOR U42621 ( .A(n41608), .B(n41609), .Z(n41615) );
  NANDN U42622 ( .A(n41559), .B(n42093), .Z(n41561) );
  XOR U42623 ( .A(n42134), .B(a[1010]), .Z(n41600) );
  NANDN U42624 ( .A(n41600), .B(n42095), .Z(n41560) );
  NAND U42625 ( .A(n41561), .B(n41560), .Z(n41613) );
  NANDN U42626 ( .A(n41562), .B(n42231), .Z(n41564) );
  XOR U42627 ( .A(n245), .B(a[1006]), .Z(n41603) );
  NANDN U42628 ( .A(n41603), .B(n42234), .Z(n41563) );
  AND U42629 ( .A(n41564), .B(n41563), .Z(n41612) );
  XNOR U42630 ( .A(n41613), .B(n41612), .Z(n41614) );
  XNOR U42631 ( .A(n41615), .B(n41614), .Z(n41619) );
  NANDN U42632 ( .A(n41566), .B(n41565), .Z(n41570) );
  NAND U42633 ( .A(n41568), .B(n41567), .Z(n41569) );
  AND U42634 ( .A(n41570), .B(n41569), .Z(n41618) );
  XOR U42635 ( .A(n41619), .B(n41618), .Z(n41620) );
  NANDN U42636 ( .A(n41572), .B(n41571), .Z(n41576) );
  NANDN U42637 ( .A(n41574), .B(n41573), .Z(n41575) );
  NAND U42638 ( .A(n41576), .B(n41575), .Z(n41621) );
  XOR U42639 ( .A(n41620), .B(n41621), .Z(n41588) );
  OR U42640 ( .A(n41578), .B(n41577), .Z(n41582) );
  NANDN U42641 ( .A(n41580), .B(n41579), .Z(n41581) );
  NAND U42642 ( .A(n41582), .B(n41581), .Z(n41589) );
  XNOR U42643 ( .A(n41588), .B(n41589), .Z(n41590) );
  XNOR U42644 ( .A(n41591), .B(n41590), .Z(n41624) );
  XNOR U42645 ( .A(n41624), .B(sreg[2028]), .Z(n41626) );
  NAND U42646 ( .A(n41583), .B(sreg[2027]), .Z(n41587) );
  OR U42647 ( .A(n41585), .B(n41584), .Z(n41586) );
  AND U42648 ( .A(n41587), .B(n41586), .Z(n41625) );
  XOR U42649 ( .A(n41626), .B(n41625), .Z(c[2028]) );
  NANDN U42650 ( .A(n41589), .B(n41588), .Z(n41593) );
  NAND U42651 ( .A(n41591), .B(n41590), .Z(n41592) );
  NAND U42652 ( .A(n41593), .B(n41592), .Z(n41632) );
  NAND U42653 ( .A(b[0]), .B(a[1013]), .Z(n41594) );
  XNOR U42654 ( .A(b[1]), .B(n41594), .Z(n41596) );
  NAND U42655 ( .A(n159), .B(a[1012]), .Z(n41595) );
  AND U42656 ( .A(n41596), .B(n41595), .Z(n41649) );
  XOR U42657 ( .A(a[1009]), .B(n42197), .Z(n41638) );
  NANDN U42658 ( .A(n41638), .B(n42173), .Z(n41599) );
  NANDN U42659 ( .A(n41597), .B(n42172), .Z(n41598) );
  NAND U42660 ( .A(n41599), .B(n41598), .Z(n41647) );
  NAND U42661 ( .A(b[7]), .B(a[1005]), .Z(n41648) );
  XNOR U42662 ( .A(n41647), .B(n41648), .Z(n41650) );
  XOR U42663 ( .A(n41649), .B(n41650), .Z(n41656) );
  NANDN U42664 ( .A(n41600), .B(n42093), .Z(n41602) );
  XOR U42665 ( .A(n42134), .B(a[1011]), .Z(n41641) );
  NANDN U42666 ( .A(n41641), .B(n42095), .Z(n41601) );
  NAND U42667 ( .A(n41602), .B(n41601), .Z(n41654) );
  NANDN U42668 ( .A(n41603), .B(n42231), .Z(n41605) );
  XOR U42669 ( .A(n246), .B(a[1007]), .Z(n41644) );
  NANDN U42670 ( .A(n41644), .B(n42234), .Z(n41604) );
  AND U42671 ( .A(n41605), .B(n41604), .Z(n41653) );
  XNOR U42672 ( .A(n41654), .B(n41653), .Z(n41655) );
  XNOR U42673 ( .A(n41656), .B(n41655), .Z(n41660) );
  NANDN U42674 ( .A(n41607), .B(n41606), .Z(n41611) );
  NAND U42675 ( .A(n41609), .B(n41608), .Z(n41610) );
  AND U42676 ( .A(n41611), .B(n41610), .Z(n41659) );
  XOR U42677 ( .A(n41660), .B(n41659), .Z(n41661) );
  NANDN U42678 ( .A(n41613), .B(n41612), .Z(n41617) );
  NANDN U42679 ( .A(n41615), .B(n41614), .Z(n41616) );
  NAND U42680 ( .A(n41617), .B(n41616), .Z(n41662) );
  XOR U42681 ( .A(n41661), .B(n41662), .Z(n41629) );
  OR U42682 ( .A(n41619), .B(n41618), .Z(n41623) );
  NANDN U42683 ( .A(n41621), .B(n41620), .Z(n41622) );
  NAND U42684 ( .A(n41623), .B(n41622), .Z(n41630) );
  XNOR U42685 ( .A(n41629), .B(n41630), .Z(n41631) );
  XNOR U42686 ( .A(n41632), .B(n41631), .Z(n41665) );
  XNOR U42687 ( .A(n41665), .B(sreg[2029]), .Z(n41667) );
  NAND U42688 ( .A(n41624), .B(sreg[2028]), .Z(n41628) );
  OR U42689 ( .A(n41626), .B(n41625), .Z(n41627) );
  AND U42690 ( .A(n41628), .B(n41627), .Z(n41666) );
  XOR U42691 ( .A(n41667), .B(n41666), .Z(c[2029]) );
  NANDN U42692 ( .A(n41630), .B(n41629), .Z(n41634) );
  NAND U42693 ( .A(n41632), .B(n41631), .Z(n41633) );
  NAND U42694 ( .A(n41634), .B(n41633), .Z(n41673) );
  NAND U42695 ( .A(b[0]), .B(a[1014]), .Z(n41635) );
  XNOR U42696 ( .A(b[1]), .B(n41635), .Z(n41637) );
  NAND U42697 ( .A(n159), .B(a[1013]), .Z(n41636) );
  AND U42698 ( .A(n41637), .B(n41636), .Z(n41690) );
  XOR U42699 ( .A(a[1010]), .B(n42197), .Z(n41679) );
  NANDN U42700 ( .A(n41679), .B(n42173), .Z(n41640) );
  NANDN U42701 ( .A(n41638), .B(n42172), .Z(n41639) );
  NAND U42702 ( .A(n41640), .B(n41639), .Z(n41688) );
  NAND U42703 ( .A(b[7]), .B(a[1006]), .Z(n41689) );
  XNOR U42704 ( .A(n41688), .B(n41689), .Z(n41691) );
  XOR U42705 ( .A(n41690), .B(n41691), .Z(n41697) );
  NANDN U42706 ( .A(n41641), .B(n42093), .Z(n41643) );
  XOR U42707 ( .A(n42134), .B(a[1012]), .Z(n41682) );
  NANDN U42708 ( .A(n41682), .B(n42095), .Z(n41642) );
  NAND U42709 ( .A(n41643), .B(n41642), .Z(n41695) );
  NANDN U42710 ( .A(n41644), .B(n42231), .Z(n41646) );
  XOR U42711 ( .A(n246), .B(a[1008]), .Z(n41685) );
  NANDN U42712 ( .A(n41685), .B(n42234), .Z(n41645) );
  AND U42713 ( .A(n41646), .B(n41645), .Z(n41694) );
  XNOR U42714 ( .A(n41695), .B(n41694), .Z(n41696) );
  XNOR U42715 ( .A(n41697), .B(n41696), .Z(n41701) );
  NANDN U42716 ( .A(n41648), .B(n41647), .Z(n41652) );
  NAND U42717 ( .A(n41650), .B(n41649), .Z(n41651) );
  AND U42718 ( .A(n41652), .B(n41651), .Z(n41700) );
  XOR U42719 ( .A(n41701), .B(n41700), .Z(n41702) );
  NANDN U42720 ( .A(n41654), .B(n41653), .Z(n41658) );
  NANDN U42721 ( .A(n41656), .B(n41655), .Z(n41657) );
  NAND U42722 ( .A(n41658), .B(n41657), .Z(n41703) );
  XOR U42723 ( .A(n41702), .B(n41703), .Z(n41670) );
  OR U42724 ( .A(n41660), .B(n41659), .Z(n41664) );
  NANDN U42725 ( .A(n41662), .B(n41661), .Z(n41663) );
  NAND U42726 ( .A(n41664), .B(n41663), .Z(n41671) );
  XNOR U42727 ( .A(n41670), .B(n41671), .Z(n41672) );
  XNOR U42728 ( .A(n41673), .B(n41672), .Z(n41706) );
  XNOR U42729 ( .A(n41706), .B(sreg[2030]), .Z(n41708) );
  NAND U42730 ( .A(n41665), .B(sreg[2029]), .Z(n41669) );
  OR U42731 ( .A(n41667), .B(n41666), .Z(n41668) );
  AND U42732 ( .A(n41669), .B(n41668), .Z(n41707) );
  XOR U42733 ( .A(n41708), .B(n41707), .Z(c[2030]) );
  NANDN U42734 ( .A(n41671), .B(n41670), .Z(n41675) );
  NAND U42735 ( .A(n41673), .B(n41672), .Z(n41674) );
  NAND U42736 ( .A(n41675), .B(n41674), .Z(n41714) );
  NAND U42737 ( .A(b[0]), .B(a[1015]), .Z(n41676) );
  XNOR U42738 ( .A(b[1]), .B(n41676), .Z(n41678) );
  NAND U42739 ( .A(n160), .B(a[1014]), .Z(n41677) );
  AND U42740 ( .A(n41678), .B(n41677), .Z(n41731) );
  XOR U42741 ( .A(a[1011]), .B(n42197), .Z(n41720) );
  NANDN U42742 ( .A(n41720), .B(n42173), .Z(n41681) );
  NANDN U42743 ( .A(n41679), .B(n42172), .Z(n41680) );
  NAND U42744 ( .A(n41681), .B(n41680), .Z(n41729) );
  NAND U42745 ( .A(b[7]), .B(a[1007]), .Z(n41730) );
  XNOR U42746 ( .A(n41729), .B(n41730), .Z(n41732) );
  XOR U42747 ( .A(n41731), .B(n41732), .Z(n41738) );
  NANDN U42748 ( .A(n41682), .B(n42093), .Z(n41684) );
  XOR U42749 ( .A(n42134), .B(a[1013]), .Z(n41723) );
  NANDN U42750 ( .A(n41723), .B(n42095), .Z(n41683) );
  NAND U42751 ( .A(n41684), .B(n41683), .Z(n41736) );
  NANDN U42752 ( .A(n41685), .B(n42231), .Z(n41687) );
  XOR U42753 ( .A(n246), .B(a[1009]), .Z(n41726) );
  NANDN U42754 ( .A(n41726), .B(n42234), .Z(n41686) );
  AND U42755 ( .A(n41687), .B(n41686), .Z(n41735) );
  XNOR U42756 ( .A(n41736), .B(n41735), .Z(n41737) );
  XNOR U42757 ( .A(n41738), .B(n41737), .Z(n41742) );
  NANDN U42758 ( .A(n41689), .B(n41688), .Z(n41693) );
  NAND U42759 ( .A(n41691), .B(n41690), .Z(n41692) );
  AND U42760 ( .A(n41693), .B(n41692), .Z(n41741) );
  XOR U42761 ( .A(n41742), .B(n41741), .Z(n41743) );
  NANDN U42762 ( .A(n41695), .B(n41694), .Z(n41699) );
  NANDN U42763 ( .A(n41697), .B(n41696), .Z(n41698) );
  NAND U42764 ( .A(n41699), .B(n41698), .Z(n41744) );
  XOR U42765 ( .A(n41743), .B(n41744), .Z(n41711) );
  OR U42766 ( .A(n41701), .B(n41700), .Z(n41705) );
  NANDN U42767 ( .A(n41703), .B(n41702), .Z(n41704) );
  NAND U42768 ( .A(n41705), .B(n41704), .Z(n41712) );
  XNOR U42769 ( .A(n41711), .B(n41712), .Z(n41713) );
  XNOR U42770 ( .A(n41714), .B(n41713), .Z(n41747) );
  XNOR U42771 ( .A(n41747), .B(sreg[2031]), .Z(n41749) );
  NAND U42772 ( .A(n41706), .B(sreg[2030]), .Z(n41710) );
  OR U42773 ( .A(n41708), .B(n41707), .Z(n41709) );
  AND U42774 ( .A(n41710), .B(n41709), .Z(n41748) );
  XOR U42775 ( .A(n41749), .B(n41748), .Z(c[2031]) );
  NANDN U42776 ( .A(n41712), .B(n41711), .Z(n41716) );
  NAND U42777 ( .A(n41714), .B(n41713), .Z(n41715) );
  NAND U42778 ( .A(n41716), .B(n41715), .Z(n41755) );
  NAND U42779 ( .A(b[0]), .B(a[1016]), .Z(n41717) );
  XNOR U42780 ( .A(b[1]), .B(n41717), .Z(n41719) );
  NAND U42781 ( .A(a[1015]), .B(n160), .Z(n41718) );
  AND U42782 ( .A(n41719), .B(n41718), .Z(n41772) );
  XOR U42783 ( .A(a[1012]), .B(n42197), .Z(n41761) );
  NANDN U42784 ( .A(n41761), .B(n42173), .Z(n41722) );
  NANDN U42785 ( .A(n41720), .B(n42172), .Z(n41721) );
  NAND U42786 ( .A(n41722), .B(n41721), .Z(n41770) );
  NAND U42787 ( .A(b[7]), .B(a[1008]), .Z(n41771) );
  XNOR U42788 ( .A(n41770), .B(n41771), .Z(n41773) );
  XOR U42789 ( .A(n41772), .B(n41773), .Z(n41779) );
  NANDN U42790 ( .A(n41723), .B(n42093), .Z(n41725) );
  XOR U42791 ( .A(n42134), .B(a[1014]), .Z(n41764) );
  NANDN U42792 ( .A(n41764), .B(n42095), .Z(n41724) );
  NAND U42793 ( .A(n41725), .B(n41724), .Z(n41777) );
  NANDN U42794 ( .A(n41726), .B(n42231), .Z(n41728) );
  XOR U42795 ( .A(n246), .B(a[1010]), .Z(n41767) );
  NANDN U42796 ( .A(n41767), .B(n42234), .Z(n41727) );
  AND U42797 ( .A(n41728), .B(n41727), .Z(n41776) );
  XNOR U42798 ( .A(n41777), .B(n41776), .Z(n41778) );
  XNOR U42799 ( .A(n41779), .B(n41778), .Z(n41783) );
  NANDN U42800 ( .A(n41730), .B(n41729), .Z(n41734) );
  NAND U42801 ( .A(n41732), .B(n41731), .Z(n41733) );
  AND U42802 ( .A(n41734), .B(n41733), .Z(n41782) );
  XOR U42803 ( .A(n41783), .B(n41782), .Z(n41784) );
  NANDN U42804 ( .A(n41736), .B(n41735), .Z(n41740) );
  NANDN U42805 ( .A(n41738), .B(n41737), .Z(n41739) );
  NAND U42806 ( .A(n41740), .B(n41739), .Z(n41785) );
  XOR U42807 ( .A(n41784), .B(n41785), .Z(n41752) );
  OR U42808 ( .A(n41742), .B(n41741), .Z(n41746) );
  NANDN U42809 ( .A(n41744), .B(n41743), .Z(n41745) );
  NAND U42810 ( .A(n41746), .B(n41745), .Z(n41753) );
  XNOR U42811 ( .A(n41752), .B(n41753), .Z(n41754) );
  XNOR U42812 ( .A(n41755), .B(n41754), .Z(n41788) );
  XNOR U42813 ( .A(n41788), .B(sreg[2032]), .Z(n41790) );
  NAND U42814 ( .A(n41747), .B(sreg[2031]), .Z(n41751) );
  OR U42815 ( .A(n41749), .B(n41748), .Z(n41750) );
  AND U42816 ( .A(n41751), .B(n41750), .Z(n41789) );
  XOR U42817 ( .A(n41790), .B(n41789), .Z(c[2032]) );
  NANDN U42818 ( .A(n41753), .B(n41752), .Z(n41757) );
  NAND U42819 ( .A(n41755), .B(n41754), .Z(n41756) );
  NAND U42820 ( .A(n41757), .B(n41756), .Z(n41796) );
  NAND U42821 ( .A(b[0]), .B(a[1017]), .Z(n41758) );
  XNOR U42822 ( .A(b[1]), .B(n41758), .Z(n41760) );
  NAND U42823 ( .A(n160), .B(a[1016]), .Z(n41759) );
  AND U42824 ( .A(n41760), .B(n41759), .Z(n41813) );
  XOR U42825 ( .A(a[1013]), .B(n42197), .Z(n41802) );
  NANDN U42826 ( .A(n41802), .B(n42173), .Z(n41763) );
  NANDN U42827 ( .A(n41761), .B(n42172), .Z(n41762) );
  NAND U42828 ( .A(n41763), .B(n41762), .Z(n41811) );
  NAND U42829 ( .A(b[7]), .B(a[1009]), .Z(n41812) );
  XNOR U42830 ( .A(n41811), .B(n41812), .Z(n41814) );
  XOR U42831 ( .A(n41813), .B(n41814), .Z(n41820) );
  NANDN U42832 ( .A(n41764), .B(n42093), .Z(n41766) );
  IV U42833 ( .A(a[1015]), .Z(n41932) );
  XNOR U42834 ( .A(n42134), .B(n41932), .Z(n41805) );
  NANDN U42835 ( .A(n41805), .B(n42095), .Z(n41765) );
  NAND U42836 ( .A(n41766), .B(n41765), .Z(n41818) );
  NANDN U42837 ( .A(n41767), .B(n42231), .Z(n41769) );
  XOR U42838 ( .A(n246), .B(a[1011]), .Z(n41808) );
  NANDN U42839 ( .A(n41808), .B(n42234), .Z(n41768) );
  AND U42840 ( .A(n41769), .B(n41768), .Z(n41817) );
  XNOR U42841 ( .A(n41818), .B(n41817), .Z(n41819) );
  XNOR U42842 ( .A(n41820), .B(n41819), .Z(n41824) );
  NANDN U42843 ( .A(n41771), .B(n41770), .Z(n41775) );
  NAND U42844 ( .A(n41773), .B(n41772), .Z(n41774) );
  AND U42845 ( .A(n41775), .B(n41774), .Z(n41823) );
  XOR U42846 ( .A(n41824), .B(n41823), .Z(n41825) );
  NANDN U42847 ( .A(n41777), .B(n41776), .Z(n41781) );
  NANDN U42848 ( .A(n41779), .B(n41778), .Z(n41780) );
  NAND U42849 ( .A(n41781), .B(n41780), .Z(n41826) );
  XOR U42850 ( .A(n41825), .B(n41826), .Z(n41793) );
  OR U42851 ( .A(n41783), .B(n41782), .Z(n41787) );
  NANDN U42852 ( .A(n41785), .B(n41784), .Z(n41786) );
  NAND U42853 ( .A(n41787), .B(n41786), .Z(n41794) );
  XNOR U42854 ( .A(n41793), .B(n41794), .Z(n41795) );
  XNOR U42855 ( .A(n41796), .B(n41795), .Z(n41829) );
  XNOR U42856 ( .A(n41829), .B(sreg[2033]), .Z(n41831) );
  NAND U42857 ( .A(n41788), .B(sreg[2032]), .Z(n41792) );
  OR U42858 ( .A(n41790), .B(n41789), .Z(n41791) );
  AND U42859 ( .A(n41792), .B(n41791), .Z(n41830) );
  XOR U42860 ( .A(n41831), .B(n41830), .Z(c[2033]) );
  NANDN U42861 ( .A(n41794), .B(n41793), .Z(n41798) );
  NAND U42862 ( .A(n41796), .B(n41795), .Z(n41797) );
  NAND U42863 ( .A(n41798), .B(n41797), .Z(n41837) );
  NAND U42864 ( .A(b[0]), .B(a[1018]), .Z(n41799) );
  XNOR U42865 ( .A(b[1]), .B(n41799), .Z(n41801) );
  NAND U42866 ( .A(a[1017]), .B(n160), .Z(n41800) );
  AND U42867 ( .A(n41801), .B(n41800), .Z(n41854) );
  XOR U42868 ( .A(a[1014]), .B(n42197), .Z(n41843) );
  NANDN U42869 ( .A(n41843), .B(n42173), .Z(n41804) );
  NANDN U42870 ( .A(n41802), .B(n42172), .Z(n41803) );
  NAND U42871 ( .A(n41804), .B(n41803), .Z(n41852) );
  NAND U42872 ( .A(b[7]), .B(a[1010]), .Z(n41853) );
  XNOR U42873 ( .A(n41852), .B(n41853), .Z(n41855) );
  XOR U42874 ( .A(n41854), .B(n41855), .Z(n41861) );
  NANDN U42875 ( .A(n41805), .B(n42093), .Z(n41807) );
  XOR U42876 ( .A(n42134), .B(a[1016]), .Z(n41846) );
  NANDN U42877 ( .A(n41846), .B(n42095), .Z(n41806) );
  NAND U42878 ( .A(n41807), .B(n41806), .Z(n41859) );
  NANDN U42879 ( .A(n41808), .B(n42231), .Z(n41810) );
  XOR U42880 ( .A(n246), .B(a[1012]), .Z(n41849) );
  NANDN U42881 ( .A(n41849), .B(n42234), .Z(n41809) );
  AND U42882 ( .A(n41810), .B(n41809), .Z(n41858) );
  XNOR U42883 ( .A(n41859), .B(n41858), .Z(n41860) );
  XNOR U42884 ( .A(n41861), .B(n41860), .Z(n41865) );
  NANDN U42885 ( .A(n41812), .B(n41811), .Z(n41816) );
  NAND U42886 ( .A(n41814), .B(n41813), .Z(n41815) );
  AND U42887 ( .A(n41816), .B(n41815), .Z(n41864) );
  XOR U42888 ( .A(n41865), .B(n41864), .Z(n41866) );
  NANDN U42889 ( .A(n41818), .B(n41817), .Z(n41822) );
  NANDN U42890 ( .A(n41820), .B(n41819), .Z(n41821) );
  NAND U42891 ( .A(n41822), .B(n41821), .Z(n41867) );
  XOR U42892 ( .A(n41866), .B(n41867), .Z(n41834) );
  OR U42893 ( .A(n41824), .B(n41823), .Z(n41828) );
  NANDN U42894 ( .A(n41826), .B(n41825), .Z(n41827) );
  NAND U42895 ( .A(n41828), .B(n41827), .Z(n41835) );
  XNOR U42896 ( .A(n41834), .B(n41835), .Z(n41836) );
  XNOR U42897 ( .A(n41837), .B(n41836), .Z(n41870) );
  XNOR U42898 ( .A(n41870), .B(sreg[2034]), .Z(n41872) );
  NAND U42899 ( .A(n41829), .B(sreg[2033]), .Z(n41833) );
  OR U42900 ( .A(n41831), .B(n41830), .Z(n41832) );
  AND U42901 ( .A(n41833), .B(n41832), .Z(n41871) );
  XOR U42902 ( .A(n41872), .B(n41871), .Z(c[2034]) );
  NANDN U42903 ( .A(n41835), .B(n41834), .Z(n41839) );
  NAND U42904 ( .A(n41837), .B(n41836), .Z(n41838) );
  NAND U42905 ( .A(n41839), .B(n41838), .Z(n41878) );
  NAND U42906 ( .A(b[0]), .B(a[1019]), .Z(n41840) );
  XNOR U42907 ( .A(b[1]), .B(n41840), .Z(n41842) );
  NAND U42908 ( .A(a[1018]), .B(n160), .Z(n41841) );
  AND U42909 ( .A(n41842), .B(n41841), .Z(n41895) );
  XOR U42910 ( .A(a[1015]), .B(n42197), .Z(n41884) );
  NANDN U42911 ( .A(n41884), .B(n42173), .Z(n41845) );
  NANDN U42912 ( .A(n41843), .B(n42172), .Z(n41844) );
  NAND U42913 ( .A(n41845), .B(n41844), .Z(n41893) );
  NAND U42914 ( .A(b[7]), .B(a[1011]), .Z(n41894) );
  XNOR U42915 ( .A(n41893), .B(n41894), .Z(n41896) );
  XOR U42916 ( .A(n41895), .B(n41896), .Z(n41902) );
  NANDN U42917 ( .A(n41846), .B(n42093), .Z(n41848) );
  IV U42918 ( .A(a[1017]), .Z(n42098) );
  XNOR U42919 ( .A(n42134), .B(n42098), .Z(n41887) );
  NANDN U42920 ( .A(n41887), .B(n42095), .Z(n41847) );
  NAND U42921 ( .A(n41848), .B(n41847), .Z(n41900) );
  NANDN U42922 ( .A(n41849), .B(n42231), .Z(n41851) );
  XOR U42923 ( .A(n246), .B(a[1013]), .Z(n41890) );
  NANDN U42924 ( .A(n41890), .B(n42234), .Z(n41850) );
  AND U42925 ( .A(n41851), .B(n41850), .Z(n41899) );
  XNOR U42926 ( .A(n41900), .B(n41899), .Z(n41901) );
  XNOR U42927 ( .A(n41902), .B(n41901), .Z(n41906) );
  NANDN U42928 ( .A(n41853), .B(n41852), .Z(n41857) );
  NAND U42929 ( .A(n41855), .B(n41854), .Z(n41856) );
  AND U42930 ( .A(n41857), .B(n41856), .Z(n41905) );
  XOR U42931 ( .A(n41906), .B(n41905), .Z(n41907) );
  NANDN U42932 ( .A(n41859), .B(n41858), .Z(n41863) );
  NANDN U42933 ( .A(n41861), .B(n41860), .Z(n41862) );
  NAND U42934 ( .A(n41863), .B(n41862), .Z(n41908) );
  XOR U42935 ( .A(n41907), .B(n41908), .Z(n41875) );
  OR U42936 ( .A(n41865), .B(n41864), .Z(n41869) );
  NANDN U42937 ( .A(n41867), .B(n41866), .Z(n41868) );
  NAND U42938 ( .A(n41869), .B(n41868), .Z(n41876) );
  XNOR U42939 ( .A(n41875), .B(n41876), .Z(n41877) );
  XNOR U42940 ( .A(n41878), .B(n41877), .Z(n41911) );
  XNOR U42941 ( .A(n41911), .B(sreg[2035]), .Z(n41913) );
  NAND U42942 ( .A(n41870), .B(sreg[2034]), .Z(n41874) );
  OR U42943 ( .A(n41872), .B(n41871), .Z(n41873) );
  AND U42944 ( .A(n41874), .B(n41873), .Z(n41912) );
  XOR U42945 ( .A(n41913), .B(n41912), .Z(c[2035]) );
  NANDN U42946 ( .A(n41876), .B(n41875), .Z(n41880) );
  NAND U42947 ( .A(n41878), .B(n41877), .Z(n41879) );
  NAND U42948 ( .A(n41880), .B(n41879), .Z(n41919) );
  NAND U42949 ( .A(b[0]), .B(a[1020]), .Z(n41881) );
  XNOR U42950 ( .A(b[1]), .B(n41881), .Z(n41883) );
  NAND U42951 ( .A(n160), .B(a[1019]), .Z(n41882) );
  AND U42952 ( .A(n41883), .B(n41882), .Z(n41937) );
  XOR U42953 ( .A(a[1016]), .B(n42197), .Z(n41925) );
  NANDN U42954 ( .A(n41925), .B(n42173), .Z(n41886) );
  NANDN U42955 ( .A(n41884), .B(n42172), .Z(n41885) );
  NAND U42956 ( .A(n41886), .B(n41885), .Z(n41935) );
  NAND U42957 ( .A(b[7]), .B(a[1012]), .Z(n41936) );
  XNOR U42958 ( .A(n41935), .B(n41936), .Z(n41938) );
  XOR U42959 ( .A(n41937), .B(n41938), .Z(n41944) );
  NANDN U42960 ( .A(n41887), .B(n42093), .Z(n41889) );
  IV U42961 ( .A(a[1018]), .Z(n42071) );
  XNOR U42962 ( .A(n42134), .B(n42071), .Z(n41928) );
  NANDN U42963 ( .A(n41928), .B(n42095), .Z(n41888) );
  NAND U42964 ( .A(n41889), .B(n41888), .Z(n41942) );
  NANDN U42965 ( .A(n41890), .B(n42231), .Z(n41892) );
  XOR U42966 ( .A(n246), .B(a[1014]), .Z(n41931) );
  NANDN U42967 ( .A(n41931), .B(n42234), .Z(n41891) );
  AND U42968 ( .A(n41892), .B(n41891), .Z(n41941) );
  XNOR U42969 ( .A(n41942), .B(n41941), .Z(n41943) );
  XNOR U42970 ( .A(n41944), .B(n41943), .Z(n41948) );
  NANDN U42971 ( .A(n41894), .B(n41893), .Z(n41898) );
  NAND U42972 ( .A(n41896), .B(n41895), .Z(n41897) );
  AND U42973 ( .A(n41898), .B(n41897), .Z(n41947) );
  XOR U42974 ( .A(n41948), .B(n41947), .Z(n41949) );
  NANDN U42975 ( .A(n41900), .B(n41899), .Z(n41904) );
  NANDN U42976 ( .A(n41902), .B(n41901), .Z(n41903) );
  NAND U42977 ( .A(n41904), .B(n41903), .Z(n41950) );
  XOR U42978 ( .A(n41949), .B(n41950), .Z(n41916) );
  OR U42979 ( .A(n41906), .B(n41905), .Z(n41910) );
  NANDN U42980 ( .A(n41908), .B(n41907), .Z(n41909) );
  NAND U42981 ( .A(n41910), .B(n41909), .Z(n41917) );
  XNOR U42982 ( .A(n41916), .B(n41917), .Z(n41918) );
  XNOR U42983 ( .A(n41919), .B(n41918), .Z(n41953) );
  XNOR U42984 ( .A(n41953), .B(sreg[2036]), .Z(n41955) );
  NAND U42985 ( .A(n41911), .B(sreg[2035]), .Z(n41915) );
  OR U42986 ( .A(n41913), .B(n41912), .Z(n41914) );
  AND U42987 ( .A(n41915), .B(n41914), .Z(n41954) );
  XOR U42988 ( .A(n41955), .B(n41954), .Z(c[2036]) );
  NANDN U42989 ( .A(n41917), .B(n41916), .Z(n41921) );
  NAND U42990 ( .A(n41919), .B(n41918), .Z(n41920) );
  NAND U42991 ( .A(n41921), .B(n41920), .Z(n41961) );
  NAND U42992 ( .A(b[0]), .B(a[1021]), .Z(n41922) );
  XNOR U42993 ( .A(b[1]), .B(n41922), .Z(n41924) );
  NAND U42994 ( .A(a[1020]), .B(n160), .Z(n41923) );
  AND U42995 ( .A(n41924), .B(n41923), .Z(n41978) );
  XOR U42996 ( .A(a[1017]), .B(n42197), .Z(n41967) );
  NANDN U42997 ( .A(n41967), .B(n42173), .Z(n41927) );
  NANDN U42998 ( .A(n41925), .B(n42172), .Z(n41926) );
  NAND U42999 ( .A(n41927), .B(n41926), .Z(n41976) );
  NAND U43000 ( .A(b[7]), .B(a[1013]), .Z(n41977) );
  XNOR U43001 ( .A(n41976), .B(n41977), .Z(n41979) );
  XOR U43002 ( .A(n41978), .B(n41979), .Z(n41985) );
  NANDN U43003 ( .A(n41928), .B(n42093), .Z(n41930) );
  XOR U43004 ( .A(n42134), .B(a[1019]), .Z(n41970) );
  NANDN U43005 ( .A(n41970), .B(n42095), .Z(n41929) );
  NAND U43006 ( .A(n41930), .B(n41929), .Z(n41983) );
  NANDN U43007 ( .A(n41931), .B(n42231), .Z(n41934) );
  XNOR U43008 ( .A(n246), .B(n41932), .Z(n41973) );
  NANDN U43009 ( .A(n41973), .B(n42234), .Z(n41933) );
  AND U43010 ( .A(n41934), .B(n41933), .Z(n41982) );
  XNOR U43011 ( .A(n41983), .B(n41982), .Z(n41984) );
  XNOR U43012 ( .A(n41985), .B(n41984), .Z(n41989) );
  NANDN U43013 ( .A(n41936), .B(n41935), .Z(n41940) );
  NAND U43014 ( .A(n41938), .B(n41937), .Z(n41939) );
  AND U43015 ( .A(n41940), .B(n41939), .Z(n41988) );
  XOR U43016 ( .A(n41989), .B(n41988), .Z(n41990) );
  NANDN U43017 ( .A(n41942), .B(n41941), .Z(n41946) );
  NANDN U43018 ( .A(n41944), .B(n41943), .Z(n41945) );
  NAND U43019 ( .A(n41946), .B(n41945), .Z(n41991) );
  XOR U43020 ( .A(n41990), .B(n41991), .Z(n41958) );
  OR U43021 ( .A(n41948), .B(n41947), .Z(n41952) );
  NANDN U43022 ( .A(n41950), .B(n41949), .Z(n41951) );
  NAND U43023 ( .A(n41952), .B(n41951), .Z(n41959) );
  XNOR U43024 ( .A(n41958), .B(n41959), .Z(n41960) );
  XNOR U43025 ( .A(n41961), .B(n41960), .Z(n41994) );
  XNOR U43026 ( .A(n41994), .B(sreg[2037]), .Z(n41996) );
  NAND U43027 ( .A(n41953), .B(sreg[2036]), .Z(n41957) );
  OR U43028 ( .A(n41955), .B(n41954), .Z(n41956) );
  AND U43029 ( .A(n41957), .B(n41956), .Z(n41995) );
  XOR U43030 ( .A(n41996), .B(n41995), .Z(c[2037]) );
  NANDN U43031 ( .A(n41959), .B(n41958), .Z(n41963) );
  NAND U43032 ( .A(n41961), .B(n41960), .Z(n41962) );
  NAND U43033 ( .A(n41963), .B(n41962), .Z(n42002) );
  NAND U43034 ( .A(b[0]), .B(a[1022]), .Z(n41964) );
  XNOR U43035 ( .A(b[1]), .B(n41964), .Z(n41966) );
  NAND U43036 ( .A(a[1021]), .B(n161), .Z(n41965) );
  AND U43037 ( .A(n41966), .B(n41965), .Z(n42031) );
  XNOR U43038 ( .A(n42197), .B(n42071), .Z(n42014) );
  NANDN U43039 ( .A(n42014), .B(n42173), .Z(n41969) );
  NANDN U43040 ( .A(n41967), .B(n42172), .Z(n41968) );
  NAND U43041 ( .A(n41969), .B(n41968), .Z(n42029) );
  NAND U43042 ( .A(b[7]), .B(a[1014]), .Z(n42030) );
  XOR U43043 ( .A(n42031), .B(n42032), .Z(n42026) );
  NANDN U43044 ( .A(n41970), .B(n42093), .Z(n41972) );
  IV U43045 ( .A(a[1020]), .Z(n42143) );
  XNOR U43046 ( .A(n42143), .B(b[3]), .Z(n42017) );
  NAND U43047 ( .A(n42017), .B(n42095), .Z(n41971) );
  NAND U43048 ( .A(n41972), .B(n41971), .Z(n42024) );
  NANDN U43049 ( .A(n41973), .B(n42231), .Z(n41975) );
  XOR U43050 ( .A(a[1016]), .B(b[7]), .Z(n42020) );
  NAND U43051 ( .A(n42234), .B(n42020), .Z(n41974) );
  AND U43052 ( .A(n41975), .B(n41974), .Z(n42023) );
  XNOR U43053 ( .A(n42024), .B(n42023), .Z(n42025) );
  XNOR U43054 ( .A(n42026), .B(n42025), .Z(n42006) );
  NANDN U43055 ( .A(n41977), .B(n41976), .Z(n41981) );
  NAND U43056 ( .A(n41979), .B(n41978), .Z(n41980) );
  AND U43057 ( .A(n41981), .B(n41980), .Z(n42005) );
  XOR U43058 ( .A(n42006), .B(n42005), .Z(n42007) );
  NANDN U43059 ( .A(n41983), .B(n41982), .Z(n41987) );
  NANDN U43060 ( .A(n41985), .B(n41984), .Z(n41986) );
  NAND U43061 ( .A(n41987), .B(n41986), .Z(n42008) );
  XOR U43062 ( .A(n42007), .B(n42008), .Z(n41999) );
  OR U43063 ( .A(n41989), .B(n41988), .Z(n41993) );
  NANDN U43064 ( .A(n41991), .B(n41990), .Z(n41992) );
  NAND U43065 ( .A(n41993), .B(n41992), .Z(n42000) );
  XNOR U43066 ( .A(n41999), .B(n42000), .Z(n42001) );
  XNOR U43067 ( .A(n42002), .B(n42001), .Z(n42035) );
  XNOR U43068 ( .A(n42035), .B(sreg[2038]), .Z(n42037) );
  NAND U43069 ( .A(n41994), .B(sreg[2037]), .Z(n41998) );
  OR U43070 ( .A(n41996), .B(n41995), .Z(n41997) );
  AND U43071 ( .A(n41998), .B(n41997), .Z(n42036) );
  XOR U43072 ( .A(n42037), .B(n42036), .Z(c[2038]) );
  NANDN U43073 ( .A(n42000), .B(n41999), .Z(n42004) );
  NAND U43074 ( .A(n42002), .B(n42001), .Z(n42003) );
  NAND U43075 ( .A(n42004), .B(n42003), .Z(n42043) );
  OR U43076 ( .A(n42006), .B(n42005), .Z(n42010) );
  NANDN U43077 ( .A(n42008), .B(n42007), .Z(n42009) );
  NAND U43078 ( .A(n42010), .B(n42009), .Z(n42040) );
  AND U43079 ( .A(b[7]), .B(a[1015]), .Z(n42061) );
  NAND U43080 ( .A(b[0]), .B(a[1023]), .Z(n42011) );
  XNOR U43081 ( .A(b[1]), .B(n42011), .Z(n42013) );
  NAND U43082 ( .A(a[1022]), .B(n161), .Z(n42012) );
  AND U43083 ( .A(n42013), .B(n42012), .Z(n42059) );
  NANDN U43084 ( .A(n42014), .B(n42172), .Z(n42016) );
  XOR U43085 ( .A(a[1019]), .B(b[5]), .Z(n42064) );
  NAND U43086 ( .A(n42173), .B(n42064), .Z(n42015) );
  AND U43087 ( .A(n42016), .B(n42015), .Z(n42058) );
  XNOR U43088 ( .A(n42059), .B(n42058), .Z(n42060) );
  XOR U43089 ( .A(n42061), .B(n42060), .Z(n42055) );
  IV U43090 ( .A(a[1021]), .Z(n42168) );
  XNOR U43091 ( .A(n42134), .B(n42168), .Z(n42067) );
  NANDN U43092 ( .A(n42067), .B(n42095), .Z(n42019) );
  NAND U43093 ( .A(n42093), .B(n42017), .Z(n42018) );
  NAND U43094 ( .A(n42019), .B(n42018), .Z(n42052) );
  NAND U43095 ( .A(n42231), .B(n42020), .Z(n42022) );
  XNOR U43096 ( .A(n246), .B(n42098), .Z(n42070) );
  NANDN U43097 ( .A(n42070), .B(n42234), .Z(n42021) );
  AND U43098 ( .A(n42022), .B(n42021), .Z(n42053) );
  XNOR U43099 ( .A(n42052), .B(n42053), .Z(n42054) );
  XOR U43100 ( .A(n42055), .B(n42054), .Z(n42049) );
  NANDN U43101 ( .A(n42024), .B(n42023), .Z(n42028) );
  NANDN U43102 ( .A(n42026), .B(n42025), .Z(n42027) );
  NAND U43103 ( .A(n42028), .B(n42027), .Z(n42046) );
  NANDN U43104 ( .A(n42030), .B(n42029), .Z(n42034) );
  NAND U43105 ( .A(n42032), .B(n42031), .Z(n42033) );
  NAND U43106 ( .A(n42034), .B(n42033), .Z(n42047) );
  XNOR U43107 ( .A(n42046), .B(n42047), .Z(n42048) );
  XOR U43108 ( .A(n42049), .B(n42048), .Z(n42041) );
  XOR U43109 ( .A(n42040), .B(n42041), .Z(n42042) );
  XNOR U43110 ( .A(n42043), .B(n42042), .Z(n42074) );
  XNOR U43111 ( .A(n42074), .B(sreg[2039]), .Z(n42076) );
  NAND U43112 ( .A(n42035), .B(sreg[2038]), .Z(n42039) );
  OR U43113 ( .A(n42037), .B(n42036), .Z(n42038) );
  AND U43114 ( .A(n42039), .B(n42038), .Z(n42075) );
  XOR U43115 ( .A(n42076), .B(n42075), .Z(c[2039]) );
  OR U43116 ( .A(n42041), .B(n42040), .Z(n42045) );
  NAND U43117 ( .A(n42043), .B(n42042), .Z(n42044) );
  NAND U43118 ( .A(n42045), .B(n42044), .Z(n42084) );
  NANDN U43119 ( .A(n42047), .B(n42046), .Z(n42051) );
  NANDN U43120 ( .A(n42049), .B(n42048), .Z(n42050) );
  NAND U43121 ( .A(n42051), .B(n42050), .Z(n42081) );
  NANDN U43122 ( .A(n42053), .B(n42052), .Z(n42057) );
  NAND U43123 ( .A(n42055), .B(n42054), .Z(n42056) );
  NAND U43124 ( .A(n42057), .B(n42056), .Z(n42090) );
  NANDN U43125 ( .A(n42059), .B(n42058), .Z(n42063) );
  NANDN U43126 ( .A(n42061), .B(n42060), .Z(n42062) );
  NAND U43127 ( .A(n42063), .B(n42062), .Z(n42087) );
  NAND U43128 ( .A(b[7]), .B(a[1016]), .Z(n42114) );
  XNOR U43129 ( .A(n42197), .B(n42143), .Z(n42102) );
  NANDN U43130 ( .A(n42102), .B(n42173), .Z(n42066) );
  NAND U43131 ( .A(n42172), .B(n42064), .Z(n42065) );
  NAND U43132 ( .A(n42066), .B(n42065), .Z(n42111) );
  IV U43133 ( .A(a[1023]), .Z(n42233) );
  XOR U43134 ( .A(n42114), .B(n42113), .Z(n42108) );
  NANDN U43135 ( .A(n42067), .B(n42093), .Z(n42069) );
  IV U43136 ( .A(a[1022]), .Z(n42203) );
  XNOR U43137 ( .A(n42134), .B(n42203), .Z(n42094) );
  NANDN U43138 ( .A(n42094), .B(n42095), .Z(n42068) );
  NAND U43139 ( .A(n42069), .B(n42068), .Z(n42106) );
  NANDN U43140 ( .A(n42070), .B(n42231), .Z(n42073) );
  XNOR U43141 ( .A(n246), .B(n42071), .Z(n42099) );
  NANDN U43142 ( .A(n42099), .B(n42234), .Z(n42072) );
  AND U43143 ( .A(n42073), .B(n42072), .Z(n42105) );
  XNOR U43144 ( .A(n42106), .B(n42105), .Z(n42107) );
  XNOR U43145 ( .A(n42108), .B(n42107), .Z(n42088) );
  XNOR U43146 ( .A(n42087), .B(n42088), .Z(n42089) );
  XOR U43147 ( .A(n42090), .B(n42089), .Z(n42082) );
  XNOR U43148 ( .A(n42081), .B(n42082), .Z(n42083) );
  XOR U43149 ( .A(n42084), .B(n42083), .Z(n42080) );
  NAND U43150 ( .A(n42074), .B(sreg[2039]), .Z(n42078) );
  OR U43151 ( .A(n42076), .B(n42075), .Z(n42077) );
  AND U43152 ( .A(n42078), .B(n42077), .Z(n42079) );
  XOR U43153 ( .A(n42080), .B(n42079), .Z(c[2040]) );
  OR U43154 ( .A(n42080), .B(n42079), .Z(n42152) );
  NANDN U43155 ( .A(n42082), .B(n42081), .Z(n42086) );
  NAND U43156 ( .A(n42084), .B(n42083), .Z(n42085) );
  NAND U43157 ( .A(n42086), .B(n42085), .Z(n42120) );
  NANDN U43158 ( .A(n42088), .B(n42087), .Z(n42092) );
  NANDN U43159 ( .A(n42090), .B(n42089), .Z(n42091) );
  NAND U43160 ( .A(n42092), .B(n42091), .Z(n42118) );
  NANDN U43161 ( .A(n42094), .B(n42093), .Z(n42097) );
  XNOR U43162 ( .A(n42233), .B(n42134), .Z(n42135) );
  NANDN U43163 ( .A(n42135), .B(n42095), .Z(n42096) );
  AND U43164 ( .A(n42097), .B(n42096), .Z(n42123) );
  XNOR U43165 ( .A(b[1]), .B(n42123), .Z(n42125) );
  NOR U43166 ( .A(n42098), .B(n246), .Z(n42208) );
  NANDN U43167 ( .A(n42099), .B(n42231), .Z(n42101) );
  XOR U43168 ( .A(n247), .B(a[1019]), .Z(n42142) );
  NANDN U43169 ( .A(n42142), .B(n42234), .Z(n42100) );
  AND U43170 ( .A(n42101), .B(n42100), .Z(n42128) );
  XNOR U43171 ( .A(n42208), .B(n42128), .Z(n42130) );
  NANDN U43172 ( .A(n42102), .B(n42172), .Z(n42104) );
  XNOR U43173 ( .A(n42197), .B(n42168), .Z(n42139) );
  NANDN U43174 ( .A(n42139), .B(n42173), .Z(n42103) );
  AND U43175 ( .A(n42104), .B(n42103), .Z(n42129) );
  XNOR U43176 ( .A(n42130), .B(n42129), .Z(n42124) );
  XOR U43177 ( .A(n42125), .B(n42124), .Z(n42148) );
  NANDN U43178 ( .A(n42106), .B(n42105), .Z(n42110) );
  NAND U43179 ( .A(n42108), .B(n42107), .Z(n42109) );
  NAND U43180 ( .A(n42110), .B(n42109), .Z(n42146) );
  NANDN U43181 ( .A(n42112), .B(n42111), .Z(n42116) );
  NANDN U43182 ( .A(n42114), .B(n42113), .Z(n42115) );
  NAND U43183 ( .A(n42116), .B(n42115), .Z(n42147) );
  XNOR U43184 ( .A(n42146), .B(n42147), .Z(n42149) );
  XNOR U43185 ( .A(n42148), .B(n42149), .Z(n42117) );
  XOR U43186 ( .A(n42118), .B(n42117), .Z(n42119) );
  XOR U43187 ( .A(n42120), .B(n42119), .Z(n42151) );
  XOR U43188 ( .A(n42152), .B(n42151), .Z(c[2041]) );
  NAND U43189 ( .A(n42118), .B(n42117), .Z(n42122) );
  NAND U43190 ( .A(n42120), .B(n42119), .Z(n42121) );
  AND U43191 ( .A(n42122), .B(n42121), .Z(n42157) );
  NAND U43192 ( .A(b[1]), .B(n42123), .Z(n42127) );
  NANDN U43193 ( .A(n42125), .B(n42124), .Z(n42126) );
  NAND U43194 ( .A(n42127), .B(n42126), .Z(n42178) );
  NAND U43195 ( .A(n42208), .B(n42128), .Z(n42132) );
  NANDN U43196 ( .A(n42130), .B(n42129), .Z(n42131) );
  NAND U43197 ( .A(n42132), .B(n42131), .Z(n42177) );
  AND U43198 ( .A(b[2]), .B(b[1]), .Z(n42133) );
  XNOR U43199 ( .A(n42134), .B(n42133), .Z(n42138) );
  XNOR U43200 ( .A(b[1]), .B(b[2]), .Z(n42136) );
  NAND U43201 ( .A(n42136), .B(n42135), .Z(n42137) );
  AND U43202 ( .A(n42138), .B(n42137), .Z(n42159) );
  ANDN U43203 ( .B(a[1018]), .A(n247), .Z(n42158) );
  XNOR U43204 ( .A(n42159), .B(n42158), .Z(n42160) );
  XOR U43205 ( .A(n42208), .B(n42160), .Z(n42164) );
  NANDN U43206 ( .A(n42139), .B(n42172), .Z(n42141) );
  XNOR U43207 ( .A(n42203), .B(b[5]), .Z(n42171) );
  NAND U43208 ( .A(n42173), .B(n42171), .Z(n42140) );
  NAND U43209 ( .A(n42141), .B(n42140), .Z(n42162) );
  NANDN U43210 ( .A(n42142), .B(n42231), .Z(n42145) );
  XNOR U43211 ( .A(n42143), .B(b[7]), .Z(n42167) );
  NAND U43212 ( .A(n42234), .B(n42167), .Z(n42144) );
  AND U43213 ( .A(n42145), .B(n42144), .Z(n42161) );
  XNOR U43214 ( .A(n42162), .B(n42161), .Z(n42163) );
  XNOR U43215 ( .A(n42164), .B(n42163), .Z(n42176) );
  XNOR U43216 ( .A(n42177), .B(n42176), .Z(n42179) );
  XOR U43217 ( .A(n42178), .B(n42179), .Z(n42155) );
  XOR U43218 ( .A(n42155), .B(n42156), .Z(n42150) );
  XOR U43219 ( .A(n42157), .B(n42150), .Z(n42153) );
  OR U43220 ( .A(n42152), .B(n42151), .Z(n42154) );
  XNOR U43221 ( .A(n42153), .B(n42154), .Z(c[2042]) );
  NANDN U43222 ( .A(n42154), .B(n42153), .Z(n42183) );
  NANDN U43223 ( .A(n42162), .B(n42161), .Z(n42166) );
  NANDN U43224 ( .A(n42164), .B(n42163), .Z(n42165) );
  NAND U43225 ( .A(n42166), .B(n42165), .Z(n42213) );
  XNOR U43226 ( .A(n42212), .B(n42213), .Z(n42214) );
  NAND U43227 ( .A(n42231), .B(n42167), .Z(n42170) );
  XNOR U43228 ( .A(n247), .B(n42168), .Z(n42202) );
  NANDN U43229 ( .A(n42202), .B(n42234), .Z(n42169) );
  NAND U43230 ( .A(n42170), .B(n42169), .Z(n42190) );
  NAND U43231 ( .A(n42172), .B(n42171), .Z(n42175) );
  XNOR U43232 ( .A(n42197), .B(n42233), .Z(n42198) );
  NANDN U43233 ( .A(n42198), .B(n42173), .Z(n42174) );
  AND U43234 ( .A(n42175), .B(n42174), .Z(n42191) );
  XNOR U43235 ( .A(n42190), .B(n42191), .Z(n42192) );
  NAND U43236 ( .A(b[7]), .B(a[1019]), .Z(n42207) );
  XOR U43237 ( .A(n42206), .B(n42207), .Z(n42209) );
  XOR U43238 ( .A(n42208), .B(n42209), .Z(n42193) );
  XOR U43239 ( .A(n42192), .B(n42193), .Z(n42215) );
  XOR U43240 ( .A(n42214), .B(n42215), .Z(n42184) );
  NAND U43241 ( .A(n42177), .B(n42176), .Z(n42181) );
  NANDN U43242 ( .A(n42179), .B(n42178), .Z(n42180) );
  AND U43243 ( .A(n42181), .B(n42180), .Z(n42185) );
  XNOR U43244 ( .A(n42184), .B(n42185), .Z(n42186) );
  XNOR U43245 ( .A(n42187), .B(n42186), .Z(n42182) );
  XOR U43246 ( .A(n42183), .B(n42182), .Z(c[2043]) );
  OR U43247 ( .A(n42183), .B(n42182), .Z(n42219) );
  NANDN U43248 ( .A(n42185), .B(n42184), .Z(n42189) );
  NANDN U43249 ( .A(n42187), .B(n42186), .Z(n42188) );
  NAND U43250 ( .A(n42189), .B(n42188), .Z(n42223) );
  NANDN U43251 ( .A(n42191), .B(n42190), .Z(n42195) );
  NANDN U43252 ( .A(n42193), .B(n42192), .Z(n42194) );
  NAND U43253 ( .A(n42195), .B(n42194), .Z(n42240) );
  AND U43254 ( .A(b[4]), .B(b[3]), .Z(n42196) );
  XNOR U43255 ( .A(n42197), .B(n42196), .Z(n42201) );
  XNOR U43256 ( .A(b[3]), .B(b[4]), .Z(n42199) );
  NAND U43257 ( .A(n42199), .B(n42198), .Z(n42200) );
  AND U43258 ( .A(n42201), .B(n42200), .Z(n42226) );
  ANDN U43259 ( .B(a[1020]), .A(n247), .Z(n42252) );
  XOR U43260 ( .A(n42226), .B(n42252), .Z(n42228) );
  NANDN U43261 ( .A(n42202), .B(n42231), .Z(n42205) );
  XNOR U43262 ( .A(b[7]), .B(n42203), .Z(n42232) );
  NAND U43263 ( .A(n42234), .B(n42232), .Z(n42204) );
  NAND U43264 ( .A(n42205), .B(n42204), .Z(n42227) );
  XNOR U43265 ( .A(n42228), .B(n42227), .Z(n42237) );
  NANDN U43266 ( .A(n42207), .B(n42206), .Z(n42211) );
  NANDN U43267 ( .A(n42209), .B(n42208), .Z(n42210) );
  AND U43268 ( .A(n42211), .B(n42210), .Z(n42238) );
  XNOR U43269 ( .A(n42237), .B(n42238), .Z(n42239) );
  XNOR U43270 ( .A(n42240), .B(n42239), .Z(n42220) );
  NANDN U43271 ( .A(n42213), .B(n42212), .Z(n42217) );
  NANDN U43272 ( .A(n42215), .B(n42214), .Z(n42216) );
  NAND U43273 ( .A(n42217), .B(n42216), .Z(n42221) );
  XNOR U43274 ( .A(n42220), .B(n42221), .Z(n42222) );
  XOR U43275 ( .A(n42223), .B(n42222), .Z(n42218) );
  XOR U43276 ( .A(n42219), .B(n42218), .Z(c[2044]) );
  OR U43277 ( .A(n42219), .B(n42218), .Z(n42244) );
  NANDN U43278 ( .A(n42221), .B(n42220), .Z(n42225) );
  NAND U43279 ( .A(n42223), .B(n42222), .Z(n42224) );
  NAND U43280 ( .A(n42225), .B(n42224), .Z(n42260) );
  NANDN U43281 ( .A(n42226), .B(n42252), .Z(n42230) );
  OR U43282 ( .A(n42228), .B(n42227), .Z(n42229) );
  NAND U43283 ( .A(n42230), .B(n42229), .Z(n42264) );
  NAND U43284 ( .A(n42232), .B(n42231), .Z(n42236) );
  XOR U43285 ( .A(n42233), .B(n247), .Z(n42247) );
  NAND U43286 ( .A(n42234), .B(n42247), .Z(n42235) );
  NAND U43287 ( .A(n42236), .B(n42235), .Z(n42263) );
  XNOR U43288 ( .A(n42264), .B(n42263), .Z(n42265) );
  NAND U43289 ( .A(a[1021]), .B(b[7]), .Z(n42251) );
  XNOR U43290 ( .A(n42250), .B(n42251), .Z(n42253) );
  XNOR U43291 ( .A(n42252), .B(n42253), .Z(n42266) );
  XOR U43292 ( .A(n42265), .B(n42266), .Z(n42257) );
  NANDN U43293 ( .A(n42238), .B(n42237), .Z(n42242) );
  NAND U43294 ( .A(n42240), .B(n42239), .Z(n42241) );
  NAND U43295 ( .A(n42242), .B(n42241), .Z(n42258) );
  XNOR U43296 ( .A(n42257), .B(n42258), .Z(n42259) );
  XOR U43297 ( .A(n42260), .B(n42259), .Z(n42243) );
  XOR U43298 ( .A(n42244), .B(n42243), .Z(c[2045]) );
  OR U43299 ( .A(n42244), .B(n42243), .Z(n42284) );
  ANDN U43300 ( .B(a[1022]), .A(n247), .Z(n42270) );
  AND U43301 ( .A(b[6]), .B(b[5]), .Z(n42245) );
  XNOR U43302 ( .A(n247), .B(n42245), .Z(n42249) );
  XNOR U43303 ( .A(b[6]), .B(b[5]), .Z(n42246) );
  NANDN U43304 ( .A(n42247), .B(n42246), .Z(n42248) );
  AND U43305 ( .A(n42249), .B(n42248), .Z(n42269) );
  NANDN U43306 ( .A(n42251), .B(n42250), .Z(n42255) );
  NAND U43307 ( .A(n42253), .B(n42252), .Z(n42254) );
  NAND U43308 ( .A(n42255), .B(n42254), .Z(n42256) );
  XNOR U43309 ( .A(n42269), .B(n42256), .Z(n42271) );
  XNOR U43310 ( .A(n42270), .B(n42271), .Z(n42280) );
  NANDN U43311 ( .A(n42258), .B(n42257), .Z(n42262) );
  NAND U43312 ( .A(n42260), .B(n42259), .Z(n42261) );
  NAND U43313 ( .A(n42262), .B(n42261), .Z(n42277) );
  NANDN U43314 ( .A(n42264), .B(n42263), .Z(n42268) );
  NANDN U43315 ( .A(n42266), .B(n42265), .Z(n42267) );
  AND U43316 ( .A(n42268), .B(n42267), .Z(n42278) );
  XOR U43317 ( .A(n42277), .B(n42278), .Z(n42279) );
  XOR U43318 ( .A(n42280), .B(n42279), .Z(n42283) );
  XOR U43319 ( .A(n42284), .B(n42283), .Z(c[2046]) );
  XNOR U43320 ( .A(n42270), .B(n42269), .Z(n42272) );
  NAND U43321 ( .A(n42272), .B(n42271), .Z(n42276) );
  XNOR U43322 ( .A(a[1023]), .B(n42273), .Z(n42274) );
  AND U43323 ( .A(n42274), .B(b[7]), .Z(n42275) );
  XNOR U43324 ( .A(n42276), .B(n42275), .Z(n42288) );
  AND U43325 ( .A(n42278), .B(n42277), .Z(n42282) );
  AND U43326 ( .A(n42280), .B(n42279), .Z(n42281) );
  OR U43327 ( .A(n42282), .B(n42281), .Z(n42286) );
  OR U43328 ( .A(n42284), .B(n42283), .Z(n42285) );
  NAND U43329 ( .A(n42286), .B(n42285), .Z(n42287) );
  XOR U43330 ( .A(n42288), .B(n42287), .Z(c[2047]) );
endmodule

