
module hamming_N1600_CC8 ( clk, rst, x, y, o );
  input [199:0] x;
  input [199:0] y;
  output [10:0] o;
  input clk, rst;
  wire   n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029;
  wire   [10:0] oglobal;

  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[0]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[1]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[2]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[3]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[4]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[5]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[6]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[7]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[8]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[9]) );
  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[10]) );
  XNOR U214 ( .A(n328), .B(n329), .Z(n341) );
  XNOR U215 ( .A(n309), .B(n560), .Z(n315) );
  XNOR U216 ( .A(n359), .B(n636), .Z(n365) );
  XNOR U217 ( .A(n377), .B(n378), .Z(n390) );
  XNOR U218 ( .A(n218), .B(n219), .Z(n227) );
  XNOR U219 ( .A(n291), .B(n503), .Z(n274) );
  XNOR U220 ( .A(n411), .B(n413), .Z(n432) );
  XNOR U221 ( .A(n148), .B(n245), .Z(n131) );
  XNOR U222 ( .A(n34), .B(n47), .Z(n36) );
  XNOR U223 ( .A(n181), .B(n293), .Z(n155) );
  XNOR U224 ( .A(n261), .B(n484), .Z(n267) );
  XNOR U225 ( .A(n110), .B(n112), .Z(n124) );
  XNOR U226 ( .A(n487), .B(n489), .Z(n508) );
  XNOR U227 ( .A(n639), .B(n641), .Z(n660) );
  XNOR U228 ( .A(n96), .B(n176), .Z(n102) );
  XNOR U229 ( .A(n226), .B(n227), .Z(n251) );
  XNOR U230 ( .A(n430), .B(n432), .Z(n470) );
  XNOR U231 ( .A(n582), .B(n584), .Z(n622) );
  XNOR U232 ( .A(n51), .B(n80), .Z(n57) );
  XNOR U233 ( .A(n348), .B(n541), .Z(n298) );
  XOR U234 ( .A(oglobal[7]), .B(n31), .Z(n12) );
  XOR U235 ( .A(oglobal[4]), .B(n105), .Z(n18) );
  ANDN U236 ( .B(n1009), .A(n680), .Z(n682) );
  XNOR U237 ( .A(n134), .B(n257), .Z(n136) );
  XNOR U238 ( .A(n353), .B(n354), .Z(n366) );
  XNOR U239 ( .A(n997), .B(n996), .Z(n1016) );
  XNOR U240 ( .A(n976), .B(n975), .Z(n973) );
  XNOR U241 ( .A(n934), .B(n933), .Z(n931) );
  XNOR U242 ( .A(n892), .B(n891), .Z(n889) );
  XNOR U243 ( .A(n852), .B(n851), .Z(n849) );
  XNOR U244 ( .A(n808), .B(n807), .Z(n805) );
  XNOR U245 ( .A(n768), .B(n767), .Z(n765) );
  XNOR U246 ( .A(n726), .B(n725), .Z(n723) );
  XNOR U247 ( .A(n142), .B(n269), .Z(n148) );
  XNOR U248 ( .A(n243), .B(n427), .Z(n226) );
  XNOR U249 ( .A(n389), .B(n655), .Z(n372) );
  XNOR U250 ( .A(n563), .B(n565), .Z(n584) );
  XNOR U251 ( .A(n65), .B(n67), .Z(n79) );
  XNOR U252 ( .A(n123), .B(n124), .Z(n132) );
  XNOR U253 ( .A(n274), .B(n465), .Z(n250) );
  XNOR U254 ( .A(n323), .B(n324), .Z(n349) );
  XNOR U255 ( .A(n658), .B(n945), .Z(n620) );
  XNOR U256 ( .A(n102), .B(n150), .Z(n85) );
  XNOR U257 ( .A(n468), .B(n470), .Z(n546) );
  XOR U258 ( .A(oglobal[6]), .B(n39), .Z(n14) );
  XOR U259 ( .A(oglobal[3]), .B(n201), .Z(n20) );
  ANDN U260 ( .B(n841), .A(n528), .Z(n530) );
  ANDN U261 ( .B(n923), .A(n604), .Z(n606) );
  XNOR U262 ( .A(n184), .B(n355), .Z(n186) );
  XNOR U263 ( .A(n237), .B(n446), .Z(n243) );
  XNOR U264 ( .A(n255), .B(n256), .Z(n268) );
  XNOR U265 ( .A(n279), .B(n280), .Z(n292) );
  XNOR U266 ( .A(n303), .B(n304), .Z(n316) );
  XNOR U267 ( .A(n1020), .B(n1019), .Z(n1017) );
  XNOR U268 ( .A(n955), .B(n954), .Z(n972) );
  XNOR U269 ( .A(n911), .B(n910), .Z(n930) );
  XNOR U270 ( .A(n871), .B(n870), .Z(n888) );
  XNOR U271 ( .A(n829), .B(n828), .Z(n848) );
  XNOR U272 ( .A(n787), .B(n786), .Z(n804) );
  XNOR U273 ( .A(n192), .B(n367), .Z(n198) );
  XNOR U274 ( .A(n340), .B(n579), .Z(n323) );
  XNOR U275 ( .A(n449), .B(n735), .Z(n430) );
  XNOR U276 ( .A(n90), .B(n91), .Z(n103) );
  XNOR U277 ( .A(n174), .B(n175), .Z(n182) );
  XNOR U278 ( .A(n372), .B(n617), .Z(n348) );
  XNOR U279 ( .A(n506), .B(n777), .Z(n468) );
  XNOR U280 ( .A(n44), .B(n46), .Z(n58) );
  XNOR U281 ( .A(n78), .B(n79), .Z(n86) );
  XNOR U282 ( .A(n131), .B(n132), .Z(n156) );
  XNOR U283 ( .A(n250), .B(n251), .Z(n299) );
  XNOR U284 ( .A(n620), .B(n861), .Z(n544) );
  XOR U285 ( .A(oglobal[5]), .B(n60), .Z(n16) );
  XOR U286 ( .A(oglobal[2]), .B(n392), .Z(n22) );
  ANDN U287 ( .B(n715), .A(n414), .Z(n416) );
  ANDN U288 ( .B(n757), .A(n452), .Z(n454) );
  ANDN U289 ( .B(n797), .A(n490), .Z(n492) );
  ANDN U290 ( .B(n881), .A(n566), .Z(n568) );
  ANDN U291 ( .B(n965), .A(n642), .Z(n644) );
  XNOR U292 ( .A(n206), .B(n207), .Z(n219) );
  XNOR U293 ( .A(n231), .B(n232), .Z(n244) );
  XNOR U294 ( .A(n285), .B(n522), .Z(n291) );
  XNOR U295 ( .A(n334), .B(n598), .Z(n340) );
  XNOR U296 ( .A(n383), .B(n674), .Z(n389) );
  XNOR U297 ( .A(n745), .B(n744), .Z(n764) );
  XNOR U298 ( .A(n705), .B(n704), .Z(n722) );
  XNOR U299 ( .A(n136), .B(n137), .Z(n149) );
  XNOR U300 ( .A(n160), .B(n162), .Z(n175) );
  XNOR U301 ( .A(n186), .B(n187), .Z(n199) );
  XNOR U302 ( .A(n267), .B(n268), .Z(n275) );
  XNOR U303 ( .A(n315), .B(n316), .Z(n324) );
  XNOR U304 ( .A(n365), .B(n366), .Z(n373) );
  XNOR U305 ( .A(n525), .B(n819), .Z(n506) );
  XNOR U306 ( .A(n601), .B(n901), .Z(n582) );
  XNOR U307 ( .A(n677), .B(n987), .Z(n658) );
  XNOR U308 ( .A(n36), .B(n37), .Z(n15) );
  XNOR U309 ( .A(n57), .B(n58), .Z(n17) );
  XNOR U310 ( .A(n85), .B(n86), .Z(n19) );
  XNOR U311 ( .A(n155), .B(n156), .Z(n21) );
  XNOR U312 ( .A(n298), .B(n299), .Z(n23) );
  XNOR U313 ( .A(n544), .B(n546), .Z(n25) );
  XNOR U314 ( .A(n12), .B(n13), .Z(o[7]) );
  XOR U315 ( .A(n14), .B(n15), .Z(o[6]) );
  XOR U316 ( .A(n16), .B(n17), .Z(o[5]) );
  XOR U317 ( .A(n18), .B(n19), .Z(o[4]) );
  XOR U318 ( .A(n20), .B(n21), .Z(o[3]) );
  XOR U319 ( .A(n22), .B(n23), .Z(o[2]) );
  XOR U320 ( .A(n24), .B(n25), .Z(o[1]) );
  XOR U321 ( .A(n26), .B(n27), .Z(o[10]) );
  XOR U322 ( .A(oglobal[10]), .B(n28), .Z(n27) );
  AND U323 ( .A(n26), .B(o[9]), .Z(n28) );
  XOR U324 ( .A(oglobal[9]), .B(n26), .Z(o[9]) );
  ANDN U325 ( .B(n29), .A(o[8]), .Z(n26) );
  XOR U326 ( .A(oglobal[8]), .B(n29), .Z(o[8]) );
  XNOR U327 ( .A(n30), .B(n31), .Z(n29) );
  ANDN U328 ( .B(n32), .A(n12), .Z(n30) );
  XNOR U329 ( .A(n31), .B(n13), .Z(n32) );
  XNOR U330 ( .A(n33), .B(n34), .Z(n13) );
  ANDN U331 ( .B(n35), .A(n36), .Z(n33) );
  XOR U332 ( .A(n34), .B(n37), .Z(n35) );
  XOR U333 ( .A(n38), .B(n39), .Z(n31) );
  ANDN U334 ( .B(n40), .A(n14), .Z(n38) );
  XOR U335 ( .A(n39), .B(n15), .Z(n40) );
  XNOR U336 ( .A(n41), .B(n42), .Z(n37) );
  ANDN U337 ( .B(n43), .A(n44), .Z(n41) );
  XOR U338 ( .A(n45), .B(n46), .Z(n43) );
  XNOR U339 ( .A(n48), .B(n49), .Z(n47) );
  ANDN U340 ( .B(n50), .A(n51), .Z(n48) );
  XNOR U341 ( .A(n52), .B(n53), .Z(n50) );
  XOR U342 ( .A(n54), .B(n55), .Z(n34) );
  ANDN U343 ( .B(n56), .A(n57), .Z(n54) );
  XOR U344 ( .A(n55), .B(n58), .Z(n56) );
  XOR U345 ( .A(n59), .B(n60), .Z(n39) );
  ANDN U346 ( .B(n61), .A(n16), .Z(n59) );
  XOR U347 ( .A(n60), .B(n17), .Z(n61) );
  XNOR U348 ( .A(n62), .B(n63), .Z(n46) );
  ANDN U349 ( .B(n64), .A(n65), .Z(n62) );
  XOR U350 ( .A(n66), .B(n67), .Z(n64) );
  XOR U351 ( .A(n42), .B(n68), .Z(n44) );
  XNOR U352 ( .A(n69), .B(n70), .Z(n68) );
  ANDN U353 ( .B(n71), .A(n72), .Z(n69) );
  XNOR U354 ( .A(n73), .B(n74), .Z(n71) );
  IV U355 ( .A(n45), .Z(n42) );
  XOR U356 ( .A(n75), .B(n76), .Z(n45) );
  ANDN U357 ( .B(n77), .A(n78), .Z(n75) );
  XOR U358 ( .A(n76), .B(n79), .Z(n77) );
  XNOR U359 ( .A(n52), .B(n81), .Z(n80) );
  IV U360 ( .A(n55), .Z(n81) );
  XOR U361 ( .A(n82), .B(n83), .Z(n55) );
  ANDN U362 ( .B(n84), .A(n85), .Z(n82) );
  XOR U363 ( .A(n83), .B(n86), .Z(n84) );
  XNOR U364 ( .A(n87), .B(n88), .Z(n52) );
  ANDN U365 ( .B(n89), .A(n90), .Z(n87) );
  XOR U366 ( .A(n88), .B(n91), .Z(n89) );
  XOR U367 ( .A(n49), .B(n92), .Z(n51) );
  XNOR U368 ( .A(n93), .B(n94), .Z(n92) );
  ANDN U369 ( .B(n95), .A(n96), .Z(n93) );
  XNOR U370 ( .A(n97), .B(n98), .Z(n95) );
  IV U371 ( .A(n53), .Z(n49) );
  XOR U372 ( .A(n99), .B(n100), .Z(n53) );
  ANDN U373 ( .B(n101), .A(n102), .Z(n99) );
  XOR U374 ( .A(n103), .B(n100), .Z(n101) );
  XOR U375 ( .A(n104), .B(n105), .Z(n60) );
  ANDN U376 ( .B(n106), .A(n18), .Z(n104) );
  XOR U377 ( .A(n105), .B(n19), .Z(n106) );
  XNOR U378 ( .A(n107), .B(n108), .Z(n67) );
  ANDN U379 ( .B(n109), .A(n110), .Z(n107) );
  XOR U380 ( .A(n111), .B(n112), .Z(n109) );
  XOR U381 ( .A(n63), .B(n113), .Z(n65) );
  XNOR U382 ( .A(n114), .B(n115), .Z(n113) );
  ANDN U383 ( .B(n116), .A(n117), .Z(n114) );
  XNOR U384 ( .A(n118), .B(n119), .Z(n116) );
  IV U385 ( .A(n66), .Z(n63) );
  XOR U386 ( .A(n120), .B(n121), .Z(n66) );
  ANDN U387 ( .B(n122), .A(n123), .Z(n120) );
  XOR U388 ( .A(n121), .B(n124), .Z(n122) );
  XOR U389 ( .A(n125), .B(n126), .Z(n78) );
  XNOR U390 ( .A(n73), .B(n127), .Z(n126) );
  IV U391 ( .A(n76), .Z(n127) );
  XOR U392 ( .A(n128), .B(n129), .Z(n76) );
  ANDN U393 ( .B(n130), .A(n131), .Z(n128) );
  XOR U394 ( .A(n129), .B(n132), .Z(n130) );
  XNOR U395 ( .A(n133), .B(n134), .Z(n73) );
  ANDN U396 ( .B(n135), .A(n136), .Z(n133) );
  XOR U397 ( .A(n134), .B(n137), .Z(n135) );
  IV U398 ( .A(n72), .Z(n125) );
  XOR U399 ( .A(n70), .B(n138), .Z(n72) );
  XNOR U400 ( .A(n139), .B(n140), .Z(n138) );
  ANDN U401 ( .B(n141), .A(n142), .Z(n139) );
  XNOR U402 ( .A(n143), .B(n144), .Z(n141) );
  IV U403 ( .A(n74), .Z(n70) );
  XOR U404 ( .A(n145), .B(n146), .Z(n74) );
  ANDN U405 ( .B(n147), .A(n148), .Z(n145) );
  XOR U406 ( .A(n149), .B(n146), .Z(n147) );
  XOR U407 ( .A(n103), .B(n151), .Z(n150) );
  IV U408 ( .A(n83), .Z(n151) );
  XOR U409 ( .A(n152), .B(n153), .Z(n83) );
  ANDN U410 ( .B(n154), .A(n155), .Z(n152) );
  XOR U411 ( .A(n153), .B(n156), .Z(n154) );
  XNOR U412 ( .A(n157), .B(n158), .Z(n91) );
  ANDN U413 ( .B(n159), .A(n160), .Z(n157) );
  XOR U414 ( .A(n161), .B(n162), .Z(n159) );
  XOR U415 ( .A(n163), .B(n164), .Z(n90) );
  XNOR U416 ( .A(n165), .B(n166), .Z(n164) );
  ANDN U417 ( .B(n167), .A(n168), .Z(n165) );
  XNOR U418 ( .A(n169), .B(n170), .Z(n167) );
  IV U419 ( .A(n88), .Z(n163) );
  XOR U420 ( .A(n171), .B(n172), .Z(n88) );
  ANDN U421 ( .B(n173), .A(n174), .Z(n171) );
  XOR U422 ( .A(n172), .B(n175), .Z(n173) );
  XNOR U423 ( .A(n97), .B(n177), .Z(n176) );
  IV U424 ( .A(n100), .Z(n177) );
  XOR U425 ( .A(n178), .B(n179), .Z(n100) );
  ANDN U426 ( .B(n180), .A(n181), .Z(n178) );
  XOR U427 ( .A(n182), .B(n179), .Z(n180) );
  XNOR U428 ( .A(n183), .B(n184), .Z(n97) );
  ANDN U429 ( .B(n185), .A(n186), .Z(n183) );
  XOR U430 ( .A(n184), .B(n187), .Z(n185) );
  XOR U431 ( .A(n94), .B(n188), .Z(n96) );
  XNOR U432 ( .A(n189), .B(n190), .Z(n188) );
  ANDN U433 ( .B(n191), .A(n192), .Z(n189) );
  XNOR U434 ( .A(n193), .B(n194), .Z(n191) );
  IV U435 ( .A(n98), .Z(n94) );
  XOR U436 ( .A(n195), .B(n196), .Z(n98) );
  ANDN U437 ( .B(n197), .A(n198), .Z(n195) );
  XOR U438 ( .A(n199), .B(n196), .Z(n197) );
  XOR U439 ( .A(n200), .B(n201), .Z(n105) );
  ANDN U440 ( .B(n202), .A(n20), .Z(n200) );
  XOR U441 ( .A(n201), .B(n21), .Z(n202) );
  XNOR U442 ( .A(n203), .B(n204), .Z(n112) );
  ANDN U443 ( .B(n205), .A(n206), .Z(n203) );
  XNOR U444 ( .A(n204), .B(n207), .Z(n205) );
  XOR U445 ( .A(n108), .B(n208), .Z(n110) );
  XNOR U446 ( .A(n209), .B(n210), .Z(n208) );
  ANDN U447 ( .B(n211), .A(n212), .Z(n209) );
  XNOR U448 ( .A(n213), .B(n214), .Z(n211) );
  IV U449 ( .A(n111), .Z(n108) );
  XOR U450 ( .A(n215), .B(n216), .Z(n111) );
  ANDN U451 ( .B(n217), .A(n218), .Z(n215) );
  XOR U452 ( .A(n216), .B(n219), .Z(n217) );
  XOR U453 ( .A(n220), .B(n221), .Z(n123) );
  XNOR U454 ( .A(n118), .B(n222), .Z(n221) );
  IV U455 ( .A(n121), .Z(n222) );
  XOR U456 ( .A(n223), .B(n224), .Z(n121) );
  ANDN U457 ( .B(n225), .A(n226), .Z(n223) );
  XOR U458 ( .A(n224), .B(n227), .Z(n225) );
  XOR U459 ( .A(n228), .B(n229), .Z(n118) );
  ANDN U460 ( .B(n230), .A(n231), .Z(n228) );
  XNOR U461 ( .A(n229), .B(n232), .Z(n230) );
  IV U462 ( .A(n117), .Z(n220) );
  XOR U463 ( .A(n115), .B(n233), .Z(n117) );
  XNOR U464 ( .A(n234), .B(n235), .Z(n233) );
  ANDN U465 ( .B(n236), .A(n237), .Z(n234) );
  XNOR U466 ( .A(n238), .B(n239), .Z(n236) );
  IV U467 ( .A(n119), .Z(n115) );
  XOR U468 ( .A(n240), .B(n241), .Z(n119) );
  ANDN U469 ( .B(n242), .A(n243), .Z(n240) );
  XOR U470 ( .A(n244), .B(n241), .Z(n242) );
  XOR U471 ( .A(n149), .B(n246), .Z(n245) );
  IV U472 ( .A(n129), .Z(n246) );
  XOR U473 ( .A(n247), .B(n248), .Z(n129) );
  ANDN U474 ( .B(n249), .A(n250), .Z(n247) );
  XOR U475 ( .A(n248), .B(n251), .Z(n249) );
  XNOR U476 ( .A(n252), .B(n253), .Z(n137) );
  ANDN U477 ( .B(n254), .A(n255), .Z(n252) );
  XNOR U478 ( .A(n253), .B(n256), .Z(n254) );
  XNOR U479 ( .A(n258), .B(n259), .Z(n257) );
  ANDN U480 ( .B(n260), .A(n261), .Z(n258) );
  XNOR U481 ( .A(n262), .B(n263), .Z(n260) );
  XOR U482 ( .A(n264), .B(n265), .Z(n134) );
  ANDN U483 ( .B(n266), .A(n267), .Z(n264) );
  XOR U484 ( .A(n265), .B(n268), .Z(n266) );
  XNOR U485 ( .A(n143), .B(n270), .Z(n269) );
  IV U486 ( .A(n146), .Z(n270) );
  XOR U487 ( .A(n271), .B(n272), .Z(n146) );
  ANDN U488 ( .B(n273), .A(n274), .Z(n271) );
  XOR U489 ( .A(n275), .B(n272), .Z(n273) );
  XOR U490 ( .A(n276), .B(n277), .Z(n143) );
  ANDN U491 ( .B(n278), .A(n279), .Z(n276) );
  XNOR U492 ( .A(n277), .B(n280), .Z(n278) );
  XOR U493 ( .A(n140), .B(n281), .Z(n142) );
  XNOR U494 ( .A(n282), .B(n283), .Z(n281) );
  ANDN U495 ( .B(n284), .A(n285), .Z(n282) );
  XNOR U496 ( .A(n286), .B(n287), .Z(n284) );
  IV U497 ( .A(n144), .Z(n140) );
  XOR U498 ( .A(n288), .B(n289), .Z(n144) );
  ANDN U499 ( .B(n290), .A(n291), .Z(n288) );
  XOR U500 ( .A(n292), .B(n289), .Z(n290) );
  XOR U501 ( .A(n182), .B(n294), .Z(n293) );
  IV U502 ( .A(n153), .Z(n294) );
  XOR U503 ( .A(n295), .B(n296), .Z(n153) );
  ANDN U504 ( .B(n297), .A(n298), .Z(n295) );
  XOR U505 ( .A(n296), .B(n299), .Z(n297) );
  XNOR U506 ( .A(n300), .B(n301), .Z(n162) );
  ANDN U507 ( .B(n302), .A(n303), .Z(n300) );
  XNOR U508 ( .A(n301), .B(n304), .Z(n302) );
  XOR U509 ( .A(n158), .B(n305), .Z(n160) );
  XNOR U510 ( .A(n306), .B(n307), .Z(n305) );
  ANDN U511 ( .B(n308), .A(n309), .Z(n306) );
  XNOR U512 ( .A(n310), .B(n311), .Z(n308) );
  IV U513 ( .A(n161), .Z(n158) );
  XOR U514 ( .A(n312), .B(n313), .Z(n161) );
  ANDN U515 ( .B(n314), .A(n315), .Z(n312) );
  XOR U516 ( .A(n313), .B(n316), .Z(n314) );
  XOR U517 ( .A(n317), .B(n318), .Z(n174) );
  XNOR U518 ( .A(n169), .B(n319), .Z(n318) );
  IV U519 ( .A(n172), .Z(n319) );
  XOR U520 ( .A(n320), .B(n321), .Z(n172) );
  ANDN U521 ( .B(n322), .A(n323), .Z(n320) );
  XOR U522 ( .A(n321), .B(n324), .Z(n322) );
  XOR U523 ( .A(n325), .B(n326), .Z(n169) );
  ANDN U524 ( .B(n327), .A(n328), .Z(n325) );
  XNOR U525 ( .A(n326), .B(n329), .Z(n327) );
  IV U526 ( .A(n168), .Z(n317) );
  XOR U527 ( .A(n166), .B(n330), .Z(n168) );
  XNOR U528 ( .A(n331), .B(n332), .Z(n330) );
  ANDN U529 ( .B(n333), .A(n334), .Z(n331) );
  XNOR U530 ( .A(n335), .B(n336), .Z(n333) );
  IV U531 ( .A(n170), .Z(n166) );
  XOR U532 ( .A(n337), .B(n338), .Z(n170) );
  ANDN U533 ( .B(n339), .A(n340), .Z(n337) );
  XOR U534 ( .A(n341), .B(n338), .Z(n339) );
  XOR U535 ( .A(n342), .B(n343), .Z(n181) );
  XOR U536 ( .A(n199), .B(n344), .Z(n343) );
  IV U537 ( .A(n179), .Z(n344) );
  XOR U538 ( .A(n345), .B(n346), .Z(n179) );
  ANDN U539 ( .B(n347), .A(n348), .Z(n345) );
  XOR U540 ( .A(n349), .B(n346), .Z(n347) );
  XNOR U541 ( .A(n350), .B(n351), .Z(n187) );
  ANDN U542 ( .B(n352), .A(n353), .Z(n350) );
  XNOR U543 ( .A(n351), .B(n354), .Z(n352) );
  XNOR U544 ( .A(n356), .B(n357), .Z(n355) );
  ANDN U545 ( .B(n358), .A(n359), .Z(n356) );
  XNOR U546 ( .A(n360), .B(n361), .Z(n358) );
  XOR U547 ( .A(n362), .B(n363), .Z(n184) );
  ANDN U548 ( .B(n364), .A(n365), .Z(n362) );
  XOR U549 ( .A(n363), .B(n366), .Z(n364) );
  IV U550 ( .A(n198), .Z(n342) );
  XNOR U551 ( .A(n193), .B(n368), .Z(n367) );
  IV U552 ( .A(n196), .Z(n368) );
  XOR U553 ( .A(n369), .B(n370), .Z(n196) );
  ANDN U554 ( .B(n371), .A(n372), .Z(n369) );
  XOR U555 ( .A(n373), .B(n370), .Z(n371) );
  XOR U556 ( .A(n374), .B(n375), .Z(n193) );
  ANDN U557 ( .B(n376), .A(n377), .Z(n374) );
  XNOR U558 ( .A(n375), .B(n378), .Z(n376) );
  XOR U559 ( .A(n190), .B(n379), .Z(n192) );
  XNOR U560 ( .A(n380), .B(n381), .Z(n379) );
  ANDN U561 ( .B(n382), .A(n383), .Z(n380) );
  XNOR U562 ( .A(n384), .B(n385), .Z(n382) );
  IV U563 ( .A(n194), .Z(n190) );
  XOR U564 ( .A(n386), .B(n387), .Z(n194) );
  ANDN U565 ( .B(n388), .A(n389), .Z(n386) );
  XOR U566 ( .A(n390), .B(n387), .Z(n388) );
  XOR U567 ( .A(n391), .B(n392), .Z(n201) );
  ANDN U568 ( .B(n393), .A(n22), .Z(n391) );
  XOR U569 ( .A(n392), .B(n23), .Z(n393) );
  XNOR U570 ( .A(n394), .B(n395), .Z(n207) );
  NANDN U571 ( .A(n396), .B(n397), .Z(n395) );
  NANDN U572 ( .A(n398), .B(n394), .Z(n397) );
  XNOR U573 ( .A(n399), .B(n204), .Z(n206) );
  XNOR U574 ( .A(n400), .B(n401), .Z(n204) );
  NAND U575 ( .A(n402), .B(n403), .Z(n401) );
  XNOR U576 ( .A(n400), .B(n404), .Z(n402) );
  NOR U577 ( .A(n405), .B(n406), .Z(n399) );
  XOR U578 ( .A(n407), .B(n408), .Z(n218) );
  XOR U579 ( .A(n213), .B(n216), .Z(n408) );
  XNOR U580 ( .A(n409), .B(n410), .Z(n216) );
  NANDN U581 ( .A(n411), .B(n412), .Z(n410) );
  XOR U582 ( .A(n409), .B(n413), .Z(n412) );
  XNOR U583 ( .A(n414), .B(n415), .Z(n213) );
  NANDN U584 ( .A(n416), .B(n417), .Z(n415) );
  NANDN U585 ( .A(n414), .B(n418), .Z(n417) );
  IV U586 ( .A(n212), .Z(n407) );
  XOR U587 ( .A(n419), .B(n214), .Z(n212) );
  IV U588 ( .A(n210), .Z(n214) );
  XNOR U589 ( .A(n420), .B(n421), .Z(n210) );
  NAND U590 ( .A(n422), .B(n423), .Z(n421) );
  XOR U591 ( .A(n420), .B(n424), .Z(n422) );
  NOR U592 ( .A(n425), .B(n426), .Z(n419) );
  XNOR U593 ( .A(n244), .B(n224), .Z(n427) );
  XNOR U594 ( .A(n428), .B(n429), .Z(n224) );
  NANDN U595 ( .A(n430), .B(n431), .Z(n429) );
  XOR U596 ( .A(n428), .B(n432), .Z(n431) );
  XNOR U597 ( .A(n433), .B(n434), .Z(n232) );
  NANDN U598 ( .A(n435), .B(n436), .Z(n434) );
  NANDN U599 ( .A(n437), .B(n433), .Z(n436) );
  XNOR U600 ( .A(n438), .B(n229), .Z(n231) );
  XNOR U601 ( .A(n439), .B(n440), .Z(n229) );
  NAND U602 ( .A(n441), .B(n442), .Z(n440) );
  XNOR U603 ( .A(n439), .B(n443), .Z(n441) );
  NOR U604 ( .A(n444), .B(n445), .Z(n438) );
  XOR U605 ( .A(n238), .B(n241), .Z(n446) );
  XNOR U606 ( .A(n447), .B(n448), .Z(n241) );
  NANDN U607 ( .A(n449), .B(n450), .Z(n448) );
  XNOR U608 ( .A(n447), .B(n451), .Z(n450) );
  XNOR U609 ( .A(n452), .B(n453), .Z(n238) );
  NANDN U610 ( .A(n454), .B(n455), .Z(n453) );
  NANDN U611 ( .A(n452), .B(n456), .Z(n455) );
  XOR U612 ( .A(n457), .B(n239), .Z(n237) );
  IV U613 ( .A(n235), .Z(n239) );
  XNOR U614 ( .A(n458), .B(n459), .Z(n235) );
  NAND U615 ( .A(n460), .B(n461), .Z(n459) );
  XOR U616 ( .A(n458), .B(n462), .Z(n460) );
  NOR U617 ( .A(n463), .B(n464), .Z(n457) );
  XNOR U618 ( .A(n275), .B(n248), .Z(n465) );
  XNOR U619 ( .A(n466), .B(n467), .Z(n248) );
  NANDN U620 ( .A(n468), .B(n469), .Z(n467) );
  XOR U621 ( .A(n466), .B(n470), .Z(n469) );
  XNOR U622 ( .A(n471), .B(n472), .Z(n256) );
  NANDN U623 ( .A(n473), .B(n474), .Z(n472) );
  NANDN U624 ( .A(n475), .B(n471), .Z(n474) );
  XNOR U625 ( .A(n476), .B(n253), .Z(n255) );
  XNOR U626 ( .A(n477), .B(n478), .Z(n253) );
  NAND U627 ( .A(n479), .B(n480), .Z(n478) );
  XNOR U628 ( .A(n477), .B(n481), .Z(n479) );
  NOR U629 ( .A(n482), .B(n483), .Z(n476) );
  XOR U630 ( .A(n262), .B(n265), .Z(n484) );
  XNOR U631 ( .A(n485), .B(n486), .Z(n265) );
  NANDN U632 ( .A(n487), .B(n488), .Z(n486) );
  XOR U633 ( .A(n485), .B(n489), .Z(n488) );
  XNOR U634 ( .A(n490), .B(n491), .Z(n262) );
  NANDN U635 ( .A(n492), .B(n493), .Z(n491) );
  NANDN U636 ( .A(n490), .B(n494), .Z(n493) );
  XOR U637 ( .A(n495), .B(n263), .Z(n261) );
  IV U638 ( .A(n259), .Z(n263) );
  XNOR U639 ( .A(n496), .B(n497), .Z(n259) );
  NAND U640 ( .A(n498), .B(n499), .Z(n497) );
  XOR U641 ( .A(n496), .B(n500), .Z(n498) );
  NOR U642 ( .A(n501), .B(n502), .Z(n495) );
  XNOR U643 ( .A(n292), .B(n272), .Z(n503) );
  XNOR U644 ( .A(n504), .B(n505), .Z(n272) );
  NANDN U645 ( .A(n506), .B(n507), .Z(n505) );
  XOR U646 ( .A(n504), .B(n508), .Z(n507) );
  XNOR U647 ( .A(n509), .B(n510), .Z(n280) );
  NANDN U648 ( .A(n511), .B(n512), .Z(n510) );
  NANDN U649 ( .A(n513), .B(n509), .Z(n512) );
  XNOR U650 ( .A(n514), .B(n277), .Z(n279) );
  XNOR U651 ( .A(n515), .B(n516), .Z(n277) );
  NAND U652 ( .A(n517), .B(n518), .Z(n516) );
  XNOR U653 ( .A(n515), .B(n519), .Z(n517) );
  NOR U654 ( .A(n520), .B(n521), .Z(n514) );
  XOR U655 ( .A(n286), .B(n289), .Z(n522) );
  XNOR U656 ( .A(n523), .B(n524), .Z(n289) );
  NANDN U657 ( .A(n525), .B(n526), .Z(n524) );
  XNOR U658 ( .A(n523), .B(n527), .Z(n526) );
  XNOR U659 ( .A(n528), .B(n529), .Z(n286) );
  NANDN U660 ( .A(n530), .B(n531), .Z(n529) );
  NANDN U661 ( .A(n528), .B(n532), .Z(n531) );
  XOR U662 ( .A(n533), .B(n287), .Z(n285) );
  IV U663 ( .A(n283), .Z(n287) );
  XNOR U664 ( .A(n534), .B(n535), .Z(n283) );
  NAND U665 ( .A(n536), .B(n537), .Z(n535) );
  XOR U666 ( .A(n534), .B(n538), .Z(n536) );
  NOR U667 ( .A(n539), .B(n540), .Z(n533) );
  XNOR U668 ( .A(n349), .B(n296), .Z(n541) );
  XNOR U669 ( .A(n542), .B(n543), .Z(n296) );
  NANDN U670 ( .A(n544), .B(n545), .Z(n543) );
  XOR U671 ( .A(n542), .B(n546), .Z(n545) );
  XNOR U672 ( .A(n547), .B(n548), .Z(n304) );
  NANDN U673 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U674 ( .A(n551), .B(n547), .Z(n550) );
  XNOR U675 ( .A(n552), .B(n301), .Z(n303) );
  XNOR U676 ( .A(n553), .B(n554), .Z(n301) );
  NAND U677 ( .A(n555), .B(n556), .Z(n554) );
  XNOR U678 ( .A(n553), .B(n557), .Z(n555) );
  NOR U679 ( .A(n558), .B(n559), .Z(n552) );
  XOR U680 ( .A(n310), .B(n313), .Z(n560) );
  XNOR U681 ( .A(n561), .B(n562), .Z(n313) );
  NANDN U682 ( .A(n563), .B(n564), .Z(n562) );
  XOR U683 ( .A(n561), .B(n565), .Z(n564) );
  XNOR U684 ( .A(n566), .B(n567), .Z(n310) );
  NANDN U685 ( .A(n568), .B(n569), .Z(n567) );
  NANDN U686 ( .A(n566), .B(n570), .Z(n569) );
  XOR U687 ( .A(n571), .B(n311), .Z(n309) );
  IV U688 ( .A(n307), .Z(n311) );
  XNOR U689 ( .A(n572), .B(n573), .Z(n307) );
  NAND U690 ( .A(n574), .B(n575), .Z(n573) );
  XOR U691 ( .A(n572), .B(n576), .Z(n574) );
  NOR U692 ( .A(n577), .B(n578), .Z(n571) );
  XNOR U693 ( .A(n341), .B(n321), .Z(n579) );
  XNOR U694 ( .A(n580), .B(n581), .Z(n321) );
  NANDN U695 ( .A(n582), .B(n583), .Z(n581) );
  XOR U696 ( .A(n580), .B(n584), .Z(n583) );
  XNOR U697 ( .A(n585), .B(n586), .Z(n329) );
  NANDN U698 ( .A(n587), .B(n588), .Z(n586) );
  NANDN U699 ( .A(n589), .B(n585), .Z(n588) );
  XNOR U700 ( .A(n590), .B(n326), .Z(n328) );
  XNOR U701 ( .A(n591), .B(n592), .Z(n326) );
  NAND U702 ( .A(n593), .B(n594), .Z(n592) );
  XNOR U703 ( .A(n591), .B(n595), .Z(n593) );
  NOR U704 ( .A(n596), .B(n597), .Z(n590) );
  XOR U705 ( .A(n335), .B(n338), .Z(n598) );
  XNOR U706 ( .A(n599), .B(n600), .Z(n338) );
  NANDN U707 ( .A(n601), .B(n602), .Z(n600) );
  XNOR U708 ( .A(n599), .B(n603), .Z(n602) );
  XNOR U709 ( .A(n604), .B(n605), .Z(n335) );
  NANDN U710 ( .A(n606), .B(n607), .Z(n605) );
  NANDN U711 ( .A(n604), .B(n608), .Z(n607) );
  XOR U712 ( .A(n609), .B(n336), .Z(n334) );
  IV U713 ( .A(n332), .Z(n336) );
  XNOR U714 ( .A(n610), .B(n611), .Z(n332) );
  NAND U715 ( .A(n612), .B(n613), .Z(n611) );
  XOR U716 ( .A(n610), .B(n614), .Z(n612) );
  NOR U717 ( .A(n615), .B(n616), .Z(n609) );
  XNOR U718 ( .A(n373), .B(n346), .Z(n617) );
  XNOR U719 ( .A(n618), .B(n619), .Z(n346) );
  NANDN U720 ( .A(n620), .B(n621), .Z(n619) );
  XOR U721 ( .A(n618), .B(n622), .Z(n621) );
  XNOR U722 ( .A(n623), .B(n624), .Z(n354) );
  NANDN U723 ( .A(n625), .B(n626), .Z(n624) );
  NANDN U724 ( .A(n627), .B(n623), .Z(n626) );
  XNOR U725 ( .A(n628), .B(n351), .Z(n353) );
  XNOR U726 ( .A(n629), .B(n630), .Z(n351) );
  NAND U727 ( .A(n631), .B(n632), .Z(n630) );
  XNOR U728 ( .A(n629), .B(n633), .Z(n631) );
  NOR U729 ( .A(n634), .B(n635), .Z(n628) );
  XOR U730 ( .A(n360), .B(n363), .Z(n636) );
  XNOR U731 ( .A(n637), .B(n638), .Z(n363) );
  NANDN U732 ( .A(n639), .B(n640), .Z(n638) );
  XOR U733 ( .A(n637), .B(n641), .Z(n640) );
  XNOR U734 ( .A(n642), .B(n643), .Z(n360) );
  NANDN U735 ( .A(n644), .B(n645), .Z(n643) );
  NANDN U736 ( .A(n642), .B(n646), .Z(n645) );
  XOR U737 ( .A(n647), .B(n361), .Z(n359) );
  IV U738 ( .A(n357), .Z(n361) );
  XNOR U739 ( .A(n648), .B(n649), .Z(n357) );
  NAND U740 ( .A(n650), .B(n651), .Z(n649) );
  XOR U741 ( .A(n648), .B(n652), .Z(n650) );
  NOR U742 ( .A(n653), .B(n654), .Z(n647) );
  XNOR U743 ( .A(n390), .B(n370), .Z(n655) );
  XNOR U744 ( .A(n656), .B(n657), .Z(n370) );
  NANDN U745 ( .A(n658), .B(n659), .Z(n657) );
  XOR U746 ( .A(n656), .B(n660), .Z(n659) );
  XNOR U747 ( .A(n661), .B(n662), .Z(n378) );
  NANDN U748 ( .A(n663), .B(n664), .Z(n662) );
  NANDN U749 ( .A(n665), .B(n661), .Z(n664) );
  XNOR U750 ( .A(n666), .B(n375), .Z(n377) );
  XNOR U751 ( .A(n667), .B(n668), .Z(n375) );
  NAND U752 ( .A(n669), .B(n670), .Z(n668) );
  XNOR U753 ( .A(n667), .B(n671), .Z(n669) );
  NOR U754 ( .A(n672), .B(n673), .Z(n666) );
  XOR U755 ( .A(n384), .B(n387), .Z(n674) );
  XNOR U756 ( .A(n675), .B(n676), .Z(n387) );
  NANDN U757 ( .A(n677), .B(n678), .Z(n676) );
  XNOR U758 ( .A(n675), .B(n679), .Z(n678) );
  XNOR U759 ( .A(n680), .B(n681), .Z(n384) );
  NANDN U760 ( .A(n682), .B(n683), .Z(n681) );
  NANDN U761 ( .A(n680), .B(n684), .Z(n683) );
  XOR U762 ( .A(n685), .B(n385), .Z(n383) );
  IV U763 ( .A(n381), .Z(n385) );
  XNOR U764 ( .A(n686), .B(n687), .Z(n381) );
  NAND U765 ( .A(n688), .B(n689), .Z(n687) );
  XOR U766 ( .A(n686), .B(n690), .Z(n688) );
  NOR U767 ( .A(n691), .B(n692), .Z(n685) );
  XOR U768 ( .A(n693), .B(n694), .Z(n392) );
  NANDN U769 ( .A(n24), .B(n695), .Z(n694) );
  XNOR U770 ( .A(n693), .B(n25), .Z(n695) );
  XOR U771 ( .A(n403), .B(n404), .Z(n413) );
  XOR U772 ( .A(n398), .B(n396), .Z(n404) );
  AND U773 ( .A(n696), .B(n394), .Z(n396) );
  OR U774 ( .A(n697), .B(n698), .Z(n394) );
  OR U775 ( .A(n699), .B(n700), .Z(n696) );
  NOR U776 ( .A(n701), .B(n702), .Z(n398) );
  XOR U777 ( .A(n405), .B(n703), .Z(n403) );
  XOR U778 ( .A(n406), .B(n400), .Z(n703) );
  NOR U779 ( .A(n704), .B(n705), .Z(n400) );
  OR U780 ( .A(n706), .B(n707), .Z(n406) );
  AND U781 ( .A(n708), .B(n709), .Z(n405) );
  OR U782 ( .A(n710), .B(n711), .Z(n709) );
  OR U783 ( .A(n712), .B(n713), .Z(n708) );
  XNOR U784 ( .A(n423), .B(n714), .Z(n411) );
  XNOR U785 ( .A(n409), .B(n424), .Z(n714) );
  XOR U786 ( .A(n418), .B(n416), .Z(n424) );
  NOR U787 ( .A(n716), .B(n717), .Z(n414) );
  OR U788 ( .A(n718), .B(n719), .Z(n715) );
  OR U789 ( .A(n720), .B(n721), .Z(n418) );
  OR U790 ( .A(n722), .B(n723), .Z(n409) );
  XOR U791 ( .A(n425), .B(n724), .Z(n423) );
  XOR U792 ( .A(n426), .B(n420), .Z(n724) );
  NOR U793 ( .A(n725), .B(n726), .Z(n420) );
  OR U794 ( .A(n727), .B(n728), .Z(n426) );
  AND U795 ( .A(n729), .B(n730), .Z(n425) );
  OR U796 ( .A(n731), .B(n732), .Z(n730) );
  OR U797 ( .A(n733), .B(n734), .Z(n729) );
  XOR U798 ( .A(n428), .B(n451), .Z(n735) );
  XNOR U799 ( .A(n442), .B(n443), .Z(n451) );
  XOR U800 ( .A(n437), .B(n435), .Z(n443) );
  AND U801 ( .A(n736), .B(n433), .Z(n435) );
  OR U802 ( .A(n737), .B(n738), .Z(n433) );
  OR U803 ( .A(n739), .B(n740), .Z(n736) );
  NOR U804 ( .A(n741), .B(n742), .Z(n437) );
  XOR U805 ( .A(n444), .B(n743), .Z(n442) );
  XOR U806 ( .A(n445), .B(n439), .Z(n743) );
  NOR U807 ( .A(n744), .B(n745), .Z(n439) );
  OR U808 ( .A(n746), .B(n747), .Z(n445) );
  AND U809 ( .A(n748), .B(n749), .Z(n444) );
  OR U810 ( .A(n750), .B(n751), .Z(n749) );
  OR U811 ( .A(n752), .B(n753), .Z(n748) );
  OR U812 ( .A(n754), .B(n755), .Z(n428) );
  XNOR U813 ( .A(n461), .B(n756), .Z(n449) );
  XNOR U814 ( .A(n447), .B(n462), .Z(n756) );
  XOR U815 ( .A(n456), .B(n454), .Z(n462) );
  NOR U816 ( .A(n758), .B(n759), .Z(n452) );
  OR U817 ( .A(n760), .B(n761), .Z(n757) );
  OR U818 ( .A(n762), .B(n763), .Z(n456) );
  OR U819 ( .A(n764), .B(n765), .Z(n447) );
  XOR U820 ( .A(n463), .B(n766), .Z(n461) );
  XOR U821 ( .A(n464), .B(n458), .Z(n766) );
  NOR U822 ( .A(n767), .B(n768), .Z(n458) );
  OR U823 ( .A(n769), .B(n770), .Z(n464) );
  AND U824 ( .A(n771), .B(n772), .Z(n463) );
  OR U825 ( .A(n773), .B(n774), .Z(n772) );
  OR U826 ( .A(n775), .B(n776), .Z(n771) );
  XNOR U827 ( .A(n466), .B(n508), .Z(n777) );
  XOR U828 ( .A(n480), .B(n481), .Z(n489) );
  XOR U829 ( .A(n475), .B(n473), .Z(n481) );
  AND U830 ( .A(n778), .B(n471), .Z(n473) );
  OR U831 ( .A(n779), .B(n780), .Z(n471) );
  OR U832 ( .A(n781), .B(n782), .Z(n778) );
  NOR U833 ( .A(n783), .B(n784), .Z(n475) );
  XOR U834 ( .A(n482), .B(n785), .Z(n480) );
  XOR U835 ( .A(n483), .B(n477), .Z(n785) );
  NOR U836 ( .A(n786), .B(n787), .Z(n477) );
  OR U837 ( .A(n788), .B(n789), .Z(n483) );
  AND U838 ( .A(n790), .B(n791), .Z(n482) );
  OR U839 ( .A(n792), .B(n793), .Z(n791) );
  OR U840 ( .A(n794), .B(n795), .Z(n790) );
  XNOR U841 ( .A(n499), .B(n796), .Z(n487) );
  XNOR U842 ( .A(n485), .B(n500), .Z(n796) );
  XOR U843 ( .A(n494), .B(n492), .Z(n500) );
  NOR U844 ( .A(n798), .B(n799), .Z(n490) );
  OR U845 ( .A(n800), .B(n801), .Z(n797) );
  OR U846 ( .A(n802), .B(n803), .Z(n494) );
  OR U847 ( .A(n804), .B(n805), .Z(n485) );
  XOR U848 ( .A(n501), .B(n806), .Z(n499) );
  XOR U849 ( .A(n502), .B(n496), .Z(n806) );
  NOR U850 ( .A(n807), .B(n808), .Z(n496) );
  OR U851 ( .A(n809), .B(n810), .Z(n502) );
  AND U852 ( .A(n811), .B(n812), .Z(n501) );
  OR U853 ( .A(n813), .B(n814), .Z(n812) );
  OR U854 ( .A(n815), .B(n816), .Z(n811) );
  OR U855 ( .A(n817), .B(n818), .Z(n466) );
  XOR U856 ( .A(n504), .B(n527), .Z(n819) );
  XNOR U857 ( .A(n518), .B(n519), .Z(n527) );
  XOR U858 ( .A(n513), .B(n511), .Z(n519) );
  AND U859 ( .A(n820), .B(n509), .Z(n511) );
  OR U860 ( .A(n821), .B(n822), .Z(n509) );
  OR U861 ( .A(n823), .B(n824), .Z(n820) );
  NOR U862 ( .A(n825), .B(n826), .Z(n513) );
  XOR U863 ( .A(n520), .B(n827), .Z(n518) );
  XOR U864 ( .A(n521), .B(n515), .Z(n827) );
  NOR U865 ( .A(n828), .B(n829), .Z(n515) );
  OR U866 ( .A(n830), .B(n831), .Z(n521) );
  AND U867 ( .A(n832), .B(n833), .Z(n520) );
  OR U868 ( .A(n834), .B(n835), .Z(n833) );
  OR U869 ( .A(n836), .B(n837), .Z(n832) );
  OR U870 ( .A(n838), .B(n839), .Z(n504) );
  XNOR U871 ( .A(n537), .B(n840), .Z(n525) );
  XNOR U872 ( .A(n523), .B(n538), .Z(n840) );
  XOR U873 ( .A(n532), .B(n530), .Z(n538) );
  NOR U874 ( .A(n842), .B(n843), .Z(n528) );
  OR U875 ( .A(n844), .B(n845), .Z(n841) );
  OR U876 ( .A(n846), .B(n847), .Z(n532) );
  OR U877 ( .A(n848), .B(n849), .Z(n523) );
  XOR U878 ( .A(n539), .B(n850), .Z(n537) );
  XOR U879 ( .A(n540), .B(n534), .Z(n850) );
  NOR U880 ( .A(n851), .B(n852), .Z(n534) );
  OR U881 ( .A(n853), .B(n854), .Z(n540) );
  AND U882 ( .A(n855), .B(n856), .Z(n539) );
  OR U883 ( .A(n857), .B(n858), .Z(n856) );
  OR U884 ( .A(n859), .B(n860), .Z(n855) );
  XNOR U885 ( .A(n542), .B(n622), .Z(n861) );
  XOR U886 ( .A(n556), .B(n557), .Z(n565) );
  XOR U887 ( .A(n551), .B(n549), .Z(n557) );
  AND U888 ( .A(n862), .B(n547), .Z(n549) );
  OR U889 ( .A(n863), .B(n864), .Z(n547) );
  OR U890 ( .A(n865), .B(n866), .Z(n862) );
  NOR U891 ( .A(n867), .B(n868), .Z(n551) );
  XOR U892 ( .A(n558), .B(n869), .Z(n556) );
  XOR U893 ( .A(n559), .B(n553), .Z(n869) );
  NOR U894 ( .A(n870), .B(n871), .Z(n553) );
  OR U895 ( .A(n872), .B(n873), .Z(n559) );
  AND U896 ( .A(n874), .B(n875), .Z(n558) );
  OR U897 ( .A(n876), .B(n877), .Z(n875) );
  OR U898 ( .A(n878), .B(n879), .Z(n874) );
  XNOR U899 ( .A(n575), .B(n880), .Z(n563) );
  XNOR U900 ( .A(n561), .B(n576), .Z(n880) );
  XOR U901 ( .A(n570), .B(n568), .Z(n576) );
  NOR U902 ( .A(n882), .B(n883), .Z(n566) );
  OR U903 ( .A(n884), .B(n885), .Z(n881) );
  OR U904 ( .A(n886), .B(n887), .Z(n570) );
  OR U905 ( .A(n888), .B(n889), .Z(n561) );
  XOR U906 ( .A(n577), .B(n890), .Z(n575) );
  XOR U907 ( .A(n578), .B(n572), .Z(n890) );
  NOR U908 ( .A(n891), .B(n892), .Z(n572) );
  OR U909 ( .A(n893), .B(n894), .Z(n578) );
  AND U910 ( .A(n895), .B(n896), .Z(n577) );
  OR U911 ( .A(n897), .B(n898), .Z(n896) );
  OR U912 ( .A(n899), .B(n900), .Z(n895) );
  XOR U913 ( .A(n580), .B(n603), .Z(n901) );
  XNOR U914 ( .A(n594), .B(n595), .Z(n603) );
  XOR U915 ( .A(n589), .B(n587), .Z(n595) );
  AND U916 ( .A(n902), .B(n585), .Z(n587) );
  OR U917 ( .A(n903), .B(n904), .Z(n585) );
  OR U918 ( .A(n905), .B(n906), .Z(n902) );
  NOR U919 ( .A(n907), .B(n908), .Z(n589) );
  XOR U920 ( .A(n596), .B(n909), .Z(n594) );
  XOR U921 ( .A(n597), .B(n591), .Z(n909) );
  NOR U922 ( .A(n910), .B(n911), .Z(n591) );
  OR U923 ( .A(n912), .B(n913), .Z(n597) );
  AND U924 ( .A(n914), .B(n915), .Z(n596) );
  OR U925 ( .A(n916), .B(n917), .Z(n915) );
  OR U926 ( .A(n918), .B(n919), .Z(n914) );
  OR U927 ( .A(n920), .B(n921), .Z(n580) );
  XNOR U928 ( .A(n613), .B(n922), .Z(n601) );
  XNOR U929 ( .A(n599), .B(n614), .Z(n922) );
  XOR U930 ( .A(n608), .B(n606), .Z(n614) );
  NOR U931 ( .A(n924), .B(n925), .Z(n604) );
  OR U932 ( .A(n926), .B(n927), .Z(n923) );
  OR U933 ( .A(n928), .B(n929), .Z(n608) );
  OR U934 ( .A(n930), .B(n931), .Z(n599) );
  XOR U935 ( .A(n615), .B(n932), .Z(n613) );
  XOR U936 ( .A(n616), .B(n610), .Z(n932) );
  NOR U937 ( .A(n933), .B(n934), .Z(n610) );
  OR U938 ( .A(n935), .B(n936), .Z(n616) );
  AND U939 ( .A(n937), .B(n938), .Z(n615) );
  OR U940 ( .A(n939), .B(n940), .Z(n938) );
  OR U941 ( .A(n941), .B(n942), .Z(n937) );
  OR U942 ( .A(n943), .B(n944), .Z(n542) );
  XNOR U943 ( .A(n618), .B(n660), .Z(n945) );
  XOR U944 ( .A(n632), .B(n633), .Z(n641) );
  XOR U945 ( .A(n627), .B(n625), .Z(n633) );
  AND U946 ( .A(n946), .B(n623), .Z(n625) );
  OR U947 ( .A(n947), .B(n948), .Z(n623) );
  OR U948 ( .A(n949), .B(n950), .Z(n946) );
  NOR U949 ( .A(n951), .B(n952), .Z(n627) );
  XOR U950 ( .A(n634), .B(n953), .Z(n632) );
  XOR U951 ( .A(n635), .B(n629), .Z(n953) );
  NOR U952 ( .A(n954), .B(n955), .Z(n629) );
  OR U953 ( .A(n956), .B(n957), .Z(n635) );
  AND U954 ( .A(n958), .B(n959), .Z(n634) );
  OR U955 ( .A(n960), .B(n961), .Z(n959) );
  OR U956 ( .A(n962), .B(n963), .Z(n958) );
  XNOR U957 ( .A(n651), .B(n964), .Z(n639) );
  XNOR U958 ( .A(n637), .B(n652), .Z(n964) );
  XOR U959 ( .A(n646), .B(n644), .Z(n652) );
  NOR U960 ( .A(n966), .B(n967), .Z(n642) );
  OR U961 ( .A(n968), .B(n969), .Z(n965) );
  OR U962 ( .A(n970), .B(n971), .Z(n646) );
  OR U963 ( .A(n972), .B(n973), .Z(n637) );
  XOR U964 ( .A(n653), .B(n974), .Z(n651) );
  XOR U965 ( .A(n654), .B(n648), .Z(n974) );
  NOR U966 ( .A(n975), .B(n976), .Z(n648) );
  OR U967 ( .A(n977), .B(n978), .Z(n654) );
  AND U968 ( .A(n979), .B(n980), .Z(n653) );
  OR U969 ( .A(n981), .B(n982), .Z(n980) );
  OR U970 ( .A(n983), .B(n984), .Z(n979) );
  OR U971 ( .A(n985), .B(n986), .Z(n618) );
  XOR U972 ( .A(n656), .B(n679), .Z(n987) );
  XNOR U973 ( .A(n670), .B(n671), .Z(n679) );
  XOR U974 ( .A(n665), .B(n663), .Z(n671) );
  AND U975 ( .A(n988), .B(n661), .Z(n663) );
  OR U976 ( .A(n989), .B(n990), .Z(n661) );
  OR U977 ( .A(n991), .B(n992), .Z(n988) );
  NOR U978 ( .A(n993), .B(n994), .Z(n665) );
  XOR U979 ( .A(n672), .B(n995), .Z(n670) );
  XOR U980 ( .A(n673), .B(n667), .Z(n995) );
  NOR U981 ( .A(n996), .B(n997), .Z(n667) );
  OR U982 ( .A(n998), .B(n999), .Z(n673) );
  AND U983 ( .A(n1000), .B(n1001), .Z(n672) );
  OR U984 ( .A(n1002), .B(n1003), .Z(n1001) );
  OR U985 ( .A(n1004), .B(n1005), .Z(n1000) );
  OR U986 ( .A(n1006), .B(n1007), .Z(n656) );
  XNOR U987 ( .A(n689), .B(n1008), .Z(n677) );
  XNOR U988 ( .A(n675), .B(n690), .Z(n1008) );
  XOR U989 ( .A(n684), .B(n682), .Z(n690) );
  NOR U990 ( .A(n1010), .B(n1011), .Z(n680) );
  OR U991 ( .A(n1012), .B(n1013), .Z(n1009) );
  OR U992 ( .A(n1014), .B(n1015), .Z(n684) );
  OR U993 ( .A(n1016), .B(n1017), .Z(n675) );
  XOR U994 ( .A(n691), .B(n1018), .Z(n689) );
  XOR U995 ( .A(n692), .B(n686), .Z(n1018) );
  NOR U996 ( .A(n1019), .B(n1020), .Z(n686) );
  OR U997 ( .A(n1021), .B(n1022), .Z(n692) );
  AND U998 ( .A(n1023), .B(n1024), .Z(n691) );
  OR U999 ( .A(n1025), .B(n1026), .Z(n1024) );
  OR U1000 ( .A(n1027), .B(n1028), .Z(n1023) );
  XNOR U1001 ( .A(oglobal[1]), .B(n693), .Z(n24) );
  ANDN U1002 ( .B(oglobal[0]), .A(n1029), .Z(n693) );
  XNOR U1003 ( .A(oglobal[0]), .B(n1029), .Z(o[0]) );
  XNOR U1004 ( .A(n944), .B(n943), .Z(n1029) );
  XNOR U1005 ( .A(n818), .B(n817), .Z(n943) );
  XNOR U1006 ( .A(n755), .B(n754), .Z(n817) );
  XNOR U1007 ( .A(n723), .B(n722), .Z(n754) );
  XNOR U1008 ( .A(n697), .B(n698), .Z(n704) );
  XNOR U1009 ( .A(n701), .B(n702), .Z(n698) );
  XNOR U1010 ( .A(y[127]), .B(x[127]), .Z(n702) );
  XNOR U1011 ( .A(y[126]), .B(x[126]), .Z(n701) );
  XNOR U1012 ( .A(n699), .B(n700), .Z(n697) );
  XNOR U1013 ( .A(y[125]), .B(x[125]), .Z(n700) );
  XNOR U1014 ( .A(y[124]), .B(x[124]), .Z(n699) );
  XNOR U1015 ( .A(n712), .B(n713), .Z(n705) );
  XNOR U1016 ( .A(n707), .B(n706), .Z(n713) );
  XNOR U1017 ( .A(y[123]), .B(x[123]), .Z(n706) );
  XNOR U1018 ( .A(y[122]), .B(x[122]), .Z(n707) );
  XNOR U1019 ( .A(n710), .B(n711), .Z(n712) );
  XNOR U1020 ( .A(y[121]), .B(x[121]), .Z(n711) );
  XNOR U1021 ( .A(y[120]), .B(x[120]), .Z(n710) );
  XNOR U1022 ( .A(n716), .B(n717), .Z(n725) );
  XNOR U1023 ( .A(n720), .B(n721), .Z(n717) );
  XNOR U1024 ( .A(y[119]), .B(x[119]), .Z(n721) );
  XNOR U1025 ( .A(y[118]), .B(x[118]), .Z(n720) );
  XNOR U1026 ( .A(n718), .B(n719), .Z(n716) );
  XNOR U1027 ( .A(y[117]), .B(x[117]), .Z(n719) );
  XNOR U1028 ( .A(y[116]), .B(x[116]), .Z(n718) );
  XNOR U1029 ( .A(n733), .B(n734), .Z(n726) );
  XNOR U1030 ( .A(n728), .B(n727), .Z(n734) );
  XNOR U1031 ( .A(y[115]), .B(x[115]), .Z(n727) );
  XNOR U1032 ( .A(y[114]), .B(x[114]), .Z(n728) );
  XNOR U1033 ( .A(n731), .B(n732), .Z(n733) );
  XNOR U1034 ( .A(y[113]), .B(x[113]), .Z(n732) );
  XNOR U1035 ( .A(y[112]), .B(x[112]), .Z(n731) );
  XNOR U1036 ( .A(n765), .B(n764), .Z(n755) );
  XNOR U1037 ( .A(n737), .B(n738), .Z(n744) );
  XNOR U1038 ( .A(n741), .B(n742), .Z(n738) );
  XNOR U1039 ( .A(y[111]), .B(x[111]), .Z(n742) );
  XNOR U1040 ( .A(y[110]), .B(x[110]), .Z(n741) );
  XNOR U1041 ( .A(n739), .B(n740), .Z(n737) );
  XNOR U1042 ( .A(y[109]), .B(x[109]), .Z(n740) );
  XNOR U1043 ( .A(y[108]), .B(x[108]), .Z(n739) );
  XNOR U1044 ( .A(n752), .B(n753), .Z(n745) );
  XNOR U1045 ( .A(n747), .B(n746), .Z(n753) );
  XNOR U1046 ( .A(y[107]), .B(x[107]), .Z(n746) );
  XNOR U1047 ( .A(y[106]), .B(x[106]), .Z(n747) );
  XNOR U1048 ( .A(n750), .B(n751), .Z(n752) );
  XNOR U1049 ( .A(y[105]), .B(x[105]), .Z(n751) );
  XNOR U1050 ( .A(y[104]), .B(x[104]), .Z(n750) );
  XNOR U1051 ( .A(n758), .B(n759), .Z(n767) );
  XNOR U1052 ( .A(n762), .B(n763), .Z(n759) );
  XNOR U1053 ( .A(y[103]), .B(x[103]), .Z(n763) );
  XNOR U1054 ( .A(y[102]), .B(x[102]), .Z(n762) );
  XNOR U1055 ( .A(n760), .B(n761), .Z(n758) );
  XNOR U1056 ( .A(y[101]), .B(x[101]), .Z(n761) );
  XNOR U1057 ( .A(y[100]), .B(x[100]), .Z(n760) );
  XNOR U1058 ( .A(n775), .B(n776), .Z(n768) );
  XNOR U1059 ( .A(n770), .B(n769), .Z(n776) );
  XNOR U1060 ( .A(y[99]), .B(x[99]), .Z(n769) );
  XNOR U1061 ( .A(y[98]), .B(x[98]), .Z(n770) );
  XNOR U1062 ( .A(n773), .B(n774), .Z(n775) );
  XNOR U1063 ( .A(y[97]), .B(x[97]), .Z(n774) );
  XNOR U1064 ( .A(y[96]), .B(x[96]), .Z(n773) );
  XNOR U1065 ( .A(n839), .B(n838), .Z(n818) );
  XNOR U1066 ( .A(n805), .B(n804), .Z(n838) );
  XNOR U1067 ( .A(n779), .B(n780), .Z(n786) );
  XNOR U1068 ( .A(n783), .B(n784), .Z(n780) );
  XNOR U1069 ( .A(y[95]), .B(x[95]), .Z(n784) );
  XNOR U1070 ( .A(y[94]), .B(x[94]), .Z(n783) );
  XNOR U1071 ( .A(n781), .B(n782), .Z(n779) );
  XNOR U1072 ( .A(y[93]), .B(x[93]), .Z(n782) );
  XNOR U1073 ( .A(y[92]), .B(x[92]), .Z(n781) );
  XNOR U1074 ( .A(n794), .B(n795), .Z(n787) );
  XNOR U1075 ( .A(n789), .B(n788), .Z(n795) );
  XNOR U1076 ( .A(y[91]), .B(x[91]), .Z(n788) );
  XNOR U1077 ( .A(y[90]), .B(x[90]), .Z(n789) );
  XNOR U1078 ( .A(n792), .B(n793), .Z(n794) );
  XNOR U1079 ( .A(y[89]), .B(x[89]), .Z(n793) );
  XNOR U1080 ( .A(y[88]), .B(x[88]), .Z(n792) );
  XNOR U1081 ( .A(n798), .B(n799), .Z(n807) );
  XNOR U1082 ( .A(n802), .B(n803), .Z(n799) );
  XNOR U1083 ( .A(y[87]), .B(x[87]), .Z(n803) );
  XNOR U1084 ( .A(y[86]), .B(x[86]), .Z(n802) );
  XNOR U1085 ( .A(n800), .B(n801), .Z(n798) );
  XNOR U1086 ( .A(y[85]), .B(x[85]), .Z(n801) );
  XNOR U1087 ( .A(y[84]), .B(x[84]), .Z(n800) );
  XNOR U1088 ( .A(n815), .B(n816), .Z(n808) );
  XNOR U1089 ( .A(n810), .B(n809), .Z(n816) );
  XNOR U1090 ( .A(y[83]), .B(x[83]), .Z(n809) );
  XNOR U1091 ( .A(y[82]), .B(x[82]), .Z(n810) );
  XNOR U1092 ( .A(n813), .B(n814), .Z(n815) );
  XNOR U1093 ( .A(y[81]), .B(x[81]), .Z(n814) );
  XNOR U1094 ( .A(y[80]), .B(x[80]), .Z(n813) );
  XNOR U1095 ( .A(n849), .B(n848), .Z(n839) );
  XNOR U1096 ( .A(n821), .B(n822), .Z(n828) );
  XNOR U1097 ( .A(n825), .B(n826), .Z(n822) );
  XNOR U1098 ( .A(y[79]), .B(x[79]), .Z(n826) );
  XNOR U1099 ( .A(y[78]), .B(x[78]), .Z(n825) );
  XNOR U1100 ( .A(n823), .B(n824), .Z(n821) );
  XNOR U1101 ( .A(y[77]), .B(x[77]), .Z(n824) );
  XNOR U1102 ( .A(y[76]), .B(x[76]), .Z(n823) );
  XNOR U1103 ( .A(n836), .B(n837), .Z(n829) );
  XNOR U1104 ( .A(n831), .B(n830), .Z(n837) );
  XNOR U1105 ( .A(y[75]), .B(x[75]), .Z(n830) );
  XNOR U1106 ( .A(y[74]), .B(x[74]), .Z(n831) );
  XNOR U1107 ( .A(n834), .B(n835), .Z(n836) );
  XNOR U1108 ( .A(y[73]), .B(x[73]), .Z(n835) );
  XNOR U1109 ( .A(y[72]), .B(x[72]), .Z(n834) );
  XNOR U1110 ( .A(n842), .B(n843), .Z(n851) );
  XNOR U1111 ( .A(n846), .B(n847), .Z(n843) );
  XNOR U1112 ( .A(y[71]), .B(x[71]), .Z(n847) );
  XNOR U1113 ( .A(y[70]), .B(x[70]), .Z(n846) );
  XNOR U1114 ( .A(n844), .B(n845), .Z(n842) );
  XNOR U1115 ( .A(y[69]), .B(x[69]), .Z(n845) );
  XNOR U1116 ( .A(y[68]), .B(x[68]), .Z(n844) );
  XNOR U1117 ( .A(n859), .B(n860), .Z(n852) );
  XNOR U1118 ( .A(n854), .B(n853), .Z(n860) );
  XNOR U1119 ( .A(y[67]), .B(x[67]), .Z(n853) );
  XNOR U1120 ( .A(y[66]), .B(x[66]), .Z(n854) );
  XNOR U1121 ( .A(n857), .B(n858), .Z(n859) );
  XNOR U1122 ( .A(y[65]), .B(x[65]), .Z(n858) );
  XNOR U1123 ( .A(y[64]), .B(x[64]), .Z(n857) );
  XNOR U1124 ( .A(n986), .B(n985), .Z(n944) );
  XNOR U1125 ( .A(n921), .B(n920), .Z(n985) );
  XNOR U1126 ( .A(n889), .B(n888), .Z(n920) );
  XNOR U1127 ( .A(n863), .B(n864), .Z(n870) );
  XNOR U1128 ( .A(n867), .B(n868), .Z(n864) );
  XNOR U1129 ( .A(y[63]), .B(x[63]), .Z(n868) );
  XNOR U1130 ( .A(y[62]), .B(x[62]), .Z(n867) );
  XNOR U1131 ( .A(n865), .B(n866), .Z(n863) );
  XNOR U1132 ( .A(y[61]), .B(x[61]), .Z(n866) );
  XNOR U1133 ( .A(y[60]), .B(x[60]), .Z(n865) );
  XNOR U1134 ( .A(n878), .B(n879), .Z(n871) );
  XNOR U1135 ( .A(n873), .B(n872), .Z(n879) );
  XNOR U1136 ( .A(y[59]), .B(x[59]), .Z(n872) );
  XNOR U1137 ( .A(y[58]), .B(x[58]), .Z(n873) );
  XNOR U1138 ( .A(n876), .B(n877), .Z(n878) );
  XNOR U1139 ( .A(y[57]), .B(x[57]), .Z(n877) );
  XNOR U1140 ( .A(y[56]), .B(x[56]), .Z(n876) );
  XNOR U1141 ( .A(n882), .B(n883), .Z(n891) );
  XNOR U1142 ( .A(n886), .B(n887), .Z(n883) );
  XNOR U1143 ( .A(y[55]), .B(x[55]), .Z(n887) );
  XNOR U1144 ( .A(y[54]), .B(x[54]), .Z(n886) );
  XNOR U1145 ( .A(n884), .B(n885), .Z(n882) );
  XNOR U1146 ( .A(y[53]), .B(x[53]), .Z(n885) );
  XNOR U1147 ( .A(y[52]), .B(x[52]), .Z(n884) );
  XNOR U1148 ( .A(n899), .B(n900), .Z(n892) );
  XNOR U1149 ( .A(n894), .B(n893), .Z(n900) );
  XNOR U1150 ( .A(y[51]), .B(x[51]), .Z(n893) );
  XNOR U1151 ( .A(y[50]), .B(x[50]), .Z(n894) );
  XNOR U1152 ( .A(n897), .B(n898), .Z(n899) );
  XNOR U1153 ( .A(y[49]), .B(x[49]), .Z(n898) );
  XNOR U1154 ( .A(y[48]), .B(x[48]), .Z(n897) );
  XNOR U1155 ( .A(n931), .B(n930), .Z(n921) );
  XNOR U1156 ( .A(n903), .B(n904), .Z(n910) );
  XNOR U1157 ( .A(n907), .B(n908), .Z(n904) );
  XNOR U1158 ( .A(y[47]), .B(x[47]), .Z(n908) );
  XNOR U1159 ( .A(y[46]), .B(x[46]), .Z(n907) );
  XNOR U1160 ( .A(n905), .B(n906), .Z(n903) );
  XNOR U1161 ( .A(y[45]), .B(x[45]), .Z(n906) );
  XNOR U1162 ( .A(y[44]), .B(x[44]), .Z(n905) );
  XNOR U1163 ( .A(n918), .B(n919), .Z(n911) );
  XNOR U1164 ( .A(n913), .B(n912), .Z(n919) );
  XNOR U1165 ( .A(y[43]), .B(x[43]), .Z(n912) );
  XNOR U1166 ( .A(y[42]), .B(x[42]), .Z(n913) );
  XNOR U1167 ( .A(n916), .B(n917), .Z(n918) );
  XNOR U1168 ( .A(y[41]), .B(x[41]), .Z(n917) );
  XNOR U1169 ( .A(y[40]), .B(x[40]), .Z(n916) );
  XNOR U1170 ( .A(n924), .B(n925), .Z(n933) );
  XNOR U1171 ( .A(n928), .B(n929), .Z(n925) );
  XNOR U1172 ( .A(y[39]), .B(x[39]), .Z(n929) );
  XNOR U1173 ( .A(y[38]), .B(x[38]), .Z(n928) );
  XNOR U1174 ( .A(n926), .B(n927), .Z(n924) );
  XNOR U1175 ( .A(y[37]), .B(x[37]), .Z(n927) );
  XNOR U1176 ( .A(y[36]), .B(x[36]), .Z(n926) );
  XNOR U1177 ( .A(n941), .B(n942), .Z(n934) );
  XNOR U1178 ( .A(n936), .B(n935), .Z(n942) );
  XNOR U1179 ( .A(y[35]), .B(x[35]), .Z(n935) );
  XNOR U1180 ( .A(y[34]), .B(x[34]), .Z(n936) );
  XNOR U1181 ( .A(n939), .B(n940), .Z(n941) );
  XNOR U1182 ( .A(y[33]), .B(x[33]), .Z(n940) );
  XNOR U1183 ( .A(y[32]), .B(x[32]), .Z(n939) );
  XNOR U1184 ( .A(n1007), .B(n1006), .Z(n986) );
  XNOR U1185 ( .A(n973), .B(n972), .Z(n1006) );
  XNOR U1186 ( .A(n947), .B(n948), .Z(n954) );
  XNOR U1187 ( .A(n951), .B(n952), .Z(n948) );
  XNOR U1188 ( .A(y[31]), .B(x[31]), .Z(n952) );
  XNOR U1189 ( .A(y[30]), .B(x[30]), .Z(n951) );
  XNOR U1190 ( .A(n949), .B(n950), .Z(n947) );
  XNOR U1191 ( .A(y[29]), .B(x[29]), .Z(n950) );
  XNOR U1192 ( .A(y[28]), .B(x[28]), .Z(n949) );
  XNOR U1193 ( .A(n962), .B(n963), .Z(n955) );
  XNOR U1194 ( .A(n957), .B(n956), .Z(n963) );
  XNOR U1195 ( .A(y[27]), .B(x[27]), .Z(n956) );
  XNOR U1196 ( .A(y[26]), .B(x[26]), .Z(n957) );
  XNOR U1197 ( .A(n960), .B(n961), .Z(n962) );
  XNOR U1198 ( .A(y[25]), .B(x[25]), .Z(n961) );
  XNOR U1199 ( .A(y[24]), .B(x[24]), .Z(n960) );
  XNOR U1200 ( .A(n966), .B(n967), .Z(n975) );
  XNOR U1201 ( .A(n970), .B(n971), .Z(n967) );
  XNOR U1202 ( .A(y[23]), .B(x[23]), .Z(n971) );
  XNOR U1203 ( .A(y[22]), .B(x[22]), .Z(n970) );
  XNOR U1204 ( .A(n968), .B(n969), .Z(n966) );
  XNOR U1205 ( .A(y[21]), .B(x[21]), .Z(n969) );
  XNOR U1206 ( .A(y[20]), .B(x[20]), .Z(n968) );
  XNOR U1207 ( .A(n983), .B(n984), .Z(n976) );
  XNOR U1208 ( .A(n978), .B(n977), .Z(n984) );
  XNOR U1209 ( .A(y[19]), .B(x[19]), .Z(n977) );
  XNOR U1210 ( .A(y[18]), .B(x[18]), .Z(n978) );
  XNOR U1211 ( .A(n981), .B(n982), .Z(n983) );
  XNOR U1212 ( .A(y[17]), .B(x[17]), .Z(n982) );
  XNOR U1213 ( .A(y[16]), .B(x[16]), .Z(n981) );
  XNOR U1214 ( .A(n1017), .B(n1016), .Z(n1007) );
  XNOR U1215 ( .A(n989), .B(n990), .Z(n996) );
  XNOR U1216 ( .A(n993), .B(n994), .Z(n990) );
  XNOR U1217 ( .A(y[15]), .B(x[15]), .Z(n994) );
  XNOR U1218 ( .A(y[14]), .B(x[14]), .Z(n993) );
  XNOR U1219 ( .A(n991), .B(n992), .Z(n989) );
  XNOR U1220 ( .A(y[13]), .B(x[13]), .Z(n992) );
  XNOR U1221 ( .A(y[12]), .B(x[12]), .Z(n991) );
  XNOR U1222 ( .A(n1004), .B(n1005), .Z(n997) );
  XNOR U1223 ( .A(n999), .B(n998), .Z(n1005) );
  XNOR U1224 ( .A(y[11]), .B(x[11]), .Z(n998) );
  XNOR U1225 ( .A(y[10]), .B(x[10]), .Z(n999) );
  XNOR U1226 ( .A(n1002), .B(n1003), .Z(n1004) );
  XNOR U1227 ( .A(y[9]), .B(x[9]), .Z(n1003) );
  XNOR U1228 ( .A(y[8]), .B(x[8]), .Z(n1002) );
  XNOR U1229 ( .A(n1010), .B(n1011), .Z(n1019) );
  XNOR U1230 ( .A(n1014), .B(n1015), .Z(n1011) );
  XNOR U1231 ( .A(y[7]), .B(x[7]), .Z(n1015) );
  XNOR U1232 ( .A(y[6]), .B(x[6]), .Z(n1014) );
  XNOR U1233 ( .A(n1012), .B(n1013), .Z(n1010) );
  XNOR U1234 ( .A(y[5]), .B(x[5]), .Z(n1013) );
  XNOR U1235 ( .A(y[4]), .B(x[4]), .Z(n1012) );
  XNOR U1236 ( .A(n1027), .B(n1028), .Z(n1020) );
  XNOR U1237 ( .A(n1022), .B(n1021), .Z(n1028) );
  XNOR U1238 ( .A(y[3]), .B(x[3]), .Z(n1021) );
  XNOR U1239 ( .A(y[2]), .B(x[2]), .Z(n1022) );
  XNOR U1240 ( .A(n1025), .B(n1026), .Z(n1027) );
  XNOR U1241 ( .A(y[1]), .B(x[1]), .Z(n1026) );
  XNOR U1242 ( .A(y[0]), .B(x[0]), .Z(n1025) );
endmodule

