
module hamming_N1600_CC2 ( clk, rst, x, y, o );
  input [799:0] x;
  input [799:0] y;
  output [10:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801;
  wire   [10:0] oglobal;

  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  OR U803 ( .A(n2663), .B(n2664), .Z(n1) );
  OR U804 ( .A(n2661), .B(n2662), .Z(n2) );
  NAND U805 ( .A(n1), .B(n2), .Z(n2767) );
  OR U806 ( .A(n1900), .B(n1901), .Z(n3) );
  OR U807 ( .A(n1898), .B(n1899), .Z(n4) );
  NAND U808 ( .A(n3), .B(n4), .Z(n2888) );
  OR U809 ( .A(n1919), .B(n1920), .Z(n5) );
  OR U810 ( .A(n1917), .B(n1918), .Z(n6) );
  NAND U811 ( .A(n5), .B(n6), .Z(n2891) );
  OR U812 ( .A(n1122), .B(n1123), .Z(n7) );
  NANDN U813 ( .A(n1125), .B(n1124), .Z(n8) );
  NAND U814 ( .A(n7), .B(n8), .Z(n2827) );
  OR U815 ( .A(n2713), .B(n2714), .Z(n9) );
  NANDN U816 ( .A(n2716), .B(n2715), .Z(n10) );
  NAND U817 ( .A(n9), .B(n10), .Z(n3111) );
  OR U818 ( .A(n1880), .B(n1881), .Z(n11) );
  OR U819 ( .A(n1878), .B(n1879), .Z(n12) );
  NAND U820 ( .A(n11), .B(n12), .Z(n2987) );
  OR U821 ( .A(n1949), .B(n1950), .Z(n13) );
  OR U822 ( .A(n1947), .B(n1948), .Z(n14) );
  NAND U823 ( .A(n13), .B(n14), .Z(n2977) );
  OR U824 ( .A(n2259), .B(n2260), .Z(n15) );
  NANDN U825 ( .A(n2262), .B(n2261), .Z(n16) );
  AND U826 ( .A(n15), .B(n16), .Z(n2964) );
  OR U827 ( .A(n1931), .B(n1932), .Z(n17) );
  NANDN U828 ( .A(n1934), .B(n1933), .Z(n18) );
  NAND U829 ( .A(n17), .B(n18), .Z(n2916) );
  OR U830 ( .A(n1386), .B(n1387), .Z(n19) );
  NANDN U831 ( .A(n1389), .B(n1388), .Z(n20) );
  NAND U832 ( .A(n19), .B(n20), .Z(n2869) );
  OR U833 ( .A(n2463), .B(n2464), .Z(n21) );
  OR U834 ( .A(n2461), .B(n2462), .Z(n22) );
  NAND U835 ( .A(n21), .B(n22), .Z(n2851) );
  OR U836 ( .A(n2617), .B(n2618), .Z(n23) );
  NANDN U837 ( .A(n2620), .B(n2619), .Z(n24) );
  NAND U838 ( .A(n23), .B(n24), .Z(n2941) );
  OR U839 ( .A(n2013), .B(n2014), .Z(n25) );
  OR U840 ( .A(n2011), .B(n2012), .Z(n26) );
  AND U841 ( .A(n25), .B(n26), .Z(n3592) );
  OR U842 ( .A(n1852), .B(n1853), .Z(n27) );
  OR U843 ( .A(n1850), .B(n1851), .Z(n28) );
  NAND U844 ( .A(n27), .B(n28), .Z(n2927) );
  OR U845 ( .A(n2147), .B(n2148), .Z(n29) );
  OR U846 ( .A(n2145), .B(n2146), .Z(n30) );
  NAND U847 ( .A(n29), .B(n30), .Z(n3653) );
  OR U848 ( .A(n2919), .B(n2920), .Z(n31) );
  NANDN U849 ( .A(n2922), .B(n2921), .Z(n32) );
  NAND U850 ( .A(n31), .B(n32), .Z(n3952) );
  OR U851 ( .A(n3015), .B(n3016), .Z(n33) );
  OR U852 ( .A(n3013), .B(n3014), .Z(n34) );
  NAND U853 ( .A(n33), .B(n34), .Z(n4003) );
  NANDN U854 ( .A(n3006), .B(n3005), .Z(n35) );
  NANDN U855 ( .A(n3007), .B(n3008), .Z(n36) );
  AND U856 ( .A(n35), .B(n36), .Z(n4241) );
  OR U857 ( .A(n4069), .B(n4070), .Z(n37) );
  OR U858 ( .A(n4067), .B(n4068), .Z(n38) );
  NAND U859 ( .A(n37), .B(n38), .Z(n4427) );
  OR U860 ( .A(n4034), .B(n4035), .Z(n39) );
  NANDN U861 ( .A(n4033), .B(n4032), .Z(n40) );
  AND U862 ( .A(n39), .B(n40), .Z(n4526) );
  NANDN U863 ( .A(n3958), .B(n3957), .Z(n41) );
  NANDN U864 ( .A(n3955), .B(n3956), .Z(n42) );
  NAND U865 ( .A(n41), .B(n42), .Z(n4314) );
  NANDN U866 ( .A(n4029), .B(n4028), .Z(n43) );
  NANDN U867 ( .A(n4030), .B(n4031), .Z(n44) );
  AND U868 ( .A(n43), .B(n44), .Z(n4445) );
  OR U869 ( .A(n4335), .B(n4336), .Z(n45) );
  NANDN U870 ( .A(n4337), .B(n4338), .Z(n46) );
  NAND U871 ( .A(n45), .B(n46), .Z(n4623) );
  OR U872 ( .A(n4508), .B(n4509), .Z(n47) );
  OR U873 ( .A(n4506), .B(n4507), .Z(n48) );
  AND U874 ( .A(n47), .B(n48), .Z(n4613) );
  OR U875 ( .A(n4541), .B(n4542), .Z(n49) );
  NANDN U876 ( .A(n4544), .B(n4543), .Z(n50) );
  AND U877 ( .A(n49), .B(n50), .Z(n4641) );
  OR U878 ( .A(n4719), .B(n4720), .Z(n51) );
  NANDN U879 ( .A(n4722), .B(n4721), .Z(n52) );
  NAND U880 ( .A(n51), .B(n52), .Z(n4750) );
  OR U881 ( .A(n1244), .B(n1245), .Z(n53) );
  NANDN U882 ( .A(n1247), .B(n1246), .Z(n54) );
  NAND U883 ( .A(n53), .B(n54), .Z(n3622) );
  OR U884 ( .A(n2659), .B(n2660), .Z(n55) );
  OR U885 ( .A(n2657), .B(n2658), .Z(n56) );
  NAND U886 ( .A(n55), .B(n56), .Z(n2768) );
  OR U887 ( .A(n823), .B(n824), .Z(n57) );
  NANDN U888 ( .A(n826), .B(n825), .Z(n58) );
  NAND U889 ( .A(n57), .B(n58), .Z(n2761) );
  OR U890 ( .A(n1140), .B(n1141), .Z(n59) );
  NANDN U891 ( .A(n1143), .B(n1142), .Z(n60) );
  NAND U892 ( .A(n59), .B(n60), .Z(n2895) );
  OR U893 ( .A(n1915), .B(n1916), .Z(n61) );
  OR U894 ( .A(n1913), .B(n1914), .Z(n62) );
  NAND U895 ( .A(n61), .B(n62), .Z(n2892) );
  OR U896 ( .A(n1126), .B(n1127), .Z(n63) );
  NANDN U897 ( .A(n1129), .B(n1128), .Z(n64) );
  NAND U898 ( .A(n63), .B(n64), .Z(n2829) );
  OR U899 ( .A(n1520), .B(n1521), .Z(n65) );
  NANDN U900 ( .A(n1523), .B(n1522), .Z(n66) );
  NAND U901 ( .A(n65), .B(n66), .Z(n2839) );
  OR U902 ( .A(n1170), .B(n1171), .Z(n67) );
  OR U903 ( .A(n1168), .B(n1169), .Z(n68) );
  NAND U904 ( .A(n67), .B(n68), .Z(n3106) );
  OR U905 ( .A(n1888), .B(n1889), .Z(n69) );
  OR U906 ( .A(n1886), .B(n1887), .Z(n70) );
  NAND U907 ( .A(n69), .B(n70), .Z(n2992) );
  OR U908 ( .A(n1876), .B(n1877), .Z(n71) );
  OR U909 ( .A(n1874), .B(n1875), .Z(n72) );
  NAND U910 ( .A(n71), .B(n72), .Z(n2988) );
  OR U911 ( .A(n799), .B(n800), .Z(n73) );
  NANDN U912 ( .A(n802), .B(n801), .Z(n74) );
  NAND U913 ( .A(n73), .B(n74), .Z(n2981) );
  OR U914 ( .A(n1945), .B(n1946), .Z(n75) );
  OR U915 ( .A(n1943), .B(n1944), .Z(n76) );
  NAND U916 ( .A(n75), .B(n76), .Z(n2978) );
  OR U917 ( .A(n1872), .B(n1873), .Z(n77) );
  OR U918 ( .A(n1870), .B(n1871), .Z(n78) );
  NAND U919 ( .A(n77), .B(n78), .Z(n2976) );
  OR U920 ( .A(n2001), .B(n2002), .Z(n79) );
  OR U921 ( .A(n1999), .B(n2000), .Z(n80) );
  NAND U922 ( .A(n79), .B(n80), .Z(n2815) );
  OR U923 ( .A(n1576), .B(n1577), .Z(n81) );
  NANDN U924 ( .A(n1579), .B(n1578), .Z(n82) );
  NAND U925 ( .A(n81), .B(n82), .Z(n2755) );
  OR U926 ( .A(n1438), .B(n1439), .Z(n83) );
  NANDN U927 ( .A(n1441), .B(n1440), .Z(n84) );
  NAND U928 ( .A(n83), .B(n84), .Z(n2953) );
  OR U929 ( .A(n2023), .B(n2024), .Z(n85) );
  NANDN U930 ( .A(n2026), .B(n2025), .Z(n86) );
  AND U931 ( .A(n85), .B(n86), .Z(n3371) );
  OR U932 ( .A(n2071), .B(n2072), .Z(n87) );
  OR U933 ( .A(n2069), .B(n2070), .Z(n88) );
  NAND U934 ( .A(n87), .B(n88), .Z(n3127) );
  OR U935 ( .A(n2671), .B(n2672), .Z(n89) );
  OR U936 ( .A(n2669), .B(n2670), .Z(n90) );
  NAND U937 ( .A(n89), .B(n90), .Z(n2912) );
  OR U938 ( .A(n1546), .B(n1547), .Z(n91) );
  NANDN U939 ( .A(n1549), .B(n1548), .Z(n92) );
  NAND U940 ( .A(n91), .B(n92), .Z(n2881) );
  OR U941 ( .A(n1382), .B(n1383), .Z(n93) );
  NANDN U942 ( .A(n1385), .B(n1384), .Z(n94) );
  NAND U943 ( .A(n93), .B(n94), .Z(n2870) );
  OR U944 ( .A(n1418), .B(n1419), .Z(n95) );
  NANDN U945 ( .A(n1421), .B(n1420), .Z(n96) );
  NAND U946 ( .A(n95), .B(n96), .Z(n3347) );
  OR U947 ( .A(n2039), .B(n2040), .Z(n97) );
  NANDN U948 ( .A(n2042), .B(n2041), .Z(n98) );
  AND U949 ( .A(n97), .B(n98), .Z(n3354) );
  OR U950 ( .A(n2055), .B(n2056), .Z(n99) );
  OR U951 ( .A(n2053), .B(n2054), .Z(n100) );
  NAND U952 ( .A(n99), .B(n100), .Z(n3045) );
  OR U953 ( .A(n1296), .B(n1297), .Z(n101) );
  OR U954 ( .A(n1294), .B(n1295), .Z(n102) );
  NAND U955 ( .A(n101), .B(n102), .Z(n2950) );
  OR U956 ( .A(n2613), .B(n2614), .Z(n103) );
  NANDN U957 ( .A(n2616), .B(n2615), .Z(n104) );
  NAND U958 ( .A(n103), .B(n104), .Z(n2942) );
  OR U959 ( .A(n2009), .B(n2010), .Z(n105) );
  OR U960 ( .A(n2007), .B(n2008), .Z(n106) );
  NAND U961 ( .A(n105), .B(n106), .Z(n3593) );
  OR U962 ( .A(n1848), .B(n1849), .Z(n107) );
  OR U963 ( .A(n1846), .B(n1847), .Z(n108) );
  NAND U964 ( .A(n107), .B(n108), .Z(n2928) );
  OR U965 ( .A(n1961), .B(n1962), .Z(n109) );
  OR U966 ( .A(n1959), .B(n1960), .Z(n110) );
  NAND U967 ( .A(n109), .B(n110), .Z(n2923) );
  OR U968 ( .A(n1969), .B(n1970), .Z(n111) );
  OR U969 ( .A(n1967), .B(n1968), .Z(n112) );
  NAND U970 ( .A(n111), .B(n112), .Z(n2920) );
  OR U971 ( .A(n1498), .B(n1499), .Z(n113) );
  NAND U972 ( .A(n1501), .B(n1500), .Z(n114) );
  NAND U973 ( .A(n113), .B(n114), .Z(n3499) );
  OR U974 ( .A(n2887), .B(n2888), .Z(n115) );
  NAND U975 ( .A(n2889), .B(n2890), .Z(n116) );
  AND U976 ( .A(n115), .B(n116), .Z(n4233) );
  OR U977 ( .A(n3111), .B(n3110), .Z(n117) );
  NANDN U978 ( .A(n3112), .B(n3113), .Z(n118) );
  AND U979 ( .A(n117), .B(n118), .Z(n4224) );
  OR U980 ( .A(n2963), .B(n2964), .Z(n119) );
  NANDN U981 ( .A(n2965), .B(n2966), .Z(n120) );
  NAND U982 ( .A(n119), .B(n120), .Z(n4179) );
  OR U983 ( .A(n2916), .B(n2915), .Z(n121) );
  NANDN U984 ( .A(n2917), .B(n2918), .Z(n122) );
  AND U985 ( .A(n121), .B(n122), .Z(n3951) );
  OR U986 ( .A(n3052), .B(n3053), .Z(n123) );
  NANDN U987 ( .A(n3055), .B(n3054), .Z(n124) );
  NAND U988 ( .A(n123), .B(n124), .Z(n4152) );
  OR U989 ( .A(n3011), .B(n3012), .Z(n125) );
  OR U990 ( .A(n3009), .B(n3010), .Z(n126) );
  NAND U991 ( .A(n125), .B(n126), .Z(n4005) );
  OR U992 ( .A(n3185), .B(n3186), .Z(n127) );
  NAND U993 ( .A(n3187), .B(n3188), .Z(n128) );
  AND U994 ( .A(n127), .B(n128), .Z(n4272) );
  OR U995 ( .A(n4281), .B(n4282), .Z(n129) );
  NAND U996 ( .A(n4284), .B(n4283), .Z(n130) );
  NAND U997 ( .A(n129), .B(n130), .Z(n4439) );
  OR U998 ( .A(n4083), .B(n4084), .Z(n131) );
  NANDN U999 ( .A(n4086), .B(n4085), .Z(n132) );
  AND U1000 ( .A(n131), .B(n132), .Z(n4432) );
  NANDN U1001 ( .A(n4151), .B(n4150), .Z(n133) );
  NANDN U1002 ( .A(n4148), .B(n4149), .Z(n134) );
  NAND U1003 ( .A(n133), .B(n134), .Z(n4331) );
  OR U1004 ( .A(n3935), .B(n3936), .Z(n135) );
  OR U1005 ( .A(n3933), .B(n3934), .Z(n136) );
  NAND U1006 ( .A(n135), .B(n136), .Z(n4534) );
  NANDN U1007 ( .A(n3199), .B(n3200), .Z(n137) );
  NANDN U1008 ( .A(n3202), .B(n3201), .Z(n138) );
  AND U1009 ( .A(n137), .B(n138), .Z(n4135) );
  OR U1010 ( .A(n4073), .B(n4074), .Z(n139) );
  OR U1011 ( .A(n4071), .B(n4072), .Z(n140) );
  NAND U1012 ( .A(n139), .B(n140), .Z(n4428) );
  OR U1013 ( .A(n4525), .B(n4526), .Z(n141) );
  OR U1014 ( .A(n4523), .B(n4524), .Z(n142) );
  AND U1015 ( .A(n141), .B(n142), .Z(n4638) );
  OR U1016 ( .A(n4343), .B(n4344), .Z(n143) );
  NANDN U1017 ( .A(n4345), .B(n4346), .Z(n144) );
  NAND U1018 ( .A(n143), .B(n144), .Z(n4618) );
  NANDN U1019 ( .A(n4502), .B(n4503), .Z(n145) );
  NANDN U1020 ( .A(n4504), .B(n4505), .Z(n146) );
  NAND U1021 ( .A(n145), .B(n146), .Z(n4615) );
  OR U1022 ( .A(n4539), .B(n4540), .Z(n147) );
  OR U1023 ( .A(n4537), .B(n4538), .Z(n148) );
  AND U1024 ( .A(n147), .B(n148), .Z(n4640) );
  OR U1025 ( .A(n4099), .B(n4100), .Z(n149) );
  NAND U1026 ( .A(n4102), .B(n4101), .Z(n150) );
  NAND U1027 ( .A(n149), .B(n150), .Z(n4386) );
  NANDN U1028 ( .A(n4119), .B(n4120), .Z(n151) );
  NANDN U1029 ( .A(n4121), .B(n4122), .Z(n152) );
  NAND U1030 ( .A(n151), .B(n152), .Z(n4477) );
  OR U1031 ( .A(n4627), .B(n4628), .Z(n153) );
  NAND U1032 ( .A(n4630), .B(n4629), .Z(n154) );
  NAND U1033 ( .A(n153), .B(n154), .Z(n4702) );
  OR U1034 ( .A(n4692), .B(n4693), .Z(n155) );
  NANDN U1035 ( .A(n4694), .B(n4695), .Z(n156) );
  AND U1036 ( .A(n155), .B(n156), .Z(n4769) );
  XNOR U1037 ( .A(n4454), .B(n4455), .Z(n4457) );
  OR U1038 ( .A(n4305), .B(n4306), .Z(n157) );
  NANDN U1039 ( .A(n4308), .B(n4307), .Z(n158) );
  AND U1040 ( .A(n157), .B(n158), .Z(n4675) );
  XOR U1041 ( .A(n4740), .B(n4741), .Z(n4743) );
  OR U1042 ( .A(n1240), .B(n1241), .Z(n159) );
  NANDN U1043 ( .A(n1243), .B(n1242), .Z(n160) );
  NAND U1044 ( .A(n159), .B(n160), .Z(n3623) );
  OR U1045 ( .A(n901), .B(n902), .Z(n161) );
  NANDN U1046 ( .A(n904), .B(n903), .Z(n162) );
  NAND U1047 ( .A(n161), .B(n162), .Z(n2772) );
  OR U1048 ( .A(n2667), .B(n2668), .Z(n163) );
  OR U1049 ( .A(n2665), .B(n2666), .Z(n164) );
  NAND U1050 ( .A(n163), .B(n164), .Z(n2770) );
  OR U1051 ( .A(n819), .B(n820), .Z(n165) );
  NANDN U1052 ( .A(n822), .B(n821), .Z(n166) );
  NAND U1053 ( .A(n165), .B(n166), .Z(n2762) );
  OR U1054 ( .A(n1516), .B(n1517), .Z(n167) );
  NANDN U1055 ( .A(n1519), .B(n1518), .Z(n168) );
  NAND U1056 ( .A(n167), .B(n168), .Z(n2840) );
  OR U1057 ( .A(n2721), .B(n2722), .Z(n169) );
  NANDN U1058 ( .A(n2724), .B(n2723), .Z(n170) );
  NAND U1059 ( .A(n169), .B(n170), .Z(n3112) );
  OR U1060 ( .A(n1892), .B(n1893), .Z(n171) );
  OR U1061 ( .A(n1890), .B(n1891), .Z(n172) );
  NAND U1062 ( .A(n171), .B(n172), .Z(n2991) );
  OR U1063 ( .A(n1884), .B(n1885), .Z(n173) );
  OR U1064 ( .A(n1882), .B(n1883), .Z(n174) );
  NAND U1065 ( .A(n173), .B(n174), .Z(n2990) );
  OR U1066 ( .A(n1997), .B(n1998), .Z(n175) );
  OR U1067 ( .A(n1995), .B(n1996), .Z(n176) );
  NAND U1068 ( .A(n175), .B(n176), .Z(n2816) );
  OR U1069 ( .A(n953), .B(n954), .Z(n177) );
  NANDN U1070 ( .A(n956), .B(n955), .Z(n178) );
  NAND U1071 ( .A(n177), .B(n178), .Z(n2810) );
  OR U1072 ( .A(n941), .B(n942), .Z(n179) );
  OR U1073 ( .A(n939), .B(n940), .Z(n180) );
  NAND U1074 ( .A(n179), .B(n180), .Z(n2805) );
  OR U1075 ( .A(n1564), .B(n1565), .Z(n181) );
  NANDN U1076 ( .A(n1567), .B(n1566), .Z(n182) );
  NAND U1077 ( .A(n181), .B(n182), .Z(n3580) );
  OR U1078 ( .A(n2249), .B(n2250), .Z(n183) );
  NANDN U1079 ( .A(n2252), .B(n2251), .Z(n184) );
  AND U1080 ( .A(n183), .B(n184), .Z(n2965) );
  OR U1081 ( .A(n1021), .B(n1022), .Z(n185) );
  OR U1082 ( .A(n1019), .B(n1020), .Z(n186) );
  NAND U1083 ( .A(n185), .B(n186), .Z(n2959) );
  OR U1084 ( .A(n2019), .B(n2020), .Z(n187) );
  NANDN U1085 ( .A(n2022), .B(n2021), .Z(n188) );
  NAND U1086 ( .A(n187), .B(n188), .Z(n3372) );
  OR U1087 ( .A(n1374), .B(n1375), .Z(n189) );
  NANDN U1088 ( .A(n1377), .B(n1376), .Z(n190) );
  NAND U1089 ( .A(n189), .B(n190), .Z(n3365) );
  OR U1090 ( .A(n2095), .B(n2096), .Z(n191) );
  NANDN U1091 ( .A(n2098), .B(n2097), .Z(n192) );
  AND U1092 ( .A(n191), .B(n192), .Z(n3359) );
  OR U1093 ( .A(n2075), .B(n2076), .Z(n193) );
  OR U1094 ( .A(n2073), .B(n2074), .Z(n194) );
  NAND U1095 ( .A(n193), .B(n194), .Z(n3126) );
  OR U1096 ( .A(n1390), .B(n1391), .Z(n195) );
  NANDN U1097 ( .A(n1393), .B(n1392), .Z(n196) );
  NAND U1098 ( .A(n195), .B(n196), .Z(n2871) );
  OR U1099 ( .A(n1608), .B(n1609), .Z(n197) );
  NANDN U1100 ( .A(n1611), .B(n1610), .Z(n198) );
  NAND U1101 ( .A(n197), .B(n198), .Z(n3562) );
  OR U1102 ( .A(n1594), .B(n1595), .Z(n199) );
  NANDN U1103 ( .A(n1597), .B(n1596), .Z(n200) );
  NAND U1104 ( .A(n199), .B(n200), .Z(n3558) );
  OR U1105 ( .A(n1358), .B(n1359), .Z(n201) );
  NANDN U1106 ( .A(n1361), .B(n1360), .Z(n202) );
  NAND U1107 ( .A(n201), .B(n202), .Z(n2864) );
  OR U1108 ( .A(n2459), .B(n2460), .Z(n203) );
  OR U1109 ( .A(n2457), .B(n2458), .Z(n204) );
  NAND U1110 ( .A(n203), .B(n204), .Z(n2852) );
  OR U1111 ( .A(n2057), .B(n2058), .Z(n205) );
  NANDN U1112 ( .A(n2060), .B(n2059), .Z(n206) );
  NAND U1113 ( .A(n205), .B(n206), .Z(n3044) );
  OR U1114 ( .A(n1088), .B(n1089), .Z(n207) );
  NANDN U1115 ( .A(n1091), .B(n1090), .Z(n208) );
  NAND U1116 ( .A(n207), .B(n208), .Z(n3068) );
  OR U1117 ( .A(n2621), .B(n2622), .Z(n209) );
  NANDN U1118 ( .A(n2624), .B(n2623), .Z(n210) );
  NAND U1119 ( .A(n209), .B(n210), .Z(n2943) );
  OR U1120 ( .A(n721), .B(n722), .Z(n211) );
  NANDN U1121 ( .A(n724), .B(n723), .Z(n212) );
  NAND U1122 ( .A(n211), .B(n212), .Z(n3605) );
  OR U1123 ( .A(n2693), .B(n2694), .Z(n213) );
  OR U1124 ( .A(n2691), .B(n2692), .Z(n214) );
  AND U1125 ( .A(n213), .B(n214), .Z(n3598) );
  OR U1126 ( .A(n2017), .B(n2018), .Z(n215) );
  OR U1127 ( .A(n2015), .B(n2016), .Z(n216) );
  NAND U1128 ( .A(n215), .B(n216), .Z(n3595) );
  OR U1129 ( .A(n1957), .B(n1958), .Z(n217) );
  OR U1130 ( .A(n1955), .B(n1956), .Z(n218) );
  NAND U1131 ( .A(n217), .B(n218), .Z(n2924) );
  OR U1132 ( .A(n1506), .B(n1507), .Z(n219) );
  NANDN U1133 ( .A(n1509), .B(n1508), .Z(n220) );
  NAND U1134 ( .A(n219), .B(n220), .Z(n3539) );
  OR U1135 ( .A(n2117), .B(n2118), .Z(n221) );
  NANDN U1136 ( .A(n2119), .B(n2120), .Z(n222) );
  NAND U1137 ( .A(n221), .B(n222), .Z(n2904) );
  NANDN U1138 ( .A(n1715), .B(n1714), .Z(n223) );
  NANDN U1139 ( .A(n1716), .B(n1717), .Z(n224) );
  NAND U1140 ( .A(n223), .B(n224), .Z(n3411) );
  OR U1141 ( .A(n1158), .B(n1159), .Z(n225) );
  OR U1142 ( .A(n1156), .B(n1157), .Z(n226) );
  AND U1143 ( .A(n225), .B(n226), .Z(n3658) );
  XNOR U1144 ( .A(n3652), .B(n3653), .Z(n3654) );
  OR U1145 ( .A(n969), .B(n970), .Z(n227) );
  NANDN U1146 ( .A(n972), .B(n971), .Z(n228) );
  AND U1147 ( .A(n227), .B(n228), .Z(n3460) );
  OR U1148 ( .A(n713), .B(n714), .Z(n229) );
  NANDN U1149 ( .A(n716), .B(n715), .Z(n230) );
  NAND U1150 ( .A(n229), .B(n230), .Z(n3486) );
  NANDN U1151 ( .A(n762), .B(n761), .Z(n231) );
  NANDN U1152 ( .A(n763), .B(n764), .Z(n232) );
  AND U1153 ( .A(n231), .B(n232), .Z(n3695) );
  OR U1154 ( .A(n3732), .B(n3733), .Z(n233) );
  NAND U1155 ( .A(n3734), .B(n3735), .Z(n234) );
  AND U1156 ( .A(n233), .B(n234), .Z(n4067) );
  OR U1157 ( .A(n2779), .B(n2780), .Z(n235) );
  OR U1158 ( .A(n2777), .B(n2778), .Z(n236) );
  NAND U1159 ( .A(n235), .B(n236), .Z(n4037) );
  OR U1160 ( .A(n3626), .B(n3627), .Z(n237) );
  NANDN U1161 ( .A(n3629), .B(n3628), .Z(n238) );
  NAND U1162 ( .A(n237), .B(n238), .Z(n4213) );
  OR U1163 ( .A(n3106), .B(n3107), .Z(n239) );
  NANDN U1164 ( .A(n3109), .B(n3108), .Z(n240) );
  AND U1165 ( .A(n239), .B(n240), .Z(n4223) );
  OR U1166 ( .A(n2995), .B(n2996), .Z(n241) );
  NANDN U1167 ( .A(n2998), .B(n2997), .Z(n242) );
  AND U1168 ( .A(n241), .B(n242), .Z(n3928) );
  OR U1169 ( .A(n2954), .B(n2953), .Z(n243) );
  NANDN U1170 ( .A(n2955), .B(n2956), .Z(n244) );
  AND U1171 ( .A(n243), .B(n244), .Z(n4181) );
  OR U1172 ( .A(n3048), .B(n3049), .Z(n245) );
  NANDN U1173 ( .A(n3051), .B(n3050), .Z(n246) );
  AND U1174 ( .A(n245), .B(n246), .Z(n4153) );
  OR U1175 ( .A(n2949), .B(n2950), .Z(n247) );
  NANDN U1176 ( .A(n2952), .B(n2951), .Z(n248) );
  AND U1177 ( .A(n247), .B(n248), .Z(n3908) );
  OR U1178 ( .A(n2927), .B(n2928), .Z(n249) );
  NANDN U1179 ( .A(n2930), .B(n2929), .Z(n250) );
  AND U1180 ( .A(n249), .B(n250), .Z(n3913) );
  NANDN U1181 ( .A(n3286), .B(n3285), .Z(n251) );
  NANDN U1182 ( .A(n3287), .B(n3288), .Z(n252) );
  AND U1183 ( .A(n251), .B(n252), .Z(n3986) );
  OR U1184 ( .A(n3098), .B(n3099), .Z(n253) );
  NANDN U1185 ( .A(n3101), .B(n3100), .Z(n254) );
  NAND U1186 ( .A(n253), .B(n254), .Z(n3943) );
  OR U1187 ( .A(n3181), .B(n3182), .Z(n255) );
  NANDN U1188 ( .A(n3183), .B(n3184), .Z(n256) );
  AND U1189 ( .A(n255), .B(n256), .Z(n4271) );
  OR U1190 ( .A(n4279), .B(n4280), .Z(n257) );
  OR U1191 ( .A(n4277), .B(n4278), .Z(n258) );
  AND U1192 ( .A(n257), .B(n258), .Z(n4438) );
  OR U1193 ( .A(n3939), .B(n3940), .Z(n259) );
  NANDN U1194 ( .A(n3938), .B(n3937), .Z(n260) );
  NAND U1195 ( .A(n259), .B(n260), .Z(n4419) );
  OR U1196 ( .A(n4231), .B(n4232), .Z(n261) );
  NANDN U1197 ( .A(n4233), .B(n4234), .Z(n262) );
  NAND U1198 ( .A(n261), .B(n262), .Z(n4401) );
  OR U1199 ( .A(n3925), .B(n3926), .Z(n263) );
  OR U1200 ( .A(n3923), .B(n3924), .Z(n264) );
  AND U1201 ( .A(n263), .B(n264), .Z(n4326) );
  NANDN U1202 ( .A(n4191), .B(n4190), .Z(n265) );
  NANDN U1203 ( .A(n4188), .B(n4189), .Z(n266) );
  NAND U1204 ( .A(n265), .B(n266), .Z(n4319) );
  NANDN U1205 ( .A(n3954), .B(n3953), .Z(n267) );
  NANDN U1206 ( .A(n3951), .B(n3952), .Z(n268) );
  NAND U1207 ( .A(n267), .B(n268), .Z(n4316) );
  OR U1208 ( .A(n4144), .B(n4145), .Z(n269) );
  NAND U1209 ( .A(n4147), .B(n4146), .Z(n270) );
  NAND U1210 ( .A(n269), .B(n270), .Z(n4332) );
  NANDN U1211 ( .A(n4195), .B(n4194), .Z(n271) );
  NANDN U1212 ( .A(n4192), .B(n4193), .Z(n272) );
  NAND U1213 ( .A(n271), .B(n272), .Z(n4342) );
  OR U1214 ( .A(n4004), .B(n4005), .Z(n273) );
  OR U1215 ( .A(n4002), .B(n4003), .Z(n274) );
  AND U1216 ( .A(n273), .B(n274), .Z(n4311) );
  OR U1217 ( .A(n3947), .B(n3948), .Z(n275) );
  NANDN U1218 ( .A(n3950), .B(n3949), .Z(n276) );
  NAND U1219 ( .A(n275), .B(n276), .Z(n4365) );
  NANDN U1220 ( .A(n3966), .B(n3967), .Z(n277) );
  NANDN U1221 ( .A(n3969), .B(n3968), .Z(n278) );
  AND U1222 ( .A(n277), .B(n278), .Z(n4361) );
  OR U1223 ( .A(n3984), .B(n3985), .Z(n279) );
  OR U1224 ( .A(n3982), .B(n3983), .Z(n280) );
  AND U1225 ( .A(n279), .B(n280), .Z(n4498) );
  OR U1226 ( .A(n4024), .B(n4025), .Z(n281) );
  NANDN U1227 ( .A(n4026), .B(n4027), .Z(n282) );
  AND U1228 ( .A(n281), .B(n282), .Z(n4444) );
  OR U1229 ( .A(n4136), .B(n4137), .Z(n283) );
  OR U1230 ( .A(n4134), .B(n4135), .Z(n284) );
  AND U1231 ( .A(n283), .B(n284), .Z(n4494) );
  OR U1232 ( .A(n3171), .B(n3172), .Z(n285) );
  NAND U1233 ( .A(n3174), .B(n3173), .Z(n286) );
  NAND U1234 ( .A(n285), .B(n286), .Z(n4076) );
  NANDN U1235 ( .A(n4115), .B(n4116), .Z(n287) );
  NANDN U1236 ( .A(n4117), .B(n4118), .Z(n288) );
  AND U1237 ( .A(n287), .B(n288), .Z(n4476) );
  OR U1238 ( .A(n4422), .B(n4423), .Z(n289) );
  NANDN U1239 ( .A(n4425), .B(n4424), .Z(n290) );
  AND U1240 ( .A(n289), .B(n290), .Z(n4566) );
  OR U1241 ( .A(n4638), .B(n4639), .Z(n291) );
  NANDN U1242 ( .A(n4637), .B(n4636), .Z(n292) );
  AND U1243 ( .A(n291), .B(n292), .Z(n4710) );
  OR U1244 ( .A(n4613), .B(n4614), .Z(n293) );
  NAND U1245 ( .A(n4616), .B(n4615), .Z(n294) );
  NAND U1246 ( .A(n293), .B(n294), .Z(n4708) );
  OR U1247 ( .A(n4385), .B(n4386), .Z(n295) );
  NANDN U1248 ( .A(n4388), .B(n4387), .Z(n296) );
  AND U1249 ( .A(n295), .B(n296), .Z(n4588) );
  OR U1250 ( .A(n4703), .B(n4704), .Z(n297) );
  OR U1251 ( .A(n4701), .B(n4702), .Z(n298) );
  NAND U1252 ( .A(n297), .B(n298), .Z(n4761) );
  OR U1253 ( .A(n4697), .B(n4696), .Z(n299) );
  NANDN U1254 ( .A(n4698), .B(n4699), .Z(n300) );
  AND U1255 ( .A(n299), .B(n300), .Z(n4766) );
  XOR U1256 ( .A(n4457), .B(n4456), .Z(n4304) );
  XOR U1257 ( .A(n4674), .B(n4675), .Z(n4677) );
  OR U1258 ( .A(n4729), .B(n4730), .Z(n301) );
  NANDN U1259 ( .A(n4732), .B(n4731), .Z(n302) );
  AND U1260 ( .A(n301), .B(n302), .Z(n4742) );
  OR U1261 ( .A(n4751), .B(n4752), .Z(n303) );
  OR U1262 ( .A(n4749), .B(n4750), .Z(n304) );
  NAND U1263 ( .A(n303), .B(n304), .Z(n4777) );
  OR U1264 ( .A(n1250), .B(n1251), .Z(n305) );
  OR U1265 ( .A(n1248), .B(n1249), .Z(n306) );
  NAND U1266 ( .A(n305), .B(n306), .Z(n3625) );
  OR U1267 ( .A(n911), .B(n912), .Z(n307) );
  NANDN U1268 ( .A(n914), .B(n913), .Z(n308) );
  NAND U1269 ( .A(n307), .B(n308), .Z(n2773) );
  OR U1270 ( .A(n827), .B(n828), .Z(n309) );
  NANDN U1271 ( .A(n830), .B(n829), .Z(n310) );
  NAND U1272 ( .A(n309), .B(n310), .Z(n2763) );
  OR U1273 ( .A(n1144), .B(n1145), .Z(n311) );
  NANDN U1274 ( .A(n1147), .B(n1146), .Z(n312) );
  NAND U1275 ( .A(n311), .B(n312), .Z(n2897) );
  OR U1276 ( .A(n1923), .B(n1924), .Z(n313) );
  OR U1277 ( .A(n1921), .B(n1922), .Z(n314) );
  NAND U1278 ( .A(n313), .B(n314), .Z(n2893) );
  OR U1279 ( .A(n2717), .B(n2718), .Z(n315) );
  NANDN U1280 ( .A(n2720), .B(n2719), .Z(n316) );
  NAND U1281 ( .A(n315), .B(n316), .Z(n3110) );
  OR U1282 ( .A(n1166), .B(n1167), .Z(n317) );
  OR U1283 ( .A(n1164), .B(n1165), .Z(n318) );
  NAND U1284 ( .A(n317), .B(n318), .Z(n3107) );
  OR U1285 ( .A(n795), .B(n796), .Z(n319) );
  NANDN U1286 ( .A(n798), .B(n797), .Z(n320) );
  NAND U1287 ( .A(n319), .B(n320), .Z(n2982) );
  OR U1288 ( .A(n1953), .B(n1954), .Z(n321) );
  OR U1289 ( .A(n1951), .B(n1952), .Z(n322) );
  AND U1290 ( .A(n321), .B(n322), .Z(n2979) );
  OR U1291 ( .A(n1580), .B(n1581), .Z(n323) );
  NANDN U1292 ( .A(n1583), .B(n1582), .Z(n324) );
  NAND U1293 ( .A(n323), .B(n324), .Z(n2757) );
  OR U1294 ( .A(n1664), .B(n1665), .Z(n325) );
  NANDN U1295 ( .A(n1667), .B(n1666), .Z(n326) );
  NAND U1296 ( .A(n325), .B(n326), .Z(n2750) );
  OR U1297 ( .A(n1568), .B(n1569), .Z(n327) );
  NANDN U1298 ( .A(n1571), .B(n1570), .Z(n328) );
  NAND U1299 ( .A(n327), .B(n328), .Z(n3582) );
  OR U1300 ( .A(n1378), .B(n1379), .Z(n329) );
  NANDN U1301 ( .A(n1381), .B(n1380), .Z(n330) );
  NAND U1302 ( .A(n329), .B(n330), .Z(n3367) );
  OR U1303 ( .A(n2079), .B(n2080), .Z(n331) );
  OR U1304 ( .A(n2077), .B(n2078), .Z(n332) );
  NAND U1305 ( .A(n331), .B(n332), .Z(n3129) );
  OR U1306 ( .A(n1941), .B(n1942), .Z(n333) );
  OR U1307 ( .A(n1939), .B(n1940), .Z(n334) );
  NAND U1308 ( .A(n333), .B(n334), .Z(n2917) );
  OR U1309 ( .A(n1338), .B(n1339), .Z(n335) );
  OR U1310 ( .A(n1336), .B(n1337), .Z(n336) );
  NAND U1311 ( .A(n335), .B(n336), .Z(n3038) );
  OR U1312 ( .A(n1826), .B(n1827), .Z(n337) );
  NANDN U1313 ( .A(n1829), .B(n1828), .Z(n338) );
  NAND U1314 ( .A(n337), .B(n338), .Z(n3029) );
  OR U1315 ( .A(n1550), .B(n1551), .Z(n339) );
  NANDN U1316 ( .A(n1553), .B(n1552), .Z(n340) );
  NAND U1317 ( .A(n339), .B(n340), .Z(n2883) );
  OR U1318 ( .A(n1604), .B(n1605), .Z(n341) );
  NANDN U1319 ( .A(n1607), .B(n1606), .Z(n342) );
  NAND U1320 ( .A(n341), .B(n342), .Z(n3563) );
  OR U1321 ( .A(n1590), .B(n1591), .Z(n343) );
  NANDN U1322 ( .A(n1593), .B(n1592), .Z(n344) );
  NAND U1323 ( .A(n343), .B(n344), .Z(n3559) );
  OR U1324 ( .A(n1362), .B(n1363), .Z(n345) );
  NANDN U1325 ( .A(n1365), .B(n1364), .Z(n346) );
  NAND U1326 ( .A(n345), .B(n346), .Z(n2863) );
  OR U1327 ( .A(n1400), .B(n1401), .Z(n347) );
  NANDN U1328 ( .A(n1403), .B(n1402), .Z(n348) );
  NAND U1329 ( .A(n347), .B(n348), .Z(n2857) );
  OR U1330 ( .A(n2465), .B(n2466), .Z(n349) );
  NANDN U1331 ( .A(n2468), .B(n2467), .Z(n350) );
  NAND U1332 ( .A(n349), .B(n350), .Z(n2853) );
  OR U1333 ( .A(n1422), .B(n1423), .Z(n351) );
  NANDN U1334 ( .A(n1425), .B(n1424), .Z(n352) );
  NAND U1335 ( .A(n351), .B(n352), .Z(n3349) );
  OR U1336 ( .A(n1232), .B(n1233), .Z(n353) );
  NANDN U1337 ( .A(n1235), .B(n1234), .Z(n354) );
  NAND U1338 ( .A(n353), .B(n354), .Z(n3341) );
  OR U1339 ( .A(n2035), .B(n2036), .Z(n355) );
  NANDN U1340 ( .A(n2038), .B(n2037), .Z(n356) );
  NAND U1341 ( .A(n355), .B(n356), .Z(n3353) );
  OR U1342 ( .A(n1322), .B(n1323), .Z(n357) );
  OR U1343 ( .A(n1320), .B(n1321), .Z(n358) );
  NAND U1344 ( .A(n357), .B(n358), .Z(n3048) );
  OR U1345 ( .A(n1636), .B(n1637), .Z(n359) );
  NANDN U1346 ( .A(n1639), .B(n1638), .Z(n360) );
  NAND U1347 ( .A(n359), .B(n360), .Z(n3086) );
  OR U1348 ( .A(n1084), .B(n1085), .Z(n361) );
  NANDN U1349 ( .A(n1087), .B(n1086), .Z(n362) );
  NAND U1350 ( .A(n361), .B(n362), .Z(n3066) );
  OR U1351 ( .A(n1692), .B(n1693), .Z(n363) );
  NANDN U1352 ( .A(n1695), .B(n1694), .Z(n364) );
  NAND U1353 ( .A(n363), .B(n364), .Z(n3062) );
  OR U1354 ( .A(n1300), .B(n1301), .Z(n365) );
  OR U1355 ( .A(n1298), .B(n1299), .Z(n366) );
  NAND U1356 ( .A(n365), .B(n366), .Z(n2949) );
  OR U1357 ( .A(n733), .B(n734), .Z(n367) );
  OR U1358 ( .A(n731), .B(n732), .Z(n368) );
  NAND U1359 ( .A(n367), .B(n368), .Z(n3606) );
  OR U1360 ( .A(n2697), .B(n2698), .Z(n369) );
  OR U1361 ( .A(n2695), .B(n2696), .Z(n370) );
  NAND U1362 ( .A(n369), .B(n370), .Z(n3600) );
  OR U1363 ( .A(n1963), .B(n1964), .Z(n371) );
  NANDN U1364 ( .A(n1966), .B(n1965), .Z(n372) );
  NAND U1365 ( .A(n371), .B(n372), .Z(n2925) );
  OR U1366 ( .A(n1620), .B(n1621), .Z(n373) );
  NANDN U1367 ( .A(n1623), .B(n1622), .Z(n374) );
  AND U1368 ( .A(n373), .B(n374), .Z(n3543) );
  OR U1369 ( .A(n1502), .B(n1503), .Z(n375) );
  NANDN U1370 ( .A(n1505), .B(n1504), .Z(n376) );
  NAND U1371 ( .A(n375), .B(n376), .Z(n3540) );
  OR U1372 ( .A(n881), .B(n882), .Z(n377) );
  NANDN U1373 ( .A(n884), .B(n883), .Z(n378) );
  AND U1374 ( .A(n377), .B(n378), .Z(n2799) );
  OR U1375 ( .A(n1047), .B(n1048), .Z(n379) );
  NANDN U1376 ( .A(n1050), .B(n1049), .Z(n380) );
  AND U1377 ( .A(n379), .B(n380), .Z(n3437) );
  NANDN U1378 ( .A(n2088), .B(n2087), .Z(n381) );
  NANDN U1379 ( .A(n2089), .B(n2090), .Z(n382) );
  NAND U1380 ( .A(n381), .B(n382), .Z(n3262) );
  OR U1381 ( .A(n1152), .B(n1153), .Z(n383) );
  NANDN U1382 ( .A(n1155), .B(n1154), .Z(n384) );
  NAND U1383 ( .A(n383), .B(n384), .Z(n3659) );
  OR U1384 ( .A(n2155), .B(n2156), .Z(n385) );
  NANDN U1385 ( .A(n2158), .B(n2157), .Z(n386) );
  NAND U1386 ( .A(n385), .B(n386), .Z(n3655) );
  OR U1387 ( .A(n838), .B(n837), .Z(n387) );
  NANDN U1388 ( .A(n839), .B(n840), .Z(n388) );
  AND U1389 ( .A(n387), .B(n388), .Z(n3468) );
  OR U1390 ( .A(n949), .B(n950), .Z(n389) );
  NANDN U1391 ( .A(n952), .B(n951), .Z(n390) );
  NAND U1392 ( .A(n389), .B(n390), .Z(n3462) );
  OR U1393 ( .A(n2709), .B(n2710), .Z(n391) );
  NANDN U1394 ( .A(n2712), .B(n2711), .Z(n392) );
  NAND U1395 ( .A(n391), .B(n392), .Z(n3393) );
  OR U1396 ( .A(n2487), .B(n2488), .Z(n393) );
  NANDN U1397 ( .A(n2490), .B(n2489), .Z(n394) );
  NAND U1398 ( .A(n393), .B(n394), .Z(n3072) );
  NANDN U1399 ( .A(n2066), .B(n2065), .Z(n395) );
  NANDN U1400 ( .A(n2067), .B(n2068), .Z(n396) );
  NAND U1401 ( .A(n395), .B(n396), .Z(n3250) );
  OR U1402 ( .A(n2005), .B(n2006), .Z(n397) );
  OR U1403 ( .A(n2003), .B(n2004), .Z(n398) );
  NAND U1404 ( .A(n397), .B(n398), .Z(n2817) );
  OR U1405 ( .A(n1973), .B(n1974), .Z(n399) );
  OR U1406 ( .A(n1971), .B(n1972), .Z(n400) );
  NAND U1407 ( .A(n399), .B(n400), .Z(n2919) );
  OR U1408 ( .A(n1896), .B(n1897), .Z(n401) );
  OR U1409 ( .A(n1894), .B(n1895), .Z(n402) );
  NAND U1410 ( .A(n401), .B(n402), .Z(n2993) );
  OR U1411 ( .A(n1856), .B(n1857), .Z(n403) );
  OR U1412 ( .A(n1854), .B(n1855), .Z(n404) );
  NAND U1413 ( .A(n403), .B(n404), .Z(n2930) );
  NANDN U1414 ( .A(n794), .B(n793), .Z(n405) );
  NANDN U1415 ( .A(n791), .B(n792), .Z(n406) );
  NAND U1416 ( .A(n405), .B(n406), .Z(n3717) );
  OR U1417 ( .A(n1496), .B(n1497), .Z(n407) );
  NANDN U1418 ( .A(n1495), .B(n1494), .Z(n408) );
  NAND U1419 ( .A(n407), .B(n408), .Z(n3502) );
  NANDN U1420 ( .A(n3695), .B(n3694), .Z(n409) );
  NANDN U1421 ( .A(n3696), .B(n3697), .Z(n410) );
  AND U1422 ( .A(n409), .B(n410), .Z(n4287) );
  OR U1423 ( .A(n3548), .B(n3549), .Z(n411) );
  NANDN U1424 ( .A(n3551), .B(n3550), .Z(n412) );
  AND U1425 ( .A(n411), .B(n412), .Z(n4084) );
  OR U1426 ( .A(n2767), .B(n2768), .Z(n413) );
  NANDN U1427 ( .A(n2770), .B(n2769), .Z(n414) );
  AND U1428 ( .A(n413), .B(n414), .Z(n4219) );
  OR U1429 ( .A(n3102), .B(n3103), .Z(n415) );
  NANDN U1430 ( .A(n3105), .B(n3104), .Z(n416) );
  AND U1431 ( .A(n415), .B(n416), .Z(n4225) );
  OR U1432 ( .A(n2987), .B(n2988), .Z(n417) );
  NANDN U1433 ( .A(n2990), .B(n2989), .Z(n418) );
  AND U1434 ( .A(n417), .B(n418), .Z(n3930) );
  OR U1435 ( .A(n2973), .B(n2974), .Z(n419) );
  NANDN U1436 ( .A(n2976), .B(n2975), .Z(n420) );
  AND U1437 ( .A(n419), .B(n420), .Z(n3926) );
  OR U1438 ( .A(n2911), .B(n2912), .Z(n421) );
  NANDN U1439 ( .A(n2914), .B(n2913), .Z(n422) );
  NAND U1440 ( .A(n421), .B(n422), .Z(n3953) );
  OR U1441 ( .A(n3044), .B(n3045), .Z(n423) );
  NANDN U1442 ( .A(n3047), .B(n3046), .Z(n424) );
  NAND U1443 ( .A(n423), .B(n424), .Z(n4154) );
  OR U1444 ( .A(n2942), .B(n2941), .Z(n425) );
  NANDN U1445 ( .A(n2943), .B(n2944), .Z(n426) );
  AND U1446 ( .A(n425), .B(n426), .Z(n3910) );
  NANDN U1447 ( .A(n3444), .B(n3443), .Z(n427) );
  NANDN U1448 ( .A(n3445), .B(n3446), .Z(n428) );
  AND U1449 ( .A(n427), .B(n428), .Z(n3897) );
  OR U1450 ( .A(n3154), .B(n3155), .Z(n429) );
  OR U1451 ( .A(n3152), .B(n3153), .Z(n430) );
  AND U1452 ( .A(n429), .B(n430), .Z(n3849) );
  NANDN U1453 ( .A(n3411), .B(n3412), .Z(n431) );
  NANDN U1454 ( .A(n3414), .B(n3413), .Z(n432) );
  AND U1455 ( .A(n431), .B(n432), .Z(n3882) );
  NANDN U1456 ( .A(n3518), .B(n3517), .Z(n433) );
  NANDN U1457 ( .A(n3519), .B(n3520), .Z(n434) );
  AND U1458 ( .A(n433), .B(n434), .Z(n3947) );
  NANDN U1459 ( .A(n3390), .B(n3389), .Z(n435) );
  NANDN U1460 ( .A(n3391), .B(n3392), .Z(n436) );
  AND U1461 ( .A(n435), .B(n436), .Z(n3996) );
  OR U1462 ( .A(n3415), .B(n3416), .Z(n437) );
  NAND U1463 ( .A(n3417), .B(n3418), .Z(n438) );
  AND U1464 ( .A(n437), .B(n438), .Z(n3877) );
  OR U1465 ( .A(n1781), .B(n1780), .Z(n439) );
  NANDN U1466 ( .A(n1782), .B(n1783), .Z(n440) );
  AND U1467 ( .A(n439), .B(n440), .Z(n2732) );
  NANDN U1468 ( .A(n3858), .B(n3857), .Z(n441) );
  NANDN U1469 ( .A(n3855), .B(n3856), .Z(n442) );
  NAND U1470 ( .A(n441), .B(n442), .Z(n4528) );
  OR U1471 ( .A(n4036), .B(n4037), .Z(n443) );
  NANDN U1472 ( .A(n4039), .B(n4038), .Z(n444) );
  AND U1473 ( .A(n443), .B(n444), .Z(n4523) );
  OR U1474 ( .A(n4227), .B(n4228), .Z(n445) );
  NANDN U1475 ( .A(n4229), .B(n4230), .Z(n446) );
  NAND U1476 ( .A(n445), .B(n446), .Z(n4402) );
  OR U1477 ( .A(n4178), .B(n4179), .Z(n447) );
  NANDN U1478 ( .A(n4181), .B(n4180), .Z(n448) );
  NAND U1479 ( .A(n447), .B(n448), .Z(n4322) );
  OR U1480 ( .A(n4249), .B(n4250), .Z(n449) );
  NANDN U1481 ( .A(n4251), .B(n4252), .Z(n450) );
  NAND U1482 ( .A(n449), .B(n450), .Z(n4512) );
  OR U1483 ( .A(n3817), .B(n3818), .Z(n451) );
  NANDN U1484 ( .A(n3819), .B(n3820), .Z(n452) );
  NAND U1485 ( .A(n451), .B(n452), .Z(n4542) );
  OR U1486 ( .A(n4158), .B(n4159), .Z(n453) );
  NAND U1487 ( .A(n4161), .B(n4160), .Z(n454) );
  NAND U1488 ( .A(n453), .B(n454), .Z(n4354) );
  OR U1489 ( .A(n3865), .B(n3866), .Z(n455) );
  NANDN U1490 ( .A(n3868), .B(n3867), .Z(n456) );
  NAND U1491 ( .A(n455), .B(n456), .Z(n4412) );
  OR U1492 ( .A(n1148), .B(n1149), .Z(n457) );
  NANDN U1493 ( .A(n1151), .B(n1150), .Z(n458) );
  NAND U1494 ( .A(n457), .B(n458), .Z(n3001) );
  NANDN U1495 ( .A(n4241), .B(n4242), .Z(n459) );
  NANDN U1496 ( .A(n4243), .B(n4244), .Z(n460) );
  NAND U1497 ( .A(n459), .B(n460), .Z(n4390) );
  OR U1498 ( .A(n4053), .B(n4054), .Z(n461) );
  NANDN U1499 ( .A(n4056), .B(n4055), .Z(n462) );
  AND U1500 ( .A(n461), .B(n462), .Z(n4545) );
  NANDN U1501 ( .A(n4419), .B(n4418), .Z(n463) );
  NANDN U1502 ( .A(n4420), .B(n4421), .Z(n464) );
  NAND U1503 ( .A(n463), .B(n464), .Z(n4594) );
  OR U1504 ( .A(n4339), .B(n4340), .Z(n465) );
  NANDN U1505 ( .A(n4342), .B(n4341), .Z(n466) );
  NAND U1506 ( .A(n465), .B(n466), .Z(n4620) );
  OR U1507 ( .A(n4533), .B(n4534), .Z(n467) );
  NANDN U1508 ( .A(n4535), .B(n4536), .Z(n468) );
  NAND U1509 ( .A(n467), .B(n468), .Z(n4643) );
  OR U1510 ( .A(n4081), .B(n4082), .Z(n469) );
  OR U1511 ( .A(n4079), .B(n4080), .Z(n470) );
  NAND U1512 ( .A(n469), .B(n470), .Z(n4388) );
  OR U1513 ( .A(n4075), .B(n4076), .Z(n471) );
  NAND U1514 ( .A(n4077), .B(n4078), .Z(n472) );
  AND U1515 ( .A(n471), .B(n472), .Z(n4467) );
  OR U1516 ( .A(n4500), .B(n4501), .Z(n473) );
  OR U1517 ( .A(n4498), .B(n4499), .Z(n474) );
  NAND U1518 ( .A(n473), .B(n474), .Z(n4610) );
  OR U1519 ( .A(n4603), .B(n4604), .Z(n475) );
  NANDN U1520 ( .A(n4606), .B(n4605), .Z(n476) );
  AND U1521 ( .A(n475), .B(n476), .Z(n4714) );
  OR U1522 ( .A(n4623), .B(n4624), .Z(n477) );
  NANDN U1523 ( .A(n4626), .B(n4625), .Z(n478) );
  AND U1524 ( .A(n477), .B(n478), .Z(n4701) );
  OR U1525 ( .A(n4125), .B(n4126), .Z(n479) );
  OR U1526 ( .A(n4123), .B(n4124), .Z(n480) );
  NAND U1527 ( .A(n479), .B(n480), .Z(n4478) );
  OR U1528 ( .A(n4709), .B(n4710), .Z(n481) );
  NANDN U1529 ( .A(n4712), .B(n4711), .Z(n482) );
  NAND U1530 ( .A(n481), .B(n482), .Z(n4753) );
  OR U1531 ( .A(n4130), .B(n4131), .Z(n483) );
  NANDN U1532 ( .A(n4132), .B(n4133), .Z(n484) );
  NAND U1533 ( .A(n483), .B(n484), .Z(n4308) );
  OR U1534 ( .A(n4557), .B(n4558), .Z(n485) );
  OR U1535 ( .A(n4555), .B(n4556), .Z(n486) );
  AND U1536 ( .A(n485), .B(n486), .Z(n4732) );
  OR U1537 ( .A(n4766), .B(n4767), .Z(n487) );
  NANDN U1538 ( .A(n4769), .B(n4768), .Z(n488) );
  NAND U1539 ( .A(n487), .B(n488), .Z(n4780) );
  OR U1540 ( .A(n1812), .B(n1813), .Z(n489) );
  NAND U1541 ( .A(n1814), .B(n1815), .Z(n490) );
  AND U1542 ( .A(n489), .B(n490), .Z(n3222) );
  XOR U1543 ( .A(n4554), .B(n4553), .Z(n491) );
  NANDN U1544 ( .A(n4552), .B(n491), .Z(n492) );
  NAND U1545 ( .A(n4554), .B(n4553), .Z(n493) );
  AND U1546 ( .A(n492), .B(n493), .Z(n4681) );
  NAND U1547 ( .A(n4773), .B(n4771), .Z(n494) );
  XOR U1548 ( .A(n4771), .B(n4773), .Z(n495) );
  NANDN U1549 ( .A(n4772), .B(n495), .Z(n496) );
  NAND U1550 ( .A(n494), .B(n496), .Z(n4786) );
  OR U1551 ( .A(n1981), .B(n1982), .Z(n497) );
  OR U1552 ( .A(n1979), .B(n1980), .Z(n498) );
  NAND U1553 ( .A(n497), .B(n498), .Z(n3627) );
  OR U1554 ( .A(n2447), .B(n2448), .Z(n499) );
  NANDN U1555 ( .A(n2450), .B(n2449), .Z(n500) );
  AND U1556 ( .A(n499), .B(n500), .Z(n3616) );
  OR U1557 ( .A(n1911), .B(n1912), .Z(n501) );
  OR U1558 ( .A(n1909), .B(n1910), .Z(n502) );
  AND U1559 ( .A(n501), .B(n502), .Z(n2889) );
  OR U1560 ( .A(n1136), .B(n1137), .Z(n503) );
  NANDN U1561 ( .A(n1139), .B(n1138), .Z(n504) );
  NAND U1562 ( .A(n503), .B(n504), .Z(n2896) );
  OR U1563 ( .A(n1524), .B(n1525), .Z(n505) );
  NANDN U1564 ( .A(n1527), .B(n1526), .Z(n506) );
  NAND U1565 ( .A(n505), .B(n506), .Z(n2841) );
  OR U1566 ( .A(n767), .B(n768), .Z(n507) );
  OR U1567 ( .A(n765), .B(n766), .Z(n508) );
  NAND U1568 ( .A(n507), .B(n508), .Z(n2996) );
  OR U1569 ( .A(n805), .B(n806), .Z(n509) );
  OR U1570 ( .A(n803), .B(n804), .Z(n510) );
  NAND U1571 ( .A(n509), .B(n510), .Z(n2983) );
  OR U1572 ( .A(n1572), .B(n1573), .Z(n511) );
  NANDN U1573 ( .A(n1575), .B(n1574), .Z(n512) );
  NAND U1574 ( .A(n511), .B(n512), .Z(n2756) );
  OR U1575 ( .A(n1560), .B(n1561), .Z(n513) );
  NANDN U1576 ( .A(n1563), .B(n1562), .Z(n514) );
  NAND U1577 ( .A(n513), .B(n514), .Z(n3581) );
  OR U1578 ( .A(n1644), .B(n1645), .Z(n515) );
  NANDN U1579 ( .A(n1647), .B(n1646), .Z(n516) );
  NAND U1580 ( .A(n515), .B(n516), .Z(n3575) );
  OR U1581 ( .A(n1017), .B(n1018), .Z(n517) );
  OR U1582 ( .A(n1015), .B(n1016), .Z(n518) );
  NAND U1583 ( .A(n517), .B(n518), .Z(n2957) );
  OR U1584 ( .A(n2027), .B(n2028), .Z(n519) );
  NANDN U1585 ( .A(n2030), .B(n2029), .Z(n520) );
  NAND U1586 ( .A(n519), .B(n520), .Z(n3374) );
  OR U1587 ( .A(n1370), .B(n1371), .Z(n521) );
  NANDN U1588 ( .A(n1373), .B(n1372), .Z(n522) );
  NAND U1589 ( .A(n521), .B(n522), .Z(n3366) );
  OR U1590 ( .A(n2091), .B(n2092), .Z(n523) );
  NANDN U1591 ( .A(n2094), .B(n2093), .Z(n524) );
  NAND U1592 ( .A(n523), .B(n524), .Z(n3360) );
  OR U1593 ( .A(n1937), .B(n1938), .Z(n525) );
  OR U1594 ( .A(n1935), .B(n1936), .Z(n526) );
  NAND U1595 ( .A(n525), .B(n526), .Z(n2915) );
  OR U1596 ( .A(n1836), .B(n1837), .Z(n527) );
  NANDN U1597 ( .A(n1839), .B(n1838), .Z(n528) );
  NAND U1598 ( .A(n527), .B(n528), .Z(n3030) );
  OR U1599 ( .A(n1612), .B(n1613), .Z(n529) );
  NANDN U1600 ( .A(n1615), .B(n1614), .Z(n530) );
  NAND U1601 ( .A(n529), .B(n530), .Z(n3564) );
  OR U1602 ( .A(n1366), .B(n1367), .Z(n531) );
  NANDN U1603 ( .A(n1369), .B(n1368), .Z(n532) );
  NAND U1604 ( .A(n531), .B(n532), .Z(n2865) );
  OR U1605 ( .A(n1404), .B(n1405), .Z(n533) );
  NANDN U1606 ( .A(n1407), .B(n1406), .Z(n534) );
  NAND U1607 ( .A(n533), .B(n534), .Z(n2859) );
  OR U1608 ( .A(n1414), .B(n1415), .Z(n535) );
  NANDN U1609 ( .A(n1417), .B(n1416), .Z(n536) );
  NAND U1610 ( .A(n535), .B(n536), .Z(n3348) );
  OR U1611 ( .A(n1236), .B(n1237), .Z(n537) );
  NANDN U1612 ( .A(n1239), .B(n1238), .Z(n538) );
  NAND U1613 ( .A(n537), .B(n538), .Z(n3343) );
  OR U1614 ( .A(n2063), .B(n2064), .Z(n539) );
  OR U1615 ( .A(n2061), .B(n2062), .Z(n540) );
  NAND U1616 ( .A(n539), .B(n540), .Z(n3047) );
  OR U1617 ( .A(n2337), .B(n2338), .Z(n541) );
  NANDN U1618 ( .A(n2340), .B(n2339), .Z(n542) );
  NAND U1619 ( .A(n541), .B(n542), .Z(n3636) );
  OR U1620 ( .A(n1640), .B(n1641), .Z(n543) );
  NANDN U1621 ( .A(n1643), .B(n1642), .Z(n544) );
  NAND U1622 ( .A(n543), .B(n544), .Z(n3088) );
  OR U1623 ( .A(n741), .B(n742), .Z(n545) );
  OR U1624 ( .A(n739), .B(n740), .Z(n546) );
  NAND U1625 ( .A(n545), .B(n546), .Z(n2932) );
  OR U1626 ( .A(n1616), .B(n1617), .Z(n547) );
  NANDN U1627 ( .A(n1619), .B(n1618), .Z(n548) );
  AND U1628 ( .A(n547), .B(n548), .Z(n3544) );
  OR U1629 ( .A(n2539), .B(n2540), .Z(n549) );
  NANDN U1630 ( .A(n2542), .B(n2541), .Z(n550) );
  NAND U1631 ( .A(n549), .B(n550), .Z(n3527) );
  OR U1632 ( .A(n2365), .B(n2366), .Z(n551) );
  NANDN U1633 ( .A(n2368), .B(n2367), .Z(n552) );
  NAND U1634 ( .A(n551), .B(n552), .Z(n3523) );
  OR U1635 ( .A(n885), .B(n886), .Z(n553) );
  NANDN U1636 ( .A(n888), .B(n887), .Z(n554) );
  AND U1637 ( .A(n553), .B(n554), .Z(n2797) );
  OR U1638 ( .A(n717), .B(n718), .Z(n555) );
  NANDN U1639 ( .A(n720), .B(n719), .Z(n556) );
  NAND U1640 ( .A(n555), .B(n556), .Z(n3483) );
  OR U1641 ( .A(n871), .B(n872), .Z(n557) );
  NANDN U1642 ( .A(n874), .B(n873), .Z(n558) );
  NAND U1643 ( .A(n557), .B(n558), .Z(n3480) );
  NANDN U1644 ( .A(n735), .B(n736), .Z(n559) );
  NANDN U1645 ( .A(n738), .B(n737), .Z(n560) );
  AND U1646 ( .A(n559), .B(n560), .Z(n3021) );
  OR U1647 ( .A(n787), .B(n788), .Z(n561) );
  NANDN U1648 ( .A(n790), .B(n789), .Z(n562) );
  NAND U1649 ( .A(n561), .B(n562), .Z(n3137) );
  OR U1650 ( .A(n1160), .B(n1161), .Z(n563) );
  NANDN U1651 ( .A(n1163), .B(n1162), .Z(n564) );
  NAND U1652 ( .A(n563), .B(n564), .Z(n3661) );
  XNOR U1653 ( .A(n3646), .B(n3647), .Z(n3648) );
  OR U1654 ( .A(n2293), .B(n2294), .Z(n565) );
  NAND U1655 ( .A(n2296), .B(n2295), .Z(n566) );
  NAND U1656 ( .A(n565), .B(n566), .Z(n3307) );
  OR U1657 ( .A(n1660), .B(n1661), .Z(n567) );
  NANDN U1658 ( .A(n1662), .B(n1663), .Z(n568) );
  NAND U1659 ( .A(n567), .B(n568), .Z(n3300) );
  OR U1660 ( .A(n2321), .B(n2322), .Z(n569) );
  NANDN U1661 ( .A(n2324), .B(n2323), .Z(n570) );
  NAND U1662 ( .A(n569), .B(n570), .Z(n2970) );
  OR U1663 ( .A(n2031), .B(n2032), .Z(n571) );
  NANDN U1664 ( .A(n2034), .B(n2033), .Z(n572) );
  NAND U1665 ( .A(n571), .B(n572), .Z(n3356) );
  NANDN U1666 ( .A(n1823), .B(n1822), .Z(n573) );
  NANDN U1667 ( .A(n1824), .B(n1825), .Z(n574) );
  NAND U1668 ( .A(n573), .B(n574), .Z(n3407) );
  OR U1669 ( .A(n2705), .B(n2706), .Z(n575) );
  NANDN U1670 ( .A(n2708), .B(n2707), .Z(n576) );
  NAND U1671 ( .A(n575), .B(n576), .Z(n3396) );
  OR U1672 ( .A(n1802), .B(n1803), .Z(n577) );
  NAND U1673 ( .A(n1805), .B(n1804), .Z(n578) );
  NAND U1674 ( .A(n577), .B(n578), .Z(n3471) );
  NANDN U1675 ( .A(n1719), .B(n1718), .Z(n579) );
  NANDN U1676 ( .A(n1720), .B(n1721), .Z(n580) );
  AND U1677 ( .A(n579), .B(n580), .Z(n3330) );
  OR U1678 ( .A(n2653), .B(n2654), .Z(n581) );
  NAND U1679 ( .A(n2655), .B(n2656), .Z(n582) );
  AND U1680 ( .A(n581), .B(n582), .Z(n3512) );
  OR U1681 ( .A(n3495), .B(n3496), .Z(n583) );
  NANDN U1682 ( .A(n3497), .B(n3498), .Z(n584) );
  AND U1683 ( .A(n583), .B(n584), .Z(n3938) );
  OR U1684 ( .A(n3622), .B(n3623), .Z(n585) );
  NANDN U1685 ( .A(n3625), .B(n3624), .Z(n586) );
  AND U1686 ( .A(n585), .B(n586), .Z(n4214) );
  OR U1687 ( .A(n2892), .B(n2891), .Z(n587) );
  NANDN U1688 ( .A(n2893), .B(n2894), .Z(n588) );
  AND U1689 ( .A(n587), .B(n588), .Z(n4231) );
  OR U1690 ( .A(n2992), .B(n2991), .Z(n589) );
  NANDN U1691 ( .A(n2993), .B(n2994), .Z(n590) );
  AND U1692 ( .A(n589), .B(n590), .Z(n3927) );
  OR U1693 ( .A(n2977), .B(n2978), .Z(n591) );
  NAND U1694 ( .A(n2979), .B(n2980), .Z(n592) );
  AND U1695 ( .A(n591), .B(n592), .Z(n3923) );
  OR U1696 ( .A(n3126), .B(n3127), .Z(n593) );
  NANDN U1697 ( .A(n3129), .B(n3128), .Z(n594) );
  NAND U1698 ( .A(n593), .B(n594), .Z(n3956) );
  OR U1699 ( .A(n3034), .B(n3035), .Z(n595) );
  NANDN U1700 ( .A(n3037), .B(n3036), .Z(n596) );
  AND U1701 ( .A(n595), .B(n596), .Z(n3837) );
  OR U1702 ( .A(n3558), .B(n3559), .Z(n597) );
  NANDN U1703 ( .A(n3561), .B(n3560), .Z(n598) );
  AND U1704 ( .A(n597), .B(n598), .Z(n3843) );
  OR U1705 ( .A(n3630), .B(n3631), .Z(n599) );
  NANDN U1706 ( .A(n3633), .B(n3632), .Z(n600) );
  AND U1707 ( .A(n599), .B(n600), .Z(n4268) );
  OR U1708 ( .A(n3083), .B(n3082), .Z(n601) );
  NANDN U1709 ( .A(n3084), .B(n3085), .Z(n602) );
  AND U1710 ( .A(n601), .B(n602), .Z(n4261) );
  OR U1711 ( .A(n3067), .B(n3066), .Z(n603) );
  NANDN U1712 ( .A(n3068), .B(n3069), .Z(n604) );
  AND U1713 ( .A(n603), .B(n604), .Z(n4253) );
  OR U1714 ( .A(n2945), .B(n2946), .Z(n605) );
  NANDN U1715 ( .A(n2948), .B(n2947), .Z(n606) );
  AND U1716 ( .A(n605), .B(n606), .Z(n3907) );
  OR U1717 ( .A(n2924), .B(n2923), .Z(n607) );
  NANDN U1718 ( .A(n2925), .B(n2926), .Z(n608) );
  AND U1719 ( .A(n607), .B(n608), .Z(n3915) );
  OR U1720 ( .A(n3540), .B(n3539), .Z(n609) );
  NANDN U1721 ( .A(n3541), .B(n3542), .Z(n610) );
  AND U1722 ( .A(n609), .B(n610), .Z(n4201) );
  OR U1723 ( .A(n2901), .B(n2902), .Z(n611) );
  NANDN U1724 ( .A(n2904), .B(n2903), .Z(n612) );
  NAND U1725 ( .A(n611), .B(n612), .Z(n4250) );
  OR U1726 ( .A(n2937), .B(n2938), .Z(n613) );
  NANDN U1727 ( .A(n2940), .B(n2939), .Z(n614) );
  NAND U1728 ( .A(n613), .B(n614), .Z(n3888) );
  OR U1729 ( .A(n3163), .B(n3164), .Z(n615) );
  NAND U1730 ( .A(n3166), .B(n3165), .Z(n616) );
  NAND U1731 ( .A(n615), .B(n616), .Z(n3851) );
  OR U1732 ( .A(n2781), .B(n2782), .Z(n617) );
  NAND U1733 ( .A(n2784), .B(n2783), .Z(n618) );
  NAND U1734 ( .A(n617), .B(n618), .Z(n3828) );
  OR U1735 ( .A(n3142), .B(n3143), .Z(n619) );
  NANDN U1736 ( .A(n3145), .B(n3144), .Z(n620) );
  NAND U1737 ( .A(n619), .B(n620), .Z(n3812) );
  OR U1738 ( .A(n3057), .B(n3056), .Z(n621) );
  NANDN U1739 ( .A(n3058), .B(n3059), .Z(n622) );
  AND U1740 ( .A(n621), .B(n622), .Z(n3822) );
  NANDN U1741 ( .A(n3239), .B(n3240), .Z(n623) );
  NANDN U1742 ( .A(n3241), .B(n3242), .Z(n624) );
  NAND U1743 ( .A(n623), .B(n624), .Z(n3967) );
  NANDN U1744 ( .A(n3292), .B(n3291), .Z(n625) );
  NANDN U1745 ( .A(n3289), .B(n3290), .Z(n626) );
  NAND U1746 ( .A(n625), .B(n626), .Z(n3987) );
  OR U1747 ( .A(n1977), .B(n1978), .Z(n627) );
  OR U1748 ( .A(n1975), .B(n1976), .Z(n628) );
  NAND U1749 ( .A(n627), .B(n628), .Z(n2922) );
  OR U1750 ( .A(n1492), .B(n1493), .Z(n629) );
  OR U1751 ( .A(n1490), .B(n1491), .Z(n630) );
  AND U1752 ( .A(n629), .B(n630), .Z(n3181) );
  NAND U1753 ( .A(n1057), .B(n1058), .Z(n631) );
  NANDN U1754 ( .A(n1059), .B(n1060), .Z(n632) );
  AND U1755 ( .A(n631), .B(n632), .Z(n3000) );
  OR U1756 ( .A(n3728), .B(n3729), .Z(n633) );
  NANDN U1757 ( .A(n3731), .B(n3730), .Z(n634) );
  AND U1758 ( .A(n633), .B(n634), .Z(n4070) );
  OR U1759 ( .A(n3750), .B(n3751), .Z(n635) );
  NANDN U1760 ( .A(n3749), .B(n3748), .Z(n636) );
  AND U1761 ( .A(n635), .B(n636), .Z(n4074) );
  OR U1762 ( .A(n3026), .B(n3027), .Z(n637) );
  NAND U1763 ( .A(n3024), .B(n3025), .Z(n638) );
  AND U1764 ( .A(n637), .B(n638), .Z(n4244) );
  OR U1765 ( .A(n3169), .B(n3170), .Z(n639) );
  NANDN U1766 ( .A(n3167), .B(n3168), .Z(n640) );
  NAND U1767 ( .A(n639), .B(n640), .Z(n3982) );
  OR U1768 ( .A(n4063), .B(n4064), .Z(n641) );
  NANDN U1769 ( .A(n4066), .B(n4065), .Z(n642) );
  AND U1770 ( .A(n641), .B(n642), .Z(n4426) );
  NANDN U1771 ( .A(n4219), .B(n4220), .Z(n643) );
  NANDN U1772 ( .A(n4222), .B(n4221), .Z(n644) );
  AND U1773 ( .A(n643), .B(n644), .Z(n4408) );
  OR U1774 ( .A(n4223), .B(n4224), .Z(n645) );
  NANDN U1775 ( .A(n4225), .B(n4226), .Z(n646) );
  NAND U1776 ( .A(n645), .B(n646), .Z(n4404) );
  NANDN U1777 ( .A(n3922), .B(n3921), .Z(n647) );
  NANDN U1778 ( .A(n3919), .B(n3920), .Z(n648) );
  NAND U1779 ( .A(n647), .B(n648), .Z(n4327) );
  OR U1780 ( .A(n3833), .B(n3834), .Z(n649) );
  NANDN U1781 ( .A(n3835), .B(n3836), .Z(n650) );
  NAND U1782 ( .A(n649), .B(n650), .Z(n4336) );
  NANDN U1783 ( .A(n3906), .B(n3905), .Z(n651) );
  NANDN U1784 ( .A(n3903), .B(n3904), .Z(n652) );
  NAND U1785 ( .A(n651), .B(n652), .Z(n4344) );
  OR U1786 ( .A(n4247), .B(n4248), .Z(n653) );
  NANDN U1787 ( .A(n4245), .B(n4246), .Z(n654) );
  NAND U1788 ( .A(n653), .B(n654), .Z(n4514) );
  OR U1789 ( .A(n3894), .B(n3893), .Z(n655) );
  NANDN U1790 ( .A(n3895), .B(n3896), .Z(n656) );
  AND U1791 ( .A(n655), .B(n656), .Z(n4506) );
  OR U1792 ( .A(n4162), .B(n4163), .Z(n657) );
  NAND U1793 ( .A(n4165), .B(n4164), .Z(n658) );
  NAND U1794 ( .A(n657), .B(n658), .Z(n4355) );
  OR U1795 ( .A(n3992), .B(n3993), .Z(n659) );
  NANDN U1796 ( .A(n3995), .B(n3994), .Z(n660) );
  AND U1797 ( .A(n659), .B(n660), .Z(n4396) );
  OR U1798 ( .A(n2043), .B(n2044), .Z(n661) );
  NANDN U1799 ( .A(n2046), .B(n2045), .Z(n662) );
  AND U1800 ( .A(n661), .B(n662), .Z(n3753) );
  NAND U1801 ( .A(n2570), .B(n2569), .Z(n663) );
  NANDN U1802 ( .A(n2567), .B(n2568), .Z(n664) );
  NAND U1803 ( .A(n663), .B(n664), .Z(n3782) );
  OR U1804 ( .A(n3807), .B(n3808), .Z(n665) );
  NAND U1805 ( .A(n3809), .B(n3810), .Z(n666) );
  AND U1806 ( .A(n665), .B(n666), .Z(n4486) );
  OR U1807 ( .A(n4331), .B(n4332), .Z(n667) );
  NAND U1808 ( .A(n4334), .B(n4333), .Z(n668) );
  NAND U1809 ( .A(n667), .B(n668), .Z(n4624) );
  OR U1810 ( .A(n4310), .B(n4309), .Z(n669) );
  NANDN U1811 ( .A(n4311), .B(n4312), .Z(n670) );
  AND U1812 ( .A(n669), .B(n670), .Z(n4644) );
  OR U1813 ( .A(n4375), .B(n4376), .Z(n671) );
  NAND U1814 ( .A(n4378), .B(n4377), .Z(n672) );
  NAND U1815 ( .A(n671), .B(n672), .Z(n4651) );
  OR U1816 ( .A(n4367), .B(n4368), .Z(n673) );
  OR U1817 ( .A(n4365), .B(n4366), .Z(n674) );
  AND U1818 ( .A(n673), .B(n674), .Z(n4663) );
  OR U1819 ( .A(n1760), .B(n1761), .Z(n675) );
  NANDN U1820 ( .A(n1759), .B(n1758), .Z(n676) );
  AND U1821 ( .A(n675), .B(n676), .Z(n3210) );
  NANDN U1822 ( .A(n2640), .B(n2639), .Z(n677) );
  NANDN U1823 ( .A(n2637), .B(n2638), .Z(n678) );
  NAND U1824 ( .A(n677), .B(n678), .Z(n3684) );
  OR U1825 ( .A(n3191), .B(n3192), .Z(n679) );
  NANDN U1826 ( .A(n3190), .B(n3189), .Z(n680) );
  NAND U1827 ( .A(n679), .B(n680), .Z(n4137) );
  XOR U1828 ( .A(n4449), .B(n4448), .Z(n4450) );
  OR U1829 ( .A(n4446), .B(n4447), .Z(n681) );
  OR U1830 ( .A(n4444), .B(n4445), .Z(n682) );
  NAND U1831 ( .A(n681), .B(n682), .Z(n4567) );
  OR U1832 ( .A(n4484), .B(n4485), .Z(n683) );
  OR U1833 ( .A(n4482), .B(n4483), .Z(n684) );
  AND U1834 ( .A(n683), .B(n684), .Z(n4577) );
  OR U1835 ( .A(n4593), .B(n4594), .Z(n685) );
  NANDN U1836 ( .A(n4596), .B(n4595), .Z(n686) );
  NAND U1837 ( .A(n685), .B(n686), .Z(n4716) );
  OR U1838 ( .A(n4640), .B(n4641), .Z(n687) );
  NANDN U1839 ( .A(n4643), .B(n4642), .Z(n688) );
  AND U1840 ( .A(n687), .B(n688), .Z(n4696) );
  OR U1841 ( .A(n4292), .B(n4291), .Z(n689) );
  NANDN U1842 ( .A(n4293), .B(n4294), .Z(n690) );
  AND U1843 ( .A(n689), .B(n690), .Z(n4306) );
  OR U1844 ( .A(n4468), .B(n4469), .Z(n691) );
  NANDN U1845 ( .A(n4467), .B(n4466), .Z(n692) );
  AND U1846 ( .A(n691), .B(n692), .Z(n4581) );
  OR U1847 ( .A(n4573), .B(n4574), .Z(n693) );
  NANDN U1848 ( .A(n4572), .B(n4571), .Z(n694) );
  NAND U1849 ( .A(n693), .B(n694), .Z(n4687) );
  OR U1850 ( .A(n4705), .B(n4706), .Z(n695) );
  NANDN U1851 ( .A(n4708), .B(n4707), .Z(n696) );
  AND U1852 ( .A(n695), .B(n696), .Z(n4763) );
  OR U1853 ( .A(n4301), .B(n4302), .Z(n697) );
  NANDN U1854 ( .A(n4304), .B(n4303), .Z(n698) );
  AND U1855 ( .A(n697), .B(n698), .Z(n4676) );
  XOR U1856 ( .A(n4129), .B(n4128), .Z(n699) );
  NANDN U1857 ( .A(n4127), .B(n699), .Z(n700) );
  NAND U1858 ( .A(n4129), .B(n4128), .Z(n701) );
  AND U1859 ( .A(n700), .B(n701), .Z(n4296) );
  OR U1860 ( .A(n4774), .B(n4775), .Z(n702) );
  NANDN U1861 ( .A(n4777), .B(n4776), .Z(n703) );
  AND U1862 ( .A(n702), .B(n703), .Z(n4785) );
  NAND U1863 ( .A(n4748), .B(n4746), .Z(n704) );
  XOR U1864 ( .A(n4746), .B(n4748), .Z(n705) );
  NANDN U1865 ( .A(n4747), .B(n705), .Z(n706) );
  NAND U1866 ( .A(n704), .B(n706), .Z(n4771) );
  XNOR U1867 ( .A(x[518]), .B(y[518]), .Z(n1950) );
  XNOR U1868 ( .A(x[520]), .B(y[520]), .Z(n1948) );
  XNOR U1869 ( .A(x[522]), .B(y[522]), .Z(n1947) );
  XNOR U1870 ( .A(n1948), .B(n1947), .Z(n1949) );
  XOR U1871 ( .A(n1950), .B(n1949), .Z(n1746) );
  XNOR U1872 ( .A(x[694]), .B(y[694]), .Z(n1916) );
  XNOR U1873 ( .A(x[308]), .B(y[308]), .Z(n1914) );
  XNOR U1874 ( .A(x[696]), .B(y[696]), .Z(n1913) );
  XNOR U1875 ( .A(n1914), .B(n1913), .Z(n1915) );
  XOR U1876 ( .A(n1916), .B(n1915), .Z(n1747) );
  XOR U1877 ( .A(n1746), .B(n1747), .Z(n1748) );
  XNOR U1878 ( .A(x[524]), .B(y[524]), .Z(n1893) );
  XNOR U1879 ( .A(x[526]), .B(y[526]), .Z(n1891) );
  XNOR U1880 ( .A(x[528]), .B(y[528]), .Z(n1890) );
  XNOR U1881 ( .A(n1891), .B(n1890), .Z(n1892) );
  XOR U1882 ( .A(n1893), .B(n1892), .Z(n1749) );
  XNOR U1883 ( .A(n1748), .B(n1749), .Z(n1501) );
  XNOR U1884 ( .A(x[690]), .B(y[690]), .Z(n1924) );
  XNOR U1885 ( .A(x[304]), .B(y[304]), .Z(n1922) );
  XNOR U1886 ( .A(x[692]), .B(y[692]), .Z(n1921) );
  XNOR U1887 ( .A(n1922), .B(n1921), .Z(n1923) );
  XOR U1888 ( .A(n1924), .B(n1923), .Z(n1728) );
  XNOR U1889 ( .A(x[534]), .B(y[534]), .Z(n1906) );
  XNOR U1890 ( .A(x[158]), .B(y[158]), .Z(n1903) );
  XNOR U1891 ( .A(x[536]), .B(y[536]), .Z(n1902) );
  XNOR U1892 ( .A(n1903), .B(n1902), .Z(n1904) );
  XOR U1893 ( .A(n1906), .B(n1904), .Z(n1729) );
  XOR U1894 ( .A(n1728), .B(n1729), .Z(n1730) );
  XNOR U1895 ( .A(x[530]), .B(y[530]), .Z(n1897) );
  XNOR U1896 ( .A(x[154]), .B(y[154]), .Z(n1895) );
  XNOR U1897 ( .A(x[532]), .B(y[532]), .Z(n1894) );
  XNOR U1898 ( .A(n1895), .B(n1894), .Z(n1896) );
  XOR U1899 ( .A(n1897), .B(n1896), .Z(n1731) );
  XOR U1900 ( .A(n1730), .B(n1731), .Z(n1498) );
  XNOR U1901 ( .A(x[538]), .B(y[538]), .Z(n1912) );
  XNOR U1902 ( .A(x[540]), .B(y[540]), .Z(n1910) );
  XNOR U1903 ( .A(x[542]), .B(y[542]), .Z(n1909) );
  XNOR U1904 ( .A(n1910), .B(n1909), .Z(n1911) );
  XOR U1905 ( .A(n1912), .B(n1911), .Z(n1702) );
  XNOR U1906 ( .A(x[684]), .B(y[684]), .Z(n2204) );
  XNOR U1907 ( .A(x[686]), .B(y[686]), .Z(n2202) );
  XNOR U1908 ( .A(x[688]), .B(y[688]), .Z(n2201) );
  XNOR U1909 ( .A(n2202), .B(n2201), .Z(n2203) );
  XNOR U1910 ( .A(n2204), .B(n2203), .Z(n1703) );
  XNOR U1911 ( .A(n1702), .B(n1703), .Z(n1704) );
  XNOR U1912 ( .A(x[544]), .B(y[544]), .Z(n1920) );
  XNOR U1913 ( .A(x[546]), .B(y[546]), .Z(n1918) );
  XNOR U1914 ( .A(x[548]), .B(y[548]), .Z(n1917) );
  XNOR U1915 ( .A(n1918), .B(n1917), .Z(n1919) );
  XOR U1916 ( .A(n1920), .B(n1919), .Z(n1705) );
  XOR U1917 ( .A(n1704), .B(n1705), .Z(n1499) );
  XOR U1918 ( .A(n1498), .B(n1499), .Z(n1500) );
  XNOR U1919 ( .A(n1501), .B(n1500), .Z(n1151) );
  XNOR U1920 ( .A(x[604]), .B(y[604]), .Z(n2368) );
  XNOR U1921 ( .A(x[606]), .B(y[606]), .Z(n2366) );
  XNOR U1922 ( .A(x[608]), .B(y[608]), .Z(n2365) );
  XOR U1923 ( .A(n2366), .B(n2365), .Z(n2367) );
  XOR U1924 ( .A(n2368), .B(n2367), .Z(n2551) );
  XNOR U1925 ( .A(x[654]), .B(y[654]), .Z(n2490) );
  XNOR U1926 ( .A(x[272]), .B(y[272]), .Z(n2488) );
  XNOR U1927 ( .A(x[656]), .B(y[656]), .Z(n2487) );
  XOR U1928 ( .A(n2488), .B(n2487), .Z(n2489) );
  XOR U1929 ( .A(n2490), .B(n2489), .Z(n2550) );
  XNOR U1930 ( .A(x[598]), .B(y[598]), .Z(n2542) );
  XNOR U1931 ( .A(x[600]), .B(y[600]), .Z(n2540) );
  XNOR U1932 ( .A(x[602]), .B(y[602]), .Z(n2539) );
  XOR U1933 ( .A(n2540), .B(n2539), .Z(n2541) );
  XOR U1934 ( .A(n2542), .B(n2541), .Z(n2549) );
  XOR U1935 ( .A(n2550), .B(n2549), .Z(n2552) );
  XNOR U1936 ( .A(n2551), .B(n2552), .Z(n2558) );
  XNOR U1937 ( .A(x[614]), .B(y[614]), .Z(n2216) );
  XNOR U1938 ( .A(x[236]), .B(y[236]), .Z(n2214) );
  XNOR U1939 ( .A(x[616]), .B(y[616]), .Z(n2213) );
  XNOR U1940 ( .A(n2214), .B(n2213), .Z(n2215) );
  XNOR U1941 ( .A(n2216), .B(n2215), .Z(n1469) );
  XNOR U1942 ( .A(x[630]), .B(y[630]), .Z(n2362) );
  XNOR U1943 ( .A(x[250]), .B(y[250]), .Z(n2360) );
  XNOR U1944 ( .A(x[632]), .B(y[632]), .Z(n2359) );
  XNOR U1945 ( .A(n2360), .B(n2359), .Z(n2361) );
  XNOR U1946 ( .A(n2362), .B(n2361), .Z(n1466) );
  XNOR U1947 ( .A(x[610]), .B(y[610]), .Z(n2124) );
  XNOR U1948 ( .A(x[232]), .B(y[232]), .Z(n2122) );
  XNOR U1949 ( .A(x[612]), .B(y[612]), .Z(n2121) );
  XNOR U1950 ( .A(n2122), .B(n2121), .Z(n2123) );
  XOR U1951 ( .A(n2124), .B(n2123), .Z(n1467) );
  XNOR U1952 ( .A(n1466), .B(n1467), .Z(n1468) );
  XOR U1953 ( .A(n1469), .B(n1468), .Z(n2555) );
  XNOR U1954 ( .A(x[644]), .B(y[644]), .Z(n2530) );
  XNOR U1955 ( .A(x[646]), .B(y[646]), .Z(n2528) );
  XNOR U1956 ( .A(x[648]), .B(y[648]), .Z(n2527) );
  XNOR U1957 ( .A(n2528), .B(n2527), .Z(n2529) );
  XNOR U1958 ( .A(n2530), .B(n2529), .Z(n1099) );
  XNOR U1959 ( .A(x[650]), .B(y[650]), .Z(n2524) );
  XNOR U1960 ( .A(x[268]), .B(y[268]), .Z(n2522) );
  XNOR U1961 ( .A(x[652]), .B(y[652]), .Z(n2521) );
  XNOR U1962 ( .A(n2522), .B(n2521), .Z(n2523) );
  XNOR U1963 ( .A(n2524), .B(n2523), .Z(n1098) );
  XOR U1964 ( .A(n1099), .B(n1098), .Z(n1100) );
  XNOR U1965 ( .A(x[618]), .B(y[618]), .Z(n2372) );
  XNOR U1966 ( .A(x[620]), .B(y[620]), .Z(n2370) );
  XNOR U1967 ( .A(x[622]), .B(y[622]), .Z(n2369) );
  XNOR U1968 ( .A(n2370), .B(n2369), .Z(n2371) );
  XNOR U1969 ( .A(n2372), .B(n2371), .Z(n1101) );
  XOR U1970 ( .A(n1100), .B(n1101), .Z(n2556) );
  XOR U1971 ( .A(n2555), .B(n2556), .Z(n2557) );
  XOR U1972 ( .A(n2558), .B(n2557), .Z(n1148) );
  XNOR U1973 ( .A(x[490]), .B(y[490]), .Z(n1938) );
  XNOR U1974 ( .A(x[118]), .B(y[118]), .Z(n1936) );
  XNOR U1975 ( .A(x[492]), .B(y[492]), .Z(n1935) );
  XNOR U1976 ( .A(n1936), .B(n1935), .Z(n1937) );
  XOR U1977 ( .A(n1938), .B(n1937), .Z(n1740) );
  XNOR U1978 ( .A(x[710]), .B(y[710]), .Z(n1954) );
  XNOR U1979 ( .A(x[322]), .B(y[322]), .Z(n1952) );
  XNOR U1980 ( .A(x[712]), .B(y[712]), .Z(n1951) );
  XNOR U1981 ( .A(n1952), .B(n1951), .Z(n1953) );
  XOR U1982 ( .A(n1954), .B(n1953), .Z(n1741) );
  XOR U1983 ( .A(n1740), .B(n1741), .Z(n1742) );
  XNOR U1984 ( .A(x[494]), .B(y[494]), .Z(n1942) );
  XNOR U1985 ( .A(x[122]), .B(y[122]), .Z(n1940) );
  XNOR U1986 ( .A(x[496]), .B(y[496]), .Z(n1939) );
  XNOR U1987 ( .A(n1940), .B(n1939), .Z(n1941) );
  XOR U1988 ( .A(n1942), .B(n1941), .Z(n1743) );
  XOR U1989 ( .A(n1742), .B(n1743), .Z(n1537) );
  XNOR U1990 ( .A(x[498]), .B(y[498]), .Z(n1958) );
  XNOR U1991 ( .A(x[500]), .B(y[500]), .Z(n1956) );
  XNOR U1992 ( .A(x[502]), .B(y[502]), .Z(n1955) );
  XNOR U1993 ( .A(n1956), .B(n1955), .Z(n1957) );
  XOR U1994 ( .A(n1958), .B(n1957), .Z(n1708) );
  XNOR U1995 ( .A(x[704]), .B(y[704]), .Z(n1889) );
  XNOR U1996 ( .A(x[706]), .B(y[706]), .Z(n1887) );
  XNOR U1997 ( .A(x[708]), .B(y[708]), .Z(n1886) );
  XNOR U1998 ( .A(n1887), .B(n1886), .Z(n1888) );
  XOR U1999 ( .A(n1889), .B(n1888), .Z(n1709) );
  XOR U2000 ( .A(n1708), .B(n1709), .Z(n1710) );
  XNOR U2001 ( .A(x[504]), .B(y[504]), .Z(n1962) );
  XNOR U2002 ( .A(x[506]), .B(y[506]), .Z(n1960) );
  XNOR U2003 ( .A(x[508]), .B(y[508]), .Z(n1959) );
  XNOR U2004 ( .A(n1960), .B(n1959), .Z(n1961) );
  XOR U2005 ( .A(n1962), .B(n1961), .Z(n1711) );
  XOR U2006 ( .A(n1710), .B(n1711), .Z(n1534) );
  XNOR U2007 ( .A(x[698]), .B(y[698]), .Z(n1901) );
  XNOR U2008 ( .A(x[700]), .B(y[700]), .Z(n1899) );
  XNOR U2009 ( .A(x[702]), .B(y[702]), .Z(n1898) );
  XNOR U2010 ( .A(n1899), .B(n1898), .Z(n1900) );
  XOR U2011 ( .A(n1901), .B(n1900), .Z(n1734) );
  XNOR U2012 ( .A(x[514]), .B(y[514]), .Z(n1946) );
  XNOR U2013 ( .A(x[140]), .B(y[140]), .Z(n1944) );
  XNOR U2014 ( .A(x[516]), .B(y[516]), .Z(n1943) );
  XNOR U2015 ( .A(n1944), .B(n1943), .Z(n1945) );
  XOR U2016 ( .A(n1946), .B(n1945), .Z(n1735) );
  XOR U2017 ( .A(n1734), .B(n1735), .Z(n1736) );
  XNOR U2018 ( .A(x[510]), .B(y[510]), .Z(n966) );
  XNOR U2019 ( .A(x[136]), .B(y[136]), .Z(n964) );
  XNOR U2020 ( .A(x[512]), .B(y[512]), .Z(n963) );
  XNOR U2021 ( .A(n964), .B(n963), .Z(n965) );
  XNOR U2022 ( .A(n966), .B(n965), .Z(n1737) );
  XOR U2023 ( .A(n1736), .B(n1737), .Z(n1535) );
  XNOR U2024 ( .A(n1534), .B(n1535), .Z(n1536) );
  XOR U2025 ( .A(n1537), .B(n1536), .Z(n1149) );
  XOR U2026 ( .A(n1148), .B(n1149), .Z(n1150) );
  XNOR U2027 ( .A(n1151), .B(n1150), .Z(n1758) );
  XNOR U2028 ( .A(x[320]), .B(y[320]), .Z(n2026) );
  XNOR U2029 ( .A(x[324]), .B(y[324]), .Z(n2024) );
  XNOR U2030 ( .A(x[328]), .B(y[328]), .Z(n2023) );
  XOR U2031 ( .A(n2024), .B(n2023), .Z(n2025) );
  XOR U2032 ( .A(n2026), .B(n2025), .Z(n1047) );
  XNOR U2033 ( .A(x[330]), .B(y[330]), .Z(n2022) );
  XNOR U2034 ( .A(x[332]), .B(y[332]), .Z(n2020) );
  XNOR U2035 ( .A(x[334]), .B(y[334]), .Z(n2019) );
  XOR U2036 ( .A(n2020), .B(n2019), .Z(n2021) );
  XOR U2037 ( .A(n2022), .B(n2021), .Z(n1048) );
  XOR U2038 ( .A(n1047), .B(n1048), .Z(n1049) );
  XNOR U2039 ( .A(x[336]), .B(y[336]), .Z(n2030) );
  XNOR U2040 ( .A(x[7]), .B(y[7]), .Z(n2028) );
  XNOR U2041 ( .A(x[338]), .B(y[338]), .Z(n2027) );
  XOR U2042 ( .A(n2028), .B(n2027), .Z(n2029) );
  XOR U2043 ( .A(n2030), .B(n2029), .Z(n1050) );
  XNOR U2044 ( .A(n1049), .B(n1050), .Z(n2471) );
  XNOR U2045 ( .A(x[372]), .B(y[372]), .Z(n1861) );
  XNOR U2046 ( .A(x[374]), .B(y[374]), .Z(n1859) );
  XNOR U2047 ( .A(x[378]), .B(y[378]), .Z(n1858) );
  XNOR U2048 ( .A(n1859), .B(n1858), .Z(n1860) );
  XNOR U2049 ( .A(n1861), .B(n1860), .Z(n1531) );
  XNOR U2050 ( .A(x[368]), .B(y[368]), .Z(n1867) );
  XNOR U2051 ( .A(x[14]), .B(y[14]), .Z(n1865) );
  XNOR U2052 ( .A(x[370]), .B(y[370]), .Z(n1864) );
  XNOR U2053 ( .A(n1865), .B(n1864), .Z(n1866) );
  XNOR U2054 ( .A(n1867), .B(n1866), .Z(n1528) );
  XNOR U2055 ( .A(x[364]), .B(y[364]), .Z(n1333) );
  XNOR U2056 ( .A(x[10]), .B(y[10]), .Z(n1331) );
  XNOR U2057 ( .A(x[366]), .B(y[366]), .Z(n1330) );
  XNOR U2058 ( .A(n1331), .B(n1330), .Z(n1332) );
  XOR U2059 ( .A(n1333), .B(n1332), .Z(n1529) );
  XNOR U2060 ( .A(n1528), .B(n1529), .Z(n1530) );
  XOR U2061 ( .A(n1531), .B(n1530), .Z(n2470) );
  XNOR U2062 ( .A(x[342]), .B(y[342]), .Z(n1339) );
  XNOR U2063 ( .A(x[3]), .B(y[3]), .Z(n1337) );
  XNOR U2064 ( .A(x[346]), .B(y[346]), .Z(n1336) );
  XNOR U2065 ( .A(n1337), .B(n1336), .Z(n1338) );
  XOR U2066 ( .A(n1339), .B(n1338), .Z(n1130) );
  XNOR U2067 ( .A(x[348]), .B(y[348]), .Z(n1297) );
  XNOR U2068 ( .A(x[350]), .B(y[350]), .Z(n1295) );
  XNOR U2069 ( .A(x[352]), .B(y[352]), .Z(n1294) );
  XNOR U2070 ( .A(n1295), .B(n1294), .Z(n1296) );
  XOR U2071 ( .A(n1297), .B(n1296), .Z(n1131) );
  XOR U2072 ( .A(n1130), .B(n1131), .Z(n1132) );
  XNOR U2073 ( .A(x[354]), .B(y[354]), .Z(n1301) );
  XNOR U2074 ( .A(x[356]), .B(y[356]), .Z(n1299) );
  XNOR U2075 ( .A(x[360]), .B(y[360]), .Z(n1298) );
  XNOR U2076 ( .A(n1299), .B(n1298), .Z(n1300) );
  XOR U2077 ( .A(n1301), .B(n1300), .Z(n1133) );
  XOR U2078 ( .A(n1132), .B(n1133), .Z(n2469) );
  XOR U2079 ( .A(n2470), .B(n2469), .Z(n2472) );
  XNOR U2080 ( .A(n2471), .B(n2472), .Z(n710) );
  XNOR U2081 ( .A(x[240]), .B(y[240]), .Z(n724) );
  XNOR U2082 ( .A(x[75]), .B(y[75]), .Z(n722) );
  XNOR U2083 ( .A(x[242]), .B(y[242]), .Z(n721) );
  XOR U2084 ( .A(n722), .B(n721), .Z(n723) );
  XNOR U2085 ( .A(n724), .B(n723), .Z(n2324) );
  XNOR U2086 ( .A(x[234]), .B(y[234]), .Z(n752) );
  XNOR U2087 ( .A(x[79]), .B(y[79]), .Z(n750) );
  XNOR U2088 ( .A(x[238]), .B(y[238]), .Z(n749) );
  XNOR U2089 ( .A(n750), .B(n749), .Z(n751) );
  XOR U2090 ( .A(n752), .B(n751), .Z(n2321) );
  XNOR U2091 ( .A(x[226]), .B(y[226]), .Z(n746) );
  XNOR U2092 ( .A(x[228]), .B(y[228]), .Z(n744) );
  XNOR U2093 ( .A(x[230]), .B(y[230]), .Z(n743) );
  XNOR U2094 ( .A(n744), .B(n743), .Z(n745) );
  XOR U2095 ( .A(n746), .B(n745), .Z(n2322) );
  XOR U2096 ( .A(n2321), .B(n2322), .Z(n2323) );
  XOR U2097 ( .A(n2324), .B(n2323), .Z(n1817) );
  XNOR U2098 ( .A(x[260]), .B(y[260]), .Z(n908) );
  XNOR U2099 ( .A(x[61]), .B(y[61]), .Z(n906) );
  XNOR U2100 ( .A(x[262]), .B(y[262]), .Z(n905) );
  XNOR U2101 ( .A(n906), .B(n905), .Z(n907) );
  XNOR U2102 ( .A(n908), .B(n907), .Z(n1825) );
  XNOR U2103 ( .A(x[252]), .B(y[252]), .Z(n930) );
  XNOR U2104 ( .A(x[256]), .B(y[256]), .Z(n928) );
  XNOR U2105 ( .A(x[258]), .B(y[258]), .Z(n927) );
  XNOR U2106 ( .A(n928), .B(n927), .Z(n929) );
  XNOR U2107 ( .A(n930), .B(n929), .Z(n1822) );
  XNOR U2108 ( .A(x[244]), .B(y[244]), .Z(n960) );
  XNOR U2109 ( .A(x[246]), .B(y[246]), .Z(n958) );
  XNOR U2110 ( .A(x[248]), .B(y[248]), .Z(n957) );
  XNOR U2111 ( .A(n958), .B(n957), .Z(n959) );
  XOR U2112 ( .A(n960), .B(n959), .Z(n1823) );
  XOR U2113 ( .A(n1822), .B(n1823), .Z(n1824) );
  XNOR U2114 ( .A(n1825), .B(n1824), .Z(n1816) );
  XOR U2115 ( .A(n1817), .B(n1816), .Z(n1819) );
  XNOR U2116 ( .A(x[220]), .B(y[220]), .Z(n802) );
  XNOR U2117 ( .A(x[222]), .B(y[222]), .Z(n800) );
  XNOR U2118 ( .A(x[224]), .B(y[224]), .Z(n799) );
  XOR U2119 ( .A(n800), .B(n799), .Z(n801) );
  XNOR U2120 ( .A(n802), .B(n801), .Z(n2343) );
  XNOR U2121 ( .A(x[212]), .B(y[212]), .Z(n2098) );
  XNOR U2122 ( .A(x[93]), .B(y[93]), .Z(n2096) );
  XNOR U2123 ( .A(x[216]), .B(y[216]), .Z(n2095) );
  XOR U2124 ( .A(n2096), .B(n2095), .Z(n2097) );
  XNOR U2125 ( .A(n2098), .B(n2097), .Z(n2341) );
  XNOR U2126 ( .A(x[208]), .B(y[208]), .Z(n1381) );
  XNOR U2127 ( .A(x[97]), .B(y[97]), .Z(n1379) );
  XNOR U2128 ( .A(x[210]), .B(y[210]), .Z(n1378) );
  XOR U2129 ( .A(n1379), .B(n1378), .Z(n1380) );
  XNOR U2130 ( .A(n1381), .B(n1380), .Z(n2342) );
  XNOR U2131 ( .A(n2341), .B(n2342), .Z(n2344) );
  XNOR U2132 ( .A(n2343), .B(n2344), .Z(n1818) );
  XOR U2133 ( .A(n1819), .B(n1818), .Z(n707) );
  XNOR U2134 ( .A(x[264]), .B(y[264]), .Z(n830) );
  XNOR U2135 ( .A(x[57]), .B(y[57]), .Z(n828) );
  XNOR U2136 ( .A(x[266]), .B(y[266]), .Z(n827) );
  XOR U2137 ( .A(n828), .B(n827), .Z(n829) );
  XOR U2138 ( .A(n830), .B(n829), .Z(n998) );
  XNOR U2139 ( .A(x[270]), .B(y[270]), .Z(n914) );
  XNOR U2140 ( .A(x[274]), .B(y[274]), .Z(n912) );
  XNOR U2141 ( .A(x[276]), .B(y[276]), .Z(n911) );
  XOR U2142 ( .A(n912), .B(n911), .Z(n913) );
  XNOR U2143 ( .A(n914), .B(n913), .Z(n997) );
  XNOR U2144 ( .A(n998), .B(n997), .Z(n1000) );
  XNOR U2145 ( .A(x[278]), .B(y[278]), .Z(n826) );
  XNOR U2146 ( .A(x[280]), .B(y[280]), .Z(n824) );
  XNOR U2147 ( .A(x[282]), .B(y[282]), .Z(n823) );
  XOR U2148 ( .A(n824), .B(n823), .Z(n825) );
  XNOR U2149 ( .A(n826), .B(n825), .Z(n999) );
  XOR U2150 ( .A(n1000), .B(n999), .Z(n2046) );
  XNOR U2151 ( .A(x[302]), .B(y[302]), .Z(n2010) );
  XNOR U2152 ( .A(x[306]), .B(y[306]), .Z(n2008) );
  XNOR U2153 ( .A(x[310]), .B(y[310]), .Z(n2007) );
  XNOR U2154 ( .A(n2008), .B(n2007), .Z(n2009) );
  XOR U2155 ( .A(n2010), .B(n2009), .Z(n1092) );
  XNOR U2156 ( .A(x[312]), .B(y[312]), .Z(n2018) );
  XNOR U2157 ( .A(x[25]), .B(y[25]), .Z(n2016) );
  XNOR U2158 ( .A(x[314]), .B(y[314]), .Z(n2015) );
  XNOR U2159 ( .A(n2016), .B(n2015), .Z(n2017) );
  XOR U2160 ( .A(n2018), .B(n2017), .Z(n1093) );
  XOR U2161 ( .A(n1092), .B(n1093), .Z(n1094) );
  XNOR U2162 ( .A(x[316]), .B(y[316]), .Z(n2014) );
  XNOR U2163 ( .A(x[21]), .B(y[21]), .Z(n2012) );
  XNOR U2164 ( .A(x[318]), .B(y[318]), .Z(n2011) );
  XNOR U2165 ( .A(n2012), .B(n2011), .Z(n2013) );
  XOR U2166 ( .A(n2014), .B(n2013), .Z(n1095) );
  XOR U2167 ( .A(n1094), .B(n1095), .Z(n2043) );
  XNOR U2168 ( .A(x[284]), .B(y[284]), .Z(n888) );
  XNOR U2169 ( .A(x[43]), .B(y[43]), .Z(n886) );
  XNOR U2170 ( .A(x[288]), .B(y[288]), .Z(n885) );
  XOR U2171 ( .A(n886), .B(n885), .Z(n887) );
  XOR U2172 ( .A(n888), .B(n887), .Z(n974) );
  XNOR U2173 ( .A(x[292]), .B(y[292]), .Z(n2034) );
  XNOR U2174 ( .A(x[39]), .B(y[39]), .Z(n2032) );
  XNOR U2175 ( .A(x[294]), .B(y[294]), .Z(n2031) );
  XOR U2176 ( .A(n2032), .B(n2031), .Z(n2033) );
  XNOR U2177 ( .A(n2034), .B(n2033), .Z(n973) );
  XNOR U2178 ( .A(n974), .B(n973), .Z(n976) );
  XNOR U2179 ( .A(x[296]), .B(y[296]), .Z(n2038) );
  XNOR U2180 ( .A(x[298]), .B(y[298]), .Z(n2036) );
  XNOR U2181 ( .A(x[300]), .B(y[300]), .Z(n2035) );
  XOR U2182 ( .A(n2036), .B(n2035), .Z(n2037) );
  XNOR U2183 ( .A(n2038), .B(n2037), .Z(n975) );
  XOR U2184 ( .A(n976), .B(n975), .Z(n2044) );
  XOR U2185 ( .A(n2043), .B(n2044), .Z(n2045) );
  XOR U2186 ( .A(n2046), .B(n2045), .Z(n708) );
  XNOR U2187 ( .A(n707), .B(n708), .Z(n709) );
  XOR U2188 ( .A(n710), .B(n709), .Z(n1759) );
  XOR U2189 ( .A(n1758), .B(n1759), .Z(n1760) );
  XNOR U2190 ( .A(x[167]), .B(y[167]), .Z(n2256) );
  XNOR U2191 ( .A(x[163]), .B(y[163]), .Z(n2254) );
  XNOR U2192 ( .A(x[483]), .B(y[483]), .Z(n2253) );
  XOR U2193 ( .A(n2254), .B(n2253), .Z(n2255) );
  XOR U2194 ( .A(n2256), .B(n2255), .Z(n1427) );
  XNOR U2195 ( .A(x[161]), .B(y[161]), .Z(n2278) );
  XNOR U2196 ( .A(x[159]), .B(y[159]), .Z(n2276) );
  XNOR U2197 ( .A(x[755]), .B(y[755]), .Z(n2275) );
  XNOR U2198 ( .A(n2276), .B(n2275), .Z(n2277) );
  XNOR U2199 ( .A(n2278), .B(n2277), .Z(n1426) );
  XOR U2200 ( .A(n1427), .B(n1426), .Z(n1428) );
  XNOR U2201 ( .A(x[157]), .B(y[157]), .Z(n2272) );
  XNOR U2202 ( .A(x[155]), .B(y[155]), .Z(n2270) );
  XNOR U2203 ( .A(x[479]), .B(y[479]), .Z(n2269) );
  XNOR U2204 ( .A(n2270), .B(n2269), .Z(n2271) );
  XNOR U2205 ( .A(n2272), .B(n2271), .Z(n1429) );
  XOR U2206 ( .A(n1428), .B(n1429), .Z(n1793) );
  XNOR U2207 ( .A(x[153]), .B(y[153]), .Z(n2284) );
  XNOR U2208 ( .A(x[149]), .B(y[149]), .Z(n2282) );
  XNOR U2209 ( .A(x[757]), .B(y[757]), .Z(n2281) );
  XNOR U2210 ( .A(n2282), .B(n2281), .Z(n2283) );
  XNOR U2211 ( .A(n2284), .B(n2283), .Z(n2082) );
  XNOR U2212 ( .A(x[145]), .B(y[145]), .Z(n2306) );
  XNOR U2213 ( .A(x[143]), .B(y[143]), .Z(n2304) );
  XNOR U2214 ( .A(x[475]), .B(y[475]), .Z(n2303) );
  XNOR U2215 ( .A(n2304), .B(n2303), .Z(n2305) );
  XNOR U2216 ( .A(n2306), .B(n2305), .Z(n2081) );
  XOR U2217 ( .A(n2082), .B(n2081), .Z(n2083) );
  XNOR U2218 ( .A(x[141]), .B(y[141]), .Z(n2300) );
  XNOR U2219 ( .A(x[139]), .B(y[139]), .Z(n2298) );
  XNOR U2220 ( .A(x[759]), .B(y[759]), .Z(n2297) );
  XNOR U2221 ( .A(n2298), .B(n2297), .Z(n2299) );
  XNOR U2222 ( .A(n2300), .B(n2299), .Z(n2084) );
  XOR U2223 ( .A(n2083), .B(n2084), .Z(n1790) );
  XNOR U2224 ( .A(x[137]), .B(y[137]), .Z(n2312) );
  XNOR U2225 ( .A(x[135]), .B(y[135]), .Z(n2310) );
  XNOR U2226 ( .A(x[471]), .B(y[471]), .Z(n2309) );
  XOR U2227 ( .A(n2310), .B(n2309), .Z(n2311) );
  XOR U2228 ( .A(n2312), .B(n2311), .Z(n1277) );
  XNOR U2229 ( .A(x[131]), .B(y[131]), .Z(n2616) );
  XNOR U2230 ( .A(x[127]), .B(y[127]), .Z(n2614) );
  XNOR U2231 ( .A(x[761]), .B(y[761]), .Z(n2613) );
  XOR U2232 ( .A(n2614), .B(n2613), .Z(n2615) );
  XNOR U2233 ( .A(n2616), .B(n2615), .Z(n1276) );
  XNOR U2234 ( .A(n1277), .B(n1276), .Z(n1279) );
  XNOR U2235 ( .A(x[125]), .B(y[125]), .Z(n2624) );
  XNOR U2236 ( .A(x[123]), .B(y[123]), .Z(n2622) );
  XNOR U2237 ( .A(x[467]), .B(y[467]), .Z(n2621) );
  XOR U2238 ( .A(n2622), .B(n2621), .Z(n2623) );
  XNOR U2239 ( .A(n2624), .B(n2623), .Z(n1278) );
  XOR U2240 ( .A(n1279), .B(n1278), .Z(n1791) );
  XNOR U2241 ( .A(n1790), .B(n1791), .Z(n1792) );
  XNOR U2242 ( .A(n1793), .B(n1792), .Z(n1781) );
  XNOR U2243 ( .A(x[121]), .B(y[121]), .Z(n2620) );
  XNOR U2244 ( .A(x[119]), .B(y[119]), .Z(n2618) );
  XNOR U2245 ( .A(x[763]), .B(y[763]), .Z(n2617) );
  XOR U2246 ( .A(n2618), .B(n2617), .Z(n2619) );
  XOR U2247 ( .A(n2620), .B(n2619), .Z(n1283) );
  XNOR U2248 ( .A(x[117]), .B(y[117]), .Z(n2720) );
  XNOR U2249 ( .A(x[113]), .B(y[113]), .Z(n2718) );
  XNOR U2250 ( .A(x[463]), .B(y[463]), .Z(n2717) );
  XOR U2251 ( .A(n2718), .B(n2717), .Z(n2719) );
  XNOR U2252 ( .A(n2720), .B(n2719), .Z(n1282) );
  XNOR U2253 ( .A(n1283), .B(n1282), .Z(n1285) );
  XNOR U2254 ( .A(x[109]), .B(y[109]), .Z(n2716) );
  XNOR U2255 ( .A(x[107]), .B(y[107]), .Z(n2714) );
  XNOR U2256 ( .A(x[765]), .B(y[765]), .Z(n2713) );
  XOR U2257 ( .A(n2714), .B(n2713), .Z(n2715) );
  XNOR U2258 ( .A(n2716), .B(n2715), .Z(n1284) );
  XOR U2259 ( .A(n1285), .B(n1284), .Z(n1771) );
  XNOR U2260 ( .A(x[89]), .B(y[89]), .Z(n1833) );
  XNOR U2261 ( .A(x[87]), .B(y[87]), .Z(n1831) );
  XNOR U2262 ( .A(x[769]), .B(y[769]), .Z(n1830) );
  XNOR U2263 ( .A(n1831), .B(n1830), .Z(n1832) );
  XNOR U2264 ( .A(n1833), .B(n1832), .Z(n1409) );
  XNOR U2265 ( .A(x[85]), .B(y[85]), .Z(n2408) );
  XNOR U2266 ( .A(x[83]), .B(y[83]), .Z(n2406) );
  XNOR U2267 ( .A(x[451]), .B(y[451]), .Z(n2405) );
  XNOR U2268 ( .A(n2406), .B(n2405), .Z(n2407) );
  XNOR U2269 ( .A(n2408), .B(n2407), .Z(n1408) );
  XOR U2270 ( .A(n1409), .B(n1408), .Z(n1410) );
  XNOR U2271 ( .A(x[81]), .B(y[81]), .Z(n2402) );
  XNOR U2272 ( .A(x[77]), .B(y[77]), .Z(n2400) );
  XNOR U2273 ( .A(x[771]), .B(y[771]), .Z(n2399) );
  XNOR U2274 ( .A(n2400), .B(n2399), .Z(n2401) );
  XNOR U2275 ( .A(n2402), .B(n2401), .Z(n1411) );
  XOR U2276 ( .A(n1410), .B(n1411), .Z(n1768) );
  XNOR U2277 ( .A(x[95]), .B(y[95]), .Z(n1839) );
  XNOR U2278 ( .A(x[91]), .B(y[91]), .Z(n1837) );
  XNOR U2279 ( .A(x[455]), .B(y[455]), .Z(n1836) );
  XOR U2280 ( .A(n1837), .B(n1836), .Z(n1838) );
  XNOR U2281 ( .A(n1839), .B(n1838), .Z(n1310) );
  XNOR U2282 ( .A(x[101]), .B(y[101]), .Z(n1829) );
  XNOR U2283 ( .A(x[99]), .B(y[99]), .Z(n1827) );
  XNOR U2284 ( .A(x[767]), .B(y[767]), .Z(n1826) );
  XOR U2285 ( .A(n1827), .B(n1826), .Z(n1828) );
  XNOR U2286 ( .A(n1829), .B(n1828), .Z(n1308) );
  XNOR U2287 ( .A(x[105]), .B(y[105]), .Z(n2724) );
  XNOR U2288 ( .A(x[103]), .B(y[103]), .Z(n2722) );
  XNOR U2289 ( .A(x[459]), .B(y[459]), .Z(n2721) );
  XOR U2290 ( .A(n2722), .B(n2721), .Z(n2723) );
  XNOR U2291 ( .A(n2724), .B(n2723), .Z(n1309) );
  XNOR U2292 ( .A(n1308), .B(n1309), .Z(n1311) );
  XNOR U2293 ( .A(n1310), .B(n1311), .Z(n1769) );
  XNOR U2294 ( .A(n1768), .B(n1769), .Z(n1770) );
  XOR U2295 ( .A(n1771), .B(n1770), .Z(n1780) );
  XOR U2296 ( .A(n1781), .B(n1780), .Z(n1783) );
  XNOR U2297 ( .A(x[73]), .B(y[73]), .Z(n2414) );
  XNOR U2298 ( .A(x[71]), .B(y[71]), .Z(n2412) );
  XNOR U2299 ( .A(x[447]), .B(y[447]), .Z(n2411) );
  XNOR U2300 ( .A(n2412), .B(n2411), .Z(n2413) );
  XNOR U2301 ( .A(n2414), .B(n2413), .Z(n1585) );
  XNOR U2302 ( .A(x[69]), .B(y[69]), .Z(n2334) );
  XNOR U2303 ( .A(x[67]), .B(y[67]), .Z(n2332) );
  XNOR U2304 ( .A(x[773]), .B(y[773]), .Z(n2331) );
  XNOR U2305 ( .A(n2332), .B(n2331), .Z(n2333) );
  XNOR U2306 ( .A(n2334), .B(n2333), .Z(n1584) );
  XOR U2307 ( .A(n1585), .B(n1584), .Z(n1586) );
  XNOR U2308 ( .A(x[65]), .B(y[65]), .Z(n2328) );
  XNOR U2309 ( .A(x[63]), .B(y[63]), .Z(n2326) );
  XNOR U2310 ( .A(x[443]), .B(y[443]), .Z(n2325) );
  XNOR U2311 ( .A(n2326), .B(n2325), .Z(n2327) );
  XNOR U2312 ( .A(n2328), .B(n2327), .Z(n1587) );
  XOR U2313 ( .A(n1586), .B(n1587), .Z(n2574) );
  XNOR U2314 ( .A(x[45]), .B(y[45]), .Z(n1159) );
  XNOR U2315 ( .A(x[41]), .B(y[41]), .Z(n1157) );
  XNOR U2316 ( .A(x[435]), .B(y[435]), .Z(n1156) );
  XNOR U2317 ( .A(n1157), .B(n1156), .Z(n1158) );
  XOR U2318 ( .A(n1159), .B(n1158), .Z(n1554) );
  XNOR U2319 ( .A(x[37]), .B(y[37]), .Z(n2152) );
  XNOR U2320 ( .A(x[35]), .B(y[35]), .Z(n2150) );
  XNOR U2321 ( .A(x[779]), .B(y[779]), .Z(n2149) );
  XNOR U2322 ( .A(n2150), .B(n2149), .Z(n2151) );
  XOR U2323 ( .A(n2152), .B(n2151), .Z(n1555) );
  XNOR U2324 ( .A(n1554), .B(n1555), .Z(n1557) );
  XNOR U2325 ( .A(x[33]), .B(y[33]), .Z(n2148) );
  XNOR U2326 ( .A(x[31]), .B(y[31]), .Z(n2146) );
  XNOR U2327 ( .A(x[431]), .B(y[431]), .Z(n2145) );
  XNOR U2328 ( .A(n2146), .B(n2145), .Z(n2147) );
  XOR U2329 ( .A(n2148), .B(n2147), .Z(n1556) );
  XOR U2330 ( .A(n1557), .B(n1556), .Z(n2571) );
  XNOR U2331 ( .A(x[49]), .B(y[49]), .Z(n1163) );
  XNOR U2332 ( .A(x[47]), .B(y[47]), .Z(n1161) );
  XNOR U2333 ( .A(x[777]), .B(y[777]), .Z(n1160) );
  XOR U2334 ( .A(n1161), .B(n1160), .Z(n1162) );
  XOR U2335 ( .A(n1163), .B(n1162), .Z(n1291) );
  XNOR U2336 ( .A(x[53]), .B(y[53]), .Z(n1155) );
  XNOR U2337 ( .A(x[51]), .B(y[51]), .Z(n1153) );
  XNOR U2338 ( .A(x[439]), .B(y[439]), .Z(n1152) );
  XOR U2339 ( .A(n1153), .B(n1152), .Z(n1154) );
  XOR U2340 ( .A(n1155), .B(n1154), .Z(n1288) );
  XNOR U2341 ( .A(x[59]), .B(y[59]), .Z(n2340) );
  XNOR U2342 ( .A(x[55]), .B(y[55]), .Z(n2338) );
  XNOR U2343 ( .A(x[775]), .B(y[775]), .Z(n2337) );
  XOR U2344 ( .A(n2338), .B(n2337), .Z(n2339) );
  XNOR U2345 ( .A(n2340), .B(n2339), .Z(n1289) );
  XNOR U2346 ( .A(n1288), .B(n1289), .Z(n1290) );
  XNOR U2347 ( .A(n1291), .B(n1290), .Z(n2572) );
  XNOR U2348 ( .A(n2571), .B(n2572), .Z(n2573) );
  XNOR U2349 ( .A(n2574), .B(n2573), .Z(n1782) );
  XOR U2350 ( .A(n1783), .B(n1782), .Z(n1761) );
  XOR U2351 ( .A(n1760), .B(n1761), .Z(n1812) );
  XNOR U2352 ( .A(x[485]), .B(y[485]), .Z(n1421) );
  XNOR U2353 ( .A(x[477]), .B(y[477]), .Z(n1419) );
  XNOR U2354 ( .A(x[481]), .B(y[481]), .Z(n1418) );
  XOR U2355 ( .A(n1419), .B(n1418), .Z(n1420) );
  XOR U2356 ( .A(n1421), .B(n1420), .Z(n918) );
  XNOR U2357 ( .A(x[168]), .B(y[168]), .Z(n1377) );
  XNOR U2358 ( .A(x[170]), .B(y[170]), .Z(n1375) );
  XNOR U2359 ( .A(x[174]), .B(y[174]), .Z(n1374) );
  XOR U2360 ( .A(n1375), .B(n1374), .Z(n1376) );
  XOR U2361 ( .A(n1377), .B(n1376), .Z(n915) );
  XNOR U2362 ( .A(x[497]), .B(y[497]), .Z(n1417) );
  XNOR U2363 ( .A(x[489]), .B(y[489]), .Z(n1415) );
  XNOR U2364 ( .A(x[493]), .B(y[493]), .Z(n1414) );
  XOR U2365 ( .A(n1415), .B(n1414), .Z(n1416) );
  XNOR U2366 ( .A(n1417), .B(n1416), .Z(n916) );
  XNOR U2367 ( .A(n915), .B(n916), .Z(n917) );
  XNOR U2368 ( .A(n918), .B(n917), .Z(n1797) );
  XNOR U2369 ( .A(x[54]), .B(y[54]), .Z(n1619) );
  XNOR U2370 ( .A(x[56]), .B(y[56]), .Z(n1617) );
  XNOR U2371 ( .A(x[201]), .B(y[201]), .Z(n1616) );
  XOR U2372 ( .A(n1617), .B(n1616), .Z(n1618) );
  XNOR U2373 ( .A(n1619), .B(n1618), .Z(n1180) );
  XNOR U2374 ( .A(x[200]), .B(y[200]), .Z(n1623) );
  XNOR U2375 ( .A(x[202]), .B(y[202]), .Z(n1621) );
  XNOR U2376 ( .A(x[799]), .B(y[799]), .Z(n1620) );
  XOR U2377 ( .A(n1621), .B(n1620), .Z(n1622) );
  XNOR U2378 ( .A(n1623), .B(n1622), .Z(n1178) );
  XNOR U2379 ( .A(x[798]), .B(y[798]), .Z(n1063) );
  XOR U2380 ( .A(x[204]), .B(y[204]), .Z(n1061) );
  XNOR U2381 ( .A(oglobal[0]), .B(n1061), .Z(n1062) );
  XOR U2382 ( .A(n1063), .B(n1062), .Z(n1179) );
  XNOR U2383 ( .A(n1178), .B(n1179), .Z(n1181) );
  XNOR U2384 ( .A(n1180), .B(n1181), .Z(n1796) );
  XOR U2385 ( .A(n1797), .B(n1796), .Z(n1798) );
  XNOR U2386 ( .A(x[509]), .B(y[509]), .Z(n1407) );
  XNOR U2387 ( .A(x[501]), .B(y[501]), .Z(n1405) );
  XNOR U2388 ( .A(x[505]), .B(y[505]), .Z(n1404) );
  XOR U2389 ( .A(n1405), .B(n1404), .Z(n1406) );
  XNOR U2390 ( .A(n1407), .B(n1406), .Z(n923) );
  XNOR U2391 ( .A(x[754]), .B(y[754]), .Z(n1425) );
  XNOR U2392 ( .A(x[362]), .B(y[362]), .Z(n1423) );
  XNOR U2393 ( .A(x[756]), .B(y[756]), .Z(n1422) );
  XOR U2394 ( .A(n1423), .B(n1422), .Z(n1424) );
  XNOR U2395 ( .A(n1425), .B(n1424), .Z(n921) );
  XNOR U2396 ( .A(x[521]), .B(y[521]), .Z(n1403) );
  XNOR U2397 ( .A(x[513]), .B(y[513]), .Z(n1401) );
  XNOR U2398 ( .A(x[517]), .B(y[517]), .Z(n1400) );
  XOR U2399 ( .A(n1401), .B(n1400), .Z(n1402) );
  XNOR U2400 ( .A(n1403), .B(n1402), .Z(n922) );
  XNOR U2401 ( .A(n921), .B(n922), .Z(n924) );
  XNOR U2402 ( .A(n923), .B(n924), .Z(n1799) );
  XOR U2403 ( .A(n1798), .B(n1799), .Z(n2637) );
  XNOR U2404 ( .A(x[573]), .B(y[573]), .Z(n1143) );
  XNOR U2405 ( .A(x[569]), .B(y[569]), .Z(n1141) );
  XNOR U2406 ( .A(x[571]), .B(y[571]), .Z(n1140) );
  XOR U2407 ( .A(n1141), .B(n1140), .Z(n1142) );
  XOR U2408 ( .A(n1143), .B(n1142), .Z(n735) );
  XNOR U2409 ( .A(x[764]), .B(y[764]), .Z(n1519) );
  XNOR U2410 ( .A(x[766]), .B(y[766]), .Z(n1517) );
  XNOR U2411 ( .A(x[768]), .B(y[768]), .Z(n1516) );
  XOR U2412 ( .A(n1517), .B(n1516), .Z(n1518) );
  XNOR U2413 ( .A(n1519), .B(n1518), .Z(n736) );
  XOR U2414 ( .A(n735), .B(n736), .Z(n738) );
  XNOR U2415 ( .A(x[567]), .B(y[567]), .Z(n1147) );
  XNOR U2416 ( .A(x[563]), .B(y[563]), .Z(n1145) );
  XNOR U2417 ( .A(x[565]), .B(y[565]), .Z(n1144) );
  XOR U2418 ( .A(n1145), .B(n1144), .Z(n1146) );
  XNOR U2419 ( .A(n1147), .B(n1146), .Z(n737) );
  XOR U2420 ( .A(n738), .B(n737), .Z(n1776) );
  XNOR U2421 ( .A(x[561]), .B(y[561]), .Z(n1523) );
  XNOR U2422 ( .A(x[557]), .B(y[557]), .Z(n1521) );
  XNOR U2423 ( .A(x[559]), .B(y[559]), .Z(n1520) );
  XOR U2424 ( .A(n1521), .B(n1520), .Z(n1522) );
  XOR U2425 ( .A(n1523), .B(n1522), .Z(n969) );
  XNOR U2426 ( .A(x[555]), .B(y[555]), .Z(n1527) );
  XNOR U2427 ( .A(x[551]), .B(y[551]), .Z(n1525) );
  XNOR U2428 ( .A(x[553]), .B(y[553]), .Z(n1524) );
  XOR U2429 ( .A(n1525), .B(n1524), .Z(n1526) );
  XOR U2430 ( .A(n1527), .B(n1526), .Z(n970) );
  XOR U2431 ( .A(n969), .B(n970), .Z(n971) );
  XNOR U2432 ( .A(x[144]), .B(y[144]), .Z(n2094) );
  XNOR U2433 ( .A(x[146]), .B(y[146]), .Z(n2092) );
  XNOR U2434 ( .A(x[148]), .B(y[148]), .Z(n2091) );
  XOR U2435 ( .A(n2092), .B(n2091), .Z(n2093) );
  XOR U2436 ( .A(n2094), .B(n2093), .Z(n972) );
  XNOR U2437 ( .A(n971), .B(n972), .Z(n1774) );
  XNOR U2438 ( .A(x[669]), .B(y[669]), .Z(n1513) );
  XNOR U2439 ( .A(x[667]), .B(y[667]), .Z(n1511) );
  XNOR U2440 ( .A(x[679]), .B(y[679]), .Z(n1510) );
  XOR U2441 ( .A(n1511), .B(n1510), .Z(n1512) );
  XOR U2442 ( .A(n1513), .B(n1512), .Z(n834) );
  XNOR U2443 ( .A(x[794]), .B(y[794]), .Z(n1633) );
  XNOR U2444 ( .A(x[796]), .B(y[796]), .Z(n1631) );
  XNOR U2445 ( .A(x[797]), .B(y[797]), .Z(n1630) );
  XOR U2446 ( .A(n1631), .B(n1630), .Z(n1632) );
  XOR U2447 ( .A(n1633), .B(n1632), .Z(n831) );
  XNOR U2448 ( .A(x[691]), .B(y[691]), .Z(n1509) );
  XNOR U2449 ( .A(x[673]), .B(y[673]), .Z(n1507) );
  XNOR U2450 ( .A(x[677]), .B(y[677]), .Z(n1506) );
  XOR U2451 ( .A(n1507), .B(n1506), .Z(n1508) );
  XNOR U2452 ( .A(n1509), .B(n1508), .Z(n832) );
  XNOR U2453 ( .A(n831), .B(n832), .Z(n833) );
  XNOR U2454 ( .A(n834), .B(n833), .Z(n1775) );
  XNOR U2455 ( .A(n1774), .B(n1775), .Z(n1777) );
  XNOR U2456 ( .A(n1776), .B(n1777), .Z(n2638) );
  XNOR U2457 ( .A(n2637), .B(n2638), .Z(n2639) );
  XNOR U2458 ( .A(x[633]), .B(y[633]), .Z(n1579) );
  XNOR U2459 ( .A(x[631]), .B(y[631]), .Z(n1577) );
  XNOR U2460 ( .A(x[719]), .B(y[719]), .Z(n1576) );
  XOR U2461 ( .A(n1577), .B(n1576), .Z(n1578) );
  XOR U2462 ( .A(n1579), .B(n1578), .Z(n717) );
  XNOR U2463 ( .A(x[778]), .B(y[778]), .Z(n1667) );
  XNOR U2464 ( .A(x[780]), .B(y[780]), .Z(n1665) );
  XNOR U2465 ( .A(x[782]), .B(y[782]), .Z(n1664) );
  XOR U2466 ( .A(n1665), .B(n1664), .Z(n1666) );
  XOR U2467 ( .A(n1667), .B(n1666), .Z(n718) );
  XOR U2468 ( .A(n717), .B(n718), .Z(n719) );
  XNOR U2469 ( .A(x[629]), .B(y[629]), .Z(n1583) );
  XNOR U2470 ( .A(x[627]), .B(y[627]), .Z(n1581) );
  XNOR U2471 ( .A(x[721]), .B(y[721]), .Z(n1580) );
  XOR U2472 ( .A(n1581), .B(n1580), .Z(n1582) );
  XOR U2473 ( .A(n1583), .B(n1582), .Z(n720) );
  XOR U2474 ( .A(n719), .B(n720), .Z(n1484) );
  XNOR U2475 ( .A(x[641]), .B(y[641]), .Z(n1563) );
  XNOR U2476 ( .A(x[639]), .B(y[639]), .Z(n1561) );
  XNOR U2477 ( .A(x[715]), .B(y[715]), .Z(n1560) );
  XOR U2478 ( .A(n1561), .B(n1560), .Z(n1562) );
  XOR U2479 ( .A(n1563), .B(n1562), .Z(n1054) );
  XNOR U2480 ( .A(x[637]), .B(y[637]), .Z(n1567) );
  XNOR U2481 ( .A(x[635]), .B(y[635]), .Z(n1565) );
  XNOR U2482 ( .A(x[717]), .B(y[717]), .Z(n1564) );
  XOR U2483 ( .A(n1565), .B(n1564), .Z(n1566) );
  XOR U2484 ( .A(n1567), .B(n1566), .Z(n1051) );
  XNOR U2485 ( .A(x[92]), .B(y[92]), .Z(n936) );
  XNOR U2486 ( .A(x[94]), .B(y[94]), .Z(n934) );
  XNOR U2487 ( .A(x[96]), .B(y[96]), .Z(n933) );
  XNOR U2488 ( .A(n934), .B(n933), .Z(n935) );
  XOR U2489 ( .A(n936), .B(n935), .Z(n1052) );
  XNOR U2490 ( .A(n1051), .B(n1052), .Z(n1053) );
  XNOR U2491 ( .A(n1054), .B(n1053), .Z(n1485) );
  XNOR U2492 ( .A(n1484), .B(n1485), .Z(n1486) );
  XNOR U2493 ( .A(x[617]), .B(y[617]), .Z(n1549) );
  XNOR U2494 ( .A(x[615]), .B(y[615]), .Z(n1547) );
  XNOR U2495 ( .A(x[727]), .B(y[727]), .Z(n1546) );
  XOR U2496 ( .A(n1547), .B(n1546), .Z(n1548) );
  XOR U2497 ( .A(n1549), .B(n1548), .Z(n713) );
  XNOR U2498 ( .A(x[774]), .B(y[774]), .Z(n1385) );
  XNOR U2499 ( .A(x[380]), .B(y[380]), .Z(n1383) );
  XNOR U2500 ( .A(x[776]), .B(y[776]), .Z(n1382) );
  XOR U2501 ( .A(n1383), .B(n1382), .Z(n1384) );
  XOR U2502 ( .A(n1385), .B(n1384), .Z(n714) );
  XOR U2503 ( .A(n713), .B(n714), .Z(n715) );
  XNOR U2504 ( .A(x[613]), .B(y[613]), .Z(n1553) );
  XNOR U2505 ( .A(x[611]), .B(y[611]), .Z(n1551) );
  XNOR U2506 ( .A(x[729]), .B(y[729]), .Z(n1550) );
  XOR U2507 ( .A(n1551), .B(n1550), .Z(n1552) );
  XOR U2508 ( .A(n1553), .B(n1552), .Z(n716) );
  XNOR U2509 ( .A(n715), .B(n716), .Z(n2585) );
  XNOR U2510 ( .A(x[116]), .B(y[116]), .Z(n806) );
  XNOR U2511 ( .A(x[120]), .B(y[120]), .Z(n804) );
  XNOR U2512 ( .A(x[124]), .B(y[124]), .Z(n803) );
  XNOR U2513 ( .A(n804), .B(n803), .Z(n805) );
  XOR U2514 ( .A(n806), .B(n805), .Z(n807) );
  XNOR U2515 ( .A(x[603]), .B(y[603]), .Z(n1393) );
  XNOR U2516 ( .A(x[599]), .B(y[599]), .Z(n1391) );
  XNOR U2517 ( .A(x[601]), .B(y[601]), .Z(n1390) );
  XOR U2518 ( .A(n1391), .B(n1390), .Z(n1392) );
  XOR U2519 ( .A(n1393), .B(n1392), .Z(n808) );
  XNOR U2520 ( .A(n807), .B(n808), .Z(n809) );
  XNOR U2521 ( .A(x[609]), .B(y[609]), .Z(n1389) );
  XNOR U2522 ( .A(x[605]), .B(y[605]), .Z(n1387) );
  XNOR U2523 ( .A(x[607]), .B(y[607]), .Z(n1386) );
  XOR U2524 ( .A(n1387), .B(n1386), .Z(n1388) );
  XOR U2525 ( .A(n1389), .B(n1388), .Z(n810) );
  XNOR U2526 ( .A(n809), .B(n810), .Z(n2583) );
  XNOR U2527 ( .A(x[649]), .B(y[649]), .Z(n1091) );
  XNOR U2528 ( .A(x[647]), .B(y[647]), .Z(n1089) );
  XNOR U2529 ( .A(x[659]), .B(y[659]), .Z(n1088) );
  XOR U2530 ( .A(n1089), .B(n1088), .Z(n1090) );
  XNOR U2531 ( .A(n1091), .B(n1090), .Z(n2113) );
  XNOR U2532 ( .A(x[790]), .B(y[790]), .Z(n1647) );
  XNOR U2533 ( .A(x[394]), .B(y[394]), .Z(n1645) );
  XNOR U2534 ( .A(x[792]), .B(y[792]), .Z(n1644) );
  XOR U2535 ( .A(n1645), .B(n1644), .Z(n1646) );
  XNOR U2536 ( .A(n1647), .B(n1646), .Z(n2111) );
  XNOR U2537 ( .A(x[699]), .B(y[699]), .Z(n1087) );
  XNOR U2538 ( .A(x[661]), .B(y[661]), .Z(n1085) );
  XNOR U2539 ( .A(x[701]), .B(y[701]), .Z(n1084) );
  XOR U2540 ( .A(n1085), .B(n1084), .Z(n1086) );
  XNOR U2541 ( .A(n1087), .B(n1086), .Z(n2112) );
  XNOR U2542 ( .A(n2111), .B(n2112), .Z(n2114) );
  XNOR U2543 ( .A(n2113), .B(n2114), .Z(n2584) );
  XNOR U2544 ( .A(n2583), .B(n2584), .Z(n2586) );
  XNOR U2545 ( .A(n2585), .B(n2586), .Z(n1487) );
  XOR U2546 ( .A(n1486), .B(n1487), .Z(n2640) );
  XNOR U2547 ( .A(n2639), .B(n2640), .Z(n1754) );
  XNOR U2548 ( .A(x[449]), .B(y[449]), .Z(n742) );
  XNOR U2549 ( .A(x[441]), .B(y[441]), .Z(n740) );
  XNOR U2550 ( .A(x[445]), .B(y[445]), .Z(n739) );
  XNOR U2551 ( .A(n740), .B(n739), .Z(n741) );
  XOR U2552 ( .A(n742), .B(n741), .Z(n875) );
  XNOR U2553 ( .A(x[182]), .B(y[182]), .Z(n1235) );
  XNOR U2554 ( .A(x[111]), .B(y[111]), .Z(n1233) );
  XNOR U2555 ( .A(x[184]), .B(y[184]), .Z(n1232) );
  XOR U2556 ( .A(n1233), .B(n1232), .Z(n1234) );
  XOR U2557 ( .A(n1235), .B(n1234), .Z(n876) );
  XNOR U2558 ( .A(n875), .B(n876), .Z(n878) );
  XNOR U2559 ( .A(x[437]), .B(y[437]), .Z(n734) );
  XNOR U2560 ( .A(x[429]), .B(y[429]), .Z(n732) );
  XNOR U2561 ( .A(x[433]), .B(y[433]), .Z(n731) );
  XNOR U2562 ( .A(n732), .B(n731), .Z(n733) );
  XOR U2563 ( .A(n734), .B(n733), .Z(n877) );
  XOR U2564 ( .A(n878), .B(n877), .Z(n1784) );
  XNOR U2565 ( .A(x[461]), .B(y[461]), .Z(n798) );
  XNOR U2566 ( .A(x[453]), .B(y[453]), .Z(n796) );
  XNOR U2567 ( .A(x[457]), .B(y[457]), .Z(n795) );
  XOR U2568 ( .A(n796), .B(n795), .Z(n797) );
  XOR U2569 ( .A(n798), .B(n797), .Z(n898) );
  XNOR U2570 ( .A(x[750]), .B(y[750]), .Z(n1373) );
  XNOR U2571 ( .A(x[358]), .B(y[358]), .Z(n1371) );
  XNOR U2572 ( .A(x[752]), .B(y[752]), .Z(n1370) );
  XOR U2573 ( .A(n1371), .B(n1370), .Z(n1372) );
  XOR U2574 ( .A(n1373), .B(n1372), .Z(n895) );
  XNOR U2575 ( .A(x[473]), .B(y[473]), .Z(n856) );
  XNOR U2576 ( .A(x[465]), .B(y[465]), .Z(n854) );
  XNOR U2577 ( .A(x[469]), .B(y[469]), .Z(n853) );
  XNOR U2578 ( .A(n854), .B(n853), .Z(n855) );
  XOR U2579 ( .A(n856), .B(n855), .Z(n896) );
  XNOR U2580 ( .A(n895), .B(n896), .Z(n897) );
  XNOR U2581 ( .A(n898), .B(n897), .Z(n1785) );
  XOR U2582 ( .A(n1784), .B(n1785), .Z(n1786) );
  XNOR U2583 ( .A(x[413]), .B(y[413]), .Z(n942) );
  XNOR U2584 ( .A(x[405]), .B(y[405]), .Z(n940) );
  XNOR U2585 ( .A(x[409]), .B(y[409]), .Z(n939) );
  XNOR U2586 ( .A(n940), .B(n939), .Z(n941) );
  XOR U2587 ( .A(n942), .B(n941), .Z(n839) );
  XNOR U2588 ( .A(x[744]), .B(y[744]), .Z(n768) );
  XNOR U2589 ( .A(x[746]), .B(y[746]), .Z(n766) );
  XNOR U2590 ( .A(x[748]), .B(y[748]), .Z(n765) );
  XNOR U2591 ( .A(n766), .B(n765), .Z(n767) );
  XOR U2592 ( .A(n768), .B(n767), .Z(n837) );
  XNOR U2593 ( .A(x[425]), .B(y[425]), .Z(n956) );
  XNOR U2594 ( .A(x[417]), .B(y[417]), .Z(n954) );
  XNOR U2595 ( .A(x[421]), .B(y[421]), .Z(n953) );
  XOR U2596 ( .A(n954), .B(n953), .Z(n955) );
  XNOR U2597 ( .A(n956), .B(n955), .Z(n838) );
  XOR U2598 ( .A(n837), .B(n838), .Z(n840) );
  XOR U2599 ( .A(n839), .B(n840), .Z(n1787) );
  XNOR U2600 ( .A(n1786), .B(n1787), .Z(n2631) );
  XNOR U2601 ( .A(x[401]), .B(y[401]), .Z(n904) );
  XNOR U2602 ( .A(x[395]), .B(y[395]), .Z(n902) );
  XNOR U2603 ( .A(x[397]), .B(y[397]), .Z(n901) );
  XOR U2604 ( .A(n902), .B(n901), .Z(n903) );
  XOR U2605 ( .A(n904), .B(n903), .Z(n871) );
  XNOR U2606 ( .A(x[393]), .B(y[393]), .Z(n822) );
  XNOR U2607 ( .A(x[389]), .B(y[389]), .Z(n820) );
  XNOR U2608 ( .A(x[391]), .B(y[391]), .Z(n819) );
  XOR U2609 ( .A(n820), .B(n819), .Z(n821) );
  XOR U2610 ( .A(n822), .B(n821), .Z(n872) );
  XOR U2611 ( .A(n871), .B(n872), .Z(n873) );
  XNOR U2612 ( .A(x[387]), .B(y[387]), .Z(n884) );
  XNOR U2613 ( .A(x[383]), .B(y[383]), .Z(n882) );
  XNOR U2614 ( .A(x[385]), .B(y[385]), .Z(n881) );
  XOR U2615 ( .A(n882), .B(n881), .Z(n883) );
  XOR U2616 ( .A(n884), .B(n883), .Z(n874) );
  XOR U2617 ( .A(n873), .B(n874), .Z(n2649) );
  XNOR U2618 ( .A(x[381]), .B(y[381]), .Z(n868) );
  XNOR U2619 ( .A(x[377]), .B(y[377]), .Z(n866) );
  XNOR U2620 ( .A(x[379]), .B(y[379]), .Z(n865) );
  XNOR U2621 ( .A(n866), .B(n865), .Z(n867) );
  XNOR U2622 ( .A(n868), .B(n867), .Z(n1353) );
  XNOR U2623 ( .A(x[375]), .B(y[375]), .Z(n862) );
  XNOR U2624 ( .A(x[371]), .B(y[371]), .Z(n860) );
  XNOR U2625 ( .A(x[373]), .B(y[373]), .Z(n859) );
  XNOR U2626 ( .A(n860), .B(n859), .Z(n861) );
  XNOR U2627 ( .A(n862), .B(n861), .Z(n1352) );
  XOR U2628 ( .A(n1353), .B(n1352), .Z(n1354) );
  XNOR U2629 ( .A(x[369]), .B(y[369]), .Z(n988) );
  XNOR U2630 ( .A(x[365]), .B(y[365]), .Z(n986) );
  XNOR U2631 ( .A(x[367]), .B(y[367]), .Z(n985) );
  XNOR U2632 ( .A(n986), .B(n985), .Z(n987) );
  XNOR U2633 ( .A(n988), .B(n987), .Z(n1355) );
  XOR U2634 ( .A(n1354), .B(n1355), .Z(n2648) );
  XNOR U2635 ( .A(x[351]), .B(y[351]), .Z(n1038) );
  XNOR U2636 ( .A(x[347]), .B(y[347]), .Z(n1036) );
  XNOR U2637 ( .A(x[349]), .B(y[349]), .Z(n1035) );
  XNOR U2638 ( .A(n1036), .B(n1035), .Z(n1037) );
  XNOR U2639 ( .A(n1038), .B(n1037), .Z(n2090) );
  XNOR U2640 ( .A(x[357]), .B(y[357]), .Z(n994) );
  XNOR U2641 ( .A(x[353]), .B(y[353]), .Z(n992) );
  XNOR U2642 ( .A(x[355]), .B(y[355]), .Z(n991) );
  XNOR U2643 ( .A(n992), .B(n991), .Z(n993) );
  XNOR U2644 ( .A(n994), .B(n993), .Z(n2087) );
  XNOR U2645 ( .A(x[363]), .B(y[363]), .Z(n982) );
  XNOR U2646 ( .A(x[359]), .B(y[359]), .Z(n980) );
  XNOR U2647 ( .A(x[361]), .B(y[361]), .Z(n979) );
  XNOR U2648 ( .A(n980), .B(n979), .Z(n981) );
  XOR U2649 ( .A(n982), .B(n981), .Z(n2088) );
  XOR U2650 ( .A(n2087), .B(n2088), .Z(n2089) );
  XNOR U2651 ( .A(n2090), .B(n2089), .Z(n2647) );
  XNOR U2652 ( .A(n2648), .B(n2647), .Z(n2650) );
  XNOR U2653 ( .A(n2649), .B(n2650), .Z(n2632) );
  XOR U2654 ( .A(n2631), .B(n2632), .Z(n2633) );
  XNOR U2655 ( .A(x[309]), .B(y[309]), .Z(n1435) );
  XNOR U2656 ( .A(x[305]), .B(y[305]), .Z(n1433) );
  XNOR U2657 ( .A(x[307]), .B(y[307]), .Z(n1432) );
  XOR U2658 ( .A(n1433), .B(n1432), .Z(n1434) );
  XOR U2659 ( .A(n1435), .B(n1434), .Z(n2709) );
  XNOR U2660 ( .A(x[303]), .B(y[303]), .Z(n1445) );
  XNOR U2661 ( .A(x[299]), .B(y[299]), .Z(n1443) );
  XNOR U2662 ( .A(x[301]), .B(y[301]), .Z(n1442) );
  XOR U2663 ( .A(n1443), .B(n1442), .Z(n1444) );
  XOR U2664 ( .A(n1445), .B(n1444), .Z(n2710) );
  XOR U2665 ( .A(n2709), .B(n2710), .Z(n2711) );
  XNOR U2666 ( .A(x[297]), .B(y[297]), .Z(n1261) );
  XNOR U2667 ( .A(x[293]), .B(y[293]), .Z(n1259) );
  XNOR U2668 ( .A(x[295]), .B(y[295]), .Z(n1258) );
  XNOR U2669 ( .A(n1259), .B(n1258), .Z(n1260) );
  XNOR U2670 ( .A(n1261), .B(n1260), .Z(n2712) );
  XOR U2671 ( .A(n2711), .B(n2712), .Z(n2644) );
  XNOR U2672 ( .A(x[333]), .B(y[333]), .Z(n1018) );
  XNOR U2673 ( .A(x[329]), .B(y[329]), .Z(n1016) );
  XNOR U2674 ( .A(x[331]), .B(y[331]), .Z(n1015) );
  XNOR U2675 ( .A(n1016), .B(n1015), .Z(n1017) );
  XOR U2676 ( .A(n1018), .B(n1017), .Z(n2315) );
  XNOR U2677 ( .A(x[339]), .B(y[339]), .Z(n1044) );
  XNOR U2678 ( .A(x[335]), .B(y[335]), .Z(n1042) );
  XNOR U2679 ( .A(x[337]), .B(y[337]), .Z(n1041) );
  XNOR U2680 ( .A(n1042), .B(n1041), .Z(n1043) );
  XOR U2681 ( .A(n1044), .B(n1043), .Z(n2316) );
  XNOR U2682 ( .A(n2315), .B(n2316), .Z(n2318) );
  XNOR U2683 ( .A(x[345]), .B(y[345]), .Z(n1032) );
  XNOR U2684 ( .A(x[341]), .B(y[341]), .Z(n1030) );
  XNOR U2685 ( .A(x[343]), .B(y[343]), .Z(n1029) );
  XNOR U2686 ( .A(n1030), .B(n1029), .Z(n1031) );
  XNOR U2687 ( .A(n1032), .B(n1031), .Z(n2317) );
  XNOR U2688 ( .A(n2318), .B(n2317), .Z(n2641) );
  XNOR U2689 ( .A(x[315]), .B(y[315]), .Z(n1441) );
  XNOR U2690 ( .A(x[311]), .B(y[311]), .Z(n1439) );
  XNOR U2691 ( .A(x[313]), .B(y[313]), .Z(n1438) );
  XOR U2692 ( .A(n1439), .B(n1438), .Z(n1440) );
  XOR U2693 ( .A(n1441), .B(n1440), .Z(n2296) );
  XNOR U2694 ( .A(x[321]), .B(y[321]), .Z(n1022) );
  XNOR U2695 ( .A(x[317]), .B(y[317]), .Z(n1020) );
  XNOR U2696 ( .A(x[319]), .B(y[319]), .Z(n1019) );
  XNOR U2697 ( .A(n1020), .B(n1019), .Z(n1021) );
  XOR U2698 ( .A(n1022), .B(n1021), .Z(n2293) );
  XNOR U2699 ( .A(x[327]), .B(y[327]), .Z(n1012) );
  XNOR U2700 ( .A(x[323]), .B(y[323]), .Z(n1010) );
  XNOR U2701 ( .A(x[325]), .B(y[325]), .Z(n1009) );
  XNOR U2702 ( .A(n1010), .B(n1009), .Z(n1011) );
  XOR U2703 ( .A(n1012), .B(n1011), .Z(n2294) );
  XOR U2704 ( .A(n2293), .B(n2294), .Z(n2295) );
  XNOR U2705 ( .A(n2296), .B(n2295), .Z(n2642) );
  XNOR U2706 ( .A(n2641), .B(n2642), .Z(n2643) );
  XOR U2707 ( .A(n2644), .B(n2643), .Z(n2634) );
  XOR U2708 ( .A(n2633), .B(n2634), .Z(n1752) );
  XNOR U2709 ( .A(x[549]), .B(y[549]), .Z(n1125) );
  XNOR U2710 ( .A(x[545]), .B(y[545]), .Z(n1123) );
  XNOR U2711 ( .A(x[547]), .B(y[547]), .Z(n1122) );
  XOR U2712 ( .A(n1123), .B(n1122), .Z(n1124) );
  XOR U2713 ( .A(n1125), .B(n1124), .Z(n949) );
  XNOR U2714 ( .A(x[758]), .B(y[758]), .Z(n1361) );
  XNOR U2715 ( .A(x[760]), .B(y[760]), .Z(n1359) );
  XNOR U2716 ( .A(x[762]), .B(y[762]), .Z(n1358) );
  XOR U2717 ( .A(n1359), .B(n1358), .Z(n1360) );
  XOR U2718 ( .A(n1361), .B(n1360), .Z(n950) );
  XOR U2719 ( .A(n949), .B(n950), .Z(n951) );
  XNOR U2720 ( .A(x[543]), .B(y[543]), .Z(n1129) );
  XNOR U2721 ( .A(x[539]), .B(y[539]), .Z(n1127) );
  XNOR U2722 ( .A(x[541]), .B(y[541]), .Z(n1126) );
  XOR U2723 ( .A(n1127), .B(n1126), .Z(n1128) );
  XOR U2724 ( .A(n1129), .B(n1128), .Z(n952) );
  XOR U2725 ( .A(n951), .B(n952), .Z(n1765) );
  XNOR U2726 ( .A(x[687]), .B(y[687]), .Z(n1069) );
  XNOR U2727 ( .A(x[683]), .B(y[683]), .Z(n1067) );
  XNOR U2728 ( .A(x[685]), .B(y[685]), .Z(n1066) );
  XNOR U2729 ( .A(n1067), .B(n1066), .Z(n1068) );
  XNOR U2730 ( .A(n1069), .B(n1068), .Z(n1203) );
  XNOR U2731 ( .A(x[48]), .B(y[48]), .Z(n2454) );
  XNOR U2732 ( .A(x[52]), .B(y[52]), .Z(n2452) );
  XNOR U2733 ( .A(x[399]), .B(y[399]), .Z(n2451) );
  XNOR U2734 ( .A(n2452), .B(n2451), .Z(n2453) );
  XNOR U2735 ( .A(n2454), .B(n2453), .Z(n1202) );
  XOR U2736 ( .A(n1203), .B(n1202), .Z(n1204) );
  XNOR U2737 ( .A(x[681]), .B(y[681]), .Z(n1075) );
  XNOR U2738 ( .A(x[675]), .B(y[675]), .Z(n1073) );
  XNOR U2739 ( .A(x[689]), .B(y[689]), .Z(n1072) );
  XNOR U2740 ( .A(n1073), .B(n1072), .Z(n1074) );
  XNOR U2741 ( .A(n1075), .B(n1074), .Z(n1205) );
  XOR U2742 ( .A(n1204), .B(n1205), .Z(n1762) );
  XNOR U2743 ( .A(x[537]), .B(y[537]), .Z(n1365) );
  XNOR U2744 ( .A(x[533]), .B(y[533]), .Z(n1363) );
  XNOR U2745 ( .A(x[535]), .B(y[535]), .Z(n1362) );
  XOR U2746 ( .A(n1363), .B(n1362), .Z(n1364) );
  XNOR U2747 ( .A(n1365), .B(n1364), .Z(n943) );
  XNOR U2748 ( .A(x[156]), .B(y[156]), .Z(n778) );
  XNOR U2749 ( .A(x[129]), .B(y[129]), .Z(n776) );
  XNOR U2750 ( .A(x[160]), .B(y[160]), .Z(n775) );
  XNOR U2751 ( .A(n776), .B(n775), .Z(n777) );
  XOR U2752 ( .A(n778), .B(n777), .Z(n944) );
  XNOR U2753 ( .A(n943), .B(n944), .Z(n945) );
  XNOR U2754 ( .A(x[531]), .B(y[531]), .Z(n1369) );
  XNOR U2755 ( .A(x[525]), .B(y[525]), .Z(n1367) );
  XNOR U2756 ( .A(x[529]), .B(y[529]), .Z(n1366) );
  XOR U2757 ( .A(n1367), .B(n1366), .Z(n1368) );
  XOR U2758 ( .A(n1369), .B(n1368), .Z(n946) );
  XOR U2759 ( .A(n945), .B(n946), .Z(n1763) );
  XNOR U2760 ( .A(n1762), .B(n1763), .Z(n1764) );
  XNOR U2761 ( .A(n1765), .B(n1764), .Z(n1493) );
  XNOR U2762 ( .A(x[707]), .B(y[707]), .Z(n1689) );
  XNOR U2763 ( .A(x[671]), .B(y[671]), .Z(n1687) );
  XNOR U2764 ( .A(x[709]), .B(y[709]), .Z(n1686) );
  XOR U2765 ( .A(n1687), .B(n1686), .Z(n1688) );
  XOR U2766 ( .A(n1689), .B(n1688), .Z(n787) );
  XNOR U2767 ( .A(x[784]), .B(y[784]), .Z(n1571) );
  XNOR U2768 ( .A(x[786]), .B(y[786]), .Z(n1569) );
  XNOR U2769 ( .A(x[788]), .B(y[788]), .Z(n1568) );
  XOR U2770 ( .A(n1569), .B(n1568), .Z(n1570) );
  XOR U2771 ( .A(n1571), .B(n1570), .Z(n788) );
  XOR U2772 ( .A(n787), .B(n788), .Z(n789) );
  XNOR U2773 ( .A(x[711]), .B(y[711]), .Z(n1695) );
  XNOR U2774 ( .A(x[653]), .B(y[653]), .Z(n1693) );
  XNOR U2775 ( .A(x[713]), .B(y[713]), .Z(n1692) );
  XOR U2776 ( .A(n1693), .B(n1692), .Z(n1694) );
  XOR U2777 ( .A(n1695), .B(n1694), .Z(n790) );
  XNOR U2778 ( .A(n789), .B(n790), .Z(n2597) );
  XNOR U2779 ( .A(x[703]), .B(y[703]), .Z(n1651) );
  XNOR U2780 ( .A(x[645]), .B(y[645]), .Z(n1649) );
  XNOR U2781 ( .A(x[663]), .B(y[663]), .Z(n1648) );
  XOR U2782 ( .A(n1649), .B(n1648), .Z(n1650) );
  XOR U2783 ( .A(n1651), .B(n1650), .Z(n783) );
  XNOR U2784 ( .A(x[78]), .B(y[78]), .Z(n892) );
  XNOR U2785 ( .A(x[80]), .B(y[80]), .Z(n890) );
  XNOR U2786 ( .A(x[183]), .B(y[183]), .Z(n889) );
  XOR U2787 ( .A(n890), .B(n889), .Z(n891) );
  XOR U2788 ( .A(n892), .B(n891), .Z(n782) );
  XNOR U2789 ( .A(x[643]), .B(y[643]), .Z(n1657) );
  XNOR U2790 ( .A(x[665]), .B(y[665]), .Z(n1655) );
  XNOR U2791 ( .A(x[705]), .B(y[705]), .Z(n1654) );
  XOR U2792 ( .A(n1655), .B(n1654), .Z(n1656) );
  XOR U2793 ( .A(n1657), .B(n1656), .Z(n781) );
  XOR U2794 ( .A(n782), .B(n781), .Z(n784) );
  XNOR U2795 ( .A(n783), .B(n784), .Z(n2595) );
  XNOR U2796 ( .A(x[625]), .B(y[625]), .Z(n1671) );
  XNOR U2797 ( .A(x[623]), .B(y[623]), .Z(n1669) );
  XNOR U2798 ( .A(x[723]), .B(y[723]), .Z(n1668) );
  XNOR U2799 ( .A(n1669), .B(n1668), .Z(n1670) );
  XNOR U2800 ( .A(n1671), .B(n1670), .Z(n1253) );
  XNOR U2801 ( .A(x[106]), .B(y[106]), .Z(n728) );
  XNOR U2802 ( .A(x[108]), .B(y[108]), .Z(n726) );
  XNOR U2803 ( .A(x[165]), .B(y[165]), .Z(n725) );
  XNOR U2804 ( .A(n726), .B(n725), .Z(n727) );
  XOR U2805 ( .A(n728), .B(n727), .Z(n1252) );
  XNOR U2806 ( .A(n1253), .B(n1252), .Z(n1254) );
  XNOR U2807 ( .A(x[621]), .B(y[621]), .Z(n1677) );
  XNOR U2808 ( .A(x[619]), .B(y[619]), .Z(n1675) );
  XNOR U2809 ( .A(x[725]), .B(y[725]), .Z(n1674) );
  XNOR U2810 ( .A(n1675), .B(n1674), .Z(n1676) );
  XOR U2811 ( .A(n1677), .B(n1676), .Z(n1255) );
  XNOR U2812 ( .A(n1254), .B(n1255), .Z(n2596) );
  XOR U2813 ( .A(n2595), .B(n2596), .Z(n2598) );
  XNOR U2814 ( .A(n2597), .B(n2598), .Z(n1490) );
  XNOR U2815 ( .A(x[585]), .B(y[585]), .Z(n1611) );
  XNOR U2816 ( .A(x[581]), .B(y[581]), .Z(n1609) );
  XNOR U2817 ( .A(x[583]), .B(y[583]), .Z(n1608) );
  XOR U2818 ( .A(n1609), .B(n1608), .Z(n1610) );
  XNOR U2819 ( .A(n1611), .B(n1610), .Z(n755) );
  XNOR U2820 ( .A(x[130]), .B(y[130]), .Z(n772) );
  XNOR U2821 ( .A(x[132]), .B(y[132]), .Z(n770) );
  XNOR U2822 ( .A(x[147]), .B(y[147]), .Z(n769) );
  XNOR U2823 ( .A(n770), .B(n769), .Z(n771) );
  XOR U2824 ( .A(n772), .B(n771), .Z(n756) );
  XNOR U2825 ( .A(n755), .B(n756), .Z(n757) );
  XNOR U2826 ( .A(x[579]), .B(y[579]), .Z(n1615) );
  XNOR U2827 ( .A(x[575]), .B(y[575]), .Z(n1613) );
  XNOR U2828 ( .A(x[577]), .B(y[577]), .Z(n1612) );
  XOR U2829 ( .A(n1613), .B(n1612), .Z(n1614) );
  XOR U2830 ( .A(n1615), .B(n1614), .Z(n758) );
  XNOR U2831 ( .A(n757), .B(n758), .Z(n2580) );
  XNOR U2832 ( .A(x[651]), .B(y[651]), .Z(n1643) );
  XNOR U2833 ( .A(x[655]), .B(y[655]), .Z(n1641) );
  XNOR U2834 ( .A(x[697]), .B(y[697]), .Z(n1640) );
  XOR U2835 ( .A(n1641), .B(n1640), .Z(n1642) );
  XOR U2836 ( .A(n1643), .B(n1642), .Z(n2108) );
  XNOR U2837 ( .A(x[66]), .B(y[66]), .Z(n2042) );
  XNOR U2838 ( .A(x[70]), .B(y[70]), .Z(n2040) );
  XNOR U2839 ( .A(x[72]), .B(y[72]), .Z(n2039) );
  XOR U2840 ( .A(n2040), .B(n2039), .Z(n2041) );
  XOR U2841 ( .A(n2042), .B(n2041), .Z(n2105) );
  XNOR U2842 ( .A(x[693]), .B(y[693]), .Z(n1639) );
  XNOR U2843 ( .A(x[657]), .B(y[657]), .Z(n1637) );
  XNOR U2844 ( .A(x[695]), .B(y[695]), .Z(n1636) );
  XOR U2845 ( .A(n1637), .B(n1636), .Z(n1638) );
  XNOR U2846 ( .A(n1639), .B(n1638), .Z(n2106) );
  XNOR U2847 ( .A(n2105), .B(n2106), .Z(n2107) );
  XNOR U2848 ( .A(n2108), .B(n2107), .Z(n2578) );
  XNOR U2849 ( .A(x[591]), .B(y[591]), .Z(n1597) );
  XNOR U2850 ( .A(x[587]), .B(y[587]), .Z(n1595) );
  XNOR U2851 ( .A(x[589]), .B(y[589]), .Z(n1594) );
  XOR U2852 ( .A(n1595), .B(n1594), .Z(n1596) );
  XOR U2853 ( .A(n1597), .B(n1596), .Z(n816) );
  XNOR U2854 ( .A(x[770]), .B(y[770]), .Z(n1607) );
  XNOR U2855 ( .A(x[376]), .B(y[376]), .Z(n1605) );
  XNOR U2856 ( .A(x[772]), .B(y[772]), .Z(n1604) );
  XOR U2857 ( .A(n1605), .B(n1604), .Z(n1606) );
  XOR U2858 ( .A(n1607), .B(n1606), .Z(n813) );
  XNOR U2859 ( .A(x[597]), .B(y[597]), .Z(n1593) );
  XNOR U2860 ( .A(x[593]), .B(y[593]), .Z(n1591) );
  XNOR U2861 ( .A(x[595]), .B(y[595]), .Z(n1590) );
  XOR U2862 ( .A(n1591), .B(n1590), .Z(n1592) );
  XNOR U2863 ( .A(n1593), .B(n1592), .Z(n814) );
  XNOR U2864 ( .A(n813), .B(n814), .Z(n815) );
  XOR U2865 ( .A(n816), .B(n815), .Z(n2577) );
  XNOR U2866 ( .A(n2578), .B(n2577), .Z(n2579) );
  XNOR U2867 ( .A(n2580), .B(n2579), .Z(n1491) );
  XNOR U2868 ( .A(n1490), .B(n1491), .Z(n1492) );
  XOR U2869 ( .A(n1493), .B(n1492), .Z(n1753) );
  XOR U2870 ( .A(n1752), .B(n1753), .Z(n1755) );
  XOR U2871 ( .A(n1754), .B(n1755), .Z(n1813) );
  XOR U2872 ( .A(n1812), .B(n1813), .Z(n1814) );
  XNOR U2873 ( .A(x[458]), .B(y[458]), .Z(n2664) );
  XNOR U2874 ( .A(x[460]), .B(y[460]), .Z(n2662) );
  XNOR U2875 ( .A(x[462]), .B(y[462]), .Z(n2661) );
  XNOR U2876 ( .A(n2662), .B(n2661), .Z(n2663) );
  XOR U2877 ( .A(n2664), .B(n2663), .Z(n1460) );
  XNOR U2878 ( .A(x[724]), .B(y[724]), .Z(n2672) );
  XNOR U2879 ( .A(x[726]), .B(y[726]), .Z(n2670) );
  XNOR U2880 ( .A(x[728]), .B(y[728]), .Z(n2669) );
  XNOR U2881 ( .A(n2670), .B(n2669), .Z(n2671) );
  XOR U2882 ( .A(n2672), .B(n2671), .Z(n1461) );
  XOR U2883 ( .A(n1460), .B(n1461), .Z(n1462) );
  XNOR U2884 ( .A(x[464]), .B(y[464]), .Z(n2668) );
  XNOR U2885 ( .A(x[466]), .B(y[466]), .Z(n2666) );
  XNOR U2886 ( .A(x[468]), .B(y[468]), .Z(n2665) );
  XNOR U2887 ( .A(n2666), .B(n2665), .Z(n2667) );
  XOR U2888 ( .A(n2668), .B(n2667), .Z(n1463) );
  XOR U2889 ( .A(n1462), .B(n1463), .Z(n794) );
  XNOR U2890 ( .A(x[470]), .B(y[470]), .Z(n2694) );
  XNOR U2891 ( .A(x[100]), .B(y[100]), .Z(n2692) );
  XNOR U2892 ( .A(x[472]), .B(y[472]), .Z(n2691) );
  XNOR U2893 ( .A(n2692), .B(n2691), .Z(n2693) );
  XOR U2894 ( .A(n2694), .B(n2693), .Z(n1454) );
  XNOR U2895 ( .A(x[718]), .B(y[718]), .Z(n1934) );
  XNOR U2896 ( .A(x[720]), .B(y[720]), .Z(n1932) );
  XNOR U2897 ( .A(x[722]), .B(y[722]), .Z(n1931) );
  XOR U2898 ( .A(n1932), .B(n1931), .Z(n1933) );
  XOR U2899 ( .A(n1934), .B(n1933), .Z(n1455) );
  XNOR U2900 ( .A(n1454), .B(n1455), .Z(n1456) );
  XNOR U2901 ( .A(x[474]), .B(y[474]), .Z(n2698) );
  XNOR U2902 ( .A(x[104]), .B(y[104]), .Z(n2696) );
  XNOR U2903 ( .A(x[476]), .B(y[476]), .Z(n2695) );
  XNOR U2904 ( .A(n2696), .B(n2695), .Z(n2697) );
  XOR U2905 ( .A(n2698), .B(n2697), .Z(n1457) );
  XOR U2906 ( .A(n1456), .B(n1457), .Z(n791) );
  XNOR U2907 ( .A(x[484]), .B(y[484]), .Z(n2682) );
  XNOR U2908 ( .A(x[486]), .B(y[486]), .Z(n2680) );
  XNOR U2909 ( .A(x[488]), .B(y[488]), .Z(n2679) );
  XNOR U2910 ( .A(n2680), .B(n2679), .Z(n2681) );
  XNOR U2911 ( .A(n2682), .B(n2681), .Z(n1451) );
  XNOR U2912 ( .A(x[714]), .B(y[714]), .Z(n1966) );
  XNOR U2913 ( .A(x[326]), .B(y[326]), .Z(n1964) );
  XNOR U2914 ( .A(x[716]), .B(y[716]), .Z(n1963) );
  XOR U2915 ( .A(n1964), .B(n1963), .Z(n1965) );
  XOR U2916 ( .A(n1966), .B(n1965), .Z(n1448) );
  XNOR U2917 ( .A(x[478]), .B(y[478]), .Z(n2676) );
  XNOR U2918 ( .A(x[480]), .B(y[480]), .Z(n2674) );
  XNOR U2919 ( .A(x[482]), .B(y[482]), .Z(n2673) );
  XNOR U2920 ( .A(n2674), .B(n2673), .Z(n2675) );
  XOR U2921 ( .A(n2676), .B(n2675), .Z(n1449) );
  XNOR U2922 ( .A(n1448), .B(n1449), .Z(n1450) );
  XOR U2923 ( .A(n1451), .B(n1450), .Z(n792) );
  XNOR U2924 ( .A(n791), .B(n792), .Z(n793) );
  XOR U2925 ( .A(n794), .B(n793), .Z(n1060) );
  XNOR U2926 ( .A(x[430]), .B(y[430]), .Z(n1978) );
  XNOR U2927 ( .A(x[64]), .B(y[64]), .Z(n1976) );
  XNOR U2928 ( .A(x[432]), .B(y[432]), .Z(n1975) );
  XNOR U2929 ( .A(n1976), .B(n1975), .Z(n1977) );
  XOR U2930 ( .A(n1978), .B(n1977), .Z(n1478) );
  XNOR U2931 ( .A(x[738]), .B(y[738]), .Z(n1982) );
  XNOR U2932 ( .A(x[740]), .B(y[740]), .Z(n1980) );
  XNOR U2933 ( .A(x[742]), .B(y[742]), .Z(n1979) );
  XNOR U2934 ( .A(n1980), .B(n1979), .Z(n1981) );
  XOR U2935 ( .A(n1982), .B(n1981), .Z(n1479) );
  XOR U2936 ( .A(n1478), .B(n1479), .Z(n1480) );
  XNOR U2937 ( .A(x[434]), .B(y[434]), .Z(n1998) );
  XNOR U2938 ( .A(x[68]), .B(y[68]), .Z(n1996) );
  XNOR U2939 ( .A(x[436]), .B(y[436]), .Z(n1995) );
  XNOR U2940 ( .A(n1996), .B(n1995), .Z(n1997) );
  XOR U2941 ( .A(n1998), .B(n1997), .Z(n1481) );
  XOR U2942 ( .A(n1480), .B(n1481), .Z(n763) );
  XNOR U2943 ( .A(x[450]), .B(y[450]), .Z(n1986) );
  XNOR U2944 ( .A(x[82]), .B(y[82]), .Z(n1984) );
  XNOR U2945 ( .A(x[452]), .B(y[452]), .Z(n1983) );
  XNOR U2946 ( .A(n1984), .B(n1983), .Z(n1985) );
  XNOR U2947 ( .A(n1986), .B(n1985), .Z(n1723) );
  XNOR U2948 ( .A(x[730]), .B(y[730]), .Z(n2688) );
  XNOR U2949 ( .A(x[340]), .B(y[340]), .Z(n2686) );
  XNOR U2950 ( .A(x[732]), .B(y[732]), .Z(n2685) );
  XNOR U2951 ( .A(n2686), .B(n2685), .Z(n2687) );
  XNOR U2952 ( .A(n2688), .B(n2687), .Z(n1722) );
  XOR U2953 ( .A(n1723), .B(n1722), .Z(n1724) );
  XNOR U2954 ( .A(x[454]), .B(y[454]), .Z(n1992) );
  XNOR U2955 ( .A(x[86]), .B(y[86]), .Z(n1990) );
  XNOR U2956 ( .A(x[456]), .B(y[456]), .Z(n1989) );
  XNOR U2957 ( .A(n1990), .B(n1989), .Z(n1991) );
  XNOR U2958 ( .A(n1992), .B(n1991), .Z(n1725) );
  XOR U2959 ( .A(n1724), .B(n1725), .Z(n761) );
  XNOR U2960 ( .A(x[438]), .B(y[438]), .Z(n2006) );
  XNOR U2961 ( .A(x[440]), .B(y[440]), .Z(n2004) );
  XNOR U2962 ( .A(x[442]), .B(y[442]), .Z(n2003) );
  XNOR U2963 ( .A(n2004), .B(n2003), .Z(n2005) );
  XOR U2964 ( .A(n2006), .B(n2005), .Z(n1472) );
  XNOR U2965 ( .A(x[734]), .B(y[734]), .Z(n2660) );
  XNOR U2966 ( .A(x[344]), .B(y[344]), .Z(n2658) );
  XNOR U2967 ( .A(x[736]), .B(y[736]), .Z(n2657) );
  XNOR U2968 ( .A(n2658), .B(n2657), .Z(n2659) );
  XOR U2969 ( .A(n2660), .B(n2659), .Z(n1473) );
  XOR U2970 ( .A(n1472), .B(n1473), .Z(n1474) );
  XNOR U2971 ( .A(x[444]), .B(y[444]), .Z(n2002) );
  XNOR U2972 ( .A(x[446]), .B(y[446]), .Z(n2000) );
  XNOR U2973 ( .A(x[448]), .B(y[448]), .Z(n1999) );
  XNOR U2974 ( .A(n2000), .B(n1999), .Z(n2001) );
  XOR U2975 ( .A(n2002), .B(n2001), .Z(n1475) );
  XOR U2976 ( .A(n1474), .B(n1475), .Z(n762) );
  XNOR U2977 ( .A(n761), .B(n762), .Z(n764) );
  XOR U2978 ( .A(n763), .B(n764), .Z(n1057) );
  XNOR U2979 ( .A(x[392]), .B(y[392]), .Z(n1877) );
  XNOR U2980 ( .A(x[32]), .B(y[32]), .Z(n1875) );
  XNOR U2981 ( .A(x[396]), .B(y[396]), .Z(n1874) );
  XNOR U2982 ( .A(n1875), .B(n1874), .Z(n1876) );
  XOR U2983 ( .A(n1877), .B(n1876), .Z(n1023) );
  XNOR U2984 ( .A(x[388]), .B(y[388]), .Z(n1881) );
  XNOR U2985 ( .A(x[28]), .B(y[28]), .Z(n1879) );
  XNOR U2986 ( .A(x[390]), .B(y[390]), .Z(n1878) );
  XNOR U2987 ( .A(n1879), .B(n1878), .Z(n1880) );
  XOR U2988 ( .A(n1881), .B(n1880), .Z(n1024) );
  XOR U2989 ( .A(n1023), .B(n1024), .Z(n1025) );
  XNOR U2990 ( .A(x[382]), .B(y[382]), .Z(n1873) );
  XNOR U2991 ( .A(x[384]), .B(y[384]), .Z(n1871) );
  XNOR U2992 ( .A(x[386]), .B(y[386]), .Z(n1870) );
  XNOR U2993 ( .A(n1871), .B(n1870), .Z(n1872) );
  XOR U2994 ( .A(n1873), .B(n1872), .Z(n1026) );
  XOR U2995 ( .A(n1025), .B(n1026), .Z(n2349) );
  XNOR U2996 ( .A(x[398]), .B(y[398]), .Z(n1885) );
  XNOR U2997 ( .A(x[400]), .B(y[400]), .Z(n1883) );
  XNOR U2998 ( .A(x[402]), .B(y[402]), .Z(n1882) );
  XNOR U2999 ( .A(n1883), .B(n1882), .Z(n1884) );
  XOR U3000 ( .A(n1885), .B(n1884), .Z(n1003) );
  XNOR U3001 ( .A(x[410]), .B(y[410]), .Z(n1857) );
  XNOR U3002 ( .A(x[46]), .B(y[46]), .Z(n1855) );
  XNOR U3003 ( .A(x[412]), .B(y[412]), .Z(n1854) );
  XNOR U3004 ( .A(n1855), .B(n1854), .Z(n1856) );
  XOR U3005 ( .A(n1857), .B(n1856), .Z(n1004) );
  XOR U3006 ( .A(n1003), .B(n1004), .Z(n1005) );
  XNOR U3007 ( .A(x[404]), .B(y[404]), .Z(n1849) );
  XNOR U3008 ( .A(x[406]), .B(y[406]), .Z(n1847) );
  XNOR U3009 ( .A(x[408]), .B(y[408]), .Z(n1846) );
  XNOR U3010 ( .A(n1847), .B(n1846), .Z(n1848) );
  XOR U3011 ( .A(n1849), .B(n1848), .Z(n1006) );
  XOR U3012 ( .A(n1005), .B(n1006), .Z(n2347) );
  XNOR U3013 ( .A(x[418]), .B(y[418]), .Z(n1974) );
  XNOR U3014 ( .A(x[420]), .B(y[420]), .Z(n1972) );
  XNOR U3015 ( .A(x[422]), .B(y[422]), .Z(n1971) );
  XNOR U3016 ( .A(n1972), .B(n1971), .Z(n1973) );
  XOR U3017 ( .A(n1974), .B(n1973), .Z(n1104) );
  XNOR U3018 ( .A(x[414]), .B(y[414]), .Z(n1853) );
  XNOR U3019 ( .A(x[50]), .B(y[50]), .Z(n1851) );
  XNOR U3020 ( .A(x[416]), .B(y[416]), .Z(n1850) );
  XNOR U3021 ( .A(n1851), .B(n1850), .Z(n1852) );
  XOR U3022 ( .A(n1853), .B(n1852), .Z(n1105) );
  XOR U3023 ( .A(n1104), .B(n1105), .Z(n1106) );
  XNOR U3024 ( .A(x[424]), .B(y[424]), .Z(n1970) );
  XNOR U3025 ( .A(x[426]), .B(y[426]), .Z(n1968) );
  XNOR U3026 ( .A(x[428]), .B(y[428]), .Z(n1967) );
  XNOR U3027 ( .A(n1968), .B(n1967), .Z(n1969) );
  XOR U3028 ( .A(n1970), .B(n1969), .Z(n1107) );
  XOR U3029 ( .A(n1106), .B(n1107), .Z(n2348) );
  XOR U3030 ( .A(n2347), .B(n2348), .Z(n2350) );
  XOR U3031 ( .A(n2349), .B(n2350), .Z(n1058) );
  XNOR U3032 ( .A(n1057), .B(n1058), .Z(n1059) );
  XOR U3033 ( .A(n1060), .B(n1059), .Z(n2564) );
  XNOR U3034 ( .A(x[550]), .B(y[550]), .Z(n2210) );
  XNOR U3035 ( .A(x[172]), .B(y[172]), .Z(n2208) );
  XNOR U3036 ( .A(x[552]), .B(y[552]), .Z(n2207) );
  XNOR U3037 ( .A(n2208), .B(n2207), .Z(n2209) );
  XNOR U3038 ( .A(n2210), .B(n2209), .Z(n2196) );
  XNOR U3039 ( .A(x[678]), .B(y[678]), .Z(n2130) );
  XNOR U3040 ( .A(x[680]), .B(y[680]), .Z(n2128) );
  XNOR U3041 ( .A(x[682]), .B(y[682]), .Z(n2127) );
  XNOR U3042 ( .A(n2128), .B(n2127), .Z(n2129) );
  XNOR U3043 ( .A(n2130), .B(n2129), .Z(n2195) );
  XNOR U3044 ( .A(n2196), .B(n2195), .Z(n2198) );
  XNOR U3045 ( .A(x[554]), .B(y[554]), .Z(n2136) );
  XNOR U3046 ( .A(x[176]), .B(y[176]), .Z(n2134) );
  XNOR U3047 ( .A(x[556]), .B(y[556]), .Z(n2133) );
  XNOR U3048 ( .A(n2134), .B(n2133), .Z(n2135) );
  XNOR U3049 ( .A(n2136), .B(n2135), .Z(n2197) );
  XNOR U3050 ( .A(n2198), .B(n2197), .Z(n1721) );
  XNOR U3051 ( .A(x[574]), .B(y[574]), .Z(n2518) );
  XNOR U3052 ( .A(x[194]), .B(y[194]), .Z(n2516) );
  XNOR U3053 ( .A(x[576]), .B(y[576]), .Z(n2515) );
  XNOR U3054 ( .A(n2516), .B(n2515), .Z(n2517) );
  XNOR U3055 ( .A(n2518), .B(n2517), .Z(n2141) );
  XNOR U3056 ( .A(x[670]), .B(y[670]), .Z(n2234) );
  XNOR U3057 ( .A(x[286]), .B(y[286]), .Z(n2232) );
  XNOR U3058 ( .A(x[672]), .B(y[672]), .Z(n2231) );
  XNOR U3059 ( .A(n2232), .B(n2231), .Z(n2233) );
  XNOR U3060 ( .A(n2234), .B(n2233), .Z(n2139) );
  XNOR U3061 ( .A(x[570]), .B(y[570]), .Z(n2378) );
  XNOR U3062 ( .A(x[190]), .B(y[190]), .Z(n2376) );
  XNOR U3063 ( .A(x[572]), .B(y[572]), .Z(n2375) );
  XNOR U3064 ( .A(n2376), .B(n2375), .Z(n2377) );
  XOR U3065 ( .A(n2378), .B(n2377), .Z(n2140) );
  XOR U3066 ( .A(n2139), .B(n2140), .Z(n2142) );
  XOR U3067 ( .A(n2141), .B(n2142), .Z(n1719) );
  XNOR U3068 ( .A(x[564]), .B(y[564]), .Z(n2484) );
  XNOR U3069 ( .A(x[566]), .B(y[566]), .Z(n2482) );
  XNOR U3070 ( .A(x[568]), .B(y[568]), .Z(n2481) );
  XNOR U3071 ( .A(n2482), .B(n2481), .Z(n2483) );
  XNOR U3072 ( .A(n2484), .B(n2483), .Z(n1717) );
  XNOR U3073 ( .A(x[674]), .B(y[674]), .Z(n2222) );
  XNOR U3074 ( .A(x[290]), .B(y[290]), .Z(n2220) );
  XNOR U3075 ( .A(x[676]), .B(y[676]), .Z(n2219) );
  XNOR U3076 ( .A(n2220), .B(n2219), .Z(n2221) );
  XNOR U3077 ( .A(n2222), .B(n2221), .Z(n1714) );
  XNOR U3078 ( .A(x[558]), .B(y[558]), .Z(n2228) );
  XNOR U3079 ( .A(x[560]), .B(y[560]), .Z(n2226) );
  XNOR U3080 ( .A(x[562]), .B(y[562]), .Z(n2225) );
  XNOR U3081 ( .A(n2226), .B(n2225), .Z(n2227) );
  XOR U3082 ( .A(n2228), .B(n2227), .Z(n1715) );
  XOR U3083 ( .A(n1714), .B(n1715), .Z(n1716) );
  XNOR U3084 ( .A(n1717), .B(n1716), .Z(n1718) );
  XOR U3085 ( .A(n1719), .B(n1718), .Z(n1720) );
  XNOR U3086 ( .A(n1721), .B(n1720), .Z(n2561) );
  XNOR U3087 ( .A(x[590]), .B(y[590]), .Z(n2536) );
  XNOR U3088 ( .A(x[214]), .B(y[214]), .Z(n2534) );
  XNOR U3089 ( .A(x[592]), .B(y[592]), .Z(n2533) );
  XNOR U3090 ( .A(n2534), .B(n2533), .Z(n2535) );
  XNOR U3091 ( .A(n2536), .B(n2535), .Z(n2510) );
  XNOR U3092 ( .A(x[658]), .B(y[658]), .Z(n2500) );
  XNOR U3093 ( .A(x[660]), .B(y[660]), .Z(n2498) );
  XNOR U3094 ( .A(x[662]), .B(y[662]), .Z(n2497) );
  XNOR U3095 ( .A(n2498), .B(n2497), .Z(n2499) );
  XNOR U3096 ( .A(n2500), .B(n2499), .Z(n2509) );
  XNOR U3097 ( .A(n2510), .B(n2509), .Z(n2512) );
  XNOR U3098 ( .A(x[594]), .B(y[594]), .Z(n2506) );
  XNOR U3099 ( .A(x[218]), .B(y[218]), .Z(n2504) );
  XNOR U3100 ( .A(x[596]), .B(y[596]), .Z(n2503) );
  XNOR U3101 ( .A(n2504), .B(n2503), .Z(n2505) );
  XNOR U3102 ( .A(n2506), .B(n2505), .Z(n2511) );
  XNOR U3103 ( .A(n2512), .B(n2511), .Z(n1494) );
  XNOR U3104 ( .A(x[624]), .B(y[624]), .Z(n2546) );
  XNOR U3105 ( .A(x[626]), .B(y[626]), .Z(n2544) );
  XNOR U3106 ( .A(x[628]), .B(y[628]), .Z(n2543) );
  XNOR U3107 ( .A(n2544), .B(n2543), .Z(n2545) );
  XNOR U3108 ( .A(n2546), .B(n2545), .Z(n1113) );
  XNOR U3109 ( .A(x[638]), .B(y[638]), .Z(n2384) );
  XNOR U3110 ( .A(x[640]), .B(y[640]), .Z(n2382) );
  XNOR U3111 ( .A(x[642]), .B(y[642]), .Z(n2381) );
  XNOR U3112 ( .A(n2382), .B(n2381), .Z(n2383) );
  XNOR U3113 ( .A(n2384), .B(n2383), .Z(n1110) );
  XNOR U3114 ( .A(x[634]), .B(y[634]), .Z(n2390) );
  XNOR U3115 ( .A(x[254]), .B(y[254]), .Z(n2388) );
  XNOR U3116 ( .A(x[636]), .B(y[636]), .Z(n2387) );
  XNOR U3117 ( .A(n2388), .B(n2387), .Z(n2389) );
  XOR U3118 ( .A(n2390), .B(n2389), .Z(n1111) );
  XNOR U3119 ( .A(n1110), .B(n1111), .Z(n1112) );
  XNOR U3120 ( .A(n1113), .B(n1112), .Z(n1495) );
  XOR U3121 ( .A(n1494), .B(n1495), .Z(n1496) );
  XNOR U3122 ( .A(x[584]), .B(y[584]), .Z(n2478) );
  XNOR U3123 ( .A(x[586]), .B(y[586]), .Z(n2476) );
  XNOR U3124 ( .A(x[588]), .B(y[588]), .Z(n2475) );
  XNOR U3125 ( .A(n2476), .B(n2475), .Z(n2477) );
  XOR U3126 ( .A(n2478), .B(n2477), .Z(n2119) );
  XNOR U3127 ( .A(x[664]), .B(y[664]), .Z(n2494) );
  XNOR U3128 ( .A(x[666]), .B(y[666]), .Z(n2492) );
  XNOR U3129 ( .A(x[668]), .B(y[668]), .Z(n2491) );
  XNOR U3130 ( .A(n2492), .B(n2491), .Z(n2493) );
  XOR U3131 ( .A(n2494), .B(n2493), .Z(n2117) );
  XNOR U3132 ( .A(x[578]), .B(y[578]), .Z(n2356) );
  XNOR U3133 ( .A(x[580]), .B(y[580]), .Z(n2354) );
  XNOR U3134 ( .A(x[582]), .B(y[582]), .Z(n2353) );
  XNOR U3135 ( .A(n2354), .B(n2353), .Z(n2355) );
  XOR U3136 ( .A(n2356), .B(n2355), .Z(n2118) );
  XOR U3137 ( .A(n2117), .B(n2118), .Z(n2120) );
  XOR U3138 ( .A(n2119), .B(n2120), .Z(n1497) );
  XOR U3139 ( .A(n1496), .B(n1497), .Z(n2562) );
  XOR U3140 ( .A(n2561), .B(n2562), .Z(n2563) );
  XNOR U3141 ( .A(n2564), .B(n2563), .Z(n2728) );
  XNOR U3142 ( .A(x[197]), .B(y[197]), .Z(n2080) );
  XNOR U3143 ( .A(x[195]), .B(y[195]), .Z(n2078) );
  XNOR U3144 ( .A(x[495]), .B(y[495]), .Z(n2077) );
  XNOR U3145 ( .A(n2078), .B(n2077), .Z(n2079) );
  XOR U3146 ( .A(n2080), .B(n2079), .Z(n2243) );
  XNOR U3147 ( .A(x[193]), .B(y[193]), .Z(n2056) );
  XNOR U3148 ( .A(x[191]), .B(y[191]), .Z(n2054) );
  XNOR U3149 ( .A(x[749]), .B(y[749]), .Z(n2053) );
  XNOR U3150 ( .A(n2054), .B(n2053), .Z(n2055) );
  XOR U3151 ( .A(n2056), .B(n2055), .Z(n2244) );
  XOR U3152 ( .A(n2243), .B(n2244), .Z(n2245) );
  XNOR U3153 ( .A(x[189]), .B(y[189]), .Z(n2064) );
  XNOR U3154 ( .A(x[185]), .B(y[185]), .Z(n2062) );
  XNOR U3155 ( .A(x[491]), .B(y[491]), .Z(n2061) );
  XNOR U3156 ( .A(n2062), .B(n2061), .Z(n2063) );
  XOR U3157 ( .A(n2064), .B(n2063), .Z(n2246) );
  XOR U3158 ( .A(n2245), .B(n2246), .Z(n2653) );
  XNOR U3159 ( .A(x[207]), .B(y[207]), .Z(n2076) );
  XNOR U3160 ( .A(x[205]), .B(y[205]), .Z(n2074) );
  XNOR U3161 ( .A(x[499]), .B(y[499]), .Z(n2073) );
  XNOR U3162 ( .A(n2074), .B(n2073), .Z(n2075) );
  XOR U3163 ( .A(n2076), .B(n2075), .Z(n2237) );
  XNOR U3164 ( .A(x[211]), .B(y[211]), .Z(n1251) );
  XNOR U3165 ( .A(x[209]), .B(y[209]), .Z(n1249) );
  XNOR U3166 ( .A(x[745]), .B(y[745]), .Z(n1248) );
  XNOR U3167 ( .A(n1249), .B(n1248), .Z(n1250) );
  XOR U3168 ( .A(n1251), .B(n1250), .Z(n2238) );
  XOR U3169 ( .A(n2237), .B(n2238), .Z(n2239) );
  XNOR U3170 ( .A(x[203]), .B(y[203]), .Z(n2072) );
  XNOR U3171 ( .A(x[199]), .B(y[199]), .Z(n2070) );
  XNOR U3172 ( .A(x[747]), .B(y[747]), .Z(n2069) );
  XNOR U3173 ( .A(n2070), .B(n2069), .Z(n2071) );
  XOR U3174 ( .A(n2072), .B(n2071), .Z(n2240) );
  XOR U3175 ( .A(n2239), .B(n2240), .Z(n2654) );
  XOR U3176 ( .A(n2653), .B(n2654), .Z(n2655) );
  XNOR U3177 ( .A(x[173]), .B(y[173]), .Z(n2252) );
  XNOR U3178 ( .A(x[171]), .B(y[171]), .Z(n2250) );
  XNOR U3179 ( .A(x[753]), .B(y[753]), .Z(n2249) );
  XOR U3180 ( .A(n2250), .B(n2249), .Z(n2251) );
  XOR U3181 ( .A(n2252), .B(n2251), .Z(n2050) );
  XNOR U3182 ( .A(x[177]), .B(y[177]), .Z(n2262) );
  XNOR U3183 ( .A(x[175]), .B(y[175]), .Z(n2260) );
  XNOR U3184 ( .A(x[487]), .B(y[487]), .Z(n2259) );
  XOR U3185 ( .A(n2260), .B(n2259), .Z(n2261) );
  XOR U3186 ( .A(n2262), .B(n2261), .Z(n2047) );
  XNOR U3187 ( .A(x[181]), .B(y[181]), .Z(n2060) );
  XNOR U3188 ( .A(x[179]), .B(y[179]), .Z(n2058) );
  XNOR U3189 ( .A(x[751]), .B(y[751]), .Z(n2057) );
  XOR U3190 ( .A(n2058), .B(n2057), .Z(n2059) );
  XNOR U3191 ( .A(n2060), .B(n2059), .Z(n2048) );
  XNOR U3192 ( .A(n2047), .B(n2048), .Z(n2049) );
  XOR U3193 ( .A(n2050), .B(n2049), .Z(n2656) );
  XOR U3194 ( .A(n2655), .B(n2656), .Z(n2591) );
  XNOR U3195 ( .A(x[259]), .B(y[259]), .Z(n1193) );
  XNOR U3196 ( .A(x[257]), .B(y[257]), .Z(n1191) );
  XNOR U3197 ( .A(x[733]), .B(y[733]), .Z(n1190) );
  XOR U3198 ( .A(n1191), .B(n1190), .Z(n1192) );
  XOR U3199 ( .A(n1193), .B(n1192), .Z(n2705) );
  XNOR U3200 ( .A(x[255]), .B(y[255]), .Z(n1211) );
  XNOR U3201 ( .A(x[253]), .B(y[253]), .Z(n1209) );
  XNOR U3202 ( .A(x[523]), .B(y[523]), .Z(n1208) );
  XOR U3203 ( .A(n1209), .B(n1208), .Z(n1210) );
  XOR U3204 ( .A(n1211), .B(n1210), .Z(n2706) );
  XOR U3205 ( .A(n2705), .B(n2706), .Z(n2707) );
  XNOR U3206 ( .A(x[251]), .B(y[251]), .Z(n1223) );
  XNOR U3207 ( .A(x[249]), .B(y[249]), .Z(n1221) );
  XNOR U3208 ( .A(x[735]), .B(y[735]), .Z(n1220) );
  XOR U3209 ( .A(n1221), .B(n1220), .Z(n1222) );
  XOR U3210 ( .A(n1223), .B(n1222), .Z(n2708) );
  XNOR U3211 ( .A(n2707), .B(n2708), .Z(n1808) );
  XNOR U3212 ( .A(x[279]), .B(y[279]), .Z(n1305) );
  XNOR U3213 ( .A(x[275]), .B(y[275]), .Z(n1303) );
  XNOR U3214 ( .A(x[277]), .B(y[277]), .Z(n1302) );
  XNOR U3215 ( .A(n1303), .B(n1302), .Z(n1304) );
  XNOR U3216 ( .A(n1305), .B(n1304), .Z(n2610) );
  XNOR U3217 ( .A(x[285]), .B(y[285]), .Z(n1267) );
  XNOR U3218 ( .A(x[281]), .B(y[281]), .Z(n1265) );
  XNOR U3219 ( .A(x[283]), .B(y[283]), .Z(n1264) );
  XNOR U3220 ( .A(n1265), .B(n1264), .Z(n1266) );
  XNOR U3221 ( .A(n1267), .B(n1266), .Z(n2607) );
  XNOR U3222 ( .A(x[291]), .B(y[291]), .Z(n1273) );
  XNOR U3223 ( .A(x[287]), .B(y[287]), .Z(n1271) );
  XNOR U3224 ( .A(x[289]), .B(y[289]), .Z(n1270) );
  XNOR U3225 ( .A(n1271), .B(n1270), .Z(n1272) );
  XOR U3226 ( .A(n1273), .B(n1272), .Z(n2608) );
  XNOR U3227 ( .A(n2607), .B(n2608), .Z(n2609) );
  XOR U3228 ( .A(n2610), .B(n2609), .Z(n1807) );
  XNOR U3229 ( .A(x[273]), .B(y[273]), .Z(n1343) );
  XNOR U3230 ( .A(x[269]), .B(y[269]), .Z(n1341) );
  XNOR U3231 ( .A(x[271]), .B(y[271]), .Z(n1340) );
  XNOR U3232 ( .A(n1341), .B(n1340), .Z(n1342) );
  XNOR U3233 ( .A(n1343), .B(n1342), .Z(n2601) );
  XNOR U3234 ( .A(x[267]), .B(y[267]), .Z(n1199) );
  XNOR U3235 ( .A(x[265]), .B(y[265]), .Z(n1197) );
  XNOR U3236 ( .A(x[731]), .B(y[731]), .Z(n1196) );
  XOR U3237 ( .A(n1197), .B(n1196), .Z(n1198) );
  XOR U3238 ( .A(n1199), .B(n1198), .Z(n2602) );
  XOR U3239 ( .A(n2601), .B(n2602), .Z(n2603) );
  XNOR U3240 ( .A(x[263]), .B(y[263]), .Z(n1187) );
  XNOR U3241 ( .A(x[261]), .B(y[261]), .Z(n1185) );
  XNOR U3242 ( .A(x[527]), .B(y[527]), .Z(n1184) );
  XOR U3243 ( .A(n1185), .B(n1184), .Z(n1186) );
  XOR U3244 ( .A(n1187), .B(n1186), .Z(n2604) );
  XNOR U3245 ( .A(n2603), .B(n2604), .Z(n1806) );
  XOR U3246 ( .A(n1807), .B(n1806), .Z(n1809) );
  XOR U3247 ( .A(n1808), .B(n1809), .Z(n2590) );
  XNOR U3248 ( .A(x[239]), .B(y[239]), .Z(n1327) );
  XNOR U3249 ( .A(x[237]), .B(y[237]), .Z(n1325) );
  XNOR U3250 ( .A(x[515]), .B(y[515]), .Z(n1324) );
  XNOR U3251 ( .A(n1325), .B(n1324), .Z(n1326) );
  XNOR U3252 ( .A(n1327), .B(n1326), .Z(n2068) );
  XNOR U3253 ( .A(x[243]), .B(y[243]), .Z(n1317) );
  XNOR U3254 ( .A(x[241]), .B(y[241]), .Z(n1315) );
  XNOR U3255 ( .A(x[737]), .B(y[737]), .Z(n1314) );
  XNOR U3256 ( .A(n1315), .B(n1314), .Z(n1316) );
  XNOR U3257 ( .A(n1317), .B(n1316), .Z(n2065) );
  XNOR U3258 ( .A(x[247]), .B(y[247]), .Z(n1217) );
  XNOR U3259 ( .A(x[245]), .B(y[245]), .Z(n1215) );
  XNOR U3260 ( .A(x[519]), .B(y[519]), .Z(n1214) );
  XNOR U3261 ( .A(n1215), .B(n1214), .Z(n1216) );
  XOR U3262 ( .A(n1217), .B(n1216), .Z(n2066) );
  XOR U3263 ( .A(n2065), .B(n2066), .Z(n2067) );
  XNOR U3264 ( .A(n2068), .B(n2067), .Z(n1804) );
  XNOR U3265 ( .A(x[235]), .B(y[235]), .Z(n1323) );
  XNOR U3266 ( .A(x[233]), .B(y[233]), .Z(n1321) );
  XNOR U3267 ( .A(x[739]), .B(y[739]), .Z(n1320) );
  XNOR U3268 ( .A(n1321), .B(n1320), .Z(n1322) );
  XOR U3269 ( .A(n1323), .B(n1322), .Z(n2287) );
  XNOR U3270 ( .A(x[231]), .B(y[231]), .Z(n1171) );
  XNOR U3271 ( .A(x[229]), .B(y[229]), .Z(n1169) );
  XNOR U3272 ( .A(x[511]), .B(y[511]), .Z(n1168) );
  XNOR U3273 ( .A(n1169), .B(n1168), .Z(n1170) );
  XOR U3274 ( .A(n1171), .B(n1170), .Z(n2288) );
  XOR U3275 ( .A(n2287), .B(n2288), .Z(n2289) );
  XNOR U3276 ( .A(x[227]), .B(y[227]), .Z(n1167) );
  XNOR U3277 ( .A(x[225]), .B(y[225]), .Z(n1165) );
  XNOR U3278 ( .A(x[741]), .B(y[741]), .Z(n1164) );
  XNOR U3279 ( .A(n1165), .B(n1164), .Z(n1166) );
  XOR U3280 ( .A(n1167), .B(n1166), .Z(n2290) );
  XOR U3281 ( .A(n2289), .B(n2290), .Z(n1802) );
  XNOR U3282 ( .A(x[215]), .B(y[215]), .Z(n1243) );
  XNOR U3283 ( .A(x[213]), .B(y[213]), .Z(n1241) );
  XNOR U3284 ( .A(x[503]), .B(y[503]), .Z(n1240) );
  XOR U3285 ( .A(n1241), .B(n1240), .Z(n1242) );
  XOR U3286 ( .A(n1243), .B(n1242), .Z(n2266) );
  XNOR U3287 ( .A(x[219]), .B(y[219]), .Z(n1247) );
  XNOR U3288 ( .A(x[217]), .B(y[217]), .Z(n1245) );
  XNOR U3289 ( .A(x[743]), .B(y[743]), .Z(n1244) );
  XOR U3290 ( .A(n1245), .B(n1244), .Z(n1246) );
  XOR U3291 ( .A(n1247), .B(n1246), .Z(n2263) );
  XNOR U3292 ( .A(x[223]), .B(y[223]), .Z(n1175) );
  XNOR U3293 ( .A(x[221]), .B(y[221]), .Z(n1173) );
  XNOR U3294 ( .A(x[507]), .B(y[507]), .Z(n1172) );
  XNOR U3295 ( .A(n1173), .B(n1172), .Z(n1174) );
  XOR U3296 ( .A(n1175), .B(n1174), .Z(n2264) );
  XNOR U3297 ( .A(n2263), .B(n2264), .Z(n2265) );
  XNOR U3298 ( .A(n2266), .B(n2265), .Z(n1803) );
  XOR U3299 ( .A(n1802), .B(n1803), .Z(n1805) );
  XOR U3300 ( .A(n1804), .B(n1805), .Z(n2589) );
  XNOR U3301 ( .A(n2590), .B(n2589), .Z(n2592) );
  XOR U3302 ( .A(n2591), .B(n2592), .Z(n2725) );
  XNOR U3303 ( .A(x[196]), .B(y[196]), .Z(n2102) );
  XNOR U3304 ( .A(x[198]), .B(y[198]), .Z(n2100) );
  XNOR U3305 ( .A(x[206]), .B(y[206]), .Z(n2099) );
  XNOR U3306 ( .A(n2100), .B(n2099), .Z(n2101) );
  XNOR U3307 ( .A(n2102), .B(n2101), .Z(n2419) );
  XNOR U3308 ( .A(x[186]), .B(y[186]), .Z(n1229) );
  XNOR U3309 ( .A(x[188]), .B(y[188]), .Z(n1227) );
  XNOR U3310 ( .A(x[192]), .B(y[192]), .Z(n1226) );
  XOR U3311 ( .A(n1227), .B(n1226), .Z(n1228) );
  XNOR U3312 ( .A(n1229), .B(n1228), .Z(n2417) );
  XNOR U3313 ( .A(x[178]), .B(y[178]), .Z(n1239) );
  XNOR U3314 ( .A(x[115]), .B(y[115]), .Z(n1237) );
  XNOR U3315 ( .A(x[180]), .B(y[180]), .Z(n1236) );
  XOR U3316 ( .A(n1237), .B(n1236), .Z(n1238) );
  XNOR U3317 ( .A(n1239), .B(n1238), .Z(n2418) );
  XNOR U3318 ( .A(n2417), .B(n2418), .Z(n2420) );
  XOR U3319 ( .A(n2419), .B(n2420), .Z(n1926) );
  XNOR U3320 ( .A(x[162]), .B(y[162]), .Z(n1397) );
  XNOR U3321 ( .A(x[164]), .B(y[164]), .Z(n1395) );
  XNOR U3322 ( .A(x[166]), .B(y[166]), .Z(n1394) );
  XOR U3323 ( .A(n1395), .B(n1394), .Z(n1396) );
  XNOR U3324 ( .A(n1397), .B(n1396), .Z(n2395) );
  XNOR U3325 ( .A(x[150]), .B(y[150]), .Z(n1119) );
  XNOR U3326 ( .A(x[133]), .B(y[133]), .Z(n1117) );
  XNOR U3327 ( .A(x[152]), .B(y[152]), .Z(n1116) );
  XOR U3328 ( .A(n1117), .B(n1116), .Z(n1118) );
  XNOR U3329 ( .A(n1119), .B(n1118), .Z(n2393) );
  XNOR U3330 ( .A(x[134]), .B(y[134]), .Z(n1139) );
  XNOR U3331 ( .A(x[138]), .B(y[138]), .Z(n1137) );
  XNOR U3332 ( .A(x[142]), .B(y[142]), .Z(n1136) );
  XOR U3333 ( .A(n1137), .B(n1136), .Z(n1138) );
  XNOR U3334 ( .A(n1139), .B(n1138), .Z(n2394) );
  XNOR U3335 ( .A(n2393), .B(n2394), .Z(n2396) );
  XNOR U3336 ( .A(n2395), .B(n2396), .Z(n1925) );
  XOR U3337 ( .A(n1926), .B(n1925), .Z(n1927) );
  XNOR U3338 ( .A(x[126]), .B(y[126]), .Z(n1601) );
  XNOR U3339 ( .A(x[128]), .B(y[128]), .Z(n1599) );
  XNOR U3340 ( .A(x[151]), .B(y[151]), .Z(n1598) );
  XOR U3341 ( .A(n1599), .B(n1598), .Z(n1600) );
  XNOR U3342 ( .A(n1601), .B(n1600), .Z(n1842) );
  XNOR U3343 ( .A(x[110]), .B(y[110]), .Z(n1543) );
  XNOR U3344 ( .A(x[112]), .B(y[112]), .Z(n1541) );
  XNOR U3345 ( .A(x[114]), .B(y[114]), .Z(n1540) );
  XOR U3346 ( .A(n1541), .B(n1540), .Z(n1542) );
  XNOR U3347 ( .A(n1543), .B(n1542), .Z(n1840) );
  XNOR U3348 ( .A(x[98]), .B(y[98]), .Z(n1575) );
  XNOR U3349 ( .A(x[102]), .B(y[102]), .Z(n1573) );
  XNOR U3350 ( .A(x[169]), .B(y[169]), .Z(n1572) );
  XOR U3351 ( .A(n1573), .B(n1572), .Z(n1574) );
  XNOR U3352 ( .A(n1575), .B(n1574), .Z(n1841) );
  XNOR U3353 ( .A(n1840), .B(n1841), .Z(n1843) );
  XNOR U3354 ( .A(n1842), .B(n1843), .Z(n1928) );
  XNOR U3355 ( .A(n1927), .B(n1928), .Z(n2569) );
  XNOR U3356 ( .A(x[2]), .B(y[2]), .Z(n2192) );
  XNOR U3357 ( .A(x[4]), .B(y[4]), .Z(n2190) );
  XNOR U3358 ( .A(x[787]), .B(y[787]), .Z(n2189) );
  XNOR U3359 ( .A(n2190), .B(n2189), .Z(n2191) );
  XNOR U3360 ( .A(n2192), .B(n2191), .Z(n1625) );
  XNOR U3361 ( .A(x[6]), .B(y[6]), .Z(n2432) );
  XNOR U3362 ( .A(x[8]), .B(y[8]), .Z(n2430) );
  XNOR U3363 ( .A(x[415]), .B(y[415]), .Z(n2429) );
  XNOR U3364 ( .A(n2430), .B(n2429), .Z(n2431) );
  XOR U3365 ( .A(n2432), .B(n2431), .Z(n1624) );
  XNOR U3366 ( .A(n1625), .B(n1624), .Z(n1626) );
  XNOR U3367 ( .A(x[12]), .B(y[12]), .Z(n2426) );
  XNOR U3368 ( .A(x[16]), .B(y[16]), .Z(n2424) );
  XNOR U3369 ( .A(x[789]), .B(y[789]), .Z(n2423) );
  XNOR U3370 ( .A(n2424), .B(n2423), .Z(n2425) );
  XNOR U3371 ( .A(n2426), .B(n2425), .Z(n1627) );
  XOR U3372 ( .A(n1626), .B(n1627), .Z(n2625) );
  XNOR U3373 ( .A(x[13]), .B(y[13]), .Z(n2174) );
  XNOR U3374 ( .A(x[11]), .B(y[11]), .Z(n2172) );
  XNOR U3375 ( .A(x[423]), .B(y[423]), .Z(n2171) );
  XNOR U3376 ( .A(n2172), .B(n2171), .Z(n2173) );
  XNOR U3377 ( .A(n2174), .B(n2173), .Z(n1697) );
  XNOR U3378 ( .A(x[9]), .B(y[9]), .Z(n2186) );
  XNOR U3379 ( .A(x[5]), .B(y[5]), .Z(n2184) );
  XNOR U3380 ( .A(x[785]), .B(y[785]), .Z(n2183) );
  XNOR U3381 ( .A(n2184), .B(n2183), .Z(n2185) );
  XOR U3382 ( .A(n2186), .B(n2185), .Z(n1696) );
  XNOR U3383 ( .A(n1697), .B(n1696), .Z(n1698) );
  XNOR U3384 ( .A(x[1]), .B(y[1]), .Z(n2180) );
  XNOR U3385 ( .A(x[0]), .B(y[0]), .Z(n2178) );
  XNOR U3386 ( .A(x[419]), .B(y[419]), .Z(n2177) );
  XNOR U3387 ( .A(n2178), .B(n2177), .Z(n2179) );
  XNOR U3388 ( .A(n2180), .B(n2179), .Z(n1699) );
  XNOR U3389 ( .A(n1698), .B(n1699), .Z(n2626) );
  XNOR U3390 ( .A(n2625), .B(n2626), .Z(n2627) );
  XNOR U3391 ( .A(x[17]), .B(y[17]), .Z(n2162) );
  XNOR U3392 ( .A(x[15]), .B(y[15]), .Z(n2160) );
  XNOR U3393 ( .A(x[783]), .B(y[783]), .Z(n2159) );
  XOR U3394 ( .A(n2160), .B(n2159), .Z(n2161) );
  XNOR U3395 ( .A(n2162), .B(n2161), .Z(n1348) );
  XNOR U3396 ( .A(x[23]), .B(y[23]), .Z(n2168) );
  XNOR U3397 ( .A(x[19]), .B(y[19]), .Z(n2166) );
  XNOR U3398 ( .A(x[427]), .B(y[427]), .Z(n2165) );
  XOR U3399 ( .A(n2166), .B(n2165), .Z(n2167) );
  XNOR U3400 ( .A(n2168), .B(n2167), .Z(n1346) );
  XNOR U3401 ( .A(x[29]), .B(y[29]), .Z(n2158) );
  XNOR U3402 ( .A(x[27]), .B(y[27]), .Z(n2156) );
  XNOR U3403 ( .A(x[781]), .B(y[781]), .Z(n2155) );
  XOR U3404 ( .A(n2156), .B(n2155), .Z(n2157) );
  XNOR U3405 ( .A(n2158), .B(n2157), .Z(n1347) );
  XNOR U3406 ( .A(n1346), .B(n1347), .Z(n1349) );
  XNOR U3407 ( .A(n1348), .B(n1349), .Z(n2628) );
  XOR U3408 ( .A(n2627), .B(n2628), .Z(n2567) );
  XNOR U3409 ( .A(x[34]), .B(y[34]), .Z(n2468) );
  XNOR U3410 ( .A(x[36]), .B(y[36]), .Z(n2466) );
  XNOR U3411 ( .A(x[793]), .B(y[793]), .Z(n2465) );
  XOR U3412 ( .A(n2466), .B(n2465), .Z(n2467) );
  XOR U3413 ( .A(n2468), .B(n2467), .Z(n848) );
  XNOR U3414 ( .A(x[38]), .B(y[38]), .Z(n2450) );
  XNOR U3415 ( .A(x[40]), .B(y[40]), .Z(n2448) );
  XNOR U3416 ( .A(x[403]), .B(y[403]), .Z(n2447) );
  XOR U3417 ( .A(n2448), .B(n2447), .Z(n2449) );
  XNOR U3418 ( .A(n2450), .B(n2449), .Z(n847) );
  XNOR U3419 ( .A(n848), .B(n847), .Z(n850) );
  XNOR U3420 ( .A(x[42]), .B(y[42]), .Z(n2444) );
  XNOR U3421 ( .A(x[44]), .B(y[44]), .Z(n2442) );
  XNOR U3422 ( .A(x[795]), .B(y[795]), .Z(n2441) );
  XOR U3423 ( .A(n2442), .B(n2441), .Z(n2443) );
  XNOR U3424 ( .A(n2444), .B(n2443), .Z(n849) );
  XOR U3425 ( .A(n850), .B(n849), .Z(n2699) );
  XNOR U3426 ( .A(x[84]), .B(y[84]), .Z(n1683) );
  XNOR U3427 ( .A(x[88]), .B(y[88]), .Z(n1681) );
  XNOR U3428 ( .A(x[90]), .B(y[90]), .Z(n1680) );
  XOR U3429 ( .A(n1681), .B(n1680), .Z(n1682) );
  XNOR U3430 ( .A(n1683), .B(n1682), .Z(n843) );
  XNOR U3431 ( .A(x[74]), .B(y[74]), .Z(n1081) );
  XNOR U3432 ( .A(x[76]), .B(y[76]), .Z(n1079) );
  XNOR U3433 ( .A(x[187]), .B(y[187]), .Z(n1078) );
  XOR U3434 ( .A(n1079), .B(n1078), .Z(n1080) );
  XNOR U3435 ( .A(n1081), .B(n1080), .Z(n841) );
  XNOR U3436 ( .A(x[58]), .B(y[58]), .Z(n1505) );
  XNOR U3437 ( .A(x[60]), .B(y[60]), .Z(n1503) );
  XNOR U3438 ( .A(x[62]), .B(y[62]), .Z(n1502) );
  XOR U3439 ( .A(n1503), .B(n1502), .Z(n1504) );
  XNOR U3440 ( .A(n1505), .B(n1504), .Z(n842) );
  XNOR U3441 ( .A(n841), .B(n842), .Z(n844) );
  XNOR U3442 ( .A(n843), .B(n844), .Z(n2700) );
  XOR U3443 ( .A(n2699), .B(n2700), .Z(n2701) );
  XNOR U3444 ( .A(x[26]), .B(y[26]), .Z(n2460) );
  XNOR U3445 ( .A(x[30]), .B(y[30]), .Z(n2458) );
  XNOR U3446 ( .A(x[407]), .B(y[407]), .Z(n2457) );
  XNOR U3447 ( .A(n2458), .B(n2457), .Z(n2459) );
  XOR U3448 ( .A(n2460), .B(n2459), .Z(n1662) );
  XNOR U3449 ( .A(x[22]), .B(y[22]), .Z(n2464) );
  XNOR U3450 ( .A(x[24]), .B(y[24]), .Z(n2462) );
  XNOR U3451 ( .A(x[791]), .B(y[791]), .Z(n2461) );
  XNOR U3452 ( .A(n2462), .B(n2461), .Z(n2463) );
  XOR U3453 ( .A(n2464), .B(n2463), .Z(n1660) );
  XNOR U3454 ( .A(x[18]), .B(y[18]), .Z(n2438) );
  XNOR U3455 ( .A(x[20]), .B(y[20]), .Z(n2436) );
  XNOR U3456 ( .A(x[411]), .B(y[411]), .Z(n2435) );
  XNOR U3457 ( .A(n2436), .B(n2435), .Z(n2437) );
  XOR U3458 ( .A(n2438), .B(n2437), .Z(n1661) );
  XOR U3459 ( .A(n1660), .B(n1661), .Z(n1663) );
  XOR U3460 ( .A(n1662), .B(n1663), .Z(n2702) );
  XNOR U3461 ( .A(n2701), .B(n2702), .Z(n2568) );
  XNOR U3462 ( .A(n2567), .B(n2568), .Z(n2570) );
  XOR U3463 ( .A(n2569), .B(n2570), .Z(n2726) );
  XNOR U3464 ( .A(n2725), .B(n2726), .Z(n2727) );
  XOR U3465 ( .A(n2728), .B(n2727), .Z(n1815) );
  XOR U3466 ( .A(n1814), .B(n1815), .Z(o[0]) );
  NANDN U3467 ( .A(n708), .B(n707), .Z(n712) );
  NANDN U3468 ( .A(n710), .B(n709), .Z(n711) );
  NAND U3469 ( .A(n712), .B(n711), .Z(n3192) );
  OR U3470 ( .A(n726), .B(n725), .Z(n730) );
  OR U3471 ( .A(n728), .B(n727), .Z(n729) );
  NAND U3472 ( .A(n730), .B(n729), .Z(n3604) );
  XNOR U3473 ( .A(n3605), .B(n3604), .Z(n3607) );
  XOR U3474 ( .A(n3607), .B(n3606), .Z(n3484) );
  XNOR U3475 ( .A(n3483), .B(n3484), .Z(n3485) );
  XNOR U3476 ( .A(n3486), .B(n3485), .Z(n3697) );
  OR U3477 ( .A(n744), .B(n743), .Z(n748) );
  OR U3478 ( .A(n746), .B(n745), .Z(n747) );
  NAND U3479 ( .A(n748), .B(n747), .Z(n2931) );
  XNOR U3480 ( .A(n2932), .B(n2931), .Z(n2934) );
  OR U3481 ( .A(n750), .B(n749), .Z(n754) );
  OR U3482 ( .A(n752), .B(n751), .Z(n753) );
  NAND U3483 ( .A(n754), .B(n753), .Z(n2933) );
  XOR U3484 ( .A(n2934), .B(n2933), .Z(n3017) );
  NAND U3485 ( .A(n756), .B(n755), .Z(n760) );
  OR U3486 ( .A(n758), .B(n757), .Z(n759) );
  AND U3487 ( .A(n760), .B(n759), .Z(n3019) );
  XOR U3488 ( .A(n3017), .B(n3019), .Z(n3020) );
  XOR U3489 ( .A(n3021), .B(n3020), .Z(n3694) );
  XOR U3490 ( .A(n3694), .B(n3695), .Z(n3696) );
  XNOR U3491 ( .A(n3697), .B(n3696), .Z(n3190) );
  OR U3492 ( .A(n770), .B(n769), .Z(n774) );
  OR U3493 ( .A(n772), .B(n771), .Z(n773) );
  NAND U3494 ( .A(n774), .B(n773), .Z(n2995) );
  XOR U3495 ( .A(n2996), .B(n2995), .Z(n2997) );
  OR U3496 ( .A(n776), .B(n775), .Z(n780) );
  OR U3497 ( .A(n778), .B(n777), .Z(n779) );
  NAND U3498 ( .A(n780), .B(n779), .Z(n2998) );
  XNOR U3499 ( .A(n2997), .B(n2998), .Z(n3138) );
  NAND U3500 ( .A(n782), .B(n781), .Z(n786) );
  NAND U3501 ( .A(n784), .B(n783), .Z(n785) );
  AND U3502 ( .A(n786), .B(n785), .Z(n3136) );
  XNOR U3503 ( .A(n3136), .B(n3137), .Z(n3139) );
  XNOR U3504 ( .A(n3138), .B(n3139), .Z(n3716) );
  XOR U3505 ( .A(n3716), .B(n3717), .Z(n3718) );
  XNOR U3506 ( .A(n2982), .B(n2981), .Z(n2984) );
  XNOR U3507 ( .A(n2984), .B(n2983), .Z(n3450) );
  NANDN U3508 ( .A(n808), .B(n807), .Z(n812) );
  NANDN U3509 ( .A(n810), .B(n809), .Z(n811) );
  NAND U3510 ( .A(n812), .B(n811), .Z(n3447) );
  NANDN U3511 ( .A(n814), .B(n813), .Z(n818) );
  NAND U3512 ( .A(n816), .B(n815), .Z(n817) );
  NAND U3513 ( .A(n818), .B(n817), .Z(n3448) );
  XNOR U3514 ( .A(n3447), .B(n3448), .Z(n3449) );
  XOR U3515 ( .A(n3450), .B(n3449), .Z(n3719) );
  XOR U3516 ( .A(n3718), .B(n3719), .Z(n3189) );
  XOR U3517 ( .A(n3190), .B(n3189), .Z(n3191) );
  XOR U3518 ( .A(n3192), .B(n3191), .Z(n3174) );
  XNOR U3519 ( .A(n2762), .B(n2761), .Z(n2764) );
  XNOR U3520 ( .A(n2764), .B(n2763), .Z(n3465) );
  NANDN U3521 ( .A(n832), .B(n831), .Z(n836) );
  NAND U3522 ( .A(n834), .B(n833), .Z(n835) );
  NAND U3523 ( .A(n836), .B(n835), .Z(n3466) );
  XNOR U3524 ( .A(n3465), .B(n3466), .Z(n3467) );
  XNOR U3525 ( .A(n3467), .B(n3468), .Z(n3739) );
  OR U3526 ( .A(n842), .B(n841), .Z(n846) );
  OR U3527 ( .A(n844), .B(n843), .Z(n845) );
  NAND U3528 ( .A(n846), .B(n845), .Z(n3012) );
  NANDN U3529 ( .A(n848), .B(n847), .Z(n852) );
  NAND U3530 ( .A(n850), .B(n849), .Z(n851) );
  AND U3531 ( .A(n852), .B(n851), .Z(n3009) );
  OR U3532 ( .A(n854), .B(n853), .Z(n858) );
  OR U3533 ( .A(n856), .B(n855), .Z(n857) );
  NAND U3534 ( .A(n858), .B(n857), .Z(n3647) );
  OR U3535 ( .A(n860), .B(n859), .Z(n864) );
  OR U3536 ( .A(n862), .B(n861), .Z(n863) );
  AND U3537 ( .A(n864), .B(n863), .Z(n3646) );
  OR U3538 ( .A(n866), .B(n865), .Z(n870) );
  OR U3539 ( .A(n868), .B(n867), .Z(n869) );
  NAND U3540 ( .A(n870), .B(n869), .Z(n3649) );
  XNOR U3541 ( .A(n3648), .B(n3649), .Z(n3010) );
  XNOR U3542 ( .A(n3009), .B(n3010), .Z(n3011) );
  XOR U3543 ( .A(n3012), .B(n3011), .Z(n3736) );
  NANDN U3544 ( .A(n876), .B(n875), .Z(n880) );
  NAND U3545 ( .A(n878), .B(n877), .Z(n879) );
  NAND U3546 ( .A(n880), .B(n879), .Z(n3477) );
  OR U3547 ( .A(n890), .B(n889), .Z(n894) );
  NANDN U3548 ( .A(n892), .B(n891), .Z(n893) );
  AND U3549 ( .A(n894), .B(n893), .Z(n2798) );
  XNOR U3550 ( .A(n2797), .B(n2798), .Z(n2800) );
  XNOR U3551 ( .A(n2799), .B(n2800), .Z(n3478) );
  XNOR U3552 ( .A(n3477), .B(n3478), .Z(n3479) );
  XOR U3553 ( .A(n3480), .B(n3479), .Z(n3737) );
  XOR U3554 ( .A(n3736), .B(n3737), .Z(n3738) );
  XNOR U3555 ( .A(n3739), .B(n3738), .Z(n3193) );
  NANDN U3556 ( .A(n896), .B(n895), .Z(n900) );
  NAND U3557 ( .A(n898), .B(n897), .Z(n899) );
  NAND U3558 ( .A(n900), .B(n899), .Z(n3455) );
  OR U3559 ( .A(n906), .B(n905), .Z(n910) );
  OR U3560 ( .A(n908), .B(n907), .Z(n909) );
  NAND U3561 ( .A(n910), .B(n909), .Z(n2771) );
  XNOR U3562 ( .A(n2772), .B(n2771), .Z(n2774) );
  XNOR U3563 ( .A(n2774), .B(n2773), .Z(n3453) );
  NANDN U3564 ( .A(n916), .B(n915), .Z(n920) );
  NAND U3565 ( .A(n918), .B(n917), .Z(n919) );
  NAND U3566 ( .A(n920), .B(n919), .Z(n3454) );
  XOR U3567 ( .A(n3453), .B(n3454), .Z(n3456) );
  XOR U3568 ( .A(n3455), .B(n3456), .Z(n3698) );
  OR U3569 ( .A(n922), .B(n921), .Z(n926) );
  OR U3570 ( .A(n924), .B(n923), .Z(n925) );
  NAND U3571 ( .A(n926), .B(n925), .Z(n3491) );
  OR U3572 ( .A(n928), .B(n927), .Z(n932) );
  OR U3573 ( .A(n930), .B(n929), .Z(n931) );
  NAND U3574 ( .A(n932), .B(n931), .Z(n2804) );
  OR U3575 ( .A(n934), .B(n933), .Z(n938) );
  OR U3576 ( .A(n936), .B(n935), .Z(n937) );
  NAND U3577 ( .A(n938), .B(n937), .Z(n2803) );
  XNOR U3578 ( .A(n2804), .B(n2803), .Z(n2806) );
  XNOR U3579 ( .A(n2806), .B(n2805), .Z(n3489) );
  NAND U3580 ( .A(n944), .B(n943), .Z(n948) );
  OR U3581 ( .A(n946), .B(n945), .Z(n947) );
  AND U3582 ( .A(n948), .B(n947), .Z(n3490) );
  XOR U3583 ( .A(n3489), .B(n3490), .Z(n3492) );
  XOR U3584 ( .A(n3491), .B(n3492), .Z(n3699) );
  XOR U3585 ( .A(n3698), .B(n3699), .Z(n3700) );
  OR U3586 ( .A(n958), .B(n957), .Z(n962) );
  OR U3587 ( .A(n960), .B(n959), .Z(n961) );
  NAND U3588 ( .A(n962), .B(n961), .Z(n2809) );
  XNOR U3589 ( .A(n2810), .B(n2809), .Z(n2812) );
  OR U3590 ( .A(n964), .B(n963), .Z(n968) );
  OR U3591 ( .A(n966), .B(n965), .Z(n967) );
  NAND U3592 ( .A(n968), .B(n967), .Z(n2811) );
  XNOR U3593 ( .A(n2812), .B(n2811), .Z(n3459) );
  XNOR U3594 ( .A(n3459), .B(n3460), .Z(n3461) );
  XNOR U3595 ( .A(n3462), .B(n3461), .Z(n3701) );
  XNOR U3596 ( .A(n3700), .B(n3701), .Z(n3194) );
  XNOR U3597 ( .A(n3193), .B(n3194), .Z(n3196) );
  NANDN U3598 ( .A(n974), .B(n973), .Z(n978) );
  NAND U3599 ( .A(n976), .B(n975), .Z(n977) );
  AND U3600 ( .A(n978), .B(n977), .Z(n3016) );
  OR U3601 ( .A(n980), .B(n979), .Z(n984) );
  OR U3602 ( .A(n982), .B(n981), .Z(n983) );
  NAND U3603 ( .A(n984), .B(n983), .Z(n3641) );
  OR U3604 ( .A(n986), .B(n985), .Z(n990) );
  OR U3605 ( .A(n988), .B(n987), .Z(n989) );
  AND U3606 ( .A(n990), .B(n989), .Z(n3640) );
  XOR U3607 ( .A(n3641), .B(n3640), .Z(n3643) );
  OR U3608 ( .A(n992), .B(n991), .Z(n996) );
  OR U3609 ( .A(n994), .B(n993), .Z(n995) );
  NAND U3610 ( .A(n996), .B(n995), .Z(n3642) );
  XOR U3611 ( .A(n3643), .B(n3642), .Z(n3013) );
  NANDN U3612 ( .A(n998), .B(n997), .Z(n1002) );
  NAND U3613 ( .A(n1000), .B(n999), .Z(n1001) );
  AND U3614 ( .A(n1002), .B(n1001), .Z(n3014) );
  XNOR U3615 ( .A(n3013), .B(n3014), .Z(n3015) );
  XOR U3616 ( .A(n3016), .B(n3015), .Z(n3751) );
  NAND U3617 ( .A(n1004), .B(n1003), .Z(n1008) );
  NAND U3618 ( .A(n1006), .B(n1005), .Z(n1007) );
  NAND U3619 ( .A(n1008), .B(n1007), .Z(n3446) );
  OR U3620 ( .A(n1010), .B(n1009), .Z(n1014) );
  OR U3621 ( .A(n1012), .B(n1011), .Z(n1013) );
  NAND U3622 ( .A(n1014), .B(n1013), .Z(n2958) );
  XNOR U3623 ( .A(n2958), .B(n2957), .Z(n2960) );
  XNOR U3624 ( .A(n2960), .B(n2959), .Z(n3443) );
  NAND U3625 ( .A(n1024), .B(n1023), .Z(n1028) );
  NAND U3626 ( .A(n1026), .B(n1025), .Z(n1027) );
  AND U3627 ( .A(n1028), .B(n1027), .Z(n3444) );
  XOR U3628 ( .A(n3443), .B(n3444), .Z(n3445) );
  XOR U3629 ( .A(n3446), .B(n3445), .Z(n3748) );
  OR U3630 ( .A(n1030), .B(n1029), .Z(n1034) );
  OR U3631 ( .A(n1032), .B(n1031), .Z(n1033) );
  NAND U3632 ( .A(n1034), .B(n1033), .Z(n3631) );
  OR U3633 ( .A(n1036), .B(n1035), .Z(n1040) );
  OR U3634 ( .A(n1038), .B(n1037), .Z(n1039) );
  NAND U3635 ( .A(n1040), .B(n1039), .Z(n3630) );
  XOR U3636 ( .A(n3631), .B(n3630), .Z(n3632) );
  OR U3637 ( .A(n1042), .B(n1041), .Z(n1046) );
  OR U3638 ( .A(n1044), .B(n1043), .Z(n1045) );
  NAND U3639 ( .A(n1046), .B(n1045), .Z(n3633) );
  XNOR U3640 ( .A(n3632), .B(n3633), .Z(n3438) );
  XOR U3641 ( .A(n3438), .B(n3437), .Z(n3439) );
  NANDN U3642 ( .A(n1052), .B(n1051), .Z(n1056) );
  NAND U3643 ( .A(n1054), .B(n1053), .Z(n1055) );
  NAND U3644 ( .A(n1056), .B(n1055), .Z(n3440) );
  XNOR U3645 ( .A(n3439), .B(n3440), .Z(n3749) );
  XOR U3646 ( .A(n3748), .B(n3749), .Z(n3750) );
  XOR U3647 ( .A(n3751), .B(n3750), .Z(n3195) );
  XNOR U3648 ( .A(n3196), .B(n3195), .Z(n3171) );
  NAND U3649 ( .A(n1061), .B(oglobal[0]), .Z(n1065) );
  OR U3650 ( .A(n1063), .B(n1062), .Z(n1064) );
  NAND U3651 ( .A(n1065), .B(n1064), .Z(n3083) );
  OR U3652 ( .A(n1067), .B(n1066), .Z(n1071) );
  OR U3653 ( .A(n1069), .B(n1068), .Z(n1070) );
  NAND U3654 ( .A(n1071), .B(n1070), .Z(n3082) );
  XOR U3655 ( .A(n3083), .B(n3082), .Z(n3085) );
  OR U3656 ( .A(n1073), .B(n1072), .Z(n1077) );
  OR U3657 ( .A(n1075), .B(n1074), .Z(n1076) );
  NAND U3658 ( .A(n1077), .B(n1076), .Z(n3084) );
  XOR U3659 ( .A(n3085), .B(n3084), .Z(n3282) );
  OR U3660 ( .A(n1079), .B(n1078), .Z(n1083) );
  NANDN U3661 ( .A(n1081), .B(n1080), .Z(n1082) );
  NAND U3662 ( .A(n1083), .B(n1082), .Z(n3067) );
  XOR U3663 ( .A(n3067), .B(n3066), .Z(n3069) );
  XOR U3664 ( .A(n3069), .B(n3068), .Z(n3279) );
  NAND U3665 ( .A(n1093), .B(n1092), .Z(n1097) );
  NAND U3666 ( .A(n1095), .B(n1094), .Z(n1096) );
  AND U3667 ( .A(n1097), .B(n1096), .Z(n3280) );
  XNOR U3668 ( .A(n3279), .B(n3280), .Z(n3281) );
  XNOR U3669 ( .A(n3282), .B(n3281), .Z(n3170) );
  OR U3670 ( .A(n1099), .B(n1098), .Z(n1103) );
  NANDN U3671 ( .A(n1101), .B(n1100), .Z(n1102) );
  NAND U3672 ( .A(n1103), .B(n1102), .Z(n3392) );
  NAND U3673 ( .A(n1105), .B(n1104), .Z(n1109) );
  NAND U3674 ( .A(n1107), .B(n1106), .Z(n1108) );
  NAND U3675 ( .A(n1109), .B(n1108), .Z(n3389) );
  NANDN U3676 ( .A(n1111), .B(n1110), .Z(n1115) );
  NAND U3677 ( .A(n1113), .B(n1112), .Z(n1114) );
  NAND U3678 ( .A(n1115), .B(n1114), .Z(n3390) );
  XOR U3679 ( .A(n3389), .B(n3390), .Z(n3391) );
  XNOR U3680 ( .A(n3392), .B(n3391), .Z(n3168) );
  OR U3681 ( .A(n1117), .B(n1116), .Z(n1121) );
  NANDN U3682 ( .A(n1119), .B(n1118), .Z(n1120) );
  NAND U3683 ( .A(n1121), .B(n1120), .Z(n2828) );
  XNOR U3684 ( .A(n2828), .B(n2827), .Z(n2830) );
  XNOR U3685 ( .A(n2830), .B(n2829), .Z(n3288) );
  NAND U3686 ( .A(n1131), .B(n1130), .Z(n1135) );
  NAND U3687 ( .A(n1133), .B(n1132), .Z(n1134) );
  NAND U3688 ( .A(n1135), .B(n1134), .Z(n3285) );
  XNOR U3689 ( .A(n2896), .B(n2895), .Z(n2898) );
  XOR U3690 ( .A(n2898), .B(n2897), .Z(n3286) );
  XOR U3691 ( .A(n3285), .B(n3286), .Z(n3287) );
  XOR U3692 ( .A(n3288), .B(n3287), .Z(n3167) );
  XOR U3693 ( .A(n3168), .B(n3167), .Z(n3169) );
  XOR U3694 ( .A(n3170), .B(n3169), .Z(n2999) );
  XOR U3695 ( .A(n3000), .B(n2999), .Z(n3002) );
  XNOR U3696 ( .A(n3002), .B(n3001), .Z(n3172) );
  XOR U3697 ( .A(n3171), .B(n3172), .Z(n3173) );
  XOR U3698 ( .A(n3174), .B(n3173), .Z(n3797) );
  XNOR U3699 ( .A(n3659), .B(n3658), .Z(n3660) );
  XOR U3700 ( .A(n3660), .B(n3661), .Z(n3160) );
  XOR U3701 ( .A(n3107), .B(n3106), .Z(n3108) );
  OR U3702 ( .A(n1173), .B(n1172), .Z(n1177) );
  OR U3703 ( .A(n1175), .B(n1174), .Z(n1176) );
  NAND U3704 ( .A(n1177), .B(n1176), .Z(n3109) );
  XNOR U3705 ( .A(n3108), .B(n3109), .Z(n3156) );
  OR U3706 ( .A(n1179), .B(n1178), .Z(n1183) );
  OR U3707 ( .A(n1181), .B(n1180), .Z(n1182) );
  NAND U3708 ( .A(n1183), .B(n1182), .Z(n3158) );
  XOR U3709 ( .A(n3156), .B(n3158), .Z(n3159) );
  XOR U3710 ( .A(n3160), .B(n3159), .Z(n3007) );
  OR U3711 ( .A(n1185), .B(n1184), .Z(n1189) );
  NANDN U3712 ( .A(n1187), .B(n1186), .Z(n1188) );
  NAND U3713 ( .A(n1189), .B(n1188), .Z(n3035) );
  OR U3714 ( .A(n1191), .B(n1190), .Z(n1195) );
  NANDN U3715 ( .A(n1193), .B(n1192), .Z(n1194) );
  NAND U3716 ( .A(n1195), .B(n1194), .Z(n3034) );
  XOR U3717 ( .A(n3035), .B(n3034), .Z(n3036) );
  OR U3718 ( .A(n1197), .B(n1196), .Z(n1201) );
  NANDN U3719 ( .A(n1199), .B(n1198), .Z(n1200) );
  NAND U3720 ( .A(n1201), .B(n1200), .Z(n3037) );
  XNOR U3721 ( .A(n3036), .B(n3037), .Z(n3276) );
  OR U3722 ( .A(n1203), .B(n1202), .Z(n1207) );
  NANDN U3723 ( .A(n1205), .B(n1204), .Z(n1206) );
  NAND U3724 ( .A(n1207), .B(n1206), .Z(n3273) );
  OR U3725 ( .A(n1209), .B(n1208), .Z(n1213) );
  NANDN U3726 ( .A(n1211), .B(n1210), .Z(n1212) );
  NAND U3727 ( .A(n1213), .B(n1212), .Z(n3053) );
  OR U3728 ( .A(n1215), .B(n1214), .Z(n1219) );
  OR U3729 ( .A(n1217), .B(n1216), .Z(n1218) );
  NAND U3730 ( .A(n1219), .B(n1218), .Z(n3052) );
  XOR U3731 ( .A(n3053), .B(n3052), .Z(n3054) );
  OR U3732 ( .A(n1221), .B(n1220), .Z(n1225) );
  NANDN U3733 ( .A(n1223), .B(n1222), .Z(n1224) );
  NAND U3734 ( .A(n1225), .B(n1224), .Z(n3055) );
  XNOR U3735 ( .A(n3054), .B(n3055), .Z(n3274) );
  XNOR U3736 ( .A(n3273), .B(n3274), .Z(n3275) );
  XOR U3737 ( .A(n3276), .B(n3275), .Z(n3005) );
  OR U3738 ( .A(n1227), .B(n1226), .Z(n1231) );
  NANDN U3739 ( .A(n1229), .B(n1228), .Z(n1230) );
  NAND U3740 ( .A(n1231), .B(n1230), .Z(n3342) );
  XNOR U3741 ( .A(n3342), .B(n3341), .Z(n3344) );
  XNOR U3742 ( .A(n3344), .B(n3343), .Z(n3270) );
  XOR U3743 ( .A(n3623), .B(n3622), .Z(n3624) );
  XNOR U3744 ( .A(n3624), .B(n3625), .Z(n3268) );
  NANDN U3745 ( .A(n1253), .B(n1252), .Z(n1257) );
  NAND U3746 ( .A(n1255), .B(n1254), .Z(n1256) );
  AND U3747 ( .A(n1257), .B(n1256), .Z(n3267) );
  XOR U3748 ( .A(n3268), .B(n3267), .Z(n3269) );
  XOR U3749 ( .A(n3270), .B(n3269), .Z(n3006) );
  XNOR U3750 ( .A(n3005), .B(n3006), .Z(n3008) );
  XOR U3751 ( .A(n3007), .B(n3008), .Z(n3199) );
  OR U3752 ( .A(n1259), .B(n1258), .Z(n1263) );
  OR U3753 ( .A(n1261), .B(n1260), .Z(n1262) );
  NAND U3754 ( .A(n1263), .B(n1262), .Z(n2946) );
  OR U3755 ( .A(n1265), .B(n1264), .Z(n1269) );
  OR U3756 ( .A(n1267), .B(n1266), .Z(n1268) );
  NAND U3757 ( .A(n1269), .B(n1268), .Z(n2945) );
  XOR U3758 ( .A(n2946), .B(n2945), .Z(n2947) );
  OR U3759 ( .A(n1271), .B(n1270), .Z(n1275) );
  OR U3760 ( .A(n1273), .B(n1272), .Z(n1274) );
  NAND U3761 ( .A(n1275), .B(n1274), .Z(n2948) );
  XOR U3762 ( .A(n2947), .B(n2948), .Z(n3148) );
  NANDN U3763 ( .A(n1277), .B(n1276), .Z(n1281) );
  NAND U3764 ( .A(n1279), .B(n1278), .Z(n1280) );
  AND U3765 ( .A(n1281), .B(n1280), .Z(n3146) );
  NANDN U3766 ( .A(n1283), .B(n1282), .Z(n1287) );
  NAND U3767 ( .A(n1285), .B(n1284), .Z(n1286) );
  AND U3768 ( .A(n1287), .B(n1286), .Z(n3147) );
  XNOR U3769 ( .A(n3146), .B(n3147), .Z(n3149) );
  XOR U3770 ( .A(n3148), .B(n3149), .Z(n3773) );
  NANDN U3771 ( .A(n1289), .B(n1288), .Z(n1293) );
  NAND U3772 ( .A(n1291), .B(n1290), .Z(n1292) );
  NAND U3773 ( .A(n1293), .B(n1292), .Z(n3145) );
  XOR U3774 ( .A(n2950), .B(n2949), .Z(n2951) );
  OR U3775 ( .A(n1303), .B(n1302), .Z(n1307) );
  OR U3776 ( .A(n1305), .B(n1304), .Z(n1306) );
  NAND U3777 ( .A(n1307), .B(n1306), .Z(n2952) );
  XNOR U3778 ( .A(n2951), .B(n2952), .Z(n3142) );
  OR U3779 ( .A(n1309), .B(n1308), .Z(n1313) );
  OR U3780 ( .A(n1311), .B(n1310), .Z(n1312) );
  NAND U3781 ( .A(n1313), .B(n1312), .Z(n3143) );
  XOR U3782 ( .A(n3142), .B(n3143), .Z(n3144) );
  XNOR U3783 ( .A(n3145), .B(n3144), .Z(n3771) );
  OR U3784 ( .A(n1315), .B(n1314), .Z(n1319) );
  OR U3785 ( .A(n1317), .B(n1316), .Z(n1318) );
  NAND U3786 ( .A(n1319), .B(n1318), .Z(n3049) );
  XOR U3787 ( .A(n3049), .B(n3048), .Z(n3050) );
  OR U3788 ( .A(n1325), .B(n1324), .Z(n1329) );
  OR U3789 ( .A(n1327), .B(n1326), .Z(n1328) );
  NAND U3790 ( .A(n1329), .B(n1328), .Z(n3051) );
  XOR U3791 ( .A(n3050), .B(n3051), .Z(n3165) );
  OR U3792 ( .A(n1331), .B(n1330), .Z(n1335) );
  OR U3793 ( .A(n1333), .B(n1332), .Z(n1334) );
  NAND U3794 ( .A(n1335), .B(n1334), .Z(n3039) );
  XNOR U3795 ( .A(n3039), .B(n3038), .Z(n3041) );
  OR U3796 ( .A(n1341), .B(n1340), .Z(n1345) );
  OR U3797 ( .A(n1343), .B(n1342), .Z(n1344) );
  NAND U3798 ( .A(n1345), .B(n1344), .Z(n3040) );
  XOR U3799 ( .A(n3041), .B(n3040), .Z(n3163) );
  OR U3800 ( .A(n1347), .B(n1346), .Z(n1351) );
  OR U3801 ( .A(n1349), .B(n1348), .Z(n1350) );
  NAND U3802 ( .A(n1351), .B(n1350), .Z(n3164) );
  XOR U3803 ( .A(n3163), .B(n3164), .Z(n3166) );
  XOR U3804 ( .A(n3165), .B(n3166), .Z(n3770) );
  XOR U3805 ( .A(n3771), .B(n3770), .Z(n3772) );
  XOR U3806 ( .A(n3773), .B(n3772), .Z(n3200) );
  XOR U3807 ( .A(n3199), .B(n3200), .Z(n3202) );
  OR U3808 ( .A(n1353), .B(n1352), .Z(n1357) );
  NANDN U3809 ( .A(n1355), .B(n1354), .Z(n1356) );
  NAND U3810 ( .A(n1357), .B(n1356), .Z(n3244) );
  XNOR U3811 ( .A(n2864), .B(n2863), .Z(n2866) );
  XNOR U3812 ( .A(n2866), .B(n2865), .Z(n3243) );
  XOR U3813 ( .A(n3244), .B(n3243), .Z(n3245) );
  XNOR U3814 ( .A(n3366), .B(n3365), .Z(n3368) );
  XNOR U3815 ( .A(n3368), .B(n3367), .Z(n3246) );
  XOR U3816 ( .A(n3245), .B(n3246), .Z(n3497) );
  XNOR U3817 ( .A(n2870), .B(n2869), .Z(n2872) );
  XNOR U3818 ( .A(n2872), .B(n2871), .Z(n3230) );
  OR U3819 ( .A(n1395), .B(n1394), .Z(n1399) );
  NANDN U3820 ( .A(n1397), .B(n1396), .Z(n1398) );
  NAND U3821 ( .A(n1399), .B(n1398), .Z(n2858) );
  XNOR U3822 ( .A(n2858), .B(n2857), .Z(n2860) );
  XNOR U3823 ( .A(n2860), .B(n2859), .Z(n3227) );
  OR U3824 ( .A(n1409), .B(n1408), .Z(n1413) );
  NANDN U3825 ( .A(n1411), .B(n1410), .Z(n1412) );
  AND U3826 ( .A(n1413), .B(n1412), .Z(n3228) );
  XNOR U3827 ( .A(n3227), .B(n3228), .Z(n3229) );
  XOR U3828 ( .A(n3230), .B(n3229), .Z(n3495) );
  XNOR U3829 ( .A(n3348), .B(n3347), .Z(n3350) );
  XNOR U3830 ( .A(n3350), .B(n3349), .Z(n3258) );
  OR U3831 ( .A(n1427), .B(n1426), .Z(n1431) );
  NANDN U3832 ( .A(n1429), .B(n1428), .Z(n1430) );
  NAND U3833 ( .A(n1431), .B(n1430), .Z(n3255) );
  OR U3834 ( .A(n1433), .B(n1432), .Z(n1437) );
  NANDN U3835 ( .A(n1435), .B(n1434), .Z(n1436) );
  NAND U3836 ( .A(n1437), .B(n1436), .Z(n2954) );
  XOR U3837 ( .A(n2954), .B(n2953), .Z(n2956) );
  OR U3838 ( .A(n1443), .B(n1442), .Z(n1447) );
  NANDN U3839 ( .A(n1445), .B(n1444), .Z(n1446) );
  NAND U3840 ( .A(n1447), .B(n1446), .Z(n2955) );
  XOR U3841 ( .A(n2956), .B(n2955), .Z(n3256) );
  XOR U3842 ( .A(n3255), .B(n3256), .Z(n3257) );
  XOR U3843 ( .A(n3258), .B(n3257), .Z(n3496) );
  XOR U3844 ( .A(n3495), .B(n3496), .Z(n3498) );
  XNOR U3845 ( .A(n3497), .B(n3498), .Z(n3201) );
  XOR U3846 ( .A(n3202), .B(n3201), .Z(n3217) );
  NANDN U3847 ( .A(n1449), .B(n1448), .Z(n1453) );
  NAND U3848 ( .A(n1451), .B(n1450), .Z(n1452) );
  NAND U3849 ( .A(n1453), .B(n1452), .Z(n3422) );
  NANDN U3850 ( .A(n1455), .B(n1454), .Z(n1459) );
  NAND U3851 ( .A(n1457), .B(n1456), .Z(n1458) );
  NAND U3852 ( .A(n1459), .B(n1458), .Z(n3419) );
  NAND U3853 ( .A(n1461), .B(n1460), .Z(n1465) );
  NAND U3854 ( .A(n1463), .B(n1462), .Z(n1464) );
  AND U3855 ( .A(n1465), .B(n1464), .Z(n3420) );
  XNOR U3856 ( .A(n3419), .B(n3420), .Z(n3421) );
  XOR U3857 ( .A(n3422), .B(n3421), .Z(n3548) );
  NANDN U3858 ( .A(n1467), .B(n1466), .Z(n1471) );
  NAND U3859 ( .A(n1469), .B(n1468), .Z(n1470) );
  NAND U3860 ( .A(n1471), .B(n1470), .Z(n3402) );
  NAND U3861 ( .A(n1473), .B(n1472), .Z(n1477) );
  NAND U3862 ( .A(n1475), .B(n1474), .Z(n1476) );
  NAND U3863 ( .A(n1477), .B(n1476), .Z(n3399) );
  NAND U3864 ( .A(n1479), .B(n1478), .Z(n1483) );
  NAND U3865 ( .A(n1481), .B(n1480), .Z(n1482) );
  AND U3866 ( .A(n1483), .B(n1482), .Z(n3400) );
  XNOR U3867 ( .A(n3399), .B(n3400), .Z(n3401) );
  XOR U3868 ( .A(n3402), .B(n3401), .Z(n3549) );
  XOR U3869 ( .A(n3548), .B(n3549), .Z(n3550) );
  NANDN U3870 ( .A(n1485), .B(n1484), .Z(n1489) );
  NANDN U3871 ( .A(n1487), .B(n1486), .Z(n1488) );
  NAND U3872 ( .A(n1489), .B(n1488), .Z(n3551) );
  XOR U3873 ( .A(n3550), .B(n3551), .Z(n3184) );
  XOR U3874 ( .A(n3540), .B(n3539), .Z(n3542) );
  OR U3875 ( .A(n1511), .B(n1510), .Z(n1515) );
  NANDN U3876 ( .A(n1513), .B(n1512), .Z(n1514) );
  NAND U3877 ( .A(n1515), .B(n1514), .Z(n3541) );
  XOR U3878 ( .A(n3542), .B(n3541), .Z(n3385) );
  XNOR U3879 ( .A(n2840), .B(n2839), .Z(n2842) );
  XNOR U3880 ( .A(n2842), .B(n2841), .Z(n3384) );
  NANDN U3881 ( .A(n1529), .B(n1528), .Z(n1533) );
  NAND U3882 ( .A(n1531), .B(n1530), .Z(n1532) );
  AND U3883 ( .A(n1533), .B(n1532), .Z(n3383) );
  XOR U3884 ( .A(n3384), .B(n3383), .Z(n3386) );
  XOR U3885 ( .A(n3385), .B(n3386), .Z(n3500) );
  XNOR U3886 ( .A(n3499), .B(n3500), .Z(n3501) );
  XNOR U3887 ( .A(n3502), .B(n3501), .Z(n3182) );
  XNOR U3888 ( .A(n3181), .B(n3182), .Z(n3183) );
  XNOR U3889 ( .A(n3184), .B(n3183), .Z(n3215) );
  NANDN U3890 ( .A(n1535), .B(n1534), .Z(n1539) );
  NAND U3891 ( .A(n1537), .B(n1536), .Z(n1538) );
  AND U3892 ( .A(n1539), .B(n1538), .Z(n3027) );
  OR U3893 ( .A(n1541), .B(n1540), .Z(n1545) );
  NANDN U3894 ( .A(n1543), .B(n1542), .Z(n1544) );
  NAND U3895 ( .A(n1545), .B(n1544), .Z(n2882) );
  XNOR U3896 ( .A(n2882), .B(n2881), .Z(n2884) );
  XNOR U3897 ( .A(n2884), .B(n2883), .Z(n3314) );
  NAND U3898 ( .A(n1555), .B(n1554), .Z(n1559) );
  NANDN U3899 ( .A(n1557), .B(n1556), .Z(n1558) );
  NAND U3900 ( .A(n1559), .B(n1558), .Z(n3311) );
  XNOR U3901 ( .A(n3581), .B(n3580), .Z(n3583) );
  XOR U3902 ( .A(n3583), .B(n3582), .Z(n3312) );
  XNOR U3903 ( .A(n3311), .B(n3312), .Z(n3313) );
  XOR U3904 ( .A(n3314), .B(n3313), .Z(n3025) );
  XNOR U3905 ( .A(n2756), .B(n2755), .Z(n2758) );
  XNOR U3906 ( .A(n2758), .B(n2757), .Z(n3236) );
  OR U3907 ( .A(n1585), .B(n1584), .Z(n1589) );
  NANDN U3908 ( .A(n1587), .B(n1586), .Z(n1588) );
  NAND U3909 ( .A(n1589), .B(n1588), .Z(n3233) );
  XOR U3910 ( .A(n3559), .B(n3558), .Z(n3560) );
  OR U3911 ( .A(n1599), .B(n1598), .Z(n1603) );
  NANDN U3912 ( .A(n1601), .B(n1600), .Z(n1602) );
  NAND U3913 ( .A(n1603), .B(n1602), .Z(n3561) );
  XNOR U3914 ( .A(n3560), .B(n3561), .Z(n3234) );
  XNOR U3915 ( .A(n3233), .B(n3234), .Z(n3235) );
  XOR U3916 ( .A(n3236), .B(n3235), .Z(n3024) );
  XNOR U3917 ( .A(n3025), .B(n3024), .Z(n3026) );
  XOR U3918 ( .A(n3027), .B(n3026), .Z(n3185) );
  XNOR U3919 ( .A(n3563), .B(n3562), .Z(n3565) );
  XNOR U3920 ( .A(n3565), .B(n3564), .Z(n3296) );
  XOR U3921 ( .A(n3543), .B(oglobal[1]), .Z(n3545) );
  XNOR U3922 ( .A(n3544), .B(n3545), .Z(n3293) );
  NANDN U3923 ( .A(n1625), .B(n1624), .Z(n1629) );
  NANDN U3924 ( .A(n1627), .B(n1626), .Z(n1628) );
  NAND U3925 ( .A(n1629), .B(n1628), .Z(n3294) );
  XNOR U3926 ( .A(n3293), .B(n3294), .Z(n3295) );
  XOR U3927 ( .A(n3296), .B(n3295), .Z(n3431) );
  OR U3928 ( .A(n1631), .B(n1630), .Z(n1635) );
  NANDN U3929 ( .A(n1633), .B(n1632), .Z(n1634) );
  NAND U3930 ( .A(n1635), .B(n1634), .Z(n3087) );
  XNOR U3931 ( .A(n3087), .B(n3086), .Z(n3089) );
  XNOR U3932 ( .A(n3089), .B(n3088), .Z(n3302) );
  OR U3933 ( .A(n1649), .B(n1648), .Z(n1653) );
  NANDN U3934 ( .A(n1651), .B(n1650), .Z(n1652) );
  NAND U3935 ( .A(n1653), .B(n1652), .Z(n3574) );
  XNOR U3936 ( .A(n3575), .B(n3574), .Z(n3577) );
  OR U3937 ( .A(n1655), .B(n1654), .Z(n1659) );
  NANDN U3938 ( .A(n1657), .B(n1656), .Z(n1658) );
  NAND U3939 ( .A(n1659), .B(n1658), .Z(n3576) );
  XNOR U3940 ( .A(n3577), .B(n3576), .Z(n3299) );
  XNOR U3941 ( .A(n3299), .B(n3300), .Z(n3301) );
  XNOR U3942 ( .A(n3302), .B(n3301), .Z(n3432) );
  XNOR U3943 ( .A(n3431), .B(n3432), .Z(n3433) );
  OR U3944 ( .A(n1669), .B(n1668), .Z(n1673) );
  OR U3945 ( .A(n1671), .B(n1670), .Z(n1672) );
  NAND U3946 ( .A(n1673), .B(n1672), .Z(n2749) );
  XNOR U3947 ( .A(n2750), .B(n2749), .Z(n2752) );
  OR U3948 ( .A(n1675), .B(n1674), .Z(n1679) );
  OR U3949 ( .A(n1677), .B(n1676), .Z(n1678) );
  NAND U3950 ( .A(n1679), .B(n1678), .Z(n2751) );
  XNOR U3951 ( .A(n2752), .B(n2751), .Z(n3326) );
  OR U3952 ( .A(n1681), .B(n1680), .Z(n1685) );
  NANDN U3953 ( .A(n1683), .B(n1682), .Z(n1684) );
  NAND U3954 ( .A(n1685), .B(n1684), .Z(n3061) );
  OR U3955 ( .A(n1687), .B(n1686), .Z(n1691) );
  NANDN U3956 ( .A(n1689), .B(n1688), .Z(n1690) );
  NAND U3957 ( .A(n1691), .B(n1690), .Z(n3060) );
  XNOR U3958 ( .A(n3061), .B(n3060), .Z(n3063) );
  XNOR U3959 ( .A(n3063), .B(n3062), .Z(n3323) );
  NANDN U3960 ( .A(n1697), .B(n1696), .Z(n1701) );
  NANDN U3961 ( .A(n1699), .B(n1698), .Z(n1700) );
  AND U3962 ( .A(n1701), .B(n1700), .Z(n3324) );
  XNOR U3963 ( .A(n3323), .B(n3324), .Z(n3325) );
  XNOR U3964 ( .A(n3326), .B(n3325), .Z(n3434) );
  XNOR U3965 ( .A(n3433), .B(n3434), .Z(n3186) );
  XOR U3966 ( .A(n3185), .B(n3186), .Z(n3188) );
  NANDN U3967 ( .A(n1703), .B(n1702), .Z(n1707) );
  NAND U3968 ( .A(n1705), .B(n1704), .Z(n1706) );
  NAND U3969 ( .A(n1707), .B(n1706), .Z(n3413) );
  NAND U3970 ( .A(n1709), .B(n1708), .Z(n1713) );
  NAND U3971 ( .A(n1711), .B(n1710), .Z(n1712) );
  NAND U3972 ( .A(n1713), .B(n1712), .Z(n3412) );
  XOR U3973 ( .A(n3412), .B(n3411), .Z(n3414) );
  XOR U3974 ( .A(n3413), .B(n3414), .Z(n3329) );
  XNOR U3975 ( .A(n3329), .B(n3330), .Z(n3331) );
  OR U3976 ( .A(n1723), .B(n1722), .Z(n1727) );
  NANDN U3977 ( .A(n1725), .B(n1724), .Z(n1726) );
  NAND U3978 ( .A(n1727), .B(n1726), .Z(n3417) );
  NAND U3979 ( .A(n1729), .B(n1728), .Z(n1733) );
  NAND U3980 ( .A(n1731), .B(n1730), .Z(n1732) );
  AND U3981 ( .A(n1733), .B(n1732), .Z(n3415) );
  NAND U3982 ( .A(n1735), .B(n1734), .Z(n1739) );
  NANDN U3983 ( .A(n1737), .B(n1736), .Z(n1738) );
  AND U3984 ( .A(n1739), .B(n1738), .Z(n3416) );
  XOR U3985 ( .A(n3415), .B(n3416), .Z(n3418) );
  XOR U3986 ( .A(n3417), .B(n3418), .Z(n3101) );
  NAND U3987 ( .A(n1741), .B(n1740), .Z(n1745) );
  NAND U3988 ( .A(n1743), .B(n1742), .Z(n1744) );
  NAND U3989 ( .A(n1745), .B(n1744), .Z(n3099) );
  NAND U3990 ( .A(n1747), .B(n1746), .Z(n1751) );
  NAND U3991 ( .A(n1749), .B(n1748), .Z(n1750) );
  NAND U3992 ( .A(n1751), .B(n1750), .Z(n3098) );
  XOR U3993 ( .A(n3099), .B(n3098), .Z(n3100) );
  XOR U3994 ( .A(n3101), .B(n3100), .Z(n3332) );
  XNOR U3995 ( .A(n3331), .B(n3332), .Z(n3187) );
  XOR U3996 ( .A(n3188), .B(n3187), .Z(n3216) );
  XOR U3997 ( .A(n3215), .B(n3216), .Z(n3218) );
  XNOR U3998 ( .A(n3217), .B(n3218), .Z(n3794) );
  NAND U3999 ( .A(n1753), .B(n1752), .Z(n1757) );
  NAND U4000 ( .A(n1755), .B(n1754), .Z(n1756) );
  AND U4001 ( .A(n1757), .B(n1756), .Z(n3211) );
  NANDN U4002 ( .A(n1763), .B(n1762), .Z(n1767) );
  NAND U4003 ( .A(n1765), .B(n1764), .Z(n1766) );
  NAND U4004 ( .A(n1767), .B(n1766), .Z(n3767) );
  NANDN U4005 ( .A(n1769), .B(n1768), .Z(n1773) );
  NANDN U4006 ( .A(n1771), .B(n1770), .Z(n1772) );
  NAND U4007 ( .A(n1773), .B(n1772), .Z(n3765) );
  OR U4008 ( .A(n1775), .B(n1774), .Z(n1779) );
  NANDN U4009 ( .A(n1777), .B(n1776), .Z(n1778) );
  AND U4010 ( .A(n1779), .B(n1778), .Z(n3764) );
  XNOR U4011 ( .A(n3765), .B(n3764), .Z(n3766) );
  XNOR U4012 ( .A(n3767), .B(n3766), .Z(n2731) );
  XNOR U4013 ( .A(n2731), .B(n2732), .Z(n2734) );
  OR U4014 ( .A(n1785), .B(n1784), .Z(n1789) );
  NANDN U4015 ( .A(n1787), .B(n1786), .Z(n1788) );
  NAND U4016 ( .A(n1789), .B(n1788), .Z(n3508) );
  NANDN U4017 ( .A(n1791), .B(n1790), .Z(n1795) );
  NAND U4018 ( .A(n1793), .B(n1792), .Z(n1794) );
  NAND U4019 ( .A(n1795), .B(n1794), .Z(n3506) );
  OR U4020 ( .A(n1797), .B(n1796), .Z(n1801) );
  NANDN U4021 ( .A(n1799), .B(n1798), .Z(n1800) );
  NAND U4022 ( .A(n1801), .B(n1800), .Z(n3505) );
  XNOR U4023 ( .A(n3506), .B(n3505), .Z(n3507) );
  XNOR U4024 ( .A(n3508), .B(n3507), .Z(n3474) );
  NANDN U4025 ( .A(n1807), .B(n1806), .Z(n1811) );
  NANDN U4026 ( .A(n1809), .B(n1808), .Z(n1810) );
  NAND U4027 ( .A(n1811), .B(n1810), .Z(n3472) );
  XNOR U4028 ( .A(n3471), .B(n3472), .Z(n3473) );
  XOR U4029 ( .A(n3474), .B(n3473), .Z(n2733) );
  XNOR U4030 ( .A(n2734), .B(n2733), .Z(n3209) );
  XOR U4031 ( .A(n3210), .B(n3209), .Z(n3212) );
  XNOR U4032 ( .A(n3211), .B(n3212), .Z(n3795) );
  XNOR U4033 ( .A(n3794), .B(n3795), .Z(n3796) );
  XNOR U4034 ( .A(n3797), .B(n3796), .Z(n3221) );
  XNOR U4035 ( .A(n3221), .B(n3222), .Z(n3223) );
  NANDN U4036 ( .A(n1817), .B(n1816), .Z(n1821) );
  OR U4037 ( .A(n1819), .B(n1818), .Z(n1820) );
  NAND U4038 ( .A(n1821), .B(n1820), .Z(n3671) );
  OR U4039 ( .A(n1831), .B(n1830), .Z(n1835) );
  OR U4040 ( .A(n1833), .B(n1832), .Z(n1834) );
  NAND U4041 ( .A(n1835), .B(n1834), .Z(n3028) );
  XNOR U4042 ( .A(n3029), .B(n3028), .Z(n3031) );
  XNOR U4043 ( .A(n3031), .B(n3030), .Z(n3405) );
  OR U4044 ( .A(n1841), .B(n1840), .Z(n1845) );
  OR U4045 ( .A(n1843), .B(n1842), .Z(n1844) );
  NAND U4046 ( .A(n1845), .B(n1844), .Z(n3406) );
  XOR U4047 ( .A(n3405), .B(n3406), .Z(n3408) );
  XOR U4048 ( .A(n3407), .B(n3408), .Z(n3670) );
  XNOR U4049 ( .A(n3671), .B(n3670), .Z(n3672) );
  XOR U4050 ( .A(n2928), .B(n2927), .Z(n2929) );
  XNOR U4051 ( .A(n2929), .B(n2930), .Z(n3058) );
  OR U4052 ( .A(n1859), .B(n1858), .Z(n1863) );
  OR U4053 ( .A(n1861), .B(n1860), .Z(n1862) );
  NAND U4054 ( .A(n1863), .B(n1862), .Z(n2974) );
  OR U4055 ( .A(n1865), .B(n1864), .Z(n1869) );
  OR U4056 ( .A(n1867), .B(n1866), .Z(n1868) );
  NAND U4057 ( .A(n1869), .B(n1868), .Z(n2973) );
  XOR U4058 ( .A(n2974), .B(n2973), .Z(n2975) );
  XNOR U4059 ( .A(n2975), .B(n2976), .Z(n3056) );
  XOR U4060 ( .A(n2988), .B(n2987), .Z(n2989) );
  XNOR U4061 ( .A(n2989), .B(n2990), .Z(n3057) );
  XOR U4062 ( .A(n3056), .B(n3057), .Z(n3059) );
  XOR U4063 ( .A(n3058), .B(n3059), .Z(n3673) );
  XNOR U4064 ( .A(n3672), .B(n3673), .Z(n3689) );
  XOR U4065 ( .A(n2992), .B(n2991), .Z(n2994) );
  XOR U4066 ( .A(n2994), .B(n2993), .Z(n3380) );
  OR U4067 ( .A(n1903), .B(n1902), .Z(n1908) );
  IV U4068 ( .A(n1904), .Z(n1905) );
  NANDN U4069 ( .A(n1906), .B(n1905), .Z(n1907) );
  NAND U4070 ( .A(n1908), .B(n1907), .Z(n2887) );
  XOR U4071 ( .A(n2888), .B(n2887), .Z(n2890) );
  XOR U4072 ( .A(n2890), .B(n2889), .Z(n3378) );
  XOR U4073 ( .A(n2892), .B(n2891), .Z(n2894) );
  XOR U4074 ( .A(n2894), .B(n2893), .Z(n3377) );
  XNOR U4075 ( .A(n3378), .B(n3377), .Z(n3379) );
  XOR U4076 ( .A(n3380), .B(n3379), .Z(n3338) );
  OR U4077 ( .A(n1926), .B(n1925), .Z(n1930) );
  NANDN U4078 ( .A(n1928), .B(n1927), .Z(n1929) );
  NAND U4079 ( .A(n1930), .B(n1929), .Z(n3335) );
  XOR U4080 ( .A(n2916), .B(n2915), .Z(n2918) );
  XOR U4081 ( .A(n2918), .B(n2917), .Z(n2740) );
  XOR U4082 ( .A(n2978), .B(n2977), .Z(n2980) );
  XOR U4083 ( .A(n2980), .B(n2979), .Z(n2738) );
  XOR U4084 ( .A(n2924), .B(n2923), .Z(n2926) );
  XOR U4085 ( .A(n2926), .B(n2925), .Z(n2737) );
  XNOR U4086 ( .A(n2738), .B(n2737), .Z(n2739) );
  XOR U4087 ( .A(n2740), .B(n2739), .Z(n3336) );
  XNOR U4088 ( .A(n3335), .B(n3336), .Z(n3337) );
  XNOR U4089 ( .A(n3338), .B(n3337), .Z(n3688) );
  XOR U4090 ( .A(n3689), .B(n3688), .Z(n3691) );
  XOR U4091 ( .A(n2920), .B(n2919), .Z(n2921) );
  XNOR U4092 ( .A(n2921), .B(n2922), .Z(n3613) );
  OR U4093 ( .A(n1984), .B(n1983), .Z(n1988) );
  OR U4094 ( .A(n1986), .B(n1985), .Z(n1987) );
  NAND U4095 ( .A(n1988), .B(n1987), .Z(n3626) );
  XOR U4096 ( .A(n3627), .B(n3626), .Z(n3628) );
  OR U4097 ( .A(n1990), .B(n1989), .Z(n1994) );
  OR U4098 ( .A(n1992), .B(n1991), .Z(n1993) );
  NAND U4099 ( .A(n1994), .B(n1993), .Z(n3629) );
  XNOR U4100 ( .A(n3628), .B(n3629), .Z(n3611) );
  XNOR U4101 ( .A(n2816), .B(n2815), .Z(n2818) );
  XOR U4102 ( .A(n2818), .B(n2817), .Z(n3610) );
  XOR U4103 ( .A(n3611), .B(n3610), .Z(n3612) );
  XOR U4104 ( .A(n3613), .B(n3612), .Z(n3754) );
  XNOR U4105 ( .A(n3593), .B(n3592), .Z(n3594) );
  XOR U4106 ( .A(n3594), .B(n3595), .Z(n3664) );
  XNOR U4107 ( .A(n3372), .B(n3371), .Z(n3373) );
  XNOR U4108 ( .A(n3373), .B(n3374), .Z(n3665) );
  XNOR U4109 ( .A(n3664), .B(n3665), .Z(n3666) );
  XNOR U4110 ( .A(n3353), .B(n3354), .Z(n3355) );
  XNOR U4111 ( .A(n3356), .B(n3355), .Z(n3667) );
  XNOR U4112 ( .A(n3666), .B(n3667), .Z(n3752) );
  XNOR U4113 ( .A(n3752), .B(n3753), .Z(n3755) );
  XNOR U4114 ( .A(n3754), .B(n3755), .Z(n3690) );
  XNOR U4115 ( .A(n3691), .B(n3690), .Z(n3679) );
  NANDN U4116 ( .A(n2048), .B(n2047), .Z(n2052) );
  NAND U4117 ( .A(n2050), .B(n2049), .Z(n2051) );
  NAND U4118 ( .A(n2052), .B(n2051), .Z(n3252) );
  XOR U4119 ( .A(n3045), .B(n3044), .Z(n3046) );
  XNOR U4120 ( .A(n3046), .B(n3047), .Z(n3249) );
  XOR U4121 ( .A(n3249), .B(n3250), .Z(n3251) );
  XNOR U4122 ( .A(n3252), .B(n3251), .Z(n3725) );
  XOR U4123 ( .A(n3127), .B(n3126), .Z(n3128) );
  XNOR U4124 ( .A(n3128), .B(n3129), .Z(n3264) );
  OR U4125 ( .A(n2082), .B(n2081), .Z(n2086) );
  NANDN U4126 ( .A(n2084), .B(n2083), .Z(n2085) );
  NAND U4127 ( .A(n2086), .B(n2085), .Z(n3261) );
  XNOR U4128 ( .A(n3261), .B(n3262), .Z(n3263) );
  XOR U4129 ( .A(n3264), .B(n3263), .Z(n3722) );
  XNOR U4130 ( .A(n3360), .B(n3359), .Z(n3361) );
  OR U4131 ( .A(n2100), .B(n2099), .Z(n2104) );
  OR U4132 ( .A(n2102), .B(n2101), .Z(n2103) );
  AND U4133 ( .A(n2104), .B(n2103), .Z(n3362) );
  XNOR U4134 ( .A(n3361), .B(n3362), .Z(n3155) );
  NANDN U4135 ( .A(n2106), .B(n2105), .Z(n2110) );
  NAND U4136 ( .A(n2108), .B(n2107), .Z(n2109) );
  AND U4137 ( .A(n2110), .B(n2109), .Z(n3152) );
  OR U4138 ( .A(n2112), .B(n2111), .Z(n2116) );
  OR U4139 ( .A(n2114), .B(n2113), .Z(n2115) );
  AND U4140 ( .A(n2116), .B(n2115), .Z(n3153) );
  XNOR U4141 ( .A(n3152), .B(n3153), .Z(n3154) );
  XOR U4142 ( .A(n3155), .B(n3154), .Z(n3723) );
  XOR U4143 ( .A(n3722), .B(n3723), .Z(n3724) );
  XOR U4144 ( .A(n3725), .B(n3724), .Z(n3178) );
  OR U4145 ( .A(n2122), .B(n2121), .Z(n2126) );
  OR U4146 ( .A(n2124), .B(n2123), .Z(n2125) );
  NAND U4147 ( .A(n2126), .B(n2125), .Z(n2876) );
  OR U4148 ( .A(n2128), .B(n2127), .Z(n2132) );
  OR U4149 ( .A(n2130), .B(n2129), .Z(n2131) );
  NAND U4150 ( .A(n2132), .B(n2131), .Z(n2875) );
  XNOR U4151 ( .A(n2876), .B(n2875), .Z(n2878) );
  OR U4152 ( .A(n2134), .B(n2133), .Z(n2138) );
  OR U4153 ( .A(n2136), .B(n2135), .Z(n2137) );
  NAND U4154 ( .A(n2138), .B(n2137), .Z(n2877) );
  XOR U4155 ( .A(n2878), .B(n2877), .Z(n2901) );
  NANDN U4156 ( .A(n2140), .B(n2139), .Z(n2144) );
  NANDN U4157 ( .A(n2142), .B(n2141), .Z(n2143) );
  NAND U4158 ( .A(n2144), .B(n2143), .Z(n2902) );
  XOR U4159 ( .A(n2901), .B(n2902), .Z(n2903) );
  XNOR U4160 ( .A(n2904), .B(n2903), .Z(n3704) );
  OR U4161 ( .A(n2150), .B(n2149), .Z(n2154) );
  OR U4162 ( .A(n2152), .B(n2151), .Z(n2153) );
  AND U4163 ( .A(n2154), .B(n2153), .Z(n3652) );
  XNOR U4164 ( .A(n3654), .B(n3655), .Z(n2940) );
  OR U4165 ( .A(n2160), .B(n2159), .Z(n2164) );
  NANDN U4166 ( .A(n2162), .B(n2161), .Z(n2163) );
  NAND U4167 ( .A(n2164), .B(n2163), .Z(n2786) );
  OR U4168 ( .A(n2166), .B(n2165), .Z(n2170) );
  NANDN U4169 ( .A(n2168), .B(n2167), .Z(n2169) );
  NAND U4170 ( .A(n2170), .B(n2169), .Z(n2785) );
  XNOR U4171 ( .A(n2786), .B(n2785), .Z(n2788) );
  OR U4172 ( .A(n2172), .B(n2171), .Z(n2176) );
  OR U4173 ( .A(n2174), .B(n2173), .Z(n2175) );
  NAND U4174 ( .A(n2176), .B(n2175), .Z(n2787) );
  XOR U4175 ( .A(n2788), .B(n2787), .Z(n2937) );
  OR U4176 ( .A(n2178), .B(n2177), .Z(n2182) );
  OR U4177 ( .A(n2180), .B(n2179), .Z(n2181) );
  NAND U4178 ( .A(n2182), .B(n2181), .Z(n2834) );
  OR U4179 ( .A(n2184), .B(n2183), .Z(n2188) );
  OR U4180 ( .A(n2186), .B(n2185), .Z(n2187) );
  NAND U4181 ( .A(n2188), .B(n2187), .Z(n2833) );
  XNOR U4182 ( .A(n2834), .B(n2833), .Z(n2836) );
  OR U4183 ( .A(n2190), .B(n2189), .Z(n2194) );
  OR U4184 ( .A(n2192), .B(n2191), .Z(n2193) );
  NAND U4185 ( .A(n2194), .B(n2193), .Z(n2835) );
  XOR U4186 ( .A(n2836), .B(n2835), .Z(n2938) );
  XOR U4187 ( .A(n2937), .B(n2938), .Z(n2939) );
  XOR U4188 ( .A(n2940), .B(n2939), .Z(n3705) );
  XNOR U4189 ( .A(n3704), .B(n3705), .Z(n3706) );
  OR U4190 ( .A(n2196), .B(n2195), .Z(n2200) );
  OR U4191 ( .A(n2198), .B(n2197), .Z(n2199) );
  AND U4192 ( .A(n2200), .B(n2199), .Z(n2847) );
  OR U4193 ( .A(n2202), .B(n2201), .Z(n2206) );
  OR U4194 ( .A(n2204), .B(n2203), .Z(n2205) );
  NAND U4195 ( .A(n2206), .B(n2205), .Z(n3553) );
  OR U4196 ( .A(n2208), .B(n2207), .Z(n2212) );
  OR U4197 ( .A(n2210), .B(n2209), .Z(n2211) );
  AND U4198 ( .A(n2212), .B(n2211), .Z(n3552) );
  XOR U4199 ( .A(n3553), .B(n3552), .Z(n3555) );
  OR U4200 ( .A(n2214), .B(n2213), .Z(n2218) );
  OR U4201 ( .A(n2216), .B(n2215), .Z(n2217) );
  NAND U4202 ( .A(n2218), .B(n2217), .Z(n3554) );
  XOR U4203 ( .A(n3555), .B(n3554), .Z(n2845) );
  OR U4204 ( .A(n2220), .B(n2219), .Z(n2224) );
  OR U4205 ( .A(n2222), .B(n2221), .Z(n2223) );
  NAND U4206 ( .A(n2224), .B(n2223), .Z(n2744) );
  OR U4207 ( .A(n2226), .B(n2225), .Z(n2230) );
  OR U4208 ( .A(n2228), .B(n2227), .Z(n2229) );
  NAND U4209 ( .A(n2230), .B(n2229), .Z(n2743) );
  XNOR U4210 ( .A(n2744), .B(n2743), .Z(n2746) );
  OR U4211 ( .A(n2232), .B(n2231), .Z(n2236) );
  OR U4212 ( .A(n2234), .B(n2233), .Z(n2235) );
  NAND U4213 ( .A(n2236), .B(n2235), .Z(n2745) );
  XOR U4214 ( .A(n2746), .B(n2745), .Z(n2846) );
  XNOR U4215 ( .A(n2845), .B(n2846), .Z(n2848) );
  XNOR U4216 ( .A(n2847), .B(n2848), .Z(n3707) );
  XNOR U4217 ( .A(n3706), .B(n3707), .Z(n3176) );
  NAND U4218 ( .A(n2238), .B(n2237), .Z(n2242) );
  NAND U4219 ( .A(n2240), .B(n2239), .Z(n2241) );
  NAND U4220 ( .A(n2242), .B(n2241), .Z(n3242) );
  NAND U4221 ( .A(n2244), .B(n2243), .Z(n2248) );
  NAND U4222 ( .A(n2246), .B(n2245), .Z(n2247) );
  NAND U4223 ( .A(n2248), .B(n2247), .Z(n3240) );
  OR U4224 ( .A(n2254), .B(n2253), .Z(n2258) );
  NANDN U4225 ( .A(n2256), .B(n2255), .Z(n2257) );
  AND U4226 ( .A(n2258), .B(n2257), .Z(n2963) );
  XOR U4227 ( .A(n2963), .B(n2964), .Z(n2966) );
  XOR U4228 ( .A(n2965), .B(n2966), .Z(n3239) );
  XOR U4229 ( .A(n3240), .B(n3239), .Z(n3241) );
  XOR U4230 ( .A(n3242), .B(n3241), .Z(n3712) );
  NANDN U4231 ( .A(n2264), .B(n2263), .Z(n2268) );
  NAND U4232 ( .A(n2266), .B(n2265), .Z(n2267) );
  NAND U4233 ( .A(n2268), .B(n2267), .Z(n3319) );
  OR U4234 ( .A(n2270), .B(n2269), .Z(n2274) );
  OR U4235 ( .A(n2272), .B(n2271), .Z(n2273) );
  NAND U4236 ( .A(n2274), .B(n2273), .Z(n3115) );
  OR U4237 ( .A(n2276), .B(n2275), .Z(n2280) );
  OR U4238 ( .A(n2278), .B(n2277), .Z(n2279) );
  NAND U4239 ( .A(n2280), .B(n2279), .Z(n3114) );
  XNOR U4240 ( .A(n3115), .B(n3114), .Z(n3117) );
  OR U4241 ( .A(n2282), .B(n2281), .Z(n2286) );
  OR U4242 ( .A(n2284), .B(n2283), .Z(n2285) );
  NAND U4243 ( .A(n2286), .B(n2285), .Z(n3116) );
  XNOR U4244 ( .A(n3117), .B(n3116), .Z(n3317) );
  NAND U4245 ( .A(n2288), .B(n2287), .Z(n2292) );
  NAND U4246 ( .A(n2290), .B(n2289), .Z(n2291) );
  AND U4247 ( .A(n2292), .B(n2291), .Z(n3318) );
  XOR U4248 ( .A(n3317), .B(n3318), .Z(n3320) );
  XOR U4249 ( .A(n3319), .B(n3320), .Z(n3710) );
  OR U4250 ( .A(n2298), .B(n2297), .Z(n2302) );
  OR U4251 ( .A(n2300), .B(n2299), .Z(n2301) );
  NAND U4252 ( .A(n2302), .B(n2301), .Z(n3121) );
  OR U4253 ( .A(n2304), .B(n2303), .Z(n2308) );
  OR U4254 ( .A(n2306), .B(n2305), .Z(n2307) );
  NAND U4255 ( .A(n2308), .B(n2307), .Z(n3120) );
  XNOR U4256 ( .A(n3121), .B(n3120), .Z(n3123) );
  OR U4257 ( .A(n2310), .B(n2309), .Z(n2314) );
  NANDN U4258 ( .A(n2312), .B(n2311), .Z(n2313) );
  NAND U4259 ( .A(n2314), .B(n2313), .Z(n3122) );
  XNOR U4260 ( .A(n3123), .B(n3122), .Z(n3305) );
  NAND U4261 ( .A(n2316), .B(n2315), .Z(n2320) );
  OR U4262 ( .A(n2318), .B(n2317), .Z(n2319) );
  AND U4263 ( .A(n2320), .B(n2319), .Z(n3306) );
  XOR U4264 ( .A(n3305), .B(n3306), .Z(n3308) );
  XOR U4265 ( .A(n3307), .B(n3308), .Z(n3711) );
  XNOR U4266 ( .A(n3710), .B(n3711), .Z(n3713) );
  XNOR U4267 ( .A(n3712), .B(n3713), .Z(n3175) );
  XNOR U4268 ( .A(n3176), .B(n3175), .Z(n3177) );
  XNOR U4269 ( .A(n3178), .B(n3177), .Z(n3677) );
  OR U4270 ( .A(n2326), .B(n2325), .Z(n2330) );
  OR U4271 ( .A(n2328), .B(n2327), .Z(n2329) );
  NAND U4272 ( .A(n2330), .B(n2329), .Z(n3635) );
  OR U4273 ( .A(n2332), .B(n2331), .Z(n2336) );
  OR U4274 ( .A(n2334), .B(n2333), .Z(n2335) );
  AND U4275 ( .A(n2336), .B(n2335), .Z(n3634) );
  XOR U4276 ( .A(n3635), .B(n3634), .Z(n3637) );
  XOR U4277 ( .A(n3637), .B(n3636), .Z(n2967) );
  OR U4278 ( .A(n2342), .B(n2341), .Z(n2346) );
  OR U4279 ( .A(n2344), .B(n2343), .Z(n2345) );
  NAND U4280 ( .A(n2346), .B(n2345), .Z(n2968) );
  XNOR U4281 ( .A(n2967), .B(n2968), .Z(n2969) );
  XNOR U4282 ( .A(n2970), .B(n2969), .Z(n3735) );
  NAND U4283 ( .A(n2348), .B(n2347), .Z(n2352) );
  NAND U4284 ( .A(n2350), .B(n2349), .Z(n2351) );
  NAND U4285 ( .A(n2352), .B(n2351), .Z(n3733) );
  OR U4286 ( .A(n2354), .B(n2353), .Z(n2358) );
  OR U4287 ( .A(n2356), .B(n2355), .Z(n2357) );
  NAND U4288 ( .A(n2358), .B(n2357), .Z(n3522) );
  OR U4289 ( .A(n2360), .B(n2359), .Z(n2364) );
  OR U4290 ( .A(n2362), .B(n2361), .Z(n2363) );
  NAND U4291 ( .A(n2364), .B(n2363), .Z(n3521) );
  XNOR U4292 ( .A(n3522), .B(n3521), .Z(n3524) );
  XNOR U4293 ( .A(n3524), .B(n3523), .Z(n3518) );
  OR U4294 ( .A(n2370), .B(n2369), .Z(n2374) );
  OR U4295 ( .A(n2372), .B(n2371), .Z(n2373) );
  AND U4296 ( .A(n2374), .B(n2373), .Z(n3517) );
  XOR U4297 ( .A(n3518), .B(n3517), .Z(n3519) );
  OR U4298 ( .A(n2376), .B(n2375), .Z(n2380) );
  OR U4299 ( .A(n2378), .B(n2377), .Z(n2379) );
  NAND U4300 ( .A(n2380), .B(n2379), .Z(n3534) );
  OR U4301 ( .A(n2382), .B(n2381), .Z(n2386) );
  OR U4302 ( .A(n2384), .B(n2383), .Z(n2385) );
  NAND U4303 ( .A(n2386), .B(n2385), .Z(n3533) );
  XNOR U4304 ( .A(n3534), .B(n3533), .Z(n3536) );
  OR U4305 ( .A(n2388), .B(n2387), .Z(n2392) );
  OR U4306 ( .A(n2390), .B(n2389), .Z(n2391) );
  NAND U4307 ( .A(n2392), .B(n2391), .Z(n3535) );
  XOR U4308 ( .A(n3536), .B(n3535), .Z(n3520) );
  XOR U4309 ( .A(n3519), .B(n3520), .Z(n3732) );
  XOR U4310 ( .A(n3733), .B(n3732), .Z(n3734) );
  XNOR U4311 ( .A(n3735), .B(n3734), .Z(n3131) );
  OR U4312 ( .A(n2394), .B(n2393), .Z(n2398) );
  OR U4313 ( .A(n2396), .B(n2395), .Z(n2397) );
  NAND U4314 ( .A(n2398), .B(n2397), .Z(n3428) );
  OR U4315 ( .A(n2400), .B(n2399), .Z(n2404) );
  OR U4316 ( .A(n2402), .B(n2401), .Z(n2403) );
  NAND U4317 ( .A(n2404), .B(n2403), .Z(n3103) );
  OR U4318 ( .A(n2406), .B(n2405), .Z(n2410) );
  OR U4319 ( .A(n2408), .B(n2407), .Z(n2409) );
  NAND U4320 ( .A(n2410), .B(n2409), .Z(n3102) );
  XOR U4321 ( .A(n3103), .B(n3102), .Z(n3104) );
  OR U4322 ( .A(n2412), .B(n2411), .Z(n2416) );
  OR U4323 ( .A(n2414), .B(n2413), .Z(n2415) );
  NAND U4324 ( .A(n2416), .B(n2415), .Z(n3105) );
  XNOR U4325 ( .A(n3104), .B(n3105), .Z(n3425) );
  OR U4326 ( .A(n2418), .B(n2417), .Z(n2422) );
  NANDN U4327 ( .A(n2420), .B(n2419), .Z(n2421) );
  NAND U4328 ( .A(n2422), .B(n2421), .Z(n3426) );
  XOR U4329 ( .A(n3425), .B(n3426), .Z(n3427) );
  XNOR U4330 ( .A(n3428), .B(n3427), .Z(n3760) );
  OR U4331 ( .A(n2424), .B(n2423), .Z(n2428) );
  OR U4332 ( .A(n2426), .B(n2425), .Z(n2427) );
  NAND U4333 ( .A(n2428), .B(n2427), .Z(n2792) );
  OR U4334 ( .A(n2430), .B(n2429), .Z(n2434) );
  OR U4335 ( .A(n2432), .B(n2431), .Z(n2433) );
  NAND U4336 ( .A(n2434), .B(n2433), .Z(n2791) );
  XNOR U4337 ( .A(n2792), .B(n2791), .Z(n2794) );
  OR U4338 ( .A(n2436), .B(n2435), .Z(n2440) );
  OR U4339 ( .A(n2438), .B(n2437), .Z(n2439) );
  NAND U4340 ( .A(n2440), .B(n2439), .Z(n2793) );
  XNOR U4341 ( .A(n2794), .B(n2793), .Z(n2907) );
  OR U4342 ( .A(n2442), .B(n2441), .Z(n2446) );
  NANDN U4343 ( .A(n2444), .B(n2443), .Z(n2445) );
  NAND U4344 ( .A(n2446), .B(n2445), .Z(n3617) );
  XNOR U4345 ( .A(n3617), .B(n3616), .Z(n3618) );
  OR U4346 ( .A(n2452), .B(n2451), .Z(n2456) );
  OR U4347 ( .A(n2454), .B(n2453), .Z(n2455) );
  NAND U4348 ( .A(n2456), .B(n2455), .Z(n3619) );
  XNOR U4349 ( .A(n3618), .B(n3619), .Z(n2905) );
  XNOR U4350 ( .A(n2852), .B(n2851), .Z(n2854) );
  XOR U4351 ( .A(n2854), .B(n2853), .Z(n2906) );
  XOR U4352 ( .A(n2905), .B(n2906), .Z(n2908) );
  XOR U4353 ( .A(n2907), .B(n2908), .Z(n3758) );
  NANDN U4354 ( .A(n2470), .B(n2469), .Z(n2474) );
  NANDN U4355 ( .A(n2472), .B(n2471), .Z(n2473) );
  NAND U4356 ( .A(n2474), .B(n2473), .Z(n3759) );
  XNOR U4357 ( .A(n3758), .B(n3759), .Z(n3761) );
  XOR U4358 ( .A(n3760), .B(n3761), .Z(n3130) );
  XNOR U4359 ( .A(n3131), .B(n3130), .Z(n3133) );
  OR U4360 ( .A(n2476), .B(n2475), .Z(n2480) );
  OR U4361 ( .A(n2478), .B(n2477), .Z(n2479) );
  NAND U4362 ( .A(n2480), .B(n2479), .Z(n3071) );
  OR U4363 ( .A(n2482), .B(n2481), .Z(n2486) );
  OR U4364 ( .A(n2484), .B(n2483), .Z(n2485) );
  NAND U4365 ( .A(n2486), .B(n2485), .Z(n3070) );
  XNOR U4366 ( .A(n3071), .B(n3070), .Z(n3073) );
  XNOR U4367 ( .A(n3073), .B(n3072), .Z(n3588) );
  OR U4368 ( .A(n2492), .B(n2491), .Z(n2496) );
  OR U4369 ( .A(n2494), .B(n2493), .Z(n2495) );
  NAND U4370 ( .A(n2496), .B(n2495), .Z(n3569) );
  OR U4371 ( .A(n2498), .B(n2497), .Z(n2502) );
  OR U4372 ( .A(n2500), .B(n2499), .Z(n2501) );
  AND U4373 ( .A(n2502), .B(n2501), .Z(n3568) );
  XNOR U4374 ( .A(n3569), .B(n3568), .Z(n3570) );
  OR U4375 ( .A(n2504), .B(n2503), .Z(n2508) );
  OR U4376 ( .A(n2506), .B(n2505), .Z(n2507) );
  AND U4377 ( .A(n2508), .B(n2507), .Z(n3571) );
  XNOR U4378 ( .A(n3570), .B(n3571), .Z(n3587) );
  OR U4379 ( .A(n2510), .B(n2509), .Z(n2514) );
  OR U4380 ( .A(n2512), .B(n2511), .Z(n2513) );
  NAND U4381 ( .A(n2514), .B(n2513), .Z(n3586) );
  XOR U4382 ( .A(n3587), .B(n3586), .Z(n3589) );
  XOR U4383 ( .A(n3588), .B(n3589), .Z(n3731) );
  OR U4384 ( .A(n2516), .B(n2515), .Z(n2520) );
  OR U4385 ( .A(n2518), .B(n2517), .Z(n2519) );
  NAND U4386 ( .A(n2520), .B(n2519), .Z(n3093) );
  OR U4387 ( .A(n2522), .B(n2521), .Z(n2526) );
  OR U4388 ( .A(n2524), .B(n2523), .Z(n2525) );
  NAND U4389 ( .A(n2526), .B(n2525), .Z(n3092) );
  XNOR U4390 ( .A(n3093), .B(n3092), .Z(n3095) );
  OR U4391 ( .A(n2528), .B(n2527), .Z(n2532) );
  OR U4392 ( .A(n2530), .B(n2529), .Z(n2531) );
  NAND U4393 ( .A(n2532), .B(n2531), .Z(n3094) );
  XNOR U4394 ( .A(n3095), .B(n3094), .Z(n3076) );
  OR U4395 ( .A(n2534), .B(n2533), .Z(n2538) );
  OR U4396 ( .A(n2536), .B(n2535), .Z(n2537) );
  NAND U4397 ( .A(n2538), .B(n2537), .Z(n3530) );
  OR U4398 ( .A(n2544), .B(n2543), .Z(n2548) );
  OR U4399 ( .A(n2546), .B(n2545), .Z(n2547) );
  AND U4400 ( .A(n2548), .B(n2547), .Z(n3528) );
  XNOR U4401 ( .A(n3527), .B(n3528), .Z(n3529) );
  XNOR U4402 ( .A(n3530), .B(n3529), .Z(n3077) );
  XOR U4403 ( .A(n3076), .B(n3077), .Z(n3079) );
  NAND U4404 ( .A(n2550), .B(n2549), .Z(n2554) );
  NAND U4405 ( .A(n2552), .B(n2551), .Z(n2553) );
  NAND U4406 ( .A(n2554), .B(n2553), .Z(n3078) );
  XOR U4407 ( .A(n3079), .B(n3078), .Z(n3728) );
  OR U4408 ( .A(n2556), .B(n2555), .Z(n2560) );
  NAND U4409 ( .A(n2558), .B(n2557), .Z(n2559) );
  NAND U4410 ( .A(n2560), .B(n2559), .Z(n3729) );
  XOR U4411 ( .A(n3728), .B(n3729), .Z(n3730) );
  XNOR U4412 ( .A(n3731), .B(n3730), .Z(n3132) );
  XOR U4413 ( .A(n3133), .B(n3132), .Z(n3676) );
  XOR U4414 ( .A(n3677), .B(n3676), .Z(n3678) );
  XNOR U4415 ( .A(n3679), .B(n3678), .Z(n3791) );
  NAND U4416 ( .A(n2562), .B(n2561), .Z(n2566) );
  NAND U4417 ( .A(n2564), .B(n2563), .Z(n2565) );
  NAND U4418 ( .A(n2566), .B(n2565), .Z(n3785) );
  NANDN U4419 ( .A(n2572), .B(n2571), .Z(n2576) );
  NAND U4420 ( .A(n2574), .B(n2573), .Z(n2575) );
  NAND U4421 ( .A(n2576), .B(n2575), .Z(n3779) );
  NANDN U4422 ( .A(n2578), .B(n2577), .Z(n2582) );
  NAND U4423 ( .A(n2580), .B(n2579), .Z(n2581) );
  NAND U4424 ( .A(n2582), .B(n2581), .Z(n3776) );
  OR U4425 ( .A(n2584), .B(n2583), .Z(n2588) );
  OR U4426 ( .A(n2586), .B(n2585), .Z(n2587) );
  AND U4427 ( .A(n2588), .B(n2587), .Z(n3777) );
  XNOR U4428 ( .A(n3776), .B(n3777), .Z(n3778) );
  XNOR U4429 ( .A(n3779), .B(n3778), .Z(n3783) );
  XNOR U4430 ( .A(n3782), .B(n3783), .Z(n3784) );
  XNOR U4431 ( .A(n3785), .B(n3784), .Z(n3205) );
  NAND U4432 ( .A(n2590), .B(n2589), .Z(n2594) );
  NANDN U4433 ( .A(n2592), .B(n2591), .Z(n2593) );
  NAND U4434 ( .A(n2594), .B(n2593), .Z(n3745) );
  NANDN U4435 ( .A(n2596), .B(n2595), .Z(n2600) );
  NANDN U4436 ( .A(n2598), .B(n2597), .Z(n2599) );
  AND U4437 ( .A(n2600), .B(n2599), .Z(n2780) );
  OR U4438 ( .A(n2602), .B(n2601), .Z(n2606) );
  NANDN U4439 ( .A(n2604), .B(n2603), .Z(n2605) );
  NAND U4440 ( .A(n2606), .B(n2605), .Z(n3292) );
  NANDN U4441 ( .A(n2608), .B(n2607), .Z(n2612) );
  NAND U4442 ( .A(n2610), .B(n2609), .Z(n2611) );
  NAND U4443 ( .A(n2612), .B(n2611), .Z(n3290) );
  XOR U4444 ( .A(n2942), .B(n2941), .Z(n2944) );
  XOR U4445 ( .A(n2944), .B(n2943), .Z(n3289) );
  XNOR U4446 ( .A(n3290), .B(n3289), .Z(n3291) );
  XNOR U4447 ( .A(n3292), .B(n3291), .Z(n2777) );
  NANDN U4448 ( .A(n2626), .B(n2625), .Z(n2630) );
  NANDN U4449 ( .A(n2628), .B(n2627), .Z(n2629) );
  NAND U4450 ( .A(n2630), .B(n2629), .Z(n2778) );
  XNOR U4451 ( .A(n2777), .B(n2778), .Z(n2779) );
  XOR U4452 ( .A(n2780), .B(n2779), .Z(n3743) );
  NAND U4453 ( .A(n2632), .B(n2631), .Z(n2636) );
  NAND U4454 ( .A(n2634), .B(n2633), .Z(n2635) );
  AND U4455 ( .A(n2636), .B(n2635), .Z(n3742) );
  XOR U4456 ( .A(n3743), .B(n3742), .Z(n3744) );
  XNOR U4457 ( .A(n3745), .B(n3744), .Z(n3204) );
  NANDN U4458 ( .A(n2642), .B(n2641), .Z(n2646) );
  NAND U4459 ( .A(n2644), .B(n2643), .Z(n2645) );
  NAND U4460 ( .A(n2646), .B(n2645), .Z(n3514) );
  NAND U4461 ( .A(n2648), .B(n2647), .Z(n2652) );
  NANDN U4462 ( .A(n2650), .B(n2649), .Z(n2651) );
  NAND U4463 ( .A(n2652), .B(n2651), .Z(n3511) );
  XNOR U4464 ( .A(n3511), .B(n3512), .Z(n3513) );
  XNOR U4465 ( .A(n3514), .B(n3513), .Z(n3682) );
  XOR U4466 ( .A(n2768), .B(n2767), .Z(n2769) );
  XOR U4467 ( .A(n2769), .B(n2770), .Z(n2783) );
  OR U4468 ( .A(n2674), .B(n2673), .Z(n2678) );
  OR U4469 ( .A(n2676), .B(n2675), .Z(n2677) );
  NAND U4470 ( .A(n2678), .B(n2677), .Z(n2911) );
  XOR U4471 ( .A(n2912), .B(n2911), .Z(n2913) );
  OR U4472 ( .A(n2680), .B(n2679), .Z(n2684) );
  OR U4473 ( .A(n2682), .B(n2681), .Z(n2683) );
  NAND U4474 ( .A(n2684), .B(n2683), .Z(n2914) );
  XNOR U4475 ( .A(n2913), .B(n2914), .Z(n2781) );
  OR U4476 ( .A(n2686), .B(n2685), .Z(n2690) );
  OR U4477 ( .A(n2688), .B(n2687), .Z(n2689) );
  NAND U4478 ( .A(n2690), .B(n2689), .Z(n3599) );
  XOR U4479 ( .A(n3599), .B(n3598), .Z(n3601) );
  XOR U4480 ( .A(n3601), .B(n3600), .Z(n2782) );
  XOR U4481 ( .A(n2781), .B(n2782), .Z(n2784) );
  XOR U4482 ( .A(n2783), .B(n2784), .Z(n2821) );
  OR U4483 ( .A(n2700), .B(n2699), .Z(n2704) );
  NANDN U4484 ( .A(n2702), .B(n2701), .Z(n2703) );
  AND U4485 ( .A(n2704), .B(n2703), .Z(n2822) );
  XNOR U4486 ( .A(n2821), .B(n2822), .Z(n2824) );
  XOR U4487 ( .A(n3111), .B(n3110), .Z(n3113) );
  XOR U4488 ( .A(n3113), .B(n3112), .Z(n3394) );
  XOR U4489 ( .A(n3393), .B(n3394), .Z(n3395) );
  XNOR U4490 ( .A(n3396), .B(n3395), .Z(n2823) );
  XNOR U4491 ( .A(n2824), .B(n2823), .Z(n3683) );
  XOR U4492 ( .A(n3682), .B(n3683), .Z(n3685) );
  XOR U4493 ( .A(n3684), .B(n3685), .Z(n3203) );
  XNOR U4494 ( .A(n3204), .B(n3203), .Z(n3206) );
  XOR U4495 ( .A(n3205), .B(n3206), .Z(n3788) );
  NANDN U4496 ( .A(n2726), .B(n2725), .Z(n2730) );
  NAND U4497 ( .A(n2728), .B(n2727), .Z(n2729) );
  NAND U4498 ( .A(n2730), .B(n2729), .Z(n3789) );
  XNOR U4499 ( .A(n3788), .B(n3789), .Z(n3790) );
  XOR U4500 ( .A(n3791), .B(n3790), .Z(n3224) );
  XNOR U4501 ( .A(n3223), .B(n3224), .Z(o[1]) );
  OR U4502 ( .A(n2732), .B(n2731), .Z(n2736) );
  NANDN U4503 ( .A(n2734), .B(n2733), .Z(n2735) );
  AND U4504 ( .A(n2736), .B(n2735), .Z(n4208) );
  NANDN U4505 ( .A(n2738), .B(n2737), .Z(n2742) );
  NAND U4506 ( .A(n2740), .B(n2739), .Z(n2741) );
  NAND U4507 ( .A(n2742), .B(n2741), .Z(n4236) );
  OR U4508 ( .A(n2744), .B(n2743), .Z(n2748) );
  OR U4509 ( .A(n2746), .B(n2745), .Z(n2747) );
  NAND U4510 ( .A(n2748), .B(n2747), .Z(n4190) );
  OR U4511 ( .A(n2750), .B(n2749), .Z(n2754) );
  OR U4512 ( .A(n2752), .B(n2751), .Z(n2753) );
  AND U4513 ( .A(n2754), .B(n2753), .Z(n4188) );
  OR U4514 ( .A(n2756), .B(n2755), .Z(n2760) );
  OR U4515 ( .A(n2758), .B(n2757), .Z(n2759) );
  NAND U4516 ( .A(n2760), .B(n2759), .Z(n4189) );
  XOR U4517 ( .A(n4188), .B(n4189), .Z(n4191) );
  XOR U4518 ( .A(n4190), .B(n4191), .Z(n4235) );
  XOR U4519 ( .A(n4236), .B(n4235), .Z(n4237) );
  OR U4520 ( .A(n2762), .B(n2761), .Z(n2766) );
  OR U4521 ( .A(n2764), .B(n2763), .Z(n2765) );
  NAND U4522 ( .A(n2766), .B(n2765), .Z(n4221) );
  OR U4523 ( .A(n2772), .B(n2771), .Z(n2776) );
  OR U4524 ( .A(n2774), .B(n2773), .Z(n2775) );
  NAND U4525 ( .A(n2776), .B(n2775), .Z(n4220) );
  XOR U4526 ( .A(n4219), .B(n4220), .Z(n4222) );
  XOR U4527 ( .A(n4221), .B(n4222), .Z(n4238) );
  XOR U4528 ( .A(n4237), .B(n4238), .Z(n4039) );
  OR U4529 ( .A(n2786), .B(n2785), .Z(n2790) );
  OR U4530 ( .A(n2788), .B(n2787), .Z(n2789) );
  NAND U4531 ( .A(n2790), .B(n2789), .Z(n4194) );
  OR U4532 ( .A(n2792), .B(n2791), .Z(n2796) );
  OR U4533 ( .A(n2794), .B(n2793), .Z(n2795) );
  NAND U4534 ( .A(n2796), .B(n2795), .Z(n4193) );
  OR U4535 ( .A(n2798), .B(n2797), .Z(n2802) );
  OR U4536 ( .A(n2800), .B(n2799), .Z(n2801) );
  NAND U4537 ( .A(n2802), .B(n2801), .Z(n4192) );
  XOR U4538 ( .A(n4193), .B(n4192), .Z(n4195) );
  XOR U4539 ( .A(n4194), .B(n4195), .Z(n3827) );
  XOR U4540 ( .A(n3828), .B(n3827), .Z(n3829) );
  OR U4541 ( .A(n2804), .B(n2803), .Z(n2808) );
  OR U4542 ( .A(n2806), .B(n2805), .Z(n2807) );
  NAND U4543 ( .A(n2808), .B(n2807), .Z(n3921) );
  OR U4544 ( .A(n2810), .B(n2809), .Z(n2814) );
  OR U4545 ( .A(n2812), .B(n2811), .Z(n2813) );
  AND U4546 ( .A(n2814), .B(n2813), .Z(n3919) );
  OR U4547 ( .A(n2816), .B(n2815), .Z(n2820) );
  OR U4548 ( .A(n2818), .B(n2817), .Z(n2819) );
  NAND U4549 ( .A(n2820), .B(n2819), .Z(n3920) );
  XOR U4550 ( .A(n3919), .B(n3920), .Z(n3922) );
  XOR U4551 ( .A(n3921), .B(n3922), .Z(n3830) );
  XOR U4552 ( .A(n3829), .B(n3830), .Z(n4036) );
  XOR U4553 ( .A(n4037), .B(n4036), .Z(n4038) );
  XNOR U4554 ( .A(n4039), .B(n4038), .Z(n4207) );
  XOR U4555 ( .A(n4208), .B(n4207), .Z(n4210) );
  OR U4556 ( .A(n2822), .B(n2821), .Z(n2826) );
  NANDN U4557 ( .A(n2824), .B(n2823), .Z(n2825) );
  AND U4558 ( .A(n2826), .B(n2825), .Z(n4033) );
  OR U4559 ( .A(n2828), .B(n2827), .Z(n2832) );
  OR U4560 ( .A(n2830), .B(n2829), .Z(n2831) );
  AND U4561 ( .A(n2832), .B(n2831), .Z(n4229) );
  OR U4562 ( .A(n2834), .B(n2833), .Z(n2838) );
  OR U4563 ( .A(n2836), .B(n2835), .Z(n2837) );
  AND U4564 ( .A(n2838), .B(n2837), .Z(n4227) );
  OR U4565 ( .A(n2840), .B(n2839), .Z(n2844) );
  OR U4566 ( .A(n2842), .B(n2841), .Z(n2843) );
  AND U4567 ( .A(n2844), .B(n2843), .Z(n4228) );
  XOR U4568 ( .A(n4227), .B(n4228), .Z(n4230) );
  XOR U4569 ( .A(n4229), .B(n4230), .Z(n4245) );
  OR U4570 ( .A(n2846), .B(n2845), .Z(n2850) );
  OR U4571 ( .A(n2848), .B(n2847), .Z(n2849) );
  AND U4572 ( .A(n2850), .B(n2849), .Z(n4246) );
  XOR U4573 ( .A(n4245), .B(n4246), .Z(n4248) );
  OR U4574 ( .A(n2852), .B(n2851), .Z(n2856) );
  OR U4575 ( .A(n2854), .B(n2853), .Z(n2855) );
  NAND U4576 ( .A(n2856), .B(n2855), .Z(n4150) );
  OR U4577 ( .A(n2858), .B(n2857), .Z(n2862) );
  OR U4578 ( .A(n2860), .B(n2859), .Z(n2861) );
  AND U4579 ( .A(n2862), .B(n2861), .Z(n4148) );
  OR U4580 ( .A(n2864), .B(n2863), .Z(n2868) );
  OR U4581 ( .A(n2866), .B(n2865), .Z(n2867) );
  NAND U4582 ( .A(n2868), .B(n2867), .Z(n4149) );
  XOR U4583 ( .A(n4148), .B(n4149), .Z(n4151) );
  XOR U4584 ( .A(n4150), .B(n4151), .Z(n4247) );
  XOR U4585 ( .A(n4248), .B(n4247), .Z(n4032) );
  XOR U4586 ( .A(n4033), .B(n4032), .Z(n4035) );
  OR U4587 ( .A(n2870), .B(n2869), .Z(n2874) );
  OR U4588 ( .A(n2872), .B(n2871), .Z(n2873) );
  AND U4589 ( .A(n2874), .B(n2873), .Z(n3835) );
  OR U4590 ( .A(n2876), .B(n2875), .Z(n2880) );
  OR U4591 ( .A(n2878), .B(n2877), .Z(n2879) );
  AND U4592 ( .A(n2880), .B(n2879), .Z(n3833) );
  OR U4593 ( .A(n2882), .B(n2881), .Z(n2886) );
  OR U4594 ( .A(n2884), .B(n2883), .Z(n2885) );
  AND U4595 ( .A(n2886), .B(n2885), .Z(n3834) );
  XOR U4596 ( .A(n3833), .B(n3834), .Z(n3836) );
  XOR U4597 ( .A(n3835), .B(n3836), .Z(n4251) );
  OR U4598 ( .A(n2896), .B(n2895), .Z(n2900) );
  OR U4599 ( .A(n2898), .B(n2897), .Z(n2899) );
  AND U4600 ( .A(n2900), .B(n2899), .Z(n4232) );
  XOR U4601 ( .A(n4231), .B(n4232), .Z(n4234) );
  XOR U4602 ( .A(n4233), .B(n4234), .Z(n4249) );
  XOR U4603 ( .A(n4249), .B(n4250), .Z(n4252) );
  XOR U4604 ( .A(n4251), .B(n4252), .Z(n4034) );
  XOR U4605 ( .A(n4035), .B(n4034), .Z(n4209) );
  XNOR U4606 ( .A(n4210), .B(n4209), .Z(n4120) );
  OR U4607 ( .A(n2906), .B(n2905), .Z(n2910) );
  NAND U4608 ( .A(n2908), .B(n2907), .Z(n2909) );
  NAND U4609 ( .A(n2910), .B(n2909), .Z(n4007) );
  XOR U4610 ( .A(n3951), .B(n3952), .Z(n3954) );
  XOR U4611 ( .A(n3953), .B(n3954), .Z(n4006) );
  XOR U4612 ( .A(n4007), .B(n4006), .Z(n4008) );
  OR U4613 ( .A(n2932), .B(n2931), .Z(n2936) );
  OR U4614 ( .A(n2934), .B(n2933), .Z(n2935) );
  AND U4615 ( .A(n2936), .B(n2935), .Z(n3914) );
  XNOR U4616 ( .A(n3913), .B(n3914), .Z(n3916) );
  XNOR U4617 ( .A(n3915), .B(n3916), .Z(n4009) );
  XNOR U4618 ( .A(n4008), .B(n4009), .Z(n4053) );
  XOR U4619 ( .A(n3907), .B(n3908), .Z(n3909) );
  XOR U4620 ( .A(n3910), .B(n3909), .Z(n3887) );
  XNOR U4621 ( .A(n3888), .B(n3887), .Z(n3890) );
  OR U4622 ( .A(n2958), .B(n2957), .Z(n2962) );
  OR U4623 ( .A(n2960), .B(n2959), .Z(n2961) );
  AND U4624 ( .A(n2962), .B(n2961), .Z(n4178) );
  XOR U4625 ( .A(n4178), .B(n4179), .Z(n4180) );
  XNOR U4626 ( .A(n4181), .B(n4180), .Z(n3889) );
  XNOR U4627 ( .A(n3890), .B(n3889), .Z(n4054) );
  XOR U4628 ( .A(n4053), .B(n4054), .Z(n4055) );
  OR U4629 ( .A(n2968), .B(n2967), .Z(n2972) );
  OR U4630 ( .A(n2970), .B(n2969), .Z(n2971) );
  AND U4631 ( .A(n2972), .B(n2971), .Z(n3872) );
  OR U4632 ( .A(n2982), .B(n2981), .Z(n2986) );
  OR U4633 ( .A(n2984), .B(n2983), .Z(n2985) );
  AND U4634 ( .A(n2986), .B(n2985), .Z(n3924) );
  XNOR U4635 ( .A(n3923), .B(n3924), .Z(n3925) );
  XNOR U4636 ( .A(n3926), .B(n3925), .Z(n3869) );
  XOR U4637 ( .A(n3927), .B(n3928), .Z(n3929) );
  XNOR U4638 ( .A(n3930), .B(n3929), .Z(n3870) );
  XNOR U4639 ( .A(n3869), .B(n3870), .Z(n3871) );
  XOR U4640 ( .A(n3872), .B(n3871), .Z(n4056) );
  XNOR U4641 ( .A(n4055), .B(n4056), .Z(n4026) );
  NANDN U4642 ( .A(n3000), .B(n2999), .Z(n3004) );
  OR U4643 ( .A(n3002), .B(n3001), .Z(n3003) );
  NAND U4644 ( .A(n3004), .B(n3003), .Z(n4025) );
  IV U4645 ( .A(n3017), .Z(n3018) );
  NANDN U4646 ( .A(n3019), .B(n3018), .Z(n3023) );
  NANDN U4647 ( .A(n3021), .B(n3020), .Z(n3022) );
  NAND U4648 ( .A(n3023), .B(n3022), .Z(n4002) );
  XNOR U4649 ( .A(n4003), .B(n4002), .Z(n4004) );
  XOR U4650 ( .A(n4005), .B(n4004), .Z(n4242) );
  XOR U4651 ( .A(n4241), .B(n4242), .Z(n4243) );
  XOR U4652 ( .A(n4243), .B(n4244), .Z(n4024) );
  XOR U4653 ( .A(n4025), .B(n4024), .Z(n4027) );
  XOR U4654 ( .A(n4026), .B(n4027), .Z(n4119) );
  XOR U4655 ( .A(n4120), .B(n4119), .Z(n4121) );
  OR U4656 ( .A(n3029), .B(n3028), .Z(n3033) );
  OR U4657 ( .A(n3031), .B(n3030), .Z(n3032) );
  AND U4658 ( .A(n3033), .B(n3032), .Z(n3840) );
  OR U4659 ( .A(n3039), .B(n3038), .Z(n3043) );
  OR U4660 ( .A(n3041), .B(n3040), .Z(n3042) );
  AND U4661 ( .A(n3043), .B(n3042), .Z(n3838) );
  XNOR U4662 ( .A(n3837), .B(n3838), .Z(n3839) );
  XNOR U4663 ( .A(n3840), .B(n3839), .Z(n3823) );
  XNOR U4664 ( .A(n4153), .B(n4152), .Z(n4155) );
  XOR U4665 ( .A(n4154), .B(n4155), .Z(n3821) );
  XOR U4666 ( .A(n3821), .B(n3822), .Z(n3824) );
  XOR U4667 ( .A(n3823), .B(n3824), .Z(n4087) );
  OR U4668 ( .A(n3061), .B(n3060), .Z(n3065) );
  OR U4669 ( .A(n3063), .B(n3062), .Z(n3064) );
  AND U4670 ( .A(n3065), .B(n3064), .Z(n4255) );
  OR U4671 ( .A(n3071), .B(n3070), .Z(n3075) );
  OR U4672 ( .A(n3073), .B(n3072), .Z(n3074) );
  AND U4673 ( .A(n3075), .B(n3074), .Z(n4254) );
  XNOR U4674 ( .A(n4253), .B(n4254), .Z(n4256) );
  XNOR U4675 ( .A(n4255), .B(n4256), .Z(n3978) );
  NANDN U4676 ( .A(n3077), .B(n3076), .Z(n3081) );
  OR U4677 ( .A(n3079), .B(n3078), .Z(n3080) );
  NAND U4678 ( .A(n3081), .B(n3080), .Z(n3976) );
  OR U4679 ( .A(n3087), .B(n3086), .Z(n3091) );
  OR U4680 ( .A(n3089), .B(n3088), .Z(n3090) );
  AND U4681 ( .A(n3091), .B(n3090), .Z(n4259) );
  OR U4682 ( .A(n3093), .B(n3092), .Z(n3097) );
  OR U4683 ( .A(n3095), .B(n3094), .Z(n3096) );
  AND U4684 ( .A(n3097), .B(n3096), .Z(n4260) );
  XNOR U4685 ( .A(n4259), .B(n4260), .Z(n4262) );
  XNOR U4686 ( .A(n4261), .B(n4262), .Z(n3977) );
  XNOR U4687 ( .A(n3976), .B(n3977), .Z(n3979) );
  XNOR U4688 ( .A(n3978), .B(n3979), .Z(n4088) );
  XNOR U4689 ( .A(n4087), .B(n4088), .Z(n4090) );
  XOR U4690 ( .A(n4223), .B(n4224), .Z(n4226) );
  XNOR U4691 ( .A(n4225), .B(n4226), .Z(n3941) );
  OR U4692 ( .A(n3115), .B(n3114), .Z(n3119) );
  OR U4693 ( .A(n3117), .B(n3116), .Z(n3118) );
  NAND U4694 ( .A(n3119), .B(n3118), .Z(n3957) );
  OR U4695 ( .A(n3121), .B(n3120), .Z(n3125) );
  OR U4696 ( .A(n3123), .B(n3122), .Z(n3124) );
  AND U4697 ( .A(n3125), .B(n3124), .Z(n3955) );
  XOR U4698 ( .A(n3955), .B(n3956), .Z(n3958) );
  XOR U4699 ( .A(n3957), .B(n3958), .Z(n3942) );
  XOR U4700 ( .A(n3941), .B(n3942), .Z(n3944) );
  XOR U4701 ( .A(n3943), .B(n3944), .Z(n4089) );
  XOR U4702 ( .A(n4090), .B(n4089), .Z(n4031) );
  NANDN U4703 ( .A(n3131), .B(n3130), .Z(n3135) );
  NAND U4704 ( .A(n3133), .B(n3132), .Z(n3134) );
  AND U4705 ( .A(n3135), .B(n3134), .Z(n4029) );
  OR U4706 ( .A(n3137), .B(n3136), .Z(n3141) );
  NANDN U4707 ( .A(n3139), .B(n3138), .Z(n3140) );
  AND U4708 ( .A(n3141), .B(n3140), .Z(n3813) );
  OR U4709 ( .A(n3147), .B(n3146), .Z(n3151) );
  NANDN U4710 ( .A(n3149), .B(n3148), .Z(n3150) );
  NAND U4711 ( .A(n3151), .B(n3150), .Z(n3811) );
  XNOR U4712 ( .A(n3812), .B(n3811), .Z(n3814) );
  XNOR U4713 ( .A(n3813), .B(n3814), .Z(n3985) );
  IV U4714 ( .A(n3156), .Z(n3157) );
  NANDN U4715 ( .A(n3158), .B(n3157), .Z(n3162) );
  NAND U4716 ( .A(n3160), .B(n3159), .Z(n3161) );
  NAND U4717 ( .A(n3162), .B(n3161), .Z(n3850) );
  XNOR U4718 ( .A(n3849), .B(n3850), .Z(n3852) );
  XNOR U4719 ( .A(n3852), .B(n3851), .Z(n3983) );
  XNOR U4720 ( .A(n3983), .B(n3982), .Z(n3984) );
  XOR U4721 ( .A(n3985), .B(n3984), .Z(n4028) );
  XOR U4722 ( .A(n4029), .B(n4028), .Z(n4030) );
  XNOR U4723 ( .A(n4031), .B(n4030), .Z(n4122) );
  XOR U4724 ( .A(n4121), .B(n4122), .Z(n4110) );
  NANDN U4725 ( .A(n3176), .B(n3175), .Z(n3180) );
  NANDN U4726 ( .A(n3178), .B(n3177), .Z(n3179) );
  AND U4727 ( .A(n3180), .B(n3179), .Z(n4273) );
  XNOR U4728 ( .A(n4271), .B(n4272), .Z(n4274) );
  XNOR U4729 ( .A(n4273), .B(n4274), .Z(n4075) );
  XOR U4730 ( .A(n4076), .B(n4075), .Z(n4078) );
  OR U4731 ( .A(n3194), .B(n3193), .Z(n3198) );
  NANDN U4732 ( .A(n3196), .B(n3195), .Z(n3197) );
  AND U4733 ( .A(n3198), .B(n3197), .Z(n4134) );
  XNOR U4734 ( .A(n4134), .B(n4135), .Z(n4136) );
  XOR U4735 ( .A(n4137), .B(n4136), .Z(n4077) );
  XOR U4736 ( .A(n4078), .B(n4077), .Z(n4109) );
  XOR U4737 ( .A(n4110), .B(n4109), .Z(n4112) );
  NAND U4738 ( .A(n3204), .B(n3203), .Z(n3208) );
  NANDN U4739 ( .A(n3206), .B(n3205), .Z(n3207) );
  NAND U4740 ( .A(n3208), .B(n3207), .Z(n4126) );
  NANDN U4741 ( .A(n3210), .B(n3209), .Z(n3214) );
  OR U4742 ( .A(n3212), .B(n3211), .Z(n3213) );
  AND U4743 ( .A(n3214), .B(n3213), .Z(n4123) );
  OR U4744 ( .A(n3216), .B(n3215), .Z(n3220) );
  NAND U4745 ( .A(n3218), .B(n3217), .Z(n3219) );
  NAND U4746 ( .A(n3220), .B(n3219), .Z(n4124) );
  XNOR U4747 ( .A(n4123), .B(n4124), .Z(n4125) );
  XOR U4748 ( .A(n4126), .B(n4125), .Z(n4111) );
  XOR U4749 ( .A(n4112), .B(n4111), .Z(n4129) );
  NAND U4750 ( .A(n3222), .B(n3221), .Z(n3226) );
  OR U4751 ( .A(n3224), .B(n3223), .Z(n3225) );
  NAND U4752 ( .A(n3226), .B(n3225), .Z(n4127) );
  NANDN U4753 ( .A(n3228), .B(n3227), .Z(n3232) );
  NAND U4754 ( .A(n3230), .B(n3229), .Z(n3231) );
  NAND U4755 ( .A(n3232), .B(n3231), .Z(n3968) );
  NANDN U4756 ( .A(n3234), .B(n3233), .Z(n3238) );
  NAND U4757 ( .A(n3236), .B(n3235), .Z(n3237) );
  AND U4758 ( .A(n3238), .B(n3237), .Z(n3966) );
  XOR U4759 ( .A(n3966), .B(n3967), .Z(n3969) );
  XOR U4760 ( .A(n3968), .B(n3969), .Z(n3857) );
  OR U4761 ( .A(n3244), .B(n3243), .Z(n3248) );
  NANDN U4762 ( .A(n3246), .B(n3245), .Z(n3247) );
  NAND U4763 ( .A(n3248), .B(n3247), .Z(n3995) );
  OR U4764 ( .A(n3250), .B(n3249), .Z(n3254) );
  NANDN U4765 ( .A(n3252), .B(n3251), .Z(n3253) );
  AND U4766 ( .A(n3254), .B(n3253), .Z(n3992) );
  OR U4767 ( .A(n3256), .B(n3255), .Z(n3260) );
  NANDN U4768 ( .A(n3258), .B(n3257), .Z(n3259) );
  NAND U4769 ( .A(n3260), .B(n3259), .Z(n3993) );
  XOR U4770 ( .A(n3992), .B(n3993), .Z(n3994) );
  XOR U4771 ( .A(n3995), .B(n3994), .Z(n3856) );
  NANDN U4772 ( .A(n3262), .B(n3261), .Z(n3266) );
  NANDN U4773 ( .A(n3264), .B(n3263), .Z(n3265) );
  NAND U4774 ( .A(n3266), .B(n3265), .Z(n3894) );
  OR U4775 ( .A(n3268), .B(n3267), .Z(n3272) );
  NAND U4776 ( .A(n3270), .B(n3269), .Z(n3271) );
  NAND U4777 ( .A(n3272), .B(n3271), .Z(n3893) );
  XOR U4778 ( .A(n3894), .B(n3893), .Z(n3896) );
  NANDN U4779 ( .A(n3274), .B(n3273), .Z(n3278) );
  NANDN U4780 ( .A(n3276), .B(n3275), .Z(n3277) );
  NAND U4781 ( .A(n3278), .B(n3277), .Z(n3895) );
  XOR U4782 ( .A(n3896), .B(n3895), .Z(n3855) );
  XOR U4783 ( .A(n3856), .B(n3855), .Z(n3858) );
  XOR U4784 ( .A(n3857), .B(n3858), .Z(n3803) );
  NANDN U4785 ( .A(n3280), .B(n3279), .Z(n3284) );
  NAND U4786 ( .A(n3282), .B(n3281), .Z(n3283) );
  AND U4787 ( .A(n3284), .B(n3283), .Z(n3989) );
  XNOR U4788 ( .A(n3986), .B(n3987), .Z(n3988) );
  XNOR U4789 ( .A(n3989), .B(n3988), .Z(n4283) );
  NANDN U4790 ( .A(n3294), .B(n3293), .Z(n3298) );
  NANDN U4791 ( .A(n3296), .B(n3295), .Z(n3297) );
  NAND U4792 ( .A(n3298), .B(n3297), .Z(n3868) );
  NANDN U4793 ( .A(n3300), .B(n3299), .Z(n3304) );
  NAND U4794 ( .A(n3302), .B(n3301), .Z(n3303) );
  AND U4795 ( .A(n3304), .B(n3303), .Z(n3865) );
  NANDN U4796 ( .A(n3306), .B(n3305), .Z(n3310) );
  OR U4797 ( .A(n3308), .B(n3307), .Z(n3309) );
  AND U4798 ( .A(n3310), .B(n3309), .Z(n3866) );
  XOR U4799 ( .A(n3865), .B(n3866), .Z(n3867) );
  XNOR U4800 ( .A(n3868), .B(n3867), .Z(n4281) );
  NANDN U4801 ( .A(n3312), .B(n3311), .Z(n3316) );
  NAND U4802 ( .A(n3314), .B(n3313), .Z(n3315) );
  NAND U4803 ( .A(n3316), .B(n3315), .Z(n3861) );
  NANDN U4804 ( .A(n3318), .B(n3317), .Z(n3322) );
  OR U4805 ( .A(n3320), .B(n3319), .Z(n3321) );
  AND U4806 ( .A(n3322), .B(n3321), .Z(n3860) );
  NANDN U4807 ( .A(n3324), .B(n3323), .Z(n3328) );
  NAND U4808 ( .A(n3326), .B(n3325), .Z(n3327) );
  NAND U4809 ( .A(n3328), .B(n3327), .Z(n3859) );
  XNOR U4810 ( .A(n3860), .B(n3859), .Z(n3862) );
  XOR U4811 ( .A(n3861), .B(n3862), .Z(n4282) );
  XOR U4812 ( .A(n4281), .B(n4282), .Z(n4284) );
  XOR U4813 ( .A(n4283), .B(n4284), .Z(n3802) );
  NANDN U4814 ( .A(n3330), .B(n3329), .Z(n3334) );
  NANDN U4815 ( .A(n3332), .B(n3331), .Z(n3333) );
  NAND U4816 ( .A(n3334), .B(n3333), .Z(n4044) );
  NANDN U4817 ( .A(n3336), .B(n3335), .Z(n3340) );
  NANDN U4818 ( .A(n3338), .B(n3337), .Z(n3339) );
  NAND U4819 ( .A(n3340), .B(n3339), .Z(n4042) );
  OR U4820 ( .A(n3342), .B(n3341), .Z(n3346) );
  OR U4821 ( .A(n3344), .B(n3343), .Z(n3345) );
  AND U4822 ( .A(n3346), .B(n3345), .Z(n4144) );
  OR U4823 ( .A(n3348), .B(n3347), .Z(n3352) );
  OR U4824 ( .A(n3350), .B(n3349), .Z(n3351) );
  AND U4825 ( .A(n3352), .B(n3351), .Z(n4145) );
  XOR U4826 ( .A(n4144), .B(n4145), .Z(n4147) );
  NANDN U4827 ( .A(n3354), .B(n3353), .Z(n3358) );
  NAND U4828 ( .A(n3356), .B(n3355), .Z(n3357) );
  AND U4829 ( .A(n3358), .B(n3357), .Z(n4146) );
  XOR U4830 ( .A(n4147), .B(n4146), .Z(n4174) );
  NANDN U4831 ( .A(n3360), .B(n3359), .Z(n3364) );
  NAND U4832 ( .A(n3362), .B(n3361), .Z(n3363) );
  NAND U4833 ( .A(n3364), .B(n3363), .Z(n3962) );
  OR U4834 ( .A(n3366), .B(n3365), .Z(n3370) );
  OR U4835 ( .A(n3368), .B(n3367), .Z(n3369) );
  AND U4836 ( .A(n3370), .B(n3369), .Z(n3959) );
  NANDN U4837 ( .A(n3372), .B(n3371), .Z(n3376) );
  NANDN U4838 ( .A(n3374), .B(n3373), .Z(n3375) );
  AND U4839 ( .A(n3376), .B(n3375), .Z(n3961) );
  XOR U4840 ( .A(n3959), .B(n3961), .Z(n3963) );
  XOR U4841 ( .A(n3962), .B(n3963), .Z(n4172) );
  NANDN U4842 ( .A(n3378), .B(n3377), .Z(n3382) );
  NAND U4843 ( .A(n3380), .B(n3379), .Z(n3381) );
  AND U4844 ( .A(n3382), .B(n3381), .Z(n4173) );
  XNOR U4845 ( .A(n4172), .B(n4173), .Z(n4175) );
  XNOR U4846 ( .A(n4174), .B(n4175), .Z(n4040) );
  XOR U4847 ( .A(n4042), .B(n4040), .Z(n4043) );
  XNOR U4848 ( .A(n4044), .B(n4043), .Z(n3801) );
  XNOR U4849 ( .A(n3802), .B(n3801), .Z(n3804) );
  XOR U4850 ( .A(n3803), .B(n3804), .Z(n4104) );
  NAND U4851 ( .A(n3384), .B(n3383), .Z(n3388) );
  NAND U4852 ( .A(n3386), .B(n3385), .Z(n3387) );
  AND U4853 ( .A(n3388), .B(n3387), .Z(n3998) );
  OR U4854 ( .A(n3394), .B(n3393), .Z(n3398) );
  NANDN U4855 ( .A(n3396), .B(n3395), .Z(n3397) );
  NAND U4856 ( .A(n3398), .B(n3397), .Z(n3997) );
  XNOR U4857 ( .A(n3996), .B(n3997), .Z(n3999) );
  XNOR U4858 ( .A(n3998), .B(n3999), .Z(n4064) );
  NANDN U4859 ( .A(n3400), .B(n3399), .Z(n3404) );
  NANDN U4860 ( .A(n3402), .B(n3401), .Z(n3403) );
  AND U4861 ( .A(n3404), .B(n3403), .Z(n3883) );
  NANDN U4862 ( .A(n3406), .B(n3405), .Z(n3410) );
  OR U4863 ( .A(n3408), .B(n3407), .Z(n3409) );
  AND U4864 ( .A(n3410), .B(n3409), .Z(n3881) );
  XNOR U4865 ( .A(n3881), .B(n3882), .Z(n3884) );
  XNOR U4866 ( .A(n3883), .B(n3884), .Z(n4063) );
  XOR U4867 ( .A(n4064), .B(n4063), .Z(n4065) );
  NANDN U4868 ( .A(n3420), .B(n3419), .Z(n3424) );
  NANDN U4869 ( .A(n3422), .B(n3421), .Z(n3423) );
  AND U4870 ( .A(n3424), .B(n3423), .Z(n3875) );
  OR U4871 ( .A(n3426), .B(n3425), .Z(n3430) );
  NANDN U4872 ( .A(n3428), .B(n3427), .Z(n3429) );
  AND U4873 ( .A(n3430), .B(n3429), .Z(n3876) );
  XNOR U4874 ( .A(n3875), .B(n3876), .Z(n3878) );
  XNOR U4875 ( .A(n3877), .B(n3878), .Z(n4066) );
  XOR U4876 ( .A(n4065), .B(n4066), .Z(n4020) );
  NANDN U4877 ( .A(n3432), .B(n3431), .Z(n3436) );
  NANDN U4878 ( .A(n3434), .B(n3433), .Z(n3435) );
  AND U4879 ( .A(n3436), .B(n3435), .Z(n4166) );
  OR U4880 ( .A(n3438), .B(n3437), .Z(n3442) );
  NANDN U4881 ( .A(n3440), .B(n3439), .Z(n3441) );
  AND U4882 ( .A(n3442), .B(n3441), .Z(n3899) );
  NANDN U4883 ( .A(n3448), .B(n3447), .Z(n3452) );
  NAND U4884 ( .A(n3450), .B(n3449), .Z(n3451) );
  AND U4885 ( .A(n3452), .B(n3451), .Z(n3898) );
  XNOR U4886 ( .A(n3897), .B(n3898), .Z(n3900) );
  XNOR U4887 ( .A(n3899), .B(n3900), .Z(n4167) );
  XNOR U4888 ( .A(n4166), .B(n4167), .Z(n4169) );
  NANDN U4889 ( .A(n3454), .B(n3453), .Z(n3458) );
  OR U4890 ( .A(n3456), .B(n3455), .Z(n3457) );
  NAND U4891 ( .A(n3458), .B(n3457), .Z(n4165) );
  NANDN U4892 ( .A(n3460), .B(n3459), .Z(n3464) );
  NAND U4893 ( .A(n3462), .B(n3461), .Z(n3463) );
  AND U4894 ( .A(n3464), .B(n3463), .Z(n4162) );
  NANDN U4895 ( .A(n3466), .B(n3465), .Z(n3470) );
  NAND U4896 ( .A(n3468), .B(n3467), .Z(n3469) );
  AND U4897 ( .A(n3470), .B(n3469), .Z(n4163) );
  XOR U4898 ( .A(n4162), .B(n4163), .Z(n4164) );
  XNOR U4899 ( .A(n4165), .B(n4164), .Z(n4168) );
  XNOR U4900 ( .A(n4169), .B(n4168), .Z(n4019) );
  NANDN U4901 ( .A(n3472), .B(n3471), .Z(n3476) );
  NAND U4902 ( .A(n3474), .B(n3473), .Z(n3475) );
  AND U4903 ( .A(n3476), .B(n3475), .Z(n3939) );
  NANDN U4904 ( .A(n3478), .B(n3477), .Z(n3482) );
  NAND U4905 ( .A(n3480), .B(n3479), .Z(n3481) );
  AND U4906 ( .A(n3482), .B(n3481), .Z(n4014) );
  NANDN U4907 ( .A(n3484), .B(n3483), .Z(n3488) );
  NAND U4908 ( .A(n3486), .B(n3485), .Z(n3487) );
  AND U4909 ( .A(n3488), .B(n3487), .Z(n4012) );
  NANDN U4910 ( .A(n3490), .B(n3489), .Z(n3494) );
  OR U4911 ( .A(n3492), .B(n3491), .Z(n3493) );
  AND U4912 ( .A(n3494), .B(n3493), .Z(n4013) );
  XNOR U4913 ( .A(n4012), .B(n4013), .Z(n4015) );
  XNOR U4914 ( .A(n4014), .B(n4015), .Z(n3937) );
  XOR U4915 ( .A(n3937), .B(n3938), .Z(n3940) );
  XOR U4916 ( .A(n3939), .B(n3940), .Z(n4018) );
  XNOR U4917 ( .A(n4019), .B(n4018), .Z(n4021) );
  XNOR U4918 ( .A(n4020), .B(n4021), .Z(n4103) );
  XOR U4919 ( .A(n4104), .B(n4103), .Z(n4106) );
  NANDN U4920 ( .A(n3500), .B(n3499), .Z(n3504) );
  NAND U4921 ( .A(n3502), .B(n3501), .Z(n3503) );
  NAND U4922 ( .A(n3504), .B(n3503), .Z(n4050) );
  OR U4923 ( .A(n3506), .B(n3505), .Z(n3510) );
  OR U4924 ( .A(n3508), .B(n3507), .Z(n3509) );
  AND U4925 ( .A(n3510), .B(n3509), .Z(n4047) );
  NANDN U4926 ( .A(n3512), .B(n3511), .Z(n3516) );
  NAND U4927 ( .A(n3514), .B(n3513), .Z(n3515) );
  NAND U4928 ( .A(n3516), .B(n3515), .Z(n4048) );
  XNOR U4929 ( .A(n4047), .B(n4048), .Z(n4049) );
  XOR U4930 ( .A(n4050), .B(n4049), .Z(n3807) );
  OR U4931 ( .A(n3522), .B(n3521), .Z(n3526) );
  OR U4932 ( .A(n3524), .B(n3523), .Z(n3525) );
  AND U4933 ( .A(n3526), .B(n3525), .Z(n4197) );
  NANDN U4934 ( .A(n3528), .B(n3527), .Z(n3532) );
  NAND U4935 ( .A(n3530), .B(n3529), .Z(n3531) );
  NAND U4936 ( .A(n3532), .B(n3531), .Z(n4196) );
  XNOR U4937 ( .A(oglobal[2]), .B(n4196), .Z(n4198) );
  XNOR U4938 ( .A(n4197), .B(n4198), .Z(n3948) );
  XOR U4939 ( .A(n3947), .B(n3948), .Z(n3949) );
  OR U4940 ( .A(n3534), .B(n3533), .Z(n3538) );
  OR U4941 ( .A(n3536), .B(n3535), .Z(n3537) );
  AND U4942 ( .A(n3538), .B(n3537), .Z(n4203) );
  NANDN U4943 ( .A(n3543), .B(oglobal[1]), .Z(n3547) );
  OR U4944 ( .A(n3545), .B(n3544), .Z(n3546) );
  NAND U4945 ( .A(n3547), .B(n3546), .Z(n4202) );
  XNOR U4946 ( .A(n4201), .B(n4202), .Z(n4204) );
  XNOR U4947 ( .A(n4203), .B(n4204), .Z(n3950) );
  XNOR U4948 ( .A(n3949), .B(n3950), .Z(n4083) );
  XOR U4949 ( .A(n4083), .B(n4084), .Z(n4085) );
  NANDN U4950 ( .A(n3553), .B(n3552), .Z(n3557) );
  OR U4951 ( .A(n3555), .B(n3554), .Z(n3556) );
  AND U4952 ( .A(n3557), .B(n3556), .Z(n3845) );
  OR U4953 ( .A(n3563), .B(n3562), .Z(n3567) );
  OR U4954 ( .A(n3565), .B(n3564), .Z(n3566) );
  AND U4955 ( .A(n3567), .B(n3566), .Z(n3844) );
  XNOR U4956 ( .A(n3843), .B(n3844), .Z(n3846) );
  XNOR U4957 ( .A(n3845), .B(n3846), .Z(n3972) );
  NANDN U4958 ( .A(n3569), .B(n3568), .Z(n3573) );
  NAND U4959 ( .A(n3571), .B(n3570), .Z(n3572) );
  AND U4960 ( .A(n3573), .B(n3572), .Z(n4184) );
  OR U4961 ( .A(n3575), .B(n3574), .Z(n3579) );
  OR U4962 ( .A(n3577), .B(n3576), .Z(n3578) );
  AND U4963 ( .A(n3579), .B(n3578), .Z(n4182) );
  OR U4964 ( .A(n3581), .B(n3580), .Z(n3585) );
  OR U4965 ( .A(n3583), .B(n3582), .Z(n3584) );
  AND U4966 ( .A(n3585), .B(n3584), .Z(n4183) );
  XNOR U4967 ( .A(n4182), .B(n4183), .Z(n4185) );
  XNOR U4968 ( .A(n4184), .B(n4185), .Z(n3970) );
  NAND U4969 ( .A(n3587), .B(n3586), .Z(n3591) );
  NAND U4970 ( .A(n3589), .B(n3588), .Z(n3590) );
  AND U4971 ( .A(n3591), .B(n3590), .Z(n3971) );
  XOR U4972 ( .A(n3970), .B(n3971), .Z(n3973) );
  XOR U4973 ( .A(n3972), .B(n3973), .Z(n4086) );
  XNOR U4974 ( .A(n4085), .B(n4086), .Z(n3808) );
  XOR U4975 ( .A(n3807), .B(n3808), .Z(n3810) );
  NANDN U4976 ( .A(n3593), .B(n3592), .Z(n3597) );
  NANDN U4977 ( .A(n3595), .B(n3594), .Z(n3596) );
  NAND U4978 ( .A(n3597), .B(n3596), .Z(n3905) );
  NANDN U4979 ( .A(n3599), .B(n3598), .Z(n3603) );
  OR U4980 ( .A(n3601), .B(n3600), .Z(n3602) );
  AND U4981 ( .A(n3603), .B(n3602), .Z(n3903) );
  OR U4982 ( .A(n3605), .B(n3604), .Z(n3609) );
  OR U4983 ( .A(n3607), .B(n3606), .Z(n3608) );
  NAND U4984 ( .A(n3609), .B(n3608), .Z(n3904) );
  XOR U4985 ( .A(n3903), .B(n3904), .Z(n3906) );
  XOR U4986 ( .A(n3905), .B(n3906), .Z(n3820) );
  OR U4987 ( .A(n3611), .B(n3610), .Z(n3615) );
  NANDN U4988 ( .A(n3613), .B(n3612), .Z(n3614) );
  AND U4989 ( .A(n3615), .B(n3614), .Z(n3817) );
  NANDN U4990 ( .A(n3617), .B(n3616), .Z(n3621) );
  NANDN U4991 ( .A(n3619), .B(n3618), .Z(n3620) );
  NAND U4992 ( .A(n3621), .B(n3620), .Z(n4215) );
  XNOR U4993 ( .A(n4214), .B(n4213), .Z(n4216) );
  XOR U4994 ( .A(n4215), .B(n4216), .Z(n3818) );
  XNOR U4995 ( .A(n3817), .B(n3818), .Z(n3819) );
  XNOR U4996 ( .A(n3820), .B(n3819), .Z(n4095) );
  NANDN U4997 ( .A(n3635), .B(n3634), .Z(n3639) );
  OR U4998 ( .A(n3637), .B(n3636), .Z(n3638) );
  AND U4999 ( .A(n3639), .B(n3638), .Z(n4265) );
  NANDN U5000 ( .A(n3641), .B(n3640), .Z(n3645) );
  OR U5001 ( .A(n3643), .B(n3642), .Z(n3644) );
  AND U5002 ( .A(n3645), .B(n3644), .Z(n4266) );
  XNOR U5003 ( .A(n4265), .B(n4266), .Z(n4267) );
  XNOR U5004 ( .A(n4268), .B(n4267), .Z(n4160) );
  NANDN U5005 ( .A(n3647), .B(n3646), .Z(n3651) );
  NANDN U5006 ( .A(n3649), .B(n3648), .Z(n3650) );
  AND U5007 ( .A(n3651), .B(n3650), .Z(n3936) );
  NANDN U5008 ( .A(n3653), .B(n3652), .Z(n3657) );
  NANDN U5009 ( .A(n3655), .B(n3654), .Z(n3656) );
  AND U5010 ( .A(n3657), .B(n3656), .Z(n3933) );
  NANDN U5011 ( .A(n3659), .B(n3658), .Z(n3663) );
  NANDN U5012 ( .A(n3661), .B(n3660), .Z(n3662) );
  AND U5013 ( .A(n3663), .B(n3662), .Z(n3934) );
  XNOR U5014 ( .A(n3933), .B(n3934), .Z(n3935) );
  XOR U5015 ( .A(n3936), .B(n3935), .Z(n4158) );
  NANDN U5016 ( .A(n3665), .B(n3664), .Z(n3669) );
  NANDN U5017 ( .A(n3667), .B(n3666), .Z(n3668) );
  AND U5018 ( .A(n3669), .B(n3668), .Z(n4159) );
  XOR U5019 ( .A(n4158), .B(n4159), .Z(n4161) );
  XOR U5020 ( .A(n4160), .B(n4161), .Z(n4093) );
  NANDN U5021 ( .A(n3671), .B(n3670), .Z(n3675) );
  NANDN U5022 ( .A(n3673), .B(n3672), .Z(n3674) );
  NAND U5023 ( .A(n3675), .B(n3674), .Z(n4094) );
  XNOR U5024 ( .A(n4093), .B(n4094), .Z(n4096) );
  XOR U5025 ( .A(n4095), .B(n4096), .Z(n3809) );
  XOR U5026 ( .A(n3810), .B(n3809), .Z(n4105) );
  XNOR U5027 ( .A(n4106), .B(n4105), .Z(n4293) );
  OR U5028 ( .A(n3677), .B(n3676), .Z(n3681) );
  NANDN U5029 ( .A(n3679), .B(n3678), .Z(n3680) );
  AND U5030 ( .A(n3681), .B(n3680), .Z(n4292) );
  NANDN U5031 ( .A(n3683), .B(n3682), .Z(n3687) );
  OR U5032 ( .A(n3685), .B(n3684), .Z(n3686) );
  NAND U5033 ( .A(n3687), .B(n3686), .Z(n4141) );
  NANDN U5034 ( .A(n3689), .B(n3688), .Z(n3693) );
  NANDN U5035 ( .A(n3691), .B(n3690), .Z(n3692) );
  AND U5036 ( .A(n3693), .B(n3692), .Z(n4138) );
  NAND U5037 ( .A(n3699), .B(n3698), .Z(n3703) );
  NANDN U5038 ( .A(n3701), .B(n3700), .Z(n3702) );
  NAND U5039 ( .A(n3703), .B(n3702), .Z(n4286) );
  NANDN U5040 ( .A(n3705), .B(n3704), .Z(n3709) );
  NANDN U5041 ( .A(n3707), .B(n3706), .Z(n3708) );
  NAND U5042 ( .A(n3709), .B(n3708), .Z(n4285) );
  XNOR U5043 ( .A(n4286), .B(n4285), .Z(n4288) );
  XNOR U5044 ( .A(n4287), .B(n4288), .Z(n4139) );
  XNOR U5045 ( .A(n4138), .B(n4139), .Z(n4140) );
  XOR U5046 ( .A(n4141), .B(n4140), .Z(n4115) );
  OR U5047 ( .A(n3711), .B(n3710), .Z(n3715) );
  NANDN U5048 ( .A(n3713), .B(n3712), .Z(n3714) );
  NAND U5049 ( .A(n3715), .B(n3714), .Z(n4280) );
  OR U5050 ( .A(n3717), .B(n3716), .Z(n3721) );
  NAND U5051 ( .A(n3719), .B(n3718), .Z(n3720) );
  AND U5052 ( .A(n3721), .B(n3720), .Z(n4277) );
  NAND U5053 ( .A(n3723), .B(n3722), .Z(n3727) );
  NANDN U5054 ( .A(n3725), .B(n3724), .Z(n3726) );
  NAND U5055 ( .A(n3727), .B(n3726), .Z(n4278) );
  XNOR U5056 ( .A(n4277), .B(n4278), .Z(n4279) );
  XOR U5057 ( .A(n4280), .B(n4279), .Z(n4102) );
  NAND U5058 ( .A(n3737), .B(n3736), .Z(n3741) );
  NANDN U5059 ( .A(n3739), .B(n3738), .Z(n3740) );
  NAND U5060 ( .A(n3741), .B(n3740), .Z(n4068) );
  XNOR U5061 ( .A(n4067), .B(n4068), .Z(n4069) );
  XOR U5062 ( .A(n4070), .B(n4069), .Z(n4099) );
  OR U5063 ( .A(n3743), .B(n3742), .Z(n3747) );
  NAND U5064 ( .A(n3745), .B(n3744), .Z(n3746) );
  NAND U5065 ( .A(n3747), .B(n3746), .Z(n4100) );
  XOR U5066 ( .A(n4099), .B(n4100), .Z(n4101) );
  XOR U5067 ( .A(n4102), .B(n4101), .Z(n4116) );
  XOR U5068 ( .A(n4115), .B(n4116), .Z(n4117) );
  OR U5069 ( .A(n3753), .B(n3752), .Z(n3757) );
  NANDN U5070 ( .A(n3755), .B(n3754), .Z(n3756) );
  AND U5071 ( .A(n3757), .B(n3756), .Z(n4071) );
  OR U5072 ( .A(n3759), .B(n3758), .Z(n3763) );
  OR U5073 ( .A(n3761), .B(n3760), .Z(n3762) );
  AND U5074 ( .A(n3763), .B(n3762), .Z(n4072) );
  XNOR U5075 ( .A(n4071), .B(n4072), .Z(n4073) );
  XOR U5076 ( .A(n4074), .B(n4073), .Z(n4081) );
  NANDN U5077 ( .A(n3765), .B(n3764), .Z(n3769) );
  NANDN U5078 ( .A(n3767), .B(n3766), .Z(n3768) );
  AND U5079 ( .A(n3769), .B(n3768), .Z(n4057) );
  OR U5080 ( .A(n3771), .B(n3770), .Z(n3775) );
  NAND U5081 ( .A(n3773), .B(n3772), .Z(n3774) );
  NAND U5082 ( .A(n3775), .B(n3774), .Z(n4058) );
  XNOR U5083 ( .A(n4057), .B(n4058), .Z(n4060) );
  NANDN U5084 ( .A(n3777), .B(n3776), .Z(n3781) );
  NAND U5085 ( .A(n3779), .B(n3778), .Z(n3780) );
  NAND U5086 ( .A(n3781), .B(n3780), .Z(n4059) );
  XNOR U5087 ( .A(n4060), .B(n4059), .Z(n4080) );
  NANDN U5088 ( .A(n3783), .B(n3782), .Z(n3787) );
  NAND U5089 ( .A(n3785), .B(n3784), .Z(n3786) );
  NAND U5090 ( .A(n3787), .B(n3786), .Z(n4079) );
  XNOR U5091 ( .A(n4080), .B(n4079), .Z(n4082) );
  XOR U5092 ( .A(n4081), .B(n4082), .Z(n4118) );
  XOR U5093 ( .A(n4117), .B(n4118), .Z(n4291) );
  XOR U5094 ( .A(n4292), .B(n4291), .Z(n4294) );
  XOR U5095 ( .A(n4293), .B(n4294), .Z(n4133) );
  NANDN U5096 ( .A(n3789), .B(n3788), .Z(n3793) );
  NANDN U5097 ( .A(n3791), .B(n3790), .Z(n3792) );
  AND U5098 ( .A(n3793), .B(n3792), .Z(n4130) );
  NANDN U5099 ( .A(n3795), .B(n3794), .Z(n3799) );
  NANDN U5100 ( .A(n3797), .B(n3796), .Z(n3798) );
  AND U5101 ( .A(n3799), .B(n3798), .Z(n4131) );
  XNOR U5102 ( .A(n4130), .B(n4131), .Z(n4132) );
  XOR U5103 ( .A(n4133), .B(n4132), .Z(n4128) );
  XOR U5104 ( .A(n4127), .B(n4128), .Z(n3800) );
  XNOR U5105 ( .A(n4129), .B(n3800), .Z(o[2]) );
  NANDN U5106 ( .A(n3802), .B(n3801), .Z(n3806) );
  NAND U5107 ( .A(n3804), .B(n3803), .Z(n3805) );
  NAND U5108 ( .A(n3806), .B(n3805), .Z(n4489) );
  OR U5109 ( .A(n3812), .B(n3811), .Z(n3816) );
  OR U5110 ( .A(n3814), .B(n3813), .Z(n3815) );
  AND U5111 ( .A(n3816), .B(n3815), .Z(n4541) );
  XOR U5112 ( .A(n4541), .B(n4542), .Z(n4543) );
  OR U5113 ( .A(n3822), .B(n3821), .Z(n3826) );
  NAND U5114 ( .A(n3824), .B(n3823), .Z(n3825) );
  NAND U5115 ( .A(n3826), .B(n3825), .Z(n4544) );
  XOR U5116 ( .A(n4543), .B(n4544), .Z(n4529) );
  OR U5117 ( .A(n3828), .B(n3827), .Z(n3832) );
  NANDN U5118 ( .A(n3830), .B(n3829), .Z(n3831) );
  AND U5119 ( .A(n3832), .B(n3831), .Z(n4504) );
  OR U5120 ( .A(n3838), .B(n3837), .Z(n3842) );
  OR U5121 ( .A(n3840), .B(n3839), .Z(n3841) );
  NAND U5122 ( .A(n3842), .B(n3841), .Z(n4335) );
  XOR U5123 ( .A(n4336), .B(n4335), .Z(n4338) );
  OR U5124 ( .A(n3844), .B(n3843), .Z(n3848) );
  OR U5125 ( .A(n3846), .B(n3845), .Z(n3847) );
  NAND U5126 ( .A(n3848), .B(n3847), .Z(n4337) );
  XOR U5127 ( .A(n4338), .B(n4337), .Z(n4503) );
  OR U5128 ( .A(n3850), .B(n3849), .Z(n3854) );
  OR U5129 ( .A(n3852), .B(n3851), .Z(n3853) );
  AND U5130 ( .A(n3854), .B(n3853), .Z(n4502) );
  XNOR U5131 ( .A(n4503), .B(n4502), .Z(n4505) );
  XNOR U5132 ( .A(n4504), .B(n4505), .Z(n4527) );
  XOR U5133 ( .A(n4527), .B(n4528), .Z(n4530) );
  XOR U5134 ( .A(n4529), .B(n4530), .Z(n4487) );
  XNOR U5135 ( .A(n4486), .B(n4487), .Z(n4488) );
  XNOR U5136 ( .A(n4489), .B(n4488), .Z(n4462) );
  NANDN U5137 ( .A(n3860), .B(n3859), .Z(n3864) );
  NAND U5138 ( .A(n3862), .B(n3861), .Z(n3863) );
  NAND U5139 ( .A(n3864), .B(n3863), .Z(n4413) );
  XNOR U5140 ( .A(n4413), .B(n4412), .Z(n4415) );
  NANDN U5141 ( .A(n3870), .B(n3869), .Z(n3874) );
  NANDN U5142 ( .A(n3872), .B(n3871), .Z(n3873) );
  NAND U5143 ( .A(n3874), .B(n3873), .Z(n4540) );
  OR U5144 ( .A(n3876), .B(n3875), .Z(n3880) );
  OR U5145 ( .A(n3878), .B(n3877), .Z(n3879) );
  NAND U5146 ( .A(n3880), .B(n3879), .Z(n4538) );
  OR U5147 ( .A(n3882), .B(n3881), .Z(n3886) );
  OR U5148 ( .A(n3884), .B(n3883), .Z(n3885) );
  NAND U5149 ( .A(n3886), .B(n3885), .Z(n4537) );
  XNOR U5150 ( .A(n4538), .B(n4537), .Z(n4539) );
  XOR U5151 ( .A(n4540), .B(n4539), .Z(n4414) );
  XOR U5152 ( .A(n4415), .B(n4414), .Z(n4381) );
  OR U5153 ( .A(n3888), .B(n3887), .Z(n3892) );
  NANDN U5154 ( .A(n3890), .B(n3889), .Z(n3891) );
  AND U5155 ( .A(n3892), .B(n3891), .Z(n4509) );
  OR U5156 ( .A(n3898), .B(n3897), .Z(n3902) );
  OR U5157 ( .A(n3900), .B(n3899), .Z(n3901) );
  NAND U5158 ( .A(n3902), .B(n3901), .Z(n4507) );
  XNOR U5159 ( .A(n4506), .B(n4507), .Z(n4508) );
  XNOR U5160 ( .A(n4509), .B(n4508), .Z(n4379) );
  OR U5161 ( .A(n3908), .B(n3907), .Z(n3912) );
  NANDN U5162 ( .A(n3910), .B(n3909), .Z(n3911) );
  NAND U5163 ( .A(n3912), .B(n3911), .Z(n4343) );
  XOR U5164 ( .A(n4344), .B(n4343), .Z(n4346) );
  OR U5165 ( .A(n3914), .B(n3913), .Z(n3918) );
  OR U5166 ( .A(n3916), .B(n3915), .Z(n3917) );
  NAND U5167 ( .A(n3918), .B(n3917), .Z(n4345) );
  XOR U5168 ( .A(n4346), .B(n4345), .Z(n4535) );
  OR U5169 ( .A(n3928), .B(n3927), .Z(n3932) );
  NANDN U5170 ( .A(n3930), .B(n3929), .Z(n3931) );
  NAND U5171 ( .A(n3932), .B(n3931), .Z(n4325) );
  XNOR U5172 ( .A(n4326), .B(n4325), .Z(n4328) );
  XOR U5173 ( .A(n4327), .B(n4328), .Z(n4533) );
  XOR U5174 ( .A(n4533), .B(n4534), .Z(n4536) );
  XOR U5175 ( .A(n4535), .B(n4536), .Z(n4380) );
  XOR U5176 ( .A(n4379), .B(n4380), .Z(n4382) );
  XOR U5177 ( .A(n4381), .B(n4382), .Z(n4451) );
  NANDN U5178 ( .A(n3942), .B(n3941), .Z(n3946) );
  NANDN U5179 ( .A(n3944), .B(n3943), .Z(n3945) );
  NAND U5180 ( .A(n3946), .B(n3945), .Z(n4366) );
  XNOR U5181 ( .A(n4366), .B(n4365), .Z(n4368) );
  IV U5182 ( .A(n3959), .Z(n3960) );
  NANDN U5183 ( .A(n3961), .B(n3960), .Z(n3965) );
  NAND U5184 ( .A(n3963), .B(n3962), .Z(n3964) );
  NAND U5185 ( .A(n3965), .B(n3964), .Z(n4313) );
  XNOR U5186 ( .A(n4314), .B(n4313), .Z(n4315) );
  XNOR U5187 ( .A(n4316), .B(n4315), .Z(n4367) );
  XOR U5188 ( .A(n4368), .B(n4367), .Z(n4418) );
  XNOR U5189 ( .A(n4419), .B(n4418), .Z(n4421) );
  NANDN U5190 ( .A(n3971), .B(n3970), .Z(n3975) );
  NANDN U5191 ( .A(n3973), .B(n3972), .Z(n3974) );
  AND U5192 ( .A(n3975), .B(n3974), .Z(n4359) );
  NAND U5193 ( .A(n3977), .B(n3976), .Z(n3981) );
  NANDN U5194 ( .A(n3979), .B(n3978), .Z(n3980) );
  AND U5195 ( .A(n3981), .B(n3980), .Z(n4360) );
  XNOR U5196 ( .A(n4359), .B(n4360), .Z(n4362) );
  XNOR U5197 ( .A(n4361), .B(n4362), .Z(n4420) );
  XOR U5198 ( .A(n4421), .B(n4420), .Z(n4448) );
  OR U5199 ( .A(n3987), .B(n3986), .Z(n3991) );
  OR U5200 ( .A(n3989), .B(n3988), .Z(n3990) );
  NAND U5201 ( .A(n3991), .B(n3990), .Z(n4397) );
  OR U5202 ( .A(n3997), .B(n3996), .Z(n4001) );
  OR U5203 ( .A(n3999), .B(n3998), .Z(n4000) );
  NAND U5204 ( .A(n4001), .B(n4000), .Z(n4395) );
  XNOR U5205 ( .A(n4396), .B(n4395), .Z(n4398) );
  XOR U5206 ( .A(n4397), .B(n4398), .Z(n4499) );
  XNOR U5207 ( .A(n4498), .B(n4499), .Z(n4501) );
  OR U5208 ( .A(n4007), .B(n4006), .Z(n4011) );
  NANDN U5209 ( .A(n4009), .B(n4008), .Z(n4010) );
  AND U5210 ( .A(n4011), .B(n4010), .Z(n4309) );
  OR U5211 ( .A(n4013), .B(n4012), .Z(n4017) );
  OR U5212 ( .A(n4015), .B(n4014), .Z(n4016) );
  NAND U5213 ( .A(n4017), .B(n4016), .Z(n4310) );
  XOR U5214 ( .A(n4309), .B(n4310), .Z(n4312) );
  XOR U5215 ( .A(n4311), .B(n4312), .Z(n4500) );
  XOR U5216 ( .A(n4501), .B(n4500), .Z(n4449) );
  XOR U5217 ( .A(n4451), .B(n4450), .Z(n4461) );
  NAND U5218 ( .A(n4019), .B(n4018), .Z(n4023) );
  NANDN U5219 ( .A(n4021), .B(n4020), .Z(n4022) );
  AND U5220 ( .A(n4023), .B(n4022), .Z(n4447) );
  XNOR U5221 ( .A(n4444), .B(n4445), .Z(n4446) );
  XNOR U5222 ( .A(n4447), .B(n4446), .Z(n4460) );
  XOR U5223 ( .A(n4461), .B(n4460), .Z(n4463) );
  XOR U5224 ( .A(n4462), .B(n4463), .Z(n4456) );
  IV U5225 ( .A(n4040), .Z(n4041) );
  NANDN U5226 ( .A(n4042), .B(n4041), .Z(n4046) );
  NANDN U5227 ( .A(n4044), .B(n4043), .Z(n4045) );
  NAND U5228 ( .A(n4046), .B(n4045), .Z(n4524) );
  XNOR U5229 ( .A(n4523), .B(n4524), .Z(n4525) );
  XOR U5230 ( .A(n4526), .B(n4525), .Z(n4422) );
  OR U5231 ( .A(n4048), .B(n4047), .Z(n4052) );
  OR U5232 ( .A(n4050), .B(n4049), .Z(n4051) );
  AND U5233 ( .A(n4052), .B(n4051), .Z(n4547) );
  OR U5234 ( .A(n4058), .B(n4057), .Z(n4062) );
  OR U5235 ( .A(n4060), .B(n4059), .Z(n4061) );
  AND U5236 ( .A(n4062), .B(n4061), .Z(n4546) );
  XNOR U5237 ( .A(n4545), .B(n4546), .Z(n4548) );
  XNOR U5238 ( .A(n4547), .B(n4548), .Z(n4423) );
  XOR U5239 ( .A(n4422), .B(n4423), .Z(n4424) );
  XNOR U5240 ( .A(n4426), .B(n4427), .Z(n4429) );
  XNOR U5241 ( .A(n4429), .B(n4428), .Z(n4425) );
  XNOR U5242 ( .A(n4424), .B(n4425), .Z(n4468) );
  OR U5243 ( .A(n4088), .B(n4087), .Z(n4092) );
  OR U5244 ( .A(n4090), .B(n4089), .Z(n4091) );
  NAND U5245 ( .A(n4092), .B(n4091), .Z(n4433) );
  XNOR U5246 ( .A(n4432), .B(n4433), .Z(n4435) );
  OR U5247 ( .A(n4094), .B(n4093), .Z(n4098) );
  OR U5248 ( .A(n4096), .B(n4095), .Z(n4097) );
  NAND U5249 ( .A(n4098), .B(n4097), .Z(n4434) );
  XOR U5250 ( .A(n4435), .B(n4434), .Z(n4385) );
  XOR U5251 ( .A(n4385), .B(n4386), .Z(n4387) );
  XNOR U5252 ( .A(n4388), .B(n4387), .Z(n4466) );
  XOR U5253 ( .A(n4467), .B(n4466), .Z(n4469) );
  XOR U5254 ( .A(n4468), .B(n4469), .Z(n4454) );
  NANDN U5255 ( .A(n4104), .B(n4103), .Z(n4108) );
  NANDN U5256 ( .A(n4106), .B(n4105), .Z(n4107) );
  AND U5257 ( .A(n4108), .B(n4107), .Z(n4455) );
  NANDN U5258 ( .A(n4110), .B(n4109), .Z(n4114) );
  NANDN U5259 ( .A(n4112), .B(n4111), .Z(n4113) );
  NAND U5260 ( .A(n4114), .B(n4113), .Z(n4302) );
  XNOR U5261 ( .A(n4476), .B(n4477), .Z(n4479) );
  XNOR U5262 ( .A(n4479), .B(n4478), .Z(n4301) );
  XOR U5263 ( .A(n4302), .B(n4301), .Z(n4303) );
  XNOR U5264 ( .A(n4304), .B(n4303), .Z(n4297) );
  OR U5265 ( .A(n4139), .B(n4138), .Z(n4143) );
  OR U5266 ( .A(n4141), .B(n4140), .Z(n4142) );
  AND U5267 ( .A(n4143), .B(n4142), .Z(n4492) );
  XOR U5268 ( .A(n4332), .B(n4331), .Z(n4334) );
  NANDN U5269 ( .A(n4153), .B(n4152), .Z(n4157) );
  NAND U5270 ( .A(n4155), .B(n4154), .Z(n4156) );
  AND U5271 ( .A(n4157), .B(n4156), .Z(n4333) );
  XOR U5272 ( .A(n4334), .B(n4333), .Z(n4353) );
  XNOR U5273 ( .A(n4353), .B(n4354), .Z(n4356) );
  XNOR U5274 ( .A(n4356), .B(n4355), .Z(n4519) );
  OR U5275 ( .A(n4167), .B(n4166), .Z(n4171) );
  OR U5276 ( .A(n4169), .B(n4168), .Z(n4170) );
  AND U5277 ( .A(n4171), .B(n4170), .Z(n4517) );
  OR U5278 ( .A(n4173), .B(n4172), .Z(n4177) );
  OR U5279 ( .A(n4175), .B(n4174), .Z(n4176) );
  AND U5280 ( .A(n4177), .B(n4176), .Z(n4375) );
  OR U5281 ( .A(n4183), .B(n4182), .Z(n4187) );
  OR U5282 ( .A(n4185), .B(n4184), .Z(n4186) );
  NAND U5283 ( .A(n4187), .B(n4186), .Z(n4320) );
  XNOR U5284 ( .A(n4320), .B(n4319), .Z(n4321) );
  XNOR U5285 ( .A(n4322), .B(n4321), .Z(n4376) );
  XOR U5286 ( .A(n4375), .B(n4376), .Z(n4378) );
  OR U5287 ( .A(n4196), .B(oglobal[2]), .Z(n4200) );
  OR U5288 ( .A(n4198), .B(n4197), .Z(n4199) );
  NAND U5289 ( .A(n4200), .B(n4199), .Z(n4340) );
  OR U5290 ( .A(n4202), .B(n4201), .Z(n4206) );
  OR U5291 ( .A(n4204), .B(n4203), .Z(n4205) );
  NAND U5292 ( .A(n4206), .B(n4205), .Z(n4339) );
  XOR U5293 ( .A(n4340), .B(n4339), .Z(n4341) );
  XNOR U5294 ( .A(n4342), .B(n4341), .Z(n4377) );
  XNOR U5295 ( .A(n4378), .B(n4377), .Z(n4518) );
  XOR U5296 ( .A(n4517), .B(n4518), .Z(n4520) );
  XOR U5297 ( .A(n4519), .B(n4520), .Z(n4493) );
  XNOR U5298 ( .A(n4492), .B(n4493), .Z(n4495) );
  XNOR U5299 ( .A(n4494), .B(n4495), .Z(n4473) );
  NANDN U5300 ( .A(n4208), .B(n4207), .Z(n4212) );
  NANDN U5301 ( .A(n4210), .B(n4209), .Z(n4211) );
  AND U5302 ( .A(n4212), .B(n4211), .Z(n4471) );
  NANDN U5303 ( .A(n4214), .B(n4213), .Z(n4218) );
  NAND U5304 ( .A(n4216), .B(n4215), .Z(n4217) );
  NAND U5305 ( .A(n4218), .B(n4217), .Z(n4407) );
  XNOR U5306 ( .A(oglobal[3]), .B(n4407), .Z(n4409) );
  XOR U5307 ( .A(n4409), .B(n4408), .Z(n4371) );
  XNOR U5308 ( .A(n4402), .B(n4401), .Z(n4403) );
  XNOR U5309 ( .A(n4404), .B(n4403), .Z(n4369) );
  OR U5310 ( .A(n4236), .B(n4235), .Z(n4240) );
  NANDN U5311 ( .A(n4238), .B(n4237), .Z(n4239) );
  AND U5312 ( .A(n4240), .B(n4239), .Z(n4370) );
  XOR U5313 ( .A(n4369), .B(n4370), .Z(n4372) );
  XNOR U5314 ( .A(n4371), .B(n4372), .Z(n4392) );
  OR U5315 ( .A(n4254), .B(n4253), .Z(n4258) );
  OR U5316 ( .A(n4256), .B(n4255), .Z(n4257) );
  NAND U5317 ( .A(n4258), .B(n4257), .Z(n4350) );
  OR U5318 ( .A(n4260), .B(n4259), .Z(n4264) );
  OR U5319 ( .A(n4262), .B(n4261), .Z(n4263) );
  NAND U5320 ( .A(n4264), .B(n4263), .Z(n4348) );
  OR U5321 ( .A(n4266), .B(n4265), .Z(n4270) );
  OR U5322 ( .A(n4268), .B(n4267), .Z(n4269) );
  NAND U5323 ( .A(n4270), .B(n4269), .Z(n4347) );
  XNOR U5324 ( .A(n4348), .B(n4347), .Z(n4349) );
  XNOR U5325 ( .A(n4350), .B(n4349), .Z(n4510) );
  XOR U5326 ( .A(n4512), .B(n4510), .Z(n4513) );
  XNOR U5327 ( .A(n4514), .B(n4513), .Z(n4389) );
  XNOR U5328 ( .A(n4390), .B(n4389), .Z(n4391) );
  XOR U5329 ( .A(n4392), .B(n4391), .Z(n4484) );
  OR U5330 ( .A(n4272), .B(n4271), .Z(n4276) );
  OR U5331 ( .A(n4274), .B(n4273), .Z(n4275) );
  AND U5332 ( .A(n4276), .B(n4275), .Z(n4482) );
  XNOR U5333 ( .A(n4438), .B(n4439), .Z(n4441) );
  OR U5334 ( .A(n4286), .B(n4285), .Z(n4290) );
  OR U5335 ( .A(n4288), .B(n4287), .Z(n4289) );
  NAND U5336 ( .A(n4290), .B(n4289), .Z(n4440) );
  XOR U5337 ( .A(n4441), .B(n4440), .Z(n4483) );
  XNOR U5338 ( .A(n4482), .B(n4483), .Z(n4485) );
  XOR U5339 ( .A(n4484), .B(n4485), .Z(n4470) );
  XOR U5340 ( .A(n4471), .B(n4470), .Z(n4472) );
  XOR U5341 ( .A(n4473), .B(n4472), .Z(n4305) );
  XOR U5342 ( .A(n4305), .B(n4306), .Z(n4307) );
  XNOR U5343 ( .A(n4308), .B(n4307), .Z(n4295) );
  XOR U5344 ( .A(n4296), .B(n4295), .Z(n4298) );
  XNOR U5345 ( .A(n4297), .B(n4298), .Z(o[3]) );
  NANDN U5346 ( .A(n4296), .B(n4295), .Z(n4300) );
  NANDN U5347 ( .A(n4298), .B(n4297), .Z(n4299) );
  NAND U5348 ( .A(n4300), .B(n4299), .Z(n4553) );
  OR U5349 ( .A(n4314), .B(n4313), .Z(n4318) );
  OR U5350 ( .A(n4316), .B(n4315), .Z(n4317) );
  NAND U5351 ( .A(n4318), .B(n4317), .Z(n4629) );
  OR U5352 ( .A(n4320), .B(n4319), .Z(n4324) );
  OR U5353 ( .A(n4322), .B(n4321), .Z(n4323) );
  AND U5354 ( .A(n4324), .B(n4323), .Z(n4627) );
  NANDN U5355 ( .A(n4326), .B(n4325), .Z(n4330) );
  NAND U5356 ( .A(n4328), .B(n4327), .Z(n4329) );
  NAND U5357 ( .A(n4330), .B(n4329), .Z(n4628) );
  XOR U5358 ( .A(n4627), .B(n4628), .Z(n4630) );
  XOR U5359 ( .A(n4629), .B(n4630), .Z(n4626) );
  XOR U5360 ( .A(n4624), .B(n4623), .Z(n4625) );
  XOR U5361 ( .A(n4626), .B(n4625), .Z(n4645) );
  XNOR U5362 ( .A(n4644), .B(n4645), .Z(n4647) );
  OR U5363 ( .A(n4348), .B(n4347), .Z(n4352) );
  OR U5364 ( .A(n4350), .B(n4349), .Z(n4351) );
  NAND U5365 ( .A(n4352), .B(n4351), .Z(n4617) );
  XNOR U5366 ( .A(n4618), .B(n4617), .Z(n4619) );
  XNOR U5367 ( .A(n4620), .B(n4619), .Z(n4646) );
  XNOR U5368 ( .A(n4647), .B(n4646), .Z(n4599) );
  OR U5369 ( .A(n4354), .B(n4353), .Z(n4358) );
  OR U5370 ( .A(n4356), .B(n4355), .Z(n4357) );
  NAND U5371 ( .A(n4358), .B(n4357), .Z(n4665) );
  OR U5372 ( .A(n4360), .B(n4359), .Z(n4364) );
  OR U5373 ( .A(n4362), .B(n4361), .Z(n4363) );
  AND U5374 ( .A(n4364), .B(n4363), .Z(n4662) );
  XNOR U5375 ( .A(n4662), .B(n4663), .Z(n4664) );
  XNOR U5376 ( .A(n4665), .B(n4664), .Z(n4652) );
  NANDN U5377 ( .A(n4370), .B(n4369), .Z(n4374) );
  OR U5378 ( .A(n4372), .B(n4371), .Z(n4373) );
  AND U5379 ( .A(n4374), .B(n4373), .Z(n4650) );
  XOR U5380 ( .A(n4650), .B(n4651), .Z(n4653) );
  XOR U5381 ( .A(n4652), .B(n4653), .Z(n4597) );
  NANDN U5382 ( .A(n4380), .B(n4379), .Z(n4384) );
  NANDN U5383 ( .A(n4382), .B(n4381), .Z(n4383) );
  AND U5384 ( .A(n4384), .B(n4383), .Z(n4598) );
  XOR U5385 ( .A(n4597), .B(n4598), .Z(n4600) );
  XOR U5386 ( .A(n4599), .B(n4600), .Z(n4587) );
  XNOR U5387 ( .A(n4587), .B(n4588), .Z(n4590) );
  NANDN U5388 ( .A(n4390), .B(n4389), .Z(n4394) );
  NAND U5389 ( .A(n4392), .B(n4391), .Z(n4393) );
  NAND U5390 ( .A(n4394), .B(n4393), .Z(n4596) );
  NANDN U5391 ( .A(n4396), .B(n4395), .Z(n4400) );
  NAND U5392 ( .A(n4398), .B(n4397), .Z(n4399) );
  AND U5393 ( .A(n4400), .B(n4399), .Z(n4657) );
  OR U5394 ( .A(n4402), .B(n4401), .Z(n4406) );
  OR U5395 ( .A(n4404), .B(n4403), .Z(n4405) );
  NAND U5396 ( .A(n4406), .B(n4405), .Z(n4632) );
  NANDN U5397 ( .A(n4407), .B(oglobal[3]), .Z(n4411) );
  NAND U5398 ( .A(n4409), .B(n4408), .Z(n4410) );
  NAND U5399 ( .A(n4411), .B(n4410), .Z(n4631) );
  XNOR U5400 ( .A(n4631), .B(oglobal[4]), .Z(n4633) );
  XNOR U5401 ( .A(n4632), .B(n4633), .Z(n4656) );
  XOR U5402 ( .A(n4657), .B(n4656), .Z(n4659) );
  OR U5403 ( .A(n4413), .B(n4412), .Z(n4417) );
  NANDN U5404 ( .A(n4415), .B(n4414), .Z(n4416) );
  NAND U5405 ( .A(n4417), .B(n4416), .Z(n4658) );
  XOR U5406 ( .A(n4659), .B(n4658), .Z(n4593) );
  XOR U5407 ( .A(n4593), .B(n4594), .Z(n4595) );
  XNOR U5408 ( .A(n4596), .B(n4595), .Z(n4589) );
  XNOR U5409 ( .A(n4590), .B(n4589), .Z(n4557) );
  OR U5410 ( .A(n4427), .B(n4426), .Z(n4431) );
  OR U5411 ( .A(n4429), .B(n4428), .Z(n4430) );
  AND U5412 ( .A(n4431), .B(n4430), .Z(n4606) );
  OR U5413 ( .A(n4433), .B(n4432), .Z(n4437) );
  OR U5414 ( .A(n4435), .B(n4434), .Z(n4436) );
  AND U5415 ( .A(n4437), .B(n4436), .Z(n4603) );
  OR U5416 ( .A(n4439), .B(n4438), .Z(n4443) );
  OR U5417 ( .A(n4441), .B(n4440), .Z(n4442) );
  AND U5418 ( .A(n4443), .B(n4442), .Z(n4604) );
  XOR U5419 ( .A(n4603), .B(n4604), .Z(n4605) );
  XNOR U5420 ( .A(n4606), .B(n4605), .Z(n4565) );
  XOR U5421 ( .A(n4566), .B(n4565), .Z(n4568) );
  XNOR U5422 ( .A(n4568), .B(n4567), .Z(n4556) );
  NAND U5423 ( .A(n4449), .B(n4448), .Z(n4453) );
  NAND U5424 ( .A(n4451), .B(n4450), .Z(n4452) );
  NAND U5425 ( .A(n4453), .B(n4452), .Z(n4555) );
  XNOR U5426 ( .A(n4556), .B(n4555), .Z(n4558) );
  XOR U5427 ( .A(n4557), .B(n4558), .Z(n4674) );
  XNOR U5428 ( .A(n4676), .B(n4677), .Z(n4552) );
  NANDN U5429 ( .A(n4455), .B(n4454), .Z(n4459) );
  NAND U5430 ( .A(n4457), .B(n4456), .Z(n4458) );
  NAND U5431 ( .A(n4459), .B(n4458), .Z(n4671) );
  NANDN U5432 ( .A(n4461), .B(n4460), .Z(n4465) );
  NANDN U5433 ( .A(n4463), .B(n4462), .Z(n4464) );
  NAND U5434 ( .A(n4465), .B(n4464), .Z(n4584) );
  NANDN U5435 ( .A(n4471), .B(n4470), .Z(n4475) );
  OR U5436 ( .A(n4473), .B(n4472), .Z(n4474) );
  AND U5437 ( .A(n4475), .B(n4474), .Z(n4582) );
  XOR U5438 ( .A(n4581), .B(n4582), .Z(n4583) );
  XNOR U5439 ( .A(n4584), .B(n4583), .Z(n4669) );
  OR U5440 ( .A(n4477), .B(n4476), .Z(n4481) );
  OR U5441 ( .A(n4479), .B(n4478), .Z(n4480) );
  NAND U5442 ( .A(n4481), .B(n4480), .Z(n4562) );
  OR U5443 ( .A(n4487), .B(n4486), .Z(n4491) );
  OR U5444 ( .A(n4489), .B(n4488), .Z(n4490) );
  AND U5445 ( .A(n4491), .B(n4490), .Z(n4575) );
  OR U5446 ( .A(n4493), .B(n4492), .Z(n4497) );
  OR U5447 ( .A(n4495), .B(n4494), .Z(n4496) );
  AND U5448 ( .A(n4497), .B(n4496), .Z(n4576) );
  XNOR U5449 ( .A(n4575), .B(n4576), .Z(n4578) );
  XNOR U5450 ( .A(n4577), .B(n4578), .Z(n4560) );
  IV U5451 ( .A(n4510), .Z(n4511) );
  NANDN U5452 ( .A(n4512), .B(n4511), .Z(n4516) );
  NANDN U5453 ( .A(n4514), .B(n4513), .Z(n4515) );
  NAND U5454 ( .A(n4516), .B(n4515), .Z(n4614) );
  XOR U5455 ( .A(n4613), .B(n4614), .Z(n4616) );
  XOR U5456 ( .A(n4615), .B(n4616), .Z(n4607) );
  OR U5457 ( .A(n4518), .B(n4517), .Z(n4522) );
  NAND U5458 ( .A(n4520), .B(n4519), .Z(n4521) );
  AND U5459 ( .A(n4522), .B(n4521), .Z(n4608) );
  XNOR U5460 ( .A(n4607), .B(n4608), .Z(n4609) );
  XOR U5461 ( .A(n4610), .B(n4609), .Z(n4573) );
  OR U5462 ( .A(n4528), .B(n4527), .Z(n4532) );
  NAND U5463 ( .A(n4530), .B(n4529), .Z(n4531) );
  NAND U5464 ( .A(n4532), .B(n4531), .Z(n4637) );
  XOR U5465 ( .A(n4640), .B(n4641), .Z(n4642) );
  XNOR U5466 ( .A(n4643), .B(n4642), .Z(n4636) );
  XOR U5467 ( .A(n4637), .B(n4636), .Z(n4639) );
  XOR U5468 ( .A(n4638), .B(n4639), .Z(n4571) );
  OR U5469 ( .A(n4546), .B(n4545), .Z(n4550) );
  OR U5470 ( .A(n4548), .B(n4547), .Z(n4549) );
  NAND U5471 ( .A(n4550), .B(n4549), .Z(n4572) );
  XOR U5472 ( .A(n4571), .B(n4572), .Z(n4574) );
  XOR U5473 ( .A(n4573), .B(n4574), .Z(n4559) );
  XOR U5474 ( .A(n4560), .B(n4559), .Z(n4561) );
  XNOR U5475 ( .A(n4562), .B(n4561), .Z(n4668) );
  XOR U5476 ( .A(n4669), .B(n4668), .Z(n4670) );
  XOR U5477 ( .A(n4671), .B(n4670), .Z(n4554) );
  XOR U5478 ( .A(n4552), .B(n4554), .Z(n4551) );
  XNOR U5479 ( .A(n4553), .B(n4551), .Z(o[4]) );
  NANDN U5480 ( .A(n4560), .B(n4559), .Z(n4564) );
  OR U5481 ( .A(n4562), .B(n4561), .Z(n4563) );
  NAND U5482 ( .A(n4564), .B(n4563), .Z(n4730) );
  NANDN U5483 ( .A(n4566), .B(n4565), .Z(n4570) );
  OR U5484 ( .A(n4568), .B(n4567), .Z(n4569) );
  AND U5485 ( .A(n4570), .B(n4569), .Z(n4686) );
  XNOR U5486 ( .A(n4686), .B(n4687), .Z(n4689) );
  OR U5487 ( .A(n4576), .B(n4575), .Z(n4580) );
  OR U5488 ( .A(n4578), .B(n4577), .Z(n4579) );
  NAND U5489 ( .A(n4580), .B(n4579), .Z(n4688) );
  XNOR U5490 ( .A(n4689), .B(n4688), .Z(n4729) );
  XOR U5491 ( .A(n4730), .B(n4729), .Z(n4731) );
  XOR U5492 ( .A(n4732), .B(n4731), .Z(n4680) );
  XOR U5493 ( .A(n4681), .B(n4680), .Z(n4682) );
  OR U5494 ( .A(n4582), .B(n4581), .Z(n4586) );
  NANDN U5495 ( .A(n4584), .B(n4583), .Z(n4585) );
  AND U5496 ( .A(n4586), .B(n4585), .Z(n4725) );
  OR U5497 ( .A(n4588), .B(n4587), .Z(n4592) );
  NANDN U5498 ( .A(n4590), .B(n4589), .Z(n4591) );
  AND U5499 ( .A(n4592), .B(n4591), .Z(n4724) );
  OR U5500 ( .A(n4598), .B(n4597), .Z(n4602) );
  NAND U5501 ( .A(n4600), .B(n4599), .Z(n4601) );
  AND U5502 ( .A(n4602), .B(n4601), .Z(n4713) );
  XNOR U5503 ( .A(n4713), .B(n4714), .Z(n4715) );
  XOR U5504 ( .A(n4716), .B(n4715), .Z(n4722) );
  OR U5505 ( .A(n4608), .B(n4607), .Z(n4612) );
  OR U5506 ( .A(n4610), .B(n4609), .Z(n4611) );
  NAND U5507 ( .A(n4612), .B(n4611), .Z(n4720) );
  OR U5508 ( .A(n4618), .B(n4617), .Z(n4622) );
  OR U5509 ( .A(n4620), .B(n4619), .Z(n4621) );
  AND U5510 ( .A(n4622), .B(n4621), .Z(n4704) );
  XNOR U5511 ( .A(n4701), .B(n4702), .Z(n4703) );
  XOR U5512 ( .A(n4704), .B(n4703), .Z(n4705) );
  NAND U5513 ( .A(n4631), .B(oglobal[4]), .Z(n4635) );
  NANDN U5514 ( .A(n4633), .B(n4632), .Z(n4634) );
  AND U5515 ( .A(n4635), .B(n4634), .Z(n4700) );
  XOR U5516 ( .A(n4700), .B(oglobal[5]), .Z(n4706) );
  XOR U5517 ( .A(n4705), .B(n4706), .Z(n4707) );
  XNOR U5518 ( .A(n4708), .B(n4707), .Z(n4709) );
  XOR U5519 ( .A(n4709), .B(n4710), .Z(n4711) );
  OR U5520 ( .A(n4645), .B(n4644), .Z(n4649) );
  OR U5521 ( .A(n4647), .B(n4646), .Z(n4648) );
  AND U5522 ( .A(n4649), .B(n4648), .Z(n4697) );
  XOR U5523 ( .A(n4696), .B(n4697), .Z(n4699) );
  OR U5524 ( .A(n4651), .B(n4650), .Z(n4655) );
  NAND U5525 ( .A(n4653), .B(n4652), .Z(n4654) );
  AND U5526 ( .A(n4655), .B(n4654), .Z(n4698) );
  XOR U5527 ( .A(n4699), .B(n4698), .Z(n4694) );
  NANDN U5528 ( .A(n4657), .B(n4656), .Z(n4661) );
  OR U5529 ( .A(n4659), .B(n4658), .Z(n4660) );
  NAND U5530 ( .A(n4661), .B(n4660), .Z(n4693) );
  OR U5531 ( .A(n4663), .B(n4662), .Z(n4667) );
  OR U5532 ( .A(n4665), .B(n4664), .Z(n4666) );
  NAND U5533 ( .A(n4667), .B(n4666), .Z(n4692) );
  XOR U5534 ( .A(n4693), .B(n4692), .Z(n4695) );
  XOR U5535 ( .A(n4694), .B(n4695), .Z(n4712) );
  XOR U5536 ( .A(n4711), .B(n4712), .Z(n4719) );
  XOR U5537 ( .A(n4720), .B(n4719), .Z(n4721) );
  XNOR U5538 ( .A(n4722), .B(n4721), .Z(n4723) );
  XOR U5539 ( .A(n4724), .B(n4723), .Z(n4726) );
  XNOR U5540 ( .A(n4725), .B(n4726), .Z(n4734) );
  NANDN U5541 ( .A(n4669), .B(n4668), .Z(n4673) );
  OR U5542 ( .A(n4671), .B(n4670), .Z(n4672) );
  NAND U5543 ( .A(n4673), .B(n4672), .Z(n4733) );
  XOR U5544 ( .A(n4734), .B(n4733), .Z(n4735) );
  NANDN U5545 ( .A(n4675), .B(n4674), .Z(n4679) );
  OR U5546 ( .A(n4677), .B(n4676), .Z(n4678) );
  NAND U5547 ( .A(n4679), .B(n4678), .Z(n4736) );
  XNOR U5548 ( .A(n4735), .B(n4736), .Z(n4683) );
  XNOR U5549 ( .A(n4682), .B(n4683), .Z(o[5]) );
  OR U5550 ( .A(n4681), .B(n4680), .Z(n4685) );
  NANDN U5551 ( .A(n4683), .B(n4682), .Z(n4684) );
  NAND U5552 ( .A(n4685), .B(n4684), .Z(n4747) );
  OR U5553 ( .A(n4687), .B(n4686), .Z(n4691) );
  OR U5554 ( .A(n4689), .B(n4688), .Z(n4690) );
  AND U5555 ( .A(n4691), .B(n4690), .Z(n4751) );
  ANDN U5556 ( .B(oglobal[5]), .A(n4700), .Z(n4759) );
  XOR U5557 ( .A(oglobal[6]), .B(n4759), .Z(n4760) );
  XNOR U5558 ( .A(n4760), .B(n4761), .Z(n4762) );
  XNOR U5559 ( .A(n4762), .B(n4763), .Z(n4767) );
  XOR U5560 ( .A(n4766), .B(n4767), .Z(n4768) );
  XNOR U5561 ( .A(n4769), .B(n4768), .Z(n4756) );
  OR U5562 ( .A(n4714), .B(n4713), .Z(n4718) );
  OR U5563 ( .A(n4716), .B(n4715), .Z(n4717) );
  NAND U5564 ( .A(n4718), .B(n4717), .Z(n4754) );
  XNOR U5565 ( .A(n4753), .B(n4754), .Z(n4755) );
  XOR U5566 ( .A(n4756), .B(n4755), .Z(n4749) );
  XNOR U5567 ( .A(n4749), .B(n4750), .Z(n4752) );
  XOR U5568 ( .A(n4751), .B(n4752), .Z(n4740) );
  NANDN U5569 ( .A(n4724), .B(n4723), .Z(n4728) );
  OR U5570 ( .A(n4726), .B(n4725), .Z(n4727) );
  NAND U5571 ( .A(n4728), .B(n4727), .Z(n4741) );
  XNOR U5572 ( .A(n4743), .B(n4742), .Z(n4746) );
  OR U5573 ( .A(n4734), .B(n4733), .Z(n4738) );
  NANDN U5574 ( .A(n4736), .B(n4735), .Z(n4737) );
  NAND U5575 ( .A(n4738), .B(n4737), .Z(n4748) );
  XNOR U5576 ( .A(n4746), .B(n4748), .Z(n4739) );
  XNOR U5577 ( .A(n4747), .B(n4739), .Z(o[6]) );
  NANDN U5578 ( .A(n4741), .B(n4740), .Z(n4745) );
  OR U5579 ( .A(n4743), .B(n4742), .Z(n4744) );
  AND U5580 ( .A(n4745), .B(n4744), .Z(n4773) );
  NANDN U5581 ( .A(n4754), .B(n4753), .Z(n4758) );
  NAND U5582 ( .A(n4756), .B(n4755), .Z(n4757) );
  AND U5583 ( .A(n4758), .B(n4757), .Z(n4774) );
  NAND U5584 ( .A(n4759), .B(oglobal[6]), .Z(n4784) );
  XOR U5585 ( .A(oglobal[7]), .B(n4784), .Z(n4779) );
  NANDN U5586 ( .A(n4761), .B(n4760), .Z(n4765) );
  NANDN U5587 ( .A(n4763), .B(n4762), .Z(n4764) );
  AND U5588 ( .A(n4765), .B(n4764), .Z(n4778) );
  XNOR U5589 ( .A(n4779), .B(n4778), .Z(n4781) );
  XOR U5590 ( .A(n4781), .B(n4780), .Z(n4775) );
  XOR U5591 ( .A(n4774), .B(n4775), .Z(n4776) );
  XOR U5592 ( .A(n4777), .B(n4776), .Z(n4772) );
  XOR U5593 ( .A(n4771), .B(n4772), .Z(n4770) );
  XOR U5594 ( .A(n4773), .B(n4770), .Z(o[7]) );
  XNOR U5595 ( .A(n4786), .B(n4785), .Z(n4787) );
  OR U5596 ( .A(n4779), .B(n4778), .Z(n4783) );
  OR U5597 ( .A(n4781), .B(n4780), .Z(n4782) );
  AND U5598 ( .A(n4783), .B(n4782), .Z(n4792) );
  NANDN U5599 ( .A(n4784), .B(oglobal[7]), .Z(n4791) );
  XOR U5600 ( .A(oglobal[8]), .B(n4791), .Z(n4793) );
  XNOR U5601 ( .A(n4792), .B(n4793), .Z(n4788) );
  XNOR U5602 ( .A(n4787), .B(n4788), .Z(o[8]) );
  NANDN U5603 ( .A(n4786), .B(n4785), .Z(n4790) );
  NANDN U5604 ( .A(n4788), .B(n4787), .Z(n4789) );
  NAND U5605 ( .A(n4790), .B(n4789), .Z(n4796) );
  XNOR U5606 ( .A(n4796), .B(oglobal[9]), .Z(n4798) );
  NANDN U5607 ( .A(n4791), .B(oglobal[8]), .Z(n4795) );
  OR U5608 ( .A(n4793), .B(n4792), .Z(n4794) );
  AND U5609 ( .A(n4795), .B(n4794), .Z(n4797) );
  XOR U5610 ( .A(n4798), .B(n4797), .Z(o[9]) );
  AND U5611 ( .A(oglobal[9]), .B(n4796), .Z(n4800) );
  NOR U5612 ( .A(n4798), .B(n4797), .Z(n4799) );
  NOR U5613 ( .A(n4800), .B(n4799), .Z(n4801) );
  XNOR U5614 ( .A(oglobal[10]), .B(n4801), .Z(o[10]) );
endmodule

